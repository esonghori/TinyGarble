
module FA_2048 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  AND U1 ( .A(A), .B(B), .Z(CO) );
  XOR U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_3071 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3070 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3069 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3068 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3067 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3066 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3065 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3064 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3063 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3062 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3061 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3060 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3059 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3058 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3057 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3056 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3055 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3054 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3053 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3052 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3051 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3050 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3049 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3048 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3047 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3046 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3045 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3044 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3043 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3042 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3041 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3040 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3039 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3038 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3037 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3036 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3035 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3034 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3033 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3032 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3031 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3030 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3029 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3028 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3027 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3026 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3025 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3024 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3023 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3022 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3021 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3020 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3019 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3018 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3017 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3016 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3015 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3014 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3013 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3012 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3011 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3010 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3009 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3008 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3007 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3006 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3005 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3004 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3003 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3002 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3001 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_3000 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2999 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2998 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2997 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2996 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2995 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2994 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2993 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2992 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2991 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2990 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2989 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2988 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2987 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2986 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2985 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2984 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2983 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2982 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2981 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2980 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2979 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2978 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2977 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2976 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2975 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2974 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2973 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2972 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2971 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2970 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2969 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2968 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2967 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2966 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2965 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2964 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2963 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2962 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2961 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2960 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2959 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2958 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2957 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2956 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2955 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2954 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2953 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2952 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2951 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2950 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2949 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2948 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2947 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2946 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2945 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2944 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2943 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2942 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2941 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2940 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2939 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2938 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2937 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2936 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2935 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2934 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2933 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2932 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2931 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2930 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2929 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2928 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2927 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2926 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2925 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2924 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2923 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2922 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2921 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2920 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2919 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2918 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2917 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2916 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2915 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2914 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2913 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2912 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2911 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2910 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2909 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2908 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2907 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2906 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2905 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2904 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2903 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2902 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2901 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2900 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2899 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2898 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2897 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2896 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2895 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2894 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2893 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2892 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2891 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2890 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2889 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2888 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2887 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2886 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2885 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2884 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2883 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2882 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2881 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2880 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2879 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2878 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2877 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2876 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2875 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2874 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2873 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2872 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2871 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2870 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2869 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2868 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2867 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2866 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2865 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2864 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2863 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2862 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2861 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2860 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2859 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2858 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2857 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2856 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2855 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2854 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2853 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2852 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2851 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2850 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2849 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2848 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2847 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2846 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2845 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2844 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2843 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2842 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2841 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2840 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2839 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2838 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2837 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2836 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2835 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2834 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2833 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2832 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2831 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2830 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2829 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2828 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2827 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2826 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2825 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2824 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2823 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2822 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2821 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2820 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2819 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2818 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2817 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2816 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2815 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2814 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2813 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2812 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2811 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2810 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2809 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2808 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2807 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2806 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2805 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2804 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2803 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2802 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2801 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2800 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2799 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2798 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2797 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2796 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2795 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2794 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2793 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2792 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2791 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2790 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2789 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2788 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2787 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2786 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2785 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2784 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2783 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2782 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2781 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2780 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2779 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2778 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2777 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2776 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2775 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2774 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2773 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2772 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2771 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2770 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2769 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2768 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2767 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2766 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2765 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2764 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2763 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2762 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2761 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2760 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2759 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2758 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2757 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2756 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2755 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2754 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2753 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2752 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2751 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2750 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2749 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2748 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2747 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2746 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2745 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2744 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2743 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2742 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2741 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2740 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2739 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2738 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2737 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2736 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2735 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2734 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2733 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2732 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2731 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2730 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2729 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2728 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2727 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2726 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2725 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2724 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2723 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2722 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2721 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2720 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2719 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2718 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2717 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2716 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2715 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2714 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2713 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2712 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2711 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2710 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2709 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2708 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2707 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2706 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2705 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2704 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2703 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2702 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2701 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2700 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2699 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2698 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2697 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2696 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2695 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2694 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2693 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2692 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2691 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2690 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2689 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2688 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2687 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2686 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2685 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2684 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2683 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2682 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2681 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2680 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2679 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2678 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2677 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2676 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2675 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2674 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2673 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2672 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2671 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2670 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2669 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2668 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2667 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2666 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2665 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2664 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2663 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2662 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2661 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2660 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2659 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2658 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2657 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2656 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2655 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2654 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2653 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2652 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2651 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2650 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2649 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2648 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2647 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2646 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2645 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2644 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2643 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2642 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2641 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2640 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2639 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2638 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2637 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2636 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2635 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2634 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2633 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2632 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2631 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2630 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2629 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2628 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2627 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2626 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2625 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2624 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2623 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2622 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2621 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2620 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2619 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2618 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2617 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2616 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2615 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2614 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2613 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2612 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2611 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2610 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2609 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2608 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2607 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2606 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2605 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2604 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2603 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2602 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2601 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2600 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2599 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2598 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2597 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2596 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2595 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2594 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2593 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2592 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2591 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2590 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2589 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2588 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2587 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2586 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2585 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2584 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2583 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2582 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2581 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2580 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2579 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2578 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2577 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2576 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2575 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2574 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2573 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2572 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2571 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2570 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2569 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2568 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2567 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2566 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2565 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2564 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2563 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2562 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2561 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2560 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2559 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2558 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2557 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2556 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2555 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2554 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2553 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2552 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2551 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2550 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2549 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2548 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2547 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2546 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2545 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2544 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2543 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2542 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2541 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2540 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2539 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2538 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2537 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2536 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2535 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2534 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2533 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2532 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2531 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2530 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2529 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2528 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2527 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2526 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2525 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2524 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2523 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2522 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2521 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2520 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2519 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2518 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2517 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2516 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2515 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2514 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2513 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2512 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2511 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2510 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2509 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2508 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2507 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2506 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2505 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2504 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2503 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2502 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2501 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2500 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2499 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2498 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2497 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2496 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2495 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2494 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2493 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2492 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2491 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2490 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2489 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2488 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2487 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2486 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2485 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2484 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2483 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2482 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2481 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2480 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2479 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2478 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2477 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2476 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2475 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2474 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2473 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2472 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2471 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2470 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2469 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2468 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2467 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2466 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2465 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2464 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2463 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2462 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2461 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2460 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2459 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2458 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2457 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2456 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2455 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2454 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2453 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2452 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2451 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2450 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2449 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2448 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2447 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2446 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2445 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2444 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2443 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2442 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2441 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2440 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2439 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2438 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2437 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2436 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2435 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2434 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2433 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2432 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2431 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2430 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2429 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2428 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2427 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2426 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2425 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2424 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2423 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2422 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2421 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2420 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2419 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2418 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2417 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2416 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2415 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2414 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2413 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2412 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2411 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2410 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2409 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2408 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2407 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2406 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2405 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2404 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2403 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2402 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2401 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2400 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2399 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2398 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2397 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2396 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2395 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2394 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2393 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2392 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2391 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2390 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2389 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2388 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2387 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2386 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2385 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2384 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2383 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2382 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2381 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2380 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2379 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2378 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2377 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2376 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2375 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2374 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2373 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2372 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2371 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2370 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2369 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2368 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2367 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2366 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2365 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2364 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2363 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2362 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2361 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2360 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2359 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2358 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2357 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2356 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2355 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2354 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2353 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2352 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2351 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2350 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2349 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2348 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2347 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2346 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2345 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2344 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2343 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2342 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2341 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2340 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2339 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2338 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2337 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2336 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2335 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2334 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2333 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2332 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2331 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2330 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2329 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2328 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2327 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2326 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2325 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2324 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2323 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2322 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2321 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2320 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2319 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2318 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2317 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2316 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2315 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2314 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2313 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2312 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2311 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2310 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2309 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2308 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2307 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2306 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2305 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2304 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2303 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2302 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2301 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2300 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2299 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2298 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2297 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2296 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2295 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2294 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2293 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2292 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2291 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2290 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2289 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2288 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2287 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2286 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2285 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2284 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2283 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2282 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2281 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2280 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2279 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2278 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2277 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2276 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2275 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2274 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2273 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2272 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2271 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2270 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2269 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2268 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2267 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2266 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2265 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2264 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2263 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2262 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2261 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2260 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2259 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2258 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2257 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2256 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2255 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2254 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2253 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2252 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2251 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2250 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2249 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2248 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2247 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2246 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2245 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2244 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2243 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2242 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2241 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2240 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2239 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2238 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2237 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2236 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2235 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2234 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2233 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2232 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2231 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2230 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2229 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2228 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2227 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2226 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2225 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2224 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2223 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2222 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2221 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2220 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2219 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2218 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2217 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2216 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2215 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2214 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2213 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2212 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2211 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2210 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2209 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2208 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2207 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2206 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2205 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2204 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2203 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2202 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2201 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2200 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2199 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2198 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2197 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2196 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2195 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2194 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2193 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2192 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2191 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2190 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2189 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2188 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2187 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2186 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2185 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2184 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2183 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2182 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2181 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2180 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2179 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2178 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2177 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2176 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2175 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2174 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2173 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2172 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2171 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2170 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2169 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2168 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2167 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2166 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2165 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2164 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2163 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2162 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2161 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2160 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2159 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2158 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2157 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2156 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2155 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2154 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2153 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2152 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2151 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2150 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2149 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2148 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2147 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2146 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2145 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2144 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2143 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2142 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2141 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2140 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2139 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2138 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2137 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2136 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2135 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2134 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2133 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2132 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2131 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2130 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2129 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2128 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2127 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2126 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2125 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2124 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2123 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2122 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2121 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2120 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2119 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2118 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2117 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2116 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2115 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2114 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2113 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2112 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2111 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2110 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2109 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2108 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2107 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2106 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2105 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2104 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2103 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2102 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2101 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2100 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2099 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2098 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2097 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2096 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2095 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2094 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2093 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2092 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2091 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2090 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2089 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2088 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2087 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2086 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2085 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2084 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2083 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2082 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2081 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2080 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2079 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2078 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2077 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2076 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2075 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2074 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2073 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2072 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2071 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2070 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2069 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2068 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2067 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2066 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2065 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2064 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2063 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2062 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2061 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2060 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2059 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2058 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2057 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2056 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2055 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2054 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2053 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_2052 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(CI), .B(n1), .Z(S) );
  ANDN U2 ( .B(CI), .A(n1), .Z(CO) );
  XOR U3 ( .A(B), .B(CI), .Z(n1) );
endmodule


module FA_2051 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(CI), .B(n1), .Z(S) );
  ANDN U2 ( .B(CI), .A(n1), .Z(CO) );
  XOR U3 ( .A(B), .B(CI), .Z(n1) );
endmodule


module FA_2050 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(CI), .B(n1), .Z(S) );
  XOR U2 ( .A(B), .B(CI), .Z(n1) );
endmodule


module FA_2049 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N1024_2 ( A, B, CI, S, CO );
  input [1023:0] A;
  input [1023:0] B;
  output [1023:0] S;
  input CI;
  output CO;

  wire   [1023:1] C;

  FA_2048 \FA_INST_0[0].FA_INST_1[0].FA_  ( .A(A[0]), .B(B[0]), .CI(1'b0), .S(
        S[0]), .CO(C[1]) );
  FA_3071 \FA_INST_0[0].FA_INST_1[1].FA_  ( .A(A[1]), .B(B[1]), .CI(C[1]), .S(
        S[1]), .CO(C[2]) );
  FA_3070 \FA_INST_0[0].FA_INST_1[2].FA_  ( .A(A[2]), .B(B[2]), .CI(C[2]), .S(
        S[2]), .CO(C[3]) );
  FA_3069 \FA_INST_0[0].FA_INST_1[3].FA_  ( .A(A[3]), .B(B[3]), .CI(C[3]), .S(
        S[3]), .CO(C[4]) );
  FA_3068 \FA_INST_0[0].FA_INST_1[4].FA_  ( .A(A[4]), .B(B[4]), .CI(C[4]), .S(
        S[4]), .CO(C[5]) );
  FA_3067 \FA_INST_0[0].FA_INST_1[5].FA_  ( .A(A[5]), .B(B[5]), .CI(C[5]), .S(
        S[5]), .CO(C[6]) );
  FA_3066 \FA_INST_0[0].FA_INST_1[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(
        S[6]), .CO(C[7]) );
  FA_3065 \FA_INST_0[0].FA_INST_1[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(
        S[7]), .CO(C[8]) );
  FA_3064 \FA_INST_0[0].FA_INST_1[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(
        S[8]), .CO(C[9]) );
  FA_3063 \FA_INST_0[0].FA_INST_1[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(
        S[9]), .CO(C[10]) );
  FA_3062 \FA_INST_0[0].FA_INST_1[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), 
        .S(S[10]), .CO(C[11]) );
  FA_3061 \FA_INST_0[0].FA_INST_1[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), 
        .S(S[11]), .CO(C[12]) );
  FA_3060 \FA_INST_0[0].FA_INST_1[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), 
        .S(S[12]), .CO(C[13]) );
  FA_3059 \FA_INST_0[0].FA_INST_1[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), 
        .S(S[13]), .CO(C[14]) );
  FA_3058 \FA_INST_0[0].FA_INST_1[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), 
        .S(S[14]), .CO(C[15]) );
  FA_3057 \FA_INST_0[0].FA_INST_1[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), 
        .S(S[15]), .CO(C[16]) );
  FA_3056 \FA_INST_0[0].FA_INST_1[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), 
        .S(S[16]), .CO(C[17]) );
  FA_3055 \FA_INST_0[0].FA_INST_1[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), 
        .S(S[17]), .CO(C[18]) );
  FA_3054 \FA_INST_0[0].FA_INST_1[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), 
        .S(S[18]), .CO(C[19]) );
  FA_3053 \FA_INST_0[0].FA_INST_1[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), 
        .S(S[19]), .CO(C[20]) );
  FA_3052 \FA_INST_0[0].FA_INST_1[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), 
        .S(S[20]), .CO(C[21]) );
  FA_3051 \FA_INST_0[0].FA_INST_1[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), 
        .S(S[21]), .CO(C[22]) );
  FA_3050 \FA_INST_0[0].FA_INST_1[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), 
        .S(S[22]), .CO(C[23]) );
  FA_3049 \FA_INST_0[0].FA_INST_1[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), 
        .S(S[23]), .CO(C[24]) );
  FA_3048 \FA_INST_0[0].FA_INST_1[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), 
        .S(S[24]), .CO(C[25]) );
  FA_3047 \FA_INST_0[0].FA_INST_1[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), 
        .S(S[25]), .CO(C[26]) );
  FA_3046 \FA_INST_0[0].FA_INST_1[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), 
        .S(S[26]), .CO(C[27]) );
  FA_3045 \FA_INST_0[0].FA_INST_1[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), 
        .S(S[27]), .CO(C[28]) );
  FA_3044 \FA_INST_0[0].FA_INST_1[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), 
        .S(S[28]), .CO(C[29]) );
  FA_3043 \FA_INST_0[0].FA_INST_1[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), 
        .S(S[29]), .CO(C[30]) );
  FA_3042 \FA_INST_0[0].FA_INST_1[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), 
        .S(S[30]), .CO(C[31]) );
  FA_3041 \FA_INST_0[0].FA_INST_1[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), 
        .S(S[31]), .CO(C[32]) );
  FA_3040 \FA_INST_0[0].FA_INST_1[32].FA_  ( .A(A[32]), .B(B[32]), .CI(C[32]), 
        .S(S[32]), .CO(C[33]) );
  FA_3039 \FA_INST_0[0].FA_INST_1[33].FA_  ( .A(A[33]), .B(B[33]), .CI(C[33]), 
        .S(S[33]), .CO(C[34]) );
  FA_3038 \FA_INST_0[0].FA_INST_1[34].FA_  ( .A(A[34]), .B(B[34]), .CI(C[34]), 
        .S(S[34]), .CO(C[35]) );
  FA_3037 \FA_INST_0[0].FA_INST_1[35].FA_  ( .A(A[35]), .B(B[35]), .CI(C[35]), 
        .S(S[35]), .CO(C[36]) );
  FA_3036 \FA_INST_0[0].FA_INST_1[36].FA_  ( .A(A[36]), .B(B[36]), .CI(C[36]), 
        .S(S[36]), .CO(C[37]) );
  FA_3035 \FA_INST_0[0].FA_INST_1[37].FA_  ( .A(A[37]), .B(B[37]), .CI(C[37]), 
        .S(S[37]), .CO(C[38]) );
  FA_3034 \FA_INST_0[0].FA_INST_1[38].FA_  ( .A(A[38]), .B(B[38]), .CI(C[38]), 
        .S(S[38]), .CO(C[39]) );
  FA_3033 \FA_INST_0[0].FA_INST_1[39].FA_  ( .A(A[39]), .B(B[39]), .CI(C[39]), 
        .S(S[39]), .CO(C[40]) );
  FA_3032 \FA_INST_0[0].FA_INST_1[40].FA_  ( .A(A[40]), .B(B[40]), .CI(C[40]), 
        .S(S[40]), .CO(C[41]) );
  FA_3031 \FA_INST_0[0].FA_INST_1[41].FA_  ( .A(A[41]), .B(B[41]), .CI(C[41]), 
        .S(S[41]), .CO(C[42]) );
  FA_3030 \FA_INST_0[0].FA_INST_1[42].FA_  ( .A(A[42]), .B(B[42]), .CI(C[42]), 
        .S(S[42]), .CO(C[43]) );
  FA_3029 \FA_INST_0[0].FA_INST_1[43].FA_  ( .A(A[43]), .B(B[43]), .CI(C[43]), 
        .S(S[43]), .CO(C[44]) );
  FA_3028 \FA_INST_0[0].FA_INST_1[44].FA_  ( .A(A[44]), .B(B[44]), .CI(C[44]), 
        .S(S[44]), .CO(C[45]) );
  FA_3027 \FA_INST_0[0].FA_INST_1[45].FA_  ( .A(A[45]), .B(B[45]), .CI(C[45]), 
        .S(S[45]), .CO(C[46]) );
  FA_3026 \FA_INST_0[0].FA_INST_1[46].FA_  ( .A(A[46]), .B(B[46]), .CI(C[46]), 
        .S(S[46]), .CO(C[47]) );
  FA_3025 \FA_INST_0[0].FA_INST_1[47].FA_  ( .A(A[47]), .B(B[47]), .CI(C[47]), 
        .S(S[47]), .CO(C[48]) );
  FA_3024 \FA_INST_0[0].FA_INST_1[48].FA_  ( .A(A[48]), .B(B[48]), .CI(C[48]), 
        .S(S[48]), .CO(C[49]) );
  FA_3023 \FA_INST_0[0].FA_INST_1[49].FA_  ( .A(A[49]), .B(B[49]), .CI(C[49]), 
        .S(S[49]), .CO(C[50]) );
  FA_3022 \FA_INST_0[0].FA_INST_1[50].FA_  ( .A(A[50]), .B(B[50]), .CI(C[50]), 
        .S(S[50]), .CO(C[51]) );
  FA_3021 \FA_INST_0[0].FA_INST_1[51].FA_  ( .A(A[51]), .B(B[51]), .CI(C[51]), 
        .S(S[51]), .CO(C[52]) );
  FA_3020 \FA_INST_0[0].FA_INST_1[52].FA_  ( .A(A[52]), .B(B[52]), .CI(C[52]), 
        .S(S[52]), .CO(C[53]) );
  FA_3019 \FA_INST_0[0].FA_INST_1[53].FA_  ( .A(A[53]), .B(B[53]), .CI(C[53]), 
        .S(S[53]), .CO(C[54]) );
  FA_3018 \FA_INST_0[0].FA_INST_1[54].FA_  ( .A(A[54]), .B(B[54]), .CI(C[54]), 
        .S(S[54]), .CO(C[55]) );
  FA_3017 \FA_INST_0[0].FA_INST_1[55].FA_  ( .A(A[55]), .B(B[55]), .CI(C[55]), 
        .S(S[55]), .CO(C[56]) );
  FA_3016 \FA_INST_0[0].FA_INST_1[56].FA_  ( .A(A[56]), .B(B[56]), .CI(C[56]), 
        .S(S[56]), .CO(C[57]) );
  FA_3015 \FA_INST_0[0].FA_INST_1[57].FA_  ( .A(A[57]), .B(B[57]), .CI(C[57]), 
        .S(S[57]), .CO(C[58]) );
  FA_3014 \FA_INST_0[0].FA_INST_1[58].FA_  ( .A(A[58]), .B(B[58]), .CI(C[58]), 
        .S(S[58]), .CO(C[59]) );
  FA_3013 \FA_INST_0[0].FA_INST_1[59].FA_  ( .A(A[59]), .B(B[59]), .CI(C[59]), 
        .S(S[59]), .CO(C[60]) );
  FA_3012 \FA_INST_0[0].FA_INST_1[60].FA_  ( .A(A[60]), .B(B[60]), .CI(C[60]), 
        .S(S[60]), .CO(C[61]) );
  FA_3011 \FA_INST_0[0].FA_INST_1[61].FA_  ( .A(A[61]), .B(B[61]), .CI(C[61]), 
        .S(S[61]), .CO(C[62]) );
  FA_3010 \FA_INST_0[0].FA_INST_1[62].FA_  ( .A(A[62]), .B(B[62]), .CI(C[62]), 
        .S(S[62]), .CO(C[63]) );
  FA_3009 \FA_INST_0[0].FA_INST_1[63].FA_  ( .A(A[63]), .B(B[63]), .CI(C[63]), 
        .S(S[63]), .CO(C[64]) );
  FA_3008 \FA_INST_0[0].FA_INST_1[64].FA_  ( .A(A[64]), .B(B[64]), .CI(C[64]), 
        .S(S[64]), .CO(C[65]) );
  FA_3007 \FA_INST_0[0].FA_INST_1[65].FA_  ( .A(A[65]), .B(B[65]), .CI(C[65]), 
        .S(S[65]), .CO(C[66]) );
  FA_3006 \FA_INST_0[0].FA_INST_1[66].FA_  ( .A(A[66]), .B(B[66]), .CI(C[66]), 
        .S(S[66]), .CO(C[67]) );
  FA_3005 \FA_INST_0[0].FA_INST_1[67].FA_  ( .A(A[67]), .B(B[67]), .CI(C[67]), 
        .S(S[67]), .CO(C[68]) );
  FA_3004 \FA_INST_0[0].FA_INST_1[68].FA_  ( .A(A[68]), .B(B[68]), .CI(C[68]), 
        .S(S[68]), .CO(C[69]) );
  FA_3003 \FA_INST_0[0].FA_INST_1[69].FA_  ( .A(A[69]), .B(B[69]), .CI(C[69]), 
        .S(S[69]), .CO(C[70]) );
  FA_3002 \FA_INST_0[0].FA_INST_1[70].FA_  ( .A(A[70]), .B(B[70]), .CI(C[70]), 
        .S(S[70]), .CO(C[71]) );
  FA_3001 \FA_INST_0[0].FA_INST_1[71].FA_  ( .A(A[71]), .B(B[71]), .CI(C[71]), 
        .S(S[71]), .CO(C[72]) );
  FA_3000 \FA_INST_0[0].FA_INST_1[72].FA_  ( .A(A[72]), .B(B[72]), .CI(C[72]), 
        .S(S[72]), .CO(C[73]) );
  FA_2999 \FA_INST_0[0].FA_INST_1[73].FA_  ( .A(A[73]), .B(B[73]), .CI(C[73]), 
        .S(S[73]), .CO(C[74]) );
  FA_2998 \FA_INST_0[0].FA_INST_1[74].FA_  ( .A(A[74]), .B(B[74]), .CI(C[74]), 
        .S(S[74]), .CO(C[75]) );
  FA_2997 \FA_INST_0[0].FA_INST_1[75].FA_  ( .A(A[75]), .B(B[75]), .CI(C[75]), 
        .S(S[75]), .CO(C[76]) );
  FA_2996 \FA_INST_0[0].FA_INST_1[76].FA_  ( .A(A[76]), .B(B[76]), .CI(C[76]), 
        .S(S[76]), .CO(C[77]) );
  FA_2995 \FA_INST_0[0].FA_INST_1[77].FA_  ( .A(A[77]), .B(B[77]), .CI(C[77]), 
        .S(S[77]), .CO(C[78]) );
  FA_2994 \FA_INST_0[0].FA_INST_1[78].FA_  ( .A(A[78]), .B(B[78]), .CI(C[78]), 
        .S(S[78]), .CO(C[79]) );
  FA_2993 \FA_INST_0[0].FA_INST_1[79].FA_  ( .A(A[79]), .B(B[79]), .CI(C[79]), 
        .S(S[79]), .CO(C[80]) );
  FA_2992 \FA_INST_0[0].FA_INST_1[80].FA_  ( .A(A[80]), .B(B[80]), .CI(C[80]), 
        .S(S[80]), .CO(C[81]) );
  FA_2991 \FA_INST_0[0].FA_INST_1[81].FA_  ( .A(A[81]), .B(B[81]), .CI(C[81]), 
        .S(S[81]), .CO(C[82]) );
  FA_2990 \FA_INST_0[0].FA_INST_1[82].FA_  ( .A(A[82]), .B(B[82]), .CI(C[82]), 
        .S(S[82]), .CO(C[83]) );
  FA_2989 \FA_INST_0[0].FA_INST_1[83].FA_  ( .A(A[83]), .B(B[83]), .CI(C[83]), 
        .S(S[83]), .CO(C[84]) );
  FA_2988 \FA_INST_0[0].FA_INST_1[84].FA_  ( .A(A[84]), .B(B[84]), .CI(C[84]), 
        .S(S[84]), .CO(C[85]) );
  FA_2987 \FA_INST_0[0].FA_INST_1[85].FA_  ( .A(A[85]), .B(B[85]), .CI(C[85]), 
        .S(S[85]), .CO(C[86]) );
  FA_2986 \FA_INST_0[0].FA_INST_1[86].FA_  ( .A(A[86]), .B(B[86]), .CI(C[86]), 
        .S(S[86]), .CO(C[87]) );
  FA_2985 \FA_INST_0[0].FA_INST_1[87].FA_  ( .A(A[87]), .B(B[87]), .CI(C[87]), 
        .S(S[87]), .CO(C[88]) );
  FA_2984 \FA_INST_0[0].FA_INST_1[88].FA_  ( .A(A[88]), .B(B[88]), .CI(C[88]), 
        .S(S[88]), .CO(C[89]) );
  FA_2983 \FA_INST_0[0].FA_INST_1[89].FA_  ( .A(A[89]), .B(B[89]), .CI(C[89]), 
        .S(S[89]), .CO(C[90]) );
  FA_2982 \FA_INST_0[0].FA_INST_1[90].FA_  ( .A(A[90]), .B(B[90]), .CI(C[90]), 
        .S(S[90]), .CO(C[91]) );
  FA_2981 \FA_INST_0[0].FA_INST_1[91].FA_  ( .A(A[91]), .B(B[91]), .CI(C[91]), 
        .S(S[91]), .CO(C[92]) );
  FA_2980 \FA_INST_0[0].FA_INST_1[92].FA_  ( .A(A[92]), .B(B[92]), .CI(C[92]), 
        .S(S[92]), .CO(C[93]) );
  FA_2979 \FA_INST_0[0].FA_INST_1[93].FA_  ( .A(A[93]), .B(B[93]), .CI(C[93]), 
        .S(S[93]), .CO(C[94]) );
  FA_2978 \FA_INST_0[0].FA_INST_1[94].FA_  ( .A(A[94]), .B(B[94]), .CI(C[94]), 
        .S(S[94]), .CO(C[95]) );
  FA_2977 \FA_INST_0[0].FA_INST_1[95].FA_  ( .A(A[95]), .B(B[95]), .CI(C[95]), 
        .S(S[95]), .CO(C[96]) );
  FA_2976 \FA_INST_0[0].FA_INST_1[96].FA_  ( .A(A[96]), .B(B[96]), .CI(C[96]), 
        .S(S[96]), .CO(C[97]) );
  FA_2975 \FA_INST_0[0].FA_INST_1[97].FA_  ( .A(A[97]), .B(B[97]), .CI(C[97]), 
        .S(S[97]), .CO(C[98]) );
  FA_2974 \FA_INST_0[0].FA_INST_1[98].FA_  ( .A(A[98]), .B(B[98]), .CI(C[98]), 
        .S(S[98]), .CO(C[99]) );
  FA_2973 \FA_INST_0[0].FA_INST_1[99].FA_  ( .A(A[99]), .B(B[99]), .CI(C[99]), 
        .S(S[99]), .CO(C[100]) );
  FA_2972 \FA_INST_0[0].FA_INST_1[100].FA_  ( .A(A[100]), .B(B[100]), .CI(
        C[100]), .S(S[100]), .CO(C[101]) );
  FA_2971 \FA_INST_0[0].FA_INST_1[101].FA_  ( .A(A[101]), .B(B[101]), .CI(
        C[101]), .S(S[101]), .CO(C[102]) );
  FA_2970 \FA_INST_0[0].FA_INST_1[102].FA_  ( .A(A[102]), .B(B[102]), .CI(
        C[102]), .S(S[102]), .CO(C[103]) );
  FA_2969 \FA_INST_0[0].FA_INST_1[103].FA_  ( .A(A[103]), .B(B[103]), .CI(
        C[103]), .S(S[103]), .CO(C[104]) );
  FA_2968 \FA_INST_0[0].FA_INST_1[104].FA_  ( .A(A[104]), .B(B[104]), .CI(
        C[104]), .S(S[104]), .CO(C[105]) );
  FA_2967 \FA_INST_0[0].FA_INST_1[105].FA_  ( .A(A[105]), .B(B[105]), .CI(
        C[105]), .S(S[105]), .CO(C[106]) );
  FA_2966 \FA_INST_0[0].FA_INST_1[106].FA_  ( .A(A[106]), .B(B[106]), .CI(
        C[106]), .S(S[106]), .CO(C[107]) );
  FA_2965 \FA_INST_0[0].FA_INST_1[107].FA_  ( .A(A[107]), .B(B[107]), .CI(
        C[107]), .S(S[107]), .CO(C[108]) );
  FA_2964 \FA_INST_0[0].FA_INST_1[108].FA_  ( .A(A[108]), .B(B[108]), .CI(
        C[108]), .S(S[108]), .CO(C[109]) );
  FA_2963 \FA_INST_0[0].FA_INST_1[109].FA_  ( .A(A[109]), .B(B[109]), .CI(
        C[109]), .S(S[109]), .CO(C[110]) );
  FA_2962 \FA_INST_0[0].FA_INST_1[110].FA_  ( .A(A[110]), .B(B[110]), .CI(
        C[110]), .S(S[110]), .CO(C[111]) );
  FA_2961 \FA_INST_0[0].FA_INST_1[111].FA_  ( .A(A[111]), .B(B[111]), .CI(
        C[111]), .S(S[111]), .CO(C[112]) );
  FA_2960 \FA_INST_0[0].FA_INST_1[112].FA_  ( .A(A[112]), .B(B[112]), .CI(
        C[112]), .S(S[112]), .CO(C[113]) );
  FA_2959 \FA_INST_0[0].FA_INST_1[113].FA_  ( .A(A[113]), .B(B[113]), .CI(
        C[113]), .S(S[113]), .CO(C[114]) );
  FA_2958 \FA_INST_0[0].FA_INST_1[114].FA_  ( .A(A[114]), .B(B[114]), .CI(
        C[114]), .S(S[114]), .CO(C[115]) );
  FA_2957 \FA_INST_0[0].FA_INST_1[115].FA_  ( .A(A[115]), .B(B[115]), .CI(
        C[115]), .S(S[115]), .CO(C[116]) );
  FA_2956 \FA_INST_0[0].FA_INST_1[116].FA_  ( .A(A[116]), .B(B[116]), .CI(
        C[116]), .S(S[116]), .CO(C[117]) );
  FA_2955 \FA_INST_0[0].FA_INST_1[117].FA_  ( .A(A[117]), .B(B[117]), .CI(
        C[117]), .S(S[117]), .CO(C[118]) );
  FA_2954 \FA_INST_0[0].FA_INST_1[118].FA_  ( .A(A[118]), .B(B[118]), .CI(
        C[118]), .S(S[118]), .CO(C[119]) );
  FA_2953 \FA_INST_0[0].FA_INST_1[119].FA_  ( .A(A[119]), .B(B[119]), .CI(
        C[119]), .S(S[119]), .CO(C[120]) );
  FA_2952 \FA_INST_0[0].FA_INST_1[120].FA_  ( .A(A[120]), .B(B[120]), .CI(
        C[120]), .S(S[120]), .CO(C[121]) );
  FA_2951 \FA_INST_0[0].FA_INST_1[121].FA_  ( .A(A[121]), .B(B[121]), .CI(
        C[121]), .S(S[121]), .CO(C[122]) );
  FA_2950 \FA_INST_0[0].FA_INST_1[122].FA_  ( .A(A[122]), .B(B[122]), .CI(
        C[122]), .S(S[122]), .CO(C[123]) );
  FA_2949 \FA_INST_0[0].FA_INST_1[123].FA_  ( .A(A[123]), .B(B[123]), .CI(
        C[123]), .S(S[123]), .CO(C[124]) );
  FA_2948 \FA_INST_0[0].FA_INST_1[124].FA_  ( .A(A[124]), .B(B[124]), .CI(
        C[124]), .S(S[124]), .CO(C[125]) );
  FA_2947 \FA_INST_0[0].FA_INST_1[125].FA_  ( .A(A[125]), .B(B[125]), .CI(
        C[125]), .S(S[125]), .CO(C[126]) );
  FA_2946 \FA_INST_0[0].FA_INST_1[126].FA_  ( .A(A[126]), .B(B[126]), .CI(
        C[126]), .S(S[126]), .CO(C[127]) );
  FA_2945 \FA_INST_0[0].FA_INST_1[127].FA_  ( .A(A[127]), .B(B[127]), .CI(
        C[127]), .S(S[127]), .CO(C[128]) );
  FA_2944 \FA_INST_0[0].FA_INST_1[128].FA_  ( .A(A[128]), .B(B[128]), .CI(
        C[128]), .S(S[128]), .CO(C[129]) );
  FA_2943 \FA_INST_0[0].FA_INST_1[129].FA_  ( .A(A[129]), .B(B[129]), .CI(
        C[129]), .S(S[129]), .CO(C[130]) );
  FA_2942 \FA_INST_0[0].FA_INST_1[130].FA_  ( .A(A[130]), .B(B[130]), .CI(
        C[130]), .S(S[130]), .CO(C[131]) );
  FA_2941 \FA_INST_0[0].FA_INST_1[131].FA_  ( .A(A[131]), .B(B[131]), .CI(
        C[131]), .S(S[131]), .CO(C[132]) );
  FA_2940 \FA_INST_0[0].FA_INST_1[132].FA_  ( .A(A[132]), .B(B[132]), .CI(
        C[132]), .S(S[132]), .CO(C[133]) );
  FA_2939 \FA_INST_0[0].FA_INST_1[133].FA_  ( .A(A[133]), .B(B[133]), .CI(
        C[133]), .S(S[133]), .CO(C[134]) );
  FA_2938 \FA_INST_0[0].FA_INST_1[134].FA_  ( .A(A[134]), .B(B[134]), .CI(
        C[134]), .S(S[134]), .CO(C[135]) );
  FA_2937 \FA_INST_0[0].FA_INST_1[135].FA_  ( .A(A[135]), .B(B[135]), .CI(
        C[135]), .S(S[135]), .CO(C[136]) );
  FA_2936 \FA_INST_0[0].FA_INST_1[136].FA_  ( .A(A[136]), .B(B[136]), .CI(
        C[136]), .S(S[136]), .CO(C[137]) );
  FA_2935 \FA_INST_0[0].FA_INST_1[137].FA_  ( .A(A[137]), .B(B[137]), .CI(
        C[137]), .S(S[137]), .CO(C[138]) );
  FA_2934 \FA_INST_0[0].FA_INST_1[138].FA_  ( .A(A[138]), .B(B[138]), .CI(
        C[138]), .S(S[138]), .CO(C[139]) );
  FA_2933 \FA_INST_0[0].FA_INST_1[139].FA_  ( .A(A[139]), .B(B[139]), .CI(
        C[139]), .S(S[139]), .CO(C[140]) );
  FA_2932 \FA_INST_0[0].FA_INST_1[140].FA_  ( .A(A[140]), .B(B[140]), .CI(
        C[140]), .S(S[140]), .CO(C[141]) );
  FA_2931 \FA_INST_0[0].FA_INST_1[141].FA_  ( .A(A[141]), .B(B[141]), .CI(
        C[141]), .S(S[141]), .CO(C[142]) );
  FA_2930 \FA_INST_0[0].FA_INST_1[142].FA_  ( .A(A[142]), .B(B[142]), .CI(
        C[142]), .S(S[142]), .CO(C[143]) );
  FA_2929 \FA_INST_0[0].FA_INST_1[143].FA_  ( .A(A[143]), .B(B[143]), .CI(
        C[143]), .S(S[143]), .CO(C[144]) );
  FA_2928 \FA_INST_0[0].FA_INST_1[144].FA_  ( .A(A[144]), .B(B[144]), .CI(
        C[144]), .S(S[144]), .CO(C[145]) );
  FA_2927 \FA_INST_0[0].FA_INST_1[145].FA_  ( .A(A[145]), .B(B[145]), .CI(
        C[145]), .S(S[145]), .CO(C[146]) );
  FA_2926 \FA_INST_0[0].FA_INST_1[146].FA_  ( .A(A[146]), .B(B[146]), .CI(
        C[146]), .S(S[146]), .CO(C[147]) );
  FA_2925 \FA_INST_0[0].FA_INST_1[147].FA_  ( .A(A[147]), .B(B[147]), .CI(
        C[147]), .S(S[147]), .CO(C[148]) );
  FA_2924 \FA_INST_0[0].FA_INST_1[148].FA_  ( .A(A[148]), .B(B[148]), .CI(
        C[148]), .S(S[148]), .CO(C[149]) );
  FA_2923 \FA_INST_0[0].FA_INST_1[149].FA_  ( .A(A[149]), .B(B[149]), .CI(
        C[149]), .S(S[149]), .CO(C[150]) );
  FA_2922 \FA_INST_0[0].FA_INST_1[150].FA_  ( .A(A[150]), .B(B[150]), .CI(
        C[150]), .S(S[150]), .CO(C[151]) );
  FA_2921 \FA_INST_0[0].FA_INST_1[151].FA_  ( .A(A[151]), .B(B[151]), .CI(
        C[151]), .S(S[151]), .CO(C[152]) );
  FA_2920 \FA_INST_0[0].FA_INST_1[152].FA_  ( .A(A[152]), .B(B[152]), .CI(
        C[152]), .S(S[152]), .CO(C[153]) );
  FA_2919 \FA_INST_0[0].FA_INST_1[153].FA_  ( .A(A[153]), .B(B[153]), .CI(
        C[153]), .S(S[153]), .CO(C[154]) );
  FA_2918 \FA_INST_0[0].FA_INST_1[154].FA_  ( .A(A[154]), .B(B[154]), .CI(
        C[154]), .S(S[154]), .CO(C[155]) );
  FA_2917 \FA_INST_0[0].FA_INST_1[155].FA_  ( .A(A[155]), .B(B[155]), .CI(
        C[155]), .S(S[155]), .CO(C[156]) );
  FA_2916 \FA_INST_0[0].FA_INST_1[156].FA_  ( .A(A[156]), .B(B[156]), .CI(
        C[156]), .S(S[156]), .CO(C[157]) );
  FA_2915 \FA_INST_0[0].FA_INST_1[157].FA_  ( .A(A[157]), .B(B[157]), .CI(
        C[157]), .S(S[157]), .CO(C[158]) );
  FA_2914 \FA_INST_0[0].FA_INST_1[158].FA_  ( .A(A[158]), .B(B[158]), .CI(
        C[158]), .S(S[158]), .CO(C[159]) );
  FA_2913 \FA_INST_0[0].FA_INST_1[159].FA_  ( .A(A[159]), .B(B[159]), .CI(
        C[159]), .S(S[159]), .CO(C[160]) );
  FA_2912 \FA_INST_0[0].FA_INST_1[160].FA_  ( .A(A[160]), .B(B[160]), .CI(
        C[160]), .S(S[160]), .CO(C[161]) );
  FA_2911 \FA_INST_0[0].FA_INST_1[161].FA_  ( .A(A[161]), .B(B[161]), .CI(
        C[161]), .S(S[161]), .CO(C[162]) );
  FA_2910 \FA_INST_0[0].FA_INST_1[162].FA_  ( .A(A[162]), .B(B[162]), .CI(
        C[162]), .S(S[162]), .CO(C[163]) );
  FA_2909 \FA_INST_0[0].FA_INST_1[163].FA_  ( .A(A[163]), .B(B[163]), .CI(
        C[163]), .S(S[163]), .CO(C[164]) );
  FA_2908 \FA_INST_0[0].FA_INST_1[164].FA_  ( .A(A[164]), .B(B[164]), .CI(
        C[164]), .S(S[164]), .CO(C[165]) );
  FA_2907 \FA_INST_0[0].FA_INST_1[165].FA_  ( .A(A[165]), .B(B[165]), .CI(
        C[165]), .S(S[165]), .CO(C[166]) );
  FA_2906 \FA_INST_0[0].FA_INST_1[166].FA_  ( .A(A[166]), .B(B[166]), .CI(
        C[166]), .S(S[166]), .CO(C[167]) );
  FA_2905 \FA_INST_0[0].FA_INST_1[167].FA_  ( .A(A[167]), .B(B[167]), .CI(
        C[167]), .S(S[167]), .CO(C[168]) );
  FA_2904 \FA_INST_0[0].FA_INST_1[168].FA_  ( .A(A[168]), .B(B[168]), .CI(
        C[168]), .S(S[168]), .CO(C[169]) );
  FA_2903 \FA_INST_0[0].FA_INST_1[169].FA_  ( .A(A[169]), .B(B[169]), .CI(
        C[169]), .S(S[169]), .CO(C[170]) );
  FA_2902 \FA_INST_0[0].FA_INST_1[170].FA_  ( .A(A[170]), .B(B[170]), .CI(
        C[170]), .S(S[170]), .CO(C[171]) );
  FA_2901 \FA_INST_0[0].FA_INST_1[171].FA_  ( .A(A[171]), .B(B[171]), .CI(
        C[171]), .S(S[171]), .CO(C[172]) );
  FA_2900 \FA_INST_0[0].FA_INST_1[172].FA_  ( .A(A[172]), .B(B[172]), .CI(
        C[172]), .S(S[172]), .CO(C[173]) );
  FA_2899 \FA_INST_0[0].FA_INST_1[173].FA_  ( .A(A[173]), .B(B[173]), .CI(
        C[173]), .S(S[173]), .CO(C[174]) );
  FA_2898 \FA_INST_0[0].FA_INST_1[174].FA_  ( .A(A[174]), .B(B[174]), .CI(
        C[174]), .S(S[174]), .CO(C[175]) );
  FA_2897 \FA_INST_0[0].FA_INST_1[175].FA_  ( .A(A[175]), .B(B[175]), .CI(
        C[175]), .S(S[175]), .CO(C[176]) );
  FA_2896 \FA_INST_0[0].FA_INST_1[176].FA_  ( .A(A[176]), .B(B[176]), .CI(
        C[176]), .S(S[176]), .CO(C[177]) );
  FA_2895 \FA_INST_0[0].FA_INST_1[177].FA_  ( .A(A[177]), .B(B[177]), .CI(
        C[177]), .S(S[177]), .CO(C[178]) );
  FA_2894 \FA_INST_0[0].FA_INST_1[178].FA_  ( .A(A[178]), .B(B[178]), .CI(
        C[178]), .S(S[178]), .CO(C[179]) );
  FA_2893 \FA_INST_0[0].FA_INST_1[179].FA_  ( .A(A[179]), .B(B[179]), .CI(
        C[179]), .S(S[179]), .CO(C[180]) );
  FA_2892 \FA_INST_0[0].FA_INST_1[180].FA_  ( .A(A[180]), .B(B[180]), .CI(
        C[180]), .S(S[180]), .CO(C[181]) );
  FA_2891 \FA_INST_0[0].FA_INST_1[181].FA_  ( .A(A[181]), .B(B[181]), .CI(
        C[181]), .S(S[181]), .CO(C[182]) );
  FA_2890 \FA_INST_0[0].FA_INST_1[182].FA_  ( .A(A[182]), .B(B[182]), .CI(
        C[182]), .S(S[182]), .CO(C[183]) );
  FA_2889 \FA_INST_0[0].FA_INST_1[183].FA_  ( .A(A[183]), .B(B[183]), .CI(
        C[183]), .S(S[183]), .CO(C[184]) );
  FA_2888 \FA_INST_0[0].FA_INST_1[184].FA_  ( .A(A[184]), .B(B[184]), .CI(
        C[184]), .S(S[184]), .CO(C[185]) );
  FA_2887 \FA_INST_0[0].FA_INST_1[185].FA_  ( .A(A[185]), .B(B[185]), .CI(
        C[185]), .S(S[185]), .CO(C[186]) );
  FA_2886 \FA_INST_0[0].FA_INST_1[186].FA_  ( .A(A[186]), .B(B[186]), .CI(
        C[186]), .S(S[186]), .CO(C[187]) );
  FA_2885 \FA_INST_0[0].FA_INST_1[187].FA_  ( .A(A[187]), .B(B[187]), .CI(
        C[187]), .S(S[187]), .CO(C[188]) );
  FA_2884 \FA_INST_0[0].FA_INST_1[188].FA_  ( .A(A[188]), .B(B[188]), .CI(
        C[188]), .S(S[188]), .CO(C[189]) );
  FA_2883 \FA_INST_0[0].FA_INST_1[189].FA_  ( .A(A[189]), .B(B[189]), .CI(
        C[189]), .S(S[189]), .CO(C[190]) );
  FA_2882 \FA_INST_0[0].FA_INST_1[190].FA_  ( .A(A[190]), .B(B[190]), .CI(
        C[190]), .S(S[190]), .CO(C[191]) );
  FA_2881 \FA_INST_0[0].FA_INST_1[191].FA_  ( .A(A[191]), .B(B[191]), .CI(
        C[191]), .S(S[191]), .CO(C[192]) );
  FA_2880 \FA_INST_0[0].FA_INST_1[192].FA_  ( .A(A[192]), .B(B[192]), .CI(
        C[192]), .S(S[192]), .CO(C[193]) );
  FA_2879 \FA_INST_0[0].FA_INST_1[193].FA_  ( .A(A[193]), .B(B[193]), .CI(
        C[193]), .S(S[193]), .CO(C[194]) );
  FA_2878 \FA_INST_0[0].FA_INST_1[194].FA_  ( .A(A[194]), .B(B[194]), .CI(
        C[194]), .S(S[194]), .CO(C[195]) );
  FA_2877 \FA_INST_0[0].FA_INST_1[195].FA_  ( .A(A[195]), .B(B[195]), .CI(
        C[195]), .S(S[195]), .CO(C[196]) );
  FA_2876 \FA_INST_0[0].FA_INST_1[196].FA_  ( .A(A[196]), .B(B[196]), .CI(
        C[196]), .S(S[196]), .CO(C[197]) );
  FA_2875 \FA_INST_0[0].FA_INST_1[197].FA_  ( .A(A[197]), .B(B[197]), .CI(
        C[197]), .S(S[197]), .CO(C[198]) );
  FA_2874 \FA_INST_0[0].FA_INST_1[198].FA_  ( .A(A[198]), .B(B[198]), .CI(
        C[198]), .S(S[198]), .CO(C[199]) );
  FA_2873 \FA_INST_0[0].FA_INST_1[199].FA_  ( .A(A[199]), .B(B[199]), .CI(
        C[199]), .S(S[199]), .CO(C[200]) );
  FA_2872 \FA_INST_0[0].FA_INST_1[200].FA_  ( .A(A[200]), .B(B[200]), .CI(
        C[200]), .S(S[200]), .CO(C[201]) );
  FA_2871 \FA_INST_0[0].FA_INST_1[201].FA_  ( .A(A[201]), .B(B[201]), .CI(
        C[201]), .S(S[201]), .CO(C[202]) );
  FA_2870 \FA_INST_0[0].FA_INST_1[202].FA_  ( .A(A[202]), .B(B[202]), .CI(
        C[202]), .S(S[202]), .CO(C[203]) );
  FA_2869 \FA_INST_0[0].FA_INST_1[203].FA_  ( .A(A[203]), .B(B[203]), .CI(
        C[203]), .S(S[203]), .CO(C[204]) );
  FA_2868 \FA_INST_0[0].FA_INST_1[204].FA_  ( .A(A[204]), .B(B[204]), .CI(
        C[204]), .S(S[204]), .CO(C[205]) );
  FA_2867 \FA_INST_0[0].FA_INST_1[205].FA_  ( .A(A[205]), .B(B[205]), .CI(
        C[205]), .S(S[205]), .CO(C[206]) );
  FA_2866 \FA_INST_0[0].FA_INST_1[206].FA_  ( .A(A[206]), .B(B[206]), .CI(
        C[206]), .S(S[206]), .CO(C[207]) );
  FA_2865 \FA_INST_0[0].FA_INST_1[207].FA_  ( .A(A[207]), .B(B[207]), .CI(
        C[207]), .S(S[207]), .CO(C[208]) );
  FA_2864 \FA_INST_0[0].FA_INST_1[208].FA_  ( .A(A[208]), .B(B[208]), .CI(
        C[208]), .S(S[208]), .CO(C[209]) );
  FA_2863 \FA_INST_0[0].FA_INST_1[209].FA_  ( .A(A[209]), .B(B[209]), .CI(
        C[209]), .S(S[209]), .CO(C[210]) );
  FA_2862 \FA_INST_0[0].FA_INST_1[210].FA_  ( .A(A[210]), .B(B[210]), .CI(
        C[210]), .S(S[210]), .CO(C[211]) );
  FA_2861 \FA_INST_0[0].FA_INST_1[211].FA_  ( .A(A[211]), .B(B[211]), .CI(
        C[211]), .S(S[211]), .CO(C[212]) );
  FA_2860 \FA_INST_0[0].FA_INST_1[212].FA_  ( .A(A[212]), .B(B[212]), .CI(
        C[212]), .S(S[212]), .CO(C[213]) );
  FA_2859 \FA_INST_0[0].FA_INST_1[213].FA_  ( .A(A[213]), .B(B[213]), .CI(
        C[213]), .S(S[213]), .CO(C[214]) );
  FA_2858 \FA_INST_0[0].FA_INST_1[214].FA_  ( .A(A[214]), .B(B[214]), .CI(
        C[214]), .S(S[214]), .CO(C[215]) );
  FA_2857 \FA_INST_0[0].FA_INST_1[215].FA_  ( .A(A[215]), .B(B[215]), .CI(
        C[215]), .S(S[215]), .CO(C[216]) );
  FA_2856 \FA_INST_0[0].FA_INST_1[216].FA_  ( .A(A[216]), .B(B[216]), .CI(
        C[216]), .S(S[216]), .CO(C[217]) );
  FA_2855 \FA_INST_0[0].FA_INST_1[217].FA_  ( .A(A[217]), .B(B[217]), .CI(
        C[217]), .S(S[217]), .CO(C[218]) );
  FA_2854 \FA_INST_0[0].FA_INST_1[218].FA_  ( .A(A[218]), .B(B[218]), .CI(
        C[218]), .S(S[218]), .CO(C[219]) );
  FA_2853 \FA_INST_0[0].FA_INST_1[219].FA_  ( .A(A[219]), .B(B[219]), .CI(
        C[219]), .S(S[219]), .CO(C[220]) );
  FA_2852 \FA_INST_0[0].FA_INST_1[220].FA_  ( .A(A[220]), .B(B[220]), .CI(
        C[220]), .S(S[220]), .CO(C[221]) );
  FA_2851 \FA_INST_0[0].FA_INST_1[221].FA_  ( .A(A[221]), .B(B[221]), .CI(
        C[221]), .S(S[221]), .CO(C[222]) );
  FA_2850 \FA_INST_0[0].FA_INST_1[222].FA_  ( .A(A[222]), .B(B[222]), .CI(
        C[222]), .S(S[222]), .CO(C[223]) );
  FA_2849 \FA_INST_0[0].FA_INST_1[223].FA_  ( .A(A[223]), .B(B[223]), .CI(
        C[223]), .S(S[223]), .CO(C[224]) );
  FA_2848 \FA_INST_0[0].FA_INST_1[224].FA_  ( .A(A[224]), .B(B[224]), .CI(
        C[224]), .S(S[224]), .CO(C[225]) );
  FA_2847 \FA_INST_0[0].FA_INST_1[225].FA_  ( .A(A[225]), .B(B[225]), .CI(
        C[225]), .S(S[225]), .CO(C[226]) );
  FA_2846 \FA_INST_0[0].FA_INST_1[226].FA_  ( .A(A[226]), .B(B[226]), .CI(
        C[226]), .S(S[226]), .CO(C[227]) );
  FA_2845 \FA_INST_0[0].FA_INST_1[227].FA_  ( .A(A[227]), .B(B[227]), .CI(
        C[227]), .S(S[227]), .CO(C[228]) );
  FA_2844 \FA_INST_0[0].FA_INST_1[228].FA_  ( .A(A[228]), .B(B[228]), .CI(
        C[228]), .S(S[228]), .CO(C[229]) );
  FA_2843 \FA_INST_0[0].FA_INST_1[229].FA_  ( .A(A[229]), .B(B[229]), .CI(
        C[229]), .S(S[229]), .CO(C[230]) );
  FA_2842 \FA_INST_0[0].FA_INST_1[230].FA_  ( .A(A[230]), .B(B[230]), .CI(
        C[230]), .S(S[230]), .CO(C[231]) );
  FA_2841 \FA_INST_0[0].FA_INST_1[231].FA_  ( .A(A[231]), .B(B[231]), .CI(
        C[231]), .S(S[231]), .CO(C[232]) );
  FA_2840 \FA_INST_0[0].FA_INST_1[232].FA_  ( .A(A[232]), .B(B[232]), .CI(
        C[232]), .S(S[232]), .CO(C[233]) );
  FA_2839 \FA_INST_0[0].FA_INST_1[233].FA_  ( .A(A[233]), .B(B[233]), .CI(
        C[233]), .S(S[233]), .CO(C[234]) );
  FA_2838 \FA_INST_0[0].FA_INST_1[234].FA_  ( .A(A[234]), .B(B[234]), .CI(
        C[234]), .S(S[234]), .CO(C[235]) );
  FA_2837 \FA_INST_0[0].FA_INST_1[235].FA_  ( .A(A[235]), .B(B[235]), .CI(
        C[235]), .S(S[235]), .CO(C[236]) );
  FA_2836 \FA_INST_0[0].FA_INST_1[236].FA_  ( .A(A[236]), .B(B[236]), .CI(
        C[236]), .S(S[236]), .CO(C[237]) );
  FA_2835 \FA_INST_0[0].FA_INST_1[237].FA_  ( .A(A[237]), .B(B[237]), .CI(
        C[237]), .S(S[237]), .CO(C[238]) );
  FA_2834 \FA_INST_0[0].FA_INST_1[238].FA_  ( .A(A[238]), .B(B[238]), .CI(
        C[238]), .S(S[238]), .CO(C[239]) );
  FA_2833 \FA_INST_0[0].FA_INST_1[239].FA_  ( .A(A[239]), .B(B[239]), .CI(
        C[239]), .S(S[239]), .CO(C[240]) );
  FA_2832 \FA_INST_0[0].FA_INST_1[240].FA_  ( .A(A[240]), .B(B[240]), .CI(
        C[240]), .S(S[240]), .CO(C[241]) );
  FA_2831 \FA_INST_0[0].FA_INST_1[241].FA_  ( .A(A[241]), .B(B[241]), .CI(
        C[241]), .S(S[241]), .CO(C[242]) );
  FA_2830 \FA_INST_0[0].FA_INST_1[242].FA_  ( .A(A[242]), .B(B[242]), .CI(
        C[242]), .S(S[242]), .CO(C[243]) );
  FA_2829 \FA_INST_0[0].FA_INST_1[243].FA_  ( .A(A[243]), .B(B[243]), .CI(
        C[243]), .S(S[243]), .CO(C[244]) );
  FA_2828 \FA_INST_0[0].FA_INST_1[244].FA_  ( .A(A[244]), .B(B[244]), .CI(
        C[244]), .S(S[244]), .CO(C[245]) );
  FA_2827 \FA_INST_0[0].FA_INST_1[245].FA_  ( .A(A[245]), .B(B[245]), .CI(
        C[245]), .S(S[245]), .CO(C[246]) );
  FA_2826 \FA_INST_0[0].FA_INST_1[246].FA_  ( .A(A[246]), .B(B[246]), .CI(
        C[246]), .S(S[246]), .CO(C[247]) );
  FA_2825 \FA_INST_0[0].FA_INST_1[247].FA_  ( .A(A[247]), .B(B[247]), .CI(
        C[247]), .S(S[247]), .CO(C[248]) );
  FA_2824 \FA_INST_0[0].FA_INST_1[248].FA_  ( .A(A[248]), .B(B[248]), .CI(
        C[248]), .S(S[248]), .CO(C[249]) );
  FA_2823 \FA_INST_0[0].FA_INST_1[249].FA_  ( .A(A[249]), .B(B[249]), .CI(
        C[249]), .S(S[249]), .CO(C[250]) );
  FA_2822 \FA_INST_0[0].FA_INST_1[250].FA_  ( .A(A[250]), .B(B[250]), .CI(
        C[250]), .S(S[250]), .CO(C[251]) );
  FA_2821 \FA_INST_0[0].FA_INST_1[251].FA_  ( .A(A[251]), .B(B[251]), .CI(
        C[251]), .S(S[251]), .CO(C[252]) );
  FA_2820 \FA_INST_0[0].FA_INST_1[252].FA_  ( .A(A[252]), .B(B[252]), .CI(
        C[252]), .S(S[252]), .CO(C[253]) );
  FA_2819 \FA_INST_0[0].FA_INST_1[253].FA_  ( .A(A[253]), .B(B[253]), .CI(
        C[253]), .S(S[253]), .CO(C[254]) );
  FA_2818 \FA_INST_0[0].FA_INST_1[254].FA_  ( .A(A[254]), .B(B[254]), .CI(
        C[254]), .S(S[254]), .CO(C[255]) );
  FA_2817 \FA_INST_0[0].FA_INST_1[255].FA_  ( .A(A[255]), .B(B[255]), .CI(
        C[255]), .S(S[255]), .CO(C[256]) );
  FA_2816 \FA_INST_0[0].FA_INST_1[256].FA_  ( .A(A[256]), .B(B[256]), .CI(
        C[256]), .S(S[256]), .CO(C[257]) );
  FA_2815 \FA_INST_0[0].FA_INST_1[257].FA_  ( .A(A[257]), .B(B[257]), .CI(
        C[257]), .S(S[257]), .CO(C[258]) );
  FA_2814 \FA_INST_0[0].FA_INST_1[258].FA_  ( .A(A[258]), .B(B[258]), .CI(
        C[258]), .S(S[258]), .CO(C[259]) );
  FA_2813 \FA_INST_0[0].FA_INST_1[259].FA_  ( .A(A[259]), .B(B[259]), .CI(
        C[259]), .S(S[259]), .CO(C[260]) );
  FA_2812 \FA_INST_0[0].FA_INST_1[260].FA_  ( .A(A[260]), .B(B[260]), .CI(
        C[260]), .S(S[260]), .CO(C[261]) );
  FA_2811 \FA_INST_0[0].FA_INST_1[261].FA_  ( .A(A[261]), .B(B[261]), .CI(
        C[261]), .S(S[261]), .CO(C[262]) );
  FA_2810 \FA_INST_0[0].FA_INST_1[262].FA_  ( .A(A[262]), .B(B[262]), .CI(
        C[262]), .S(S[262]), .CO(C[263]) );
  FA_2809 \FA_INST_0[0].FA_INST_1[263].FA_  ( .A(A[263]), .B(B[263]), .CI(
        C[263]), .S(S[263]), .CO(C[264]) );
  FA_2808 \FA_INST_0[0].FA_INST_1[264].FA_  ( .A(A[264]), .B(B[264]), .CI(
        C[264]), .S(S[264]), .CO(C[265]) );
  FA_2807 \FA_INST_0[0].FA_INST_1[265].FA_  ( .A(A[265]), .B(B[265]), .CI(
        C[265]), .S(S[265]), .CO(C[266]) );
  FA_2806 \FA_INST_0[0].FA_INST_1[266].FA_  ( .A(A[266]), .B(B[266]), .CI(
        C[266]), .S(S[266]), .CO(C[267]) );
  FA_2805 \FA_INST_0[0].FA_INST_1[267].FA_  ( .A(A[267]), .B(B[267]), .CI(
        C[267]), .S(S[267]), .CO(C[268]) );
  FA_2804 \FA_INST_0[0].FA_INST_1[268].FA_  ( .A(A[268]), .B(B[268]), .CI(
        C[268]), .S(S[268]), .CO(C[269]) );
  FA_2803 \FA_INST_0[0].FA_INST_1[269].FA_  ( .A(A[269]), .B(B[269]), .CI(
        C[269]), .S(S[269]), .CO(C[270]) );
  FA_2802 \FA_INST_0[0].FA_INST_1[270].FA_  ( .A(A[270]), .B(B[270]), .CI(
        C[270]), .S(S[270]), .CO(C[271]) );
  FA_2801 \FA_INST_0[0].FA_INST_1[271].FA_  ( .A(A[271]), .B(B[271]), .CI(
        C[271]), .S(S[271]), .CO(C[272]) );
  FA_2800 \FA_INST_0[0].FA_INST_1[272].FA_  ( .A(A[272]), .B(B[272]), .CI(
        C[272]), .S(S[272]), .CO(C[273]) );
  FA_2799 \FA_INST_0[0].FA_INST_1[273].FA_  ( .A(A[273]), .B(B[273]), .CI(
        C[273]), .S(S[273]), .CO(C[274]) );
  FA_2798 \FA_INST_0[0].FA_INST_1[274].FA_  ( .A(A[274]), .B(B[274]), .CI(
        C[274]), .S(S[274]), .CO(C[275]) );
  FA_2797 \FA_INST_0[0].FA_INST_1[275].FA_  ( .A(A[275]), .B(B[275]), .CI(
        C[275]), .S(S[275]), .CO(C[276]) );
  FA_2796 \FA_INST_0[0].FA_INST_1[276].FA_  ( .A(A[276]), .B(B[276]), .CI(
        C[276]), .S(S[276]), .CO(C[277]) );
  FA_2795 \FA_INST_0[0].FA_INST_1[277].FA_  ( .A(A[277]), .B(B[277]), .CI(
        C[277]), .S(S[277]), .CO(C[278]) );
  FA_2794 \FA_INST_0[0].FA_INST_1[278].FA_  ( .A(A[278]), .B(B[278]), .CI(
        C[278]), .S(S[278]), .CO(C[279]) );
  FA_2793 \FA_INST_0[0].FA_INST_1[279].FA_  ( .A(A[279]), .B(B[279]), .CI(
        C[279]), .S(S[279]), .CO(C[280]) );
  FA_2792 \FA_INST_0[0].FA_INST_1[280].FA_  ( .A(A[280]), .B(B[280]), .CI(
        C[280]), .S(S[280]), .CO(C[281]) );
  FA_2791 \FA_INST_0[0].FA_INST_1[281].FA_  ( .A(A[281]), .B(B[281]), .CI(
        C[281]), .S(S[281]), .CO(C[282]) );
  FA_2790 \FA_INST_0[0].FA_INST_1[282].FA_  ( .A(A[282]), .B(B[282]), .CI(
        C[282]), .S(S[282]), .CO(C[283]) );
  FA_2789 \FA_INST_0[0].FA_INST_1[283].FA_  ( .A(A[283]), .B(B[283]), .CI(
        C[283]), .S(S[283]), .CO(C[284]) );
  FA_2788 \FA_INST_0[0].FA_INST_1[284].FA_  ( .A(A[284]), .B(B[284]), .CI(
        C[284]), .S(S[284]), .CO(C[285]) );
  FA_2787 \FA_INST_0[0].FA_INST_1[285].FA_  ( .A(A[285]), .B(B[285]), .CI(
        C[285]), .S(S[285]), .CO(C[286]) );
  FA_2786 \FA_INST_0[0].FA_INST_1[286].FA_  ( .A(A[286]), .B(B[286]), .CI(
        C[286]), .S(S[286]), .CO(C[287]) );
  FA_2785 \FA_INST_0[0].FA_INST_1[287].FA_  ( .A(A[287]), .B(B[287]), .CI(
        C[287]), .S(S[287]), .CO(C[288]) );
  FA_2784 \FA_INST_0[0].FA_INST_1[288].FA_  ( .A(A[288]), .B(B[288]), .CI(
        C[288]), .S(S[288]), .CO(C[289]) );
  FA_2783 \FA_INST_0[0].FA_INST_1[289].FA_  ( .A(A[289]), .B(B[289]), .CI(
        C[289]), .S(S[289]), .CO(C[290]) );
  FA_2782 \FA_INST_0[0].FA_INST_1[290].FA_  ( .A(A[290]), .B(B[290]), .CI(
        C[290]), .S(S[290]), .CO(C[291]) );
  FA_2781 \FA_INST_0[0].FA_INST_1[291].FA_  ( .A(A[291]), .B(B[291]), .CI(
        C[291]), .S(S[291]), .CO(C[292]) );
  FA_2780 \FA_INST_0[0].FA_INST_1[292].FA_  ( .A(A[292]), .B(B[292]), .CI(
        C[292]), .S(S[292]), .CO(C[293]) );
  FA_2779 \FA_INST_0[0].FA_INST_1[293].FA_  ( .A(A[293]), .B(B[293]), .CI(
        C[293]), .S(S[293]), .CO(C[294]) );
  FA_2778 \FA_INST_0[0].FA_INST_1[294].FA_  ( .A(A[294]), .B(B[294]), .CI(
        C[294]), .S(S[294]), .CO(C[295]) );
  FA_2777 \FA_INST_0[0].FA_INST_1[295].FA_  ( .A(A[295]), .B(B[295]), .CI(
        C[295]), .S(S[295]), .CO(C[296]) );
  FA_2776 \FA_INST_0[0].FA_INST_1[296].FA_  ( .A(A[296]), .B(B[296]), .CI(
        C[296]), .S(S[296]), .CO(C[297]) );
  FA_2775 \FA_INST_0[0].FA_INST_1[297].FA_  ( .A(A[297]), .B(B[297]), .CI(
        C[297]), .S(S[297]), .CO(C[298]) );
  FA_2774 \FA_INST_0[0].FA_INST_1[298].FA_  ( .A(A[298]), .B(B[298]), .CI(
        C[298]), .S(S[298]), .CO(C[299]) );
  FA_2773 \FA_INST_0[0].FA_INST_1[299].FA_  ( .A(A[299]), .B(B[299]), .CI(
        C[299]), .S(S[299]), .CO(C[300]) );
  FA_2772 \FA_INST_0[0].FA_INST_1[300].FA_  ( .A(A[300]), .B(B[300]), .CI(
        C[300]), .S(S[300]), .CO(C[301]) );
  FA_2771 \FA_INST_0[0].FA_INST_1[301].FA_  ( .A(A[301]), .B(B[301]), .CI(
        C[301]), .S(S[301]), .CO(C[302]) );
  FA_2770 \FA_INST_0[0].FA_INST_1[302].FA_  ( .A(A[302]), .B(B[302]), .CI(
        C[302]), .S(S[302]), .CO(C[303]) );
  FA_2769 \FA_INST_0[0].FA_INST_1[303].FA_  ( .A(A[303]), .B(B[303]), .CI(
        C[303]), .S(S[303]), .CO(C[304]) );
  FA_2768 \FA_INST_0[0].FA_INST_1[304].FA_  ( .A(A[304]), .B(B[304]), .CI(
        C[304]), .S(S[304]), .CO(C[305]) );
  FA_2767 \FA_INST_0[0].FA_INST_1[305].FA_  ( .A(A[305]), .B(B[305]), .CI(
        C[305]), .S(S[305]), .CO(C[306]) );
  FA_2766 \FA_INST_0[0].FA_INST_1[306].FA_  ( .A(A[306]), .B(B[306]), .CI(
        C[306]), .S(S[306]), .CO(C[307]) );
  FA_2765 \FA_INST_0[0].FA_INST_1[307].FA_  ( .A(A[307]), .B(B[307]), .CI(
        C[307]), .S(S[307]), .CO(C[308]) );
  FA_2764 \FA_INST_0[0].FA_INST_1[308].FA_  ( .A(A[308]), .B(B[308]), .CI(
        C[308]), .S(S[308]), .CO(C[309]) );
  FA_2763 \FA_INST_0[0].FA_INST_1[309].FA_  ( .A(A[309]), .B(B[309]), .CI(
        C[309]), .S(S[309]), .CO(C[310]) );
  FA_2762 \FA_INST_0[0].FA_INST_1[310].FA_  ( .A(A[310]), .B(B[310]), .CI(
        C[310]), .S(S[310]), .CO(C[311]) );
  FA_2761 \FA_INST_0[0].FA_INST_1[311].FA_  ( .A(A[311]), .B(B[311]), .CI(
        C[311]), .S(S[311]), .CO(C[312]) );
  FA_2760 \FA_INST_0[0].FA_INST_1[312].FA_  ( .A(A[312]), .B(B[312]), .CI(
        C[312]), .S(S[312]), .CO(C[313]) );
  FA_2759 \FA_INST_0[0].FA_INST_1[313].FA_  ( .A(A[313]), .B(B[313]), .CI(
        C[313]), .S(S[313]), .CO(C[314]) );
  FA_2758 \FA_INST_0[0].FA_INST_1[314].FA_  ( .A(A[314]), .B(B[314]), .CI(
        C[314]), .S(S[314]), .CO(C[315]) );
  FA_2757 \FA_INST_0[0].FA_INST_1[315].FA_  ( .A(A[315]), .B(B[315]), .CI(
        C[315]), .S(S[315]), .CO(C[316]) );
  FA_2756 \FA_INST_0[0].FA_INST_1[316].FA_  ( .A(A[316]), .B(B[316]), .CI(
        C[316]), .S(S[316]), .CO(C[317]) );
  FA_2755 \FA_INST_0[0].FA_INST_1[317].FA_  ( .A(A[317]), .B(B[317]), .CI(
        C[317]), .S(S[317]), .CO(C[318]) );
  FA_2754 \FA_INST_0[0].FA_INST_1[318].FA_  ( .A(A[318]), .B(B[318]), .CI(
        C[318]), .S(S[318]), .CO(C[319]) );
  FA_2753 \FA_INST_0[0].FA_INST_1[319].FA_  ( .A(A[319]), .B(B[319]), .CI(
        C[319]), .S(S[319]), .CO(C[320]) );
  FA_2752 \FA_INST_0[0].FA_INST_1[320].FA_  ( .A(A[320]), .B(B[320]), .CI(
        C[320]), .S(S[320]), .CO(C[321]) );
  FA_2751 \FA_INST_0[0].FA_INST_1[321].FA_  ( .A(A[321]), .B(B[321]), .CI(
        C[321]), .S(S[321]), .CO(C[322]) );
  FA_2750 \FA_INST_0[0].FA_INST_1[322].FA_  ( .A(A[322]), .B(B[322]), .CI(
        C[322]), .S(S[322]), .CO(C[323]) );
  FA_2749 \FA_INST_0[0].FA_INST_1[323].FA_  ( .A(A[323]), .B(B[323]), .CI(
        C[323]), .S(S[323]), .CO(C[324]) );
  FA_2748 \FA_INST_0[0].FA_INST_1[324].FA_  ( .A(A[324]), .B(B[324]), .CI(
        C[324]), .S(S[324]), .CO(C[325]) );
  FA_2747 \FA_INST_0[0].FA_INST_1[325].FA_  ( .A(A[325]), .B(B[325]), .CI(
        C[325]), .S(S[325]), .CO(C[326]) );
  FA_2746 \FA_INST_0[0].FA_INST_1[326].FA_  ( .A(A[326]), .B(B[326]), .CI(
        C[326]), .S(S[326]), .CO(C[327]) );
  FA_2745 \FA_INST_0[0].FA_INST_1[327].FA_  ( .A(A[327]), .B(B[327]), .CI(
        C[327]), .S(S[327]), .CO(C[328]) );
  FA_2744 \FA_INST_0[0].FA_INST_1[328].FA_  ( .A(A[328]), .B(B[328]), .CI(
        C[328]), .S(S[328]), .CO(C[329]) );
  FA_2743 \FA_INST_0[0].FA_INST_1[329].FA_  ( .A(A[329]), .B(B[329]), .CI(
        C[329]), .S(S[329]), .CO(C[330]) );
  FA_2742 \FA_INST_0[0].FA_INST_1[330].FA_  ( .A(A[330]), .B(B[330]), .CI(
        C[330]), .S(S[330]), .CO(C[331]) );
  FA_2741 \FA_INST_0[0].FA_INST_1[331].FA_  ( .A(A[331]), .B(B[331]), .CI(
        C[331]), .S(S[331]), .CO(C[332]) );
  FA_2740 \FA_INST_0[0].FA_INST_1[332].FA_  ( .A(A[332]), .B(B[332]), .CI(
        C[332]), .S(S[332]), .CO(C[333]) );
  FA_2739 \FA_INST_0[0].FA_INST_1[333].FA_  ( .A(A[333]), .B(B[333]), .CI(
        C[333]), .S(S[333]), .CO(C[334]) );
  FA_2738 \FA_INST_0[0].FA_INST_1[334].FA_  ( .A(A[334]), .B(B[334]), .CI(
        C[334]), .S(S[334]), .CO(C[335]) );
  FA_2737 \FA_INST_0[0].FA_INST_1[335].FA_  ( .A(A[335]), .B(B[335]), .CI(
        C[335]), .S(S[335]), .CO(C[336]) );
  FA_2736 \FA_INST_0[0].FA_INST_1[336].FA_  ( .A(A[336]), .B(B[336]), .CI(
        C[336]), .S(S[336]), .CO(C[337]) );
  FA_2735 \FA_INST_0[0].FA_INST_1[337].FA_  ( .A(A[337]), .B(B[337]), .CI(
        C[337]), .S(S[337]), .CO(C[338]) );
  FA_2734 \FA_INST_0[0].FA_INST_1[338].FA_  ( .A(A[338]), .B(B[338]), .CI(
        C[338]), .S(S[338]), .CO(C[339]) );
  FA_2733 \FA_INST_0[0].FA_INST_1[339].FA_  ( .A(A[339]), .B(B[339]), .CI(
        C[339]), .S(S[339]), .CO(C[340]) );
  FA_2732 \FA_INST_0[0].FA_INST_1[340].FA_  ( .A(A[340]), .B(B[340]), .CI(
        C[340]), .S(S[340]), .CO(C[341]) );
  FA_2731 \FA_INST_0[0].FA_INST_1[341].FA_  ( .A(A[341]), .B(B[341]), .CI(
        C[341]), .S(S[341]), .CO(C[342]) );
  FA_2730 \FA_INST_0[0].FA_INST_1[342].FA_  ( .A(A[342]), .B(B[342]), .CI(
        C[342]), .S(S[342]), .CO(C[343]) );
  FA_2729 \FA_INST_0[0].FA_INST_1[343].FA_  ( .A(A[343]), .B(B[343]), .CI(
        C[343]), .S(S[343]), .CO(C[344]) );
  FA_2728 \FA_INST_0[0].FA_INST_1[344].FA_  ( .A(A[344]), .B(B[344]), .CI(
        C[344]), .S(S[344]), .CO(C[345]) );
  FA_2727 \FA_INST_0[0].FA_INST_1[345].FA_  ( .A(A[345]), .B(B[345]), .CI(
        C[345]), .S(S[345]), .CO(C[346]) );
  FA_2726 \FA_INST_0[0].FA_INST_1[346].FA_  ( .A(A[346]), .B(B[346]), .CI(
        C[346]), .S(S[346]), .CO(C[347]) );
  FA_2725 \FA_INST_0[0].FA_INST_1[347].FA_  ( .A(A[347]), .B(B[347]), .CI(
        C[347]), .S(S[347]), .CO(C[348]) );
  FA_2724 \FA_INST_0[0].FA_INST_1[348].FA_  ( .A(A[348]), .B(B[348]), .CI(
        C[348]), .S(S[348]), .CO(C[349]) );
  FA_2723 \FA_INST_0[0].FA_INST_1[349].FA_  ( .A(A[349]), .B(B[349]), .CI(
        C[349]), .S(S[349]), .CO(C[350]) );
  FA_2722 \FA_INST_0[0].FA_INST_1[350].FA_  ( .A(A[350]), .B(B[350]), .CI(
        C[350]), .S(S[350]), .CO(C[351]) );
  FA_2721 \FA_INST_0[0].FA_INST_1[351].FA_  ( .A(A[351]), .B(B[351]), .CI(
        C[351]), .S(S[351]), .CO(C[352]) );
  FA_2720 \FA_INST_0[0].FA_INST_1[352].FA_  ( .A(A[352]), .B(B[352]), .CI(
        C[352]), .S(S[352]), .CO(C[353]) );
  FA_2719 \FA_INST_0[0].FA_INST_1[353].FA_  ( .A(A[353]), .B(B[353]), .CI(
        C[353]), .S(S[353]), .CO(C[354]) );
  FA_2718 \FA_INST_0[0].FA_INST_1[354].FA_  ( .A(A[354]), .B(B[354]), .CI(
        C[354]), .S(S[354]), .CO(C[355]) );
  FA_2717 \FA_INST_0[0].FA_INST_1[355].FA_  ( .A(A[355]), .B(B[355]), .CI(
        C[355]), .S(S[355]), .CO(C[356]) );
  FA_2716 \FA_INST_0[0].FA_INST_1[356].FA_  ( .A(A[356]), .B(B[356]), .CI(
        C[356]), .S(S[356]), .CO(C[357]) );
  FA_2715 \FA_INST_0[0].FA_INST_1[357].FA_  ( .A(A[357]), .B(B[357]), .CI(
        C[357]), .S(S[357]), .CO(C[358]) );
  FA_2714 \FA_INST_0[0].FA_INST_1[358].FA_  ( .A(A[358]), .B(B[358]), .CI(
        C[358]), .S(S[358]), .CO(C[359]) );
  FA_2713 \FA_INST_0[0].FA_INST_1[359].FA_  ( .A(A[359]), .B(B[359]), .CI(
        C[359]), .S(S[359]), .CO(C[360]) );
  FA_2712 \FA_INST_0[0].FA_INST_1[360].FA_  ( .A(A[360]), .B(B[360]), .CI(
        C[360]), .S(S[360]), .CO(C[361]) );
  FA_2711 \FA_INST_0[0].FA_INST_1[361].FA_  ( .A(A[361]), .B(B[361]), .CI(
        C[361]), .S(S[361]), .CO(C[362]) );
  FA_2710 \FA_INST_0[0].FA_INST_1[362].FA_  ( .A(A[362]), .B(B[362]), .CI(
        C[362]), .S(S[362]), .CO(C[363]) );
  FA_2709 \FA_INST_0[0].FA_INST_1[363].FA_  ( .A(A[363]), .B(B[363]), .CI(
        C[363]), .S(S[363]), .CO(C[364]) );
  FA_2708 \FA_INST_0[0].FA_INST_1[364].FA_  ( .A(A[364]), .B(B[364]), .CI(
        C[364]), .S(S[364]), .CO(C[365]) );
  FA_2707 \FA_INST_0[0].FA_INST_1[365].FA_  ( .A(A[365]), .B(B[365]), .CI(
        C[365]), .S(S[365]), .CO(C[366]) );
  FA_2706 \FA_INST_0[0].FA_INST_1[366].FA_  ( .A(A[366]), .B(B[366]), .CI(
        C[366]), .S(S[366]), .CO(C[367]) );
  FA_2705 \FA_INST_0[0].FA_INST_1[367].FA_  ( .A(A[367]), .B(B[367]), .CI(
        C[367]), .S(S[367]), .CO(C[368]) );
  FA_2704 \FA_INST_0[0].FA_INST_1[368].FA_  ( .A(A[368]), .B(B[368]), .CI(
        C[368]), .S(S[368]), .CO(C[369]) );
  FA_2703 \FA_INST_0[0].FA_INST_1[369].FA_  ( .A(A[369]), .B(B[369]), .CI(
        C[369]), .S(S[369]), .CO(C[370]) );
  FA_2702 \FA_INST_0[0].FA_INST_1[370].FA_  ( .A(A[370]), .B(B[370]), .CI(
        C[370]), .S(S[370]), .CO(C[371]) );
  FA_2701 \FA_INST_0[0].FA_INST_1[371].FA_  ( .A(A[371]), .B(B[371]), .CI(
        C[371]), .S(S[371]), .CO(C[372]) );
  FA_2700 \FA_INST_0[0].FA_INST_1[372].FA_  ( .A(A[372]), .B(B[372]), .CI(
        C[372]), .S(S[372]), .CO(C[373]) );
  FA_2699 \FA_INST_0[0].FA_INST_1[373].FA_  ( .A(A[373]), .B(B[373]), .CI(
        C[373]), .S(S[373]), .CO(C[374]) );
  FA_2698 \FA_INST_0[0].FA_INST_1[374].FA_  ( .A(A[374]), .B(B[374]), .CI(
        C[374]), .S(S[374]), .CO(C[375]) );
  FA_2697 \FA_INST_0[0].FA_INST_1[375].FA_  ( .A(A[375]), .B(B[375]), .CI(
        C[375]), .S(S[375]), .CO(C[376]) );
  FA_2696 \FA_INST_0[0].FA_INST_1[376].FA_  ( .A(A[376]), .B(B[376]), .CI(
        C[376]), .S(S[376]), .CO(C[377]) );
  FA_2695 \FA_INST_0[0].FA_INST_1[377].FA_  ( .A(A[377]), .B(B[377]), .CI(
        C[377]), .S(S[377]), .CO(C[378]) );
  FA_2694 \FA_INST_0[0].FA_INST_1[378].FA_  ( .A(A[378]), .B(B[378]), .CI(
        C[378]), .S(S[378]), .CO(C[379]) );
  FA_2693 \FA_INST_0[0].FA_INST_1[379].FA_  ( .A(A[379]), .B(B[379]), .CI(
        C[379]), .S(S[379]), .CO(C[380]) );
  FA_2692 \FA_INST_0[0].FA_INST_1[380].FA_  ( .A(A[380]), .B(B[380]), .CI(
        C[380]), .S(S[380]), .CO(C[381]) );
  FA_2691 \FA_INST_0[0].FA_INST_1[381].FA_  ( .A(A[381]), .B(B[381]), .CI(
        C[381]), .S(S[381]), .CO(C[382]) );
  FA_2690 \FA_INST_0[0].FA_INST_1[382].FA_  ( .A(A[382]), .B(B[382]), .CI(
        C[382]), .S(S[382]), .CO(C[383]) );
  FA_2689 \FA_INST_0[0].FA_INST_1[383].FA_  ( .A(A[383]), .B(B[383]), .CI(
        C[383]), .S(S[383]), .CO(C[384]) );
  FA_2688 \FA_INST_0[0].FA_INST_1[384].FA_  ( .A(A[384]), .B(B[384]), .CI(
        C[384]), .S(S[384]), .CO(C[385]) );
  FA_2687 \FA_INST_0[0].FA_INST_1[385].FA_  ( .A(A[385]), .B(B[385]), .CI(
        C[385]), .S(S[385]), .CO(C[386]) );
  FA_2686 \FA_INST_0[0].FA_INST_1[386].FA_  ( .A(A[386]), .B(B[386]), .CI(
        C[386]), .S(S[386]), .CO(C[387]) );
  FA_2685 \FA_INST_0[0].FA_INST_1[387].FA_  ( .A(A[387]), .B(B[387]), .CI(
        C[387]), .S(S[387]), .CO(C[388]) );
  FA_2684 \FA_INST_0[0].FA_INST_1[388].FA_  ( .A(A[388]), .B(B[388]), .CI(
        C[388]), .S(S[388]), .CO(C[389]) );
  FA_2683 \FA_INST_0[0].FA_INST_1[389].FA_  ( .A(A[389]), .B(B[389]), .CI(
        C[389]), .S(S[389]), .CO(C[390]) );
  FA_2682 \FA_INST_0[0].FA_INST_1[390].FA_  ( .A(A[390]), .B(B[390]), .CI(
        C[390]), .S(S[390]), .CO(C[391]) );
  FA_2681 \FA_INST_0[0].FA_INST_1[391].FA_  ( .A(A[391]), .B(B[391]), .CI(
        C[391]), .S(S[391]), .CO(C[392]) );
  FA_2680 \FA_INST_0[0].FA_INST_1[392].FA_  ( .A(A[392]), .B(B[392]), .CI(
        C[392]), .S(S[392]), .CO(C[393]) );
  FA_2679 \FA_INST_0[0].FA_INST_1[393].FA_  ( .A(A[393]), .B(B[393]), .CI(
        C[393]), .S(S[393]), .CO(C[394]) );
  FA_2678 \FA_INST_0[0].FA_INST_1[394].FA_  ( .A(A[394]), .B(B[394]), .CI(
        C[394]), .S(S[394]), .CO(C[395]) );
  FA_2677 \FA_INST_0[0].FA_INST_1[395].FA_  ( .A(A[395]), .B(B[395]), .CI(
        C[395]), .S(S[395]), .CO(C[396]) );
  FA_2676 \FA_INST_0[0].FA_INST_1[396].FA_  ( .A(A[396]), .B(B[396]), .CI(
        C[396]), .S(S[396]), .CO(C[397]) );
  FA_2675 \FA_INST_0[0].FA_INST_1[397].FA_  ( .A(A[397]), .B(B[397]), .CI(
        C[397]), .S(S[397]), .CO(C[398]) );
  FA_2674 \FA_INST_0[0].FA_INST_1[398].FA_  ( .A(A[398]), .B(B[398]), .CI(
        C[398]), .S(S[398]), .CO(C[399]) );
  FA_2673 \FA_INST_0[0].FA_INST_1[399].FA_  ( .A(A[399]), .B(B[399]), .CI(
        C[399]), .S(S[399]), .CO(C[400]) );
  FA_2672 \FA_INST_0[0].FA_INST_1[400].FA_  ( .A(A[400]), .B(B[400]), .CI(
        C[400]), .S(S[400]), .CO(C[401]) );
  FA_2671 \FA_INST_0[0].FA_INST_1[401].FA_  ( .A(A[401]), .B(B[401]), .CI(
        C[401]), .S(S[401]), .CO(C[402]) );
  FA_2670 \FA_INST_0[0].FA_INST_1[402].FA_  ( .A(A[402]), .B(B[402]), .CI(
        C[402]), .S(S[402]), .CO(C[403]) );
  FA_2669 \FA_INST_0[0].FA_INST_1[403].FA_  ( .A(A[403]), .B(B[403]), .CI(
        C[403]), .S(S[403]), .CO(C[404]) );
  FA_2668 \FA_INST_0[0].FA_INST_1[404].FA_  ( .A(A[404]), .B(B[404]), .CI(
        C[404]), .S(S[404]), .CO(C[405]) );
  FA_2667 \FA_INST_0[0].FA_INST_1[405].FA_  ( .A(A[405]), .B(B[405]), .CI(
        C[405]), .S(S[405]), .CO(C[406]) );
  FA_2666 \FA_INST_0[0].FA_INST_1[406].FA_  ( .A(A[406]), .B(B[406]), .CI(
        C[406]), .S(S[406]), .CO(C[407]) );
  FA_2665 \FA_INST_0[0].FA_INST_1[407].FA_  ( .A(A[407]), .B(B[407]), .CI(
        C[407]), .S(S[407]), .CO(C[408]) );
  FA_2664 \FA_INST_0[0].FA_INST_1[408].FA_  ( .A(A[408]), .B(B[408]), .CI(
        C[408]), .S(S[408]), .CO(C[409]) );
  FA_2663 \FA_INST_0[0].FA_INST_1[409].FA_  ( .A(A[409]), .B(B[409]), .CI(
        C[409]), .S(S[409]), .CO(C[410]) );
  FA_2662 \FA_INST_0[0].FA_INST_1[410].FA_  ( .A(A[410]), .B(B[410]), .CI(
        C[410]), .S(S[410]), .CO(C[411]) );
  FA_2661 \FA_INST_0[0].FA_INST_1[411].FA_  ( .A(A[411]), .B(B[411]), .CI(
        C[411]), .S(S[411]), .CO(C[412]) );
  FA_2660 \FA_INST_0[0].FA_INST_1[412].FA_  ( .A(A[412]), .B(B[412]), .CI(
        C[412]), .S(S[412]), .CO(C[413]) );
  FA_2659 \FA_INST_0[0].FA_INST_1[413].FA_  ( .A(A[413]), .B(B[413]), .CI(
        C[413]), .S(S[413]), .CO(C[414]) );
  FA_2658 \FA_INST_0[0].FA_INST_1[414].FA_  ( .A(A[414]), .B(B[414]), .CI(
        C[414]), .S(S[414]), .CO(C[415]) );
  FA_2657 \FA_INST_0[0].FA_INST_1[415].FA_  ( .A(A[415]), .B(B[415]), .CI(
        C[415]), .S(S[415]), .CO(C[416]) );
  FA_2656 \FA_INST_0[0].FA_INST_1[416].FA_  ( .A(A[416]), .B(B[416]), .CI(
        C[416]), .S(S[416]), .CO(C[417]) );
  FA_2655 \FA_INST_0[0].FA_INST_1[417].FA_  ( .A(A[417]), .B(B[417]), .CI(
        C[417]), .S(S[417]), .CO(C[418]) );
  FA_2654 \FA_INST_0[0].FA_INST_1[418].FA_  ( .A(A[418]), .B(B[418]), .CI(
        C[418]), .S(S[418]), .CO(C[419]) );
  FA_2653 \FA_INST_0[0].FA_INST_1[419].FA_  ( .A(A[419]), .B(B[419]), .CI(
        C[419]), .S(S[419]), .CO(C[420]) );
  FA_2652 \FA_INST_0[0].FA_INST_1[420].FA_  ( .A(A[420]), .B(B[420]), .CI(
        C[420]), .S(S[420]), .CO(C[421]) );
  FA_2651 \FA_INST_0[0].FA_INST_1[421].FA_  ( .A(A[421]), .B(B[421]), .CI(
        C[421]), .S(S[421]), .CO(C[422]) );
  FA_2650 \FA_INST_0[0].FA_INST_1[422].FA_  ( .A(A[422]), .B(B[422]), .CI(
        C[422]), .S(S[422]), .CO(C[423]) );
  FA_2649 \FA_INST_0[0].FA_INST_1[423].FA_  ( .A(A[423]), .B(B[423]), .CI(
        C[423]), .S(S[423]), .CO(C[424]) );
  FA_2648 \FA_INST_0[0].FA_INST_1[424].FA_  ( .A(A[424]), .B(B[424]), .CI(
        C[424]), .S(S[424]), .CO(C[425]) );
  FA_2647 \FA_INST_0[0].FA_INST_1[425].FA_  ( .A(A[425]), .B(B[425]), .CI(
        C[425]), .S(S[425]), .CO(C[426]) );
  FA_2646 \FA_INST_0[0].FA_INST_1[426].FA_  ( .A(A[426]), .B(B[426]), .CI(
        C[426]), .S(S[426]), .CO(C[427]) );
  FA_2645 \FA_INST_0[0].FA_INST_1[427].FA_  ( .A(A[427]), .B(B[427]), .CI(
        C[427]), .S(S[427]), .CO(C[428]) );
  FA_2644 \FA_INST_0[0].FA_INST_1[428].FA_  ( .A(A[428]), .B(B[428]), .CI(
        C[428]), .S(S[428]), .CO(C[429]) );
  FA_2643 \FA_INST_0[0].FA_INST_1[429].FA_  ( .A(A[429]), .B(B[429]), .CI(
        C[429]), .S(S[429]), .CO(C[430]) );
  FA_2642 \FA_INST_0[0].FA_INST_1[430].FA_  ( .A(A[430]), .B(B[430]), .CI(
        C[430]), .S(S[430]), .CO(C[431]) );
  FA_2641 \FA_INST_0[0].FA_INST_1[431].FA_  ( .A(A[431]), .B(B[431]), .CI(
        C[431]), .S(S[431]), .CO(C[432]) );
  FA_2640 \FA_INST_0[0].FA_INST_1[432].FA_  ( .A(A[432]), .B(B[432]), .CI(
        C[432]), .S(S[432]), .CO(C[433]) );
  FA_2639 \FA_INST_0[0].FA_INST_1[433].FA_  ( .A(A[433]), .B(B[433]), .CI(
        C[433]), .S(S[433]), .CO(C[434]) );
  FA_2638 \FA_INST_0[0].FA_INST_1[434].FA_  ( .A(A[434]), .B(B[434]), .CI(
        C[434]), .S(S[434]), .CO(C[435]) );
  FA_2637 \FA_INST_0[0].FA_INST_1[435].FA_  ( .A(A[435]), .B(B[435]), .CI(
        C[435]), .S(S[435]), .CO(C[436]) );
  FA_2636 \FA_INST_0[0].FA_INST_1[436].FA_  ( .A(A[436]), .B(B[436]), .CI(
        C[436]), .S(S[436]), .CO(C[437]) );
  FA_2635 \FA_INST_0[0].FA_INST_1[437].FA_  ( .A(A[437]), .B(B[437]), .CI(
        C[437]), .S(S[437]), .CO(C[438]) );
  FA_2634 \FA_INST_0[0].FA_INST_1[438].FA_  ( .A(A[438]), .B(B[438]), .CI(
        C[438]), .S(S[438]), .CO(C[439]) );
  FA_2633 \FA_INST_0[0].FA_INST_1[439].FA_  ( .A(A[439]), .B(B[439]), .CI(
        C[439]), .S(S[439]), .CO(C[440]) );
  FA_2632 \FA_INST_0[0].FA_INST_1[440].FA_  ( .A(A[440]), .B(B[440]), .CI(
        C[440]), .S(S[440]), .CO(C[441]) );
  FA_2631 \FA_INST_0[0].FA_INST_1[441].FA_  ( .A(A[441]), .B(B[441]), .CI(
        C[441]), .S(S[441]), .CO(C[442]) );
  FA_2630 \FA_INST_0[0].FA_INST_1[442].FA_  ( .A(A[442]), .B(B[442]), .CI(
        C[442]), .S(S[442]), .CO(C[443]) );
  FA_2629 \FA_INST_0[0].FA_INST_1[443].FA_  ( .A(A[443]), .B(B[443]), .CI(
        C[443]), .S(S[443]), .CO(C[444]) );
  FA_2628 \FA_INST_0[0].FA_INST_1[444].FA_  ( .A(A[444]), .B(B[444]), .CI(
        C[444]), .S(S[444]), .CO(C[445]) );
  FA_2627 \FA_INST_0[0].FA_INST_1[445].FA_  ( .A(A[445]), .B(B[445]), .CI(
        C[445]), .S(S[445]), .CO(C[446]) );
  FA_2626 \FA_INST_0[0].FA_INST_1[446].FA_  ( .A(A[446]), .B(B[446]), .CI(
        C[446]), .S(S[446]), .CO(C[447]) );
  FA_2625 \FA_INST_0[0].FA_INST_1[447].FA_  ( .A(A[447]), .B(B[447]), .CI(
        C[447]), .S(S[447]), .CO(C[448]) );
  FA_2624 \FA_INST_0[0].FA_INST_1[448].FA_  ( .A(A[448]), .B(B[448]), .CI(
        C[448]), .S(S[448]), .CO(C[449]) );
  FA_2623 \FA_INST_0[0].FA_INST_1[449].FA_  ( .A(A[449]), .B(B[449]), .CI(
        C[449]), .S(S[449]), .CO(C[450]) );
  FA_2622 \FA_INST_0[0].FA_INST_1[450].FA_  ( .A(A[450]), .B(B[450]), .CI(
        C[450]), .S(S[450]), .CO(C[451]) );
  FA_2621 \FA_INST_0[0].FA_INST_1[451].FA_  ( .A(A[451]), .B(B[451]), .CI(
        C[451]), .S(S[451]), .CO(C[452]) );
  FA_2620 \FA_INST_0[0].FA_INST_1[452].FA_  ( .A(A[452]), .B(B[452]), .CI(
        C[452]), .S(S[452]), .CO(C[453]) );
  FA_2619 \FA_INST_0[0].FA_INST_1[453].FA_  ( .A(A[453]), .B(B[453]), .CI(
        C[453]), .S(S[453]), .CO(C[454]) );
  FA_2618 \FA_INST_0[0].FA_INST_1[454].FA_  ( .A(A[454]), .B(B[454]), .CI(
        C[454]), .S(S[454]), .CO(C[455]) );
  FA_2617 \FA_INST_0[0].FA_INST_1[455].FA_  ( .A(A[455]), .B(B[455]), .CI(
        C[455]), .S(S[455]), .CO(C[456]) );
  FA_2616 \FA_INST_0[0].FA_INST_1[456].FA_  ( .A(A[456]), .B(B[456]), .CI(
        C[456]), .S(S[456]), .CO(C[457]) );
  FA_2615 \FA_INST_0[0].FA_INST_1[457].FA_  ( .A(A[457]), .B(B[457]), .CI(
        C[457]), .S(S[457]), .CO(C[458]) );
  FA_2614 \FA_INST_0[0].FA_INST_1[458].FA_  ( .A(A[458]), .B(B[458]), .CI(
        C[458]), .S(S[458]), .CO(C[459]) );
  FA_2613 \FA_INST_0[0].FA_INST_1[459].FA_  ( .A(A[459]), .B(B[459]), .CI(
        C[459]), .S(S[459]), .CO(C[460]) );
  FA_2612 \FA_INST_0[0].FA_INST_1[460].FA_  ( .A(A[460]), .B(B[460]), .CI(
        C[460]), .S(S[460]), .CO(C[461]) );
  FA_2611 \FA_INST_0[0].FA_INST_1[461].FA_  ( .A(A[461]), .B(B[461]), .CI(
        C[461]), .S(S[461]), .CO(C[462]) );
  FA_2610 \FA_INST_0[0].FA_INST_1[462].FA_  ( .A(A[462]), .B(B[462]), .CI(
        C[462]), .S(S[462]), .CO(C[463]) );
  FA_2609 \FA_INST_0[0].FA_INST_1[463].FA_  ( .A(A[463]), .B(B[463]), .CI(
        C[463]), .S(S[463]), .CO(C[464]) );
  FA_2608 \FA_INST_0[0].FA_INST_1[464].FA_  ( .A(A[464]), .B(B[464]), .CI(
        C[464]), .S(S[464]), .CO(C[465]) );
  FA_2607 \FA_INST_0[0].FA_INST_1[465].FA_  ( .A(A[465]), .B(B[465]), .CI(
        C[465]), .S(S[465]), .CO(C[466]) );
  FA_2606 \FA_INST_0[0].FA_INST_1[466].FA_  ( .A(A[466]), .B(B[466]), .CI(
        C[466]), .S(S[466]), .CO(C[467]) );
  FA_2605 \FA_INST_0[0].FA_INST_1[467].FA_  ( .A(A[467]), .B(B[467]), .CI(
        C[467]), .S(S[467]), .CO(C[468]) );
  FA_2604 \FA_INST_0[0].FA_INST_1[468].FA_  ( .A(A[468]), .B(B[468]), .CI(
        C[468]), .S(S[468]), .CO(C[469]) );
  FA_2603 \FA_INST_0[0].FA_INST_1[469].FA_  ( .A(A[469]), .B(B[469]), .CI(
        C[469]), .S(S[469]), .CO(C[470]) );
  FA_2602 \FA_INST_0[0].FA_INST_1[470].FA_  ( .A(A[470]), .B(B[470]), .CI(
        C[470]), .S(S[470]), .CO(C[471]) );
  FA_2601 \FA_INST_0[0].FA_INST_1[471].FA_  ( .A(A[471]), .B(B[471]), .CI(
        C[471]), .S(S[471]), .CO(C[472]) );
  FA_2600 \FA_INST_0[0].FA_INST_1[472].FA_  ( .A(A[472]), .B(B[472]), .CI(
        C[472]), .S(S[472]), .CO(C[473]) );
  FA_2599 \FA_INST_0[0].FA_INST_1[473].FA_  ( .A(A[473]), .B(B[473]), .CI(
        C[473]), .S(S[473]), .CO(C[474]) );
  FA_2598 \FA_INST_0[0].FA_INST_1[474].FA_  ( .A(A[474]), .B(B[474]), .CI(
        C[474]), .S(S[474]), .CO(C[475]) );
  FA_2597 \FA_INST_0[0].FA_INST_1[475].FA_  ( .A(A[475]), .B(B[475]), .CI(
        C[475]), .S(S[475]), .CO(C[476]) );
  FA_2596 \FA_INST_0[0].FA_INST_1[476].FA_  ( .A(A[476]), .B(B[476]), .CI(
        C[476]), .S(S[476]), .CO(C[477]) );
  FA_2595 \FA_INST_0[0].FA_INST_1[477].FA_  ( .A(A[477]), .B(B[477]), .CI(
        C[477]), .S(S[477]), .CO(C[478]) );
  FA_2594 \FA_INST_0[0].FA_INST_1[478].FA_  ( .A(A[478]), .B(B[478]), .CI(
        C[478]), .S(S[478]), .CO(C[479]) );
  FA_2593 \FA_INST_0[0].FA_INST_1[479].FA_  ( .A(A[479]), .B(B[479]), .CI(
        C[479]), .S(S[479]), .CO(C[480]) );
  FA_2592 \FA_INST_0[0].FA_INST_1[480].FA_  ( .A(A[480]), .B(B[480]), .CI(
        C[480]), .S(S[480]), .CO(C[481]) );
  FA_2591 \FA_INST_0[0].FA_INST_1[481].FA_  ( .A(A[481]), .B(B[481]), .CI(
        C[481]), .S(S[481]), .CO(C[482]) );
  FA_2590 \FA_INST_0[0].FA_INST_1[482].FA_  ( .A(A[482]), .B(B[482]), .CI(
        C[482]), .S(S[482]), .CO(C[483]) );
  FA_2589 \FA_INST_0[0].FA_INST_1[483].FA_  ( .A(A[483]), .B(B[483]), .CI(
        C[483]), .S(S[483]), .CO(C[484]) );
  FA_2588 \FA_INST_0[0].FA_INST_1[484].FA_  ( .A(A[484]), .B(B[484]), .CI(
        C[484]), .S(S[484]), .CO(C[485]) );
  FA_2587 \FA_INST_0[0].FA_INST_1[485].FA_  ( .A(A[485]), .B(B[485]), .CI(
        C[485]), .S(S[485]), .CO(C[486]) );
  FA_2586 \FA_INST_0[0].FA_INST_1[486].FA_  ( .A(A[486]), .B(B[486]), .CI(
        C[486]), .S(S[486]), .CO(C[487]) );
  FA_2585 \FA_INST_0[0].FA_INST_1[487].FA_  ( .A(A[487]), .B(B[487]), .CI(
        C[487]), .S(S[487]), .CO(C[488]) );
  FA_2584 \FA_INST_0[0].FA_INST_1[488].FA_  ( .A(A[488]), .B(B[488]), .CI(
        C[488]), .S(S[488]), .CO(C[489]) );
  FA_2583 \FA_INST_0[0].FA_INST_1[489].FA_  ( .A(A[489]), .B(B[489]), .CI(
        C[489]), .S(S[489]), .CO(C[490]) );
  FA_2582 \FA_INST_0[0].FA_INST_1[490].FA_  ( .A(A[490]), .B(B[490]), .CI(
        C[490]), .S(S[490]), .CO(C[491]) );
  FA_2581 \FA_INST_0[0].FA_INST_1[491].FA_  ( .A(A[491]), .B(B[491]), .CI(
        C[491]), .S(S[491]), .CO(C[492]) );
  FA_2580 \FA_INST_0[0].FA_INST_1[492].FA_  ( .A(A[492]), .B(B[492]), .CI(
        C[492]), .S(S[492]), .CO(C[493]) );
  FA_2579 \FA_INST_0[0].FA_INST_1[493].FA_  ( .A(A[493]), .B(B[493]), .CI(
        C[493]), .S(S[493]), .CO(C[494]) );
  FA_2578 \FA_INST_0[0].FA_INST_1[494].FA_  ( .A(A[494]), .B(B[494]), .CI(
        C[494]), .S(S[494]), .CO(C[495]) );
  FA_2577 \FA_INST_0[0].FA_INST_1[495].FA_  ( .A(A[495]), .B(B[495]), .CI(
        C[495]), .S(S[495]), .CO(C[496]) );
  FA_2576 \FA_INST_0[0].FA_INST_1[496].FA_  ( .A(A[496]), .B(B[496]), .CI(
        C[496]), .S(S[496]), .CO(C[497]) );
  FA_2575 \FA_INST_0[0].FA_INST_1[497].FA_  ( .A(A[497]), .B(B[497]), .CI(
        C[497]), .S(S[497]), .CO(C[498]) );
  FA_2574 \FA_INST_0[0].FA_INST_1[498].FA_  ( .A(A[498]), .B(B[498]), .CI(
        C[498]), .S(S[498]), .CO(C[499]) );
  FA_2573 \FA_INST_0[0].FA_INST_1[499].FA_  ( .A(A[499]), .B(B[499]), .CI(
        C[499]), .S(S[499]), .CO(C[500]) );
  FA_2572 \FA_INST_0[0].FA_INST_1[500].FA_  ( .A(A[500]), .B(B[500]), .CI(
        C[500]), .S(S[500]), .CO(C[501]) );
  FA_2571 \FA_INST_0[0].FA_INST_1[501].FA_  ( .A(A[501]), .B(B[501]), .CI(
        C[501]), .S(S[501]), .CO(C[502]) );
  FA_2570 \FA_INST_0[0].FA_INST_1[502].FA_  ( .A(A[502]), .B(B[502]), .CI(
        C[502]), .S(S[502]), .CO(C[503]) );
  FA_2569 \FA_INST_0[0].FA_INST_1[503].FA_  ( .A(A[503]), .B(B[503]), .CI(
        C[503]), .S(S[503]), .CO(C[504]) );
  FA_2568 \FA_INST_0[0].FA_INST_1[504].FA_  ( .A(A[504]), .B(B[504]), .CI(
        C[504]), .S(S[504]), .CO(C[505]) );
  FA_2567 \FA_INST_0[0].FA_INST_1[505].FA_  ( .A(A[505]), .B(B[505]), .CI(
        C[505]), .S(S[505]), .CO(C[506]) );
  FA_2566 \FA_INST_0[0].FA_INST_1[506].FA_  ( .A(A[506]), .B(B[506]), .CI(
        C[506]), .S(S[506]), .CO(C[507]) );
  FA_2565 \FA_INST_0[0].FA_INST_1[507].FA_  ( .A(A[507]), .B(B[507]), .CI(
        C[507]), .S(S[507]), .CO(C[508]) );
  FA_2564 \FA_INST_0[0].FA_INST_1[508].FA_  ( .A(A[508]), .B(B[508]), .CI(
        C[508]), .S(S[508]), .CO(C[509]) );
  FA_2563 \FA_INST_0[0].FA_INST_1[509].FA_  ( .A(A[509]), .B(B[509]), .CI(
        C[509]), .S(S[509]), .CO(C[510]) );
  FA_2562 \FA_INST_0[0].FA_INST_1[510].FA_  ( .A(A[510]), .B(B[510]), .CI(
        C[510]), .S(S[510]), .CO(C[511]) );
  FA_2561 \FA_INST_0[0].FA_INST_1[511].FA_  ( .A(A[511]), .B(B[511]), .CI(
        C[511]), .S(S[511]), .CO(C[512]) );
  FA_2560 \FA_INST_0[1].FA_INST_1[0].FA_  ( .A(A[512]), .B(B[512]), .CI(C[512]), .S(S[512]), .CO(C[513]) );
  FA_2559 \FA_INST_0[1].FA_INST_1[1].FA_  ( .A(A[513]), .B(B[513]), .CI(C[513]), .S(S[513]), .CO(C[514]) );
  FA_2558 \FA_INST_0[1].FA_INST_1[2].FA_  ( .A(A[514]), .B(B[514]), .CI(C[514]), .S(S[514]), .CO(C[515]) );
  FA_2557 \FA_INST_0[1].FA_INST_1[3].FA_  ( .A(A[515]), .B(B[515]), .CI(C[515]), .S(S[515]), .CO(C[516]) );
  FA_2556 \FA_INST_0[1].FA_INST_1[4].FA_  ( .A(A[516]), .B(B[516]), .CI(C[516]), .S(S[516]), .CO(C[517]) );
  FA_2555 \FA_INST_0[1].FA_INST_1[5].FA_  ( .A(A[517]), .B(B[517]), .CI(C[517]), .S(S[517]), .CO(C[518]) );
  FA_2554 \FA_INST_0[1].FA_INST_1[6].FA_  ( .A(A[518]), .B(B[518]), .CI(C[518]), .S(S[518]), .CO(C[519]) );
  FA_2553 \FA_INST_0[1].FA_INST_1[7].FA_  ( .A(A[519]), .B(B[519]), .CI(C[519]), .S(S[519]), .CO(C[520]) );
  FA_2552 \FA_INST_0[1].FA_INST_1[8].FA_  ( .A(A[520]), .B(B[520]), .CI(C[520]), .S(S[520]), .CO(C[521]) );
  FA_2551 \FA_INST_0[1].FA_INST_1[9].FA_  ( .A(A[521]), .B(B[521]), .CI(C[521]), .S(S[521]), .CO(C[522]) );
  FA_2550 \FA_INST_0[1].FA_INST_1[10].FA_  ( .A(A[522]), .B(B[522]), .CI(
        C[522]), .S(S[522]), .CO(C[523]) );
  FA_2549 \FA_INST_0[1].FA_INST_1[11].FA_  ( .A(A[523]), .B(B[523]), .CI(
        C[523]), .S(S[523]), .CO(C[524]) );
  FA_2548 \FA_INST_0[1].FA_INST_1[12].FA_  ( .A(A[524]), .B(B[524]), .CI(
        C[524]), .S(S[524]), .CO(C[525]) );
  FA_2547 \FA_INST_0[1].FA_INST_1[13].FA_  ( .A(A[525]), .B(B[525]), .CI(
        C[525]), .S(S[525]), .CO(C[526]) );
  FA_2546 \FA_INST_0[1].FA_INST_1[14].FA_  ( .A(A[526]), .B(B[526]), .CI(
        C[526]), .S(S[526]), .CO(C[527]) );
  FA_2545 \FA_INST_0[1].FA_INST_1[15].FA_  ( .A(A[527]), .B(B[527]), .CI(
        C[527]), .S(S[527]), .CO(C[528]) );
  FA_2544 \FA_INST_0[1].FA_INST_1[16].FA_  ( .A(A[528]), .B(B[528]), .CI(
        C[528]), .S(S[528]), .CO(C[529]) );
  FA_2543 \FA_INST_0[1].FA_INST_1[17].FA_  ( .A(A[529]), .B(B[529]), .CI(
        C[529]), .S(S[529]), .CO(C[530]) );
  FA_2542 \FA_INST_0[1].FA_INST_1[18].FA_  ( .A(A[530]), .B(B[530]), .CI(
        C[530]), .S(S[530]), .CO(C[531]) );
  FA_2541 \FA_INST_0[1].FA_INST_1[19].FA_  ( .A(A[531]), .B(B[531]), .CI(
        C[531]), .S(S[531]), .CO(C[532]) );
  FA_2540 \FA_INST_0[1].FA_INST_1[20].FA_  ( .A(A[532]), .B(B[532]), .CI(
        C[532]), .S(S[532]), .CO(C[533]) );
  FA_2539 \FA_INST_0[1].FA_INST_1[21].FA_  ( .A(A[533]), .B(B[533]), .CI(
        C[533]), .S(S[533]), .CO(C[534]) );
  FA_2538 \FA_INST_0[1].FA_INST_1[22].FA_  ( .A(A[534]), .B(B[534]), .CI(
        C[534]), .S(S[534]), .CO(C[535]) );
  FA_2537 \FA_INST_0[1].FA_INST_1[23].FA_  ( .A(A[535]), .B(B[535]), .CI(
        C[535]), .S(S[535]), .CO(C[536]) );
  FA_2536 \FA_INST_0[1].FA_INST_1[24].FA_  ( .A(A[536]), .B(B[536]), .CI(
        C[536]), .S(S[536]), .CO(C[537]) );
  FA_2535 \FA_INST_0[1].FA_INST_1[25].FA_  ( .A(A[537]), .B(B[537]), .CI(
        C[537]), .S(S[537]), .CO(C[538]) );
  FA_2534 \FA_INST_0[1].FA_INST_1[26].FA_  ( .A(A[538]), .B(B[538]), .CI(
        C[538]), .S(S[538]), .CO(C[539]) );
  FA_2533 \FA_INST_0[1].FA_INST_1[27].FA_  ( .A(A[539]), .B(B[539]), .CI(
        C[539]), .S(S[539]), .CO(C[540]) );
  FA_2532 \FA_INST_0[1].FA_INST_1[28].FA_  ( .A(A[540]), .B(B[540]), .CI(
        C[540]), .S(S[540]), .CO(C[541]) );
  FA_2531 \FA_INST_0[1].FA_INST_1[29].FA_  ( .A(A[541]), .B(B[541]), .CI(
        C[541]), .S(S[541]), .CO(C[542]) );
  FA_2530 \FA_INST_0[1].FA_INST_1[30].FA_  ( .A(A[542]), .B(B[542]), .CI(
        C[542]), .S(S[542]), .CO(C[543]) );
  FA_2529 \FA_INST_0[1].FA_INST_1[31].FA_  ( .A(A[543]), .B(B[543]), .CI(
        C[543]), .S(S[543]), .CO(C[544]) );
  FA_2528 \FA_INST_0[1].FA_INST_1[32].FA_  ( .A(A[544]), .B(B[544]), .CI(
        C[544]), .S(S[544]), .CO(C[545]) );
  FA_2527 \FA_INST_0[1].FA_INST_1[33].FA_  ( .A(A[545]), .B(B[545]), .CI(
        C[545]), .S(S[545]), .CO(C[546]) );
  FA_2526 \FA_INST_0[1].FA_INST_1[34].FA_  ( .A(A[546]), .B(B[546]), .CI(
        C[546]), .S(S[546]), .CO(C[547]) );
  FA_2525 \FA_INST_0[1].FA_INST_1[35].FA_  ( .A(A[547]), .B(B[547]), .CI(
        C[547]), .S(S[547]), .CO(C[548]) );
  FA_2524 \FA_INST_0[1].FA_INST_1[36].FA_  ( .A(A[548]), .B(B[548]), .CI(
        C[548]), .S(S[548]), .CO(C[549]) );
  FA_2523 \FA_INST_0[1].FA_INST_1[37].FA_  ( .A(A[549]), .B(B[549]), .CI(
        C[549]), .S(S[549]), .CO(C[550]) );
  FA_2522 \FA_INST_0[1].FA_INST_1[38].FA_  ( .A(A[550]), .B(B[550]), .CI(
        C[550]), .S(S[550]), .CO(C[551]) );
  FA_2521 \FA_INST_0[1].FA_INST_1[39].FA_  ( .A(A[551]), .B(B[551]), .CI(
        C[551]), .S(S[551]), .CO(C[552]) );
  FA_2520 \FA_INST_0[1].FA_INST_1[40].FA_  ( .A(A[552]), .B(B[552]), .CI(
        C[552]), .S(S[552]), .CO(C[553]) );
  FA_2519 \FA_INST_0[1].FA_INST_1[41].FA_  ( .A(A[553]), .B(B[553]), .CI(
        C[553]), .S(S[553]), .CO(C[554]) );
  FA_2518 \FA_INST_0[1].FA_INST_1[42].FA_  ( .A(A[554]), .B(B[554]), .CI(
        C[554]), .S(S[554]), .CO(C[555]) );
  FA_2517 \FA_INST_0[1].FA_INST_1[43].FA_  ( .A(A[555]), .B(B[555]), .CI(
        C[555]), .S(S[555]), .CO(C[556]) );
  FA_2516 \FA_INST_0[1].FA_INST_1[44].FA_  ( .A(A[556]), .B(B[556]), .CI(
        C[556]), .S(S[556]), .CO(C[557]) );
  FA_2515 \FA_INST_0[1].FA_INST_1[45].FA_  ( .A(A[557]), .B(B[557]), .CI(
        C[557]), .S(S[557]), .CO(C[558]) );
  FA_2514 \FA_INST_0[1].FA_INST_1[46].FA_  ( .A(A[558]), .B(B[558]), .CI(
        C[558]), .S(S[558]), .CO(C[559]) );
  FA_2513 \FA_INST_0[1].FA_INST_1[47].FA_  ( .A(A[559]), .B(B[559]), .CI(
        C[559]), .S(S[559]), .CO(C[560]) );
  FA_2512 \FA_INST_0[1].FA_INST_1[48].FA_  ( .A(A[560]), .B(B[560]), .CI(
        C[560]), .S(S[560]), .CO(C[561]) );
  FA_2511 \FA_INST_0[1].FA_INST_1[49].FA_  ( .A(A[561]), .B(B[561]), .CI(
        C[561]), .S(S[561]), .CO(C[562]) );
  FA_2510 \FA_INST_0[1].FA_INST_1[50].FA_  ( .A(A[562]), .B(B[562]), .CI(
        C[562]), .S(S[562]), .CO(C[563]) );
  FA_2509 \FA_INST_0[1].FA_INST_1[51].FA_  ( .A(A[563]), .B(B[563]), .CI(
        C[563]), .S(S[563]), .CO(C[564]) );
  FA_2508 \FA_INST_0[1].FA_INST_1[52].FA_  ( .A(A[564]), .B(B[564]), .CI(
        C[564]), .S(S[564]), .CO(C[565]) );
  FA_2507 \FA_INST_0[1].FA_INST_1[53].FA_  ( .A(A[565]), .B(B[565]), .CI(
        C[565]), .S(S[565]), .CO(C[566]) );
  FA_2506 \FA_INST_0[1].FA_INST_1[54].FA_  ( .A(A[566]), .B(B[566]), .CI(
        C[566]), .S(S[566]), .CO(C[567]) );
  FA_2505 \FA_INST_0[1].FA_INST_1[55].FA_  ( .A(A[567]), .B(B[567]), .CI(
        C[567]), .S(S[567]), .CO(C[568]) );
  FA_2504 \FA_INST_0[1].FA_INST_1[56].FA_  ( .A(A[568]), .B(B[568]), .CI(
        C[568]), .S(S[568]), .CO(C[569]) );
  FA_2503 \FA_INST_0[1].FA_INST_1[57].FA_  ( .A(A[569]), .B(B[569]), .CI(
        C[569]), .S(S[569]), .CO(C[570]) );
  FA_2502 \FA_INST_0[1].FA_INST_1[58].FA_  ( .A(A[570]), .B(B[570]), .CI(
        C[570]), .S(S[570]), .CO(C[571]) );
  FA_2501 \FA_INST_0[1].FA_INST_1[59].FA_  ( .A(A[571]), .B(B[571]), .CI(
        C[571]), .S(S[571]), .CO(C[572]) );
  FA_2500 \FA_INST_0[1].FA_INST_1[60].FA_  ( .A(A[572]), .B(B[572]), .CI(
        C[572]), .S(S[572]), .CO(C[573]) );
  FA_2499 \FA_INST_0[1].FA_INST_1[61].FA_  ( .A(A[573]), .B(B[573]), .CI(
        C[573]), .S(S[573]), .CO(C[574]) );
  FA_2498 \FA_INST_0[1].FA_INST_1[62].FA_  ( .A(A[574]), .B(B[574]), .CI(
        C[574]), .S(S[574]), .CO(C[575]) );
  FA_2497 \FA_INST_0[1].FA_INST_1[63].FA_  ( .A(A[575]), .B(B[575]), .CI(
        C[575]), .S(S[575]), .CO(C[576]) );
  FA_2496 \FA_INST_0[1].FA_INST_1[64].FA_  ( .A(A[576]), .B(B[576]), .CI(
        C[576]), .S(S[576]), .CO(C[577]) );
  FA_2495 \FA_INST_0[1].FA_INST_1[65].FA_  ( .A(A[577]), .B(B[577]), .CI(
        C[577]), .S(S[577]), .CO(C[578]) );
  FA_2494 \FA_INST_0[1].FA_INST_1[66].FA_  ( .A(A[578]), .B(B[578]), .CI(
        C[578]), .S(S[578]), .CO(C[579]) );
  FA_2493 \FA_INST_0[1].FA_INST_1[67].FA_  ( .A(A[579]), .B(B[579]), .CI(
        C[579]), .S(S[579]), .CO(C[580]) );
  FA_2492 \FA_INST_0[1].FA_INST_1[68].FA_  ( .A(A[580]), .B(B[580]), .CI(
        C[580]), .S(S[580]), .CO(C[581]) );
  FA_2491 \FA_INST_0[1].FA_INST_1[69].FA_  ( .A(A[581]), .B(B[581]), .CI(
        C[581]), .S(S[581]), .CO(C[582]) );
  FA_2490 \FA_INST_0[1].FA_INST_1[70].FA_  ( .A(A[582]), .B(B[582]), .CI(
        C[582]), .S(S[582]), .CO(C[583]) );
  FA_2489 \FA_INST_0[1].FA_INST_1[71].FA_  ( .A(A[583]), .B(B[583]), .CI(
        C[583]), .S(S[583]), .CO(C[584]) );
  FA_2488 \FA_INST_0[1].FA_INST_1[72].FA_  ( .A(A[584]), .B(B[584]), .CI(
        C[584]), .S(S[584]), .CO(C[585]) );
  FA_2487 \FA_INST_0[1].FA_INST_1[73].FA_  ( .A(A[585]), .B(B[585]), .CI(
        C[585]), .S(S[585]), .CO(C[586]) );
  FA_2486 \FA_INST_0[1].FA_INST_1[74].FA_  ( .A(A[586]), .B(B[586]), .CI(
        C[586]), .S(S[586]), .CO(C[587]) );
  FA_2485 \FA_INST_0[1].FA_INST_1[75].FA_  ( .A(A[587]), .B(B[587]), .CI(
        C[587]), .S(S[587]), .CO(C[588]) );
  FA_2484 \FA_INST_0[1].FA_INST_1[76].FA_  ( .A(A[588]), .B(B[588]), .CI(
        C[588]), .S(S[588]), .CO(C[589]) );
  FA_2483 \FA_INST_0[1].FA_INST_1[77].FA_  ( .A(A[589]), .B(B[589]), .CI(
        C[589]), .S(S[589]), .CO(C[590]) );
  FA_2482 \FA_INST_0[1].FA_INST_1[78].FA_  ( .A(A[590]), .B(B[590]), .CI(
        C[590]), .S(S[590]), .CO(C[591]) );
  FA_2481 \FA_INST_0[1].FA_INST_1[79].FA_  ( .A(A[591]), .B(B[591]), .CI(
        C[591]), .S(S[591]), .CO(C[592]) );
  FA_2480 \FA_INST_0[1].FA_INST_1[80].FA_  ( .A(A[592]), .B(B[592]), .CI(
        C[592]), .S(S[592]), .CO(C[593]) );
  FA_2479 \FA_INST_0[1].FA_INST_1[81].FA_  ( .A(A[593]), .B(B[593]), .CI(
        C[593]), .S(S[593]), .CO(C[594]) );
  FA_2478 \FA_INST_0[1].FA_INST_1[82].FA_  ( .A(A[594]), .B(B[594]), .CI(
        C[594]), .S(S[594]), .CO(C[595]) );
  FA_2477 \FA_INST_0[1].FA_INST_1[83].FA_  ( .A(A[595]), .B(B[595]), .CI(
        C[595]), .S(S[595]), .CO(C[596]) );
  FA_2476 \FA_INST_0[1].FA_INST_1[84].FA_  ( .A(A[596]), .B(B[596]), .CI(
        C[596]), .S(S[596]), .CO(C[597]) );
  FA_2475 \FA_INST_0[1].FA_INST_1[85].FA_  ( .A(A[597]), .B(B[597]), .CI(
        C[597]), .S(S[597]), .CO(C[598]) );
  FA_2474 \FA_INST_0[1].FA_INST_1[86].FA_  ( .A(A[598]), .B(B[598]), .CI(
        C[598]), .S(S[598]), .CO(C[599]) );
  FA_2473 \FA_INST_0[1].FA_INST_1[87].FA_  ( .A(A[599]), .B(B[599]), .CI(
        C[599]), .S(S[599]), .CO(C[600]) );
  FA_2472 \FA_INST_0[1].FA_INST_1[88].FA_  ( .A(A[600]), .B(B[600]), .CI(
        C[600]), .S(S[600]), .CO(C[601]) );
  FA_2471 \FA_INST_0[1].FA_INST_1[89].FA_  ( .A(A[601]), .B(B[601]), .CI(
        C[601]), .S(S[601]), .CO(C[602]) );
  FA_2470 \FA_INST_0[1].FA_INST_1[90].FA_  ( .A(A[602]), .B(B[602]), .CI(
        C[602]), .S(S[602]), .CO(C[603]) );
  FA_2469 \FA_INST_0[1].FA_INST_1[91].FA_  ( .A(A[603]), .B(B[603]), .CI(
        C[603]), .S(S[603]), .CO(C[604]) );
  FA_2468 \FA_INST_0[1].FA_INST_1[92].FA_  ( .A(A[604]), .B(B[604]), .CI(
        C[604]), .S(S[604]), .CO(C[605]) );
  FA_2467 \FA_INST_0[1].FA_INST_1[93].FA_  ( .A(A[605]), .B(B[605]), .CI(
        C[605]), .S(S[605]), .CO(C[606]) );
  FA_2466 \FA_INST_0[1].FA_INST_1[94].FA_  ( .A(A[606]), .B(B[606]), .CI(
        C[606]), .S(S[606]), .CO(C[607]) );
  FA_2465 \FA_INST_0[1].FA_INST_1[95].FA_  ( .A(A[607]), .B(B[607]), .CI(
        C[607]), .S(S[607]), .CO(C[608]) );
  FA_2464 \FA_INST_0[1].FA_INST_1[96].FA_  ( .A(A[608]), .B(B[608]), .CI(
        C[608]), .S(S[608]), .CO(C[609]) );
  FA_2463 \FA_INST_0[1].FA_INST_1[97].FA_  ( .A(A[609]), .B(B[609]), .CI(
        C[609]), .S(S[609]), .CO(C[610]) );
  FA_2462 \FA_INST_0[1].FA_INST_1[98].FA_  ( .A(A[610]), .B(B[610]), .CI(
        C[610]), .S(S[610]), .CO(C[611]) );
  FA_2461 \FA_INST_0[1].FA_INST_1[99].FA_  ( .A(A[611]), .B(B[611]), .CI(
        C[611]), .S(S[611]), .CO(C[612]) );
  FA_2460 \FA_INST_0[1].FA_INST_1[100].FA_  ( .A(A[612]), .B(B[612]), .CI(
        C[612]), .S(S[612]), .CO(C[613]) );
  FA_2459 \FA_INST_0[1].FA_INST_1[101].FA_  ( .A(A[613]), .B(B[613]), .CI(
        C[613]), .S(S[613]), .CO(C[614]) );
  FA_2458 \FA_INST_0[1].FA_INST_1[102].FA_  ( .A(A[614]), .B(B[614]), .CI(
        C[614]), .S(S[614]), .CO(C[615]) );
  FA_2457 \FA_INST_0[1].FA_INST_1[103].FA_  ( .A(A[615]), .B(B[615]), .CI(
        C[615]), .S(S[615]), .CO(C[616]) );
  FA_2456 \FA_INST_0[1].FA_INST_1[104].FA_  ( .A(A[616]), .B(B[616]), .CI(
        C[616]), .S(S[616]), .CO(C[617]) );
  FA_2455 \FA_INST_0[1].FA_INST_1[105].FA_  ( .A(A[617]), .B(B[617]), .CI(
        C[617]), .S(S[617]), .CO(C[618]) );
  FA_2454 \FA_INST_0[1].FA_INST_1[106].FA_  ( .A(A[618]), .B(B[618]), .CI(
        C[618]), .S(S[618]), .CO(C[619]) );
  FA_2453 \FA_INST_0[1].FA_INST_1[107].FA_  ( .A(A[619]), .B(B[619]), .CI(
        C[619]), .S(S[619]), .CO(C[620]) );
  FA_2452 \FA_INST_0[1].FA_INST_1[108].FA_  ( .A(A[620]), .B(B[620]), .CI(
        C[620]), .S(S[620]), .CO(C[621]) );
  FA_2451 \FA_INST_0[1].FA_INST_1[109].FA_  ( .A(A[621]), .B(B[621]), .CI(
        C[621]), .S(S[621]), .CO(C[622]) );
  FA_2450 \FA_INST_0[1].FA_INST_1[110].FA_  ( .A(A[622]), .B(B[622]), .CI(
        C[622]), .S(S[622]), .CO(C[623]) );
  FA_2449 \FA_INST_0[1].FA_INST_1[111].FA_  ( .A(A[623]), .B(B[623]), .CI(
        C[623]), .S(S[623]), .CO(C[624]) );
  FA_2448 \FA_INST_0[1].FA_INST_1[112].FA_  ( .A(A[624]), .B(B[624]), .CI(
        C[624]), .S(S[624]), .CO(C[625]) );
  FA_2447 \FA_INST_0[1].FA_INST_1[113].FA_  ( .A(A[625]), .B(B[625]), .CI(
        C[625]), .S(S[625]), .CO(C[626]) );
  FA_2446 \FA_INST_0[1].FA_INST_1[114].FA_  ( .A(A[626]), .B(B[626]), .CI(
        C[626]), .S(S[626]), .CO(C[627]) );
  FA_2445 \FA_INST_0[1].FA_INST_1[115].FA_  ( .A(A[627]), .B(B[627]), .CI(
        C[627]), .S(S[627]), .CO(C[628]) );
  FA_2444 \FA_INST_0[1].FA_INST_1[116].FA_  ( .A(A[628]), .B(B[628]), .CI(
        C[628]), .S(S[628]), .CO(C[629]) );
  FA_2443 \FA_INST_0[1].FA_INST_1[117].FA_  ( .A(A[629]), .B(B[629]), .CI(
        C[629]), .S(S[629]), .CO(C[630]) );
  FA_2442 \FA_INST_0[1].FA_INST_1[118].FA_  ( .A(A[630]), .B(B[630]), .CI(
        C[630]), .S(S[630]), .CO(C[631]) );
  FA_2441 \FA_INST_0[1].FA_INST_1[119].FA_  ( .A(A[631]), .B(B[631]), .CI(
        C[631]), .S(S[631]), .CO(C[632]) );
  FA_2440 \FA_INST_0[1].FA_INST_1[120].FA_  ( .A(A[632]), .B(B[632]), .CI(
        C[632]), .S(S[632]), .CO(C[633]) );
  FA_2439 \FA_INST_0[1].FA_INST_1[121].FA_  ( .A(A[633]), .B(B[633]), .CI(
        C[633]), .S(S[633]), .CO(C[634]) );
  FA_2438 \FA_INST_0[1].FA_INST_1[122].FA_  ( .A(A[634]), .B(B[634]), .CI(
        C[634]), .S(S[634]), .CO(C[635]) );
  FA_2437 \FA_INST_0[1].FA_INST_1[123].FA_  ( .A(A[635]), .B(B[635]), .CI(
        C[635]), .S(S[635]), .CO(C[636]) );
  FA_2436 \FA_INST_0[1].FA_INST_1[124].FA_  ( .A(A[636]), .B(B[636]), .CI(
        C[636]), .S(S[636]), .CO(C[637]) );
  FA_2435 \FA_INST_0[1].FA_INST_1[125].FA_  ( .A(A[637]), .B(B[637]), .CI(
        C[637]), .S(S[637]), .CO(C[638]) );
  FA_2434 \FA_INST_0[1].FA_INST_1[126].FA_  ( .A(A[638]), .B(B[638]), .CI(
        C[638]), .S(S[638]), .CO(C[639]) );
  FA_2433 \FA_INST_0[1].FA_INST_1[127].FA_  ( .A(A[639]), .B(B[639]), .CI(
        C[639]), .S(S[639]), .CO(C[640]) );
  FA_2432 \FA_INST_0[1].FA_INST_1[128].FA_  ( .A(A[640]), .B(B[640]), .CI(
        C[640]), .S(S[640]), .CO(C[641]) );
  FA_2431 \FA_INST_0[1].FA_INST_1[129].FA_  ( .A(A[641]), .B(B[641]), .CI(
        C[641]), .S(S[641]), .CO(C[642]) );
  FA_2430 \FA_INST_0[1].FA_INST_1[130].FA_  ( .A(A[642]), .B(B[642]), .CI(
        C[642]), .S(S[642]), .CO(C[643]) );
  FA_2429 \FA_INST_0[1].FA_INST_1[131].FA_  ( .A(A[643]), .B(B[643]), .CI(
        C[643]), .S(S[643]), .CO(C[644]) );
  FA_2428 \FA_INST_0[1].FA_INST_1[132].FA_  ( .A(A[644]), .B(B[644]), .CI(
        C[644]), .S(S[644]), .CO(C[645]) );
  FA_2427 \FA_INST_0[1].FA_INST_1[133].FA_  ( .A(A[645]), .B(B[645]), .CI(
        C[645]), .S(S[645]), .CO(C[646]) );
  FA_2426 \FA_INST_0[1].FA_INST_1[134].FA_  ( .A(A[646]), .B(B[646]), .CI(
        C[646]), .S(S[646]), .CO(C[647]) );
  FA_2425 \FA_INST_0[1].FA_INST_1[135].FA_  ( .A(A[647]), .B(B[647]), .CI(
        C[647]), .S(S[647]), .CO(C[648]) );
  FA_2424 \FA_INST_0[1].FA_INST_1[136].FA_  ( .A(A[648]), .B(B[648]), .CI(
        C[648]), .S(S[648]), .CO(C[649]) );
  FA_2423 \FA_INST_0[1].FA_INST_1[137].FA_  ( .A(A[649]), .B(B[649]), .CI(
        C[649]), .S(S[649]), .CO(C[650]) );
  FA_2422 \FA_INST_0[1].FA_INST_1[138].FA_  ( .A(A[650]), .B(B[650]), .CI(
        C[650]), .S(S[650]), .CO(C[651]) );
  FA_2421 \FA_INST_0[1].FA_INST_1[139].FA_  ( .A(A[651]), .B(B[651]), .CI(
        C[651]), .S(S[651]), .CO(C[652]) );
  FA_2420 \FA_INST_0[1].FA_INST_1[140].FA_  ( .A(A[652]), .B(B[652]), .CI(
        C[652]), .S(S[652]), .CO(C[653]) );
  FA_2419 \FA_INST_0[1].FA_INST_1[141].FA_  ( .A(A[653]), .B(B[653]), .CI(
        C[653]), .S(S[653]), .CO(C[654]) );
  FA_2418 \FA_INST_0[1].FA_INST_1[142].FA_  ( .A(A[654]), .B(B[654]), .CI(
        C[654]), .S(S[654]), .CO(C[655]) );
  FA_2417 \FA_INST_0[1].FA_INST_1[143].FA_  ( .A(A[655]), .B(B[655]), .CI(
        C[655]), .S(S[655]), .CO(C[656]) );
  FA_2416 \FA_INST_0[1].FA_INST_1[144].FA_  ( .A(A[656]), .B(B[656]), .CI(
        C[656]), .S(S[656]), .CO(C[657]) );
  FA_2415 \FA_INST_0[1].FA_INST_1[145].FA_  ( .A(A[657]), .B(B[657]), .CI(
        C[657]), .S(S[657]), .CO(C[658]) );
  FA_2414 \FA_INST_0[1].FA_INST_1[146].FA_  ( .A(A[658]), .B(B[658]), .CI(
        C[658]), .S(S[658]), .CO(C[659]) );
  FA_2413 \FA_INST_0[1].FA_INST_1[147].FA_  ( .A(A[659]), .B(B[659]), .CI(
        C[659]), .S(S[659]), .CO(C[660]) );
  FA_2412 \FA_INST_0[1].FA_INST_1[148].FA_  ( .A(A[660]), .B(B[660]), .CI(
        C[660]), .S(S[660]), .CO(C[661]) );
  FA_2411 \FA_INST_0[1].FA_INST_1[149].FA_  ( .A(A[661]), .B(B[661]), .CI(
        C[661]), .S(S[661]), .CO(C[662]) );
  FA_2410 \FA_INST_0[1].FA_INST_1[150].FA_  ( .A(A[662]), .B(B[662]), .CI(
        C[662]), .S(S[662]), .CO(C[663]) );
  FA_2409 \FA_INST_0[1].FA_INST_1[151].FA_  ( .A(A[663]), .B(B[663]), .CI(
        C[663]), .S(S[663]), .CO(C[664]) );
  FA_2408 \FA_INST_0[1].FA_INST_1[152].FA_  ( .A(A[664]), .B(B[664]), .CI(
        C[664]), .S(S[664]), .CO(C[665]) );
  FA_2407 \FA_INST_0[1].FA_INST_1[153].FA_  ( .A(A[665]), .B(B[665]), .CI(
        C[665]), .S(S[665]), .CO(C[666]) );
  FA_2406 \FA_INST_0[1].FA_INST_1[154].FA_  ( .A(A[666]), .B(B[666]), .CI(
        C[666]), .S(S[666]), .CO(C[667]) );
  FA_2405 \FA_INST_0[1].FA_INST_1[155].FA_  ( .A(A[667]), .B(B[667]), .CI(
        C[667]), .S(S[667]), .CO(C[668]) );
  FA_2404 \FA_INST_0[1].FA_INST_1[156].FA_  ( .A(A[668]), .B(B[668]), .CI(
        C[668]), .S(S[668]), .CO(C[669]) );
  FA_2403 \FA_INST_0[1].FA_INST_1[157].FA_  ( .A(A[669]), .B(B[669]), .CI(
        C[669]), .S(S[669]), .CO(C[670]) );
  FA_2402 \FA_INST_0[1].FA_INST_1[158].FA_  ( .A(A[670]), .B(B[670]), .CI(
        C[670]), .S(S[670]), .CO(C[671]) );
  FA_2401 \FA_INST_0[1].FA_INST_1[159].FA_  ( .A(A[671]), .B(B[671]), .CI(
        C[671]), .S(S[671]), .CO(C[672]) );
  FA_2400 \FA_INST_0[1].FA_INST_1[160].FA_  ( .A(A[672]), .B(B[672]), .CI(
        C[672]), .S(S[672]), .CO(C[673]) );
  FA_2399 \FA_INST_0[1].FA_INST_1[161].FA_  ( .A(A[673]), .B(B[673]), .CI(
        C[673]), .S(S[673]), .CO(C[674]) );
  FA_2398 \FA_INST_0[1].FA_INST_1[162].FA_  ( .A(A[674]), .B(B[674]), .CI(
        C[674]), .S(S[674]), .CO(C[675]) );
  FA_2397 \FA_INST_0[1].FA_INST_1[163].FA_  ( .A(A[675]), .B(B[675]), .CI(
        C[675]), .S(S[675]), .CO(C[676]) );
  FA_2396 \FA_INST_0[1].FA_INST_1[164].FA_  ( .A(A[676]), .B(B[676]), .CI(
        C[676]), .S(S[676]), .CO(C[677]) );
  FA_2395 \FA_INST_0[1].FA_INST_1[165].FA_  ( .A(A[677]), .B(B[677]), .CI(
        C[677]), .S(S[677]), .CO(C[678]) );
  FA_2394 \FA_INST_0[1].FA_INST_1[166].FA_  ( .A(A[678]), .B(B[678]), .CI(
        C[678]), .S(S[678]), .CO(C[679]) );
  FA_2393 \FA_INST_0[1].FA_INST_1[167].FA_  ( .A(A[679]), .B(B[679]), .CI(
        C[679]), .S(S[679]), .CO(C[680]) );
  FA_2392 \FA_INST_0[1].FA_INST_1[168].FA_  ( .A(A[680]), .B(B[680]), .CI(
        C[680]), .S(S[680]), .CO(C[681]) );
  FA_2391 \FA_INST_0[1].FA_INST_1[169].FA_  ( .A(A[681]), .B(B[681]), .CI(
        C[681]), .S(S[681]), .CO(C[682]) );
  FA_2390 \FA_INST_0[1].FA_INST_1[170].FA_  ( .A(A[682]), .B(B[682]), .CI(
        C[682]), .S(S[682]), .CO(C[683]) );
  FA_2389 \FA_INST_0[1].FA_INST_1[171].FA_  ( .A(A[683]), .B(B[683]), .CI(
        C[683]), .S(S[683]), .CO(C[684]) );
  FA_2388 \FA_INST_0[1].FA_INST_1[172].FA_  ( .A(A[684]), .B(B[684]), .CI(
        C[684]), .S(S[684]), .CO(C[685]) );
  FA_2387 \FA_INST_0[1].FA_INST_1[173].FA_  ( .A(A[685]), .B(B[685]), .CI(
        C[685]), .S(S[685]), .CO(C[686]) );
  FA_2386 \FA_INST_0[1].FA_INST_1[174].FA_  ( .A(A[686]), .B(B[686]), .CI(
        C[686]), .S(S[686]), .CO(C[687]) );
  FA_2385 \FA_INST_0[1].FA_INST_1[175].FA_  ( .A(A[687]), .B(B[687]), .CI(
        C[687]), .S(S[687]), .CO(C[688]) );
  FA_2384 \FA_INST_0[1].FA_INST_1[176].FA_  ( .A(A[688]), .B(B[688]), .CI(
        C[688]), .S(S[688]), .CO(C[689]) );
  FA_2383 \FA_INST_0[1].FA_INST_1[177].FA_  ( .A(A[689]), .B(B[689]), .CI(
        C[689]), .S(S[689]), .CO(C[690]) );
  FA_2382 \FA_INST_0[1].FA_INST_1[178].FA_  ( .A(A[690]), .B(B[690]), .CI(
        C[690]), .S(S[690]), .CO(C[691]) );
  FA_2381 \FA_INST_0[1].FA_INST_1[179].FA_  ( .A(A[691]), .B(B[691]), .CI(
        C[691]), .S(S[691]), .CO(C[692]) );
  FA_2380 \FA_INST_0[1].FA_INST_1[180].FA_  ( .A(A[692]), .B(B[692]), .CI(
        C[692]), .S(S[692]), .CO(C[693]) );
  FA_2379 \FA_INST_0[1].FA_INST_1[181].FA_  ( .A(A[693]), .B(B[693]), .CI(
        C[693]), .S(S[693]), .CO(C[694]) );
  FA_2378 \FA_INST_0[1].FA_INST_1[182].FA_  ( .A(A[694]), .B(B[694]), .CI(
        C[694]), .S(S[694]), .CO(C[695]) );
  FA_2377 \FA_INST_0[1].FA_INST_1[183].FA_  ( .A(A[695]), .B(B[695]), .CI(
        C[695]), .S(S[695]), .CO(C[696]) );
  FA_2376 \FA_INST_0[1].FA_INST_1[184].FA_  ( .A(A[696]), .B(B[696]), .CI(
        C[696]), .S(S[696]), .CO(C[697]) );
  FA_2375 \FA_INST_0[1].FA_INST_1[185].FA_  ( .A(A[697]), .B(B[697]), .CI(
        C[697]), .S(S[697]), .CO(C[698]) );
  FA_2374 \FA_INST_0[1].FA_INST_1[186].FA_  ( .A(A[698]), .B(B[698]), .CI(
        C[698]), .S(S[698]), .CO(C[699]) );
  FA_2373 \FA_INST_0[1].FA_INST_1[187].FA_  ( .A(A[699]), .B(B[699]), .CI(
        C[699]), .S(S[699]), .CO(C[700]) );
  FA_2372 \FA_INST_0[1].FA_INST_1[188].FA_  ( .A(A[700]), .B(B[700]), .CI(
        C[700]), .S(S[700]), .CO(C[701]) );
  FA_2371 \FA_INST_0[1].FA_INST_1[189].FA_  ( .A(A[701]), .B(B[701]), .CI(
        C[701]), .S(S[701]), .CO(C[702]) );
  FA_2370 \FA_INST_0[1].FA_INST_1[190].FA_  ( .A(A[702]), .B(B[702]), .CI(
        C[702]), .S(S[702]), .CO(C[703]) );
  FA_2369 \FA_INST_0[1].FA_INST_1[191].FA_  ( .A(A[703]), .B(B[703]), .CI(
        C[703]), .S(S[703]), .CO(C[704]) );
  FA_2368 \FA_INST_0[1].FA_INST_1[192].FA_  ( .A(A[704]), .B(B[704]), .CI(
        C[704]), .S(S[704]), .CO(C[705]) );
  FA_2367 \FA_INST_0[1].FA_INST_1[193].FA_  ( .A(A[705]), .B(B[705]), .CI(
        C[705]), .S(S[705]), .CO(C[706]) );
  FA_2366 \FA_INST_0[1].FA_INST_1[194].FA_  ( .A(A[706]), .B(B[706]), .CI(
        C[706]), .S(S[706]), .CO(C[707]) );
  FA_2365 \FA_INST_0[1].FA_INST_1[195].FA_  ( .A(A[707]), .B(B[707]), .CI(
        C[707]), .S(S[707]), .CO(C[708]) );
  FA_2364 \FA_INST_0[1].FA_INST_1[196].FA_  ( .A(A[708]), .B(B[708]), .CI(
        C[708]), .S(S[708]), .CO(C[709]) );
  FA_2363 \FA_INST_0[1].FA_INST_1[197].FA_  ( .A(A[709]), .B(B[709]), .CI(
        C[709]), .S(S[709]), .CO(C[710]) );
  FA_2362 \FA_INST_0[1].FA_INST_1[198].FA_  ( .A(A[710]), .B(B[710]), .CI(
        C[710]), .S(S[710]), .CO(C[711]) );
  FA_2361 \FA_INST_0[1].FA_INST_1[199].FA_  ( .A(A[711]), .B(B[711]), .CI(
        C[711]), .S(S[711]), .CO(C[712]) );
  FA_2360 \FA_INST_0[1].FA_INST_1[200].FA_  ( .A(A[712]), .B(B[712]), .CI(
        C[712]), .S(S[712]), .CO(C[713]) );
  FA_2359 \FA_INST_0[1].FA_INST_1[201].FA_  ( .A(A[713]), .B(B[713]), .CI(
        C[713]), .S(S[713]), .CO(C[714]) );
  FA_2358 \FA_INST_0[1].FA_INST_1[202].FA_  ( .A(A[714]), .B(B[714]), .CI(
        C[714]), .S(S[714]), .CO(C[715]) );
  FA_2357 \FA_INST_0[1].FA_INST_1[203].FA_  ( .A(A[715]), .B(B[715]), .CI(
        C[715]), .S(S[715]), .CO(C[716]) );
  FA_2356 \FA_INST_0[1].FA_INST_1[204].FA_  ( .A(A[716]), .B(B[716]), .CI(
        C[716]), .S(S[716]), .CO(C[717]) );
  FA_2355 \FA_INST_0[1].FA_INST_1[205].FA_  ( .A(A[717]), .B(B[717]), .CI(
        C[717]), .S(S[717]), .CO(C[718]) );
  FA_2354 \FA_INST_0[1].FA_INST_1[206].FA_  ( .A(A[718]), .B(B[718]), .CI(
        C[718]), .S(S[718]), .CO(C[719]) );
  FA_2353 \FA_INST_0[1].FA_INST_1[207].FA_  ( .A(A[719]), .B(B[719]), .CI(
        C[719]), .S(S[719]), .CO(C[720]) );
  FA_2352 \FA_INST_0[1].FA_INST_1[208].FA_  ( .A(A[720]), .B(B[720]), .CI(
        C[720]), .S(S[720]), .CO(C[721]) );
  FA_2351 \FA_INST_0[1].FA_INST_1[209].FA_  ( .A(A[721]), .B(B[721]), .CI(
        C[721]), .S(S[721]), .CO(C[722]) );
  FA_2350 \FA_INST_0[1].FA_INST_1[210].FA_  ( .A(A[722]), .B(B[722]), .CI(
        C[722]), .S(S[722]), .CO(C[723]) );
  FA_2349 \FA_INST_0[1].FA_INST_1[211].FA_  ( .A(A[723]), .B(B[723]), .CI(
        C[723]), .S(S[723]), .CO(C[724]) );
  FA_2348 \FA_INST_0[1].FA_INST_1[212].FA_  ( .A(A[724]), .B(B[724]), .CI(
        C[724]), .S(S[724]), .CO(C[725]) );
  FA_2347 \FA_INST_0[1].FA_INST_1[213].FA_  ( .A(A[725]), .B(B[725]), .CI(
        C[725]), .S(S[725]), .CO(C[726]) );
  FA_2346 \FA_INST_0[1].FA_INST_1[214].FA_  ( .A(A[726]), .B(B[726]), .CI(
        C[726]), .S(S[726]), .CO(C[727]) );
  FA_2345 \FA_INST_0[1].FA_INST_1[215].FA_  ( .A(A[727]), .B(B[727]), .CI(
        C[727]), .S(S[727]), .CO(C[728]) );
  FA_2344 \FA_INST_0[1].FA_INST_1[216].FA_  ( .A(A[728]), .B(B[728]), .CI(
        C[728]), .S(S[728]), .CO(C[729]) );
  FA_2343 \FA_INST_0[1].FA_INST_1[217].FA_  ( .A(A[729]), .B(B[729]), .CI(
        C[729]), .S(S[729]), .CO(C[730]) );
  FA_2342 \FA_INST_0[1].FA_INST_1[218].FA_  ( .A(A[730]), .B(B[730]), .CI(
        C[730]), .S(S[730]), .CO(C[731]) );
  FA_2341 \FA_INST_0[1].FA_INST_1[219].FA_  ( .A(A[731]), .B(B[731]), .CI(
        C[731]), .S(S[731]), .CO(C[732]) );
  FA_2340 \FA_INST_0[1].FA_INST_1[220].FA_  ( .A(A[732]), .B(B[732]), .CI(
        C[732]), .S(S[732]), .CO(C[733]) );
  FA_2339 \FA_INST_0[1].FA_INST_1[221].FA_  ( .A(A[733]), .B(B[733]), .CI(
        C[733]), .S(S[733]), .CO(C[734]) );
  FA_2338 \FA_INST_0[1].FA_INST_1[222].FA_  ( .A(A[734]), .B(B[734]), .CI(
        C[734]), .S(S[734]), .CO(C[735]) );
  FA_2337 \FA_INST_0[1].FA_INST_1[223].FA_  ( .A(A[735]), .B(B[735]), .CI(
        C[735]), .S(S[735]), .CO(C[736]) );
  FA_2336 \FA_INST_0[1].FA_INST_1[224].FA_  ( .A(A[736]), .B(B[736]), .CI(
        C[736]), .S(S[736]), .CO(C[737]) );
  FA_2335 \FA_INST_0[1].FA_INST_1[225].FA_  ( .A(A[737]), .B(B[737]), .CI(
        C[737]), .S(S[737]), .CO(C[738]) );
  FA_2334 \FA_INST_0[1].FA_INST_1[226].FA_  ( .A(A[738]), .B(B[738]), .CI(
        C[738]), .S(S[738]), .CO(C[739]) );
  FA_2333 \FA_INST_0[1].FA_INST_1[227].FA_  ( .A(A[739]), .B(B[739]), .CI(
        C[739]), .S(S[739]), .CO(C[740]) );
  FA_2332 \FA_INST_0[1].FA_INST_1[228].FA_  ( .A(A[740]), .B(B[740]), .CI(
        C[740]), .S(S[740]), .CO(C[741]) );
  FA_2331 \FA_INST_0[1].FA_INST_1[229].FA_  ( .A(A[741]), .B(B[741]), .CI(
        C[741]), .S(S[741]), .CO(C[742]) );
  FA_2330 \FA_INST_0[1].FA_INST_1[230].FA_  ( .A(A[742]), .B(B[742]), .CI(
        C[742]), .S(S[742]), .CO(C[743]) );
  FA_2329 \FA_INST_0[1].FA_INST_1[231].FA_  ( .A(A[743]), .B(B[743]), .CI(
        C[743]), .S(S[743]), .CO(C[744]) );
  FA_2328 \FA_INST_0[1].FA_INST_1[232].FA_  ( .A(A[744]), .B(B[744]), .CI(
        C[744]), .S(S[744]), .CO(C[745]) );
  FA_2327 \FA_INST_0[1].FA_INST_1[233].FA_  ( .A(A[745]), .B(B[745]), .CI(
        C[745]), .S(S[745]), .CO(C[746]) );
  FA_2326 \FA_INST_0[1].FA_INST_1[234].FA_  ( .A(A[746]), .B(B[746]), .CI(
        C[746]), .S(S[746]), .CO(C[747]) );
  FA_2325 \FA_INST_0[1].FA_INST_1[235].FA_  ( .A(A[747]), .B(B[747]), .CI(
        C[747]), .S(S[747]), .CO(C[748]) );
  FA_2324 \FA_INST_0[1].FA_INST_1[236].FA_  ( .A(A[748]), .B(B[748]), .CI(
        C[748]), .S(S[748]), .CO(C[749]) );
  FA_2323 \FA_INST_0[1].FA_INST_1[237].FA_  ( .A(A[749]), .B(B[749]), .CI(
        C[749]), .S(S[749]), .CO(C[750]) );
  FA_2322 \FA_INST_0[1].FA_INST_1[238].FA_  ( .A(A[750]), .B(B[750]), .CI(
        C[750]), .S(S[750]), .CO(C[751]) );
  FA_2321 \FA_INST_0[1].FA_INST_1[239].FA_  ( .A(A[751]), .B(B[751]), .CI(
        C[751]), .S(S[751]), .CO(C[752]) );
  FA_2320 \FA_INST_0[1].FA_INST_1[240].FA_  ( .A(A[752]), .B(B[752]), .CI(
        C[752]), .S(S[752]), .CO(C[753]) );
  FA_2319 \FA_INST_0[1].FA_INST_1[241].FA_  ( .A(A[753]), .B(B[753]), .CI(
        C[753]), .S(S[753]), .CO(C[754]) );
  FA_2318 \FA_INST_0[1].FA_INST_1[242].FA_  ( .A(A[754]), .B(B[754]), .CI(
        C[754]), .S(S[754]), .CO(C[755]) );
  FA_2317 \FA_INST_0[1].FA_INST_1[243].FA_  ( .A(A[755]), .B(B[755]), .CI(
        C[755]), .S(S[755]), .CO(C[756]) );
  FA_2316 \FA_INST_0[1].FA_INST_1[244].FA_  ( .A(A[756]), .B(B[756]), .CI(
        C[756]), .S(S[756]), .CO(C[757]) );
  FA_2315 \FA_INST_0[1].FA_INST_1[245].FA_  ( .A(A[757]), .B(B[757]), .CI(
        C[757]), .S(S[757]), .CO(C[758]) );
  FA_2314 \FA_INST_0[1].FA_INST_1[246].FA_  ( .A(A[758]), .B(B[758]), .CI(
        C[758]), .S(S[758]), .CO(C[759]) );
  FA_2313 \FA_INST_0[1].FA_INST_1[247].FA_  ( .A(A[759]), .B(B[759]), .CI(
        C[759]), .S(S[759]), .CO(C[760]) );
  FA_2312 \FA_INST_0[1].FA_INST_1[248].FA_  ( .A(A[760]), .B(B[760]), .CI(
        C[760]), .S(S[760]), .CO(C[761]) );
  FA_2311 \FA_INST_0[1].FA_INST_1[249].FA_  ( .A(A[761]), .B(B[761]), .CI(
        C[761]), .S(S[761]), .CO(C[762]) );
  FA_2310 \FA_INST_0[1].FA_INST_1[250].FA_  ( .A(A[762]), .B(B[762]), .CI(
        C[762]), .S(S[762]), .CO(C[763]) );
  FA_2309 \FA_INST_0[1].FA_INST_1[251].FA_  ( .A(A[763]), .B(B[763]), .CI(
        C[763]), .S(S[763]), .CO(C[764]) );
  FA_2308 \FA_INST_0[1].FA_INST_1[252].FA_  ( .A(A[764]), .B(B[764]), .CI(
        C[764]), .S(S[764]), .CO(C[765]) );
  FA_2307 \FA_INST_0[1].FA_INST_1[253].FA_  ( .A(A[765]), .B(B[765]), .CI(
        C[765]), .S(S[765]), .CO(C[766]) );
  FA_2306 \FA_INST_0[1].FA_INST_1[254].FA_  ( .A(A[766]), .B(B[766]), .CI(
        C[766]), .S(S[766]), .CO(C[767]) );
  FA_2305 \FA_INST_0[1].FA_INST_1[255].FA_  ( .A(A[767]), .B(B[767]), .CI(
        C[767]), .S(S[767]), .CO(C[768]) );
  FA_2304 \FA_INST_0[1].FA_INST_1[256].FA_  ( .A(A[768]), .B(B[768]), .CI(
        C[768]), .S(S[768]), .CO(C[769]) );
  FA_2303 \FA_INST_0[1].FA_INST_1[257].FA_  ( .A(A[769]), .B(B[769]), .CI(
        C[769]), .S(S[769]), .CO(C[770]) );
  FA_2302 \FA_INST_0[1].FA_INST_1[258].FA_  ( .A(A[770]), .B(B[770]), .CI(
        C[770]), .S(S[770]), .CO(C[771]) );
  FA_2301 \FA_INST_0[1].FA_INST_1[259].FA_  ( .A(A[771]), .B(B[771]), .CI(
        C[771]), .S(S[771]), .CO(C[772]) );
  FA_2300 \FA_INST_0[1].FA_INST_1[260].FA_  ( .A(A[772]), .B(B[772]), .CI(
        C[772]), .S(S[772]), .CO(C[773]) );
  FA_2299 \FA_INST_0[1].FA_INST_1[261].FA_  ( .A(A[773]), .B(B[773]), .CI(
        C[773]), .S(S[773]), .CO(C[774]) );
  FA_2298 \FA_INST_0[1].FA_INST_1[262].FA_  ( .A(A[774]), .B(B[774]), .CI(
        C[774]), .S(S[774]), .CO(C[775]) );
  FA_2297 \FA_INST_0[1].FA_INST_1[263].FA_  ( .A(A[775]), .B(B[775]), .CI(
        C[775]), .S(S[775]), .CO(C[776]) );
  FA_2296 \FA_INST_0[1].FA_INST_1[264].FA_  ( .A(A[776]), .B(B[776]), .CI(
        C[776]), .S(S[776]), .CO(C[777]) );
  FA_2295 \FA_INST_0[1].FA_INST_1[265].FA_  ( .A(A[777]), .B(B[777]), .CI(
        C[777]), .S(S[777]), .CO(C[778]) );
  FA_2294 \FA_INST_0[1].FA_INST_1[266].FA_  ( .A(A[778]), .B(B[778]), .CI(
        C[778]), .S(S[778]), .CO(C[779]) );
  FA_2293 \FA_INST_0[1].FA_INST_1[267].FA_  ( .A(A[779]), .B(B[779]), .CI(
        C[779]), .S(S[779]), .CO(C[780]) );
  FA_2292 \FA_INST_0[1].FA_INST_1[268].FA_  ( .A(A[780]), .B(B[780]), .CI(
        C[780]), .S(S[780]), .CO(C[781]) );
  FA_2291 \FA_INST_0[1].FA_INST_1[269].FA_  ( .A(A[781]), .B(B[781]), .CI(
        C[781]), .S(S[781]), .CO(C[782]) );
  FA_2290 \FA_INST_0[1].FA_INST_1[270].FA_  ( .A(A[782]), .B(B[782]), .CI(
        C[782]), .S(S[782]), .CO(C[783]) );
  FA_2289 \FA_INST_0[1].FA_INST_1[271].FA_  ( .A(A[783]), .B(B[783]), .CI(
        C[783]), .S(S[783]), .CO(C[784]) );
  FA_2288 \FA_INST_0[1].FA_INST_1[272].FA_  ( .A(A[784]), .B(B[784]), .CI(
        C[784]), .S(S[784]), .CO(C[785]) );
  FA_2287 \FA_INST_0[1].FA_INST_1[273].FA_  ( .A(A[785]), .B(B[785]), .CI(
        C[785]), .S(S[785]), .CO(C[786]) );
  FA_2286 \FA_INST_0[1].FA_INST_1[274].FA_  ( .A(A[786]), .B(B[786]), .CI(
        C[786]), .S(S[786]), .CO(C[787]) );
  FA_2285 \FA_INST_0[1].FA_INST_1[275].FA_  ( .A(A[787]), .B(B[787]), .CI(
        C[787]), .S(S[787]), .CO(C[788]) );
  FA_2284 \FA_INST_0[1].FA_INST_1[276].FA_  ( .A(A[788]), .B(B[788]), .CI(
        C[788]), .S(S[788]), .CO(C[789]) );
  FA_2283 \FA_INST_0[1].FA_INST_1[277].FA_  ( .A(A[789]), .B(B[789]), .CI(
        C[789]), .S(S[789]), .CO(C[790]) );
  FA_2282 \FA_INST_0[1].FA_INST_1[278].FA_  ( .A(A[790]), .B(B[790]), .CI(
        C[790]), .S(S[790]), .CO(C[791]) );
  FA_2281 \FA_INST_0[1].FA_INST_1[279].FA_  ( .A(A[791]), .B(B[791]), .CI(
        C[791]), .S(S[791]), .CO(C[792]) );
  FA_2280 \FA_INST_0[1].FA_INST_1[280].FA_  ( .A(A[792]), .B(B[792]), .CI(
        C[792]), .S(S[792]), .CO(C[793]) );
  FA_2279 \FA_INST_0[1].FA_INST_1[281].FA_  ( .A(A[793]), .B(B[793]), .CI(
        C[793]), .S(S[793]), .CO(C[794]) );
  FA_2278 \FA_INST_0[1].FA_INST_1[282].FA_  ( .A(A[794]), .B(B[794]), .CI(
        C[794]), .S(S[794]), .CO(C[795]) );
  FA_2277 \FA_INST_0[1].FA_INST_1[283].FA_  ( .A(A[795]), .B(B[795]), .CI(
        C[795]), .S(S[795]), .CO(C[796]) );
  FA_2276 \FA_INST_0[1].FA_INST_1[284].FA_  ( .A(A[796]), .B(B[796]), .CI(
        C[796]), .S(S[796]), .CO(C[797]) );
  FA_2275 \FA_INST_0[1].FA_INST_1[285].FA_  ( .A(A[797]), .B(B[797]), .CI(
        C[797]), .S(S[797]), .CO(C[798]) );
  FA_2274 \FA_INST_0[1].FA_INST_1[286].FA_  ( .A(A[798]), .B(B[798]), .CI(
        C[798]), .S(S[798]), .CO(C[799]) );
  FA_2273 \FA_INST_0[1].FA_INST_1[287].FA_  ( .A(A[799]), .B(B[799]), .CI(
        C[799]), .S(S[799]), .CO(C[800]) );
  FA_2272 \FA_INST_0[1].FA_INST_1[288].FA_  ( .A(A[800]), .B(B[800]), .CI(
        C[800]), .S(S[800]), .CO(C[801]) );
  FA_2271 \FA_INST_0[1].FA_INST_1[289].FA_  ( .A(A[801]), .B(B[801]), .CI(
        C[801]), .S(S[801]), .CO(C[802]) );
  FA_2270 \FA_INST_0[1].FA_INST_1[290].FA_  ( .A(A[802]), .B(B[802]), .CI(
        C[802]), .S(S[802]), .CO(C[803]) );
  FA_2269 \FA_INST_0[1].FA_INST_1[291].FA_  ( .A(A[803]), .B(B[803]), .CI(
        C[803]), .S(S[803]), .CO(C[804]) );
  FA_2268 \FA_INST_0[1].FA_INST_1[292].FA_  ( .A(A[804]), .B(B[804]), .CI(
        C[804]), .S(S[804]), .CO(C[805]) );
  FA_2267 \FA_INST_0[1].FA_INST_1[293].FA_  ( .A(A[805]), .B(B[805]), .CI(
        C[805]), .S(S[805]), .CO(C[806]) );
  FA_2266 \FA_INST_0[1].FA_INST_1[294].FA_  ( .A(A[806]), .B(B[806]), .CI(
        C[806]), .S(S[806]), .CO(C[807]) );
  FA_2265 \FA_INST_0[1].FA_INST_1[295].FA_  ( .A(A[807]), .B(B[807]), .CI(
        C[807]), .S(S[807]), .CO(C[808]) );
  FA_2264 \FA_INST_0[1].FA_INST_1[296].FA_  ( .A(A[808]), .B(B[808]), .CI(
        C[808]), .S(S[808]), .CO(C[809]) );
  FA_2263 \FA_INST_0[1].FA_INST_1[297].FA_  ( .A(A[809]), .B(B[809]), .CI(
        C[809]), .S(S[809]), .CO(C[810]) );
  FA_2262 \FA_INST_0[1].FA_INST_1[298].FA_  ( .A(A[810]), .B(B[810]), .CI(
        C[810]), .S(S[810]), .CO(C[811]) );
  FA_2261 \FA_INST_0[1].FA_INST_1[299].FA_  ( .A(A[811]), .B(B[811]), .CI(
        C[811]), .S(S[811]), .CO(C[812]) );
  FA_2260 \FA_INST_0[1].FA_INST_1[300].FA_  ( .A(A[812]), .B(B[812]), .CI(
        C[812]), .S(S[812]), .CO(C[813]) );
  FA_2259 \FA_INST_0[1].FA_INST_1[301].FA_  ( .A(A[813]), .B(B[813]), .CI(
        C[813]), .S(S[813]), .CO(C[814]) );
  FA_2258 \FA_INST_0[1].FA_INST_1[302].FA_  ( .A(A[814]), .B(B[814]), .CI(
        C[814]), .S(S[814]), .CO(C[815]) );
  FA_2257 \FA_INST_0[1].FA_INST_1[303].FA_  ( .A(A[815]), .B(B[815]), .CI(
        C[815]), .S(S[815]), .CO(C[816]) );
  FA_2256 \FA_INST_0[1].FA_INST_1[304].FA_  ( .A(A[816]), .B(B[816]), .CI(
        C[816]), .S(S[816]), .CO(C[817]) );
  FA_2255 \FA_INST_0[1].FA_INST_1[305].FA_  ( .A(A[817]), .B(B[817]), .CI(
        C[817]), .S(S[817]), .CO(C[818]) );
  FA_2254 \FA_INST_0[1].FA_INST_1[306].FA_  ( .A(A[818]), .B(B[818]), .CI(
        C[818]), .S(S[818]), .CO(C[819]) );
  FA_2253 \FA_INST_0[1].FA_INST_1[307].FA_  ( .A(A[819]), .B(B[819]), .CI(
        C[819]), .S(S[819]), .CO(C[820]) );
  FA_2252 \FA_INST_0[1].FA_INST_1[308].FA_  ( .A(A[820]), .B(B[820]), .CI(
        C[820]), .S(S[820]), .CO(C[821]) );
  FA_2251 \FA_INST_0[1].FA_INST_1[309].FA_  ( .A(A[821]), .B(B[821]), .CI(
        C[821]), .S(S[821]), .CO(C[822]) );
  FA_2250 \FA_INST_0[1].FA_INST_1[310].FA_  ( .A(A[822]), .B(B[822]), .CI(
        C[822]), .S(S[822]), .CO(C[823]) );
  FA_2249 \FA_INST_0[1].FA_INST_1[311].FA_  ( .A(A[823]), .B(B[823]), .CI(
        C[823]), .S(S[823]), .CO(C[824]) );
  FA_2248 \FA_INST_0[1].FA_INST_1[312].FA_  ( .A(A[824]), .B(B[824]), .CI(
        C[824]), .S(S[824]), .CO(C[825]) );
  FA_2247 \FA_INST_0[1].FA_INST_1[313].FA_  ( .A(A[825]), .B(B[825]), .CI(
        C[825]), .S(S[825]), .CO(C[826]) );
  FA_2246 \FA_INST_0[1].FA_INST_1[314].FA_  ( .A(A[826]), .B(B[826]), .CI(
        C[826]), .S(S[826]), .CO(C[827]) );
  FA_2245 \FA_INST_0[1].FA_INST_1[315].FA_  ( .A(A[827]), .B(B[827]), .CI(
        C[827]), .S(S[827]), .CO(C[828]) );
  FA_2244 \FA_INST_0[1].FA_INST_1[316].FA_  ( .A(A[828]), .B(B[828]), .CI(
        C[828]), .S(S[828]), .CO(C[829]) );
  FA_2243 \FA_INST_0[1].FA_INST_1[317].FA_  ( .A(A[829]), .B(B[829]), .CI(
        C[829]), .S(S[829]), .CO(C[830]) );
  FA_2242 \FA_INST_0[1].FA_INST_1[318].FA_  ( .A(A[830]), .B(B[830]), .CI(
        C[830]), .S(S[830]), .CO(C[831]) );
  FA_2241 \FA_INST_0[1].FA_INST_1[319].FA_  ( .A(A[831]), .B(B[831]), .CI(
        C[831]), .S(S[831]), .CO(C[832]) );
  FA_2240 \FA_INST_0[1].FA_INST_1[320].FA_  ( .A(A[832]), .B(B[832]), .CI(
        C[832]), .S(S[832]), .CO(C[833]) );
  FA_2239 \FA_INST_0[1].FA_INST_1[321].FA_  ( .A(A[833]), .B(B[833]), .CI(
        C[833]), .S(S[833]), .CO(C[834]) );
  FA_2238 \FA_INST_0[1].FA_INST_1[322].FA_  ( .A(A[834]), .B(B[834]), .CI(
        C[834]), .S(S[834]), .CO(C[835]) );
  FA_2237 \FA_INST_0[1].FA_INST_1[323].FA_  ( .A(A[835]), .B(B[835]), .CI(
        C[835]), .S(S[835]), .CO(C[836]) );
  FA_2236 \FA_INST_0[1].FA_INST_1[324].FA_  ( .A(A[836]), .B(B[836]), .CI(
        C[836]), .S(S[836]), .CO(C[837]) );
  FA_2235 \FA_INST_0[1].FA_INST_1[325].FA_  ( .A(A[837]), .B(B[837]), .CI(
        C[837]), .S(S[837]), .CO(C[838]) );
  FA_2234 \FA_INST_0[1].FA_INST_1[326].FA_  ( .A(A[838]), .B(B[838]), .CI(
        C[838]), .S(S[838]), .CO(C[839]) );
  FA_2233 \FA_INST_0[1].FA_INST_1[327].FA_  ( .A(A[839]), .B(B[839]), .CI(
        C[839]), .S(S[839]), .CO(C[840]) );
  FA_2232 \FA_INST_0[1].FA_INST_1[328].FA_  ( .A(A[840]), .B(B[840]), .CI(
        C[840]), .S(S[840]), .CO(C[841]) );
  FA_2231 \FA_INST_0[1].FA_INST_1[329].FA_  ( .A(A[841]), .B(B[841]), .CI(
        C[841]), .S(S[841]), .CO(C[842]) );
  FA_2230 \FA_INST_0[1].FA_INST_1[330].FA_  ( .A(A[842]), .B(B[842]), .CI(
        C[842]), .S(S[842]), .CO(C[843]) );
  FA_2229 \FA_INST_0[1].FA_INST_1[331].FA_  ( .A(A[843]), .B(B[843]), .CI(
        C[843]), .S(S[843]), .CO(C[844]) );
  FA_2228 \FA_INST_0[1].FA_INST_1[332].FA_  ( .A(A[844]), .B(B[844]), .CI(
        C[844]), .S(S[844]), .CO(C[845]) );
  FA_2227 \FA_INST_0[1].FA_INST_1[333].FA_  ( .A(A[845]), .B(B[845]), .CI(
        C[845]), .S(S[845]), .CO(C[846]) );
  FA_2226 \FA_INST_0[1].FA_INST_1[334].FA_  ( .A(A[846]), .B(B[846]), .CI(
        C[846]), .S(S[846]), .CO(C[847]) );
  FA_2225 \FA_INST_0[1].FA_INST_1[335].FA_  ( .A(A[847]), .B(B[847]), .CI(
        C[847]), .S(S[847]), .CO(C[848]) );
  FA_2224 \FA_INST_0[1].FA_INST_1[336].FA_  ( .A(A[848]), .B(B[848]), .CI(
        C[848]), .S(S[848]), .CO(C[849]) );
  FA_2223 \FA_INST_0[1].FA_INST_1[337].FA_  ( .A(A[849]), .B(B[849]), .CI(
        C[849]), .S(S[849]), .CO(C[850]) );
  FA_2222 \FA_INST_0[1].FA_INST_1[338].FA_  ( .A(A[850]), .B(B[850]), .CI(
        C[850]), .S(S[850]), .CO(C[851]) );
  FA_2221 \FA_INST_0[1].FA_INST_1[339].FA_  ( .A(A[851]), .B(B[851]), .CI(
        C[851]), .S(S[851]), .CO(C[852]) );
  FA_2220 \FA_INST_0[1].FA_INST_1[340].FA_  ( .A(A[852]), .B(B[852]), .CI(
        C[852]), .S(S[852]), .CO(C[853]) );
  FA_2219 \FA_INST_0[1].FA_INST_1[341].FA_  ( .A(A[853]), .B(B[853]), .CI(
        C[853]), .S(S[853]), .CO(C[854]) );
  FA_2218 \FA_INST_0[1].FA_INST_1[342].FA_  ( .A(A[854]), .B(B[854]), .CI(
        C[854]), .S(S[854]), .CO(C[855]) );
  FA_2217 \FA_INST_0[1].FA_INST_1[343].FA_  ( .A(A[855]), .B(B[855]), .CI(
        C[855]), .S(S[855]), .CO(C[856]) );
  FA_2216 \FA_INST_0[1].FA_INST_1[344].FA_  ( .A(A[856]), .B(B[856]), .CI(
        C[856]), .S(S[856]), .CO(C[857]) );
  FA_2215 \FA_INST_0[1].FA_INST_1[345].FA_  ( .A(A[857]), .B(B[857]), .CI(
        C[857]), .S(S[857]), .CO(C[858]) );
  FA_2214 \FA_INST_0[1].FA_INST_1[346].FA_  ( .A(A[858]), .B(B[858]), .CI(
        C[858]), .S(S[858]), .CO(C[859]) );
  FA_2213 \FA_INST_0[1].FA_INST_1[347].FA_  ( .A(A[859]), .B(B[859]), .CI(
        C[859]), .S(S[859]), .CO(C[860]) );
  FA_2212 \FA_INST_0[1].FA_INST_1[348].FA_  ( .A(A[860]), .B(B[860]), .CI(
        C[860]), .S(S[860]), .CO(C[861]) );
  FA_2211 \FA_INST_0[1].FA_INST_1[349].FA_  ( .A(A[861]), .B(B[861]), .CI(
        C[861]), .S(S[861]), .CO(C[862]) );
  FA_2210 \FA_INST_0[1].FA_INST_1[350].FA_  ( .A(A[862]), .B(B[862]), .CI(
        C[862]), .S(S[862]), .CO(C[863]) );
  FA_2209 \FA_INST_0[1].FA_INST_1[351].FA_  ( .A(A[863]), .B(B[863]), .CI(
        C[863]), .S(S[863]), .CO(C[864]) );
  FA_2208 \FA_INST_0[1].FA_INST_1[352].FA_  ( .A(A[864]), .B(B[864]), .CI(
        C[864]), .S(S[864]), .CO(C[865]) );
  FA_2207 \FA_INST_0[1].FA_INST_1[353].FA_  ( .A(A[865]), .B(B[865]), .CI(
        C[865]), .S(S[865]), .CO(C[866]) );
  FA_2206 \FA_INST_0[1].FA_INST_1[354].FA_  ( .A(A[866]), .B(B[866]), .CI(
        C[866]), .S(S[866]), .CO(C[867]) );
  FA_2205 \FA_INST_0[1].FA_INST_1[355].FA_  ( .A(A[867]), .B(B[867]), .CI(
        C[867]), .S(S[867]), .CO(C[868]) );
  FA_2204 \FA_INST_0[1].FA_INST_1[356].FA_  ( .A(A[868]), .B(B[868]), .CI(
        C[868]), .S(S[868]), .CO(C[869]) );
  FA_2203 \FA_INST_0[1].FA_INST_1[357].FA_  ( .A(A[869]), .B(B[869]), .CI(
        C[869]), .S(S[869]), .CO(C[870]) );
  FA_2202 \FA_INST_0[1].FA_INST_1[358].FA_  ( .A(A[870]), .B(B[870]), .CI(
        C[870]), .S(S[870]), .CO(C[871]) );
  FA_2201 \FA_INST_0[1].FA_INST_1[359].FA_  ( .A(A[871]), .B(B[871]), .CI(
        C[871]), .S(S[871]), .CO(C[872]) );
  FA_2200 \FA_INST_0[1].FA_INST_1[360].FA_  ( .A(A[872]), .B(B[872]), .CI(
        C[872]), .S(S[872]), .CO(C[873]) );
  FA_2199 \FA_INST_0[1].FA_INST_1[361].FA_  ( .A(A[873]), .B(B[873]), .CI(
        C[873]), .S(S[873]), .CO(C[874]) );
  FA_2198 \FA_INST_0[1].FA_INST_1[362].FA_  ( .A(A[874]), .B(B[874]), .CI(
        C[874]), .S(S[874]), .CO(C[875]) );
  FA_2197 \FA_INST_0[1].FA_INST_1[363].FA_  ( .A(A[875]), .B(B[875]), .CI(
        C[875]), .S(S[875]), .CO(C[876]) );
  FA_2196 \FA_INST_0[1].FA_INST_1[364].FA_  ( .A(A[876]), .B(B[876]), .CI(
        C[876]), .S(S[876]), .CO(C[877]) );
  FA_2195 \FA_INST_0[1].FA_INST_1[365].FA_  ( .A(A[877]), .B(B[877]), .CI(
        C[877]), .S(S[877]), .CO(C[878]) );
  FA_2194 \FA_INST_0[1].FA_INST_1[366].FA_  ( .A(A[878]), .B(B[878]), .CI(
        C[878]), .S(S[878]), .CO(C[879]) );
  FA_2193 \FA_INST_0[1].FA_INST_1[367].FA_  ( .A(A[879]), .B(B[879]), .CI(
        C[879]), .S(S[879]), .CO(C[880]) );
  FA_2192 \FA_INST_0[1].FA_INST_1[368].FA_  ( .A(A[880]), .B(B[880]), .CI(
        C[880]), .S(S[880]), .CO(C[881]) );
  FA_2191 \FA_INST_0[1].FA_INST_1[369].FA_  ( .A(A[881]), .B(B[881]), .CI(
        C[881]), .S(S[881]), .CO(C[882]) );
  FA_2190 \FA_INST_0[1].FA_INST_1[370].FA_  ( .A(A[882]), .B(B[882]), .CI(
        C[882]), .S(S[882]), .CO(C[883]) );
  FA_2189 \FA_INST_0[1].FA_INST_1[371].FA_  ( .A(A[883]), .B(B[883]), .CI(
        C[883]), .S(S[883]), .CO(C[884]) );
  FA_2188 \FA_INST_0[1].FA_INST_1[372].FA_  ( .A(A[884]), .B(B[884]), .CI(
        C[884]), .S(S[884]), .CO(C[885]) );
  FA_2187 \FA_INST_0[1].FA_INST_1[373].FA_  ( .A(A[885]), .B(B[885]), .CI(
        C[885]), .S(S[885]), .CO(C[886]) );
  FA_2186 \FA_INST_0[1].FA_INST_1[374].FA_  ( .A(A[886]), .B(B[886]), .CI(
        C[886]), .S(S[886]), .CO(C[887]) );
  FA_2185 \FA_INST_0[1].FA_INST_1[375].FA_  ( .A(A[887]), .B(B[887]), .CI(
        C[887]), .S(S[887]), .CO(C[888]) );
  FA_2184 \FA_INST_0[1].FA_INST_1[376].FA_  ( .A(A[888]), .B(B[888]), .CI(
        C[888]), .S(S[888]), .CO(C[889]) );
  FA_2183 \FA_INST_0[1].FA_INST_1[377].FA_  ( .A(A[889]), .B(B[889]), .CI(
        C[889]), .S(S[889]), .CO(C[890]) );
  FA_2182 \FA_INST_0[1].FA_INST_1[378].FA_  ( .A(A[890]), .B(B[890]), .CI(
        C[890]), .S(S[890]), .CO(C[891]) );
  FA_2181 \FA_INST_0[1].FA_INST_1[379].FA_  ( .A(A[891]), .B(B[891]), .CI(
        C[891]), .S(S[891]), .CO(C[892]) );
  FA_2180 \FA_INST_0[1].FA_INST_1[380].FA_  ( .A(A[892]), .B(B[892]), .CI(
        C[892]), .S(S[892]), .CO(C[893]) );
  FA_2179 \FA_INST_0[1].FA_INST_1[381].FA_  ( .A(A[893]), .B(B[893]), .CI(
        C[893]), .S(S[893]), .CO(C[894]) );
  FA_2178 \FA_INST_0[1].FA_INST_1[382].FA_  ( .A(A[894]), .B(B[894]), .CI(
        C[894]), .S(S[894]), .CO(C[895]) );
  FA_2177 \FA_INST_0[1].FA_INST_1[383].FA_  ( .A(A[895]), .B(B[895]), .CI(
        C[895]), .S(S[895]), .CO(C[896]) );
  FA_2176 \FA_INST_0[1].FA_INST_1[384].FA_  ( .A(A[896]), .B(B[896]), .CI(
        C[896]), .S(S[896]), .CO(C[897]) );
  FA_2175 \FA_INST_0[1].FA_INST_1[385].FA_  ( .A(A[897]), .B(B[897]), .CI(
        C[897]), .S(S[897]), .CO(C[898]) );
  FA_2174 \FA_INST_0[1].FA_INST_1[386].FA_  ( .A(A[898]), .B(B[898]), .CI(
        C[898]), .S(S[898]), .CO(C[899]) );
  FA_2173 \FA_INST_0[1].FA_INST_1[387].FA_  ( .A(A[899]), .B(B[899]), .CI(
        C[899]), .S(S[899]), .CO(C[900]) );
  FA_2172 \FA_INST_0[1].FA_INST_1[388].FA_  ( .A(A[900]), .B(B[900]), .CI(
        C[900]), .S(S[900]), .CO(C[901]) );
  FA_2171 \FA_INST_0[1].FA_INST_1[389].FA_  ( .A(A[901]), .B(B[901]), .CI(
        C[901]), .S(S[901]), .CO(C[902]) );
  FA_2170 \FA_INST_0[1].FA_INST_1[390].FA_  ( .A(A[902]), .B(B[902]), .CI(
        C[902]), .S(S[902]), .CO(C[903]) );
  FA_2169 \FA_INST_0[1].FA_INST_1[391].FA_  ( .A(A[903]), .B(B[903]), .CI(
        C[903]), .S(S[903]), .CO(C[904]) );
  FA_2168 \FA_INST_0[1].FA_INST_1[392].FA_  ( .A(A[904]), .B(B[904]), .CI(
        C[904]), .S(S[904]), .CO(C[905]) );
  FA_2167 \FA_INST_0[1].FA_INST_1[393].FA_  ( .A(A[905]), .B(B[905]), .CI(
        C[905]), .S(S[905]), .CO(C[906]) );
  FA_2166 \FA_INST_0[1].FA_INST_1[394].FA_  ( .A(A[906]), .B(B[906]), .CI(
        C[906]), .S(S[906]), .CO(C[907]) );
  FA_2165 \FA_INST_0[1].FA_INST_1[395].FA_  ( .A(A[907]), .B(B[907]), .CI(
        C[907]), .S(S[907]), .CO(C[908]) );
  FA_2164 \FA_INST_0[1].FA_INST_1[396].FA_  ( .A(A[908]), .B(B[908]), .CI(
        C[908]), .S(S[908]), .CO(C[909]) );
  FA_2163 \FA_INST_0[1].FA_INST_1[397].FA_  ( .A(A[909]), .B(B[909]), .CI(
        C[909]), .S(S[909]), .CO(C[910]) );
  FA_2162 \FA_INST_0[1].FA_INST_1[398].FA_  ( .A(A[910]), .B(B[910]), .CI(
        C[910]), .S(S[910]), .CO(C[911]) );
  FA_2161 \FA_INST_0[1].FA_INST_1[399].FA_  ( .A(A[911]), .B(B[911]), .CI(
        C[911]), .S(S[911]), .CO(C[912]) );
  FA_2160 \FA_INST_0[1].FA_INST_1[400].FA_  ( .A(A[912]), .B(B[912]), .CI(
        C[912]), .S(S[912]), .CO(C[913]) );
  FA_2159 \FA_INST_0[1].FA_INST_1[401].FA_  ( .A(A[913]), .B(B[913]), .CI(
        C[913]), .S(S[913]), .CO(C[914]) );
  FA_2158 \FA_INST_0[1].FA_INST_1[402].FA_  ( .A(A[914]), .B(B[914]), .CI(
        C[914]), .S(S[914]), .CO(C[915]) );
  FA_2157 \FA_INST_0[1].FA_INST_1[403].FA_  ( .A(A[915]), .B(B[915]), .CI(
        C[915]), .S(S[915]), .CO(C[916]) );
  FA_2156 \FA_INST_0[1].FA_INST_1[404].FA_  ( .A(A[916]), .B(B[916]), .CI(
        C[916]), .S(S[916]), .CO(C[917]) );
  FA_2155 \FA_INST_0[1].FA_INST_1[405].FA_  ( .A(A[917]), .B(B[917]), .CI(
        C[917]), .S(S[917]), .CO(C[918]) );
  FA_2154 \FA_INST_0[1].FA_INST_1[406].FA_  ( .A(A[918]), .B(B[918]), .CI(
        C[918]), .S(S[918]), .CO(C[919]) );
  FA_2153 \FA_INST_0[1].FA_INST_1[407].FA_  ( .A(A[919]), .B(B[919]), .CI(
        C[919]), .S(S[919]), .CO(C[920]) );
  FA_2152 \FA_INST_0[1].FA_INST_1[408].FA_  ( .A(A[920]), .B(B[920]), .CI(
        C[920]), .S(S[920]), .CO(C[921]) );
  FA_2151 \FA_INST_0[1].FA_INST_1[409].FA_  ( .A(A[921]), .B(B[921]), .CI(
        C[921]), .S(S[921]), .CO(C[922]) );
  FA_2150 \FA_INST_0[1].FA_INST_1[410].FA_  ( .A(A[922]), .B(B[922]), .CI(
        C[922]), .S(S[922]), .CO(C[923]) );
  FA_2149 \FA_INST_0[1].FA_INST_1[411].FA_  ( .A(A[923]), .B(B[923]), .CI(
        C[923]), .S(S[923]), .CO(C[924]) );
  FA_2148 \FA_INST_0[1].FA_INST_1[412].FA_  ( .A(A[924]), .B(B[924]), .CI(
        C[924]), .S(S[924]), .CO(C[925]) );
  FA_2147 \FA_INST_0[1].FA_INST_1[413].FA_  ( .A(A[925]), .B(B[925]), .CI(
        C[925]), .S(S[925]), .CO(C[926]) );
  FA_2146 \FA_INST_0[1].FA_INST_1[414].FA_  ( .A(A[926]), .B(B[926]), .CI(
        C[926]), .S(S[926]), .CO(C[927]) );
  FA_2145 \FA_INST_0[1].FA_INST_1[415].FA_  ( .A(A[927]), .B(B[927]), .CI(
        C[927]), .S(S[927]), .CO(C[928]) );
  FA_2144 \FA_INST_0[1].FA_INST_1[416].FA_  ( .A(A[928]), .B(B[928]), .CI(
        C[928]), .S(S[928]), .CO(C[929]) );
  FA_2143 \FA_INST_0[1].FA_INST_1[417].FA_  ( .A(A[929]), .B(B[929]), .CI(
        C[929]), .S(S[929]), .CO(C[930]) );
  FA_2142 \FA_INST_0[1].FA_INST_1[418].FA_  ( .A(A[930]), .B(B[930]), .CI(
        C[930]), .S(S[930]), .CO(C[931]) );
  FA_2141 \FA_INST_0[1].FA_INST_1[419].FA_  ( .A(A[931]), .B(B[931]), .CI(
        C[931]), .S(S[931]), .CO(C[932]) );
  FA_2140 \FA_INST_0[1].FA_INST_1[420].FA_  ( .A(A[932]), .B(B[932]), .CI(
        C[932]), .S(S[932]), .CO(C[933]) );
  FA_2139 \FA_INST_0[1].FA_INST_1[421].FA_  ( .A(A[933]), .B(B[933]), .CI(
        C[933]), .S(S[933]), .CO(C[934]) );
  FA_2138 \FA_INST_0[1].FA_INST_1[422].FA_  ( .A(A[934]), .B(B[934]), .CI(
        C[934]), .S(S[934]), .CO(C[935]) );
  FA_2137 \FA_INST_0[1].FA_INST_1[423].FA_  ( .A(A[935]), .B(B[935]), .CI(
        C[935]), .S(S[935]), .CO(C[936]) );
  FA_2136 \FA_INST_0[1].FA_INST_1[424].FA_  ( .A(A[936]), .B(B[936]), .CI(
        C[936]), .S(S[936]), .CO(C[937]) );
  FA_2135 \FA_INST_0[1].FA_INST_1[425].FA_  ( .A(A[937]), .B(B[937]), .CI(
        C[937]), .S(S[937]), .CO(C[938]) );
  FA_2134 \FA_INST_0[1].FA_INST_1[426].FA_  ( .A(A[938]), .B(B[938]), .CI(
        C[938]), .S(S[938]), .CO(C[939]) );
  FA_2133 \FA_INST_0[1].FA_INST_1[427].FA_  ( .A(A[939]), .B(B[939]), .CI(
        C[939]), .S(S[939]), .CO(C[940]) );
  FA_2132 \FA_INST_0[1].FA_INST_1[428].FA_  ( .A(A[940]), .B(B[940]), .CI(
        C[940]), .S(S[940]), .CO(C[941]) );
  FA_2131 \FA_INST_0[1].FA_INST_1[429].FA_  ( .A(A[941]), .B(B[941]), .CI(
        C[941]), .S(S[941]), .CO(C[942]) );
  FA_2130 \FA_INST_0[1].FA_INST_1[430].FA_  ( .A(A[942]), .B(B[942]), .CI(
        C[942]), .S(S[942]), .CO(C[943]) );
  FA_2129 \FA_INST_0[1].FA_INST_1[431].FA_  ( .A(A[943]), .B(B[943]), .CI(
        C[943]), .S(S[943]), .CO(C[944]) );
  FA_2128 \FA_INST_0[1].FA_INST_1[432].FA_  ( .A(A[944]), .B(B[944]), .CI(
        C[944]), .S(S[944]), .CO(C[945]) );
  FA_2127 \FA_INST_0[1].FA_INST_1[433].FA_  ( .A(A[945]), .B(B[945]), .CI(
        C[945]), .S(S[945]), .CO(C[946]) );
  FA_2126 \FA_INST_0[1].FA_INST_1[434].FA_  ( .A(A[946]), .B(B[946]), .CI(
        C[946]), .S(S[946]), .CO(C[947]) );
  FA_2125 \FA_INST_0[1].FA_INST_1[435].FA_  ( .A(A[947]), .B(B[947]), .CI(
        C[947]), .S(S[947]), .CO(C[948]) );
  FA_2124 \FA_INST_0[1].FA_INST_1[436].FA_  ( .A(A[948]), .B(B[948]), .CI(
        C[948]), .S(S[948]), .CO(C[949]) );
  FA_2123 \FA_INST_0[1].FA_INST_1[437].FA_  ( .A(A[949]), .B(B[949]), .CI(
        C[949]), .S(S[949]), .CO(C[950]) );
  FA_2122 \FA_INST_0[1].FA_INST_1[438].FA_  ( .A(A[950]), .B(B[950]), .CI(
        C[950]), .S(S[950]), .CO(C[951]) );
  FA_2121 \FA_INST_0[1].FA_INST_1[439].FA_  ( .A(A[951]), .B(B[951]), .CI(
        C[951]), .S(S[951]), .CO(C[952]) );
  FA_2120 \FA_INST_0[1].FA_INST_1[440].FA_  ( .A(A[952]), .B(B[952]), .CI(
        C[952]), .S(S[952]), .CO(C[953]) );
  FA_2119 \FA_INST_0[1].FA_INST_1[441].FA_  ( .A(A[953]), .B(B[953]), .CI(
        C[953]), .S(S[953]), .CO(C[954]) );
  FA_2118 \FA_INST_0[1].FA_INST_1[442].FA_  ( .A(A[954]), .B(B[954]), .CI(
        C[954]), .S(S[954]), .CO(C[955]) );
  FA_2117 \FA_INST_0[1].FA_INST_1[443].FA_  ( .A(A[955]), .B(B[955]), .CI(
        C[955]), .S(S[955]), .CO(C[956]) );
  FA_2116 \FA_INST_0[1].FA_INST_1[444].FA_  ( .A(A[956]), .B(B[956]), .CI(
        C[956]), .S(S[956]), .CO(C[957]) );
  FA_2115 \FA_INST_0[1].FA_INST_1[445].FA_  ( .A(A[957]), .B(B[957]), .CI(
        C[957]), .S(S[957]), .CO(C[958]) );
  FA_2114 \FA_INST_0[1].FA_INST_1[446].FA_  ( .A(A[958]), .B(B[958]), .CI(
        C[958]), .S(S[958]), .CO(C[959]) );
  FA_2113 \FA_INST_0[1].FA_INST_1[447].FA_  ( .A(A[959]), .B(B[959]), .CI(
        C[959]), .S(S[959]), .CO(C[960]) );
  FA_2112 \FA_INST_0[1].FA_INST_1[448].FA_  ( .A(A[960]), .B(B[960]), .CI(
        C[960]), .S(S[960]), .CO(C[961]) );
  FA_2111 \FA_INST_0[1].FA_INST_1[449].FA_  ( .A(A[961]), .B(B[961]), .CI(
        C[961]), .S(S[961]), .CO(C[962]) );
  FA_2110 \FA_INST_0[1].FA_INST_1[450].FA_  ( .A(A[962]), .B(B[962]), .CI(
        C[962]), .S(S[962]), .CO(C[963]) );
  FA_2109 \FA_INST_0[1].FA_INST_1[451].FA_  ( .A(A[963]), .B(B[963]), .CI(
        C[963]), .S(S[963]), .CO(C[964]) );
  FA_2108 \FA_INST_0[1].FA_INST_1[452].FA_  ( .A(A[964]), .B(B[964]), .CI(
        C[964]), .S(S[964]), .CO(C[965]) );
  FA_2107 \FA_INST_0[1].FA_INST_1[453].FA_  ( .A(A[965]), .B(B[965]), .CI(
        C[965]), .S(S[965]), .CO(C[966]) );
  FA_2106 \FA_INST_0[1].FA_INST_1[454].FA_  ( .A(A[966]), .B(B[966]), .CI(
        C[966]), .S(S[966]), .CO(C[967]) );
  FA_2105 \FA_INST_0[1].FA_INST_1[455].FA_  ( .A(A[967]), .B(B[967]), .CI(
        C[967]), .S(S[967]), .CO(C[968]) );
  FA_2104 \FA_INST_0[1].FA_INST_1[456].FA_  ( .A(A[968]), .B(B[968]), .CI(
        C[968]), .S(S[968]), .CO(C[969]) );
  FA_2103 \FA_INST_0[1].FA_INST_1[457].FA_  ( .A(A[969]), .B(B[969]), .CI(
        C[969]), .S(S[969]), .CO(C[970]) );
  FA_2102 \FA_INST_0[1].FA_INST_1[458].FA_  ( .A(A[970]), .B(B[970]), .CI(
        C[970]), .S(S[970]), .CO(C[971]) );
  FA_2101 \FA_INST_0[1].FA_INST_1[459].FA_  ( .A(A[971]), .B(B[971]), .CI(
        C[971]), .S(S[971]), .CO(C[972]) );
  FA_2100 \FA_INST_0[1].FA_INST_1[460].FA_  ( .A(A[972]), .B(B[972]), .CI(
        C[972]), .S(S[972]), .CO(C[973]) );
  FA_2099 \FA_INST_0[1].FA_INST_1[461].FA_  ( .A(A[973]), .B(B[973]), .CI(
        C[973]), .S(S[973]), .CO(C[974]) );
  FA_2098 \FA_INST_0[1].FA_INST_1[462].FA_  ( .A(A[974]), .B(B[974]), .CI(
        C[974]), .S(S[974]), .CO(C[975]) );
  FA_2097 \FA_INST_0[1].FA_INST_1[463].FA_  ( .A(A[975]), .B(B[975]), .CI(
        C[975]), .S(S[975]), .CO(C[976]) );
  FA_2096 \FA_INST_0[1].FA_INST_1[464].FA_  ( .A(A[976]), .B(B[976]), .CI(
        C[976]), .S(S[976]), .CO(C[977]) );
  FA_2095 \FA_INST_0[1].FA_INST_1[465].FA_  ( .A(A[977]), .B(B[977]), .CI(
        C[977]), .S(S[977]), .CO(C[978]) );
  FA_2094 \FA_INST_0[1].FA_INST_1[466].FA_  ( .A(A[978]), .B(B[978]), .CI(
        C[978]), .S(S[978]), .CO(C[979]) );
  FA_2093 \FA_INST_0[1].FA_INST_1[467].FA_  ( .A(A[979]), .B(B[979]), .CI(
        C[979]), .S(S[979]), .CO(C[980]) );
  FA_2092 \FA_INST_0[1].FA_INST_1[468].FA_  ( .A(A[980]), .B(B[980]), .CI(
        C[980]), .S(S[980]), .CO(C[981]) );
  FA_2091 \FA_INST_0[1].FA_INST_1[469].FA_  ( .A(A[981]), .B(B[981]), .CI(
        C[981]), .S(S[981]), .CO(C[982]) );
  FA_2090 \FA_INST_0[1].FA_INST_1[470].FA_  ( .A(A[982]), .B(B[982]), .CI(
        C[982]), .S(S[982]), .CO(C[983]) );
  FA_2089 \FA_INST_0[1].FA_INST_1[471].FA_  ( .A(A[983]), .B(B[983]), .CI(
        C[983]), .S(S[983]), .CO(C[984]) );
  FA_2088 \FA_INST_0[1].FA_INST_1[472].FA_  ( .A(A[984]), .B(B[984]), .CI(
        C[984]), .S(S[984]), .CO(C[985]) );
  FA_2087 \FA_INST_0[1].FA_INST_1[473].FA_  ( .A(A[985]), .B(B[985]), .CI(
        C[985]), .S(S[985]), .CO(C[986]) );
  FA_2086 \FA_INST_0[1].FA_INST_1[474].FA_  ( .A(A[986]), .B(B[986]), .CI(
        C[986]), .S(S[986]), .CO(C[987]) );
  FA_2085 \FA_INST_0[1].FA_INST_1[475].FA_  ( .A(A[987]), .B(B[987]), .CI(
        C[987]), .S(S[987]), .CO(C[988]) );
  FA_2084 \FA_INST_0[1].FA_INST_1[476].FA_  ( .A(A[988]), .B(B[988]), .CI(
        C[988]), .S(S[988]), .CO(C[989]) );
  FA_2083 \FA_INST_0[1].FA_INST_1[477].FA_  ( .A(A[989]), .B(B[989]), .CI(
        C[989]), .S(S[989]), .CO(C[990]) );
  FA_2082 \FA_INST_0[1].FA_INST_1[478].FA_  ( .A(A[990]), .B(B[990]), .CI(
        C[990]), .S(S[990]), .CO(C[991]) );
  FA_2081 \FA_INST_0[1].FA_INST_1[479].FA_  ( .A(A[991]), .B(B[991]), .CI(
        C[991]), .S(S[991]), .CO(C[992]) );
  FA_2080 \FA_INST_0[1].FA_INST_1[480].FA_  ( .A(A[992]), .B(B[992]), .CI(
        C[992]), .S(S[992]), .CO(C[993]) );
  FA_2079 \FA_INST_0[1].FA_INST_1[481].FA_  ( .A(A[993]), .B(B[993]), .CI(
        C[993]), .S(S[993]), .CO(C[994]) );
  FA_2078 \FA_INST_0[1].FA_INST_1[482].FA_  ( .A(A[994]), .B(B[994]), .CI(
        C[994]), .S(S[994]), .CO(C[995]) );
  FA_2077 \FA_INST_0[1].FA_INST_1[483].FA_  ( .A(A[995]), .B(B[995]), .CI(
        C[995]), .S(S[995]), .CO(C[996]) );
  FA_2076 \FA_INST_0[1].FA_INST_1[484].FA_  ( .A(A[996]), .B(B[996]), .CI(
        C[996]), .S(S[996]), .CO(C[997]) );
  FA_2075 \FA_INST_0[1].FA_INST_1[485].FA_  ( .A(A[997]), .B(B[997]), .CI(
        C[997]), .S(S[997]), .CO(C[998]) );
  FA_2074 \FA_INST_0[1].FA_INST_1[486].FA_  ( .A(A[998]), .B(B[998]), .CI(
        C[998]), .S(S[998]), .CO(C[999]) );
  FA_2073 \FA_INST_0[1].FA_INST_1[487].FA_  ( .A(A[999]), .B(B[999]), .CI(
        C[999]), .S(S[999]), .CO(C[1000]) );
  FA_2072 \FA_INST_0[1].FA_INST_1[488].FA_  ( .A(A[1000]), .B(B[1000]), .CI(
        C[1000]), .S(S[1000]), .CO(C[1001]) );
  FA_2071 \FA_INST_0[1].FA_INST_1[489].FA_  ( .A(A[1001]), .B(B[1001]), .CI(
        C[1001]), .S(S[1001]), .CO(C[1002]) );
  FA_2070 \FA_INST_0[1].FA_INST_1[490].FA_  ( .A(A[1002]), .B(B[1002]), .CI(
        C[1002]), .S(S[1002]), .CO(C[1003]) );
  FA_2069 \FA_INST_0[1].FA_INST_1[491].FA_  ( .A(A[1003]), .B(B[1003]), .CI(
        C[1003]), .S(S[1003]), .CO(C[1004]) );
  FA_2068 \FA_INST_0[1].FA_INST_1[492].FA_  ( .A(A[1004]), .B(B[1004]), .CI(
        C[1004]), .S(S[1004]), .CO(C[1005]) );
  FA_2067 \FA_INST_0[1].FA_INST_1[493].FA_  ( .A(A[1005]), .B(B[1005]), .CI(
        C[1005]), .S(S[1005]), .CO(C[1006]) );
  FA_2066 \FA_INST_0[1].FA_INST_1[494].FA_  ( .A(A[1006]), .B(B[1006]), .CI(
        C[1006]), .S(S[1006]), .CO(C[1007]) );
  FA_2065 \FA_INST_0[1].FA_INST_1[495].FA_  ( .A(A[1007]), .B(B[1007]), .CI(
        C[1007]), .S(S[1007]), .CO(C[1008]) );
  FA_2064 \FA_INST_0[1].FA_INST_1[496].FA_  ( .A(A[1008]), .B(B[1008]), .CI(
        C[1008]), .S(S[1008]), .CO(C[1009]) );
  FA_2063 \FA_INST_0[1].FA_INST_1[497].FA_  ( .A(A[1009]), .B(B[1009]), .CI(
        C[1009]), .S(S[1009]), .CO(C[1010]) );
  FA_2062 \FA_INST_0[1].FA_INST_1[498].FA_  ( .A(A[1010]), .B(B[1010]), .CI(
        C[1010]), .S(S[1010]), .CO(C[1011]) );
  FA_2061 \FA_INST_0[1].FA_INST_1[499].FA_  ( .A(A[1011]), .B(B[1011]), .CI(
        C[1011]), .S(S[1011]), .CO(C[1012]) );
  FA_2060 \FA_INST_0[1].FA_INST_1[500].FA_  ( .A(A[1012]), .B(B[1012]), .CI(
        C[1012]), .S(S[1012]), .CO(C[1013]) );
  FA_2059 \FA_INST_0[1].FA_INST_1[501].FA_  ( .A(A[1013]), .B(B[1013]), .CI(
        C[1013]), .S(S[1013]), .CO(C[1014]) );
  FA_2058 \FA_INST_0[1].FA_INST_1[502].FA_  ( .A(A[1014]), .B(B[1014]), .CI(
        C[1014]), .S(S[1014]), .CO(C[1015]) );
  FA_2057 \FA_INST_0[1].FA_INST_1[503].FA_  ( .A(A[1015]), .B(B[1015]), .CI(
        C[1015]), .S(S[1015]), .CO(C[1016]) );
  FA_2056 \FA_INST_0[1].FA_INST_1[504].FA_  ( .A(A[1016]), .B(B[1016]), .CI(
        C[1016]), .S(S[1016]), .CO(C[1017]) );
  FA_2055 \FA_INST_0[1].FA_INST_1[505].FA_  ( .A(A[1017]), .B(B[1017]), .CI(
        C[1017]), .S(S[1017]), .CO(C[1018]) );
  FA_2054 \FA_INST_0[1].FA_INST_1[506].FA_  ( .A(A[1018]), .B(B[1018]), .CI(
        C[1018]), .S(S[1018]), .CO(C[1019]) );
  FA_2053 \FA_INST_0[1].FA_INST_1[507].FA_  ( .A(A[1019]), .B(B[1019]), .CI(
        C[1019]), .S(S[1019]), .CO(C[1020]) );
  FA_2052 \FA_INST_0[1].FA_INST_1[508].FA_  ( .A(1'b0), .B(B[1020]), .CI(
        C[1020]), .S(S[1020]), .CO(C[1021]) );
  FA_2051 \FA_INST_0[1].FA_INST_1[509].FA_  ( .A(1'b0), .B(B[1021]), .CI(
        C[1021]), .S(S[1021]), .CO(C[1022]) );
  FA_2050 \FA_INST_0[1].FA_INST_1[510].FA_  ( .A(1'b0), .B(B[1022]), .CI(
        C[1022]), .S(S[1022]) );
  FA_2049 \FA_INST_0[1].FA_INST_1[511].FA_  ( .A(1'b0), .B(B[1023]), .CI(1'b0), 
        .S(S[1023]) );
endmodule


module mult_N1024_CC256_DW01_add_0 ( A, B, CI, SUM, CO );
  input [1025:0] A;
  input [1025:0] B;
  output [1025:0] SUM;
  input CI;
  output CO;
  wire   \A[2] , \A[1] , \A[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
         n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
         n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
         n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
         n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
         n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
         n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
         n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
         n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
         n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
         n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
         n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
         n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
         n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
         n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
         n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
         n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
         n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
         n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
         n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
         n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
         n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
         n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
         n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
         n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
         n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
         n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
         n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
         n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
         n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
         n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
         n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
         n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
         n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
         n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
         n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
         n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
         n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
         n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
         n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
         n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
         n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
         n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
         n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
         n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
         n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
         n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
         n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
         n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
         n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
         n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
         n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
         n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
         n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
         n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968,
         n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
         n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
         n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998,
         n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008,
         n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018,
         n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028,
         n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
         n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
         n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058,
         n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068,
         n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078,
         n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088,
         n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098,
         n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108,
         n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
         n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
         n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
         n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
         n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
         n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
         n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
         n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
         n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
         n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
         n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
         n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
         n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
         n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
         n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
         n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
         n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
         n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
         n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
         n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
         n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
         n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
         n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
         n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358,
         n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368,
         n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378,
         n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388,
         n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398,
         n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408,
         n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418,
         n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428,
         n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438,
         n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448,
         n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458,
         n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468,
         n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478,
         n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488,
         n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498,
         n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508,
         n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518,
         n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528,
         n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
         n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
         n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
         n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
         n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
         n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
         n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
         n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
         n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
         n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
         n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
         n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
         n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
         n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
         n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678,
         n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688,
         n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698,
         n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
         n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
         n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728,
         n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
         n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748,
         n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
         n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768,
         n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778,
         n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788,
         n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798,
         n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808,
         n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818,
         n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828,
         n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838,
         n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848,
         n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858,
         n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868,
         n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878,
         n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888,
         n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
         n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908,
         n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918,
         n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928,
         n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938,
         n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948,
         n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958,
         n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968,
         n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978,
         n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988,
         n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
         n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008,
         n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018,
         n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
         n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
         n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048,
         n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
         n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
         n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
         n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
         n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
         n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
         n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
         n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
         n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
         n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
         n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
         n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
         n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
         n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
         n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
         n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
         n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
         n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
         n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
         n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
         n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
         n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
         n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
         n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
         n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
         n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
         n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
         n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
         n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
         n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
         n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
         n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
         n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
         n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
         n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438,
         n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
         n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458,
         n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468,
         n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478,
         n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488,
         n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
         n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
         n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
         n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
         n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
         n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
         n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
         n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
         n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
         n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
         n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598,
         n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
         n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618,
         n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
         n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
         n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
         n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
         n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
         n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
         n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
         n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
         n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
         n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
         n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728,
         n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738,
         n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748,
         n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
         n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
         n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
         n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
         n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
         n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
         n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
         n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
         n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
         n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
         n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
         n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
         n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
         n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
         n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
         n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
         n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
         n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
         n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
         n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258,
         n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268,
         n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
         n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
         n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
         n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
         n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318,
         n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
         n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338,
         n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
         n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
         n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
         n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
         n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388,
         n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398,
         n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408,
         n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418,
         n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428,
         n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438,
         n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
         n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458,
         n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468,
         n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478,
         n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488,
         n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498,
         n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508,
         n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518,
         n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
         n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
         n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
         n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
         n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568,
         n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578,
         n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588,
         n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598,
         n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608,
         n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
         n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
         n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
         n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
         n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
         n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
         n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
         n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
         n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698,
         n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708,
         n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718,
         n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
         n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
         n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
         n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
         n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
         n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
         n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788,
         n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798,
         n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808,
         n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818,
         n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828,
         n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838,
         n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848,
         n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858,
         n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868,
         n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878,
         n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888,
         n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898,
         n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908,
         n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918,
         n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928,
         n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938,
         n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948,
         n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958,
         n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968,
         n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978,
         n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988,
         n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998,
         n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008,
         n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018,
         n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028,
         n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038,
         n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048,
         n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058,
         n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068,
         n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078,
         n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088,
         n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098,
         n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108,
         n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118,
         n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128,
         n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138,
         n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148,
         n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158,
         n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168,
         n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178,
         n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188,
         n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198,
         n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208,
         n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218,
         n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228,
         n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238,
         n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248,
         n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258,
         n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268,
         n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278,
         n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
         n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298,
         n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308,
         n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318,
         n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
         n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
         n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348,
         n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
         n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
         n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378,
         n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
         n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398,
         n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408,
         n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418,
         n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428,
         n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
         n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448,
         n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458,
         n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468,
         n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478,
         n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
         n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
         n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
         n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
         n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
         n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
         n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
         n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
         n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
         n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
         n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
         n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
         n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608,
         n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
         n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
         n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
         n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
         n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
         n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
         n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
         n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
         n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
         n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
         n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
         n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
         n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
         n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
         n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
         n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
         n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
         n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
         n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
         n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
         n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
         n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
         n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858,
         n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
         n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878,
         n7879, n7880, n7881, n7882, n7883, n7884, n7885;
  assign SUM[2] = \A[2] ;
  assign \A[2]  = A[2];
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  NAND U2 ( .A(n27), .B(n30), .Z(n31) );
  XOR U3 ( .A(n1), .B(n2), .Z(SUM[9]) );
  NANDN U4 ( .A(n3), .B(n4), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[99]) );
  NANDN U6 ( .A(n7), .B(n8), .Z(n6) );
  ANDN U7 ( .B(n9), .A(n10), .Z(n5) );
  NAND U8 ( .A(n11), .B(n12), .Z(n9) );
  XOR U9 ( .A(n13), .B(n14), .Z(SUM[999]) );
  NANDN U10 ( .A(n15), .B(n16), .Z(n14) );
  ANDN U11 ( .B(n17), .A(n18), .Z(n13) );
  NAND U12 ( .A(n19), .B(n20), .Z(n17) );
  XNOR U13 ( .A(n19), .B(n21), .Z(SUM[998]) );
  NANDN U14 ( .A(n18), .B(n20), .Z(n21) );
  NANDN U15 ( .A(n22), .B(n23), .Z(n19) );
  NAND U16 ( .A(n24), .B(n25), .Z(n23) );
  XNOR U17 ( .A(n24), .B(n26), .Z(SUM[997]) );
  NANDN U18 ( .A(n22), .B(n25), .Z(n26) );
  NAND U19 ( .A(n27), .B(n28), .Z(n24) );
  NANDN U20 ( .A(n29), .B(n30), .Z(n28) );
  XOR U21 ( .A(n29), .B(n31), .Z(SUM[996]) );
  XOR U22 ( .A(n32), .B(n33), .Z(SUM[995]) );
  NANDN U23 ( .A(n34), .B(n35), .Z(n33) );
  ANDN U24 ( .B(n36), .A(n37), .Z(n32) );
  NAND U25 ( .A(n38), .B(n39), .Z(n36) );
  XNOR U26 ( .A(n38), .B(n40), .Z(SUM[994]) );
  NANDN U27 ( .A(n37), .B(n39), .Z(n40) );
  NANDN U28 ( .A(n41), .B(n42), .Z(n38) );
  NAND U29 ( .A(n43), .B(n44), .Z(n42) );
  XNOR U30 ( .A(n43), .B(n45), .Z(SUM[993]) );
  NANDN U31 ( .A(n41), .B(n44), .Z(n45) );
  NANDN U32 ( .A(n46), .B(n47), .Z(n43) );
  OR U33 ( .A(n48), .B(n49), .Z(n47) );
  XOR U34 ( .A(n48), .B(n50), .Z(SUM[992]) );
  OR U35 ( .A(n49), .B(n46), .Z(n50) );
  XOR U36 ( .A(n51), .B(n52), .Z(SUM[991]) );
  OR U37 ( .A(n53), .B(n54), .Z(n52) );
  ANDN U38 ( .B(n55), .A(n56), .Z(n51) );
  NANDN U39 ( .A(n57), .B(n58), .Z(n55) );
  XNOR U40 ( .A(n58), .B(n59), .Z(SUM[990]) );
  OR U41 ( .A(n57), .B(n56), .Z(n59) );
  NANDN U42 ( .A(n60), .B(n61), .Z(n58) );
  NANDN U43 ( .A(n62), .B(n63), .Z(n61) );
  XNOR U44 ( .A(n11), .B(n64), .Z(SUM[98]) );
  NANDN U45 ( .A(n10), .B(n12), .Z(n64) );
  NANDN U46 ( .A(n65), .B(n66), .Z(n11) );
  NAND U47 ( .A(n67), .B(n68), .Z(n66) );
  XNOR U48 ( .A(n63), .B(n69), .Z(SUM[989]) );
  OR U49 ( .A(n62), .B(n60), .Z(n69) );
  NANDN U50 ( .A(n70), .B(n71), .Z(n63) );
  NANDN U51 ( .A(n72), .B(n73), .Z(n71) );
  XNOR U52 ( .A(n73), .B(n74), .Z(SUM[988]) );
  OR U53 ( .A(n72), .B(n70), .Z(n74) );
  NANDN U54 ( .A(n75), .B(n76), .Z(n73) );
  NANDN U55 ( .A(n77), .B(n78), .Z(n76) );
  XOR U56 ( .A(n79), .B(n80), .Z(SUM[987]) );
  NANDN U57 ( .A(n81), .B(n82), .Z(n80) );
  ANDN U58 ( .B(n83), .A(n84), .Z(n79) );
  NAND U59 ( .A(n85), .B(n86), .Z(n83) );
  XNOR U60 ( .A(n85), .B(n87), .Z(SUM[986]) );
  NANDN U61 ( .A(n84), .B(n86), .Z(n87) );
  NANDN U62 ( .A(n88), .B(n89), .Z(n85) );
  NAND U63 ( .A(n90), .B(n91), .Z(n89) );
  XNOR U64 ( .A(n90), .B(n92), .Z(SUM[985]) );
  NANDN U65 ( .A(n88), .B(n91), .Z(n92) );
  NANDN U66 ( .A(n93), .B(n94), .Z(n90) );
  NAND U67 ( .A(n78), .B(n95), .Z(n94) );
  XNOR U68 ( .A(n78), .B(n96), .Z(SUM[984]) );
  NANDN U69 ( .A(n93), .B(n95), .Z(n96) );
  NANDN U70 ( .A(n97), .B(n98), .Z(n78) );
  OR U71 ( .A(n99), .B(n100), .Z(n98) );
  XOR U72 ( .A(n101), .B(n102), .Z(SUM[983]) );
  NANDN U73 ( .A(n103), .B(n104), .Z(n102) );
  ANDN U74 ( .B(n105), .A(n106), .Z(n101) );
  NAND U75 ( .A(n107), .B(n108), .Z(n105) );
  XNOR U76 ( .A(n107), .B(n109), .Z(SUM[982]) );
  NANDN U77 ( .A(n106), .B(n108), .Z(n109) );
  NANDN U78 ( .A(n110), .B(n111), .Z(n107) );
  NAND U79 ( .A(n112), .B(n113), .Z(n111) );
  XNOR U80 ( .A(n112), .B(n114), .Z(SUM[981]) );
  NANDN U81 ( .A(n110), .B(n113), .Z(n114) );
  NANDN U82 ( .A(n115), .B(n116), .Z(n112) );
  NANDN U83 ( .A(n100), .B(n117), .Z(n116) );
  XOR U84 ( .A(n100), .B(n118), .Z(SUM[980]) );
  NANDN U85 ( .A(n115), .B(n117), .Z(n118) );
  NOR U86 ( .A(n119), .B(n120), .Z(n100) );
  XNOR U87 ( .A(n67), .B(n121), .Z(SUM[97]) );
  NANDN U88 ( .A(n65), .B(n68), .Z(n121) );
  NANDN U89 ( .A(n122), .B(n123), .Z(n67) );
  OR U90 ( .A(n124), .B(n125), .Z(n123) );
  XOR U91 ( .A(n126), .B(n127), .Z(SUM[979]) );
  NANDN U92 ( .A(n128), .B(n129), .Z(n127) );
  ANDN U93 ( .B(n130), .A(n131), .Z(n126) );
  NAND U94 ( .A(n132), .B(n133), .Z(n130) );
  XNOR U95 ( .A(n132), .B(n134), .Z(SUM[978]) );
  NANDN U96 ( .A(n131), .B(n133), .Z(n134) );
  NANDN U97 ( .A(n135), .B(n136), .Z(n132) );
  NAND U98 ( .A(n137), .B(n138), .Z(n136) );
  XNOR U99 ( .A(n137), .B(n139), .Z(SUM[977]) );
  NANDN U100 ( .A(n135), .B(n138), .Z(n139) );
  NANDN U101 ( .A(n140), .B(n141), .Z(n137) );
  OR U102 ( .A(n142), .B(n143), .Z(n141) );
  XOR U103 ( .A(n142), .B(n144), .Z(SUM[976]) );
  OR U104 ( .A(n143), .B(n140), .Z(n144) );
  XOR U105 ( .A(n145), .B(n146), .Z(SUM[975]) );
  OR U106 ( .A(n147), .B(n148), .Z(n146) );
  ANDN U107 ( .B(n149), .A(n150), .Z(n145) );
  NANDN U108 ( .A(n151), .B(n152), .Z(n149) );
  XNOR U109 ( .A(n152), .B(n153), .Z(SUM[974]) );
  OR U110 ( .A(n151), .B(n150), .Z(n153) );
  NANDN U111 ( .A(n154), .B(n155), .Z(n152) );
  NANDN U112 ( .A(n156), .B(n157), .Z(n155) );
  XNOR U113 ( .A(n157), .B(n158), .Z(SUM[973]) );
  OR U114 ( .A(n156), .B(n154), .Z(n158) );
  NANDN U115 ( .A(n159), .B(n160), .Z(n157) );
  NANDN U116 ( .A(n161), .B(n162), .Z(n160) );
  XNOR U117 ( .A(n162), .B(n163), .Z(SUM[972]) );
  OR U118 ( .A(n161), .B(n159), .Z(n163) );
  NANDN U119 ( .A(n164), .B(n165), .Z(n162) );
  NANDN U120 ( .A(n166), .B(n167), .Z(n165) );
  XOR U121 ( .A(n168), .B(n169), .Z(SUM[971]) );
  NANDN U122 ( .A(n170), .B(n171), .Z(n169) );
  ANDN U123 ( .B(n172), .A(n173), .Z(n168) );
  NAND U124 ( .A(n174), .B(n175), .Z(n172) );
  XNOR U125 ( .A(n174), .B(n176), .Z(SUM[970]) );
  NANDN U126 ( .A(n173), .B(n175), .Z(n176) );
  NANDN U127 ( .A(n177), .B(n178), .Z(n174) );
  NAND U128 ( .A(n179), .B(n180), .Z(n178) );
  XOR U129 ( .A(n125), .B(n181), .Z(SUM[96]) );
  OR U130 ( .A(n124), .B(n122), .Z(n181) );
  XNOR U131 ( .A(n179), .B(n182), .Z(SUM[969]) );
  NANDN U132 ( .A(n177), .B(n180), .Z(n182) );
  NANDN U133 ( .A(n183), .B(n184), .Z(n179) );
  NAND U134 ( .A(n167), .B(n185), .Z(n184) );
  XNOR U135 ( .A(n167), .B(n186), .Z(SUM[968]) );
  NANDN U136 ( .A(n183), .B(n185), .Z(n186) );
  NANDN U137 ( .A(n187), .B(n188), .Z(n167) );
  OR U138 ( .A(n189), .B(n190), .Z(n188) );
  XOR U139 ( .A(n191), .B(n192), .Z(SUM[967]) );
  NANDN U140 ( .A(n193), .B(n194), .Z(n192) );
  ANDN U141 ( .B(n195), .A(n196), .Z(n191) );
  NAND U142 ( .A(n197), .B(n198), .Z(n195) );
  XNOR U143 ( .A(n197), .B(n199), .Z(SUM[966]) );
  NANDN U144 ( .A(n196), .B(n198), .Z(n199) );
  NANDN U145 ( .A(n200), .B(n201), .Z(n197) );
  NAND U146 ( .A(n202), .B(n203), .Z(n201) );
  XNOR U147 ( .A(n202), .B(n204), .Z(SUM[965]) );
  NANDN U148 ( .A(n200), .B(n203), .Z(n204) );
  NANDN U149 ( .A(n205), .B(n206), .Z(n202) );
  NANDN U150 ( .A(n190), .B(n207), .Z(n206) );
  XOR U151 ( .A(n190), .B(n208), .Z(SUM[964]) );
  NANDN U152 ( .A(n205), .B(n207), .Z(n208) );
  NOR U153 ( .A(n209), .B(n210), .Z(n190) );
  XOR U154 ( .A(n211), .B(n212), .Z(SUM[963]) );
  NANDN U155 ( .A(n213), .B(n214), .Z(n212) );
  ANDN U156 ( .B(n215), .A(n216), .Z(n211) );
  NAND U157 ( .A(n217), .B(n218), .Z(n215) );
  XNOR U158 ( .A(n217), .B(n219), .Z(SUM[962]) );
  NANDN U159 ( .A(n216), .B(n218), .Z(n219) );
  NANDN U160 ( .A(n220), .B(n221), .Z(n217) );
  NAND U161 ( .A(n222), .B(n223), .Z(n221) );
  XNOR U162 ( .A(n222), .B(n224), .Z(SUM[961]) );
  NANDN U163 ( .A(n220), .B(n223), .Z(n224) );
  NANDN U164 ( .A(n225), .B(n226), .Z(n222) );
  OR U165 ( .A(n227), .B(n228), .Z(n226) );
  XOR U166 ( .A(n227), .B(n229), .Z(SUM[960]) );
  OR U167 ( .A(n228), .B(n225), .Z(n229) );
  XOR U168 ( .A(n230), .B(n231), .Z(SUM[95]) );
  NANDN U169 ( .A(n232), .B(n233), .Z(n231) );
  ANDN U170 ( .B(n234), .A(n235), .Z(n230) );
  NANDN U171 ( .A(n236), .B(n237), .Z(n234) );
  XOR U172 ( .A(n238), .B(n239), .Z(SUM[959]) );
  OR U173 ( .A(n240), .B(n241), .Z(n239) );
  ANDN U174 ( .B(n242), .A(n243), .Z(n238) );
  NANDN U175 ( .A(n244), .B(n245), .Z(n242) );
  XNOR U176 ( .A(n245), .B(n246), .Z(SUM[958]) );
  OR U177 ( .A(n244), .B(n243), .Z(n246) );
  NANDN U178 ( .A(n247), .B(n248), .Z(n245) );
  NANDN U179 ( .A(n249), .B(n250), .Z(n248) );
  XNOR U180 ( .A(n250), .B(n251), .Z(SUM[957]) );
  OR U181 ( .A(n249), .B(n247), .Z(n251) );
  NANDN U182 ( .A(n252), .B(n253), .Z(n250) );
  NAND U183 ( .A(n254), .B(n255), .Z(n253) );
  XNOR U184 ( .A(n254), .B(n256), .Z(SUM[956]) );
  NANDN U185 ( .A(n252), .B(n255), .Z(n256) );
  NANDN U186 ( .A(n257), .B(n258), .Z(n254) );
  NANDN U187 ( .A(n259), .B(n260), .Z(n258) );
  XOR U188 ( .A(n261), .B(n262), .Z(SUM[955]) );
  NANDN U189 ( .A(n263), .B(n264), .Z(n262) );
  ANDN U190 ( .B(n265), .A(n266), .Z(n261) );
  NAND U191 ( .A(n267), .B(n268), .Z(n265) );
  XNOR U192 ( .A(n267), .B(n269), .Z(SUM[954]) );
  NANDN U193 ( .A(n266), .B(n268), .Z(n269) );
  NANDN U194 ( .A(n270), .B(n271), .Z(n267) );
  NAND U195 ( .A(n272), .B(n273), .Z(n271) );
  XNOR U196 ( .A(n272), .B(n274), .Z(SUM[953]) );
  NANDN U197 ( .A(n270), .B(n273), .Z(n274) );
  NANDN U198 ( .A(n275), .B(n276), .Z(n272) );
  NAND U199 ( .A(n260), .B(n277), .Z(n276) );
  XNOR U200 ( .A(n260), .B(n278), .Z(SUM[952]) );
  NANDN U201 ( .A(n275), .B(n277), .Z(n278) );
  NANDN U202 ( .A(n279), .B(n280), .Z(n260) );
  NANDN U203 ( .A(n281), .B(n282), .Z(n280) );
  XOR U204 ( .A(n283), .B(n284), .Z(SUM[951]) );
  NANDN U205 ( .A(n285), .B(n286), .Z(n284) );
  ANDN U206 ( .B(n287), .A(n288), .Z(n283) );
  NAND U207 ( .A(n289), .B(n290), .Z(n287) );
  XNOR U208 ( .A(n289), .B(n291), .Z(SUM[950]) );
  NANDN U209 ( .A(n288), .B(n290), .Z(n291) );
  NANDN U210 ( .A(n292), .B(n293), .Z(n289) );
  NAND U211 ( .A(n294), .B(n295), .Z(n293) );
  XNOR U212 ( .A(n237), .B(n296), .Z(SUM[94]) );
  OR U213 ( .A(n236), .B(n235), .Z(n296) );
  NANDN U214 ( .A(n297), .B(n298), .Z(n237) );
  NAND U215 ( .A(n299), .B(n300), .Z(n298) );
  XNOR U216 ( .A(n294), .B(n301), .Z(SUM[949]) );
  NANDN U217 ( .A(n292), .B(n295), .Z(n301) );
  NANDN U218 ( .A(n302), .B(n303), .Z(n294) );
  NANDN U219 ( .A(n281), .B(n304), .Z(n303) );
  XOR U220 ( .A(n281), .B(n305), .Z(SUM[948]) );
  NANDN U221 ( .A(n302), .B(n304), .Z(n305) );
  ANDN U222 ( .B(n306), .A(n307), .Z(n281) );
  OR U223 ( .A(n308), .B(n309), .Z(n306) );
  XOR U224 ( .A(n310), .B(n311), .Z(SUM[947]) );
  NANDN U225 ( .A(n312), .B(n313), .Z(n311) );
  ANDN U226 ( .B(n314), .A(n315), .Z(n310) );
  NANDN U227 ( .A(n316), .B(n317), .Z(n314) );
  XNOR U228 ( .A(n317), .B(n318), .Z(SUM[946]) );
  OR U229 ( .A(n316), .B(n315), .Z(n318) );
  NANDN U230 ( .A(n319), .B(n320), .Z(n317) );
  NAND U231 ( .A(n321), .B(n322), .Z(n320) );
  XNOR U232 ( .A(n321), .B(n323), .Z(SUM[945]) );
  NANDN U233 ( .A(n319), .B(n322), .Z(n323) );
  NANDN U234 ( .A(n324), .B(n325), .Z(n321) );
  NANDN U235 ( .A(n309), .B(n326), .Z(n325) );
  XOR U236 ( .A(n309), .B(n327), .Z(SUM[944]) );
  NANDN U237 ( .A(n324), .B(n326), .Z(n327) );
  XOR U238 ( .A(n328), .B(n329), .Z(SUM[943]) );
  OR U239 ( .A(n330), .B(n331), .Z(n329) );
  ANDN U240 ( .B(n332), .A(n333), .Z(n328) );
  NANDN U241 ( .A(n334), .B(n335), .Z(n332) );
  XNOR U242 ( .A(n335), .B(n336), .Z(SUM[942]) );
  OR U243 ( .A(n334), .B(n333), .Z(n336) );
  NANDN U244 ( .A(n337), .B(n338), .Z(n335) );
  NANDN U245 ( .A(n339), .B(n340), .Z(n338) );
  XNOR U246 ( .A(n340), .B(n341), .Z(SUM[941]) );
  OR U247 ( .A(n339), .B(n337), .Z(n341) );
  NANDN U248 ( .A(n342), .B(n343), .Z(n340) );
  NAND U249 ( .A(n344), .B(n345), .Z(n343) );
  XNOR U250 ( .A(n344), .B(n346), .Z(SUM[940]) );
  NANDN U251 ( .A(n342), .B(n345), .Z(n346) );
  NANDN U252 ( .A(n347), .B(n348), .Z(n344) );
  NANDN U253 ( .A(n349), .B(n350), .Z(n348) );
  XNOR U254 ( .A(n299), .B(n351), .Z(SUM[93]) );
  NANDN U255 ( .A(n297), .B(n300), .Z(n351) );
  NANDN U256 ( .A(n352), .B(n353), .Z(n299) );
  NANDN U257 ( .A(n354), .B(n355), .Z(n353) );
  XOR U258 ( .A(n356), .B(n357), .Z(SUM[939]) );
  NANDN U259 ( .A(n358), .B(n359), .Z(n357) );
  ANDN U260 ( .B(n360), .A(n361), .Z(n356) );
  NAND U261 ( .A(n362), .B(n363), .Z(n360) );
  XNOR U262 ( .A(n362), .B(n364), .Z(SUM[938]) );
  NANDN U263 ( .A(n361), .B(n363), .Z(n364) );
  NANDN U264 ( .A(n365), .B(n366), .Z(n362) );
  NAND U265 ( .A(n367), .B(n368), .Z(n366) );
  XNOR U266 ( .A(n367), .B(n369), .Z(SUM[937]) );
  NANDN U267 ( .A(n365), .B(n368), .Z(n369) );
  NANDN U268 ( .A(n370), .B(n371), .Z(n367) );
  NAND U269 ( .A(n350), .B(n372), .Z(n371) );
  XNOR U270 ( .A(n350), .B(n373), .Z(SUM[936]) );
  NANDN U271 ( .A(n370), .B(n372), .Z(n373) );
  NANDN U272 ( .A(n374), .B(n375), .Z(n350) );
  NANDN U273 ( .A(n376), .B(n377), .Z(n375) );
  XOR U274 ( .A(n378), .B(n379), .Z(SUM[935]) );
  NANDN U275 ( .A(n380), .B(n381), .Z(n379) );
  ANDN U276 ( .B(n382), .A(n383), .Z(n378) );
  NAND U277 ( .A(n384), .B(n385), .Z(n382) );
  XNOR U278 ( .A(n384), .B(n386), .Z(SUM[934]) );
  NANDN U279 ( .A(n383), .B(n385), .Z(n386) );
  NANDN U280 ( .A(n387), .B(n388), .Z(n384) );
  NAND U281 ( .A(n389), .B(n390), .Z(n388) );
  XNOR U282 ( .A(n389), .B(n391), .Z(SUM[933]) );
  NANDN U283 ( .A(n387), .B(n390), .Z(n391) );
  NANDN U284 ( .A(n392), .B(n393), .Z(n389) );
  NANDN U285 ( .A(n376), .B(n394), .Z(n393) );
  XOR U286 ( .A(n376), .B(n395), .Z(SUM[932]) );
  NANDN U287 ( .A(n392), .B(n394), .Z(n395) );
  ANDN U288 ( .B(n396), .A(n397), .Z(n376) );
  OR U289 ( .A(n398), .B(n399), .Z(n396) );
  XOR U290 ( .A(n400), .B(n401), .Z(SUM[931]) );
  NANDN U291 ( .A(n402), .B(n403), .Z(n401) );
  ANDN U292 ( .B(n404), .A(n405), .Z(n400) );
  NANDN U293 ( .A(n406), .B(n407), .Z(n404) );
  XNOR U294 ( .A(n407), .B(n408), .Z(SUM[930]) );
  OR U295 ( .A(n406), .B(n405), .Z(n408) );
  NANDN U296 ( .A(n409), .B(n410), .Z(n407) );
  NAND U297 ( .A(n411), .B(n412), .Z(n410) );
  XNOR U298 ( .A(n355), .B(n413), .Z(SUM[92]) );
  OR U299 ( .A(n354), .B(n352), .Z(n413) );
  NANDN U300 ( .A(n414), .B(n415), .Z(n355) );
  NANDN U301 ( .A(n416), .B(n417), .Z(n415) );
  XNOR U302 ( .A(n411), .B(n418), .Z(SUM[929]) );
  NANDN U303 ( .A(n409), .B(n412), .Z(n418) );
  NANDN U304 ( .A(n419), .B(n420), .Z(n411) );
  NANDN U305 ( .A(n399), .B(n421), .Z(n420) );
  XOR U306 ( .A(n399), .B(n422), .Z(SUM[928]) );
  NANDN U307 ( .A(n419), .B(n421), .Z(n422) );
  XOR U308 ( .A(n423), .B(n424), .Z(SUM[927]) );
  OR U309 ( .A(n425), .B(n426), .Z(n424) );
  ANDN U310 ( .B(n427), .A(n428), .Z(n423) );
  NANDN U311 ( .A(n429), .B(n430), .Z(n427) );
  XNOR U312 ( .A(n430), .B(n431), .Z(SUM[926]) );
  OR U313 ( .A(n429), .B(n428), .Z(n431) );
  NANDN U314 ( .A(n432), .B(n433), .Z(n430) );
  NANDN U315 ( .A(n434), .B(n435), .Z(n433) );
  XNOR U316 ( .A(n435), .B(n436), .Z(SUM[925]) );
  OR U317 ( .A(n434), .B(n432), .Z(n436) );
  NANDN U318 ( .A(n437), .B(n438), .Z(n435) );
  NAND U319 ( .A(n439), .B(n440), .Z(n438) );
  XNOR U320 ( .A(n439), .B(n441), .Z(SUM[924]) );
  NANDN U321 ( .A(n437), .B(n440), .Z(n441) );
  NANDN U322 ( .A(n442), .B(n443), .Z(n439) );
  NANDN U323 ( .A(n444), .B(n445), .Z(n443) );
  XOR U324 ( .A(n446), .B(n447), .Z(SUM[923]) );
  NANDN U325 ( .A(n448), .B(n449), .Z(n447) );
  ANDN U326 ( .B(n450), .A(n451), .Z(n446) );
  NAND U327 ( .A(n452), .B(n453), .Z(n450) );
  XNOR U328 ( .A(n452), .B(n454), .Z(SUM[922]) );
  NANDN U329 ( .A(n451), .B(n453), .Z(n454) );
  NANDN U330 ( .A(n455), .B(n456), .Z(n452) );
  NAND U331 ( .A(n457), .B(n458), .Z(n456) );
  XNOR U332 ( .A(n457), .B(n459), .Z(SUM[921]) );
  NANDN U333 ( .A(n455), .B(n458), .Z(n459) );
  NANDN U334 ( .A(n460), .B(n461), .Z(n457) );
  NAND U335 ( .A(n445), .B(n462), .Z(n461) );
  XNOR U336 ( .A(n445), .B(n463), .Z(SUM[920]) );
  NANDN U337 ( .A(n460), .B(n462), .Z(n463) );
  NANDN U338 ( .A(n464), .B(n465), .Z(n445) );
  NANDN U339 ( .A(n466), .B(n467), .Z(n465) );
  XOR U340 ( .A(n468), .B(n469), .Z(SUM[91]) );
  NANDN U341 ( .A(n470), .B(n471), .Z(n469) );
  ANDN U342 ( .B(n472), .A(n473), .Z(n468) );
  NAND U343 ( .A(n474), .B(n475), .Z(n472) );
  XOR U344 ( .A(n476), .B(n477), .Z(SUM[919]) );
  NANDN U345 ( .A(n478), .B(n479), .Z(n477) );
  ANDN U346 ( .B(n480), .A(n481), .Z(n476) );
  NAND U347 ( .A(n482), .B(n483), .Z(n480) );
  XNOR U348 ( .A(n482), .B(n484), .Z(SUM[918]) );
  NANDN U349 ( .A(n481), .B(n483), .Z(n484) );
  NANDN U350 ( .A(n485), .B(n486), .Z(n482) );
  NAND U351 ( .A(n487), .B(n488), .Z(n486) );
  XNOR U352 ( .A(n487), .B(n489), .Z(SUM[917]) );
  NANDN U353 ( .A(n485), .B(n488), .Z(n489) );
  NANDN U354 ( .A(n490), .B(n491), .Z(n487) );
  NANDN U355 ( .A(n466), .B(n492), .Z(n491) );
  XOR U356 ( .A(n466), .B(n493), .Z(SUM[916]) );
  NANDN U357 ( .A(n490), .B(n492), .Z(n493) );
  ANDN U358 ( .B(n494), .A(n495), .Z(n466) );
  OR U359 ( .A(n496), .B(n497), .Z(n494) );
  XOR U360 ( .A(n498), .B(n499), .Z(SUM[915]) );
  NANDN U361 ( .A(n500), .B(n501), .Z(n499) );
  ANDN U362 ( .B(n502), .A(n503), .Z(n498) );
  NANDN U363 ( .A(n504), .B(n505), .Z(n502) );
  XNOR U364 ( .A(n505), .B(n506), .Z(SUM[914]) );
  OR U365 ( .A(n504), .B(n503), .Z(n506) );
  NANDN U366 ( .A(n507), .B(n508), .Z(n505) );
  NAND U367 ( .A(n509), .B(n510), .Z(n508) );
  XNOR U368 ( .A(n509), .B(n511), .Z(SUM[913]) );
  NANDN U369 ( .A(n507), .B(n510), .Z(n511) );
  NANDN U370 ( .A(n512), .B(n513), .Z(n509) );
  NANDN U371 ( .A(n497), .B(n514), .Z(n513) );
  XOR U372 ( .A(n497), .B(n515), .Z(SUM[912]) );
  NANDN U373 ( .A(n512), .B(n514), .Z(n515) );
  XOR U374 ( .A(n516), .B(n517), .Z(SUM[911]) );
  OR U375 ( .A(n518), .B(n519), .Z(n517) );
  ANDN U376 ( .B(n520), .A(n521), .Z(n516) );
  NANDN U377 ( .A(n522), .B(n523), .Z(n520) );
  XNOR U378 ( .A(n523), .B(n524), .Z(SUM[910]) );
  OR U379 ( .A(n522), .B(n521), .Z(n524) );
  NANDN U380 ( .A(n525), .B(n526), .Z(n523) );
  NANDN U381 ( .A(n527), .B(n528), .Z(n526) );
  XNOR U382 ( .A(n474), .B(n529), .Z(SUM[90]) );
  NANDN U383 ( .A(n473), .B(n475), .Z(n529) );
  NANDN U384 ( .A(n530), .B(n531), .Z(n474) );
  NAND U385 ( .A(n532), .B(n533), .Z(n531) );
  XNOR U386 ( .A(n528), .B(n534), .Z(SUM[909]) );
  OR U387 ( .A(n527), .B(n525), .Z(n534) );
  NANDN U388 ( .A(n535), .B(n536), .Z(n528) );
  NAND U389 ( .A(n537), .B(n538), .Z(n536) );
  XNOR U390 ( .A(n537), .B(n539), .Z(SUM[908]) );
  NANDN U391 ( .A(n535), .B(n538), .Z(n539) );
  NANDN U392 ( .A(n540), .B(n541), .Z(n537) );
  NANDN U393 ( .A(n542), .B(n543), .Z(n541) );
  XOR U394 ( .A(n544), .B(n545), .Z(SUM[907]) );
  NANDN U395 ( .A(n546), .B(n547), .Z(n545) );
  ANDN U396 ( .B(n548), .A(n549), .Z(n544) );
  NAND U397 ( .A(n550), .B(n551), .Z(n548) );
  XNOR U398 ( .A(n550), .B(n552), .Z(SUM[906]) );
  NANDN U399 ( .A(n549), .B(n551), .Z(n552) );
  NANDN U400 ( .A(n553), .B(n554), .Z(n550) );
  NAND U401 ( .A(n555), .B(n556), .Z(n554) );
  XNOR U402 ( .A(n555), .B(n557), .Z(SUM[905]) );
  NANDN U403 ( .A(n553), .B(n556), .Z(n557) );
  NANDN U404 ( .A(n558), .B(n559), .Z(n555) );
  NAND U405 ( .A(n543), .B(n560), .Z(n559) );
  XNOR U406 ( .A(n543), .B(n561), .Z(SUM[904]) );
  NANDN U407 ( .A(n558), .B(n560), .Z(n561) );
  NANDN U408 ( .A(n562), .B(n563), .Z(n543) );
  NANDN U409 ( .A(n564), .B(n565), .Z(n563) );
  XOR U410 ( .A(n566), .B(n567), .Z(SUM[903]) );
  NANDN U411 ( .A(n568), .B(n569), .Z(n567) );
  ANDN U412 ( .B(n570), .A(n571), .Z(n566) );
  NAND U413 ( .A(n572), .B(n573), .Z(n570) );
  XNOR U414 ( .A(n572), .B(n574), .Z(SUM[902]) );
  NANDN U415 ( .A(n571), .B(n573), .Z(n574) );
  NANDN U416 ( .A(n575), .B(n576), .Z(n572) );
  NAND U417 ( .A(n577), .B(n578), .Z(n576) );
  XNOR U418 ( .A(n577), .B(n579), .Z(SUM[901]) );
  NANDN U419 ( .A(n575), .B(n578), .Z(n579) );
  NANDN U420 ( .A(n580), .B(n581), .Z(n577) );
  NANDN U421 ( .A(n564), .B(n582), .Z(n581) );
  XOR U422 ( .A(n564), .B(n583), .Z(SUM[900]) );
  NANDN U423 ( .A(n580), .B(n582), .Z(n583) );
  ANDN U424 ( .B(n584), .A(n585), .Z(n564) );
  OR U425 ( .A(n586), .B(n587), .Z(n584) );
  XOR U426 ( .A(n588), .B(n589), .Z(SUM[8]) );
  OR U427 ( .A(n590), .B(n591), .Z(n589) );
  XNOR U428 ( .A(n532), .B(n592), .Z(SUM[89]) );
  NANDN U429 ( .A(n530), .B(n533), .Z(n592) );
  NANDN U430 ( .A(n593), .B(n594), .Z(n532) );
  NAND U431 ( .A(n417), .B(n595), .Z(n594) );
  XOR U432 ( .A(n596), .B(n597), .Z(SUM[899]) );
  NANDN U433 ( .A(n598), .B(n599), .Z(n597) );
  ANDN U434 ( .B(n600), .A(n601), .Z(n596) );
  NANDN U435 ( .A(n602), .B(n603), .Z(n600) );
  XNOR U436 ( .A(n603), .B(n604), .Z(SUM[898]) );
  OR U437 ( .A(n602), .B(n601), .Z(n604) );
  NANDN U438 ( .A(n605), .B(n606), .Z(n603) );
  NAND U439 ( .A(n607), .B(n608), .Z(n606) );
  XNOR U440 ( .A(n607), .B(n609), .Z(SUM[897]) );
  NANDN U441 ( .A(n605), .B(n608), .Z(n609) );
  NANDN U442 ( .A(n610), .B(n611), .Z(n607) );
  NANDN U443 ( .A(n587), .B(n612), .Z(n611) );
  XOR U444 ( .A(n587), .B(n613), .Z(SUM[896]) );
  NANDN U445 ( .A(n610), .B(n612), .Z(n613) );
  XOR U446 ( .A(n614), .B(n615), .Z(SUM[895]) );
  OR U447 ( .A(n616), .B(n617), .Z(n615) );
  ANDN U448 ( .B(n618), .A(n619), .Z(n614) );
  NANDN U449 ( .A(n620), .B(n621), .Z(n618) );
  XNOR U450 ( .A(n621), .B(n622), .Z(SUM[894]) );
  OR U451 ( .A(n620), .B(n619), .Z(n622) );
  NANDN U452 ( .A(n623), .B(n624), .Z(n621) );
  NANDN U453 ( .A(n625), .B(n626), .Z(n624) );
  XNOR U454 ( .A(n626), .B(n627), .Z(SUM[893]) );
  OR U455 ( .A(n625), .B(n623), .Z(n627) );
  NANDN U456 ( .A(n628), .B(n629), .Z(n626) );
  NAND U457 ( .A(n630), .B(n631), .Z(n629) );
  XNOR U458 ( .A(n630), .B(n632), .Z(SUM[892]) );
  NANDN U459 ( .A(n628), .B(n631), .Z(n632) );
  NANDN U460 ( .A(n633), .B(n634), .Z(n630) );
  NANDN U461 ( .A(n635), .B(n636), .Z(n634) );
  XOR U462 ( .A(n637), .B(n638), .Z(SUM[891]) );
  NANDN U463 ( .A(n639), .B(n640), .Z(n638) );
  ANDN U464 ( .B(n641), .A(n642), .Z(n637) );
  NAND U465 ( .A(n643), .B(n644), .Z(n641) );
  XNOR U466 ( .A(n643), .B(n645), .Z(SUM[890]) );
  NANDN U467 ( .A(n642), .B(n644), .Z(n645) );
  NANDN U468 ( .A(n646), .B(n647), .Z(n643) );
  NAND U469 ( .A(n648), .B(n649), .Z(n647) );
  XNOR U470 ( .A(n417), .B(n650), .Z(SUM[88]) );
  NANDN U471 ( .A(n593), .B(n595), .Z(n650) );
  NANDN U472 ( .A(n651), .B(n652), .Z(n417) );
  NANDN U473 ( .A(n653), .B(n654), .Z(n652) );
  XNOR U474 ( .A(n648), .B(n655), .Z(SUM[889]) );
  NANDN U475 ( .A(n646), .B(n649), .Z(n655) );
  NANDN U476 ( .A(n656), .B(n657), .Z(n648) );
  NAND U477 ( .A(n636), .B(n658), .Z(n657) );
  XNOR U478 ( .A(n636), .B(n659), .Z(SUM[888]) );
  NANDN U479 ( .A(n656), .B(n658), .Z(n659) );
  NANDN U480 ( .A(n660), .B(n661), .Z(n636) );
  NANDN U481 ( .A(n662), .B(n663), .Z(n661) );
  XOR U482 ( .A(n664), .B(n665), .Z(SUM[887]) );
  NANDN U483 ( .A(n666), .B(n667), .Z(n665) );
  ANDN U484 ( .B(n668), .A(n669), .Z(n664) );
  NAND U485 ( .A(n670), .B(n671), .Z(n668) );
  XNOR U486 ( .A(n670), .B(n672), .Z(SUM[886]) );
  NANDN U487 ( .A(n669), .B(n671), .Z(n672) );
  NANDN U488 ( .A(n673), .B(n674), .Z(n670) );
  NAND U489 ( .A(n675), .B(n676), .Z(n674) );
  XNOR U490 ( .A(n675), .B(n677), .Z(SUM[885]) );
  NANDN U491 ( .A(n673), .B(n676), .Z(n677) );
  NANDN U492 ( .A(n678), .B(n679), .Z(n675) );
  NANDN U493 ( .A(n662), .B(n680), .Z(n679) );
  XOR U494 ( .A(n662), .B(n681), .Z(SUM[884]) );
  NANDN U495 ( .A(n678), .B(n680), .Z(n681) );
  ANDN U496 ( .B(n682), .A(n683), .Z(n662) );
  OR U497 ( .A(n684), .B(n685), .Z(n682) );
  XOR U498 ( .A(n686), .B(n687), .Z(SUM[883]) );
  NANDN U499 ( .A(n688), .B(n689), .Z(n687) );
  ANDN U500 ( .B(n690), .A(n691), .Z(n686) );
  NANDN U501 ( .A(n692), .B(n693), .Z(n690) );
  XNOR U502 ( .A(n693), .B(n694), .Z(SUM[882]) );
  OR U503 ( .A(n692), .B(n691), .Z(n694) );
  NANDN U504 ( .A(n695), .B(n696), .Z(n693) );
  NAND U505 ( .A(n697), .B(n698), .Z(n696) );
  XNOR U506 ( .A(n697), .B(n699), .Z(SUM[881]) );
  NANDN U507 ( .A(n695), .B(n698), .Z(n699) );
  NANDN U508 ( .A(n700), .B(n701), .Z(n697) );
  NANDN U509 ( .A(n685), .B(n702), .Z(n701) );
  XOR U510 ( .A(n685), .B(n703), .Z(SUM[880]) );
  NANDN U511 ( .A(n700), .B(n702), .Z(n703) );
  XOR U512 ( .A(n704), .B(n705), .Z(SUM[87]) );
  NANDN U513 ( .A(n706), .B(n707), .Z(n705) );
  ANDN U514 ( .B(n708), .A(n709), .Z(n704) );
  NAND U515 ( .A(n710), .B(n711), .Z(n708) );
  XOR U516 ( .A(n712), .B(n713), .Z(SUM[879]) );
  OR U517 ( .A(n714), .B(n715), .Z(n713) );
  ANDN U518 ( .B(n716), .A(n717), .Z(n712) );
  NANDN U519 ( .A(n718), .B(n719), .Z(n716) );
  XNOR U520 ( .A(n719), .B(n720), .Z(SUM[878]) );
  OR U521 ( .A(n718), .B(n717), .Z(n720) );
  NANDN U522 ( .A(n721), .B(n722), .Z(n719) );
  NANDN U523 ( .A(n723), .B(n724), .Z(n722) );
  XNOR U524 ( .A(n724), .B(n725), .Z(SUM[877]) );
  OR U525 ( .A(n723), .B(n721), .Z(n725) );
  NANDN U526 ( .A(n726), .B(n727), .Z(n724) );
  NAND U527 ( .A(n728), .B(n729), .Z(n727) );
  XNOR U528 ( .A(n728), .B(n730), .Z(SUM[876]) );
  NANDN U529 ( .A(n726), .B(n729), .Z(n730) );
  NANDN U530 ( .A(n731), .B(n732), .Z(n728) );
  NANDN U531 ( .A(n733), .B(n734), .Z(n732) );
  XOR U532 ( .A(n735), .B(n736), .Z(SUM[875]) );
  NANDN U533 ( .A(n737), .B(n738), .Z(n736) );
  ANDN U534 ( .B(n739), .A(n740), .Z(n735) );
  NAND U535 ( .A(n741), .B(n742), .Z(n739) );
  XNOR U536 ( .A(n741), .B(n743), .Z(SUM[874]) );
  NANDN U537 ( .A(n740), .B(n742), .Z(n743) );
  NANDN U538 ( .A(n744), .B(n745), .Z(n741) );
  NAND U539 ( .A(n746), .B(n747), .Z(n745) );
  XNOR U540 ( .A(n746), .B(n748), .Z(SUM[873]) );
  NANDN U541 ( .A(n744), .B(n747), .Z(n748) );
  NANDN U542 ( .A(n749), .B(n750), .Z(n746) );
  NAND U543 ( .A(n734), .B(n751), .Z(n750) );
  XNOR U544 ( .A(n734), .B(n752), .Z(SUM[872]) );
  NANDN U545 ( .A(n749), .B(n751), .Z(n752) );
  NANDN U546 ( .A(n753), .B(n754), .Z(n734) );
  NANDN U547 ( .A(n755), .B(n756), .Z(n754) );
  XOR U548 ( .A(n757), .B(n758), .Z(SUM[871]) );
  NANDN U549 ( .A(n759), .B(n760), .Z(n758) );
  ANDN U550 ( .B(n761), .A(n762), .Z(n757) );
  NAND U551 ( .A(n763), .B(n764), .Z(n761) );
  XNOR U552 ( .A(n763), .B(n765), .Z(SUM[870]) );
  NANDN U553 ( .A(n762), .B(n764), .Z(n765) );
  NANDN U554 ( .A(n766), .B(n767), .Z(n763) );
  NAND U555 ( .A(n768), .B(n769), .Z(n767) );
  XNOR U556 ( .A(n710), .B(n770), .Z(SUM[86]) );
  NANDN U557 ( .A(n709), .B(n711), .Z(n770) );
  NANDN U558 ( .A(n771), .B(n772), .Z(n710) );
  NAND U559 ( .A(n773), .B(n774), .Z(n772) );
  XNOR U560 ( .A(n768), .B(n775), .Z(SUM[869]) );
  NANDN U561 ( .A(n766), .B(n769), .Z(n775) );
  NANDN U562 ( .A(n776), .B(n777), .Z(n768) );
  NANDN U563 ( .A(n755), .B(n778), .Z(n777) );
  XOR U564 ( .A(n755), .B(n779), .Z(SUM[868]) );
  NANDN U565 ( .A(n776), .B(n778), .Z(n779) );
  ANDN U566 ( .B(n780), .A(n781), .Z(n755) );
  OR U567 ( .A(n782), .B(n783), .Z(n780) );
  XOR U568 ( .A(n784), .B(n785), .Z(SUM[867]) );
  NANDN U569 ( .A(n786), .B(n787), .Z(n785) );
  ANDN U570 ( .B(n788), .A(n789), .Z(n784) );
  NANDN U571 ( .A(n790), .B(n791), .Z(n788) );
  XNOR U572 ( .A(n791), .B(n792), .Z(SUM[866]) );
  OR U573 ( .A(n790), .B(n789), .Z(n792) );
  NANDN U574 ( .A(n793), .B(n794), .Z(n791) );
  NAND U575 ( .A(n795), .B(n796), .Z(n794) );
  XNOR U576 ( .A(n795), .B(n797), .Z(SUM[865]) );
  NANDN U577 ( .A(n793), .B(n796), .Z(n797) );
  NANDN U578 ( .A(n798), .B(n799), .Z(n795) );
  NANDN U579 ( .A(n783), .B(n800), .Z(n799) );
  XOR U580 ( .A(n783), .B(n801), .Z(SUM[864]) );
  NANDN U581 ( .A(n798), .B(n800), .Z(n801) );
  XOR U582 ( .A(n802), .B(n803), .Z(SUM[863]) );
  OR U583 ( .A(n804), .B(n805), .Z(n803) );
  ANDN U584 ( .B(n806), .A(n807), .Z(n802) );
  NANDN U585 ( .A(n808), .B(n809), .Z(n806) );
  XNOR U586 ( .A(n809), .B(n810), .Z(SUM[862]) );
  OR U587 ( .A(n808), .B(n807), .Z(n810) );
  NANDN U588 ( .A(n811), .B(n812), .Z(n809) );
  NANDN U589 ( .A(n813), .B(n814), .Z(n812) );
  XNOR U590 ( .A(n814), .B(n815), .Z(SUM[861]) );
  OR U591 ( .A(n813), .B(n811), .Z(n815) );
  NANDN U592 ( .A(n816), .B(n817), .Z(n814) );
  NAND U593 ( .A(n818), .B(n819), .Z(n817) );
  XNOR U594 ( .A(n818), .B(n820), .Z(SUM[860]) );
  NANDN U595 ( .A(n816), .B(n819), .Z(n820) );
  NANDN U596 ( .A(n821), .B(n822), .Z(n818) );
  NANDN U597 ( .A(n823), .B(n824), .Z(n822) );
  XNOR U598 ( .A(n773), .B(n825), .Z(SUM[85]) );
  NANDN U599 ( .A(n771), .B(n774), .Z(n825) );
  NANDN U600 ( .A(n826), .B(n827), .Z(n773) );
  NANDN U601 ( .A(n653), .B(n828), .Z(n827) );
  XOR U602 ( .A(n829), .B(n830), .Z(SUM[859]) );
  NANDN U603 ( .A(n831), .B(n832), .Z(n830) );
  ANDN U604 ( .B(n833), .A(n834), .Z(n829) );
  NAND U605 ( .A(n835), .B(n836), .Z(n833) );
  XNOR U606 ( .A(n835), .B(n837), .Z(SUM[858]) );
  NANDN U607 ( .A(n834), .B(n836), .Z(n837) );
  NANDN U608 ( .A(n838), .B(n839), .Z(n835) );
  NAND U609 ( .A(n840), .B(n841), .Z(n839) );
  XNOR U610 ( .A(n840), .B(n842), .Z(SUM[857]) );
  NANDN U611 ( .A(n838), .B(n841), .Z(n842) );
  NANDN U612 ( .A(n843), .B(n844), .Z(n840) );
  NAND U613 ( .A(n824), .B(n845), .Z(n844) );
  XNOR U614 ( .A(n824), .B(n846), .Z(SUM[856]) );
  NANDN U615 ( .A(n843), .B(n845), .Z(n846) );
  NANDN U616 ( .A(n847), .B(n848), .Z(n824) );
  NANDN U617 ( .A(n849), .B(n850), .Z(n848) );
  XOR U618 ( .A(n851), .B(n852), .Z(SUM[855]) );
  NANDN U619 ( .A(n853), .B(n854), .Z(n852) );
  ANDN U620 ( .B(n855), .A(n856), .Z(n851) );
  NAND U621 ( .A(n857), .B(n858), .Z(n855) );
  XNOR U622 ( .A(n857), .B(n859), .Z(SUM[854]) );
  NANDN U623 ( .A(n856), .B(n858), .Z(n859) );
  NANDN U624 ( .A(n860), .B(n861), .Z(n857) );
  NAND U625 ( .A(n862), .B(n863), .Z(n861) );
  XNOR U626 ( .A(n862), .B(n864), .Z(SUM[853]) );
  NANDN U627 ( .A(n860), .B(n863), .Z(n864) );
  NANDN U628 ( .A(n865), .B(n866), .Z(n862) );
  NANDN U629 ( .A(n849), .B(n867), .Z(n866) );
  XOR U630 ( .A(n849), .B(n868), .Z(SUM[852]) );
  NANDN U631 ( .A(n865), .B(n867), .Z(n868) );
  ANDN U632 ( .B(n869), .A(n870), .Z(n849) );
  OR U633 ( .A(n871), .B(n872), .Z(n869) );
  XOR U634 ( .A(n873), .B(n874), .Z(SUM[851]) );
  NANDN U635 ( .A(n875), .B(n876), .Z(n874) );
  ANDN U636 ( .B(n877), .A(n878), .Z(n873) );
  NANDN U637 ( .A(n879), .B(n880), .Z(n877) );
  XNOR U638 ( .A(n880), .B(n881), .Z(SUM[850]) );
  OR U639 ( .A(n879), .B(n878), .Z(n881) );
  NANDN U640 ( .A(n882), .B(n883), .Z(n880) );
  NAND U641 ( .A(n884), .B(n885), .Z(n883) );
  XOR U642 ( .A(n653), .B(n886), .Z(SUM[84]) );
  NANDN U643 ( .A(n826), .B(n828), .Z(n886) );
  ANDN U644 ( .B(n887), .A(n888), .Z(n653) );
  OR U645 ( .A(n889), .B(n890), .Z(n887) );
  XNOR U646 ( .A(n884), .B(n891), .Z(SUM[849]) );
  NANDN U647 ( .A(n882), .B(n885), .Z(n891) );
  NANDN U648 ( .A(n892), .B(n893), .Z(n884) );
  NANDN U649 ( .A(n872), .B(n894), .Z(n893) );
  XOR U650 ( .A(n872), .B(n895), .Z(SUM[848]) );
  NANDN U651 ( .A(n892), .B(n894), .Z(n895) );
  XOR U652 ( .A(n896), .B(n897), .Z(SUM[847]) );
  OR U653 ( .A(n898), .B(n899), .Z(n897) );
  ANDN U654 ( .B(n900), .A(n901), .Z(n896) );
  NANDN U655 ( .A(n902), .B(n903), .Z(n900) );
  XNOR U656 ( .A(n903), .B(n904), .Z(SUM[846]) );
  OR U657 ( .A(n902), .B(n901), .Z(n904) );
  NANDN U658 ( .A(n905), .B(n906), .Z(n903) );
  NANDN U659 ( .A(n907), .B(n908), .Z(n906) );
  XNOR U660 ( .A(n908), .B(n909), .Z(SUM[845]) );
  OR U661 ( .A(n907), .B(n905), .Z(n909) );
  NANDN U662 ( .A(n910), .B(n911), .Z(n908) );
  NAND U663 ( .A(n912), .B(n913), .Z(n911) );
  XNOR U664 ( .A(n912), .B(n914), .Z(SUM[844]) );
  NANDN U665 ( .A(n910), .B(n913), .Z(n914) );
  NANDN U666 ( .A(n915), .B(n916), .Z(n912) );
  NANDN U667 ( .A(n917), .B(n918), .Z(n916) );
  XOR U668 ( .A(n919), .B(n920), .Z(SUM[843]) );
  NANDN U669 ( .A(n921), .B(n922), .Z(n920) );
  ANDN U670 ( .B(n923), .A(n924), .Z(n919) );
  NAND U671 ( .A(n925), .B(n926), .Z(n923) );
  XNOR U672 ( .A(n925), .B(n927), .Z(SUM[842]) );
  NANDN U673 ( .A(n924), .B(n926), .Z(n927) );
  NANDN U674 ( .A(n928), .B(n929), .Z(n925) );
  NAND U675 ( .A(n930), .B(n931), .Z(n929) );
  XNOR U676 ( .A(n930), .B(n932), .Z(SUM[841]) );
  NANDN U677 ( .A(n928), .B(n931), .Z(n932) );
  NANDN U678 ( .A(n933), .B(n934), .Z(n930) );
  NAND U679 ( .A(n918), .B(n935), .Z(n934) );
  XNOR U680 ( .A(n918), .B(n936), .Z(SUM[840]) );
  NANDN U681 ( .A(n933), .B(n935), .Z(n936) );
  NANDN U682 ( .A(n937), .B(n938), .Z(n918) );
  NANDN U683 ( .A(n939), .B(n940), .Z(n938) );
  XOR U684 ( .A(n941), .B(n942), .Z(SUM[83]) );
  NANDN U685 ( .A(n943), .B(n944), .Z(n942) );
  ANDN U686 ( .B(n945), .A(n946), .Z(n941) );
  NANDN U687 ( .A(n947), .B(n948), .Z(n945) );
  XOR U688 ( .A(n949), .B(n950), .Z(SUM[839]) );
  NANDN U689 ( .A(n951), .B(n952), .Z(n950) );
  ANDN U690 ( .B(n953), .A(n954), .Z(n949) );
  NAND U691 ( .A(n955), .B(n956), .Z(n953) );
  XNOR U692 ( .A(n955), .B(n957), .Z(SUM[838]) );
  NANDN U693 ( .A(n954), .B(n956), .Z(n957) );
  NANDN U694 ( .A(n958), .B(n959), .Z(n955) );
  NAND U695 ( .A(n960), .B(n961), .Z(n959) );
  XNOR U696 ( .A(n960), .B(n962), .Z(SUM[837]) );
  NANDN U697 ( .A(n958), .B(n961), .Z(n962) );
  NANDN U698 ( .A(n963), .B(n964), .Z(n960) );
  NANDN U699 ( .A(n939), .B(n965), .Z(n964) );
  XOR U700 ( .A(n939), .B(n966), .Z(SUM[836]) );
  NANDN U701 ( .A(n963), .B(n965), .Z(n966) );
  ANDN U702 ( .B(n967), .A(n968), .Z(n939) );
  OR U703 ( .A(n969), .B(n970), .Z(n967) );
  XOR U704 ( .A(n971), .B(n972), .Z(SUM[835]) );
  NANDN U705 ( .A(n973), .B(n974), .Z(n972) );
  ANDN U706 ( .B(n975), .A(n976), .Z(n971) );
  NANDN U707 ( .A(n977), .B(n978), .Z(n975) );
  XNOR U708 ( .A(n978), .B(n979), .Z(SUM[834]) );
  OR U709 ( .A(n977), .B(n976), .Z(n979) );
  NANDN U710 ( .A(n980), .B(n981), .Z(n978) );
  NAND U711 ( .A(n982), .B(n983), .Z(n981) );
  XNOR U712 ( .A(n982), .B(n984), .Z(SUM[833]) );
  NANDN U713 ( .A(n980), .B(n983), .Z(n984) );
  NANDN U714 ( .A(n985), .B(n986), .Z(n982) );
  NANDN U715 ( .A(n970), .B(n987), .Z(n986) );
  XOR U716 ( .A(n970), .B(n988), .Z(SUM[832]) );
  NANDN U717 ( .A(n985), .B(n987), .Z(n988) );
  XOR U718 ( .A(n989), .B(n990), .Z(SUM[831]) );
  OR U719 ( .A(n991), .B(n992), .Z(n990) );
  ANDN U720 ( .B(n993), .A(n994), .Z(n989) );
  NANDN U721 ( .A(n995), .B(n996), .Z(n993) );
  XNOR U722 ( .A(n996), .B(n997), .Z(SUM[830]) );
  OR U723 ( .A(n995), .B(n994), .Z(n997) );
  NANDN U724 ( .A(n998), .B(n999), .Z(n996) );
  NANDN U725 ( .A(n1000), .B(n1001), .Z(n999) );
  XNOR U726 ( .A(n948), .B(n1002), .Z(SUM[82]) );
  OR U727 ( .A(n947), .B(n946), .Z(n1002) );
  NANDN U728 ( .A(n1003), .B(n1004), .Z(n948) );
  NAND U729 ( .A(n1005), .B(n1006), .Z(n1004) );
  XNOR U730 ( .A(n1001), .B(n1007), .Z(SUM[829]) );
  OR U731 ( .A(n1000), .B(n998), .Z(n1007) );
  NANDN U732 ( .A(n1008), .B(n1009), .Z(n1001) );
  NAND U733 ( .A(n1010), .B(n1011), .Z(n1009) );
  XNOR U734 ( .A(n1010), .B(n1012), .Z(SUM[828]) );
  NANDN U735 ( .A(n1008), .B(n1011), .Z(n1012) );
  NANDN U736 ( .A(n1013), .B(n1014), .Z(n1010) );
  NANDN U737 ( .A(n1015), .B(n1016), .Z(n1014) );
  XOR U738 ( .A(n1017), .B(n1018), .Z(SUM[827]) );
  NANDN U739 ( .A(n1019), .B(n1020), .Z(n1018) );
  ANDN U740 ( .B(n1021), .A(n1022), .Z(n1017) );
  NAND U741 ( .A(n1023), .B(n1024), .Z(n1021) );
  XNOR U742 ( .A(n1023), .B(n1025), .Z(SUM[826]) );
  NANDN U743 ( .A(n1022), .B(n1024), .Z(n1025) );
  NANDN U744 ( .A(n1026), .B(n1027), .Z(n1023) );
  NAND U745 ( .A(n1028), .B(n1029), .Z(n1027) );
  XNOR U746 ( .A(n1028), .B(n1030), .Z(SUM[825]) );
  NANDN U747 ( .A(n1026), .B(n1029), .Z(n1030) );
  NANDN U748 ( .A(n1031), .B(n1032), .Z(n1028) );
  NAND U749 ( .A(n1016), .B(n1033), .Z(n1032) );
  XNOR U750 ( .A(n1016), .B(n1034), .Z(SUM[824]) );
  NANDN U751 ( .A(n1031), .B(n1033), .Z(n1034) );
  NANDN U752 ( .A(n1035), .B(n1036), .Z(n1016) );
  NANDN U753 ( .A(n1037), .B(n1038), .Z(n1036) );
  XOR U754 ( .A(n1039), .B(n1040), .Z(SUM[823]) );
  NANDN U755 ( .A(n1041), .B(n1042), .Z(n1040) );
  ANDN U756 ( .B(n1043), .A(n1044), .Z(n1039) );
  NAND U757 ( .A(n1045), .B(n1046), .Z(n1043) );
  XNOR U758 ( .A(n1045), .B(n1047), .Z(SUM[822]) );
  NANDN U759 ( .A(n1044), .B(n1046), .Z(n1047) );
  NANDN U760 ( .A(n1048), .B(n1049), .Z(n1045) );
  NAND U761 ( .A(n1050), .B(n1051), .Z(n1049) );
  XNOR U762 ( .A(n1050), .B(n1052), .Z(SUM[821]) );
  NANDN U763 ( .A(n1048), .B(n1051), .Z(n1052) );
  NANDN U764 ( .A(n1053), .B(n1054), .Z(n1050) );
  NANDN U765 ( .A(n1037), .B(n1055), .Z(n1054) );
  XOR U766 ( .A(n1037), .B(n1056), .Z(SUM[820]) );
  NANDN U767 ( .A(n1053), .B(n1055), .Z(n1056) );
  ANDN U768 ( .B(n1057), .A(n1058), .Z(n1037) );
  OR U769 ( .A(n1059), .B(n1060), .Z(n1057) );
  XNOR U770 ( .A(n1005), .B(n1061), .Z(SUM[81]) );
  NANDN U771 ( .A(n1003), .B(n1006), .Z(n1061) );
  NANDN U772 ( .A(n1062), .B(n1063), .Z(n1005) );
  NANDN U773 ( .A(n890), .B(n1064), .Z(n1063) );
  XOR U774 ( .A(n1065), .B(n1066), .Z(SUM[819]) );
  NANDN U775 ( .A(n1067), .B(n1068), .Z(n1066) );
  ANDN U776 ( .B(n1069), .A(n1070), .Z(n1065) );
  NANDN U777 ( .A(n1071), .B(n1072), .Z(n1069) );
  XNOR U778 ( .A(n1072), .B(n1073), .Z(SUM[818]) );
  OR U779 ( .A(n1071), .B(n1070), .Z(n1073) );
  NANDN U780 ( .A(n1074), .B(n1075), .Z(n1072) );
  NAND U781 ( .A(n1076), .B(n1077), .Z(n1075) );
  XNOR U782 ( .A(n1076), .B(n1078), .Z(SUM[817]) );
  NANDN U783 ( .A(n1074), .B(n1077), .Z(n1078) );
  NANDN U784 ( .A(n1079), .B(n1080), .Z(n1076) );
  NANDN U785 ( .A(n1060), .B(n1081), .Z(n1080) );
  XOR U786 ( .A(n1060), .B(n1082), .Z(SUM[816]) );
  NANDN U787 ( .A(n1079), .B(n1081), .Z(n1082) );
  XOR U788 ( .A(n1083), .B(n1084), .Z(SUM[815]) );
  OR U789 ( .A(n1085), .B(n1086), .Z(n1084) );
  ANDN U790 ( .B(n1087), .A(n1088), .Z(n1083) );
  NANDN U791 ( .A(n1089), .B(n1090), .Z(n1087) );
  XNOR U792 ( .A(n1090), .B(n1091), .Z(SUM[814]) );
  OR U793 ( .A(n1089), .B(n1088), .Z(n1091) );
  NANDN U794 ( .A(n1092), .B(n1093), .Z(n1090) );
  NANDN U795 ( .A(n1094), .B(n1095), .Z(n1093) );
  XNOR U796 ( .A(n1095), .B(n1096), .Z(SUM[813]) );
  OR U797 ( .A(n1094), .B(n1092), .Z(n1096) );
  NANDN U798 ( .A(n1097), .B(n1098), .Z(n1095) );
  NAND U799 ( .A(n1099), .B(n1100), .Z(n1098) );
  XNOR U800 ( .A(n1099), .B(n1101), .Z(SUM[812]) );
  NANDN U801 ( .A(n1097), .B(n1100), .Z(n1101) );
  NANDN U802 ( .A(n1102), .B(n1103), .Z(n1099) );
  NANDN U803 ( .A(n1104), .B(n1105), .Z(n1103) );
  XOR U804 ( .A(n1106), .B(n1107), .Z(SUM[811]) );
  NANDN U805 ( .A(n1108), .B(n1109), .Z(n1107) );
  ANDN U806 ( .B(n1110), .A(n1111), .Z(n1106) );
  NAND U807 ( .A(n1112), .B(n1113), .Z(n1110) );
  XNOR U808 ( .A(n1112), .B(n1114), .Z(SUM[810]) );
  NANDN U809 ( .A(n1111), .B(n1113), .Z(n1114) );
  NANDN U810 ( .A(n1115), .B(n1116), .Z(n1112) );
  NAND U811 ( .A(n1117), .B(n1118), .Z(n1116) );
  XOR U812 ( .A(n890), .B(n1119), .Z(SUM[80]) );
  NANDN U813 ( .A(n1062), .B(n1064), .Z(n1119) );
  XNOR U814 ( .A(n1117), .B(n1120), .Z(SUM[809]) );
  NANDN U815 ( .A(n1115), .B(n1118), .Z(n1120) );
  NANDN U816 ( .A(n1121), .B(n1122), .Z(n1117) );
  NAND U817 ( .A(n1105), .B(n1123), .Z(n1122) );
  XNOR U818 ( .A(n1105), .B(n1124), .Z(SUM[808]) );
  NANDN U819 ( .A(n1121), .B(n1123), .Z(n1124) );
  NANDN U820 ( .A(n1125), .B(n1126), .Z(n1105) );
  NANDN U821 ( .A(n1127), .B(n1128), .Z(n1126) );
  XOR U822 ( .A(n1129), .B(n1130), .Z(SUM[807]) );
  NANDN U823 ( .A(n1131), .B(n1132), .Z(n1130) );
  ANDN U824 ( .B(n1133), .A(n1134), .Z(n1129) );
  NAND U825 ( .A(n1135), .B(n1136), .Z(n1133) );
  XNOR U826 ( .A(n1135), .B(n1137), .Z(SUM[806]) );
  NANDN U827 ( .A(n1134), .B(n1136), .Z(n1137) );
  NANDN U828 ( .A(n1138), .B(n1139), .Z(n1135) );
  NAND U829 ( .A(n1140), .B(n1141), .Z(n1139) );
  XNOR U830 ( .A(n1140), .B(n1142), .Z(SUM[805]) );
  NANDN U831 ( .A(n1138), .B(n1141), .Z(n1142) );
  NANDN U832 ( .A(n1143), .B(n1144), .Z(n1140) );
  NANDN U833 ( .A(n1127), .B(n1145), .Z(n1144) );
  XOR U834 ( .A(n1127), .B(n1146), .Z(SUM[804]) );
  NANDN U835 ( .A(n1143), .B(n1145), .Z(n1146) );
  ANDN U836 ( .B(n1147), .A(n1148), .Z(n1127) );
  OR U837 ( .A(n1149), .B(n1150), .Z(n1147) );
  XOR U838 ( .A(n1151), .B(n1152), .Z(SUM[803]) );
  NANDN U839 ( .A(n1153), .B(n1154), .Z(n1152) );
  ANDN U840 ( .B(n1155), .A(n1156), .Z(n1151) );
  NANDN U841 ( .A(n1157), .B(n1158), .Z(n1155) );
  XNOR U842 ( .A(n1158), .B(n1159), .Z(SUM[802]) );
  OR U843 ( .A(n1157), .B(n1156), .Z(n1159) );
  NANDN U844 ( .A(n1160), .B(n1161), .Z(n1158) );
  NAND U845 ( .A(n1162), .B(n1163), .Z(n1161) );
  XNOR U846 ( .A(n1162), .B(n1164), .Z(SUM[801]) );
  NANDN U847 ( .A(n1160), .B(n1163), .Z(n1164) );
  NANDN U848 ( .A(n1165), .B(n1166), .Z(n1162) );
  NANDN U849 ( .A(n1150), .B(n1167), .Z(n1166) );
  XOR U850 ( .A(n1150), .B(n1168), .Z(SUM[800]) );
  NANDN U851 ( .A(n1165), .B(n1167), .Z(n1168) );
  XOR U852 ( .A(n1169), .B(n1170), .Z(SUM[7]) );
  OR U853 ( .A(n1171), .B(n1172), .Z(n1170) );
  ANDN U854 ( .B(n1173), .A(n1174), .Z(n1169) );
  XOR U855 ( .A(n1175), .B(n1176), .Z(SUM[79]) );
  NANDN U856 ( .A(n1177), .B(n1178), .Z(n1176) );
  ANDN U857 ( .B(n1179), .A(n1180), .Z(n1175) );
  NANDN U858 ( .A(n1181), .B(n1182), .Z(n1179) );
  XOR U859 ( .A(n1183), .B(n1184), .Z(SUM[799]) );
  OR U860 ( .A(n1185), .B(n1186), .Z(n1184) );
  ANDN U861 ( .B(n1187), .A(n1188), .Z(n1183) );
  NANDN U862 ( .A(n1189), .B(n1190), .Z(n1187) );
  XNOR U863 ( .A(n1190), .B(n1191), .Z(SUM[798]) );
  OR U864 ( .A(n1189), .B(n1188), .Z(n1191) );
  NANDN U865 ( .A(n1192), .B(n1193), .Z(n1190) );
  NANDN U866 ( .A(n1194), .B(n1195), .Z(n1193) );
  XNOR U867 ( .A(n1195), .B(n1196), .Z(SUM[797]) );
  OR U868 ( .A(n1194), .B(n1192), .Z(n1196) );
  NANDN U869 ( .A(n1197), .B(n1198), .Z(n1195) );
  NAND U870 ( .A(n1199), .B(n1200), .Z(n1198) );
  XNOR U871 ( .A(n1199), .B(n1201), .Z(SUM[796]) );
  NANDN U872 ( .A(n1197), .B(n1200), .Z(n1201) );
  NANDN U873 ( .A(n1202), .B(n1203), .Z(n1199) );
  NANDN U874 ( .A(n1204), .B(n1205), .Z(n1203) );
  XOR U875 ( .A(n1206), .B(n1207), .Z(SUM[795]) );
  NANDN U876 ( .A(n1208), .B(n1209), .Z(n1207) );
  ANDN U877 ( .B(n1210), .A(n1211), .Z(n1206) );
  NAND U878 ( .A(n1212), .B(n1213), .Z(n1210) );
  XNOR U879 ( .A(n1212), .B(n1214), .Z(SUM[794]) );
  NANDN U880 ( .A(n1211), .B(n1213), .Z(n1214) );
  NANDN U881 ( .A(n1215), .B(n1216), .Z(n1212) );
  NAND U882 ( .A(n1217), .B(n1218), .Z(n1216) );
  XNOR U883 ( .A(n1217), .B(n1219), .Z(SUM[793]) );
  NANDN U884 ( .A(n1215), .B(n1218), .Z(n1219) );
  NANDN U885 ( .A(n1220), .B(n1221), .Z(n1217) );
  NAND U886 ( .A(n1205), .B(n1222), .Z(n1221) );
  XNOR U887 ( .A(n1205), .B(n1223), .Z(SUM[792]) );
  NANDN U888 ( .A(n1220), .B(n1222), .Z(n1223) );
  NANDN U889 ( .A(n1224), .B(n1225), .Z(n1205) );
  NANDN U890 ( .A(n1226), .B(n1227), .Z(n1225) );
  XOR U891 ( .A(n1228), .B(n1229), .Z(SUM[791]) );
  NANDN U892 ( .A(n1230), .B(n1231), .Z(n1229) );
  ANDN U893 ( .B(n1232), .A(n1233), .Z(n1228) );
  NAND U894 ( .A(n1234), .B(n1235), .Z(n1232) );
  XNOR U895 ( .A(n1234), .B(n1236), .Z(SUM[790]) );
  NANDN U896 ( .A(n1233), .B(n1235), .Z(n1236) );
  NANDN U897 ( .A(n1237), .B(n1238), .Z(n1234) );
  NAND U898 ( .A(n1239), .B(n1240), .Z(n1238) );
  XNOR U899 ( .A(n1182), .B(n1241), .Z(SUM[78]) );
  OR U900 ( .A(n1181), .B(n1180), .Z(n1241) );
  NANDN U901 ( .A(n1242), .B(n1243), .Z(n1182) );
  NAND U902 ( .A(n1244), .B(n1245), .Z(n1243) );
  XNOR U903 ( .A(n1239), .B(n1246), .Z(SUM[789]) );
  NANDN U904 ( .A(n1237), .B(n1240), .Z(n1246) );
  NANDN U905 ( .A(n1247), .B(n1248), .Z(n1239) );
  NANDN U906 ( .A(n1226), .B(n1249), .Z(n1248) );
  XOR U907 ( .A(n1226), .B(n1250), .Z(SUM[788]) );
  NANDN U908 ( .A(n1247), .B(n1249), .Z(n1250) );
  ANDN U909 ( .B(n1251), .A(n1252), .Z(n1226) );
  OR U910 ( .A(n1253), .B(n1254), .Z(n1251) );
  XOR U911 ( .A(n1255), .B(n1256), .Z(SUM[787]) );
  NANDN U912 ( .A(n1257), .B(n1258), .Z(n1256) );
  ANDN U913 ( .B(n1259), .A(n1260), .Z(n1255) );
  NANDN U914 ( .A(n1261), .B(n1262), .Z(n1259) );
  XNOR U915 ( .A(n1262), .B(n1263), .Z(SUM[786]) );
  OR U916 ( .A(n1261), .B(n1260), .Z(n1263) );
  NANDN U917 ( .A(n1264), .B(n1265), .Z(n1262) );
  NAND U918 ( .A(n1266), .B(n1267), .Z(n1265) );
  XNOR U919 ( .A(n1266), .B(n1268), .Z(SUM[785]) );
  NANDN U920 ( .A(n1264), .B(n1267), .Z(n1268) );
  NANDN U921 ( .A(n1269), .B(n1270), .Z(n1266) );
  NANDN U922 ( .A(n1254), .B(n1271), .Z(n1270) );
  XOR U923 ( .A(n1254), .B(n1272), .Z(SUM[784]) );
  NANDN U924 ( .A(n1269), .B(n1271), .Z(n1272) );
  XOR U925 ( .A(n1273), .B(n1274), .Z(SUM[783]) );
  OR U926 ( .A(n1275), .B(n1276), .Z(n1274) );
  ANDN U927 ( .B(n1277), .A(n1278), .Z(n1273) );
  NANDN U928 ( .A(n1279), .B(n1280), .Z(n1277) );
  XNOR U929 ( .A(n1280), .B(n1281), .Z(SUM[782]) );
  OR U930 ( .A(n1279), .B(n1278), .Z(n1281) );
  NANDN U931 ( .A(n1282), .B(n1283), .Z(n1280) );
  NANDN U932 ( .A(n1284), .B(n1285), .Z(n1283) );
  XNOR U933 ( .A(n1285), .B(n1286), .Z(SUM[781]) );
  OR U934 ( .A(n1284), .B(n1282), .Z(n1286) );
  NANDN U935 ( .A(n1287), .B(n1288), .Z(n1285) );
  NAND U936 ( .A(n1289), .B(n1290), .Z(n1288) );
  XNOR U937 ( .A(n1289), .B(n1291), .Z(SUM[780]) );
  NANDN U938 ( .A(n1287), .B(n1290), .Z(n1291) );
  NANDN U939 ( .A(n1292), .B(n1293), .Z(n1289) );
  NANDN U940 ( .A(n1294), .B(n1295), .Z(n1293) );
  XNOR U941 ( .A(n1244), .B(n1296), .Z(SUM[77]) );
  NANDN U942 ( .A(n1242), .B(n1245), .Z(n1296) );
  NANDN U943 ( .A(n1297), .B(n1298), .Z(n1244) );
  NANDN U944 ( .A(n1299), .B(n1300), .Z(n1298) );
  XOR U945 ( .A(n1301), .B(n1302), .Z(SUM[779]) );
  NANDN U946 ( .A(n1303), .B(n1304), .Z(n1302) );
  ANDN U947 ( .B(n1305), .A(n1306), .Z(n1301) );
  NAND U948 ( .A(n1307), .B(n1308), .Z(n1305) );
  XNOR U949 ( .A(n1307), .B(n1309), .Z(SUM[778]) );
  NANDN U950 ( .A(n1306), .B(n1308), .Z(n1309) );
  NANDN U951 ( .A(n1310), .B(n1311), .Z(n1307) );
  NAND U952 ( .A(n1312), .B(n1313), .Z(n1311) );
  XNOR U953 ( .A(n1312), .B(n1314), .Z(SUM[777]) );
  NANDN U954 ( .A(n1310), .B(n1313), .Z(n1314) );
  NANDN U955 ( .A(n1315), .B(n1316), .Z(n1312) );
  NAND U956 ( .A(n1295), .B(n1317), .Z(n1316) );
  XNOR U957 ( .A(n1295), .B(n1318), .Z(SUM[776]) );
  NANDN U958 ( .A(n1315), .B(n1317), .Z(n1318) );
  NANDN U959 ( .A(n1319), .B(n1320), .Z(n1295) );
  NANDN U960 ( .A(n1321), .B(n1322), .Z(n1320) );
  XOR U961 ( .A(n1323), .B(n1324), .Z(SUM[775]) );
  NANDN U962 ( .A(n1325), .B(n1326), .Z(n1324) );
  ANDN U963 ( .B(n1327), .A(n1328), .Z(n1323) );
  NAND U964 ( .A(n1329), .B(n1330), .Z(n1327) );
  XNOR U965 ( .A(n1329), .B(n1331), .Z(SUM[774]) );
  NANDN U966 ( .A(n1328), .B(n1330), .Z(n1331) );
  NANDN U967 ( .A(n1332), .B(n1333), .Z(n1329) );
  NAND U968 ( .A(n1334), .B(n1335), .Z(n1333) );
  XNOR U969 ( .A(n1334), .B(n1336), .Z(SUM[773]) );
  NANDN U970 ( .A(n1332), .B(n1335), .Z(n1336) );
  NANDN U971 ( .A(n1337), .B(n1338), .Z(n1334) );
  NANDN U972 ( .A(n1321), .B(n1339), .Z(n1338) );
  XOR U973 ( .A(n1321), .B(n1340), .Z(SUM[772]) );
  NANDN U974 ( .A(n1337), .B(n1339), .Z(n1340) );
  ANDN U975 ( .B(n1341), .A(n1342), .Z(n1321) );
  OR U976 ( .A(n1343), .B(n1344), .Z(n1341) );
  XOR U977 ( .A(n1345), .B(n1346), .Z(SUM[771]) );
  NANDN U978 ( .A(n1347), .B(n1348), .Z(n1346) );
  ANDN U979 ( .B(n1349), .A(n1350), .Z(n1345) );
  NANDN U980 ( .A(n1351), .B(n1352), .Z(n1349) );
  XNOR U981 ( .A(n1352), .B(n1353), .Z(SUM[770]) );
  OR U982 ( .A(n1351), .B(n1350), .Z(n1353) );
  NANDN U983 ( .A(n1354), .B(n1355), .Z(n1352) );
  NAND U984 ( .A(n1356), .B(n1357), .Z(n1355) );
  XNOR U985 ( .A(n1300), .B(n1358), .Z(SUM[76]) );
  OR U986 ( .A(n1299), .B(n1297), .Z(n1358) );
  NANDN U987 ( .A(n1359), .B(n1360), .Z(n1300) );
  NANDN U988 ( .A(n1361), .B(n1362), .Z(n1360) );
  XNOR U989 ( .A(n1356), .B(n1363), .Z(SUM[769]) );
  NANDN U990 ( .A(n1354), .B(n1357), .Z(n1363) );
  NANDN U991 ( .A(n1364), .B(n1365), .Z(n1356) );
  NANDN U992 ( .A(n1344), .B(n1366), .Z(n1365) );
  XOR U993 ( .A(n1344), .B(n1367), .Z(SUM[768]) );
  NANDN U994 ( .A(n1364), .B(n1366), .Z(n1367) );
  XOR U995 ( .A(n1368), .B(n1369), .Z(SUM[767]) );
  OR U996 ( .A(n1370), .B(n1371), .Z(n1369) );
  ANDN U997 ( .B(n1372), .A(n1373), .Z(n1368) );
  NAND U998 ( .A(n1374), .B(n1375), .Z(n1372) );
  XNOR U999 ( .A(n1374), .B(n1376), .Z(SUM[766]) );
  NANDN U1000 ( .A(n1373), .B(n1375), .Z(n1376) );
  NANDN U1001 ( .A(n1377), .B(n1378), .Z(n1374) );
  NAND U1002 ( .A(n1379), .B(n1380), .Z(n1378) );
  XNOR U1003 ( .A(n1379), .B(n1381), .Z(SUM[765]) );
  NANDN U1004 ( .A(n1377), .B(n1380), .Z(n1381) );
  NANDN U1005 ( .A(n1382), .B(n1383), .Z(n1379) );
  NANDN U1006 ( .A(n1384), .B(n1385), .Z(n1383) );
  XNOR U1007 ( .A(n1385), .B(n1386), .Z(SUM[764]) );
  OR U1008 ( .A(n1384), .B(n1382), .Z(n1386) );
  NANDN U1009 ( .A(n1387), .B(n1388), .Z(n1385) );
  NANDN U1010 ( .A(n1389), .B(n1390), .Z(n1388) );
  XOR U1011 ( .A(n1391), .B(n1392), .Z(SUM[763]) );
  NANDN U1012 ( .A(n1393), .B(n1394), .Z(n1392) );
  ANDN U1013 ( .B(n1395), .A(n1396), .Z(n1391) );
  NAND U1014 ( .A(n1397), .B(n1398), .Z(n1395) );
  XNOR U1015 ( .A(n1397), .B(n1399), .Z(SUM[762]) );
  NANDN U1016 ( .A(n1396), .B(n1398), .Z(n1399) );
  NANDN U1017 ( .A(n1400), .B(n1401), .Z(n1397) );
  NAND U1018 ( .A(n1402), .B(n1403), .Z(n1401) );
  XNOR U1019 ( .A(n1402), .B(n1404), .Z(SUM[761]) );
  NANDN U1020 ( .A(n1400), .B(n1403), .Z(n1404) );
  NANDN U1021 ( .A(n1405), .B(n1406), .Z(n1402) );
  NAND U1022 ( .A(n1390), .B(n1407), .Z(n1406) );
  XNOR U1023 ( .A(n1390), .B(n1408), .Z(SUM[760]) );
  NANDN U1024 ( .A(n1405), .B(n1407), .Z(n1408) );
  NANDN U1025 ( .A(n1409), .B(n1410), .Z(n1390) );
  NANDN U1026 ( .A(n1411), .B(n1412), .Z(n1410) );
  XOR U1027 ( .A(n1413), .B(n1414), .Z(SUM[75]) );
  NANDN U1028 ( .A(n1415), .B(n1416), .Z(n1414) );
  ANDN U1029 ( .B(n1417), .A(n1418), .Z(n1413) );
  NAND U1030 ( .A(n1419), .B(n1420), .Z(n1417) );
  XOR U1031 ( .A(n1421), .B(n1422), .Z(SUM[759]) );
  NANDN U1032 ( .A(n1423), .B(n1424), .Z(n1422) );
  ANDN U1033 ( .B(n1425), .A(n1426), .Z(n1421) );
  NAND U1034 ( .A(n1427), .B(n1428), .Z(n1425) );
  XNOR U1035 ( .A(n1427), .B(n1429), .Z(SUM[758]) );
  NANDN U1036 ( .A(n1426), .B(n1428), .Z(n1429) );
  NANDN U1037 ( .A(n1430), .B(n1431), .Z(n1427) );
  NAND U1038 ( .A(n1432), .B(n1433), .Z(n1431) );
  XNOR U1039 ( .A(n1432), .B(n1434), .Z(SUM[757]) );
  NANDN U1040 ( .A(n1430), .B(n1433), .Z(n1434) );
  NANDN U1041 ( .A(n1435), .B(n1436), .Z(n1432) );
  NANDN U1042 ( .A(n1411), .B(n1437), .Z(n1436) );
  XOR U1043 ( .A(n1411), .B(n1438), .Z(SUM[756]) );
  NANDN U1044 ( .A(n1435), .B(n1437), .Z(n1438) );
  ANDN U1045 ( .B(n1439), .A(n1440), .Z(n1411) );
  NANDN U1046 ( .A(n1441), .B(n1442), .Z(n1439) );
  XOR U1047 ( .A(n1443), .B(n1444), .Z(SUM[755]) );
  NANDN U1048 ( .A(n1445), .B(n1446), .Z(n1444) );
  ANDN U1049 ( .B(n1447), .A(n1448), .Z(n1443) );
  NANDN U1050 ( .A(n1449), .B(n1450), .Z(n1447) );
  XNOR U1051 ( .A(n1450), .B(n1451), .Z(SUM[754]) );
  OR U1052 ( .A(n1449), .B(n1448), .Z(n1451) );
  NANDN U1053 ( .A(n1452), .B(n1453), .Z(n1450) );
  NAND U1054 ( .A(n1454), .B(n1455), .Z(n1453) );
  XNOR U1055 ( .A(n1454), .B(n1456), .Z(SUM[753]) );
  NANDN U1056 ( .A(n1452), .B(n1455), .Z(n1456) );
  NANDN U1057 ( .A(n1457), .B(n1458), .Z(n1454) );
  NAND U1058 ( .A(n1442), .B(n1459), .Z(n1458) );
  XNOR U1059 ( .A(n1442), .B(n1460), .Z(SUM[752]) );
  NANDN U1060 ( .A(n1457), .B(n1459), .Z(n1460) );
  NANDN U1061 ( .A(n1461), .B(n1462), .Z(n1442) );
  NANDN U1062 ( .A(n1463), .B(n1464), .Z(n1462) );
  XOR U1063 ( .A(n1465), .B(n1466), .Z(SUM[751]) );
  NANDN U1064 ( .A(n1467), .B(n1468), .Z(n1466) );
  ANDN U1065 ( .B(n1469), .A(n1470), .Z(n1465) );
  NAND U1066 ( .A(n1471), .B(n1472), .Z(n1469) );
  XNOR U1067 ( .A(n1471), .B(n1473), .Z(SUM[750]) );
  NANDN U1068 ( .A(n1470), .B(n1472), .Z(n1473) );
  NANDN U1069 ( .A(n1474), .B(n1475), .Z(n1471) );
  NAND U1070 ( .A(n1476), .B(n1477), .Z(n1475) );
  XNOR U1071 ( .A(n1419), .B(n1478), .Z(SUM[74]) );
  NANDN U1072 ( .A(n1418), .B(n1420), .Z(n1478) );
  NANDN U1073 ( .A(n1479), .B(n1480), .Z(n1419) );
  NAND U1074 ( .A(n1481), .B(n1482), .Z(n1480) );
  XNOR U1075 ( .A(n1476), .B(n1483), .Z(SUM[749]) );
  NANDN U1076 ( .A(n1474), .B(n1477), .Z(n1483) );
  NANDN U1077 ( .A(n1484), .B(n1485), .Z(n1476) );
  NAND U1078 ( .A(n1486), .B(n1487), .Z(n1485) );
  XNOR U1079 ( .A(n1486), .B(n1488), .Z(SUM[748]) );
  NANDN U1080 ( .A(n1484), .B(n1487), .Z(n1488) );
  NANDN U1081 ( .A(n1489), .B(n1490), .Z(n1486) );
  NAND U1082 ( .A(n1491), .B(n1492), .Z(n1490) );
  XOR U1083 ( .A(n1493), .B(n1494), .Z(SUM[747]) );
  NANDN U1084 ( .A(n1495), .B(n1496), .Z(n1494) );
  ANDN U1085 ( .B(n1497), .A(n1498), .Z(n1493) );
  NAND U1086 ( .A(n1499), .B(n1500), .Z(n1497) );
  XNOR U1087 ( .A(n1499), .B(n1501), .Z(SUM[746]) );
  NANDN U1088 ( .A(n1498), .B(n1500), .Z(n1501) );
  NANDN U1089 ( .A(n1502), .B(n1503), .Z(n1499) );
  NAND U1090 ( .A(n1504), .B(n1505), .Z(n1503) );
  XNOR U1091 ( .A(n1504), .B(n1506), .Z(SUM[745]) );
  NANDN U1092 ( .A(n1502), .B(n1505), .Z(n1506) );
  NANDN U1093 ( .A(n1507), .B(n1508), .Z(n1504) );
  NAND U1094 ( .A(n1492), .B(n1509), .Z(n1508) );
  XNOR U1095 ( .A(n1492), .B(n1510), .Z(SUM[744]) );
  NANDN U1096 ( .A(n1507), .B(n1509), .Z(n1510) );
  NANDN U1097 ( .A(n1511), .B(n1512), .Z(n1492) );
  OR U1098 ( .A(n1513), .B(n1514), .Z(n1512) );
  XOR U1099 ( .A(n1515), .B(n1516), .Z(SUM[743]) );
  NANDN U1100 ( .A(n1517), .B(n1518), .Z(n1516) );
  ANDN U1101 ( .B(n1519), .A(n1520), .Z(n1515) );
  NAND U1102 ( .A(n1521), .B(n1522), .Z(n1519) );
  XNOR U1103 ( .A(n1521), .B(n1523), .Z(SUM[742]) );
  NANDN U1104 ( .A(n1520), .B(n1522), .Z(n1523) );
  NANDN U1105 ( .A(n1524), .B(n1525), .Z(n1521) );
  NAND U1106 ( .A(n1526), .B(n1527), .Z(n1525) );
  XNOR U1107 ( .A(n1526), .B(n1528), .Z(SUM[741]) );
  NANDN U1108 ( .A(n1524), .B(n1527), .Z(n1528) );
  NANDN U1109 ( .A(n1529), .B(n1530), .Z(n1526) );
  NANDN U1110 ( .A(n1514), .B(n1531), .Z(n1530) );
  XOR U1111 ( .A(n1514), .B(n1532), .Z(SUM[740]) );
  NANDN U1112 ( .A(n1529), .B(n1531), .Z(n1532) );
  ANDN U1113 ( .B(n1533), .A(n1534), .Z(n1514) );
  NANDN U1114 ( .A(n1535), .B(n1464), .Z(n1533) );
  XNOR U1115 ( .A(n1481), .B(n1536), .Z(SUM[73]) );
  NANDN U1116 ( .A(n1479), .B(n1482), .Z(n1536) );
  NANDN U1117 ( .A(n1537), .B(n1538), .Z(n1481) );
  NAND U1118 ( .A(n1362), .B(n1539), .Z(n1538) );
  XOR U1119 ( .A(n1540), .B(n1541), .Z(SUM[739]) );
  NANDN U1120 ( .A(n1542), .B(n1543), .Z(n1541) );
  ANDN U1121 ( .B(n1544), .A(n1545), .Z(n1540) );
  NAND U1122 ( .A(n1546), .B(n1547), .Z(n1544) );
  XNOR U1123 ( .A(n1546), .B(n1548), .Z(SUM[738]) );
  NANDN U1124 ( .A(n1545), .B(n1547), .Z(n1548) );
  NANDN U1125 ( .A(n1549), .B(n1550), .Z(n1546) );
  NAND U1126 ( .A(n1551), .B(n1552), .Z(n1550) );
  XNOR U1127 ( .A(n1551), .B(n1553), .Z(SUM[737]) );
  NANDN U1128 ( .A(n1549), .B(n1552), .Z(n1553) );
  NANDN U1129 ( .A(n1554), .B(n1555), .Z(n1551) );
  NAND U1130 ( .A(n1464), .B(n1556), .Z(n1555) );
  XNOR U1131 ( .A(n1464), .B(n1557), .Z(SUM[736]) );
  NANDN U1132 ( .A(n1554), .B(n1556), .Z(n1557) );
  NANDN U1133 ( .A(n1558), .B(n1559), .Z(n1464) );
  NANDN U1134 ( .A(n1560), .B(n1561), .Z(n1559) );
  XOR U1135 ( .A(n1562), .B(n1563), .Z(SUM[735]) );
  NANDN U1136 ( .A(n1564), .B(n1565), .Z(n1563) );
  ANDN U1137 ( .B(n1566), .A(n1567), .Z(n1562) );
  NAND U1138 ( .A(n1568), .B(n1569), .Z(n1566) );
  XNOR U1139 ( .A(n1568), .B(n1570), .Z(SUM[734]) );
  NANDN U1140 ( .A(n1567), .B(n1569), .Z(n1570) );
  NANDN U1141 ( .A(n1571), .B(n1572), .Z(n1568) );
  NAND U1142 ( .A(n1573), .B(n1574), .Z(n1572) );
  XNOR U1143 ( .A(n1573), .B(n1575), .Z(SUM[733]) );
  NANDN U1144 ( .A(n1571), .B(n1574), .Z(n1575) );
  NANDN U1145 ( .A(n1576), .B(n1577), .Z(n1573) );
  NAND U1146 ( .A(n1578), .B(n1579), .Z(n1577) );
  XNOR U1147 ( .A(n1578), .B(n1580), .Z(SUM[732]) );
  NANDN U1148 ( .A(n1576), .B(n1579), .Z(n1580) );
  NANDN U1149 ( .A(n1581), .B(n1582), .Z(n1578) );
  NAND U1150 ( .A(n1583), .B(n1584), .Z(n1582) );
  XOR U1151 ( .A(n1585), .B(n1586), .Z(SUM[731]) );
  NANDN U1152 ( .A(n1587), .B(n1588), .Z(n1586) );
  ANDN U1153 ( .B(n1589), .A(n1590), .Z(n1585) );
  NAND U1154 ( .A(n1591), .B(n1592), .Z(n1589) );
  XNOR U1155 ( .A(n1591), .B(n1593), .Z(SUM[730]) );
  NANDN U1156 ( .A(n1590), .B(n1592), .Z(n1593) );
  NANDN U1157 ( .A(n1594), .B(n1595), .Z(n1591) );
  NAND U1158 ( .A(n1596), .B(n1597), .Z(n1595) );
  XNOR U1159 ( .A(n1362), .B(n1598), .Z(SUM[72]) );
  NANDN U1160 ( .A(n1537), .B(n1539), .Z(n1598) );
  NANDN U1161 ( .A(n1599), .B(n1600), .Z(n1362) );
  NANDN U1162 ( .A(n1601), .B(n1602), .Z(n1600) );
  XNOR U1163 ( .A(n1596), .B(n1603), .Z(SUM[729]) );
  NANDN U1164 ( .A(n1594), .B(n1597), .Z(n1603) );
  NANDN U1165 ( .A(n1604), .B(n1605), .Z(n1596) );
  NAND U1166 ( .A(n1584), .B(n1606), .Z(n1605) );
  XNOR U1167 ( .A(n1584), .B(n1607), .Z(SUM[728]) );
  NANDN U1168 ( .A(n1604), .B(n1606), .Z(n1607) );
  NANDN U1169 ( .A(n1608), .B(n1609), .Z(n1584) );
  OR U1170 ( .A(n1610), .B(n1611), .Z(n1609) );
  XOR U1171 ( .A(n1612), .B(n1613), .Z(SUM[727]) );
  NANDN U1172 ( .A(n1614), .B(n1615), .Z(n1613) );
  ANDN U1173 ( .B(n1616), .A(n1617), .Z(n1612) );
  NAND U1174 ( .A(n1618), .B(n1619), .Z(n1616) );
  XNOR U1175 ( .A(n1618), .B(n1620), .Z(SUM[726]) );
  NANDN U1176 ( .A(n1617), .B(n1619), .Z(n1620) );
  NANDN U1177 ( .A(n1621), .B(n1622), .Z(n1618) );
  NAND U1178 ( .A(n1623), .B(n1624), .Z(n1622) );
  XNOR U1179 ( .A(n1623), .B(n1625), .Z(SUM[725]) );
  NANDN U1180 ( .A(n1621), .B(n1624), .Z(n1625) );
  NANDN U1181 ( .A(n1626), .B(n1627), .Z(n1623) );
  NANDN U1182 ( .A(n1611), .B(n1628), .Z(n1627) );
  XOR U1183 ( .A(n1611), .B(n1629), .Z(SUM[724]) );
  NANDN U1184 ( .A(n1626), .B(n1628), .Z(n1629) );
  ANDN U1185 ( .B(n1630), .A(n1631), .Z(n1611) );
  NANDN U1186 ( .A(n1632), .B(n1561), .Z(n1630) );
  XOR U1187 ( .A(n1633), .B(n1634), .Z(SUM[723]) );
  NANDN U1188 ( .A(n1635), .B(n1636), .Z(n1634) );
  ANDN U1189 ( .B(n1637), .A(n1638), .Z(n1633) );
  NAND U1190 ( .A(n1639), .B(n1640), .Z(n1637) );
  XNOR U1191 ( .A(n1639), .B(n1641), .Z(SUM[722]) );
  NANDN U1192 ( .A(n1638), .B(n1640), .Z(n1641) );
  NANDN U1193 ( .A(n1642), .B(n1643), .Z(n1639) );
  NAND U1194 ( .A(n1644), .B(n1645), .Z(n1643) );
  XNOR U1195 ( .A(n1644), .B(n1646), .Z(SUM[721]) );
  NANDN U1196 ( .A(n1642), .B(n1645), .Z(n1646) );
  NANDN U1197 ( .A(n1647), .B(n1648), .Z(n1644) );
  NAND U1198 ( .A(n1561), .B(n1649), .Z(n1648) );
  XNOR U1199 ( .A(n1561), .B(n1650), .Z(SUM[720]) );
  NANDN U1200 ( .A(n1647), .B(n1649), .Z(n1650) );
  NANDN U1201 ( .A(n1651), .B(n1652), .Z(n1561) );
  NANDN U1202 ( .A(n1653), .B(n1654), .Z(n1652) );
  XOR U1203 ( .A(n1655), .B(n1656), .Z(SUM[71]) );
  NANDN U1204 ( .A(n1657), .B(n1658), .Z(n1656) );
  ANDN U1205 ( .B(n1659), .A(n1660), .Z(n1655) );
  NAND U1206 ( .A(n1661), .B(n1662), .Z(n1659) );
  XOR U1207 ( .A(n1663), .B(n1664), .Z(SUM[719]) );
  NANDN U1208 ( .A(n1665), .B(n1666), .Z(n1664) );
  ANDN U1209 ( .B(n1667), .A(n1668), .Z(n1663) );
  NAND U1210 ( .A(n1669), .B(n1670), .Z(n1667) );
  XNOR U1211 ( .A(n1669), .B(n1671), .Z(SUM[718]) );
  NANDN U1212 ( .A(n1668), .B(n1670), .Z(n1671) );
  NANDN U1213 ( .A(n1672), .B(n1673), .Z(n1669) );
  NAND U1214 ( .A(n1674), .B(n1675), .Z(n1673) );
  XNOR U1215 ( .A(n1674), .B(n1676), .Z(SUM[717]) );
  NANDN U1216 ( .A(n1672), .B(n1675), .Z(n1676) );
  NANDN U1217 ( .A(n1677), .B(n1678), .Z(n1674) );
  NAND U1218 ( .A(n1679), .B(n1680), .Z(n1678) );
  XNOR U1219 ( .A(n1679), .B(n1681), .Z(SUM[716]) );
  NANDN U1220 ( .A(n1677), .B(n1680), .Z(n1681) );
  NANDN U1221 ( .A(n1682), .B(n1683), .Z(n1679) );
  NAND U1222 ( .A(n1684), .B(n1685), .Z(n1683) );
  XOR U1223 ( .A(n1686), .B(n1687), .Z(SUM[715]) );
  NANDN U1224 ( .A(n1688), .B(n1689), .Z(n1687) );
  ANDN U1225 ( .B(n1690), .A(n1691), .Z(n1686) );
  NAND U1226 ( .A(n1692), .B(n1693), .Z(n1690) );
  XNOR U1227 ( .A(n1692), .B(n1694), .Z(SUM[714]) );
  NANDN U1228 ( .A(n1691), .B(n1693), .Z(n1694) );
  NANDN U1229 ( .A(n1695), .B(n1696), .Z(n1692) );
  NAND U1230 ( .A(n1697), .B(n1698), .Z(n1696) );
  XNOR U1231 ( .A(n1697), .B(n1699), .Z(SUM[713]) );
  NANDN U1232 ( .A(n1695), .B(n1698), .Z(n1699) );
  NANDN U1233 ( .A(n1700), .B(n1701), .Z(n1697) );
  NAND U1234 ( .A(n1685), .B(n1702), .Z(n1701) );
  XNOR U1235 ( .A(n1685), .B(n1703), .Z(SUM[712]) );
  NANDN U1236 ( .A(n1700), .B(n1702), .Z(n1703) );
  NANDN U1237 ( .A(n1704), .B(n1705), .Z(n1685) );
  OR U1238 ( .A(n1706), .B(n1707), .Z(n1705) );
  XOR U1239 ( .A(n1708), .B(n1709), .Z(SUM[711]) );
  NANDN U1240 ( .A(n1710), .B(n1711), .Z(n1709) );
  ANDN U1241 ( .B(n1712), .A(n1713), .Z(n1708) );
  NAND U1242 ( .A(n1714), .B(n1715), .Z(n1712) );
  XNOR U1243 ( .A(n1714), .B(n1716), .Z(SUM[710]) );
  NANDN U1244 ( .A(n1713), .B(n1715), .Z(n1716) );
  NANDN U1245 ( .A(n1717), .B(n1718), .Z(n1714) );
  NAND U1246 ( .A(n1719), .B(n1720), .Z(n1718) );
  XNOR U1247 ( .A(n1661), .B(n1721), .Z(SUM[70]) );
  NANDN U1248 ( .A(n1660), .B(n1662), .Z(n1721) );
  NANDN U1249 ( .A(n1722), .B(n1723), .Z(n1661) );
  NAND U1250 ( .A(n1724), .B(n1725), .Z(n1723) );
  XNOR U1251 ( .A(n1719), .B(n1726), .Z(SUM[709]) );
  NANDN U1252 ( .A(n1717), .B(n1720), .Z(n1726) );
  NANDN U1253 ( .A(n1727), .B(n1728), .Z(n1719) );
  NANDN U1254 ( .A(n1707), .B(n1729), .Z(n1728) );
  XOR U1255 ( .A(n1707), .B(n1730), .Z(SUM[708]) );
  NANDN U1256 ( .A(n1727), .B(n1729), .Z(n1730) );
  ANDN U1257 ( .B(n1731), .A(n1732), .Z(n1707) );
  NANDN U1258 ( .A(n1733), .B(n1654), .Z(n1731) );
  XOR U1259 ( .A(n1734), .B(n1735), .Z(SUM[707]) );
  NANDN U1260 ( .A(n1736), .B(n1737), .Z(n1735) );
  ANDN U1261 ( .B(n1738), .A(n1739), .Z(n1734) );
  NAND U1262 ( .A(n1740), .B(n1741), .Z(n1738) );
  XNOR U1263 ( .A(n1740), .B(n1742), .Z(SUM[706]) );
  NANDN U1264 ( .A(n1739), .B(n1741), .Z(n1742) );
  NANDN U1265 ( .A(n1743), .B(n1744), .Z(n1740) );
  NAND U1266 ( .A(n1745), .B(n1746), .Z(n1744) );
  XNOR U1267 ( .A(n1745), .B(n1747), .Z(SUM[705]) );
  NANDN U1268 ( .A(n1743), .B(n1746), .Z(n1747) );
  NANDN U1269 ( .A(n1748), .B(n1749), .Z(n1745) );
  NAND U1270 ( .A(n1654), .B(n1750), .Z(n1749) );
  XNOR U1271 ( .A(n1654), .B(n1751), .Z(SUM[704]) );
  NANDN U1272 ( .A(n1748), .B(n1750), .Z(n1751) );
  NANDN U1273 ( .A(n1752), .B(n1753), .Z(n1654) );
  NANDN U1274 ( .A(n1754), .B(n1755), .Z(n1753) );
  XOR U1275 ( .A(n1756), .B(n1757), .Z(SUM[703]) );
  NANDN U1276 ( .A(n1758), .B(n1759), .Z(n1757) );
  ANDN U1277 ( .B(n1760), .A(n1761), .Z(n1756) );
  NAND U1278 ( .A(n1762), .B(n1763), .Z(n1760) );
  XNOR U1279 ( .A(n1762), .B(n1764), .Z(SUM[702]) );
  NANDN U1280 ( .A(n1761), .B(n1763), .Z(n1764) );
  NANDN U1281 ( .A(n1765), .B(n1766), .Z(n1762) );
  NAND U1282 ( .A(n1767), .B(n1768), .Z(n1766) );
  XNOR U1283 ( .A(n1767), .B(n1769), .Z(SUM[701]) );
  NANDN U1284 ( .A(n1765), .B(n1768), .Z(n1769) );
  NANDN U1285 ( .A(n1770), .B(n1771), .Z(n1767) );
  NAND U1286 ( .A(n1772), .B(n1773), .Z(n1771) );
  XNOR U1287 ( .A(n1772), .B(n1774), .Z(SUM[700]) );
  NANDN U1288 ( .A(n1770), .B(n1773), .Z(n1774) );
  NANDN U1289 ( .A(n1775), .B(n1776), .Z(n1772) );
  NANDN U1290 ( .A(n1777), .B(n1778), .Z(n1776) );
  XNOR U1291 ( .A(n1779), .B(n1780), .Z(SUM[6]) );
  OR U1292 ( .A(n1781), .B(n1174), .Z(n1780) );
  XNOR U1293 ( .A(n1724), .B(n1782), .Z(SUM[69]) );
  NANDN U1294 ( .A(n1722), .B(n1725), .Z(n1782) );
  NANDN U1295 ( .A(n1783), .B(n1784), .Z(n1724) );
  NANDN U1296 ( .A(n1601), .B(n1785), .Z(n1784) );
  XOR U1297 ( .A(n1786), .B(n1787), .Z(SUM[699]) );
  NANDN U1298 ( .A(n1788), .B(n1789), .Z(n1787) );
  ANDN U1299 ( .B(n1790), .A(n1791), .Z(n1786) );
  NAND U1300 ( .A(n1792), .B(n1793), .Z(n1790) );
  XNOR U1301 ( .A(n1792), .B(n1794), .Z(SUM[698]) );
  NANDN U1302 ( .A(n1791), .B(n1793), .Z(n1794) );
  NANDN U1303 ( .A(n1795), .B(n1796), .Z(n1792) );
  NAND U1304 ( .A(n1797), .B(n1798), .Z(n1796) );
  XNOR U1305 ( .A(n1797), .B(n1799), .Z(SUM[697]) );
  NANDN U1306 ( .A(n1795), .B(n1798), .Z(n1799) );
  NANDN U1307 ( .A(n1800), .B(n1801), .Z(n1797) );
  NAND U1308 ( .A(n1778), .B(n1802), .Z(n1801) );
  XNOR U1309 ( .A(n1778), .B(n1803), .Z(SUM[696]) );
  NANDN U1310 ( .A(n1800), .B(n1802), .Z(n1803) );
  NANDN U1311 ( .A(n1804), .B(n1805), .Z(n1778) );
  OR U1312 ( .A(n1806), .B(n1807), .Z(n1805) );
  XOR U1313 ( .A(n1808), .B(n1809), .Z(SUM[695]) );
  NANDN U1314 ( .A(n1810), .B(n1811), .Z(n1809) );
  ANDN U1315 ( .B(n1812), .A(n1813), .Z(n1808) );
  NAND U1316 ( .A(n1814), .B(n1815), .Z(n1812) );
  XNOR U1317 ( .A(n1814), .B(n1816), .Z(SUM[694]) );
  NANDN U1318 ( .A(n1813), .B(n1815), .Z(n1816) );
  NANDN U1319 ( .A(n1817), .B(n1818), .Z(n1814) );
  NAND U1320 ( .A(n1819), .B(n1820), .Z(n1818) );
  XNOR U1321 ( .A(n1819), .B(n1821), .Z(SUM[693]) );
  NANDN U1322 ( .A(n1817), .B(n1820), .Z(n1821) );
  NANDN U1323 ( .A(n1822), .B(n1823), .Z(n1819) );
  NANDN U1324 ( .A(n1807), .B(n1824), .Z(n1823) );
  XOR U1325 ( .A(n1807), .B(n1825), .Z(SUM[692]) );
  NANDN U1326 ( .A(n1822), .B(n1824), .Z(n1825) );
  ANDN U1327 ( .B(n1826), .A(n1827), .Z(n1807) );
  NANDN U1328 ( .A(n1828), .B(n1829), .Z(n1826) );
  XOR U1329 ( .A(n1830), .B(n1831), .Z(SUM[691]) );
  NANDN U1330 ( .A(n1832), .B(n1833), .Z(n1831) );
  ANDN U1331 ( .B(n1834), .A(n1835), .Z(n1830) );
  NAND U1332 ( .A(n1836), .B(n1837), .Z(n1834) );
  XNOR U1333 ( .A(n1836), .B(n1838), .Z(SUM[690]) );
  NANDN U1334 ( .A(n1835), .B(n1837), .Z(n1838) );
  NANDN U1335 ( .A(n1839), .B(n1840), .Z(n1836) );
  NAND U1336 ( .A(n1841), .B(n1842), .Z(n1840) );
  XOR U1337 ( .A(n1601), .B(n1843), .Z(SUM[68]) );
  NANDN U1338 ( .A(n1783), .B(n1785), .Z(n1843) );
  ANDN U1339 ( .B(n1844), .A(n1845), .Z(n1601) );
  OR U1340 ( .A(n1846), .B(n1847), .Z(n1844) );
  XNOR U1341 ( .A(n1841), .B(n1848), .Z(SUM[689]) );
  NANDN U1342 ( .A(n1839), .B(n1842), .Z(n1848) );
  NANDN U1343 ( .A(n1849), .B(n1850), .Z(n1841) );
  NAND U1344 ( .A(n1829), .B(n1851), .Z(n1850) );
  XNOR U1345 ( .A(n1829), .B(n1852), .Z(SUM[688]) );
  NANDN U1346 ( .A(n1849), .B(n1851), .Z(n1852) );
  NANDN U1347 ( .A(n1853), .B(n1854), .Z(n1829) );
  NAND U1348 ( .A(n1855), .B(n1856), .Z(n1854) );
  XOR U1349 ( .A(n1857), .B(n1858), .Z(SUM[687]) );
  NANDN U1350 ( .A(n1859), .B(n1860), .Z(n1858) );
  ANDN U1351 ( .B(n1861), .A(n1862), .Z(n1857) );
  NAND U1352 ( .A(n1863), .B(n1864), .Z(n1861) );
  XNOR U1353 ( .A(n1863), .B(n1865), .Z(SUM[686]) );
  NANDN U1354 ( .A(n1862), .B(n1864), .Z(n1865) );
  NANDN U1355 ( .A(n1866), .B(n1867), .Z(n1863) );
  NAND U1356 ( .A(n1868), .B(n1869), .Z(n1867) );
  XNOR U1357 ( .A(n1868), .B(n1870), .Z(SUM[685]) );
  NANDN U1358 ( .A(n1866), .B(n1869), .Z(n1870) );
  NANDN U1359 ( .A(n1871), .B(n1872), .Z(n1868) );
  NAND U1360 ( .A(n1873), .B(n1874), .Z(n1872) );
  XNOR U1361 ( .A(n1873), .B(n1875), .Z(SUM[684]) );
  NANDN U1362 ( .A(n1871), .B(n1874), .Z(n1875) );
  NANDN U1363 ( .A(n1876), .B(n1877), .Z(n1873) );
  NAND U1364 ( .A(n1878), .B(n1879), .Z(n1877) );
  XOR U1365 ( .A(n1880), .B(n1881), .Z(SUM[683]) );
  NANDN U1366 ( .A(n1882), .B(n1883), .Z(n1881) );
  ANDN U1367 ( .B(n1884), .A(n1885), .Z(n1880) );
  NAND U1368 ( .A(n1886), .B(n1887), .Z(n1884) );
  XNOR U1369 ( .A(n1886), .B(n1888), .Z(SUM[682]) );
  NANDN U1370 ( .A(n1885), .B(n1887), .Z(n1888) );
  NANDN U1371 ( .A(n1889), .B(n1890), .Z(n1886) );
  NAND U1372 ( .A(n1891), .B(n1892), .Z(n1890) );
  XNOR U1373 ( .A(n1891), .B(n1893), .Z(SUM[681]) );
  NANDN U1374 ( .A(n1889), .B(n1892), .Z(n1893) );
  NANDN U1375 ( .A(n1894), .B(n1895), .Z(n1891) );
  NAND U1376 ( .A(n1879), .B(n1896), .Z(n1895) );
  XNOR U1377 ( .A(n1879), .B(n1897), .Z(SUM[680]) );
  NANDN U1378 ( .A(n1894), .B(n1896), .Z(n1897) );
  NANDN U1379 ( .A(n1898), .B(n1899), .Z(n1879) );
  OR U1380 ( .A(n1900), .B(n1901), .Z(n1899) );
  XOR U1381 ( .A(n1902), .B(n1903), .Z(SUM[67]) );
  NANDN U1382 ( .A(n1904), .B(n1905), .Z(n1903) );
  ANDN U1383 ( .B(n1906), .A(n1907), .Z(n1902) );
  NANDN U1384 ( .A(n1908), .B(n1909), .Z(n1906) );
  XOR U1385 ( .A(n1910), .B(n1911), .Z(SUM[679]) );
  NANDN U1386 ( .A(n1912), .B(n1913), .Z(n1911) );
  ANDN U1387 ( .B(n1914), .A(n1915), .Z(n1910) );
  NAND U1388 ( .A(n1916), .B(n1917), .Z(n1914) );
  XNOR U1389 ( .A(n1916), .B(n1918), .Z(SUM[678]) );
  NANDN U1390 ( .A(n1915), .B(n1917), .Z(n1918) );
  NANDN U1391 ( .A(n1919), .B(n1920), .Z(n1916) );
  NAND U1392 ( .A(n1921), .B(n1922), .Z(n1920) );
  XNOR U1393 ( .A(n1921), .B(n1923), .Z(SUM[677]) );
  NANDN U1394 ( .A(n1919), .B(n1922), .Z(n1923) );
  NANDN U1395 ( .A(n1924), .B(n1925), .Z(n1921) );
  NANDN U1396 ( .A(n1901), .B(n1926), .Z(n1925) );
  XOR U1397 ( .A(n1901), .B(n1927), .Z(SUM[676]) );
  NANDN U1398 ( .A(n1924), .B(n1926), .Z(n1927) );
  ANDN U1399 ( .B(n1928), .A(n1929), .Z(n1901) );
  NANDN U1400 ( .A(n1930), .B(n1856), .Z(n1928) );
  XOR U1401 ( .A(n1931), .B(n1932), .Z(SUM[675]) );
  NANDN U1402 ( .A(n1933), .B(n1934), .Z(n1932) );
  ANDN U1403 ( .B(n1935), .A(n1936), .Z(n1931) );
  NAND U1404 ( .A(n1937), .B(n1938), .Z(n1935) );
  XNOR U1405 ( .A(n1937), .B(n1939), .Z(SUM[674]) );
  NANDN U1406 ( .A(n1936), .B(n1938), .Z(n1939) );
  NANDN U1407 ( .A(n1940), .B(n1941), .Z(n1937) );
  NAND U1408 ( .A(n1942), .B(n1943), .Z(n1941) );
  XNOR U1409 ( .A(n1942), .B(n1944), .Z(SUM[673]) );
  NANDN U1410 ( .A(n1940), .B(n1943), .Z(n1944) );
  NANDN U1411 ( .A(n1945), .B(n1946), .Z(n1942) );
  NAND U1412 ( .A(n1856), .B(n1947), .Z(n1946) );
  XNOR U1413 ( .A(n1856), .B(n1948), .Z(SUM[672]) );
  NANDN U1414 ( .A(n1945), .B(n1947), .Z(n1948) );
  NANDN U1415 ( .A(n1949), .B(n1950), .Z(n1856) );
  OR U1416 ( .A(n1951), .B(n1952), .Z(n1950) );
  XOR U1417 ( .A(n1953), .B(n1954), .Z(SUM[671]) );
  NANDN U1418 ( .A(n1955), .B(n1956), .Z(n1954) );
  ANDN U1419 ( .B(n1957), .A(n1958), .Z(n1953) );
  NAND U1420 ( .A(n1959), .B(n1960), .Z(n1957) );
  XNOR U1421 ( .A(n1959), .B(n1961), .Z(SUM[670]) );
  NANDN U1422 ( .A(n1958), .B(n1960), .Z(n1961) );
  NANDN U1423 ( .A(n1962), .B(n1963), .Z(n1959) );
  NAND U1424 ( .A(n1964), .B(n1965), .Z(n1963) );
  XNOR U1425 ( .A(n1909), .B(n1966), .Z(SUM[66]) );
  OR U1426 ( .A(n1908), .B(n1907), .Z(n1966) );
  NANDN U1427 ( .A(n1967), .B(n1968), .Z(n1909) );
  NAND U1428 ( .A(n1969), .B(n1970), .Z(n1968) );
  XNOR U1429 ( .A(n1964), .B(n1971), .Z(SUM[669]) );
  NANDN U1430 ( .A(n1962), .B(n1965), .Z(n1971) );
  NANDN U1431 ( .A(n1972), .B(n1973), .Z(n1964) );
  NAND U1432 ( .A(n1974), .B(n1975), .Z(n1973) );
  XNOR U1433 ( .A(n1974), .B(n1976), .Z(SUM[668]) );
  NANDN U1434 ( .A(n1972), .B(n1975), .Z(n1976) );
  NANDN U1435 ( .A(n1977), .B(n1978), .Z(n1974) );
  NAND U1436 ( .A(n1979), .B(n1980), .Z(n1978) );
  XOR U1437 ( .A(n1981), .B(n1982), .Z(SUM[667]) );
  NANDN U1438 ( .A(n1983), .B(n1984), .Z(n1982) );
  ANDN U1439 ( .B(n1985), .A(n1986), .Z(n1981) );
  NAND U1440 ( .A(n1987), .B(n1988), .Z(n1985) );
  XNOR U1441 ( .A(n1987), .B(n1989), .Z(SUM[666]) );
  NANDN U1442 ( .A(n1986), .B(n1988), .Z(n1989) );
  NANDN U1443 ( .A(n1990), .B(n1991), .Z(n1987) );
  NAND U1444 ( .A(n1992), .B(n1993), .Z(n1991) );
  XNOR U1445 ( .A(n1992), .B(n1994), .Z(SUM[665]) );
  NANDN U1446 ( .A(n1990), .B(n1993), .Z(n1994) );
  NANDN U1447 ( .A(n1995), .B(n1996), .Z(n1992) );
  NAND U1448 ( .A(n1980), .B(n1997), .Z(n1996) );
  XNOR U1449 ( .A(n1980), .B(n1998), .Z(SUM[664]) );
  NANDN U1450 ( .A(n1995), .B(n1997), .Z(n1998) );
  NANDN U1451 ( .A(n1999), .B(n2000), .Z(n1980) );
  OR U1452 ( .A(n2001), .B(n2002), .Z(n2000) );
  XOR U1453 ( .A(n2003), .B(n2004), .Z(SUM[663]) );
  NANDN U1454 ( .A(n2005), .B(n2006), .Z(n2004) );
  ANDN U1455 ( .B(n2007), .A(n2008), .Z(n2003) );
  NAND U1456 ( .A(n2009), .B(n2010), .Z(n2007) );
  XNOR U1457 ( .A(n2009), .B(n2011), .Z(SUM[662]) );
  NANDN U1458 ( .A(n2008), .B(n2010), .Z(n2011) );
  NANDN U1459 ( .A(n2012), .B(n2013), .Z(n2009) );
  NAND U1460 ( .A(n2014), .B(n2015), .Z(n2013) );
  XNOR U1461 ( .A(n2014), .B(n2016), .Z(SUM[661]) );
  NANDN U1462 ( .A(n2012), .B(n2015), .Z(n2016) );
  NANDN U1463 ( .A(n2017), .B(n2018), .Z(n2014) );
  NANDN U1464 ( .A(n2002), .B(n2019), .Z(n2018) );
  XOR U1465 ( .A(n2002), .B(n2020), .Z(SUM[660]) );
  NANDN U1466 ( .A(n2017), .B(n2019), .Z(n2020) );
  ANDN U1467 ( .B(n2021), .A(n2022), .Z(n2002) );
  OR U1468 ( .A(n2023), .B(n1952), .Z(n2021) );
  XNOR U1469 ( .A(n1969), .B(n2024), .Z(SUM[65]) );
  NANDN U1470 ( .A(n1967), .B(n1970), .Z(n2024) );
  NANDN U1471 ( .A(n2025), .B(n2026), .Z(n1969) );
  NANDN U1472 ( .A(n1847), .B(n2027), .Z(n2026) );
  XOR U1473 ( .A(n2028), .B(n2029), .Z(SUM[659]) );
  NANDN U1474 ( .A(n2030), .B(n2031), .Z(n2029) );
  ANDN U1475 ( .B(n2032), .A(n2033), .Z(n2028) );
  NAND U1476 ( .A(n2034), .B(n2035), .Z(n2032) );
  XNOR U1477 ( .A(n2034), .B(n2036), .Z(SUM[658]) );
  NANDN U1478 ( .A(n2033), .B(n2035), .Z(n2036) );
  NANDN U1479 ( .A(n2037), .B(n2038), .Z(n2034) );
  NAND U1480 ( .A(n2039), .B(n2040), .Z(n2038) );
  XNOR U1481 ( .A(n2039), .B(n2041), .Z(SUM[657]) );
  NANDN U1482 ( .A(n2037), .B(n2040), .Z(n2041) );
  NANDN U1483 ( .A(n2042), .B(n2043), .Z(n2039) );
  NANDN U1484 ( .A(n1952), .B(n2044), .Z(n2043) );
  XOR U1485 ( .A(n1952), .B(n2045), .Z(SUM[656]) );
  NANDN U1486 ( .A(n2042), .B(n2044), .Z(n2045) );
  ANDN U1487 ( .B(n2046), .A(n2047), .Z(n1952) );
  NANDN U1488 ( .A(n2048), .B(n1755), .Z(n2046) );
  XOR U1489 ( .A(n2049), .B(n2050), .Z(SUM[655]) );
  NANDN U1490 ( .A(n2051), .B(n2052), .Z(n2050) );
  ANDN U1491 ( .B(n2053), .A(n2054), .Z(n2049) );
  NAND U1492 ( .A(n2055), .B(n2056), .Z(n2053) );
  XNOR U1493 ( .A(n2055), .B(n2057), .Z(SUM[654]) );
  NANDN U1494 ( .A(n2054), .B(n2056), .Z(n2057) );
  NANDN U1495 ( .A(n2058), .B(n2059), .Z(n2055) );
  NAND U1496 ( .A(n2060), .B(n2061), .Z(n2059) );
  XNOR U1497 ( .A(n2060), .B(n2062), .Z(SUM[653]) );
  NANDN U1498 ( .A(n2058), .B(n2061), .Z(n2062) );
  NANDN U1499 ( .A(n2063), .B(n2064), .Z(n2060) );
  NAND U1500 ( .A(n2065), .B(n2066), .Z(n2064) );
  XNOR U1501 ( .A(n2065), .B(n2067), .Z(SUM[652]) );
  NANDN U1502 ( .A(n2063), .B(n2066), .Z(n2067) );
  NANDN U1503 ( .A(n2068), .B(n2069), .Z(n2065) );
  NAND U1504 ( .A(n2070), .B(n2071), .Z(n2069) );
  XOR U1505 ( .A(n2072), .B(n2073), .Z(SUM[651]) );
  NANDN U1506 ( .A(n2074), .B(n2075), .Z(n2073) );
  ANDN U1507 ( .B(n2076), .A(n2077), .Z(n2072) );
  NAND U1508 ( .A(n2078), .B(n2079), .Z(n2076) );
  XNOR U1509 ( .A(n2078), .B(n2080), .Z(SUM[650]) );
  NANDN U1510 ( .A(n2077), .B(n2079), .Z(n2080) );
  NANDN U1511 ( .A(n2081), .B(n2082), .Z(n2078) );
  NAND U1512 ( .A(n2083), .B(n2084), .Z(n2082) );
  XOR U1513 ( .A(n1847), .B(n2085), .Z(SUM[64]) );
  NANDN U1514 ( .A(n2025), .B(n2027), .Z(n2085) );
  XNOR U1515 ( .A(n2083), .B(n2086), .Z(SUM[649]) );
  NANDN U1516 ( .A(n2081), .B(n2084), .Z(n2086) );
  NANDN U1517 ( .A(n2087), .B(n2088), .Z(n2083) );
  NAND U1518 ( .A(n2071), .B(n2089), .Z(n2088) );
  XNOR U1519 ( .A(n2071), .B(n2090), .Z(SUM[648]) );
  NANDN U1520 ( .A(n2087), .B(n2089), .Z(n2090) );
  NANDN U1521 ( .A(n2091), .B(n2092), .Z(n2071) );
  OR U1522 ( .A(n2093), .B(n2094), .Z(n2092) );
  XOR U1523 ( .A(n2095), .B(n2096), .Z(SUM[647]) );
  NANDN U1524 ( .A(n2097), .B(n2098), .Z(n2096) );
  ANDN U1525 ( .B(n2099), .A(n2100), .Z(n2095) );
  NAND U1526 ( .A(n2101), .B(n2102), .Z(n2099) );
  XNOR U1527 ( .A(n2101), .B(n2103), .Z(SUM[646]) );
  NANDN U1528 ( .A(n2100), .B(n2102), .Z(n2103) );
  NANDN U1529 ( .A(n2104), .B(n2105), .Z(n2101) );
  NAND U1530 ( .A(n2106), .B(n2107), .Z(n2105) );
  XNOR U1531 ( .A(n2106), .B(n2108), .Z(SUM[645]) );
  NANDN U1532 ( .A(n2104), .B(n2107), .Z(n2108) );
  NANDN U1533 ( .A(n2109), .B(n2110), .Z(n2106) );
  NANDN U1534 ( .A(n2094), .B(n2111), .Z(n2110) );
  XOR U1535 ( .A(n2094), .B(n2112), .Z(SUM[644]) );
  NANDN U1536 ( .A(n2109), .B(n2111), .Z(n2112) );
  ANDN U1537 ( .B(n2113), .A(n2114), .Z(n2094) );
  NANDN U1538 ( .A(n2115), .B(n1755), .Z(n2113) );
  XOR U1539 ( .A(n2116), .B(n2117), .Z(SUM[643]) );
  NANDN U1540 ( .A(n2118), .B(n2119), .Z(n2117) );
  ANDN U1541 ( .B(n2120), .A(n2121), .Z(n2116) );
  NAND U1542 ( .A(n2122), .B(n2123), .Z(n2120) );
  XNOR U1543 ( .A(n2122), .B(n2124), .Z(SUM[642]) );
  NANDN U1544 ( .A(n2121), .B(n2123), .Z(n2124) );
  NANDN U1545 ( .A(n2125), .B(n2126), .Z(n2122) );
  NAND U1546 ( .A(n2127), .B(n2128), .Z(n2126) );
  XNOR U1547 ( .A(n2127), .B(n2129), .Z(SUM[641]) );
  NANDN U1548 ( .A(n2125), .B(n2128), .Z(n2129) );
  NANDN U1549 ( .A(n2130), .B(n2131), .Z(n2127) );
  NAND U1550 ( .A(n1755), .B(n2132), .Z(n2131) );
  XNOR U1551 ( .A(n1755), .B(n2133), .Z(SUM[640]) );
  NANDN U1552 ( .A(n2130), .B(n2132), .Z(n2133) );
  NANDN U1553 ( .A(n2134), .B(n2135), .Z(n1755) );
  OR U1554 ( .A(n2136), .B(n2137), .Z(n2135) );
  XOR U1555 ( .A(n2138), .B(n2139), .Z(SUM[63]) );
  OR U1556 ( .A(n2140), .B(n2141), .Z(n2139) );
  ANDN U1557 ( .B(n2142), .A(n2143), .Z(n2138) );
  NANDN U1558 ( .A(n2144), .B(n2145), .Z(n2142) );
  XOR U1559 ( .A(n2146), .B(n2147), .Z(SUM[639]) );
  NANDN U1560 ( .A(n2148), .B(n2149), .Z(n2147) );
  ANDN U1561 ( .B(n2150), .A(n2151), .Z(n2146) );
  NAND U1562 ( .A(n2152), .B(n2153), .Z(n2150) );
  XNOR U1563 ( .A(n2152), .B(n2154), .Z(SUM[638]) );
  NANDN U1564 ( .A(n2151), .B(n2153), .Z(n2154) );
  NANDN U1565 ( .A(n2155), .B(n2156), .Z(n2152) );
  NAND U1566 ( .A(n2157), .B(n2158), .Z(n2156) );
  XNOR U1567 ( .A(n2157), .B(n2159), .Z(SUM[637]) );
  NANDN U1568 ( .A(n2155), .B(n2158), .Z(n2159) );
  NANDN U1569 ( .A(n2160), .B(n2161), .Z(n2157) );
  NAND U1570 ( .A(n2162), .B(n2163), .Z(n2161) );
  XNOR U1571 ( .A(n2162), .B(n2164), .Z(SUM[636]) );
  NANDN U1572 ( .A(n2160), .B(n2163), .Z(n2164) );
  NANDN U1573 ( .A(n2165), .B(n2166), .Z(n2162) );
  NANDN U1574 ( .A(n2167), .B(n2168), .Z(n2166) );
  XOR U1575 ( .A(n2169), .B(n2170), .Z(SUM[635]) );
  NANDN U1576 ( .A(n2171), .B(n2172), .Z(n2170) );
  ANDN U1577 ( .B(n2173), .A(n2174), .Z(n2169) );
  NAND U1578 ( .A(n2175), .B(n2176), .Z(n2173) );
  XNOR U1579 ( .A(n2175), .B(n2177), .Z(SUM[634]) );
  NANDN U1580 ( .A(n2174), .B(n2176), .Z(n2177) );
  NANDN U1581 ( .A(n2178), .B(n2179), .Z(n2175) );
  NAND U1582 ( .A(n2180), .B(n2181), .Z(n2179) );
  XNOR U1583 ( .A(n2180), .B(n2182), .Z(SUM[633]) );
  NANDN U1584 ( .A(n2178), .B(n2181), .Z(n2182) );
  NANDN U1585 ( .A(n2183), .B(n2184), .Z(n2180) );
  NAND U1586 ( .A(n2168), .B(n2185), .Z(n2184) );
  XNOR U1587 ( .A(n2168), .B(n2186), .Z(SUM[632]) );
  NANDN U1588 ( .A(n2183), .B(n2185), .Z(n2186) );
  NANDN U1589 ( .A(n2187), .B(n2188), .Z(n2168) );
  OR U1590 ( .A(n2189), .B(n2190), .Z(n2188) );
  XOR U1591 ( .A(n2191), .B(n2192), .Z(SUM[631]) );
  NANDN U1592 ( .A(n2193), .B(n2194), .Z(n2192) );
  ANDN U1593 ( .B(n2195), .A(n2196), .Z(n2191) );
  NAND U1594 ( .A(n2197), .B(n2198), .Z(n2195) );
  XNOR U1595 ( .A(n2197), .B(n2199), .Z(SUM[630]) );
  NANDN U1596 ( .A(n2196), .B(n2198), .Z(n2199) );
  NANDN U1597 ( .A(n2200), .B(n2201), .Z(n2197) );
  NAND U1598 ( .A(n2202), .B(n2203), .Z(n2201) );
  XNOR U1599 ( .A(n2145), .B(n2204), .Z(SUM[62]) );
  OR U1600 ( .A(n2144), .B(n2143), .Z(n2204) );
  NANDN U1601 ( .A(n2205), .B(n2206), .Z(n2145) );
  NANDN U1602 ( .A(n2207), .B(n2208), .Z(n2206) );
  XNOR U1603 ( .A(n2202), .B(n2209), .Z(SUM[629]) );
  NANDN U1604 ( .A(n2200), .B(n2203), .Z(n2209) );
  NANDN U1605 ( .A(n2210), .B(n2211), .Z(n2202) );
  NANDN U1606 ( .A(n2190), .B(n2212), .Z(n2211) );
  XOR U1607 ( .A(n2190), .B(n2213), .Z(SUM[628]) );
  NANDN U1608 ( .A(n2210), .B(n2212), .Z(n2213) );
  ANDN U1609 ( .B(n2214), .A(n2215), .Z(n2190) );
  NANDN U1610 ( .A(n2216), .B(n2217), .Z(n2214) );
  XOR U1611 ( .A(n2218), .B(n2219), .Z(SUM[627]) );
  NANDN U1612 ( .A(n2220), .B(n2221), .Z(n2219) );
  ANDN U1613 ( .B(n2222), .A(n2223), .Z(n2218) );
  NAND U1614 ( .A(n2224), .B(n2225), .Z(n2222) );
  XNOR U1615 ( .A(n2224), .B(n2226), .Z(SUM[626]) );
  NANDN U1616 ( .A(n2223), .B(n2225), .Z(n2226) );
  NANDN U1617 ( .A(n2227), .B(n2228), .Z(n2224) );
  NAND U1618 ( .A(n2229), .B(n2230), .Z(n2228) );
  XNOR U1619 ( .A(n2229), .B(n2231), .Z(SUM[625]) );
  NANDN U1620 ( .A(n2227), .B(n2230), .Z(n2231) );
  NANDN U1621 ( .A(n2232), .B(n2233), .Z(n2229) );
  NAND U1622 ( .A(n2217), .B(n2234), .Z(n2233) );
  XNOR U1623 ( .A(n2217), .B(n2235), .Z(SUM[624]) );
  NANDN U1624 ( .A(n2232), .B(n2234), .Z(n2235) );
  NANDN U1625 ( .A(n2236), .B(n2237), .Z(n2217) );
  NANDN U1626 ( .A(n2238), .B(n2239), .Z(n2237) );
  XOR U1627 ( .A(n2240), .B(n2241), .Z(SUM[623]) );
  NANDN U1628 ( .A(n2242), .B(n2243), .Z(n2241) );
  ANDN U1629 ( .B(n2244), .A(n2245), .Z(n2240) );
  NAND U1630 ( .A(n2246), .B(n2247), .Z(n2244) );
  XNOR U1631 ( .A(n2246), .B(n2248), .Z(SUM[622]) );
  NANDN U1632 ( .A(n2245), .B(n2247), .Z(n2248) );
  NANDN U1633 ( .A(n2249), .B(n2250), .Z(n2246) );
  NAND U1634 ( .A(n2251), .B(n2252), .Z(n2250) );
  XNOR U1635 ( .A(n2251), .B(n2253), .Z(SUM[621]) );
  NANDN U1636 ( .A(n2249), .B(n2252), .Z(n2253) );
  NANDN U1637 ( .A(n2254), .B(n2255), .Z(n2251) );
  NAND U1638 ( .A(n2256), .B(n2257), .Z(n2255) );
  XNOR U1639 ( .A(n2256), .B(n2258), .Z(SUM[620]) );
  NANDN U1640 ( .A(n2254), .B(n2257), .Z(n2258) );
  NANDN U1641 ( .A(n2259), .B(n2260), .Z(n2256) );
  NANDN U1642 ( .A(n2261), .B(n2262), .Z(n2260) );
  XNOR U1643 ( .A(n2208), .B(n2263), .Z(SUM[61]) );
  OR U1644 ( .A(n2207), .B(n2205), .Z(n2263) );
  NANDN U1645 ( .A(n2264), .B(n2265), .Z(n2208) );
  NANDN U1646 ( .A(n2266), .B(n2267), .Z(n2265) );
  XOR U1647 ( .A(n2268), .B(n2269), .Z(SUM[619]) );
  NANDN U1648 ( .A(n2270), .B(n2271), .Z(n2269) );
  ANDN U1649 ( .B(n2272), .A(n2273), .Z(n2268) );
  NAND U1650 ( .A(n2274), .B(n2275), .Z(n2272) );
  XNOR U1651 ( .A(n2274), .B(n2276), .Z(SUM[618]) );
  NANDN U1652 ( .A(n2273), .B(n2275), .Z(n2276) );
  NANDN U1653 ( .A(n2277), .B(n2278), .Z(n2274) );
  NAND U1654 ( .A(n2279), .B(n2280), .Z(n2278) );
  XNOR U1655 ( .A(n2279), .B(n2281), .Z(SUM[617]) );
  NANDN U1656 ( .A(n2277), .B(n2280), .Z(n2281) );
  NANDN U1657 ( .A(n2282), .B(n2283), .Z(n2279) );
  NAND U1658 ( .A(n2262), .B(n2284), .Z(n2283) );
  XNOR U1659 ( .A(n2262), .B(n2285), .Z(SUM[616]) );
  NANDN U1660 ( .A(n2282), .B(n2284), .Z(n2285) );
  NANDN U1661 ( .A(n2286), .B(n2287), .Z(n2262) );
  OR U1662 ( .A(n2288), .B(n2289), .Z(n2287) );
  XOR U1663 ( .A(n2290), .B(n2291), .Z(SUM[615]) );
  NANDN U1664 ( .A(n2292), .B(n2293), .Z(n2291) );
  ANDN U1665 ( .B(n2294), .A(n2295), .Z(n2290) );
  NAND U1666 ( .A(n2296), .B(n2297), .Z(n2294) );
  XNOR U1667 ( .A(n2296), .B(n2298), .Z(SUM[614]) );
  NANDN U1668 ( .A(n2295), .B(n2297), .Z(n2298) );
  NANDN U1669 ( .A(n2299), .B(n2300), .Z(n2296) );
  NAND U1670 ( .A(n2301), .B(n2302), .Z(n2300) );
  XNOR U1671 ( .A(n2301), .B(n2303), .Z(SUM[613]) );
  NANDN U1672 ( .A(n2299), .B(n2302), .Z(n2303) );
  NANDN U1673 ( .A(n2304), .B(n2305), .Z(n2301) );
  NANDN U1674 ( .A(n2289), .B(n2306), .Z(n2305) );
  XOR U1675 ( .A(n2289), .B(n2307), .Z(SUM[612]) );
  NANDN U1676 ( .A(n2304), .B(n2306), .Z(n2307) );
  ANDN U1677 ( .B(n2308), .A(n2309), .Z(n2289) );
  NANDN U1678 ( .A(n2310), .B(n2239), .Z(n2308) );
  XOR U1679 ( .A(n2311), .B(n2312), .Z(SUM[611]) );
  NANDN U1680 ( .A(n2313), .B(n2314), .Z(n2312) );
  ANDN U1681 ( .B(n2315), .A(n2316), .Z(n2311) );
  NAND U1682 ( .A(n2317), .B(n2318), .Z(n2315) );
  XNOR U1683 ( .A(n2317), .B(n2319), .Z(SUM[610]) );
  NANDN U1684 ( .A(n2316), .B(n2318), .Z(n2319) );
  NANDN U1685 ( .A(n2320), .B(n2321), .Z(n2317) );
  NAND U1686 ( .A(n2322), .B(n2323), .Z(n2321) );
  XNOR U1687 ( .A(n2267), .B(n2324), .Z(SUM[60]) );
  OR U1688 ( .A(n2266), .B(n2264), .Z(n2324) );
  NANDN U1689 ( .A(n2325), .B(n2326), .Z(n2267) );
  NANDN U1690 ( .A(n2327), .B(n2328), .Z(n2326) );
  XNOR U1691 ( .A(n2322), .B(n2329), .Z(SUM[609]) );
  NANDN U1692 ( .A(n2320), .B(n2323), .Z(n2329) );
  NANDN U1693 ( .A(n2330), .B(n2331), .Z(n2322) );
  NAND U1694 ( .A(n2239), .B(n2332), .Z(n2331) );
  XNOR U1695 ( .A(n2239), .B(n2333), .Z(SUM[608]) );
  NANDN U1696 ( .A(n2330), .B(n2332), .Z(n2333) );
  NANDN U1697 ( .A(n2334), .B(n2335), .Z(n2239) );
  OR U1698 ( .A(n2336), .B(n2337), .Z(n2335) );
  XOR U1699 ( .A(n2338), .B(n2339), .Z(SUM[607]) );
  NANDN U1700 ( .A(n2340), .B(n2341), .Z(n2339) );
  ANDN U1701 ( .B(n2342), .A(n2343), .Z(n2338) );
  NAND U1702 ( .A(n2344), .B(n2345), .Z(n2342) );
  XNOR U1703 ( .A(n2344), .B(n2346), .Z(SUM[606]) );
  NANDN U1704 ( .A(n2343), .B(n2345), .Z(n2346) );
  NANDN U1705 ( .A(n2347), .B(n2348), .Z(n2344) );
  NAND U1706 ( .A(n2349), .B(n2350), .Z(n2348) );
  XNOR U1707 ( .A(n2349), .B(n2351), .Z(SUM[605]) );
  NANDN U1708 ( .A(n2347), .B(n2350), .Z(n2351) );
  NANDN U1709 ( .A(n2352), .B(n2353), .Z(n2349) );
  NAND U1710 ( .A(n2354), .B(n2355), .Z(n2353) );
  XNOR U1711 ( .A(n2354), .B(n2356), .Z(SUM[604]) );
  NANDN U1712 ( .A(n2352), .B(n2355), .Z(n2356) );
  NANDN U1713 ( .A(n2357), .B(n2358), .Z(n2354) );
  NANDN U1714 ( .A(n2359), .B(n2360), .Z(n2358) );
  XOR U1715 ( .A(n2361), .B(n2362), .Z(SUM[603]) );
  NANDN U1716 ( .A(n2363), .B(n2364), .Z(n2362) );
  ANDN U1717 ( .B(n2365), .A(n2366), .Z(n2361) );
  NAND U1718 ( .A(n2367), .B(n2368), .Z(n2365) );
  XNOR U1719 ( .A(n2367), .B(n2369), .Z(SUM[602]) );
  NANDN U1720 ( .A(n2366), .B(n2368), .Z(n2369) );
  NANDN U1721 ( .A(n2370), .B(n2371), .Z(n2367) );
  NAND U1722 ( .A(n2372), .B(n2373), .Z(n2371) );
  XNOR U1723 ( .A(n2372), .B(n2374), .Z(SUM[601]) );
  NANDN U1724 ( .A(n2370), .B(n2373), .Z(n2374) );
  NANDN U1725 ( .A(n2375), .B(n2376), .Z(n2372) );
  NAND U1726 ( .A(n2360), .B(n2377), .Z(n2376) );
  XNOR U1727 ( .A(n2360), .B(n2378), .Z(SUM[600]) );
  NANDN U1728 ( .A(n2375), .B(n2377), .Z(n2378) );
  NANDN U1729 ( .A(n2379), .B(n2380), .Z(n2360) );
  OR U1730 ( .A(n2381), .B(n2382), .Z(n2380) );
  XNOR U1731 ( .A(n2383), .B(n2384), .Z(SUM[5]) );
  OR U1732 ( .A(n2385), .B(n2386), .Z(n2384) );
  XOR U1733 ( .A(n2387), .B(n2388), .Z(SUM[59]) );
  NANDN U1734 ( .A(n2389), .B(n2390), .Z(n2388) );
  ANDN U1735 ( .B(n2391), .A(n2392), .Z(n2387) );
  NAND U1736 ( .A(n2393), .B(n2394), .Z(n2391) );
  XOR U1737 ( .A(n2395), .B(n2396), .Z(SUM[599]) );
  NANDN U1738 ( .A(n2397), .B(n2398), .Z(n2396) );
  ANDN U1739 ( .B(n2399), .A(n2400), .Z(n2395) );
  NAND U1740 ( .A(n2401), .B(n2402), .Z(n2399) );
  XNOR U1741 ( .A(n2401), .B(n2403), .Z(SUM[598]) );
  NANDN U1742 ( .A(n2400), .B(n2402), .Z(n2403) );
  NANDN U1743 ( .A(n2404), .B(n2405), .Z(n2401) );
  NAND U1744 ( .A(n2406), .B(n2407), .Z(n2405) );
  XNOR U1745 ( .A(n2406), .B(n2408), .Z(SUM[597]) );
  NANDN U1746 ( .A(n2404), .B(n2407), .Z(n2408) );
  NANDN U1747 ( .A(n2409), .B(n2410), .Z(n2406) );
  NANDN U1748 ( .A(n2382), .B(n2411), .Z(n2410) );
  XOR U1749 ( .A(n2382), .B(n2412), .Z(SUM[596]) );
  NANDN U1750 ( .A(n2409), .B(n2411), .Z(n2412) );
  ANDN U1751 ( .B(n2413), .A(n2414), .Z(n2382) );
  OR U1752 ( .A(n2415), .B(n2337), .Z(n2413) );
  XOR U1753 ( .A(n2416), .B(n2417), .Z(SUM[595]) );
  NANDN U1754 ( .A(n2418), .B(n2419), .Z(n2417) );
  ANDN U1755 ( .B(n2420), .A(n2421), .Z(n2416) );
  NAND U1756 ( .A(n2422), .B(n2423), .Z(n2420) );
  XNOR U1757 ( .A(n2422), .B(n2424), .Z(SUM[594]) );
  NANDN U1758 ( .A(n2421), .B(n2423), .Z(n2424) );
  NANDN U1759 ( .A(n2425), .B(n2426), .Z(n2422) );
  NAND U1760 ( .A(n2427), .B(n2428), .Z(n2426) );
  XNOR U1761 ( .A(n2427), .B(n2429), .Z(SUM[593]) );
  NANDN U1762 ( .A(n2425), .B(n2428), .Z(n2429) );
  NANDN U1763 ( .A(n2430), .B(n2431), .Z(n2427) );
  NANDN U1764 ( .A(n2337), .B(n2432), .Z(n2431) );
  XOR U1765 ( .A(n2337), .B(n2433), .Z(SUM[592]) );
  NANDN U1766 ( .A(n2430), .B(n2432), .Z(n2433) );
  ANDN U1767 ( .B(n2434), .A(n2435), .Z(n2337) );
  OR U1768 ( .A(n2436), .B(n2137), .Z(n2434) );
  XOR U1769 ( .A(n2437), .B(n2438), .Z(SUM[591]) );
  NANDN U1770 ( .A(n2439), .B(n2440), .Z(n2438) );
  ANDN U1771 ( .B(n2441), .A(n2442), .Z(n2437) );
  NAND U1772 ( .A(n2443), .B(n2444), .Z(n2441) );
  XNOR U1773 ( .A(n2443), .B(n2445), .Z(SUM[590]) );
  NANDN U1774 ( .A(n2442), .B(n2444), .Z(n2445) );
  NANDN U1775 ( .A(n2446), .B(n2447), .Z(n2443) );
  NAND U1776 ( .A(n2448), .B(n2449), .Z(n2447) );
  XNOR U1777 ( .A(n2393), .B(n2450), .Z(SUM[58]) );
  NANDN U1778 ( .A(n2392), .B(n2394), .Z(n2450) );
  NANDN U1779 ( .A(n2451), .B(n2452), .Z(n2393) );
  NAND U1780 ( .A(n2453), .B(n2454), .Z(n2452) );
  XNOR U1781 ( .A(n2448), .B(n2455), .Z(SUM[589]) );
  NANDN U1782 ( .A(n2446), .B(n2449), .Z(n2455) );
  NANDN U1783 ( .A(n2456), .B(n2457), .Z(n2448) );
  NAND U1784 ( .A(n2458), .B(n2459), .Z(n2457) );
  XNOR U1785 ( .A(n2458), .B(n2460), .Z(SUM[588]) );
  NANDN U1786 ( .A(n2456), .B(n2459), .Z(n2460) );
  NANDN U1787 ( .A(n2461), .B(n2462), .Z(n2458) );
  NANDN U1788 ( .A(n2463), .B(n2464), .Z(n2462) );
  XOR U1789 ( .A(n2465), .B(n2466), .Z(SUM[587]) );
  NANDN U1790 ( .A(n2467), .B(n2468), .Z(n2466) );
  ANDN U1791 ( .B(n2469), .A(n2470), .Z(n2465) );
  NAND U1792 ( .A(n2471), .B(n2472), .Z(n2469) );
  XNOR U1793 ( .A(n2471), .B(n2473), .Z(SUM[586]) );
  NANDN U1794 ( .A(n2470), .B(n2472), .Z(n2473) );
  NANDN U1795 ( .A(n2474), .B(n2475), .Z(n2471) );
  NAND U1796 ( .A(n2476), .B(n2477), .Z(n2475) );
  XNOR U1797 ( .A(n2476), .B(n2478), .Z(SUM[585]) );
  NANDN U1798 ( .A(n2474), .B(n2477), .Z(n2478) );
  NANDN U1799 ( .A(n2479), .B(n2480), .Z(n2476) );
  NAND U1800 ( .A(n2464), .B(n2481), .Z(n2480) );
  XNOR U1801 ( .A(n2464), .B(n2482), .Z(SUM[584]) );
  NANDN U1802 ( .A(n2479), .B(n2481), .Z(n2482) );
  NANDN U1803 ( .A(n2483), .B(n2484), .Z(n2464) );
  OR U1804 ( .A(n2485), .B(n2486), .Z(n2484) );
  XOR U1805 ( .A(n2487), .B(n2488), .Z(SUM[583]) );
  NANDN U1806 ( .A(n2489), .B(n2490), .Z(n2488) );
  ANDN U1807 ( .B(n2491), .A(n2492), .Z(n2487) );
  NAND U1808 ( .A(n2493), .B(n2494), .Z(n2491) );
  XNOR U1809 ( .A(n2493), .B(n2495), .Z(SUM[582]) );
  NANDN U1810 ( .A(n2492), .B(n2494), .Z(n2495) );
  NANDN U1811 ( .A(n2496), .B(n2497), .Z(n2493) );
  NAND U1812 ( .A(n2498), .B(n2499), .Z(n2497) );
  XNOR U1813 ( .A(n2498), .B(n2500), .Z(SUM[581]) );
  NANDN U1814 ( .A(n2496), .B(n2499), .Z(n2500) );
  NANDN U1815 ( .A(n2501), .B(n2502), .Z(n2498) );
  NANDN U1816 ( .A(n2486), .B(n2503), .Z(n2502) );
  XOR U1817 ( .A(n2486), .B(n2504), .Z(SUM[580]) );
  NANDN U1818 ( .A(n2501), .B(n2503), .Z(n2504) );
  ANDN U1819 ( .B(n2505), .A(n2506), .Z(n2486) );
  OR U1820 ( .A(n2507), .B(n2137), .Z(n2505) );
  XNOR U1821 ( .A(n2453), .B(n2508), .Z(SUM[57]) );
  NANDN U1822 ( .A(n2451), .B(n2454), .Z(n2508) );
  NANDN U1823 ( .A(n2509), .B(n2510), .Z(n2453) );
  NAND U1824 ( .A(n2328), .B(n2511), .Z(n2510) );
  XOR U1825 ( .A(n2512), .B(n2513), .Z(SUM[579]) );
  NANDN U1826 ( .A(n2514), .B(n2515), .Z(n2513) );
  ANDN U1827 ( .B(n2516), .A(n2517), .Z(n2512) );
  NAND U1828 ( .A(n2518), .B(n2519), .Z(n2516) );
  XNOR U1829 ( .A(n2518), .B(n2520), .Z(SUM[578]) );
  NANDN U1830 ( .A(n2517), .B(n2519), .Z(n2520) );
  NANDN U1831 ( .A(n2521), .B(n2522), .Z(n2518) );
  NAND U1832 ( .A(n2523), .B(n2524), .Z(n2522) );
  XNOR U1833 ( .A(n2523), .B(n2525), .Z(SUM[577]) );
  NANDN U1834 ( .A(n2521), .B(n2524), .Z(n2525) );
  NANDN U1835 ( .A(n2526), .B(n2527), .Z(n2523) );
  NANDN U1836 ( .A(n2137), .B(n2528), .Z(n2527) );
  XOR U1837 ( .A(n2137), .B(n2529), .Z(SUM[576]) );
  NANDN U1838 ( .A(n2526), .B(n2528), .Z(n2529) );
  NOR U1839 ( .A(n2530), .B(n2531), .Z(n2137) );
  XOR U1840 ( .A(n2532), .B(n2533), .Z(SUM[575]) );
  NANDN U1841 ( .A(n2534), .B(n2535), .Z(n2533) );
  ANDN U1842 ( .B(n2536), .A(n2537), .Z(n2532) );
  NAND U1843 ( .A(n2538), .B(n2539), .Z(n2536) );
  XNOR U1844 ( .A(n2538), .B(n2540), .Z(SUM[574]) );
  NANDN U1845 ( .A(n2537), .B(n2539), .Z(n2540) );
  NANDN U1846 ( .A(n2541), .B(n2542), .Z(n2538) );
  NAND U1847 ( .A(n2543), .B(n2544), .Z(n2542) );
  XNOR U1848 ( .A(n2543), .B(n2545), .Z(SUM[573]) );
  NANDN U1849 ( .A(n2541), .B(n2544), .Z(n2545) );
  NANDN U1850 ( .A(n2546), .B(n2547), .Z(n2543) );
  NAND U1851 ( .A(n2548), .B(n2549), .Z(n2547) );
  XNOR U1852 ( .A(n2548), .B(n2550), .Z(SUM[572]) );
  NANDN U1853 ( .A(n2546), .B(n2549), .Z(n2550) );
  NANDN U1854 ( .A(n2551), .B(n2552), .Z(n2548) );
  NANDN U1855 ( .A(n2553), .B(n2554), .Z(n2552) );
  XOR U1856 ( .A(n2555), .B(n2556), .Z(SUM[571]) );
  NANDN U1857 ( .A(n2557), .B(n2558), .Z(n2556) );
  ANDN U1858 ( .B(n2559), .A(n2560), .Z(n2555) );
  NAND U1859 ( .A(n2561), .B(n2562), .Z(n2559) );
  XNOR U1860 ( .A(n2561), .B(n2563), .Z(SUM[570]) );
  NANDN U1861 ( .A(n2560), .B(n2562), .Z(n2563) );
  NANDN U1862 ( .A(n2564), .B(n2565), .Z(n2561) );
  NAND U1863 ( .A(n2566), .B(n2567), .Z(n2565) );
  XNOR U1864 ( .A(n2328), .B(n2568), .Z(SUM[56]) );
  NANDN U1865 ( .A(n2509), .B(n2511), .Z(n2568) );
  NANDN U1866 ( .A(n2569), .B(n2570), .Z(n2328) );
  OR U1867 ( .A(n2571), .B(n2572), .Z(n2570) );
  XNOR U1868 ( .A(n2566), .B(n2573), .Z(SUM[569]) );
  NANDN U1869 ( .A(n2564), .B(n2567), .Z(n2573) );
  NANDN U1870 ( .A(n2574), .B(n2575), .Z(n2566) );
  NAND U1871 ( .A(n2554), .B(n2576), .Z(n2575) );
  XNOR U1872 ( .A(n2554), .B(n2577), .Z(SUM[568]) );
  NANDN U1873 ( .A(n2574), .B(n2576), .Z(n2577) );
  NANDN U1874 ( .A(n2578), .B(n2579), .Z(n2554) );
  OR U1875 ( .A(n2580), .B(n2581), .Z(n2579) );
  XOR U1876 ( .A(n2582), .B(n2583), .Z(SUM[567]) );
  NANDN U1877 ( .A(n2584), .B(n2585), .Z(n2583) );
  ANDN U1878 ( .B(n2586), .A(n2587), .Z(n2582) );
  NAND U1879 ( .A(n2588), .B(n2589), .Z(n2586) );
  XNOR U1880 ( .A(n2588), .B(n2590), .Z(SUM[566]) );
  NANDN U1881 ( .A(n2587), .B(n2589), .Z(n2590) );
  NANDN U1882 ( .A(n2591), .B(n2592), .Z(n2588) );
  NAND U1883 ( .A(n2593), .B(n2594), .Z(n2592) );
  XNOR U1884 ( .A(n2593), .B(n2595), .Z(SUM[565]) );
  NANDN U1885 ( .A(n2591), .B(n2594), .Z(n2595) );
  NANDN U1886 ( .A(n2596), .B(n2597), .Z(n2593) );
  NANDN U1887 ( .A(n2581), .B(n2598), .Z(n2597) );
  XOR U1888 ( .A(n2581), .B(n2599), .Z(SUM[564]) );
  NANDN U1889 ( .A(n2596), .B(n2598), .Z(n2599) );
  ANDN U1890 ( .B(n2600), .A(n2601), .Z(n2581) );
  NANDN U1891 ( .A(n2602), .B(n2603), .Z(n2600) );
  XOR U1892 ( .A(n2604), .B(n2605), .Z(SUM[563]) );
  NANDN U1893 ( .A(n2606), .B(n2607), .Z(n2605) );
  ANDN U1894 ( .B(n2608), .A(n2609), .Z(n2604) );
  NAND U1895 ( .A(n2610), .B(n2611), .Z(n2608) );
  XNOR U1896 ( .A(n2610), .B(n2612), .Z(SUM[562]) );
  NANDN U1897 ( .A(n2609), .B(n2611), .Z(n2612) );
  NANDN U1898 ( .A(n2613), .B(n2614), .Z(n2610) );
  NAND U1899 ( .A(n2615), .B(n2616), .Z(n2614) );
  XNOR U1900 ( .A(n2615), .B(n2617), .Z(SUM[561]) );
  NANDN U1901 ( .A(n2613), .B(n2616), .Z(n2617) );
  NANDN U1902 ( .A(n2618), .B(n2619), .Z(n2615) );
  NAND U1903 ( .A(n2603), .B(n2620), .Z(n2619) );
  XNOR U1904 ( .A(n2603), .B(n2621), .Z(SUM[560]) );
  NANDN U1905 ( .A(n2618), .B(n2620), .Z(n2621) );
  NANDN U1906 ( .A(n2622), .B(n2623), .Z(n2603) );
  NANDN U1907 ( .A(n2624), .B(n2625), .Z(n2623) );
  XOR U1908 ( .A(n2626), .B(n2627), .Z(SUM[55]) );
  NANDN U1909 ( .A(n2628), .B(n2629), .Z(n2627) );
  ANDN U1910 ( .B(n2630), .A(n2631), .Z(n2626) );
  NAND U1911 ( .A(n2632), .B(n2633), .Z(n2630) );
  XOR U1912 ( .A(n2634), .B(n2635), .Z(SUM[559]) );
  NANDN U1913 ( .A(n2636), .B(n2637), .Z(n2635) );
  ANDN U1914 ( .B(n2638), .A(n2639), .Z(n2634) );
  NAND U1915 ( .A(n2640), .B(n2641), .Z(n2638) );
  XNOR U1916 ( .A(n2640), .B(n2642), .Z(SUM[558]) );
  NANDN U1917 ( .A(n2639), .B(n2641), .Z(n2642) );
  NANDN U1918 ( .A(n2643), .B(n2644), .Z(n2640) );
  NAND U1919 ( .A(n2645), .B(n2646), .Z(n2644) );
  XNOR U1920 ( .A(n2645), .B(n2647), .Z(SUM[557]) );
  NANDN U1921 ( .A(n2643), .B(n2646), .Z(n2647) );
  NANDN U1922 ( .A(n2648), .B(n2649), .Z(n2645) );
  NAND U1923 ( .A(n2650), .B(n2651), .Z(n2649) );
  XNOR U1924 ( .A(n2650), .B(n2652), .Z(SUM[556]) );
  NANDN U1925 ( .A(n2648), .B(n2651), .Z(n2652) );
  NANDN U1926 ( .A(n2653), .B(n2654), .Z(n2650) );
  NANDN U1927 ( .A(n2655), .B(n2656), .Z(n2654) );
  XOR U1928 ( .A(n2657), .B(n2658), .Z(SUM[555]) );
  NANDN U1929 ( .A(n2659), .B(n2660), .Z(n2658) );
  ANDN U1930 ( .B(n2661), .A(n2662), .Z(n2657) );
  NAND U1931 ( .A(n2663), .B(n2664), .Z(n2661) );
  XNOR U1932 ( .A(n2663), .B(n2665), .Z(SUM[554]) );
  NANDN U1933 ( .A(n2662), .B(n2664), .Z(n2665) );
  NANDN U1934 ( .A(n2666), .B(n2667), .Z(n2663) );
  NAND U1935 ( .A(n2668), .B(n2669), .Z(n2667) );
  XNOR U1936 ( .A(n2668), .B(n2670), .Z(SUM[553]) );
  NANDN U1937 ( .A(n2666), .B(n2669), .Z(n2670) );
  NANDN U1938 ( .A(n2671), .B(n2672), .Z(n2668) );
  NAND U1939 ( .A(n2656), .B(n2673), .Z(n2672) );
  XNOR U1940 ( .A(n2656), .B(n2674), .Z(SUM[552]) );
  NANDN U1941 ( .A(n2671), .B(n2673), .Z(n2674) );
  NANDN U1942 ( .A(n2675), .B(n2676), .Z(n2656) );
  OR U1943 ( .A(n2677), .B(n2678), .Z(n2676) );
  XOR U1944 ( .A(n2679), .B(n2680), .Z(SUM[551]) );
  NANDN U1945 ( .A(n2681), .B(n2682), .Z(n2680) );
  ANDN U1946 ( .B(n2683), .A(n2684), .Z(n2679) );
  NAND U1947 ( .A(n2685), .B(n2686), .Z(n2683) );
  XNOR U1948 ( .A(n2685), .B(n2687), .Z(SUM[550]) );
  NANDN U1949 ( .A(n2684), .B(n2686), .Z(n2687) );
  NANDN U1950 ( .A(n2688), .B(n2689), .Z(n2685) );
  NAND U1951 ( .A(n2690), .B(n2691), .Z(n2689) );
  XNOR U1952 ( .A(n2632), .B(n2692), .Z(SUM[54]) );
  NANDN U1953 ( .A(n2631), .B(n2633), .Z(n2692) );
  NANDN U1954 ( .A(n2693), .B(n2694), .Z(n2632) );
  NAND U1955 ( .A(n2695), .B(n2696), .Z(n2694) );
  XNOR U1956 ( .A(n2690), .B(n2697), .Z(SUM[549]) );
  NANDN U1957 ( .A(n2688), .B(n2691), .Z(n2697) );
  NANDN U1958 ( .A(n2698), .B(n2699), .Z(n2690) );
  NANDN U1959 ( .A(n2678), .B(n2700), .Z(n2699) );
  XOR U1960 ( .A(n2678), .B(n2701), .Z(SUM[548]) );
  NANDN U1961 ( .A(n2698), .B(n2700), .Z(n2701) );
  ANDN U1962 ( .B(n2702), .A(n2703), .Z(n2678) );
  NANDN U1963 ( .A(n2704), .B(n2625), .Z(n2702) );
  XOR U1964 ( .A(n2705), .B(n2706), .Z(SUM[547]) );
  NANDN U1965 ( .A(n2707), .B(n2708), .Z(n2706) );
  ANDN U1966 ( .B(n2709), .A(n2710), .Z(n2705) );
  NAND U1967 ( .A(n2711), .B(n2712), .Z(n2709) );
  XNOR U1968 ( .A(n2711), .B(n2713), .Z(SUM[546]) );
  NANDN U1969 ( .A(n2710), .B(n2712), .Z(n2713) );
  NANDN U1970 ( .A(n2714), .B(n2715), .Z(n2711) );
  NAND U1971 ( .A(n2716), .B(n2717), .Z(n2715) );
  XNOR U1972 ( .A(n2716), .B(n2718), .Z(SUM[545]) );
  NANDN U1973 ( .A(n2714), .B(n2717), .Z(n2718) );
  NANDN U1974 ( .A(n2719), .B(n2720), .Z(n2716) );
  NAND U1975 ( .A(n2625), .B(n2721), .Z(n2720) );
  XNOR U1976 ( .A(n2625), .B(n2722), .Z(SUM[544]) );
  NANDN U1977 ( .A(n2719), .B(n2721), .Z(n2722) );
  NANDN U1978 ( .A(n2723), .B(n2724), .Z(n2625) );
  OR U1979 ( .A(n2725), .B(n2726), .Z(n2724) );
  XOR U1980 ( .A(n2727), .B(n2728), .Z(SUM[543]) );
  NANDN U1981 ( .A(n2729), .B(n2730), .Z(n2728) );
  ANDN U1982 ( .B(n2731), .A(n2732), .Z(n2727) );
  NAND U1983 ( .A(n2733), .B(n2734), .Z(n2731) );
  XNOR U1984 ( .A(n2733), .B(n2735), .Z(SUM[542]) );
  NANDN U1985 ( .A(n2732), .B(n2734), .Z(n2735) );
  NANDN U1986 ( .A(n2736), .B(n2737), .Z(n2733) );
  NAND U1987 ( .A(n2738), .B(n2739), .Z(n2737) );
  XNOR U1988 ( .A(n2738), .B(n2740), .Z(SUM[541]) );
  NANDN U1989 ( .A(n2736), .B(n2739), .Z(n2740) );
  NANDN U1990 ( .A(n2741), .B(n2742), .Z(n2738) );
  NAND U1991 ( .A(n2743), .B(n2744), .Z(n2742) );
  XNOR U1992 ( .A(n2743), .B(n2745), .Z(SUM[540]) );
  NANDN U1993 ( .A(n2741), .B(n2744), .Z(n2745) );
  NANDN U1994 ( .A(n2746), .B(n2747), .Z(n2743) );
  NANDN U1995 ( .A(n2748), .B(n2749), .Z(n2747) );
  XNOR U1996 ( .A(n2695), .B(n2750), .Z(SUM[53]) );
  NANDN U1997 ( .A(n2693), .B(n2696), .Z(n2750) );
  NANDN U1998 ( .A(n2751), .B(n2752), .Z(n2695) );
  NANDN U1999 ( .A(n2572), .B(n2753), .Z(n2752) );
  XOR U2000 ( .A(n2754), .B(n2755), .Z(SUM[539]) );
  NANDN U2001 ( .A(n2756), .B(n2757), .Z(n2755) );
  ANDN U2002 ( .B(n2758), .A(n2759), .Z(n2754) );
  NAND U2003 ( .A(n2760), .B(n2761), .Z(n2758) );
  XNOR U2004 ( .A(n2760), .B(n2762), .Z(SUM[538]) );
  NANDN U2005 ( .A(n2759), .B(n2761), .Z(n2762) );
  NANDN U2006 ( .A(n2763), .B(n2764), .Z(n2760) );
  NAND U2007 ( .A(n2765), .B(n2766), .Z(n2764) );
  XNOR U2008 ( .A(n2765), .B(n2767), .Z(SUM[537]) );
  NANDN U2009 ( .A(n2763), .B(n2766), .Z(n2767) );
  NANDN U2010 ( .A(n2768), .B(n2769), .Z(n2765) );
  NAND U2011 ( .A(n2749), .B(n2770), .Z(n2769) );
  XNOR U2012 ( .A(n2749), .B(n2771), .Z(SUM[536]) );
  NANDN U2013 ( .A(n2768), .B(n2770), .Z(n2771) );
  NANDN U2014 ( .A(n2772), .B(n2773), .Z(n2749) );
  OR U2015 ( .A(n2774), .B(n2775), .Z(n2773) );
  XOR U2016 ( .A(n2776), .B(n2777), .Z(SUM[535]) );
  NANDN U2017 ( .A(n2778), .B(n2779), .Z(n2777) );
  ANDN U2018 ( .B(n2780), .A(n2781), .Z(n2776) );
  NAND U2019 ( .A(n2782), .B(n2783), .Z(n2780) );
  XNOR U2020 ( .A(n2782), .B(n2784), .Z(SUM[534]) );
  NANDN U2021 ( .A(n2781), .B(n2783), .Z(n2784) );
  NANDN U2022 ( .A(n2785), .B(n2786), .Z(n2782) );
  NAND U2023 ( .A(n2787), .B(n2788), .Z(n2786) );
  XNOR U2024 ( .A(n2787), .B(n2789), .Z(SUM[533]) );
  NANDN U2025 ( .A(n2785), .B(n2788), .Z(n2789) );
  NANDN U2026 ( .A(n2790), .B(n2791), .Z(n2787) );
  NANDN U2027 ( .A(n2775), .B(n2792), .Z(n2791) );
  XOR U2028 ( .A(n2775), .B(n2793), .Z(SUM[532]) );
  NANDN U2029 ( .A(n2790), .B(n2792), .Z(n2793) );
  ANDN U2030 ( .B(n2794), .A(n2795), .Z(n2775) );
  OR U2031 ( .A(n2796), .B(n2726), .Z(n2794) );
  XOR U2032 ( .A(n2797), .B(n2798), .Z(SUM[531]) );
  NANDN U2033 ( .A(n2799), .B(n2800), .Z(n2798) );
  ANDN U2034 ( .B(n2801), .A(n2802), .Z(n2797) );
  NAND U2035 ( .A(n2803), .B(n2804), .Z(n2801) );
  XNOR U2036 ( .A(n2803), .B(n2805), .Z(SUM[530]) );
  NANDN U2037 ( .A(n2802), .B(n2804), .Z(n2805) );
  NANDN U2038 ( .A(n2806), .B(n2807), .Z(n2803) );
  NAND U2039 ( .A(n2808), .B(n2809), .Z(n2807) );
  XOR U2040 ( .A(n2572), .B(n2810), .Z(SUM[52]) );
  NANDN U2041 ( .A(n2751), .B(n2753), .Z(n2810) );
  NOR U2042 ( .A(n2811), .B(n2812), .Z(n2572) );
  XNOR U2043 ( .A(n2808), .B(n2813), .Z(SUM[529]) );
  NANDN U2044 ( .A(n2806), .B(n2809), .Z(n2813) );
  NANDN U2045 ( .A(n2814), .B(n2815), .Z(n2808) );
  NANDN U2046 ( .A(n2726), .B(n2816), .Z(n2815) );
  XOR U2047 ( .A(n2726), .B(n2817), .Z(SUM[528]) );
  NANDN U2048 ( .A(n2814), .B(n2816), .Z(n2817) );
  ANDN U2049 ( .B(n2818), .A(n2819), .Z(n2726) );
  OR U2050 ( .A(n2820), .B(n2821), .Z(n2818) );
  XOR U2051 ( .A(n2822), .B(n2823), .Z(SUM[527]) );
  NANDN U2052 ( .A(n2824), .B(n2825), .Z(n2823) );
  ANDN U2053 ( .B(n2826), .A(n2827), .Z(n2822) );
  NAND U2054 ( .A(n2828), .B(n2829), .Z(n2826) );
  XNOR U2055 ( .A(n2828), .B(n2830), .Z(SUM[526]) );
  NANDN U2056 ( .A(n2827), .B(n2829), .Z(n2830) );
  NANDN U2057 ( .A(n2831), .B(n2832), .Z(n2828) );
  NAND U2058 ( .A(n2833), .B(n2834), .Z(n2832) );
  XNOR U2059 ( .A(n2833), .B(n2835), .Z(SUM[525]) );
  NANDN U2060 ( .A(n2831), .B(n2834), .Z(n2835) );
  NANDN U2061 ( .A(n2836), .B(n2837), .Z(n2833) );
  NAND U2062 ( .A(n2838), .B(n2839), .Z(n2837) );
  XNOR U2063 ( .A(n2838), .B(n2840), .Z(SUM[524]) );
  NANDN U2064 ( .A(n2836), .B(n2839), .Z(n2840) );
  NANDN U2065 ( .A(n2841), .B(n2842), .Z(n2838) );
  NANDN U2066 ( .A(n2843), .B(n2844), .Z(n2842) );
  XOR U2067 ( .A(n2845), .B(n2846), .Z(SUM[523]) );
  NANDN U2068 ( .A(n2847), .B(n2848), .Z(n2846) );
  ANDN U2069 ( .B(n2849), .A(n2850), .Z(n2845) );
  NAND U2070 ( .A(n2851), .B(n2852), .Z(n2849) );
  XNOR U2071 ( .A(n2851), .B(n2853), .Z(SUM[522]) );
  NANDN U2072 ( .A(n2850), .B(n2852), .Z(n2853) );
  NANDN U2073 ( .A(n2854), .B(n2855), .Z(n2851) );
  NAND U2074 ( .A(n2856), .B(n2857), .Z(n2855) );
  XNOR U2075 ( .A(n2856), .B(n2858), .Z(SUM[521]) );
  NANDN U2076 ( .A(n2854), .B(n2857), .Z(n2858) );
  NANDN U2077 ( .A(n2859), .B(n2860), .Z(n2856) );
  NAND U2078 ( .A(n2844), .B(n2861), .Z(n2860) );
  XNOR U2079 ( .A(n2844), .B(n2862), .Z(SUM[520]) );
  NANDN U2080 ( .A(n2859), .B(n2861), .Z(n2862) );
  NANDN U2081 ( .A(n2863), .B(n2864), .Z(n2844) );
  OR U2082 ( .A(n2865), .B(n2866), .Z(n2864) );
  XOR U2083 ( .A(n2867), .B(n2868), .Z(SUM[51]) );
  NANDN U2084 ( .A(n2869), .B(n2870), .Z(n2868) );
  ANDN U2085 ( .B(n2871), .A(n2872), .Z(n2867) );
  NAND U2086 ( .A(n2873), .B(n2874), .Z(n2871) );
  XOR U2087 ( .A(n2875), .B(n2876), .Z(SUM[519]) );
  NANDN U2088 ( .A(n2877), .B(n2878), .Z(n2876) );
  ANDN U2089 ( .B(n2879), .A(n2880), .Z(n2875) );
  NAND U2090 ( .A(n2881), .B(n2882), .Z(n2879) );
  XNOR U2091 ( .A(n2881), .B(n2883), .Z(SUM[518]) );
  NANDN U2092 ( .A(n2880), .B(n2882), .Z(n2883) );
  NANDN U2093 ( .A(n2884), .B(n2885), .Z(n2881) );
  NAND U2094 ( .A(n2886), .B(n2887), .Z(n2885) );
  XNOR U2095 ( .A(n2886), .B(n2888), .Z(SUM[517]) );
  NANDN U2096 ( .A(n2884), .B(n2887), .Z(n2888) );
  NANDN U2097 ( .A(n2889), .B(n2890), .Z(n2886) );
  NANDN U2098 ( .A(n2866), .B(n2891), .Z(n2890) );
  XOR U2099 ( .A(n2866), .B(n2892), .Z(SUM[516]) );
  NANDN U2100 ( .A(n2889), .B(n2891), .Z(n2892) );
  ANDN U2101 ( .B(n2893), .A(n2894), .Z(n2866) );
  OR U2102 ( .A(n2895), .B(n2821), .Z(n2893) );
  XOR U2103 ( .A(n2896), .B(n2897), .Z(SUM[515]) );
  NANDN U2104 ( .A(n2898), .B(n2899), .Z(n2897) );
  ANDN U2105 ( .B(n2900), .A(n2901), .Z(n2896) );
  NAND U2106 ( .A(n2902), .B(n2903), .Z(n2900) );
  XNOR U2107 ( .A(n2902), .B(n2904), .Z(SUM[514]) );
  NANDN U2108 ( .A(n2901), .B(n2903), .Z(n2904) );
  NANDN U2109 ( .A(n2905), .B(n2906), .Z(n2902) );
  NAND U2110 ( .A(n2907), .B(n2908), .Z(n2906) );
  XNOR U2111 ( .A(n2907), .B(n2909), .Z(SUM[513]) );
  NANDN U2112 ( .A(n2905), .B(n2908), .Z(n2909) );
  NANDN U2113 ( .A(n2910), .B(n2911), .Z(n2907) );
  NANDN U2114 ( .A(n2821), .B(n2912), .Z(n2911) );
  XOR U2115 ( .A(n2821), .B(n2913), .Z(SUM[512]) );
  NANDN U2116 ( .A(n2910), .B(n2912), .Z(n2913) );
  XOR U2117 ( .A(n2914), .B(n2915), .Z(SUM[511]) );
  OR U2118 ( .A(n2916), .B(n2917), .Z(n2915) );
  ANDN U2119 ( .B(n2918), .A(n2919), .Z(n2914) );
  NAND U2120 ( .A(n2920), .B(n2921), .Z(n2918) );
  XNOR U2121 ( .A(n2920), .B(n2922), .Z(SUM[510]) );
  NANDN U2122 ( .A(n2919), .B(n2921), .Z(n2922) );
  NANDN U2123 ( .A(n2923), .B(n2924), .Z(n2920) );
  NAND U2124 ( .A(n2925), .B(n2926), .Z(n2924) );
  XNOR U2125 ( .A(n2873), .B(n2927), .Z(SUM[50]) );
  NANDN U2126 ( .A(n2872), .B(n2874), .Z(n2927) );
  NANDN U2127 ( .A(n2928), .B(n2929), .Z(n2873) );
  NAND U2128 ( .A(n2930), .B(n2931), .Z(n2929) );
  XNOR U2129 ( .A(n2925), .B(n2932), .Z(SUM[509]) );
  NANDN U2130 ( .A(n2923), .B(n2926), .Z(n2932) );
  NANDN U2131 ( .A(n2933), .B(n2934), .Z(n2925) );
  NANDN U2132 ( .A(n2935), .B(n2936), .Z(n2934) );
  XNOR U2133 ( .A(n2936), .B(n2937), .Z(SUM[508]) );
  OR U2134 ( .A(n2935), .B(n2933), .Z(n2937) );
  NANDN U2135 ( .A(n2938), .B(n2939), .Z(n2936) );
  NANDN U2136 ( .A(n2940), .B(n2941), .Z(n2939) );
  XOR U2137 ( .A(n2942), .B(n2943), .Z(SUM[507]) );
  NANDN U2138 ( .A(n2944), .B(n2945), .Z(n2943) );
  ANDN U2139 ( .B(n2946), .A(n2947), .Z(n2942) );
  NAND U2140 ( .A(n2948), .B(n2949), .Z(n2946) );
  XNOR U2141 ( .A(n2948), .B(n2950), .Z(SUM[506]) );
  NANDN U2142 ( .A(n2947), .B(n2949), .Z(n2950) );
  NANDN U2143 ( .A(n2951), .B(n2952), .Z(n2948) );
  NAND U2144 ( .A(n2953), .B(n2954), .Z(n2952) );
  XNOR U2145 ( .A(n2953), .B(n2955), .Z(SUM[505]) );
  NANDN U2146 ( .A(n2951), .B(n2954), .Z(n2955) );
  NANDN U2147 ( .A(n2956), .B(n2957), .Z(n2953) );
  NAND U2148 ( .A(n2941), .B(n2958), .Z(n2957) );
  XNOR U2149 ( .A(n2941), .B(n2959), .Z(SUM[504]) );
  NANDN U2150 ( .A(n2956), .B(n2958), .Z(n2959) );
  NANDN U2151 ( .A(n2960), .B(n2961), .Z(n2941) );
  NANDN U2152 ( .A(n2962), .B(n2963), .Z(n2961) );
  XOR U2153 ( .A(n2964), .B(n2965), .Z(SUM[503]) );
  NANDN U2154 ( .A(n2966), .B(n2967), .Z(n2965) );
  ANDN U2155 ( .B(n2968), .A(n2969), .Z(n2964) );
  NAND U2156 ( .A(n2970), .B(n2971), .Z(n2968) );
  XNOR U2157 ( .A(n2970), .B(n2972), .Z(SUM[502]) );
  NANDN U2158 ( .A(n2969), .B(n2971), .Z(n2972) );
  NANDN U2159 ( .A(n2973), .B(n2974), .Z(n2970) );
  NAND U2160 ( .A(n2975), .B(n2976), .Z(n2974) );
  XNOR U2161 ( .A(n2975), .B(n2977), .Z(SUM[501]) );
  NANDN U2162 ( .A(n2973), .B(n2976), .Z(n2977) );
  NANDN U2163 ( .A(n2978), .B(n2979), .Z(n2975) );
  NANDN U2164 ( .A(n2962), .B(n2980), .Z(n2979) );
  XOR U2165 ( .A(n2962), .B(n2981), .Z(SUM[500]) );
  NANDN U2166 ( .A(n2978), .B(n2980), .Z(n2981) );
  ANDN U2167 ( .B(n2982), .A(n2983), .Z(n2962) );
  NANDN U2168 ( .A(n2984), .B(n2985), .Z(n2982) );
  XOR U2169 ( .A(n2986), .B(n2987), .Z(SUM[4]) );
  ANDN U2170 ( .B(n2988), .A(n2989), .Z(n2987) );
  XNOR U2171 ( .A(n2930), .B(n2990), .Z(SUM[49]) );
  NANDN U2172 ( .A(n2928), .B(n2931), .Z(n2990) );
  NANDN U2173 ( .A(n2991), .B(n2992), .Z(n2930) );
  NANDN U2174 ( .A(n2993), .B(n2994), .Z(n2992) );
  XOR U2175 ( .A(n2995), .B(n2996), .Z(SUM[499]) );
  NANDN U2176 ( .A(n2997), .B(n2998), .Z(n2996) );
  ANDN U2177 ( .B(n2999), .A(n3000), .Z(n2995) );
  NANDN U2178 ( .A(n3001), .B(n3002), .Z(n2999) );
  XNOR U2179 ( .A(n3002), .B(n3003), .Z(SUM[498]) );
  OR U2180 ( .A(n3001), .B(n3000), .Z(n3003) );
  NANDN U2181 ( .A(n3004), .B(n3005), .Z(n3002) );
  NAND U2182 ( .A(n3006), .B(n3007), .Z(n3005) );
  XNOR U2183 ( .A(n3006), .B(n3008), .Z(SUM[497]) );
  NANDN U2184 ( .A(n3004), .B(n3007), .Z(n3008) );
  NANDN U2185 ( .A(n3009), .B(n3010), .Z(n3006) );
  NAND U2186 ( .A(n2985), .B(n3011), .Z(n3010) );
  XNOR U2187 ( .A(n2985), .B(n3012), .Z(SUM[496]) );
  NANDN U2188 ( .A(n3009), .B(n3011), .Z(n3012) );
  NANDN U2189 ( .A(n3013), .B(n3014), .Z(n2985) );
  NANDN U2190 ( .A(n3015), .B(n3016), .Z(n3014) );
  XOR U2191 ( .A(n3017), .B(n3018), .Z(SUM[495]) );
  NANDN U2192 ( .A(n3019), .B(n3020), .Z(n3018) );
  ANDN U2193 ( .B(n3021), .A(n3022), .Z(n3017) );
  NAND U2194 ( .A(n3023), .B(n3024), .Z(n3021) );
  XNOR U2195 ( .A(n3023), .B(n3025), .Z(SUM[494]) );
  NANDN U2196 ( .A(n3022), .B(n3024), .Z(n3025) );
  NANDN U2197 ( .A(n3026), .B(n3027), .Z(n3023) );
  NAND U2198 ( .A(n3028), .B(n3029), .Z(n3027) );
  XNOR U2199 ( .A(n3028), .B(n3030), .Z(SUM[493]) );
  NANDN U2200 ( .A(n3026), .B(n3029), .Z(n3030) );
  NANDN U2201 ( .A(n3031), .B(n3032), .Z(n3028) );
  NAND U2202 ( .A(n3033), .B(n3034), .Z(n3032) );
  XNOR U2203 ( .A(n3033), .B(n3035), .Z(SUM[492]) );
  NANDN U2204 ( .A(n3031), .B(n3034), .Z(n3035) );
  NANDN U2205 ( .A(n3036), .B(n3037), .Z(n3033) );
  NAND U2206 ( .A(n3038), .B(n3039), .Z(n3037) );
  XOR U2207 ( .A(n3040), .B(n3041), .Z(SUM[491]) );
  NANDN U2208 ( .A(n3042), .B(n3043), .Z(n3041) );
  ANDN U2209 ( .B(n3044), .A(n3045), .Z(n3040) );
  NAND U2210 ( .A(n3046), .B(n3047), .Z(n3044) );
  XNOR U2211 ( .A(n3046), .B(n3048), .Z(SUM[490]) );
  NANDN U2212 ( .A(n3045), .B(n3047), .Z(n3048) );
  NANDN U2213 ( .A(n3049), .B(n3050), .Z(n3046) );
  NAND U2214 ( .A(n3051), .B(n3052), .Z(n3050) );
  XOR U2215 ( .A(n2993), .B(n3053), .Z(SUM[48]) );
  NANDN U2216 ( .A(n2991), .B(n2994), .Z(n3053) );
  XNOR U2217 ( .A(n3051), .B(n3054), .Z(SUM[489]) );
  NANDN U2218 ( .A(n3049), .B(n3052), .Z(n3054) );
  NANDN U2219 ( .A(n3055), .B(n3056), .Z(n3051) );
  NAND U2220 ( .A(n3039), .B(n3057), .Z(n3056) );
  XNOR U2221 ( .A(n3039), .B(n3058), .Z(SUM[488]) );
  NANDN U2222 ( .A(n3055), .B(n3057), .Z(n3058) );
  NANDN U2223 ( .A(n3059), .B(n3060), .Z(n3039) );
  OR U2224 ( .A(n3061), .B(n3062), .Z(n3060) );
  XOR U2225 ( .A(n3063), .B(n3064), .Z(SUM[487]) );
  NANDN U2226 ( .A(n3065), .B(n3066), .Z(n3064) );
  ANDN U2227 ( .B(n3067), .A(n3068), .Z(n3063) );
  NAND U2228 ( .A(n3069), .B(n3070), .Z(n3067) );
  XNOR U2229 ( .A(n3069), .B(n3071), .Z(SUM[486]) );
  NANDN U2230 ( .A(n3068), .B(n3070), .Z(n3071) );
  NANDN U2231 ( .A(n3072), .B(n3073), .Z(n3069) );
  NAND U2232 ( .A(n3074), .B(n3075), .Z(n3073) );
  XNOR U2233 ( .A(n3074), .B(n3076), .Z(SUM[485]) );
  NANDN U2234 ( .A(n3072), .B(n3075), .Z(n3076) );
  NANDN U2235 ( .A(n3077), .B(n3078), .Z(n3074) );
  NANDN U2236 ( .A(n3062), .B(n3079), .Z(n3078) );
  XOR U2237 ( .A(n3062), .B(n3080), .Z(SUM[484]) );
  NANDN U2238 ( .A(n3077), .B(n3079), .Z(n3080) );
  ANDN U2239 ( .B(n3081), .A(n3082), .Z(n3062) );
  NANDN U2240 ( .A(n3083), .B(n3016), .Z(n3081) );
  XOR U2241 ( .A(n3084), .B(n3085), .Z(SUM[483]) );
  NANDN U2242 ( .A(n3086), .B(n3087), .Z(n3085) );
  ANDN U2243 ( .B(n3088), .A(n3089), .Z(n3084) );
  NAND U2244 ( .A(n3090), .B(n3091), .Z(n3088) );
  XNOR U2245 ( .A(n3090), .B(n3092), .Z(SUM[482]) );
  NANDN U2246 ( .A(n3089), .B(n3091), .Z(n3092) );
  NANDN U2247 ( .A(n3093), .B(n3094), .Z(n3090) );
  NAND U2248 ( .A(n3095), .B(n3096), .Z(n3094) );
  XNOR U2249 ( .A(n3095), .B(n3097), .Z(SUM[481]) );
  NANDN U2250 ( .A(n3093), .B(n3096), .Z(n3097) );
  NANDN U2251 ( .A(n3098), .B(n3099), .Z(n3095) );
  NAND U2252 ( .A(n3016), .B(n3100), .Z(n3099) );
  XNOR U2253 ( .A(n3016), .B(n3101), .Z(SUM[480]) );
  NANDN U2254 ( .A(n3098), .B(n3100), .Z(n3101) );
  NANDN U2255 ( .A(n3102), .B(n3103), .Z(n3016) );
  NANDN U2256 ( .A(n3104), .B(n3105), .Z(n3103) );
  XOR U2257 ( .A(n3106), .B(n3107), .Z(SUM[47]) );
  OR U2258 ( .A(n3108), .B(n3109), .Z(n3107) );
  ANDN U2259 ( .B(n3110), .A(n3111), .Z(n3106) );
  NANDN U2260 ( .A(n3112), .B(n3113), .Z(n3110) );
  XOR U2261 ( .A(n3114), .B(n3115), .Z(SUM[479]) );
  NANDN U2262 ( .A(n3116), .B(n3117), .Z(n3115) );
  ANDN U2263 ( .B(n3118), .A(n3119), .Z(n3114) );
  NAND U2264 ( .A(n3120), .B(n3121), .Z(n3118) );
  XNOR U2265 ( .A(n3120), .B(n3122), .Z(SUM[478]) );
  NANDN U2266 ( .A(n3119), .B(n3121), .Z(n3122) );
  NANDN U2267 ( .A(n3123), .B(n3124), .Z(n3120) );
  NAND U2268 ( .A(n3125), .B(n3126), .Z(n3124) );
  XNOR U2269 ( .A(n3125), .B(n3127), .Z(SUM[477]) );
  NANDN U2270 ( .A(n3123), .B(n3126), .Z(n3127) );
  NANDN U2271 ( .A(n3128), .B(n3129), .Z(n3125) );
  NAND U2272 ( .A(n3130), .B(n3131), .Z(n3129) );
  XNOR U2273 ( .A(n3130), .B(n3132), .Z(SUM[476]) );
  NANDN U2274 ( .A(n3128), .B(n3131), .Z(n3132) );
  NANDN U2275 ( .A(n3133), .B(n3134), .Z(n3130) );
  NAND U2276 ( .A(n3135), .B(n3136), .Z(n3134) );
  XOR U2277 ( .A(n3137), .B(n3138), .Z(SUM[475]) );
  NANDN U2278 ( .A(n3139), .B(n3140), .Z(n3138) );
  ANDN U2279 ( .B(n3141), .A(n3142), .Z(n3137) );
  NAND U2280 ( .A(n3143), .B(n3144), .Z(n3141) );
  XNOR U2281 ( .A(n3143), .B(n3145), .Z(SUM[474]) );
  NANDN U2282 ( .A(n3142), .B(n3144), .Z(n3145) );
  NANDN U2283 ( .A(n3146), .B(n3147), .Z(n3143) );
  NAND U2284 ( .A(n3148), .B(n3149), .Z(n3147) );
  XNOR U2285 ( .A(n3148), .B(n3150), .Z(SUM[473]) );
  NANDN U2286 ( .A(n3146), .B(n3149), .Z(n3150) );
  NANDN U2287 ( .A(n3151), .B(n3152), .Z(n3148) );
  NAND U2288 ( .A(n3136), .B(n3153), .Z(n3152) );
  XNOR U2289 ( .A(n3136), .B(n3154), .Z(SUM[472]) );
  NANDN U2290 ( .A(n3151), .B(n3153), .Z(n3154) );
  NANDN U2291 ( .A(n3155), .B(n3156), .Z(n3136) );
  OR U2292 ( .A(n3157), .B(n3158), .Z(n3156) );
  XOR U2293 ( .A(n3159), .B(n3160), .Z(SUM[471]) );
  NANDN U2294 ( .A(n3161), .B(n3162), .Z(n3160) );
  ANDN U2295 ( .B(n3163), .A(n3164), .Z(n3159) );
  NAND U2296 ( .A(n3165), .B(n3166), .Z(n3163) );
  XNOR U2297 ( .A(n3165), .B(n3167), .Z(SUM[470]) );
  NANDN U2298 ( .A(n3164), .B(n3166), .Z(n3167) );
  NANDN U2299 ( .A(n3168), .B(n3169), .Z(n3165) );
  NAND U2300 ( .A(n3170), .B(n3171), .Z(n3169) );
  XNOR U2301 ( .A(n3113), .B(n3172), .Z(SUM[46]) );
  OR U2302 ( .A(n3112), .B(n3111), .Z(n3172) );
  NANDN U2303 ( .A(n3173), .B(n3174), .Z(n3113) );
  NANDN U2304 ( .A(n3175), .B(n3176), .Z(n3174) );
  XNOR U2305 ( .A(n3170), .B(n3177), .Z(SUM[469]) );
  NANDN U2306 ( .A(n3168), .B(n3171), .Z(n3177) );
  NANDN U2307 ( .A(n3178), .B(n3179), .Z(n3170) );
  NANDN U2308 ( .A(n3158), .B(n3180), .Z(n3179) );
  XOR U2309 ( .A(n3158), .B(n3181), .Z(SUM[468]) );
  NANDN U2310 ( .A(n3178), .B(n3180), .Z(n3181) );
  ANDN U2311 ( .B(n3182), .A(n3183), .Z(n3158) );
  NANDN U2312 ( .A(n3184), .B(n3105), .Z(n3182) );
  XOR U2313 ( .A(n3185), .B(n3186), .Z(SUM[467]) );
  NANDN U2314 ( .A(n3187), .B(n3188), .Z(n3186) );
  ANDN U2315 ( .B(n3189), .A(n3190), .Z(n3185) );
  NAND U2316 ( .A(n3191), .B(n3192), .Z(n3189) );
  XNOR U2317 ( .A(n3191), .B(n3193), .Z(SUM[466]) );
  NANDN U2318 ( .A(n3190), .B(n3192), .Z(n3193) );
  NANDN U2319 ( .A(n3194), .B(n3195), .Z(n3191) );
  NAND U2320 ( .A(n3196), .B(n3197), .Z(n3195) );
  XNOR U2321 ( .A(n3196), .B(n3198), .Z(SUM[465]) );
  NANDN U2322 ( .A(n3194), .B(n3197), .Z(n3198) );
  NANDN U2323 ( .A(n3199), .B(n3200), .Z(n3196) );
  NAND U2324 ( .A(n3105), .B(n3201), .Z(n3200) );
  XNOR U2325 ( .A(n3105), .B(n3202), .Z(SUM[464]) );
  NANDN U2326 ( .A(n3199), .B(n3201), .Z(n3202) );
  NANDN U2327 ( .A(n3203), .B(n3204), .Z(n3105) );
  NANDN U2328 ( .A(n3205), .B(n3206), .Z(n3204) );
  XOR U2329 ( .A(n3207), .B(n3208), .Z(SUM[463]) );
  NANDN U2330 ( .A(n3209), .B(n3210), .Z(n3208) );
  ANDN U2331 ( .B(n3211), .A(n3212), .Z(n3207) );
  NAND U2332 ( .A(n3213), .B(n3214), .Z(n3211) );
  XNOR U2333 ( .A(n3213), .B(n3215), .Z(SUM[462]) );
  NANDN U2334 ( .A(n3212), .B(n3214), .Z(n3215) );
  NANDN U2335 ( .A(n3216), .B(n3217), .Z(n3213) );
  NAND U2336 ( .A(n3218), .B(n3219), .Z(n3217) );
  XNOR U2337 ( .A(n3218), .B(n3220), .Z(SUM[461]) );
  NANDN U2338 ( .A(n3216), .B(n3219), .Z(n3220) );
  NANDN U2339 ( .A(n3221), .B(n3222), .Z(n3218) );
  NAND U2340 ( .A(n3223), .B(n3224), .Z(n3222) );
  XNOR U2341 ( .A(n3223), .B(n3225), .Z(SUM[460]) );
  NANDN U2342 ( .A(n3221), .B(n3224), .Z(n3225) );
  NANDN U2343 ( .A(n3226), .B(n3227), .Z(n3223) );
  NAND U2344 ( .A(n3228), .B(n3229), .Z(n3227) );
  XNOR U2345 ( .A(n3176), .B(n3230), .Z(SUM[45]) );
  OR U2346 ( .A(n3175), .B(n3173), .Z(n3230) );
  NANDN U2347 ( .A(n3231), .B(n3232), .Z(n3176) );
  NAND U2348 ( .A(n3233), .B(n3234), .Z(n3232) );
  XOR U2349 ( .A(n3235), .B(n3236), .Z(SUM[459]) );
  NANDN U2350 ( .A(n3237), .B(n3238), .Z(n3236) );
  ANDN U2351 ( .B(n3239), .A(n3240), .Z(n3235) );
  NAND U2352 ( .A(n3241), .B(n3242), .Z(n3239) );
  XNOR U2353 ( .A(n3241), .B(n3243), .Z(SUM[458]) );
  NANDN U2354 ( .A(n3240), .B(n3242), .Z(n3243) );
  NANDN U2355 ( .A(n3244), .B(n3245), .Z(n3241) );
  NAND U2356 ( .A(n3246), .B(n3247), .Z(n3245) );
  XNOR U2357 ( .A(n3246), .B(n3248), .Z(SUM[457]) );
  NANDN U2358 ( .A(n3244), .B(n3247), .Z(n3248) );
  NANDN U2359 ( .A(n3249), .B(n3250), .Z(n3246) );
  NAND U2360 ( .A(n3229), .B(n3251), .Z(n3250) );
  XNOR U2361 ( .A(n3229), .B(n3252), .Z(SUM[456]) );
  NANDN U2362 ( .A(n3249), .B(n3251), .Z(n3252) );
  NANDN U2363 ( .A(n3253), .B(n3254), .Z(n3229) );
  OR U2364 ( .A(n3255), .B(n3256), .Z(n3254) );
  XOR U2365 ( .A(n3257), .B(n3258), .Z(SUM[455]) );
  NANDN U2366 ( .A(n3259), .B(n3260), .Z(n3258) );
  ANDN U2367 ( .B(n3261), .A(n3262), .Z(n3257) );
  NAND U2368 ( .A(n3263), .B(n3264), .Z(n3261) );
  XNOR U2369 ( .A(n3263), .B(n3265), .Z(SUM[454]) );
  NANDN U2370 ( .A(n3262), .B(n3264), .Z(n3265) );
  NANDN U2371 ( .A(n3266), .B(n3267), .Z(n3263) );
  NAND U2372 ( .A(n3268), .B(n3269), .Z(n3267) );
  XNOR U2373 ( .A(n3268), .B(n3270), .Z(SUM[453]) );
  NANDN U2374 ( .A(n3266), .B(n3269), .Z(n3270) );
  NANDN U2375 ( .A(n3271), .B(n3272), .Z(n3268) );
  NANDN U2376 ( .A(n3256), .B(n3273), .Z(n3272) );
  XOR U2377 ( .A(n3256), .B(n3274), .Z(SUM[452]) );
  NANDN U2378 ( .A(n3271), .B(n3273), .Z(n3274) );
  ANDN U2379 ( .B(n3275), .A(n3276), .Z(n3256) );
  NANDN U2380 ( .A(n3277), .B(n3206), .Z(n3275) );
  XOR U2381 ( .A(n3278), .B(n3279), .Z(SUM[451]) );
  NANDN U2382 ( .A(n3280), .B(n3281), .Z(n3279) );
  ANDN U2383 ( .B(n3282), .A(n3283), .Z(n3278) );
  NAND U2384 ( .A(n3284), .B(n3285), .Z(n3282) );
  XNOR U2385 ( .A(n3284), .B(n3286), .Z(SUM[450]) );
  NANDN U2386 ( .A(n3283), .B(n3285), .Z(n3286) );
  NANDN U2387 ( .A(n3287), .B(n3288), .Z(n3284) );
  NAND U2388 ( .A(n3289), .B(n3290), .Z(n3288) );
  XNOR U2389 ( .A(n3233), .B(n3291), .Z(SUM[44]) );
  NANDN U2390 ( .A(n3231), .B(n3234), .Z(n3291) );
  NANDN U2391 ( .A(n3292), .B(n3293), .Z(n3233) );
  NANDN U2392 ( .A(n3294), .B(n3295), .Z(n3293) );
  XNOR U2393 ( .A(n3289), .B(n3296), .Z(SUM[449]) );
  NANDN U2394 ( .A(n3287), .B(n3290), .Z(n3296) );
  NANDN U2395 ( .A(n3297), .B(n3298), .Z(n3289) );
  NAND U2396 ( .A(n3206), .B(n3299), .Z(n3298) );
  XNOR U2397 ( .A(n3206), .B(n3300), .Z(SUM[448]) );
  NANDN U2398 ( .A(n3297), .B(n3299), .Z(n3300) );
  NANDN U2399 ( .A(n3301), .B(n3302), .Z(n3206) );
  NANDN U2400 ( .A(n3303), .B(n3304), .Z(n3302) );
  XOR U2401 ( .A(n3305), .B(n3306), .Z(SUM[447]) );
  NANDN U2402 ( .A(n3307), .B(n3308), .Z(n3306) );
  ANDN U2403 ( .B(n3309), .A(n3310), .Z(n3305) );
  NAND U2404 ( .A(n3311), .B(n3312), .Z(n3309) );
  XNOR U2405 ( .A(n3311), .B(n3313), .Z(SUM[446]) );
  NANDN U2406 ( .A(n3310), .B(n3312), .Z(n3313) );
  NANDN U2407 ( .A(n3314), .B(n3315), .Z(n3311) );
  NAND U2408 ( .A(n3316), .B(n3317), .Z(n3315) );
  XNOR U2409 ( .A(n3316), .B(n3318), .Z(SUM[445]) );
  NANDN U2410 ( .A(n3314), .B(n3317), .Z(n3318) );
  NANDN U2411 ( .A(n3319), .B(n3320), .Z(n3316) );
  NAND U2412 ( .A(n3321), .B(n3322), .Z(n3320) );
  XNOR U2413 ( .A(n3321), .B(n3323), .Z(SUM[444]) );
  NANDN U2414 ( .A(n3319), .B(n3322), .Z(n3323) );
  NANDN U2415 ( .A(n3324), .B(n3325), .Z(n3321) );
  NANDN U2416 ( .A(n3326), .B(n3327), .Z(n3325) );
  XOR U2417 ( .A(n3328), .B(n3329), .Z(SUM[443]) );
  NANDN U2418 ( .A(n3330), .B(n3331), .Z(n3329) );
  ANDN U2419 ( .B(n3332), .A(n3333), .Z(n3328) );
  NAND U2420 ( .A(n3334), .B(n3335), .Z(n3332) );
  XNOR U2421 ( .A(n3334), .B(n3336), .Z(SUM[442]) );
  NANDN U2422 ( .A(n3333), .B(n3335), .Z(n3336) );
  NANDN U2423 ( .A(n3337), .B(n3338), .Z(n3334) );
  NAND U2424 ( .A(n3339), .B(n3340), .Z(n3338) );
  XNOR U2425 ( .A(n3339), .B(n3341), .Z(SUM[441]) );
  NANDN U2426 ( .A(n3337), .B(n3340), .Z(n3341) );
  NANDN U2427 ( .A(n3342), .B(n3343), .Z(n3339) );
  NAND U2428 ( .A(n3327), .B(n3344), .Z(n3343) );
  XNOR U2429 ( .A(n3327), .B(n3345), .Z(SUM[440]) );
  NANDN U2430 ( .A(n3342), .B(n3344), .Z(n3345) );
  NANDN U2431 ( .A(n3346), .B(n3347), .Z(n3327) );
  OR U2432 ( .A(n3348), .B(n3349), .Z(n3347) );
  XOR U2433 ( .A(n3350), .B(n3351), .Z(SUM[43]) );
  NANDN U2434 ( .A(n3352), .B(n3353), .Z(n3351) );
  ANDN U2435 ( .B(n3354), .A(n3355), .Z(n3350) );
  NAND U2436 ( .A(n3356), .B(n3357), .Z(n3354) );
  XOR U2437 ( .A(n3358), .B(n3359), .Z(SUM[439]) );
  NANDN U2438 ( .A(n3360), .B(n3361), .Z(n3359) );
  ANDN U2439 ( .B(n3362), .A(n3363), .Z(n3358) );
  NAND U2440 ( .A(n3364), .B(n3365), .Z(n3362) );
  XNOR U2441 ( .A(n3364), .B(n3366), .Z(SUM[438]) );
  NANDN U2442 ( .A(n3363), .B(n3365), .Z(n3366) );
  NANDN U2443 ( .A(n3367), .B(n3368), .Z(n3364) );
  NAND U2444 ( .A(n3369), .B(n3370), .Z(n3368) );
  XNOR U2445 ( .A(n3369), .B(n3371), .Z(SUM[437]) );
  NANDN U2446 ( .A(n3367), .B(n3370), .Z(n3371) );
  NANDN U2447 ( .A(n3372), .B(n3373), .Z(n3369) );
  NANDN U2448 ( .A(n3349), .B(n3374), .Z(n3373) );
  XOR U2449 ( .A(n3349), .B(n3375), .Z(SUM[436]) );
  NANDN U2450 ( .A(n3372), .B(n3374), .Z(n3375) );
  ANDN U2451 ( .B(n3376), .A(n3377), .Z(n3349) );
  NANDN U2452 ( .A(n3378), .B(n3379), .Z(n3376) );
  XOR U2453 ( .A(n3380), .B(n3381), .Z(SUM[435]) );
  NANDN U2454 ( .A(n3382), .B(n3383), .Z(n3381) );
  ANDN U2455 ( .B(n3384), .A(n3385), .Z(n3380) );
  NAND U2456 ( .A(n3386), .B(n3387), .Z(n3384) );
  XNOR U2457 ( .A(n3386), .B(n3388), .Z(SUM[434]) );
  NANDN U2458 ( .A(n3385), .B(n3387), .Z(n3388) );
  NANDN U2459 ( .A(n3389), .B(n3390), .Z(n3386) );
  NAND U2460 ( .A(n3391), .B(n3392), .Z(n3390) );
  XNOR U2461 ( .A(n3391), .B(n3393), .Z(SUM[433]) );
  NANDN U2462 ( .A(n3389), .B(n3392), .Z(n3393) );
  NANDN U2463 ( .A(n3394), .B(n3395), .Z(n3391) );
  NAND U2464 ( .A(n3379), .B(n3396), .Z(n3395) );
  XNOR U2465 ( .A(n3379), .B(n3397), .Z(SUM[432]) );
  NANDN U2466 ( .A(n3394), .B(n3396), .Z(n3397) );
  NANDN U2467 ( .A(n3398), .B(n3399), .Z(n3379) );
  NAND U2468 ( .A(n3400), .B(n3401), .Z(n3399) );
  XOR U2469 ( .A(n3402), .B(n3403), .Z(SUM[431]) );
  NANDN U2470 ( .A(n3404), .B(n3405), .Z(n3403) );
  ANDN U2471 ( .B(n3406), .A(n3407), .Z(n3402) );
  NAND U2472 ( .A(n3408), .B(n3409), .Z(n3406) );
  XNOR U2473 ( .A(n3408), .B(n3410), .Z(SUM[430]) );
  NANDN U2474 ( .A(n3407), .B(n3409), .Z(n3410) );
  NANDN U2475 ( .A(n3411), .B(n3412), .Z(n3408) );
  NAND U2476 ( .A(n3413), .B(n3414), .Z(n3412) );
  XNOR U2477 ( .A(n3356), .B(n3415), .Z(SUM[42]) );
  NANDN U2478 ( .A(n3355), .B(n3357), .Z(n3415) );
  NANDN U2479 ( .A(n3416), .B(n3417), .Z(n3356) );
  NAND U2480 ( .A(n3418), .B(n3419), .Z(n3417) );
  XNOR U2481 ( .A(n3413), .B(n3420), .Z(SUM[429]) );
  NANDN U2482 ( .A(n3411), .B(n3414), .Z(n3420) );
  NANDN U2483 ( .A(n3421), .B(n3422), .Z(n3413) );
  NAND U2484 ( .A(n3423), .B(n3424), .Z(n3422) );
  XNOR U2485 ( .A(n3423), .B(n3425), .Z(SUM[428]) );
  NANDN U2486 ( .A(n3421), .B(n3424), .Z(n3425) );
  NANDN U2487 ( .A(n3426), .B(n3427), .Z(n3423) );
  NAND U2488 ( .A(n3428), .B(n3429), .Z(n3427) );
  XOR U2489 ( .A(n3430), .B(n3431), .Z(SUM[427]) );
  NANDN U2490 ( .A(n3432), .B(n3433), .Z(n3431) );
  ANDN U2491 ( .B(n3434), .A(n3435), .Z(n3430) );
  NAND U2492 ( .A(n3436), .B(n3437), .Z(n3434) );
  XNOR U2493 ( .A(n3436), .B(n3438), .Z(SUM[426]) );
  NANDN U2494 ( .A(n3435), .B(n3437), .Z(n3438) );
  NANDN U2495 ( .A(n3439), .B(n3440), .Z(n3436) );
  NAND U2496 ( .A(n3441), .B(n3442), .Z(n3440) );
  XNOR U2497 ( .A(n3441), .B(n3443), .Z(SUM[425]) );
  NANDN U2498 ( .A(n3439), .B(n3442), .Z(n3443) );
  NANDN U2499 ( .A(n3444), .B(n3445), .Z(n3441) );
  NAND U2500 ( .A(n3429), .B(n3446), .Z(n3445) );
  XNOR U2501 ( .A(n3429), .B(n3447), .Z(SUM[424]) );
  NANDN U2502 ( .A(n3444), .B(n3446), .Z(n3447) );
  NANDN U2503 ( .A(n3448), .B(n3449), .Z(n3429) );
  OR U2504 ( .A(n3450), .B(n3451), .Z(n3449) );
  XOR U2505 ( .A(n3452), .B(n3453), .Z(SUM[423]) );
  NANDN U2506 ( .A(n3454), .B(n3455), .Z(n3453) );
  ANDN U2507 ( .B(n3456), .A(n3457), .Z(n3452) );
  NAND U2508 ( .A(n3458), .B(n3459), .Z(n3456) );
  XNOR U2509 ( .A(n3458), .B(n3460), .Z(SUM[422]) );
  NANDN U2510 ( .A(n3457), .B(n3459), .Z(n3460) );
  NANDN U2511 ( .A(n3461), .B(n3462), .Z(n3458) );
  NAND U2512 ( .A(n3463), .B(n3464), .Z(n3462) );
  XNOR U2513 ( .A(n3463), .B(n3465), .Z(SUM[421]) );
  NANDN U2514 ( .A(n3461), .B(n3464), .Z(n3465) );
  NANDN U2515 ( .A(n3466), .B(n3467), .Z(n3463) );
  NANDN U2516 ( .A(n3451), .B(n3468), .Z(n3467) );
  XOR U2517 ( .A(n3451), .B(n3469), .Z(SUM[420]) );
  NANDN U2518 ( .A(n3466), .B(n3468), .Z(n3469) );
  ANDN U2519 ( .B(n3470), .A(n3471), .Z(n3451) );
  NANDN U2520 ( .A(n3472), .B(n3401), .Z(n3470) );
  XNOR U2521 ( .A(n3418), .B(n3473), .Z(SUM[41]) );
  NANDN U2522 ( .A(n3416), .B(n3419), .Z(n3473) );
  NANDN U2523 ( .A(n3474), .B(n3475), .Z(n3418) );
  NAND U2524 ( .A(n3295), .B(n3476), .Z(n3475) );
  XOR U2525 ( .A(n3477), .B(n3478), .Z(SUM[419]) );
  NANDN U2526 ( .A(n3479), .B(n3480), .Z(n3478) );
  ANDN U2527 ( .B(n3481), .A(n3482), .Z(n3477) );
  NAND U2528 ( .A(n3483), .B(n3484), .Z(n3481) );
  XNOR U2529 ( .A(n3483), .B(n3485), .Z(SUM[418]) );
  NANDN U2530 ( .A(n3482), .B(n3484), .Z(n3485) );
  NANDN U2531 ( .A(n3486), .B(n3487), .Z(n3483) );
  NAND U2532 ( .A(n3488), .B(n3489), .Z(n3487) );
  XNOR U2533 ( .A(n3488), .B(n3490), .Z(SUM[417]) );
  NANDN U2534 ( .A(n3486), .B(n3489), .Z(n3490) );
  NANDN U2535 ( .A(n3491), .B(n3492), .Z(n3488) );
  NAND U2536 ( .A(n3401), .B(n3493), .Z(n3492) );
  XNOR U2537 ( .A(n3401), .B(n3494), .Z(SUM[416]) );
  NANDN U2538 ( .A(n3491), .B(n3493), .Z(n3494) );
  NANDN U2539 ( .A(n3495), .B(n3496), .Z(n3401) );
  OR U2540 ( .A(n3497), .B(n3498), .Z(n3496) );
  XOR U2541 ( .A(n3499), .B(n3500), .Z(SUM[415]) );
  NANDN U2542 ( .A(n3501), .B(n3502), .Z(n3500) );
  ANDN U2543 ( .B(n3503), .A(n3504), .Z(n3499) );
  NAND U2544 ( .A(n3505), .B(n3506), .Z(n3503) );
  XNOR U2545 ( .A(n3505), .B(n3507), .Z(SUM[414]) );
  NANDN U2546 ( .A(n3504), .B(n3506), .Z(n3507) );
  NANDN U2547 ( .A(n3508), .B(n3509), .Z(n3505) );
  NAND U2548 ( .A(n3510), .B(n3511), .Z(n3509) );
  XNOR U2549 ( .A(n3510), .B(n3512), .Z(SUM[413]) );
  NANDN U2550 ( .A(n3508), .B(n3511), .Z(n3512) );
  NANDN U2551 ( .A(n3513), .B(n3514), .Z(n3510) );
  NAND U2552 ( .A(n3515), .B(n3516), .Z(n3514) );
  XNOR U2553 ( .A(n3515), .B(n3517), .Z(SUM[412]) );
  NANDN U2554 ( .A(n3513), .B(n3516), .Z(n3517) );
  NANDN U2555 ( .A(n3518), .B(n3519), .Z(n3515) );
  NAND U2556 ( .A(n3520), .B(n3521), .Z(n3519) );
  XOR U2557 ( .A(n3522), .B(n3523), .Z(SUM[411]) );
  NANDN U2558 ( .A(n3524), .B(n3525), .Z(n3523) );
  ANDN U2559 ( .B(n3526), .A(n3527), .Z(n3522) );
  NAND U2560 ( .A(n3528), .B(n3529), .Z(n3526) );
  XNOR U2561 ( .A(n3528), .B(n3530), .Z(SUM[410]) );
  NANDN U2562 ( .A(n3527), .B(n3529), .Z(n3530) );
  NANDN U2563 ( .A(n3531), .B(n3532), .Z(n3528) );
  NAND U2564 ( .A(n3533), .B(n3534), .Z(n3532) );
  XNOR U2565 ( .A(n3295), .B(n3535), .Z(SUM[40]) );
  NANDN U2566 ( .A(n3474), .B(n3476), .Z(n3535) );
  NANDN U2567 ( .A(n3536), .B(n3537), .Z(n3295) );
  NANDN U2568 ( .A(n3538), .B(n3539), .Z(n3537) );
  XNOR U2569 ( .A(n3533), .B(n3540), .Z(SUM[409]) );
  NANDN U2570 ( .A(n3531), .B(n3534), .Z(n3540) );
  NANDN U2571 ( .A(n3541), .B(n3542), .Z(n3533) );
  NAND U2572 ( .A(n3521), .B(n3543), .Z(n3542) );
  XNOR U2573 ( .A(n3521), .B(n3544), .Z(SUM[408]) );
  NANDN U2574 ( .A(n3541), .B(n3543), .Z(n3544) );
  NANDN U2575 ( .A(n3545), .B(n3546), .Z(n3521) );
  OR U2576 ( .A(n3547), .B(n3548), .Z(n3546) );
  XOR U2577 ( .A(n3549), .B(n3550), .Z(SUM[407]) );
  NANDN U2578 ( .A(n3551), .B(n3552), .Z(n3550) );
  ANDN U2579 ( .B(n3553), .A(n3554), .Z(n3549) );
  NAND U2580 ( .A(n3555), .B(n3556), .Z(n3553) );
  XNOR U2581 ( .A(n3555), .B(n3557), .Z(SUM[406]) );
  NANDN U2582 ( .A(n3554), .B(n3556), .Z(n3557) );
  NANDN U2583 ( .A(n3558), .B(n3559), .Z(n3555) );
  NAND U2584 ( .A(n3560), .B(n3561), .Z(n3559) );
  XNOR U2585 ( .A(n3560), .B(n3562), .Z(SUM[405]) );
  NANDN U2586 ( .A(n3558), .B(n3561), .Z(n3562) );
  NANDN U2587 ( .A(n3563), .B(n3564), .Z(n3560) );
  NANDN U2588 ( .A(n3548), .B(n3565), .Z(n3564) );
  XOR U2589 ( .A(n3548), .B(n3566), .Z(SUM[404]) );
  NANDN U2590 ( .A(n3563), .B(n3565), .Z(n3566) );
  ANDN U2591 ( .B(n3567), .A(n3568), .Z(n3548) );
  OR U2592 ( .A(n3569), .B(n3498), .Z(n3567) );
  XOR U2593 ( .A(n3570), .B(n3571), .Z(SUM[403]) );
  NANDN U2594 ( .A(n3572), .B(n3573), .Z(n3571) );
  ANDN U2595 ( .B(n3574), .A(n3575), .Z(n3570) );
  NAND U2596 ( .A(n3576), .B(n3577), .Z(n3574) );
  XNOR U2597 ( .A(n3576), .B(n3578), .Z(SUM[402]) );
  NANDN U2598 ( .A(n3575), .B(n3577), .Z(n3578) );
  NANDN U2599 ( .A(n3579), .B(n3580), .Z(n3576) );
  NAND U2600 ( .A(n3581), .B(n3582), .Z(n3580) );
  XNOR U2601 ( .A(n3581), .B(n3583), .Z(SUM[401]) );
  NANDN U2602 ( .A(n3579), .B(n3582), .Z(n3583) );
  NANDN U2603 ( .A(n3584), .B(n3585), .Z(n3581) );
  NANDN U2604 ( .A(n3498), .B(n3586), .Z(n3585) );
  XOR U2605 ( .A(n3498), .B(n3587), .Z(SUM[400]) );
  NANDN U2606 ( .A(n3584), .B(n3586), .Z(n3587) );
  ANDN U2607 ( .B(n3588), .A(n3589), .Z(n3498) );
  NANDN U2608 ( .A(n3590), .B(n3304), .Z(n3588) );
  ANDN U2609 ( .B(n3591), .A(n2986), .Z(SUM[3]) );
  OR U2610 ( .A(A[3]), .B(B[3]), .Z(n3591) );
  XOR U2611 ( .A(n3592), .B(n3593), .Z(SUM[39]) );
  NANDN U2612 ( .A(n3594), .B(n3595), .Z(n3593) );
  ANDN U2613 ( .B(n3596), .A(n3597), .Z(n3592) );
  NAND U2614 ( .A(n3598), .B(n3599), .Z(n3596) );
  XOR U2615 ( .A(n3600), .B(n3601), .Z(SUM[399]) );
  NANDN U2616 ( .A(n3602), .B(n3603), .Z(n3601) );
  ANDN U2617 ( .B(n3604), .A(n3605), .Z(n3600) );
  NAND U2618 ( .A(n3606), .B(n3607), .Z(n3604) );
  XNOR U2619 ( .A(n3606), .B(n3608), .Z(SUM[398]) );
  NANDN U2620 ( .A(n3605), .B(n3607), .Z(n3608) );
  NANDN U2621 ( .A(n3609), .B(n3610), .Z(n3606) );
  NAND U2622 ( .A(n3611), .B(n3612), .Z(n3610) );
  XNOR U2623 ( .A(n3611), .B(n3613), .Z(SUM[397]) );
  NANDN U2624 ( .A(n3609), .B(n3612), .Z(n3613) );
  NANDN U2625 ( .A(n3614), .B(n3615), .Z(n3611) );
  NAND U2626 ( .A(n3616), .B(n3617), .Z(n3615) );
  XNOR U2627 ( .A(n3616), .B(n3618), .Z(SUM[396]) );
  NANDN U2628 ( .A(n3614), .B(n3617), .Z(n3618) );
  NANDN U2629 ( .A(n3619), .B(n3620), .Z(n3616) );
  NAND U2630 ( .A(n3621), .B(n3622), .Z(n3620) );
  XOR U2631 ( .A(n3623), .B(n3624), .Z(SUM[395]) );
  NANDN U2632 ( .A(n3625), .B(n3626), .Z(n3624) );
  ANDN U2633 ( .B(n3627), .A(n3628), .Z(n3623) );
  NAND U2634 ( .A(n3629), .B(n3630), .Z(n3627) );
  XNOR U2635 ( .A(n3629), .B(n3631), .Z(SUM[394]) );
  NANDN U2636 ( .A(n3628), .B(n3630), .Z(n3631) );
  NANDN U2637 ( .A(n3632), .B(n3633), .Z(n3629) );
  NAND U2638 ( .A(n3634), .B(n3635), .Z(n3633) );
  XNOR U2639 ( .A(n3634), .B(n3636), .Z(SUM[393]) );
  NANDN U2640 ( .A(n3632), .B(n3635), .Z(n3636) );
  NANDN U2641 ( .A(n3637), .B(n3638), .Z(n3634) );
  NAND U2642 ( .A(n3622), .B(n3639), .Z(n3638) );
  XNOR U2643 ( .A(n3622), .B(n3640), .Z(SUM[392]) );
  NANDN U2644 ( .A(n3637), .B(n3639), .Z(n3640) );
  NANDN U2645 ( .A(n3641), .B(n3642), .Z(n3622) );
  OR U2646 ( .A(n3643), .B(n3644), .Z(n3642) );
  XOR U2647 ( .A(n3645), .B(n3646), .Z(SUM[391]) );
  NANDN U2648 ( .A(n3647), .B(n3648), .Z(n3646) );
  ANDN U2649 ( .B(n3649), .A(n3650), .Z(n3645) );
  NAND U2650 ( .A(n3651), .B(n3652), .Z(n3649) );
  XNOR U2651 ( .A(n3651), .B(n3653), .Z(SUM[390]) );
  NANDN U2652 ( .A(n3650), .B(n3652), .Z(n3653) );
  NANDN U2653 ( .A(n3654), .B(n3655), .Z(n3651) );
  NAND U2654 ( .A(n3656), .B(n3657), .Z(n3655) );
  XNOR U2655 ( .A(n3598), .B(n3658), .Z(SUM[38]) );
  NANDN U2656 ( .A(n3597), .B(n3599), .Z(n3658) );
  NANDN U2657 ( .A(n3659), .B(n3660), .Z(n3598) );
  NAND U2658 ( .A(n3661), .B(n3662), .Z(n3660) );
  XNOR U2659 ( .A(n3656), .B(n3663), .Z(SUM[389]) );
  NANDN U2660 ( .A(n3654), .B(n3657), .Z(n3663) );
  NANDN U2661 ( .A(n3664), .B(n3665), .Z(n3656) );
  NANDN U2662 ( .A(n3644), .B(n3666), .Z(n3665) );
  XOR U2663 ( .A(n3644), .B(n3667), .Z(SUM[388]) );
  NANDN U2664 ( .A(n3664), .B(n3666), .Z(n3667) );
  ANDN U2665 ( .B(n3668), .A(n3669), .Z(n3644) );
  NANDN U2666 ( .A(n3670), .B(n3304), .Z(n3668) );
  XOR U2667 ( .A(n3671), .B(n3672), .Z(SUM[387]) );
  NANDN U2668 ( .A(n3673), .B(n3674), .Z(n3672) );
  ANDN U2669 ( .B(n3675), .A(n3676), .Z(n3671) );
  NAND U2670 ( .A(n3677), .B(n3678), .Z(n3675) );
  XNOR U2671 ( .A(n3677), .B(n3679), .Z(SUM[386]) );
  NANDN U2672 ( .A(n3676), .B(n3678), .Z(n3679) );
  NANDN U2673 ( .A(n3680), .B(n3681), .Z(n3677) );
  NAND U2674 ( .A(n3682), .B(n3683), .Z(n3681) );
  XNOR U2675 ( .A(n3682), .B(n3684), .Z(SUM[385]) );
  NANDN U2676 ( .A(n3680), .B(n3683), .Z(n3684) );
  NANDN U2677 ( .A(n3685), .B(n3686), .Z(n3682) );
  NAND U2678 ( .A(n3304), .B(n3687), .Z(n3686) );
  XNOR U2679 ( .A(n3304), .B(n3688), .Z(SUM[384]) );
  NANDN U2680 ( .A(n3685), .B(n3687), .Z(n3688) );
  NANDN U2681 ( .A(n3689), .B(n3690), .Z(n3304) );
  OR U2682 ( .A(n3691), .B(n3692), .Z(n3690) );
  XOR U2683 ( .A(n3693), .B(n3694), .Z(SUM[383]) );
  NANDN U2684 ( .A(n3695), .B(n3696), .Z(n3694) );
  ANDN U2685 ( .B(n3697), .A(n3698), .Z(n3693) );
  NAND U2686 ( .A(n3699), .B(n3700), .Z(n3697) );
  XNOR U2687 ( .A(n3699), .B(n3701), .Z(SUM[382]) );
  NANDN U2688 ( .A(n3698), .B(n3700), .Z(n3701) );
  NANDN U2689 ( .A(n3702), .B(n3703), .Z(n3699) );
  NAND U2690 ( .A(n3704), .B(n3705), .Z(n3703) );
  XNOR U2691 ( .A(n3704), .B(n3706), .Z(SUM[381]) );
  NANDN U2692 ( .A(n3702), .B(n3705), .Z(n3706) );
  NANDN U2693 ( .A(n3707), .B(n3708), .Z(n3704) );
  NAND U2694 ( .A(n3709), .B(n3710), .Z(n3708) );
  XNOR U2695 ( .A(n3709), .B(n3711), .Z(SUM[380]) );
  NANDN U2696 ( .A(n3707), .B(n3710), .Z(n3711) );
  NANDN U2697 ( .A(n3712), .B(n3713), .Z(n3709) );
  NANDN U2698 ( .A(n3714), .B(n3715), .Z(n3713) );
  XNOR U2699 ( .A(n3661), .B(n3716), .Z(SUM[37]) );
  NANDN U2700 ( .A(n3659), .B(n3662), .Z(n3716) );
  NANDN U2701 ( .A(n3717), .B(n3718), .Z(n3661) );
  NANDN U2702 ( .A(n3538), .B(n3719), .Z(n3718) );
  XOR U2703 ( .A(n3720), .B(n3721), .Z(SUM[379]) );
  NANDN U2704 ( .A(n3722), .B(n3723), .Z(n3721) );
  ANDN U2705 ( .B(n3724), .A(n3725), .Z(n3720) );
  NAND U2706 ( .A(n3726), .B(n3727), .Z(n3724) );
  XNOR U2707 ( .A(n3726), .B(n3728), .Z(SUM[378]) );
  NANDN U2708 ( .A(n3725), .B(n3727), .Z(n3728) );
  NANDN U2709 ( .A(n3729), .B(n3730), .Z(n3726) );
  NAND U2710 ( .A(n3731), .B(n3732), .Z(n3730) );
  XNOR U2711 ( .A(n3731), .B(n3733), .Z(SUM[377]) );
  NANDN U2712 ( .A(n3729), .B(n3732), .Z(n3733) );
  NANDN U2713 ( .A(n3734), .B(n3735), .Z(n3731) );
  NAND U2714 ( .A(n3715), .B(n3736), .Z(n3735) );
  XNOR U2715 ( .A(n3715), .B(n3737), .Z(SUM[376]) );
  NANDN U2716 ( .A(n3734), .B(n3736), .Z(n3737) );
  NANDN U2717 ( .A(n3738), .B(n3739), .Z(n3715) );
  OR U2718 ( .A(n3740), .B(n3741), .Z(n3739) );
  XOR U2719 ( .A(n3742), .B(n3743), .Z(SUM[375]) );
  NANDN U2720 ( .A(n3744), .B(n3745), .Z(n3743) );
  ANDN U2721 ( .B(n3746), .A(n3747), .Z(n3742) );
  NAND U2722 ( .A(n3748), .B(n3749), .Z(n3746) );
  XNOR U2723 ( .A(n3748), .B(n3750), .Z(SUM[374]) );
  NANDN U2724 ( .A(n3747), .B(n3749), .Z(n3750) );
  NANDN U2725 ( .A(n3751), .B(n3752), .Z(n3748) );
  NAND U2726 ( .A(n3753), .B(n3754), .Z(n3752) );
  XNOR U2727 ( .A(n3753), .B(n3755), .Z(SUM[373]) );
  NANDN U2728 ( .A(n3751), .B(n3754), .Z(n3755) );
  NANDN U2729 ( .A(n3756), .B(n3757), .Z(n3753) );
  NANDN U2730 ( .A(n3741), .B(n3758), .Z(n3757) );
  XOR U2731 ( .A(n3741), .B(n3759), .Z(SUM[372]) );
  NANDN U2732 ( .A(n3756), .B(n3758), .Z(n3759) );
  ANDN U2733 ( .B(n3760), .A(n3761), .Z(n3741) );
  NANDN U2734 ( .A(n3762), .B(n3763), .Z(n3760) );
  XOR U2735 ( .A(n3764), .B(n3765), .Z(SUM[371]) );
  NANDN U2736 ( .A(n3766), .B(n3767), .Z(n3765) );
  ANDN U2737 ( .B(n3768), .A(n3769), .Z(n3764) );
  NAND U2738 ( .A(n3770), .B(n3771), .Z(n3768) );
  XNOR U2739 ( .A(n3770), .B(n3772), .Z(SUM[370]) );
  NANDN U2740 ( .A(n3769), .B(n3771), .Z(n3772) );
  NANDN U2741 ( .A(n3773), .B(n3774), .Z(n3770) );
  NAND U2742 ( .A(n3775), .B(n3776), .Z(n3774) );
  XOR U2743 ( .A(n3538), .B(n3777), .Z(SUM[36]) );
  NANDN U2744 ( .A(n3717), .B(n3719), .Z(n3777) );
  ANDN U2745 ( .B(n3778), .A(n3779), .Z(n3538) );
  OR U2746 ( .A(n3780), .B(n3781), .Z(n3778) );
  XNOR U2747 ( .A(n3775), .B(n3782), .Z(SUM[369]) );
  NANDN U2748 ( .A(n3773), .B(n3776), .Z(n3782) );
  NANDN U2749 ( .A(n3783), .B(n3784), .Z(n3775) );
  NAND U2750 ( .A(n3763), .B(n3785), .Z(n3784) );
  XNOR U2751 ( .A(n3763), .B(n3786), .Z(SUM[368]) );
  NANDN U2752 ( .A(n3783), .B(n3785), .Z(n3786) );
  NANDN U2753 ( .A(n3787), .B(n3788), .Z(n3763) );
  NANDN U2754 ( .A(n3789), .B(n3790), .Z(n3788) );
  XOR U2755 ( .A(n3791), .B(n3792), .Z(SUM[367]) );
  NANDN U2756 ( .A(n3793), .B(n3794), .Z(n3792) );
  ANDN U2757 ( .B(n3795), .A(n3796), .Z(n3791) );
  NAND U2758 ( .A(n3797), .B(n3798), .Z(n3795) );
  XNOR U2759 ( .A(n3797), .B(n3799), .Z(SUM[366]) );
  NANDN U2760 ( .A(n3796), .B(n3798), .Z(n3799) );
  NANDN U2761 ( .A(n3800), .B(n3801), .Z(n3797) );
  NAND U2762 ( .A(n3802), .B(n3803), .Z(n3801) );
  XNOR U2763 ( .A(n3802), .B(n3804), .Z(SUM[365]) );
  NANDN U2764 ( .A(n3800), .B(n3803), .Z(n3804) );
  NANDN U2765 ( .A(n3805), .B(n3806), .Z(n3802) );
  NAND U2766 ( .A(n3807), .B(n3808), .Z(n3806) );
  XNOR U2767 ( .A(n3807), .B(n3809), .Z(SUM[364]) );
  NANDN U2768 ( .A(n3805), .B(n3808), .Z(n3809) );
  NANDN U2769 ( .A(n3810), .B(n3811), .Z(n3807) );
  NANDN U2770 ( .A(n3812), .B(n3813), .Z(n3811) );
  XOR U2771 ( .A(n3814), .B(n3815), .Z(SUM[363]) );
  NANDN U2772 ( .A(n3816), .B(n3817), .Z(n3815) );
  ANDN U2773 ( .B(n3818), .A(n3819), .Z(n3814) );
  NAND U2774 ( .A(n3820), .B(n3821), .Z(n3818) );
  XNOR U2775 ( .A(n3820), .B(n3822), .Z(SUM[362]) );
  NANDN U2776 ( .A(n3819), .B(n3821), .Z(n3822) );
  NANDN U2777 ( .A(n3823), .B(n3824), .Z(n3820) );
  NAND U2778 ( .A(n3825), .B(n3826), .Z(n3824) );
  XNOR U2779 ( .A(n3825), .B(n3827), .Z(SUM[361]) );
  NANDN U2780 ( .A(n3823), .B(n3826), .Z(n3827) );
  NANDN U2781 ( .A(n3828), .B(n3829), .Z(n3825) );
  NAND U2782 ( .A(n3813), .B(n3830), .Z(n3829) );
  XNOR U2783 ( .A(n3813), .B(n3831), .Z(SUM[360]) );
  NANDN U2784 ( .A(n3828), .B(n3830), .Z(n3831) );
  NANDN U2785 ( .A(n3832), .B(n3833), .Z(n3813) );
  OR U2786 ( .A(n3834), .B(n3835), .Z(n3833) );
  XOR U2787 ( .A(n3836), .B(n3837), .Z(SUM[35]) );
  NANDN U2788 ( .A(n3838), .B(n3839), .Z(n3837) );
  ANDN U2789 ( .B(n3840), .A(n3841), .Z(n3836) );
  NANDN U2790 ( .A(n3842), .B(n3843), .Z(n3840) );
  XOR U2791 ( .A(n3844), .B(n3845), .Z(SUM[359]) );
  NANDN U2792 ( .A(n3846), .B(n3847), .Z(n3845) );
  ANDN U2793 ( .B(n3848), .A(n3849), .Z(n3844) );
  NAND U2794 ( .A(n3850), .B(n3851), .Z(n3848) );
  XNOR U2795 ( .A(n3850), .B(n3852), .Z(SUM[358]) );
  NANDN U2796 ( .A(n3849), .B(n3851), .Z(n3852) );
  NANDN U2797 ( .A(n3853), .B(n3854), .Z(n3850) );
  NAND U2798 ( .A(n3855), .B(n3856), .Z(n3854) );
  XNOR U2799 ( .A(n3855), .B(n3857), .Z(SUM[357]) );
  NANDN U2800 ( .A(n3853), .B(n3856), .Z(n3857) );
  NANDN U2801 ( .A(n3858), .B(n3859), .Z(n3855) );
  NANDN U2802 ( .A(n3835), .B(n3860), .Z(n3859) );
  XOR U2803 ( .A(n3835), .B(n3861), .Z(SUM[356]) );
  NANDN U2804 ( .A(n3858), .B(n3860), .Z(n3861) );
  ANDN U2805 ( .B(n3862), .A(n3863), .Z(n3835) );
  NANDN U2806 ( .A(n3864), .B(n3790), .Z(n3862) );
  XOR U2807 ( .A(n3865), .B(n3866), .Z(SUM[355]) );
  NANDN U2808 ( .A(n3867), .B(n3868), .Z(n3866) );
  ANDN U2809 ( .B(n3869), .A(n3870), .Z(n3865) );
  NAND U2810 ( .A(n3871), .B(n3872), .Z(n3869) );
  XNOR U2811 ( .A(n3871), .B(n3873), .Z(SUM[354]) );
  NANDN U2812 ( .A(n3870), .B(n3872), .Z(n3873) );
  NANDN U2813 ( .A(n3874), .B(n3875), .Z(n3871) );
  NAND U2814 ( .A(n3876), .B(n3877), .Z(n3875) );
  XNOR U2815 ( .A(n3876), .B(n3878), .Z(SUM[353]) );
  NANDN U2816 ( .A(n3874), .B(n3877), .Z(n3878) );
  NANDN U2817 ( .A(n3879), .B(n3880), .Z(n3876) );
  NAND U2818 ( .A(n3790), .B(n3881), .Z(n3880) );
  XNOR U2819 ( .A(n3790), .B(n3882), .Z(SUM[352]) );
  NANDN U2820 ( .A(n3879), .B(n3881), .Z(n3882) );
  NANDN U2821 ( .A(n3883), .B(n3884), .Z(n3790) );
  OR U2822 ( .A(n3885), .B(n3886), .Z(n3884) );
  XOR U2823 ( .A(n3887), .B(n3888), .Z(SUM[351]) );
  NANDN U2824 ( .A(n3889), .B(n3890), .Z(n3888) );
  ANDN U2825 ( .B(n3891), .A(n3892), .Z(n3887) );
  NAND U2826 ( .A(n3893), .B(n3894), .Z(n3891) );
  XNOR U2827 ( .A(n3893), .B(n3895), .Z(SUM[350]) );
  NANDN U2828 ( .A(n3892), .B(n3894), .Z(n3895) );
  NANDN U2829 ( .A(n3896), .B(n3897), .Z(n3893) );
  NAND U2830 ( .A(n3898), .B(n3899), .Z(n3897) );
  XNOR U2831 ( .A(n3843), .B(n3900), .Z(SUM[34]) );
  OR U2832 ( .A(n3842), .B(n3841), .Z(n3900) );
  NANDN U2833 ( .A(n3901), .B(n3902), .Z(n3843) );
  NAND U2834 ( .A(n3903), .B(n3904), .Z(n3902) );
  XNOR U2835 ( .A(n3898), .B(n3905), .Z(SUM[349]) );
  NANDN U2836 ( .A(n3896), .B(n3899), .Z(n3905) );
  NANDN U2837 ( .A(n3906), .B(n3907), .Z(n3898) );
  NAND U2838 ( .A(n3908), .B(n3909), .Z(n3907) );
  XNOR U2839 ( .A(n3908), .B(n3910), .Z(SUM[348]) );
  NANDN U2840 ( .A(n3906), .B(n3909), .Z(n3910) );
  NANDN U2841 ( .A(n3911), .B(n3912), .Z(n3908) );
  NANDN U2842 ( .A(n3913), .B(n3914), .Z(n3912) );
  XOR U2843 ( .A(n3915), .B(n3916), .Z(SUM[347]) );
  NANDN U2844 ( .A(n3917), .B(n3918), .Z(n3916) );
  ANDN U2845 ( .B(n3919), .A(n3920), .Z(n3915) );
  NAND U2846 ( .A(n3921), .B(n3922), .Z(n3919) );
  XNOR U2847 ( .A(n3921), .B(n3923), .Z(SUM[346]) );
  NANDN U2848 ( .A(n3920), .B(n3922), .Z(n3923) );
  NANDN U2849 ( .A(n3924), .B(n3925), .Z(n3921) );
  NAND U2850 ( .A(n3926), .B(n3927), .Z(n3925) );
  XNOR U2851 ( .A(n3926), .B(n3928), .Z(SUM[345]) );
  NANDN U2852 ( .A(n3924), .B(n3927), .Z(n3928) );
  NANDN U2853 ( .A(n3929), .B(n3930), .Z(n3926) );
  NAND U2854 ( .A(n3914), .B(n3931), .Z(n3930) );
  XNOR U2855 ( .A(n3914), .B(n3932), .Z(SUM[344]) );
  NANDN U2856 ( .A(n3929), .B(n3931), .Z(n3932) );
  NANDN U2857 ( .A(n3933), .B(n3934), .Z(n3914) );
  OR U2858 ( .A(n3935), .B(n3936), .Z(n3934) );
  XOR U2859 ( .A(n3937), .B(n3938), .Z(SUM[343]) );
  NANDN U2860 ( .A(n3939), .B(n3940), .Z(n3938) );
  ANDN U2861 ( .B(n3941), .A(n3942), .Z(n3937) );
  NAND U2862 ( .A(n3943), .B(n3944), .Z(n3941) );
  XNOR U2863 ( .A(n3943), .B(n3945), .Z(SUM[342]) );
  NANDN U2864 ( .A(n3942), .B(n3944), .Z(n3945) );
  NANDN U2865 ( .A(n3946), .B(n3947), .Z(n3943) );
  NAND U2866 ( .A(n3948), .B(n3949), .Z(n3947) );
  XNOR U2867 ( .A(n3948), .B(n3950), .Z(SUM[341]) );
  NANDN U2868 ( .A(n3946), .B(n3949), .Z(n3950) );
  NANDN U2869 ( .A(n3951), .B(n3952), .Z(n3948) );
  NANDN U2870 ( .A(n3936), .B(n3953), .Z(n3952) );
  XOR U2871 ( .A(n3936), .B(n3954), .Z(SUM[340]) );
  NANDN U2872 ( .A(n3951), .B(n3953), .Z(n3954) );
  ANDN U2873 ( .B(n3955), .A(n3956), .Z(n3936) );
  OR U2874 ( .A(n3957), .B(n3886), .Z(n3955) );
  XNOR U2875 ( .A(n3903), .B(n3958), .Z(SUM[33]) );
  NANDN U2876 ( .A(n3901), .B(n3904), .Z(n3958) );
  NANDN U2877 ( .A(n3959), .B(n3960), .Z(n3903) );
  NANDN U2878 ( .A(n3781), .B(n3961), .Z(n3960) );
  XOR U2879 ( .A(n3962), .B(n3963), .Z(SUM[339]) );
  NANDN U2880 ( .A(n3964), .B(n3965), .Z(n3963) );
  ANDN U2881 ( .B(n3966), .A(n3967), .Z(n3962) );
  NAND U2882 ( .A(n3968), .B(n3969), .Z(n3966) );
  XNOR U2883 ( .A(n3968), .B(n3970), .Z(SUM[338]) );
  NANDN U2884 ( .A(n3967), .B(n3969), .Z(n3970) );
  NANDN U2885 ( .A(n3971), .B(n3972), .Z(n3968) );
  NAND U2886 ( .A(n3973), .B(n3974), .Z(n3972) );
  XNOR U2887 ( .A(n3973), .B(n3975), .Z(SUM[337]) );
  NANDN U2888 ( .A(n3971), .B(n3974), .Z(n3975) );
  NANDN U2889 ( .A(n3976), .B(n3977), .Z(n3973) );
  NANDN U2890 ( .A(n3886), .B(n3978), .Z(n3977) );
  XOR U2891 ( .A(n3886), .B(n3979), .Z(SUM[336]) );
  NANDN U2892 ( .A(n3976), .B(n3978), .Z(n3979) );
  ANDN U2893 ( .B(n3980), .A(n3981), .Z(n3886) );
  OR U2894 ( .A(n3982), .B(n3692), .Z(n3980) );
  XOR U2895 ( .A(n3983), .B(n3984), .Z(SUM[335]) );
  NANDN U2896 ( .A(n3985), .B(n3986), .Z(n3984) );
  ANDN U2897 ( .B(n3987), .A(n3988), .Z(n3983) );
  NAND U2898 ( .A(n3989), .B(n3990), .Z(n3987) );
  XNOR U2899 ( .A(n3989), .B(n3991), .Z(SUM[334]) );
  NANDN U2900 ( .A(n3988), .B(n3990), .Z(n3991) );
  NANDN U2901 ( .A(n3992), .B(n3993), .Z(n3989) );
  NAND U2902 ( .A(n3994), .B(n3995), .Z(n3993) );
  XNOR U2903 ( .A(n3994), .B(n3996), .Z(SUM[333]) );
  NANDN U2904 ( .A(n3992), .B(n3995), .Z(n3996) );
  NANDN U2905 ( .A(n3997), .B(n3998), .Z(n3994) );
  NAND U2906 ( .A(n3999), .B(n4000), .Z(n3998) );
  XNOR U2907 ( .A(n3999), .B(n4001), .Z(SUM[332]) );
  NANDN U2908 ( .A(n3997), .B(n4000), .Z(n4001) );
  NANDN U2909 ( .A(n4002), .B(n4003), .Z(n3999) );
  NANDN U2910 ( .A(n4004), .B(n4005), .Z(n4003) );
  XOR U2911 ( .A(n4006), .B(n4007), .Z(SUM[331]) );
  NANDN U2912 ( .A(n4008), .B(n4009), .Z(n4007) );
  ANDN U2913 ( .B(n4010), .A(n4011), .Z(n4006) );
  NAND U2914 ( .A(n4012), .B(n4013), .Z(n4010) );
  XNOR U2915 ( .A(n4012), .B(n4014), .Z(SUM[330]) );
  NANDN U2916 ( .A(n4011), .B(n4013), .Z(n4014) );
  NANDN U2917 ( .A(n4015), .B(n4016), .Z(n4012) );
  NAND U2918 ( .A(n4017), .B(n4018), .Z(n4016) );
  XOR U2919 ( .A(n3781), .B(n4019), .Z(SUM[32]) );
  NANDN U2920 ( .A(n3959), .B(n3961), .Z(n4019) );
  XNOR U2921 ( .A(n4017), .B(n4020), .Z(SUM[329]) );
  NANDN U2922 ( .A(n4015), .B(n4018), .Z(n4020) );
  NANDN U2923 ( .A(n4021), .B(n4022), .Z(n4017) );
  NAND U2924 ( .A(n4005), .B(n4023), .Z(n4022) );
  XNOR U2925 ( .A(n4005), .B(n4024), .Z(SUM[328]) );
  NANDN U2926 ( .A(n4021), .B(n4023), .Z(n4024) );
  NANDN U2927 ( .A(n4025), .B(n4026), .Z(n4005) );
  OR U2928 ( .A(n4027), .B(n4028), .Z(n4026) );
  XOR U2929 ( .A(n4029), .B(n4030), .Z(SUM[327]) );
  NANDN U2930 ( .A(n4031), .B(n4032), .Z(n4030) );
  ANDN U2931 ( .B(n4033), .A(n4034), .Z(n4029) );
  NAND U2932 ( .A(n4035), .B(n4036), .Z(n4033) );
  XNOR U2933 ( .A(n4035), .B(n4037), .Z(SUM[326]) );
  NANDN U2934 ( .A(n4034), .B(n4036), .Z(n4037) );
  NANDN U2935 ( .A(n4038), .B(n4039), .Z(n4035) );
  NAND U2936 ( .A(n4040), .B(n4041), .Z(n4039) );
  XNOR U2937 ( .A(n4040), .B(n4042), .Z(SUM[325]) );
  NANDN U2938 ( .A(n4038), .B(n4041), .Z(n4042) );
  NANDN U2939 ( .A(n4043), .B(n4044), .Z(n4040) );
  NANDN U2940 ( .A(n4028), .B(n4045), .Z(n4044) );
  XOR U2941 ( .A(n4028), .B(n4046), .Z(SUM[324]) );
  NANDN U2942 ( .A(n4043), .B(n4045), .Z(n4046) );
  ANDN U2943 ( .B(n4047), .A(n4048), .Z(n4028) );
  OR U2944 ( .A(n4049), .B(n3692), .Z(n4047) );
  XOR U2945 ( .A(n4050), .B(n4051), .Z(SUM[323]) );
  NANDN U2946 ( .A(n4052), .B(n4053), .Z(n4051) );
  ANDN U2947 ( .B(n4054), .A(n4055), .Z(n4050) );
  NAND U2948 ( .A(n4056), .B(n4057), .Z(n4054) );
  XNOR U2949 ( .A(n4056), .B(n4058), .Z(SUM[322]) );
  NANDN U2950 ( .A(n4055), .B(n4057), .Z(n4058) );
  NANDN U2951 ( .A(n4059), .B(n4060), .Z(n4056) );
  NAND U2952 ( .A(n4061), .B(n4062), .Z(n4060) );
  XNOR U2953 ( .A(n4061), .B(n4063), .Z(SUM[321]) );
  NANDN U2954 ( .A(n4059), .B(n4062), .Z(n4063) );
  NANDN U2955 ( .A(n4064), .B(n4065), .Z(n4061) );
  NANDN U2956 ( .A(n3692), .B(n4066), .Z(n4065) );
  XOR U2957 ( .A(n3692), .B(n4067), .Z(SUM[320]) );
  NANDN U2958 ( .A(n4064), .B(n4066), .Z(n4067) );
  NOR U2959 ( .A(n4068), .B(n4069), .Z(n3692) );
  XOR U2960 ( .A(n4070), .B(n4071), .Z(SUM[31]) );
  OR U2961 ( .A(n4072), .B(n4073), .Z(n4071) );
  ANDN U2962 ( .B(n4074), .A(n4075), .Z(n4070) );
  NANDN U2963 ( .A(n4076), .B(n4077), .Z(n4074) );
  XOR U2964 ( .A(n4078), .B(n4079), .Z(SUM[319]) );
  NANDN U2965 ( .A(n4080), .B(n4081), .Z(n4079) );
  ANDN U2966 ( .B(n4082), .A(n4083), .Z(n4078) );
  NAND U2967 ( .A(n4084), .B(n4085), .Z(n4082) );
  XNOR U2968 ( .A(n4084), .B(n4086), .Z(SUM[318]) );
  NANDN U2969 ( .A(n4083), .B(n4085), .Z(n4086) );
  NANDN U2970 ( .A(n4087), .B(n4088), .Z(n4084) );
  NAND U2971 ( .A(n4089), .B(n4090), .Z(n4088) );
  XNOR U2972 ( .A(n4089), .B(n4091), .Z(SUM[317]) );
  NANDN U2973 ( .A(n4087), .B(n4090), .Z(n4091) );
  NANDN U2974 ( .A(n4092), .B(n4093), .Z(n4089) );
  NAND U2975 ( .A(n4094), .B(n4095), .Z(n4093) );
  XNOR U2976 ( .A(n4094), .B(n4096), .Z(SUM[316]) );
  NANDN U2977 ( .A(n4092), .B(n4095), .Z(n4096) );
  NANDN U2978 ( .A(n4097), .B(n4098), .Z(n4094) );
  NANDN U2979 ( .A(n4099), .B(n4100), .Z(n4098) );
  XOR U2980 ( .A(n4101), .B(n4102), .Z(SUM[315]) );
  NANDN U2981 ( .A(n4103), .B(n4104), .Z(n4102) );
  ANDN U2982 ( .B(n4105), .A(n4106), .Z(n4101) );
  NAND U2983 ( .A(n4107), .B(n4108), .Z(n4105) );
  XNOR U2984 ( .A(n4107), .B(n4109), .Z(SUM[314]) );
  NANDN U2985 ( .A(n4106), .B(n4108), .Z(n4109) );
  NANDN U2986 ( .A(n4110), .B(n4111), .Z(n4107) );
  NAND U2987 ( .A(n4112), .B(n4113), .Z(n4111) );
  XNOR U2988 ( .A(n4112), .B(n4114), .Z(SUM[313]) );
  NANDN U2989 ( .A(n4110), .B(n4113), .Z(n4114) );
  NANDN U2990 ( .A(n4115), .B(n4116), .Z(n4112) );
  NAND U2991 ( .A(n4100), .B(n4117), .Z(n4116) );
  XNOR U2992 ( .A(n4100), .B(n4118), .Z(SUM[312]) );
  NANDN U2993 ( .A(n4115), .B(n4117), .Z(n4118) );
  NANDN U2994 ( .A(n4119), .B(n4120), .Z(n4100) );
  OR U2995 ( .A(n4121), .B(n4122), .Z(n4120) );
  XOR U2996 ( .A(n4123), .B(n4124), .Z(SUM[311]) );
  NANDN U2997 ( .A(n4125), .B(n4126), .Z(n4124) );
  ANDN U2998 ( .B(n4127), .A(n4128), .Z(n4123) );
  NAND U2999 ( .A(n4129), .B(n4130), .Z(n4127) );
  XNOR U3000 ( .A(n4129), .B(n4131), .Z(SUM[310]) );
  NANDN U3001 ( .A(n4128), .B(n4130), .Z(n4131) );
  NANDN U3002 ( .A(n4132), .B(n4133), .Z(n4129) );
  NAND U3003 ( .A(n4134), .B(n4135), .Z(n4133) );
  XNOR U3004 ( .A(n4077), .B(n4136), .Z(SUM[30]) );
  OR U3005 ( .A(n4076), .B(n4075), .Z(n4136) );
  NANDN U3006 ( .A(n4137), .B(n4138), .Z(n4077) );
  NANDN U3007 ( .A(n4139), .B(n4140), .Z(n4138) );
  XNOR U3008 ( .A(n4134), .B(n4141), .Z(SUM[309]) );
  NANDN U3009 ( .A(n4132), .B(n4135), .Z(n4141) );
  NANDN U3010 ( .A(n4142), .B(n4143), .Z(n4134) );
  NANDN U3011 ( .A(n4122), .B(n4144), .Z(n4143) );
  XOR U3012 ( .A(n4122), .B(n4145), .Z(SUM[308]) );
  NANDN U3013 ( .A(n4142), .B(n4144), .Z(n4145) );
  ANDN U3014 ( .B(n4146), .A(n4147), .Z(n4122) );
  NANDN U3015 ( .A(n4148), .B(n4149), .Z(n4146) );
  XOR U3016 ( .A(n4150), .B(n4151), .Z(SUM[307]) );
  NANDN U3017 ( .A(n4152), .B(n4153), .Z(n4151) );
  ANDN U3018 ( .B(n4154), .A(n4155), .Z(n4150) );
  NAND U3019 ( .A(n4156), .B(n4157), .Z(n4154) );
  XNOR U3020 ( .A(n4156), .B(n4158), .Z(SUM[306]) );
  NANDN U3021 ( .A(n4155), .B(n4157), .Z(n4158) );
  NANDN U3022 ( .A(n4159), .B(n4160), .Z(n4156) );
  NAND U3023 ( .A(n4161), .B(n4162), .Z(n4160) );
  XNOR U3024 ( .A(n4161), .B(n4163), .Z(SUM[305]) );
  NANDN U3025 ( .A(n4159), .B(n4162), .Z(n4163) );
  NANDN U3026 ( .A(n4164), .B(n4165), .Z(n4161) );
  NAND U3027 ( .A(n4149), .B(n4166), .Z(n4165) );
  XNOR U3028 ( .A(n4149), .B(n4167), .Z(SUM[304]) );
  NANDN U3029 ( .A(n4164), .B(n4166), .Z(n4167) );
  NANDN U3030 ( .A(n4168), .B(n4169), .Z(n4149) );
  NANDN U3031 ( .A(n4170), .B(n4171), .Z(n4169) );
  XOR U3032 ( .A(n4172), .B(n4173), .Z(SUM[303]) );
  NANDN U3033 ( .A(n4174), .B(n4175), .Z(n4173) );
  ANDN U3034 ( .B(n4176), .A(n4177), .Z(n4172) );
  NAND U3035 ( .A(n4178), .B(n4179), .Z(n4176) );
  XNOR U3036 ( .A(n4178), .B(n4180), .Z(SUM[302]) );
  NANDN U3037 ( .A(n4177), .B(n4179), .Z(n4180) );
  NANDN U3038 ( .A(n4181), .B(n4182), .Z(n4178) );
  NAND U3039 ( .A(n4183), .B(n4184), .Z(n4182) );
  XNOR U3040 ( .A(n4183), .B(n4185), .Z(SUM[301]) );
  NANDN U3041 ( .A(n4181), .B(n4184), .Z(n4185) );
  NANDN U3042 ( .A(n4186), .B(n4187), .Z(n4183) );
  NAND U3043 ( .A(n4188), .B(n4189), .Z(n4187) );
  XNOR U3044 ( .A(n4188), .B(n4190), .Z(SUM[300]) );
  NANDN U3045 ( .A(n4186), .B(n4189), .Z(n4190) );
  NANDN U3046 ( .A(n4191), .B(n4192), .Z(n4188) );
  NANDN U3047 ( .A(n4193), .B(n4194), .Z(n4192) );
  XNOR U3048 ( .A(n4140), .B(n4195), .Z(SUM[29]) );
  OR U3049 ( .A(n4139), .B(n4137), .Z(n4195) );
  NANDN U3050 ( .A(n4196), .B(n4197), .Z(n4140) );
  NAND U3051 ( .A(n4198), .B(n4199), .Z(n4197) );
  XOR U3052 ( .A(n4200), .B(n4201), .Z(SUM[299]) );
  NANDN U3053 ( .A(n4202), .B(n4203), .Z(n4201) );
  ANDN U3054 ( .B(n4204), .A(n4205), .Z(n4200) );
  NAND U3055 ( .A(n4206), .B(n4207), .Z(n4204) );
  XNOR U3056 ( .A(n4206), .B(n4208), .Z(SUM[298]) );
  NANDN U3057 ( .A(n4205), .B(n4207), .Z(n4208) );
  NANDN U3058 ( .A(n4209), .B(n4210), .Z(n4206) );
  NAND U3059 ( .A(n4211), .B(n4212), .Z(n4210) );
  XNOR U3060 ( .A(n4211), .B(n4213), .Z(SUM[297]) );
  NANDN U3061 ( .A(n4209), .B(n4212), .Z(n4213) );
  NANDN U3062 ( .A(n4214), .B(n4215), .Z(n4211) );
  NAND U3063 ( .A(n4194), .B(n4216), .Z(n4215) );
  XNOR U3064 ( .A(n4194), .B(n4217), .Z(SUM[296]) );
  NANDN U3065 ( .A(n4214), .B(n4216), .Z(n4217) );
  NANDN U3066 ( .A(n4218), .B(n4219), .Z(n4194) );
  OR U3067 ( .A(n4220), .B(n4221), .Z(n4219) );
  XOR U3068 ( .A(n4222), .B(n4223), .Z(SUM[295]) );
  NANDN U3069 ( .A(n4224), .B(n4225), .Z(n4223) );
  ANDN U3070 ( .B(n4226), .A(n4227), .Z(n4222) );
  NAND U3071 ( .A(n4228), .B(n4229), .Z(n4226) );
  XNOR U3072 ( .A(n4228), .B(n4230), .Z(SUM[294]) );
  NANDN U3073 ( .A(n4227), .B(n4229), .Z(n4230) );
  NANDN U3074 ( .A(n4231), .B(n4232), .Z(n4228) );
  NAND U3075 ( .A(n4233), .B(n4234), .Z(n4232) );
  XNOR U3076 ( .A(n4233), .B(n4235), .Z(SUM[293]) );
  NANDN U3077 ( .A(n4231), .B(n4234), .Z(n4235) );
  NANDN U3078 ( .A(n4236), .B(n4237), .Z(n4233) );
  NANDN U3079 ( .A(n4221), .B(n4238), .Z(n4237) );
  XOR U3080 ( .A(n4221), .B(n4239), .Z(SUM[292]) );
  NANDN U3081 ( .A(n4236), .B(n4238), .Z(n4239) );
  ANDN U3082 ( .B(n4240), .A(n4241), .Z(n4221) );
  NANDN U3083 ( .A(n4242), .B(n4171), .Z(n4240) );
  XOR U3084 ( .A(n4243), .B(n4244), .Z(SUM[291]) );
  NANDN U3085 ( .A(n4245), .B(n4246), .Z(n4244) );
  ANDN U3086 ( .B(n4247), .A(n4248), .Z(n4243) );
  NAND U3087 ( .A(n4249), .B(n4250), .Z(n4247) );
  XNOR U3088 ( .A(n4249), .B(n4251), .Z(SUM[290]) );
  NANDN U3089 ( .A(n4248), .B(n4250), .Z(n4251) );
  NANDN U3090 ( .A(n4252), .B(n4253), .Z(n4249) );
  NAND U3091 ( .A(n4254), .B(n4255), .Z(n4253) );
  XNOR U3092 ( .A(n4198), .B(n4256), .Z(SUM[28]) );
  NANDN U3093 ( .A(n4196), .B(n4199), .Z(n4256) );
  NANDN U3094 ( .A(n4257), .B(n4258), .Z(n4198) );
  NANDN U3095 ( .A(n4259), .B(n4260), .Z(n4258) );
  XNOR U3096 ( .A(n4254), .B(n4261), .Z(SUM[289]) );
  NANDN U3097 ( .A(n4252), .B(n4255), .Z(n4261) );
  NANDN U3098 ( .A(n4262), .B(n4263), .Z(n4254) );
  NAND U3099 ( .A(n4171), .B(n4264), .Z(n4263) );
  XNOR U3100 ( .A(n4171), .B(n4265), .Z(SUM[288]) );
  NANDN U3101 ( .A(n4262), .B(n4264), .Z(n4265) );
  NANDN U3102 ( .A(n4266), .B(n4267), .Z(n4171) );
  OR U3103 ( .A(n4268), .B(n4269), .Z(n4267) );
  XOR U3104 ( .A(n4270), .B(n4271), .Z(SUM[287]) );
  NANDN U3105 ( .A(n4272), .B(n4273), .Z(n4271) );
  ANDN U3106 ( .B(n4274), .A(n4275), .Z(n4270) );
  NAND U3107 ( .A(n4276), .B(n4277), .Z(n4274) );
  XNOR U3108 ( .A(n4276), .B(n4278), .Z(SUM[286]) );
  NANDN U3109 ( .A(n4275), .B(n4277), .Z(n4278) );
  NANDN U3110 ( .A(n4279), .B(n4280), .Z(n4276) );
  NAND U3111 ( .A(n4281), .B(n4282), .Z(n4280) );
  XNOR U3112 ( .A(n4281), .B(n4283), .Z(SUM[285]) );
  NANDN U3113 ( .A(n4279), .B(n4282), .Z(n4283) );
  NANDN U3114 ( .A(n4284), .B(n4285), .Z(n4281) );
  NAND U3115 ( .A(n4286), .B(n4287), .Z(n4285) );
  XNOR U3116 ( .A(n4286), .B(n4288), .Z(SUM[284]) );
  NANDN U3117 ( .A(n4284), .B(n4287), .Z(n4288) );
  NANDN U3118 ( .A(n4289), .B(n4290), .Z(n4286) );
  NANDN U3119 ( .A(n4291), .B(n4292), .Z(n4290) );
  XOR U3120 ( .A(n4293), .B(n4294), .Z(SUM[283]) );
  NANDN U3121 ( .A(n4295), .B(n4296), .Z(n4294) );
  ANDN U3122 ( .B(n4297), .A(n4298), .Z(n4293) );
  NAND U3123 ( .A(n4299), .B(n4300), .Z(n4297) );
  XNOR U3124 ( .A(n4299), .B(n4301), .Z(SUM[282]) );
  NANDN U3125 ( .A(n4298), .B(n4300), .Z(n4301) );
  NANDN U3126 ( .A(n4302), .B(n4303), .Z(n4299) );
  NAND U3127 ( .A(n4304), .B(n4305), .Z(n4303) );
  XNOR U3128 ( .A(n4304), .B(n4306), .Z(SUM[281]) );
  NANDN U3129 ( .A(n4302), .B(n4305), .Z(n4306) );
  NANDN U3130 ( .A(n4307), .B(n4308), .Z(n4304) );
  NAND U3131 ( .A(n4292), .B(n4309), .Z(n4308) );
  XNOR U3132 ( .A(n4292), .B(n4310), .Z(SUM[280]) );
  NANDN U3133 ( .A(n4307), .B(n4309), .Z(n4310) );
  NANDN U3134 ( .A(n4311), .B(n4312), .Z(n4292) );
  OR U3135 ( .A(n4313), .B(n4314), .Z(n4312) );
  XOR U3136 ( .A(n4315), .B(n4316), .Z(SUM[27]) );
  NANDN U3137 ( .A(n4317), .B(n4318), .Z(n4316) );
  ANDN U3138 ( .B(n4319), .A(n4320), .Z(n4315) );
  NAND U3139 ( .A(n4321), .B(n4322), .Z(n4319) );
  XOR U3140 ( .A(n4323), .B(n4324), .Z(SUM[279]) );
  NANDN U3141 ( .A(n4325), .B(n4326), .Z(n4324) );
  ANDN U3142 ( .B(n4327), .A(n4328), .Z(n4323) );
  NAND U3143 ( .A(n4329), .B(n4330), .Z(n4327) );
  XNOR U3144 ( .A(n4329), .B(n4331), .Z(SUM[278]) );
  NANDN U3145 ( .A(n4328), .B(n4330), .Z(n4331) );
  NANDN U3146 ( .A(n4332), .B(n4333), .Z(n4329) );
  NAND U3147 ( .A(n4334), .B(n4335), .Z(n4333) );
  XNOR U3148 ( .A(n4334), .B(n4336), .Z(SUM[277]) );
  NANDN U3149 ( .A(n4332), .B(n4335), .Z(n4336) );
  NANDN U3150 ( .A(n4337), .B(n4338), .Z(n4334) );
  NANDN U3151 ( .A(n4314), .B(n4339), .Z(n4338) );
  XOR U3152 ( .A(n4314), .B(n4340), .Z(SUM[276]) );
  NANDN U3153 ( .A(n4337), .B(n4339), .Z(n4340) );
  ANDN U3154 ( .B(n4341), .A(n4342), .Z(n4314) );
  OR U3155 ( .A(n4343), .B(n4269), .Z(n4341) );
  XOR U3156 ( .A(n4344), .B(n4345), .Z(SUM[275]) );
  NANDN U3157 ( .A(n4346), .B(n4347), .Z(n4345) );
  ANDN U3158 ( .B(n4348), .A(n4349), .Z(n4344) );
  NAND U3159 ( .A(n4350), .B(n4351), .Z(n4348) );
  XNOR U3160 ( .A(n4350), .B(n4352), .Z(SUM[274]) );
  NANDN U3161 ( .A(n4349), .B(n4351), .Z(n4352) );
  NANDN U3162 ( .A(n4353), .B(n4354), .Z(n4350) );
  NAND U3163 ( .A(n4355), .B(n4356), .Z(n4354) );
  XNOR U3164 ( .A(n4355), .B(n4357), .Z(SUM[273]) );
  NANDN U3165 ( .A(n4353), .B(n4356), .Z(n4357) );
  NANDN U3166 ( .A(n4358), .B(n4359), .Z(n4355) );
  NANDN U3167 ( .A(n4269), .B(n4360), .Z(n4359) );
  XOR U3168 ( .A(n4269), .B(n4361), .Z(SUM[272]) );
  NANDN U3169 ( .A(n4358), .B(n4360), .Z(n4361) );
  ANDN U3170 ( .B(n4362), .A(n4363), .Z(n4269) );
  OR U3171 ( .A(n4364), .B(n4365), .Z(n4362) );
  XOR U3172 ( .A(n4366), .B(n4367), .Z(SUM[271]) );
  NANDN U3173 ( .A(n4368), .B(n4369), .Z(n4367) );
  ANDN U3174 ( .B(n4370), .A(n4371), .Z(n4366) );
  NAND U3175 ( .A(n4372), .B(n4373), .Z(n4370) );
  XNOR U3176 ( .A(n4372), .B(n4374), .Z(SUM[270]) );
  NANDN U3177 ( .A(n4371), .B(n4373), .Z(n4374) );
  NANDN U3178 ( .A(n4375), .B(n4376), .Z(n4372) );
  NAND U3179 ( .A(n4377), .B(n4378), .Z(n4376) );
  XNOR U3180 ( .A(n4321), .B(n4379), .Z(SUM[26]) );
  NANDN U3181 ( .A(n4320), .B(n4322), .Z(n4379) );
  NANDN U3182 ( .A(n4380), .B(n4381), .Z(n4321) );
  NAND U3183 ( .A(n4382), .B(n4383), .Z(n4381) );
  XNOR U3184 ( .A(n4377), .B(n4384), .Z(SUM[269]) );
  NANDN U3185 ( .A(n4375), .B(n4378), .Z(n4384) );
  NANDN U3186 ( .A(n4385), .B(n4386), .Z(n4377) );
  NAND U3187 ( .A(n4387), .B(n4388), .Z(n4386) );
  XNOR U3188 ( .A(n4387), .B(n4389), .Z(SUM[268]) );
  NANDN U3189 ( .A(n4385), .B(n4388), .Z(n4389) );
  NANDN U3190 ( .A(n4390), .B(n4391), .Z(n4387) );
  NANDN U3191 ( .A(n4392), .B(n4393), .Z(n4391) );
  XOR U3192 ( .A(n4394), .B(n4395), .Z(SUM[267]) );
  NANDN U3193 ( .A(n4396), .B(n4397), .Z(n4395) );
  ANDN U3194 ( .B(n4398), .A(n4399), .Z(n4394) );
  NAND U3195 ( .A(n4400), .B(n4401), .Z(n4398) );
  XNOR U3196 ( .A(n4400), .B(n4402), .Z(SUM[266]) );
  NANDN U3197 ( .A(n4399), .B(n4401), .Z(n4402) );
  NANDN U3198 ( .A(n4403), .B(n4404), .Z(n4400) );
  NAND U3199 ( .A(n4405), .B(n4406), .Z(n4404) );
  XNOR U3200 ( .A(n4405), .B(n4407), .Z(SUM[265]) );
  NANDN U3201 ( .A(n4403), .B(n4406), .Z(n4407) );
  NANDN U3202 ( .A(n4408), .B(n4409), .Z(n4405) );
  NAND U3203 ( .A(n4393), .B(n4410), .Z(n4409) );
  XNOR U3204 ( .A(n4393), .B(n4411), .Z(SUM[264]) );
  NANDN U3205 ( .A(n4408), .B(n4410), .Z(n4411) );
  NANDN U3206 ( .A(n4412), .B(n4413), .Z(n4393) );
  OR U3207 ( .A(n4414), .B(n4415), .Z(n4413) );
  XOR U3208 ( .A(n4416), .B(n4417), .Z(SUM[263]) );
  NANDN U3209 ( .A(n4418), .B(n4419), .Z(n4417) );
  ANDN U3210 ( .B(n4420), .A(n4421), .Z(n4416) );
  NAND U3211 ( .A(n4422), .B(n4423), .Z(n4420) );
  XNOR U3212 ( .A(n4422), .B(n4424), .Z(SUM[262]) );
  NANDN U3213 ( .A(n4421), .B(n4423), .Z(n4424) );
  NANDN U3214 ( .A(n4425), .B(n4426), .Z(n4422) );
  NAND U3215 ( .A(n4427), .B(n4428), .Z(n4426) );
  XNOR U3216 ( .A(n4427), .B(n4429), .Z(SUM[261]) );
  NANDN U3217 ( .A(n4425), .B(n4428), .Z(n4429) );
  NANDN U3218 ( .A(n4430), .B(n4431), .Z(n4427) );
  NANDN U3219 ( .A(n4415), .B(n4432), .Z(n4431) );
  XOR U3220 ( .A(n4415), .B(n4433), .Z(SUM[260]) );
  NANDN U3221 ( .A(n4430), .B(n4432), .Z(n4433) );
  ANDN U3222 ( .B(n4434), .A(n4435), .Z(n4415) );
  OR U3223 ( .A(n4436), .B(n4365), .Z(n4434) );
  XNOR U3224 ( .A(n4382), .B(n4437), .Z(SUM[25]) );
  NANDN U3225 ( .A(n4380), .B(n4383), .Z(n4437) );
  NANDN U3226 ( .A(n4438), .B(n4439), .Z(n4382) );
  NAND U3227 ( .A(n4260), .B(n4440), .Z(n4439) );
  XOR U3228 ( .A(n4441), .B(n4442), .Z(SUM[259]) );
  NANDN U3229 ( .A(n4443), .B(n4444), .Z(n4442) );
  ANDN U3230 ( .B(n4445), .A(n4446), .Z(n4441) );
  NAND U3231 ( .A(n4447), .B(n4448), .Z(n4445) );
  XNOR U3232 ( .A(n4447), .B(n4449), .Z(SUM[258]) );
  NANDN U3233 ( .A(n4446), .B(n4448), .Z(n4449) );
  NANDN U3234 ( .A(n4450), .B(n4451), .Z(n4447) );
  NAND U3235 ( .A(n4452), .B(n4453), .Z(n4451) );
  XNOR U3236 ( .A(n4452), .B(n4454), .Z(SUM[257]) );
  NANDN U3237 ( .A(n4450), .B(n4453), .Z(n4454) );
  NANDN U3238 ( .A(n4455), .B(n4456), .Z(n4452) );
  NANDN U3239 ( .A(n4365), .B(n4457), .Z(n4456) );
  XOR U3240 ( .A(n4365), .B(n4458), .Z(SUM[256]) );
  NANDN U3241 ( .A(n4455), .B(n4457), .Z(n4458) );
  XOR U3242 ( .A(n4459), .B(n4460), .Z(SUM[255]) );
  OR U3243 ( .A(n4461), .B(n4462), .Z(n4460) );
  ANDN U3244 ( .B(n4463), .A(n4464), .Z(n4459) );
  NANDN U3245 ( .A(n4465), .B(n4466), .Z(n4463) );
  XNOR U3246 ( .A(n4466), .B(n4467), .Z(SUM[254]) );
  OR U3247 ( .A(n4465), .B(n4464), .Z(n4467) );
  NANDN U3248 ( .A(n4468), .B(n4469), .Z(n4466) );
  NANDN U3249 ( .A(n4470), .B(n4471), .Z(n4469) );
  XNOR U3250 ( .A(n4471), .B(n4472), .Z(SUM[253]) );
  OR U3251 ( .A(n4470), .B(n4468), .Z(n4472) );
  NANDN U3252 ( .A(n4473), .B(n4474), .Z(n4471) );
  NAND U3253 ( .A(n4475), .B(n4476), .Z(n4474) );
  XNOR U3254 ( .A(n4475), .B(n4477), .Z(SUM[252]) );
  NANDN U3255 ( .A(n4473), .B(n4476), .Z(n4477) );
  NANDN U3256 ( .A(n4478), .B(n4479), .Z(n4475) );
  NANDN U3257 ( .A(n4480), .B(n4481), .Z(n4479) );
  XOR U3258 ( .A(n4482), .B(n4483), .Z(SUM[251]) );
  NANDN U3259 ( .A(n4484), .B(n4485), .Z(n4483) );
  ANDN U3260 ( .B(n4486), .A(n4487), .Z(n4482) );
  NAND U3261 ( .A(n4488), .B(n4489), .Z(n4486) );
  XNOR U3262 ( .A(n4488), .B(n4490), .Z(SUM[250]) );
  NANDN U3263 ( .A(n4487), .B(n4489), .Z(n4490) );
  NANDN U3264 ( .A(n4491), .B(n4492), .Z(n4488) );
  NAND U3265 ( .A(n4493), .B(n4494), .Z(n4492) );
  XNOR U3266 ( .A(n4260), .B(n4495), .Z(SUM[24]) );
  NANDN U3267 ( .A(n4438), .B(n4440), .Z(n4495) );
  NANDN U3268 ( .A(n4496), .B(n4497), .Z(n4260) );
  NANDN U3269 ( .A(n4498), .B(n4499), .Z(n4497) );
  XNOR U3270 ( .A(n4493), .B(n4500), .Z(SUM[249]) );
  NANDN U3271 ( .A(n4491), .B(n4494), .Z(n4500) );
  NANDN U3272 ( .A(n4501), .B(n4502), .Z(n4493) );
  NAND U3273 ( .A(n4481), .B(n4503), .Z(n4502) );
  XNOR U3274 ( .A(n4481), .B(n4504), .Z(SUM[248]) );
  NANDN U3275 ( .A(n4501), .B(n4503), .Z(n4504) );
  NANDN U3276 ( .A(n4505), .B(n4506), .Z(n4481) );
  NANDN U3277 ( .A(n4507), .B(n4508), .Z(n4506) );
  XOR U3278 ( .A(n4509), .B(n4510), .Z(SUM[247]) );
  NANDN U3279 ( .A(n4511), .B(n4512), .Z(n4510) );
  ANDN U3280 ( .B(n4513), .A(n4514), .Z(n4509) );
  NAND U3281 ( .A(n4515), .B(n4516), .Z(n4513) );
  XNOR U3282 ( .A(n4515), .B(n4517), .Z(SUM[246]) );
  NANDN U3283 ( .A(n4514), .B(n4516), .Z(n4517) );
  NANDN U3284 ( .A(n4518), .B(n4519), .Z(n4515) );
  NAND U3285 ( .A(n4520), .B(n4521), .Z(n4519) );
  XNOR U3286 ( .A(n4520), .B(n4522), .Z(SUM[245]) );
  NANDN U3287 ( .A(n4518), .B(n4521), .Z(n4522) );
  NANDN U3288 ( .A(n4523), .B(n4524), .Z(n4520) );
  NANDN U3289 ( .A(n4507), .B(n4525), .Z(n4524) );
  XOR U3290 ( .A(n4507), .B(n4526), .Z(SUM[244]) );
  NANDN U3291 ( .A(n4523), .B(n4525), .Z(n4526) );
  ANDN U3292 ( .B(n4527), .A(n4528), .Z(n4507) );
  OR U3293 ( .A(n4529), .B(n4530), .Z(n4527) );
  XOR U3294 ( .A(n4531), .B(n4532), .Z(SUM[243]) );
  NANDN U3295 ( .A(n4533), .B(n4534), .Z(n4532) );
  ANDN U3296 ( .B(n4535), .A(n4536), .Z(n4531) );
  NANDN U3297 ( .A(n4537), .B(n4538), .Z(n4535) );
  XNOR U3298 ( .A(n4538), .B(n4539), .Z(SUM[242]) );
  OR U3299 ( .A(n4537), .B(n4536), .Z(n4539) );
  NANDN U3300 ( .A(n4540), .B(n4541), .Z(n4538) );
  NAND U3301 ( .A(n4542), .B(n4543), .Z(n4541) );
  XNOR U3302 ( .A(n4542), .B(n4544), .Z(SUM[241]) );
  NANDN U3303 ( .A(n4540), .B(n4543), .Z(n4544) );
  NANDN U3304 ( .A(n4545), .B(n4546), .Z(n4542) );
  NANDN U3305 ( .A(n4530), .B(n4547), .Z(n4546) );
  XOR U3306 ( .A(n4530), .B(n4548), .Z(SUM[240]) );
  NANDN U3307 ( .A(n4545), .B(n4547), .Z(n4548) );
  XOR U3308 ( .A(n4549), .B(n4550), .Z(SUM[23]) );
  NANDN U3309 ( .A(n4551), .B(n4552), .Z(n4550) );
  ANDN U3310 ( .B(n4553), .A(n4554), .Z(n4549) );
  NAND U3311 ( .A(n4555), .B(n4556), .Z(n4553) );
  XOR U3312 ( .A(n4557), .B(n4558), .Z(SUM[239]) );
  OR U3313 ( .A(n4559), .B(n4560), .Z(n4558) );
  ANDN U3314 ( .B(n4561), .A(n4562), .Z(n4557) );
  NANDN U3315 ( .A(n4563), .B(n4564), .Z(n4561) );
  XNOR U3316 ( .A(n4564), .B(n4565), .Z(SUM[238]) );
  OR U3317 ( .A(n4563), .B(n4562), .Z(n4565) );
  NANDN U3318 ( .A(n4566), .B(n4567), .Z(n4564) );
  NANDN U3319 ( .A(n4568), .B(n4569), .Z(n4567) );
  XNOR U3320 ( .A(n4569), .B(n4570), .Z(SUM[237]) );
  OR U3321 ( .A(n4568), .B(n4566), .Z(n4570) );
  NANDN U3322 ( .A(n4571), .B(n4572), .Z(n4569) );
  NAND U3323 ( .A(n4573), .B(n4574), .Z(n4572) );
  XNOR U3324 ( .A(n4573), .B(n4575), .Z(SUM[236]) );
  NANDN U3325 ( .A(n4571), .B(n4574), .Z(n4575) );
  NANDN U3326 ( .A(n4576), .B(n4577), .Z(n4573) );
  NANDN U3327 ( .A(n4578), .B(n4579), .Z(n4577) );
  XOR U3328 ( .A(n4580), .B(n4581), .Z(SUM[235]) );
  NANDN U3329 ( .A(n4582), .B(n4583), .Z(n4581) );
  ANDN U3330 ( .B(n4584), .A(n4585), .Z(n4580) );
  NAND U3331 ( .A(n4586), .B(n4587), .Z(n4584) );
  XNOR U3332 ( .A(n4586), .B(n4588), .Z(SUM[234]) );
  NANDN U3333 ( .A(n4585), .B(n4587), .Z(n4588) );
  NANDN U3334 ( .A(n4589), .B(n4590), .Z(n4586) );
  NAND U3335 ( .A(n4591), .B(n4592), .Z(n4590) );
  XNOR U3336 ( .A(n4591), .B(n4593), .Z(SUM[233]) );
  NANDN U3337 ( .A(n4589), .B(n4592), .Z(n4593) );
  NANDN U3338 ( .A(n4594), .B(n4595), .Z(n4591) );
  NAND U3339 ( .A(n4579), .B(n4596), .Z(n4595) );
  XNOR U3340 ( .A(n4579), .B(n4597), .Z(SUM[232]) );
  NANDN U3341 ( .A(n4594), .B(n4596), .Z(n4597) );
  NANDN U3342 ( .A(n4598), .B(n4599), .Z(n4579) );
  NANDN U3343 ( .A(n4600), .B(n4601), .Z(n4599) );
  XOR U3344 ( .A(n4602), .B(n4603), .Z(SUM[231]) );
  NANDN U3345 ( .A(n4604), .B(n4605), .Z(n4603) );
  ANDN U3346 ( .B(n4606), .A(n4607), .Z(n4602) );
  NAND U3347 ( .A(n4608), .B(n4609), .Z(n4606) );
  XNOR U3348 ( .A(n4608), .B(n4610), .Z(SUM[230]) );
  NANDN U3349 ( .A(n4607), .B(n4609), .Z(n4610) );
  NANDN U3350 ( .A(n4611), .B(n4612), .Z(n4608) );
  NAND U3351 ( .A(n4613), .B(n4614), .Z(n4612) );
  XNOR U3352 ( .A(n4555), .B(n4615), .Z(SUM[22]) );
  NANDN U3353 ( .A(n4554), .B(n4556), .Z(n4615) );
  NANDN U3354 ( .A(n4616), .B(n4617), .Z(n4555) );
  NAND U3355 ( .A(n4618), .B(n4619), .Z(n4617) );
  XNOR U3356 ( .A(n4613), .B(n4620), .Z(SUM[229]) );
  NANDN U3357 ( .A(n4611), .B(n4614), .Z(n4620) );
  NANDN U3358 ( .A(n4621), .B(n4622), .Z(n4613) );
  NANDN U3359 ( .A(n4600), .B(n4623), .Z(n4622) );
  XOR U3360 ( .A(n4600), .B(n4624), .Z(SUM[228]) );
  NANDN U3361 ( .A(n4621), .B(n4623), .Z(n4624) );
  ANDN U3362 ( .B(n4625), .A(n4626), .Z(n4600) );
  OR U3363 ( .A(n4627), .B(n4628), .Z(n4625) );
  XOR U3364 ( .A(n4629), .B(n4630), .Z(SUM[227]) );
  NANDN U3365 ( .A(n4631), .B(n4632), .Z(n4630) );
  ANDN U3366 ( .B(n4633), .A(n4634), .Z(n4629) );
  NANDN U3367 ( .A(n4635), .B(n4636), .Z(n4633) );
  XNOR U3368 ( .A(n4636), .B(n4637), .Z(SUM[226]) );
  OR U3369 ( .A(n4635), .B(n4634), .Z(n4637) );
  NANDN U3370 ( .A(n4638), .B(n4639), .Z(n4636) );
  NAND U3371 ( .A(n4640), .B(n4641), .Z(n4639) );
  XNOR U3372 ( .A(n4640), .B(n4642), .Z(SUM[225]) );
  NANDN U3373 ( .A(n4638), .B(n4641), .Z(n4642) );
  NANDN U3374 ( .A(n4643), .B(n4644), .Z(n4640) );
  NANDN U3375 ( .A(n4628), .B(n4645), .Z(n4644) );
  XOR U3376 ( .A(n4628), .B(n4646), .Z(SUM[224]) );
  NANDN U3377 ( .A(n4643), .B(n4645), .Z(n4646) );
  XOR U3378 ( .A(n4647), .B(n4648), .Z(SUM[223]) );
  OR U3379 ( .A(n4649), .B(n4650), .Z(n4648) );
  ANDN U3380 ( .B(n4651), .A(n4652), .Z(n4647) );
  NANDN U3381 ( .A(n4653), .B(n4654), .Z(n4651) );
  XNOR U3382 ( .A(n4654), .B(n4655), .Z(SUM[222]) );
  OR U3383 ( .A(n4653), .B(n4652), .Z(n4655) );
  NANDN U3384 ( .A(n4656), .B(n4657), .Z(n4654) );
  NANDN U3385 ( .A(n4658), .B(n4659), .Z(n4657) );
  XNOR U3386 ( .A(n4659), .B(n4660), .Z(SUM[221]) );
  OR U3387 ( .A(n4658), .B(n4656), .Z(n4660) );
  NANDN U3388 ( .A(n4661), .B(n4662), .Z(n4659) );
  NAND U3389 ( .A(n4663), .B(n4664), .Z(n4662) );
  XNOR U3390 ( .A(n4663), .B(n4665), .Z(SUM[220]) );
  NANDN U3391 ( .A(n4661), .B(n4664), .Z(n4665) );
  NANDN U3392 ( .A(n4666), .B(n4667), .Z(n4663) );
  NANDN U3393 ( .A(n4668), .B(n4669), .Z(n4667) );
  XNOR U3394 ( .A(n4618), .B(n4670), .Z(SUM[21]) );
  NANDN U3395 ( .A(n4616), .B(n4619), .Z(n4670) );
  NANDN U3396 ( .A(n4671), .B(n4672), .Z(n4618) );
  NANDN U3397 ( .A(n4498), .B(n4673), .Z(n4672) );
  XOR U3398 ( .A(n4674), .B(n4675), .Z(SUM[219]) );
  NANDN U3399 ( .A(n4676), .B(n4677), .Z(n4675) );
  ANDN U3400 ( .B(n4678), .A(n4679), .Z(n4674) );
  NAND U3401 ( .A(n4680), .B(n4681), .Z(n4678) );
  XNOR U3402 ( .A(n4680), .B(n4682), .Z(SUM[218]) );
  NANDN U3403 ( .A(n4679), .B(n4681), .Z(n4682) );
  NANDN U3404 ( .A(n4683), .B(n4684), .Z(n4680) );
  NAND U3405 ( .A(n4685), .B(n4686), .Z(n4684) );
  XNOR U3406 ( .A(n4685), .B(n4687), .Z(SUM[217]) );
  NANDN U3407 ( .A(n4683), .B(n4686), .Z(n4687) );
  NANDN U3408 ( .A(n4688), .B(n4689), .Z(n4685) );
  NAND U3409 ( .A(n4669), .B(n4690), .Z(n4689) );
  XNOR U3410 ( .A(n4669), .B(n4691), .Z(SUM[216]) );
  NANDN U3411 ( .A(n4688), .B(n4690), .Z(n4691) );
  NANDN U3412 ( .A(n4692), .B(n4693), .Z(n4669) );
  NANDN U3413 ( .A(n4694), .B(n4695), .Z(n4693) );
  XOR U3414 ( .A(n4696), .B(n4697), .Z(SUM[215]) );
  NANDN U3415 ( .A(n4698), .B(n4699), .Z(n4697) );
  ANDN U3416 ( .B(n4700), .A(n4701), .Z(n4696) );
  NAND U3417 ( .A(n4702), .B(n4703), .Z(n4700) );
  XNOR U3418 ( .A(n4702), .B(n4704), .Z(SUM[214]) );
  NANDN U3419 ( .A(n4701), .B(n4703), .Z(n4704) );
  NANDN U3420 ( .A(n4705), .B(n4706), .Z(n4702) );
  NAND U3421 ( .A(n4707), .B(n4708), .Z(n4706) );
  XNOR U3422 ( .A(n4707), .B(n4709), .Z(SUM[213]) );
  NANDN U3423 ( .A(n4705), .B(n4708), .Z(n4709) );
  NANDN U3424 ( .A(n4710), .B(n4711), .Z(n4707) );
  NANDN U3425 ( .A(n4694), .B(n4712), .Z(n4711) );
  XOR U3426 ( .A(n4694), .B(n4713), .Z(SUM[212]) );
  NANDN U3427 ( .A(n4710), .B(n4712), .Z(n4713) );
  ANDN U3428 ( .B(n4714), .A(n4715), .Z(n4694) );
  OR U3429 ( .A(n4716), .B(n4717), .Z(n4714) );
  XOR U3430 ( .A(n4718), .B(n4719), .Z(SUM[211]) );
  NANDN U3431 ( .A(n4720), .B(n4721), .Z(n4719) );
  ANDN U3432 ( .B(n4722), .A(n4723), .Z(n4718) );
  NANDN U3433 ( .A(n4724), .B(n4725), .Z(n4722) );
  XNOR U3434 ( .A(n4725), .B(n4726), .Z(SUM[210]) );
  OR U3435 ( .A(n4724), .B(n4723), .Z(n4726) );
  NANDN U3436 ( .A(n4727), .B(n4728), .Z(n4725) );
  NAND U3437 ( .A(n4729), .B(n4730), .Z(n4728) );
  XOR U3438 ( .A(n4498), .B(n4731), .Z(SUM[20]) );
  NANDN U3439 ( .A(n4671), .B(n4673), .Z(n4731) );
  ANDN U3440 ( .B(n4732), .A(n4733), .Z(n4498) );
  OR U3441 ( .A(n4734), .B(n4735), .Z(n4732) );
  XNOR U3442 ( .A(n4729), .B(n4736), .Z(SUM[209]) );
  NANDN U3443 ( .A(n4727), .B(n4730), .Z(n4736) );
  NANDN U3444 ( .A(n4737), .B(n4738), .Z(n4729) );
  NANDN U3445 ( .A(n4717), .B(n4739), .Z(n4738) );
  XOR U3446 ( .A(n4717), .B(n4740), .Z(SUM[208]) );
  NANDN U3447 ( .A(n4737), .B(n4739), .Z(n4740) );
  XOR U3448 ( .A(n4741), .B(n4742), .Z(SUM[207]) );
  OR U3449 ( .A(n4743), .B(n4744), .Z(n4742) );
  ANDN U3450 ( .B(n4745), .A(n4746), .Z(n4741) );
  NANDN U3451 ( .A(n4747), .B(n4748), .Z(n4745) );
  XNOR U3452 ( .A(n4748), .B(n4749), .Z(SUM[206]) );
  OR U3453 ( .A(n4747), .B(n4746), .Z(n4749) );
  NANDN U3454 ( .A(n4750), .B(n4751), .Z(n4748) );
  NANDN U3455 ( .A(n4752), .B(n4753), .Z(n4751) );
  XNOR U3456 ( .A(n4753), .B(n4754), .Z(SUM[205]) );
  OR U3457 ( .A(n4752), .B(n4750), .Z(n4754) );
  NANDN U3458 ( .A(n4755), .B(n4756), .Z(n4753) );
  NAND U3459 ( .A(n4757), .B(n4758), .Z(n4756) );
  XNOR U3460 ( .A(n4757), .B(n4759), .Z(SUM[204]) );
  NANDN U3461 ( .A(n4755), .B(n4758), .Z(n4759) );
  NANDN U3462 ( .A(n4760), .B(n4761), .Z(n4757) );
  NANDN U3463 ( .A(n4762), .B(n4763), .Z(n4761) );
  XOR U3464 ( .A(n4764), .B(n4765), .Z(SUM[203]) );
  NANDN U3465 ( .A(n4766), .B(n4767), .Z(n4765) );
  ANDN U3466 ( .B(n4768), .A(n4769), .Z(n4764) );
  NAND U3467 ( .A(n4770), .B(n4771), .Z(n4768) );
  XNOR U3468 ( .A(n4770), .B(n4772), .Z(SUM[202]) );
  NANDN U3469 ( .A(n4769), .B(n4771), .Z(n4772) );
  NANDN U3470 ( .A(n4773), .B(n4774), .Z(n4770) );
  NAND U3471 ( .A(n4775), .B(n4776), .Z(n4774) );
  XNOR U3472 ( .A(n4775), .B(n4777), .Z(SUM[201]) );
  NANDN U3473 ( .A(n4773), .B(n4776), .Z(n4777) );
  NANDN U3474 ( .A(n4778), .B(n4779), .Z(n4775) );
  NAND U3475 ( .A(n4763), .B(n4780), .Z(n4779) );
  XNOR U3476 ( .A(n4763), .B(n4781), .Z(SUM[200]) );
  NANDN U3477 ( .A(n4778), .B(n4780), .Z(n4781) );
  NANDN U3478 ( .A(n4782), .B(n4783), .Z(n4763) );
  NANDN U3479 ( .A(n4784), .B(n4785), .Z(n4783) );
  XOR U3480 ( .A(n4786), .B(n4787), .Z(SUM[19]) );
  NANDN U3481 ( .A(n4788), .B(n4789), .Z(n4787) );
  ANDN U3482 ( .B(n4790), .A(n4791), .Z(n4786) );
  NANDN U3483 ( .A(n4792), .B(n4793), .Z(n4790) );
  XOR U3484 ( .A(n4794), .B(n4795), .Z(SUM[199]) );
  NANDN U3485 ( .A(n4796), .B(n4797), .Z(n4795) );
  ANDN U3486 ( .B(n4798), .A(n4799), .Z(n4794) );
  NAND U3487 ( .A(n4800), .B(n4801), .Z(n4798) );
  XNOR U3488 ( .A(n4800), .B(n4802), .Z(SUM[198]) );
  NANDN U3489 ( .A(n4799), .B(n4801), .Z(n4802) );
  NANDN U3490 ( .A(n4803), .B(n4804), .Z(n4800) );
  NAND U3491 ( .A(n4805), .B(n4806), .Z(n4804) );
  XNOR U3492 ( .A(n4805), .B(n4807), .Z(SUM[197]) );
  NANDN U3493 ( .A(n4803), .B(n4806), .Z(n4807) );
  NANDN U3494 ( .A(n4808), .B(n4809), .Z(n4805) );
  NANDN U3495 ( .A(n4784), .B(n4810), .Z(n4809) );
  XOR U3496 ( .A(n4784), .B(n4811), .Z(SUM[196]) );
  NANDN U3497 ( .A(n4808), .B(n4810), .Z(n4811) );
  ANDN U3498 ( .B(n4812), .A(n4813), .Z(n4784) );
  OR U3499 ( .A(n4814), .B(n4815), .Z(n4812) );
  XOR U3500 ( .A(n4816), .B(n4817), .Z(SUM[195]) );
  NANDN U3501 ( .A(n4818), .B(n4819), .Z(n4817) );
  ANDN U3502 ( .B(n4820), .A(n4821), .Z(n4816) );
  NANDN U3503 ( .A(n4822), .B(n4823), .Z(n4820) );
  XNOR U3504 ( .A(n4823), .B(n4824), .Z(SUM[194]) );
  OR U3505 ( .A(n4822), .B(n4821), .Z(n4824) );
  NANDN U3506 ( .A(n4825), .B(n4826), .Z(n4823) );
  NAND U3507 ( .A(n4827), .B(n4828), .Z(n4826) );
  XNOR U3508 ( .A(n4827), .B(n4829), .Z(SUM[193]) );
  NANDN U3509 ( .A(n4825), .B(n4828), .Z(n4829) );
  NANDN U3510 ( .A(n4830), .B(n4831), .Z(n4827) );
  NANDN U3511 ( .A(n4815), .B(n4832), .Z(n4831) );
  XOR U3512 ( .A(n4815), .B(n4833), .Z(SUM[192]) );
  NANDN U3513 ( .A(n4830), .B(n4832), .Z(n4833) );
  XOR U3514 ( .A(n4834), .B(n4835), .Z(SUM[191]) );
  OR U3515 ( .A(n4836), .B(n4837), .Z(n4835) );
  ANDN U3516 ( .B(n4838), .A(n4839), .Z(n4834) );
  NAND U3517 ( .A(n4840), .B(n4841), .Z(n4838) );
  XNOR U3518 ( .A(n4840), .B(n4842), .Z(SUM[190]) );
  NANDN U3519 ( .A(n4839), .B(n4841), .Z(n4842) );
  NANDN U3520 ( .A(n4843), .B(n4844), .Z(n4840) );
  NAND U3521 ( .A(n4845), .B(n4846), .Z(n4844) );
  XNOR U3522 ( .A(n4793), .B(n4847), .Z(SUM[18]) );
  OR U3523 ( .A(n4792), .B(n4791), .Z(n4847) );
  NANDN U3524 ( .A(n4848), .B(n4849), .Z(n4793) );
  NAND U3525 ( .A(n4850), .B(n4851), .Z(n4849) );
  XNOR U3526 ( .A(n4845), .B(n4852), .Z(SUM[189]) );
  NANDN U3527 ( .A(n4843), .B(n4846), .Z(n4852) );
  NANDN U3528 ( .A(n4853), .B(n4854), .Z(n4845) );
  NANDN U3529 ( .A(n4855), .B(n4856), .Z(n4854) );
  XNOR U3530 ( .A(n4856), .B(n4857), .Z(SUM[188]) );
  OR U3531 ( .A(n4855), .B(n4853), .Z(n4857) );
  NANDN U3532 ( .A(n4858), .B(n4859), .Z(n4856) );
  NANDN U3533 ( .A(n4860), .B(n4861), .Z(n4859) );
  XOR U3534 ( .A(n4862), .B(n4863), .Z(SUM[187]) );
  NANDN U3535 ( .A(n4864), .B(n4865), .Z(n4863) );
  ANDN U3536 ( .B(n4866), .A(n4867), .Z(n4862) );
  NAND U3537 ( .A(n4868), .B(n4869), .Z(n4866) );
  XNOR U3538 ( .A(n4868), .B(n4870), .Z(SUM[186]) );
  NANDN U3539 ( .A(n4867), .B(n4869), .Z(n4870) );
  NANDN U3540 ( .A(n4871), .B(n4872), .Z(n4868) );
  NAND U3541 ( .A(n4873), .B(n4874), .Z(n4872) );
  XNOR U3542 ( .A(n4873), .B(n4875), .Z(SUM[185]) );
  NANDN U3543 ( .A(n4871), .B(n4874), .Z(n4875) );
  NANDN U3544 ( .A(n4876), .B(n4877), .Z(n4873) );
  NAND U3545 ( .A(n4861), .B(n4878), .Z(n4877) );
  XNOR U3546 ( .A(n4861), .B(n4879), .Z(SUM[184]) );
  NANDN U3547 ( .A(n4876), .B(n4878), .Z(n4879) );
  NANDN U3548 ( .A(n4880), .B(n4881), .Z(n4861) );
  NANDN U3549 ( .A(n4882), .B(n4883), .Z(n4881) );
  XOR U3550 ( .A(n4884), .B(n4885), .Z(SUM[183]) );
  NANDN U3551 ( .A(n4886), .B(n4887), .Z(n4885) );
  ANDN U3552 ( .B(n4888), .A(n4889), .Z(n4884) );
  NAND U3553 ( .A(n4890), .B(n4891), .Z(n4888) );
  XNOR U3554 ( .A(n4890), .B(n4892), .Z(SUM[182]) );
  NANDN U3555 ( .A(n4889), .B(n4891), .Z(n4892) );
  NANDN U3556 ( .A(n4893), .B(n4894), .Z(n4890) );
  NAND U3557 ( .A(n4895), .B(n4896), .Z(n4894) );
  XNOR U3558 ( .A(n4895), .B(n4897), .Z(SUM[181]) );
  NANDN U3559 ( .A(n4893), .B(n4896), .Z(n4897) );
  NANDN U3560 ( .A(n4898), .B(n4899), .Z(n4895) );
  NANDN U3561 ( .A(n4882), .B(n4900), .Z(n4899) );
  XOR U3562 ( .A(n4882), .B(n4901), .Z(SUM[180]) );
  NANDN U3563 ( .A(n4898), .B(n4900), .Z(n4901) );
  ANDN U3564 ( .B(n4902), .A(n4903), .Z(n4882) );
  NANDN U3565 ( .A(n4904), .B(n4905), .Z(n4902) );
  XNOR U3566 ( .A(n4850), .B(n4906), .Z(SUM[17]) );
  NANDN U3567 ( .A(n4848), .B(n4851), .Z(n4906) );
  NANDN U3568 ( .A(n4907), .B(n4908), .Z(n4850) );
  NANDN U3569 ( .A(n4735), .B(n4909), .Z(n4908) );
  XOR U3570 ( .A(n4910), .B(n4911), .Z(SUM[179]) );
  NANDN U3571 ( .A(n4912), .B(n4913), .Z(n4911) );
  ANDN U3572 ( .B(n4914), .A(n4915), .Z(n4910) );
  NANDN U3573 ( .A(n4916), .B(n4917), .Z(n4914) );
  XNOR U3574 ( .A(n4917), .B(n4918), .Z(SUM[178]) );
  OR U3575 ( .A(n4916), .B(n4915), .Z(n4918) );
  NANDN U3576 ( .A(n4919), .B(n4920), .Z(n4917) );
  NAND U3577 ( .A(n4921), .B(n4922), .Z(n4920) );
  XNOR U3578 ( .A(n4921), .B(n4923), .Z(SUM[177]) );
  NANDN U3579 ( .A(n4919), .B(n4922), .Z(n4923) );
  NANDN U3580 ( .A(n4924), .B(n4925), .Z(n4921) );
  NAND U3581 ( .A(n4905), .B(n4926), .Z(n4925) );
  XNOR U3582 ( .A(n4905), .B(n4927), .Z(SUM[176]) );
  NANDN U3583 ( .A(n4924), .B(n4926), .Z(n4927) );
  XOR U3584 ( .A(n4928), .B(n4929), .Z(SUM[175]) );
  NANDN U3585 ( .A(n4930), .B(n4931), .Z(n4929) );
  ANDN U3586 ( .B(n4932), .A(n4933), .Z(n4928) );
  NAND U3587 ( .A(n4934), .B(n4935), .Z(n4932) );
  XNOR U3588 ( .A(n4934), .B(n4936), .Z(SUM[174]) );
  NANDN U3589 ( .A(n4933), .B(n4935), .Z(n4936) );
  NANDN U3590 ( .A(n4937), .B(n4938), .Z(n4934) );
  NAND U3591 ( .A(n4939), .B(n4940), .Z(n4938) );
  XNOR U3592 ( .A(n4939), .B(n4941), .Z(SUM[173]) );
  NANDN U3593 ( .A(n4937), .B(n4940), .Z(n4941) );
  NANDN U3594 ( .A(n4942), .B(n4943), .Z(n4939) );
  NAND U3595 ( .A(n4944), .B(n4945), .Z(n4943) );
  XNOR U3596 ( .A(n4944), .B(n4946), .Z(SUM[172]) );
  NANDN U3597 ( .A(n4942), .B(n4945), .Z(n4946) );
  NANDN U3598 ( .A(n4947), .B(n4948), .Z(n4944) );
  NAND U3599 ( .A(n4949), .B(n4950), .Z(n4948) );
  XOR U3600 ( .A(n4951), .B(n4952), .Z(SUM[171]) );
  NANDN U3601 ( .A(n4953), .B(n4954), .Z(n4952) );
  ANDN U3602 ( .B(n4955), .A(n4956), .Z(n4951) );
  NAND U3603 ( .A(n4957), .B(n4958), .Z(n4955) );
  XNOR U3604 ( .A(n4957), .B(n4959), .Z(SUM[170]) );
  NANDN U3605 ( .A(n4956), .B(n4958), .Z(n4959) );
  NANDN U3606 ( .A(n4960), .B(n4961), .Z(n4957) );
  NAND U3607 ( .A(n4962), .B(n4963), .Z(n4961) );
  XOR U3608 ( .A(n4735), .B(n4964), .Z(SUM[16]) );
  NANDN U3609 ( .A(n4907), .B(n4909), .Z(n4964) );
  XNOR U3610 ( .A(n4962), .B(n4965), .Z(SUM[169]) );
  NANDN U3611 ( .A(n4960), .B(n4963), .Z(n4965) );
  NANDN U3612 ( .A(n4966), .B(n4967), .Z(n4962) );
  NAND U3613 ( .A(n4950), .B(n4968), .Z(n4967) );
  XNOR U3614 ( .A(n4950), .B(n4969), .Z(SUM[168]) );
  NANDN U3615 ( .A(n4966), .B(n4968), .Z(n4969) );
  NANDN U3616 ( .A(n4970), .B(n4971), .Z(n4950) );
  OR U3617 ( .A(n4972), .B(n4973), .Z(n4971) );
  XOR U3618 ( .A(n4974), .B(n4975), .Z(SUM[167]) );
  NANDN U3619 ( .A(n4976), .B(n4977), .Z(n4975) );
  ANDN U3620 ( .B(n4978), .A(n4979), .Z(n4974) );
  NAND U3621 ( .A(n4980), .B(n4981), .Z(n4978) );
  XNOR U3622 ( .A(n4980), .B(n4982), .Z(SUM[166]) );
  NANDN U3623 ( .A(n4979), .B(n4981), .Z(n4982) );
  NANDN U3624 ( .A(n4983), .B(n4984), .Z(n4980) );
  NAND U3625 ( .A(n4985), .B(n4986), .Z(n4984) );
  XNOR U3626 ( .A(n4985), .B(n4987), .Z(SUM[165]) );
  NANDN U3627 ( .A(n4983), .B(n4986), .Z(n4987) );
  NANDN U3628 ( .A(n4988), .B(n4989), .Z(n4985) );
  NANDN U3629 ( .A(n4973), .B(n4990), .Z(n4989) );
  XOR U3630 ( .A(n4973), .B(n4991), .Z(SUM[164]) );
  NANDN U3631 ( .A(n4988), .B(n4990), .Z(n4991) );
  ANDN U3632 ( .B(n4992), .A(n4993), .Z(n4973) );
  NANDN U3633 ( .A(n4994), .B(n4995), .Z(n4992) );
  XOR U3634 ( .A(n4996), .B(n4997), .Z(SUM[163]) );
  NANDN U3635 ( .A(n4998), .B(n4999), .Z(n4997) );
  ANDN U3636 ( .B(n5000), .A(n5001), .Z(n4996) );
  NAND U3637 ( .A(n5002), .B(n5003), .Z(n5000) );
  XNOR U3638 ( .A(n5002), .B(n5004), .Z(SUM[162]) );
  NANDN U3639 ( .A(n5001), .B(n5003), .Z(n5004) );
  NANDN U3640 ( .A(n5005), .B(n5006), .Z(n5002) );
  NAND U3641 ( .A(n5007), .B(n5008), .Z(n5006) );
  XNOR U3642 ( .A(n5007), .B(n5009), .Z(SUM[161]) );
  NANDN U3643 ( .A(n5005), .B(n5008), .Z(n5009) );
  NANDN U3644 ( .A(n5010), .B(n5011), .Z(n5007) );
  NAND U3645 ( .A(n4995), .B(n5012), .Z(n5011) );
  XNOR U3646 ( .A(n4995), .B(n5013), .Z(SUM[160]) );
  NANDN U3647 ( .A(n5010), .B(n5012), .Z(n5013) );
  XNOR U3648 ( .A(n5014), .B(n5015), .Z(SUM[15]) );
  NANDN U3649 ( .A(n5016), .B(n5017), .Z(n5015) );
  XOR U3650 ( .A(n5018), .B(n5019), .Z(SUM[159]) );
  NANDN U3651 ( .A(n5020), .B(n5021), .Z(n5019) );
  ANDN U3652 ( .B(n5022), .A(n5023), .Z(n5018) );
  NAND U3653 ( .A(n5024), .B(n5025), .Z(n5022) );
  XNOR U3654 ( .A(n5024), .B(n5026), .Z(SUM[158]) );
  NANDN U3655 ( .A(n5023), .B(n5025), .Z(n5026) );
  NANDN U3656 ( .A(n5027), .B(n5028), .Z(n5024) );
  NAND U3657 ( .A(n5029), .B(n5030), .Z(n5028) );
  XNOR U3658 ( .A(n5029), .B(n5031), .Z(SUM[157]) );
  NANDN U3659 ( .A(n5027), .B(n5030), .Z(n5031) );
  NANDN U3660 ( .A(n5032), .B(n5033), .Z(n5029) );
  NAND U3661 ( .A(n5034), .B(n5035), .Z(n5033) );
  XNOR U3662 ( .A(n5034), .B(n5036), .Z(SUM[156]) );
  NANDN U3663 ( .A(n5032), .B(n5035), .Z(n5036) );
  NANDN U3664 ( .A(n5037), .B(n5038), .Z(n5034) );
  NAND U3665 ( .A(n5039), .B(n5040), .Z(n5038) );
  XOR U3666 ( .A(n5041), .B(n5042), .Z(SUM[155]) );
  NANDN U3667 ( .A(n5043), .B(n5044), .Z(n5042) );
  ANDN U3668 ( .B(n5045), .A(n5046), .Z(n5041) );
  NAND U3669 ( .A(n5047), .B(n5048), .Z(n5045) );
  XNOR U3670 ( .A(n5047), .B(n5049), .Z(SUM[154]) );
  NANDN U3671 ( .A(n5046), .B(n5048), .Z(n5049) );
  NANDN U3672 ( .A(n5050), .B(n5051), .Z(n5047) );
  NAND U3673 ( .A(n5052), .B(n5053), .Z(n5051) );
  XNOR U3674 ( .A(n5052), .B(n5054), .Z(SUM[153]) );
  NANDN U3675 ( .A(n5050), .B(n5053), .Z(n5054) );
  NANDN U3676 ( .A(n5055), .B(n5056), .Z(n5052) );
  NAND U3677 ( .A(n5040), .B(n5057), .Z(n5056) );
  XNOR U3678 ( .A(n5040), .B(n5058), .Z(SUM[152]) );
  NANDN U3679 ( .A(n5055), .B(n5057), .Z(n5058) );
  NANDN U3680 ( .A(n5059), .B(n5060), .Z(n5040) );
  OR U3681 ( .A(n5061), .B(n5062), .Z(n5060) );
  XOR U3682 ( .A(n5063), .B(n5064), .Z(SUM[151]) );
  NANDN U3683 ( .A(n5065), .B(n5066), .Z(n5064) );
  ANDN U3684 ( .B(n5067), .A(n5068), .Z(n5063) );
  NAND U3685 ( .A(n5069), .B(n5070), .Z(n5067) );
  XNOR U3686 ( .A(n5069), .B(n5071), .Z(SUM[150]) );
  NANDN U3687 ( .A(n5068), .B(n5070), .Z(n5071) );
  NANDN U3688 ( .A(n5072), .B(n5073), .Z(n5069) );
  NAND U3689 ( .A(n5074), .B(n5075), .Z(n5073) );
  XNOR U3690 ( .A(n5076), .B(n5077), .Z(SUM[14]) );
  NANDN U3691 ( .A(n5078), .B(n5079), .Z(n5077) );
  XNOR U3692 ( .A(n5074), .B(n5080), .Z(SUM[149]) );
  NANDN U3693 ( .A(n5072), .B(n5075), .Z(n5080) );
  NANDN U3694 ( .A(n5081), .B(n5082), .Z(n5074) );
  NANDN U3695 ( .A(n5062), .B(n5083), .Z(n5082) );
  XOR U3696 ( .A(n5062), .B(n5084), .Z(SUM[148]) );
  NANDN U3697 ( .A(n5081), .B(n5083), .Z(n5084) );
  ANDN U3698 ( .B(n5085), .A(n5086), .Z(n5062) );
  NANDN U3699 ( .A(n5087), .B(n5088), .Z(n5085) );
  XOR U3700 ( .A(n5089), .B(n5090), .Z(SUM[147]) );
  NANDN U3701 ( .A(n5091), .B(n5092), .Z(n5090) );
  ANDN U3702 ( .B(n5093), .A(n5094), .Z(n5089) );
  NAND U3703 ( .A(n5095), .B(n5096), .Z(n5093) );
  XNOR U3704 ( .A(n5095), .B(n5097), .Z(SUM[146]) );
  NANDN U3705 ( .A(n5094), .B(n5096), .Z(n5097) );
  NANDN U3706 ( .A(n5098), .B(n5099), .Z(n5095) );
  NAND U3707 ( .A(n5100), .B(n5101), .Z(n5099) );
  XNOR U3708 ( .A(n5100), .B(n5102), .Z(SUM[145]) );
  NANDN U3709 ( .A(n5098), .B(n5101), .Z(n5102) );
  NANDN U3710 ( .A(n5103), .B(n5104), .Z(n5100) );
  NAND U3711 ( .A(n5088), .B(n5105), .Z(n5104) );
  XNOR U3712 ( .A(n5088), .B(n5106), .Z(SUM[144]) );
  NANDN U3713 ( .A(n5103), .B(n5105), .Z(n5106) );
  XOR U3714 ( .A(n5107), .B(n5108), .Z(SUM[143]) );
  NANDN U3715 ( .A(n5109), .B(n5110), .Z(n5108) );
  ANDN U3716 ( .B(n5111), .A(n5112), .Z(n5107) );
  NAND U3717 ( .A(n5113), .B(n5114), .Z(n5111) );
  XNOR U3718 ( .A(n5113), .B(n5115), .Z(SUM[142]) );
  NANDN U3719 ( .A(n5112), .B(n5114), .Z(n5115) );
  NANDN U3720 ( .A(n5116), .B(n5117), .Z(n5113) );
  NAND U3721 ( .A(n5118), .B(n5119), .Z(n5117) );
  XNOR U3722 ( .A(n5118), .B(n5120), .Z(SUM[141]) );
  NANDN U3723 ( .A(n5116), .B(n5119), .Z(n5120) );
  NANDN U3724 ( .A(n5121), .B(n5122), .Z(n5118) );
  NAND U3725 ( .A(n5123), .B(n5124), .Z(n5122) );
  XNOR U3726 ( .A(n5123), .B(n5125), .Z(SUM[140]) );
  NANDN U3727 ( .A(n5121), .B(n5124), .Z(n5125) );
  NANDN U3728 ( .A(n5126), .B(n5127), .Z(n5123) );
  NAND U3729 ( .A(n5128), .B(n5129), .Z(n5127) );
  XNOR U3730 ( .A(n5130), .B(n5131), .Z(SUM[13]) );
  NANDN U3731 ( .A(n5132), .B(n5133), .Z(n5131) );
  XOR U3732 ( .A(n5134), .B(n5135), .Z(SUM[139]) );
  NANDN U3733 ( .A(n5136), .B(n5137), .Z(n5135) );
  ANDN U3734 ( .B(n5138), .A(n5139), .Z(n5134) );
  NAND U3735 ( .A(n5140), .B(n5141), .Z(n5138) );
  XNOR U3736 ( .A(n5140), .B(n5142), .Z(SUM[138]) );
  NANDN U3737 ( .A(n5139), .B(n5141), .Z(n5142) );
  NANDN U3738 ( .A(n5143), .B(n5144), .Z(n5140) );
  NAND U3739 ( .A(n5145), .B(n5146), .Z(n5144) );
  XNOR U3740 ( .A(n5145), .B(n5147), .Z(SUM[137]) );
  NANDN U3741 ( .A(n5143), .B(n5146), .Z(n5147) );
  NANDN U3742 ( .A(n5148), .B(n5149), .Z(n5145) );
  NAND U3743 ( .A(n5129), .B(n5150), .Z(n5149) );
  XNOR U3744 ( .A(n5129), .B(n5151), .Z(SUM[136]) );
  NANDN U3745 ( .A(n5148), .B(n5150), .Z(n5151) );
  NANDN U3746 ( .A(n5152), .B(n5153), .Z(n5129) );
  OR U3747 ( .A(n5154), .B(n5155), .Z(n5153) );
  XOR U3748 ( .A(n5156), .B(n5157), .Z(SUM[135]) );
  NANDN U3749 ( .A(n5158), .B(n5159), .Z(n5157) );
  ANDN U3750 ( .B(n5160), .A(n5161), .Z(n5156) );
  NAND U3751 ( .A(n5162), .B(n5163), .Z(n5160) );
  XNOR U3752 ( .A(n5162), .B(n5164), .Z(SUM[134]) );
  NANDN U3753 ( .A(n5161), .B(n5163), .Z(n5164) );
  NANDN U3754 ( .A(n5165), .B(n5166), .Z(n5162) );
  NAND U3755 ( .A(n5167), .B(n5168), .Z(n5166) );
  XNOR U3756 ( .A(n5167), .B(n5169), .Z(SUM[133]) );
  NANDN U3757 ( .A(n5165), .B(n5168), .Z(n5169) );
  NANDN U3758 ( .A(n5170), .B(n5171), .Z(n5167) );
  NANDN U3759 ( .A(n5155), .B(n5172), .Z(n5171) );
  XOR U3760 ( .A(n5155), .B(n5173), .Z(SUM[132]) );
  NANDN U3761 ( .A(n5170), .B(n5172), .Z(n5173) );
  ANDN U3762 ( .B(n5174), .A(n5175), .Z(n5155) );
  OR U3763 ( .A(n5176), .B(n5177), .Z(n5174) );
  XOR U3764 ( .A(n5178), .B(n5179), .Z(SUM[131]) );
  NANDN U3765 ( .A(n5180), .B(n5181), .Z(n5179) );
  ANDN U3766 ( .B(n5182), .A(n5183), .Z(n5178) );
  NAND U3767 ( .A(n5184), .B(n5185), .Z(n5182) );
  XNOR U3768 ( .A(n5184), .B(n5186), .Z(SUM[130]) );
  NANDN U3769 ( .A(n5183), .B(n5185), .Z(n5186) );
  NANDN U3770 ( .A(n5187), .B(n5188), .Z(n5184) );
  NAND U3771 ( .A(n5189), .B(n5190), .Z(n5188) );
  XNOR U3772 ( .A(n5191), .B(n5192), .Z(SUM[12]) );
  NANDN U3773 ( .A(n5193), .B(n5194), .Z(n5192) );
  XNOR U3774 ( .A(n5189), .B(n5195), .Z(SUM[129]) );
  NANDN U3775 ( .A(n5187), .B(n5190), .Z(n5195) );
  NANDN U3776 ( .A(n5196), .B(n5197), .Z(n5189) );
  NANDN U3777 ( .A(n5177), .B(n5198), .Z(n5197) );
  XOR U3778 ( .A(n5177), .B(n5199), .Z(SUM[128]) );
  NANDN U3779 ( .A(n5196), .B(n5198), .Z(n5199) );
  XOR U3780 ( .A(n5200), .B(n5201), .Z(SUM[127]) );
  OR U3781 ( .A(n5202), .B(n5203), .Z(n5201) );
  ANDN U3782 ( .B(n5204), .A(n5205), .Z(n5200) );
  NAND U3783 ( .A(n5206), .B(n5207), .Z(n5204) );
  XNOR U3784 ( .A(n5206), .B(n5208), .Z(SUM[126]) );
  NANDN U3785 ( .A(n5205), .B(n5207), .Z(n5208) );
  NANDN U3786 ( .A(n5209), .B(n5210), .Z(n5206) );
  NAND U3787 ( .A(n5211), .B(n5212), .Z(n5210) );
  XNOR U3788 ( .A(n5211), .B(n5213), .Z(SUM[125]) );
  NANDN U3789 ( .A(n5209), .B(n5212), .Z(n5213) );
  NANDN U3790 ( .A(n5214), .B(n5215), .Z(n5211) );
  NANDN U3791 ( .A(n5216), .B(n5217), .Z(n5215) );
  XNOR U3792 ( .A(n5217), .B(n5218), .Z(SUM[124]) );
  OR U3793 ( .A(n5216), .B(n5214), .Z(n5218) );
  NANDN U3794 ( .A(n5219), .B(n5220), .Z(n5217) );
  NANDN U3795 ( .A(n5221), .B(n5222), .Z(n5220) );
  XOR U3796 ( .A(n5223), .B(n5224), .Z(SUM[123]) );
  NANDN U3797 ( .A(n5225), .B(n5226), .Z(n5224) );
  ANDN U3798 ( .B(n5227), .A(n5228), .Z(n5223) );
  NAND U3799 ( .A(n5229), .B(n5230), .Z(n5227) );
  XNOR U3800 ( .A(n5229), .B(n5231), .Z(SUM[122]) );
  NANDN U3801 ( .A(n5228), .B(n5230), .Z(n5231) );
  NANDN U3802 ( .A(n5232), .B(n5233), .Z(n5229) );
  NAND U3803 ( .A(n5234), .B(n5235), .Z(n5233) );
  XNOR U3804 ( .A(n5234), .B(n5236), .Z(SUM[121]) );
  NANDN U3805 ( .A(n5232), .B(n5235), .Z(n5236) );
  NANDN U3806 ( .A(n5237), .B(n5238), .Z(n5234) );
  NAND U3807 ( .A(n5222), .B(n5239), .Z(n5238) );
  XNOR U3808 ( .A(n5222), .B(n5240), .Z(SUM[120]) );
  NANDN U3809 ( .A(n5237), .B(n5239), .Z(n5240) );
  NANDN U3810 ( .A(n5241), .B(n5242), .Z(n5222) );
  NANDN U3811 ( .A(n5243), .B(n5244), .Z(n5242) );
  XOR U3812 ( .A(n5245), .B(n5246), .Z(SUM[11]) );
  OR U3813 ( .A(n5247), .B(n5248), .Z(n5246) );
  ANDN U3814 ( .B(n5249), .A(n5250), .Z(n5245) );
  NANDN U3815 ( .A(n5251), .B(n5252), .Z(n5249) );
  XOR U3816 ( .A(n5253), .B(n5254), .Z(SUM[119]) );
  NANDN U3817 ( .A(n5255), .B(n5256), .Z(n5254) );
  ANDN U3818 ( .B(n5257), .A(n5258), .Z(n5253) );
  NAND U3819 ( .A(n5259), .B(n5260), .Z(n5257) );
  XNOR U3820 ( .A(n5259), .B(n5261), .Z(SUM[118]) );
  NANDN U3821 ( .A(n5258), .B(n5260), .Z(n5261) );
  NANDN U3822 ( .A(n5262), .B(n5263), .Z(n5259) );
  NAND U3823 ( .A(n5264), .B(n5265), .Z(n5263) );
  XNOR U3824 ( .A(n5264), .B(n5266), .Z(SUM[117]) );
  NANDN U3825 ( .A(n5262), .B(n5265), .Z(n5266) );
  NANDN U3826 ( .A(n5267), .B(n5268), .Z(n5264) );
  NANDN U3827 ( .A(n5243), .B(n5269), .Z(n5268) );
  XOR U3828 ( .A(n5243), .B(n5270), .Z(SUM[116]) );
  NANDN U3829 ( .A(n5267), .B(n5269), .Z(n5270) );
  ANDN U3830 ( .B(n5271), .A(n5272), .Z(n5243) );
  NANDN U3831 ( .A(n5273), .B(n5274), .Z(n5271) );
  XOR U3832 ( .A(n5275), .B(n5276), .Z(SUM[115]) );
  NANDN U3833 ( .A(n5277), .B(n5278), .Z(n5276) );
  ANDN U3834 ( .B(n5279), .A(n5280), .Z(n5275) );
  NANDN U3835 ( .A(n5281), .B(n5282), .Z(n5279) );
  XNOR U3836 ( .A(n5282), .B(n5283), .Z(SUM[114]) );
  OR U3837 ( .A(n5281), .B(n5280), .Z(n5283) );
  NANDN U3838 ( .A(n5284), .B(n5285), .Z(n5282) );
  NAND U3839 ( .A(n5286), .B(n5287), .Z(n5285) );
  XNOR U3840 ( .A(n5286), .B(n5288), .Z(SUM[113]) );
  NANDN U3841 ( .A(n5284), .B(n5287), .Z(n5288) );
  NANDN U3842 ( .A(n5289), .B(n5290), .Z(n5286) );
  NAND U3843 ( .A(n5274), .B(n5291), .Z(n5290) );
  XNOR U3844 ( .A(n5274), .B(n5292), .Z(SUM[112]) );
  NANDN U3845 ( .A(n5289), .B(n5291), .Z(n5292) );
  NANDN U3846 ( .A(n5293), .B(n5294), .Z(n5274) );
  OR U3847 ( .A(n5295), .B(n125), .Z(n5294) );
  XOR U3848 ( .A(n5296), .B(n5297), .Z(SUM[111]) );
  NANDN U3849 ( .A(n5298), .B(n5299), .Z(n5297) );
  ANDN U3850 ( .B(n5300), .A(n5301), .Z(n5296) );
  NAND U3851 ( .A(n5302), .B(n5303), .Z(n5300) );
  XNOR U3852 ( .A(n5302), .B(n5304), .Z(SUM[110]) );
  NANDN U3853 ( .A(n5301), .B(n5303), .Z(n5304) );
  NANDN U3854 ( .A(n5305), .B(n5306), .Z(n5302) );
  NAND U3855 ( .A(n5307), .B(n5308), .Z(n5306) );
  XNOR U3856 ( .A(n5252), .B(n5309), .Z(SUM[10]) );
  OR U3857 ( .A(n5251), .B(n5250), .Z(n5309) );
  NANDN U3858 ( .A(n3), .B(n5310), .Z(n5252) );
  NANDN U3859 ( .A(n1), .B(n4), .Z(n5310) );
  ANDN U3860 ( .B(n5311), .A(n591), .Z(n1) );
  XNOR U3861 ( .A(n5307), .B(n5312), .Z(SUM[109]) );
  NANDN U3862 ( .A(n5305), .B(n5308), .Z(n5312) );
  NANDN U3863 ( .A(n5313), .B(n5314), .Z(n5307) );
  NAND U3864 ( .A(n5315), .B(n5316), .Z(n5314) );
  XNOR U3865 ( .A(n5315), .B(n5317), .Z(SUM[108]) );
  NANDN U3866 ( .A(n5313), .B(n5316), .Z(n5317) );
  NANDN U3867 ( .A(n5318), .B(n5319), .Z(n5315) );
  NAND U3868 ( .A(n5320), .B(n5321), .Z(n5319) );
  XOR U3869 ( .A(n5322), .B(n5323), .Z(SUM[107]) );
  NANDN U3870 ( .A(n5324), .B(n5325), .Z(n5323) );
  ANDN U3871 ( .B(n5326), .A(n5327), .Z(n5322) );
  NAND U3872 ( .A(n5328), .B(n5329), .Z(n5326) );
  XNOR U3873 ( .A(n5328), .B(n5330), .Z(SUM[106]) );
  NANDN U3874 ( .A(n5327), .B(n5329), .Z(n5330) );
  NANDN U3875 ( .A(n5331), .B(n5332), .Z(n5328) );
  NAND U3876 ( .A(n5333), .B(n5334), .Z(n5332) );
  XNOR U3877 ( .A(n5333), .B(n5335), .Z(SUM[105]) );
  NANDN U3878 ( .A(n5331), .B(n5334), .Z(n5335) );
  NANDN U3879 ( .A(n5336), .B(n5337), .Z(n5333) );
  NAND U3880 ( .A(n5321), .B(n5338), .Z(n5337) );
  XNOR U3881 ( .A(n5321), .B(n5339), .Z(SUM[104]) );
  NANDN U3882 ( .A(n5336), .B(n5338), .Z(n5339) );
  NANDN U3883 ( .A(n5340), .B(n5341), .Z(n5321) );
  OR U3884 ( .A(n5342), .B(n5343), .Z(n5341) );
  XOR U3885 ( .A(n5344), .B(n5345), .Z(SUM[103]) );
  NANDN U3886 ( .A(n5346), .B(n5347), .Z(n5345) );
  ANDN U3887 ( .B(n5348), .A(n5349), .Z(n5344) );
  NAND U3888 ( .A(n5350), .B(n5351), .Z(n5348) );
  XNOR U3889 ( .A(n5350), .B(n5352), .Z(SUM[102]) );
  NANDN U3890 ( .A(n5349), .B(n5351), .Z(n5352) );
  NANDN U3891 ( .A(n5353), .B(n5354), .Z(n5350) );
  NAND U3892 ( .A(n5355), .B(n5356), .Z(n5354) );
  XOR U3893 ( .A(n5357), .B(n5358), .Z(SUM[1021]) );
  XNOR U3894 ( .A(B[1021]), .B(A[1021]), .Z(n5358) );
  ANDN U3895 ( .B(n5359), .A(n5360), .Z(n5357) );
  NAND U3896 ( .A(n5361), .B(n5362), .Z(n5359) );
  XNOR U3897 ( .A(n5361), .B(n5363), .Z(SUM[1020]) );
  NANDN U3898 ( .A(n5360), .B(n5362), .Z(n5363) );
  OR U3899 ( .A(B[1020]), .B(A[1020]), .Z(n5362) );
  AND U3900 ( .A(B[1020]), .B(A[1020]), .Z(n5360) );
  NANDN U3901 ( .A(n5364), .B(n5365), .Z(n5361) );
  NAND U3902 ( .A(n5366), .B(n5367), .Z(n5365) );
  XNOR U3903 ( .A(n5355), .B(n5368), .Z(SUM[101]) );
  NANDN U3904 ( .A(n5353), .B(n5356), .Z(n5368) );
  NANDN U3905 ( .A(n5369), .B(n5370), .Z(n5355) );
  NANDN U3906 ( .A(n5343), .B(n5371), .Z(n5370) );
  XNOR U3907 ( .A(n5366), .B(n5372), .Z(SUM[1019]) );
  NANDN U3908 ( .A(n5364), .B(n5367), .Z(n5372) );
  OR U3909 ( .A(B[1019]), .B(A[1019]), .Z(n5367) );
  AND U3910 ( .A(B[1019]), .B(A[1019]), .Z(n5364) );
  NANDN U3911 ( .A(n5373), .B(n5374), .Z(n5366) );
  NAND U3912 ( .A(n5375), .B(n5376), .Z(n5374) );
  XNOR U3913 ( .A(n5375), .B(n5377), .Z(SUM[1018]) );
  NANDN U3914 ( .A(n5373), .B(n5376), .Z(n5377) );
  OR U3915 ( .A(B[1018]), .B(A[1018]), .Z(n5376) );
  AND U3916 ( .A(B[1018]), .B(A[1018]), .Z(n5373) );
  NANDN U3917 ( .A(n5378), .B(n5379), .Z(n5375) );
  NAND U3918 ( .A(n5380), .B(n5381), .Z(n5379) );
  XNOR U3919 ( .A(n5380), .B(n5382), .Z(SUM[1017]) );
  NANDN U3920 ( .A(n5378), .B(n5381), .Z(n5382) );
  OR U3921 ( .A(B[1017]), .B(A[1017]), .Z(n5381) );
  AND U3922 ( .A(B[1017]), .B(A[1017]), .Z(n5378) );
  NANDN U3923 ( .A(n5383), .B(n5384), .Z(n5380) );
  NAND U3924 ( .A(n5385), .B(n5386), .Z(n5384) );
  XNOR U3925 ( .A(n5385), .B(n5387), .Z(SUM[1016]) );
  NANDN U3926 ( .A(n5383), .B(n5386), .Z(n5387) );
  OR U3927 ( .A(B[1016]), .B(A[1016]), .Z(n5386) );
  AND U3928 ( .A(B[1016]), .B(A[1016]), .Z(n5383) );
  NANDN U3929 ( .A(n5388), .B(n5389), .Z(n5385) );
  NAND U3930 ( .A(n5390), .B(n5391), .Z(n5389) );
  XNOR U3931 ( .A(n5390), .B(n5392), .Z(SUM[1015]) );
  NANDN U3932 ( .A(n5388), .B(n5391), .Z(n5392) );
  OR U3933 ( .A(B[1015]), .B(A[1015]), .Z(n5391) );
  AND U3934 ( .A(B[1015]), .B(A[1015]), .Z(n5388) );
  NANDN U3935 ( .A(n5393), .B(n5394), .Z(n5390) );
  NAND U3936 ( .A(n5395), .B(n5396), .Z(n5394) );
  XNOR U3937 ( .A(n5395), .B(n5397), .Z(SUM[1014]) );
  NANDN U3938 ( .A(n5393), .B(n5396), .Z(n5397) );
  OR U3939 ( .A(B[1014]), .B(A[1014]), .Z(n5396) );
  AND U3940 ( .A(B[1014]), .B(A[1014]), .Z(n5393) );
  NANDN U3941 ( .A(n5398), .B(n5399), .Z(n5395) );
  NAND U3942 ( .A(n5400), .B(n5401), .Z(n5399) );
  XNOR U3943 ( .A(n5400), .B(n5402), .Z(SUM[1013]) );
  NANDN U3944 ( .A(n5398), .B(n5401), .Z(n5402) );
  OR U3945 ( .A(B[1013]), .B(A[1013]), .Z(n5401) );
  AND U3946 ( .A(B[1013]), .B(A[1013]), .Z(n5398) );
  NANDN U3947 ( .A(n5403), .B(n5404), .Z(n5400) );
  NAND U3948 ( .A(n5405), .B(n5406), .Z(n5404) );
  XNOR U3949 ( .A(n5405), .B(n5407), .Z(SUM[1012]) );
  NANDN U3950 ( .A(n5403), .B(n5406), .Z(n5407) );
  OR U3951 ( .A(B[1012]), .B(A[1012]), .Z(n5406) );
  AND U3952 ( .A(B[1012]), .B(A[1012]), .Z(n5403) );
  NANDN U3953 ( .A(n5408), .B(n5409), .Z(n5405) );
  NAND U3954 ( .A(n5410), .B(n5411), .Z(n5409) );
  XNOR U3955 ( .A(n5410), .B(n5412), .Z(SUM[1011]) );
  NANDN U3956 ( .A(n5408), .B(n5411), .Z(n5412) );
  OR U3957 ( .A(B[1011]), .B(A[1011]), .Z(n5411) );
  AND U3958 ( .A(B[1011]), .B(A[1011]), .Z(n5408) );
  NANDN U3959 ( .A(n5413), .B(n5414), .Z(n5410) );
  NAND U3960 ( .A(n5415), .B(n5416), .Z(n5414) );
  XNOR U3961 ( .A(n5415), .B(n5417), .Z(SUM[1010]) );
  NANDN U3962 ( .A(n5413), .B(n5416), .Z(n5417) );
  OR U3963 ( .A(B[1010]), .B(A[1010]), .Z(n5416) );
  AND U3964 ( .A(B[1010]), .B(A[1010]), .Z(n5413) );
  NANDN U3965 ( .A(n5418), .B(n5419), .Z(n5415) );
  NAND U3966 ( .A(n5420), .B(n5421), .Z(n5419) );
  XOR U3967 ( .A(n5343), .B(n5422), .Z(SUM[100]) );
  NANDN U3968 ( .A(n5369), .B(n5371), .Z(n5422) );
  ANDN U3969 ( .B(n5423), .A(n5424), .Z(n5343) );
  OR U3970 ( .A(n5425), .B(n125), .Z(n5423) );
  ANDN U3971 ( .B(n5426), .A(n5427), .Z(n125) );
  OR U3972 ( .A(n890), .B(n5428), .Z(n5426) );
  ANDN U3973 ( .B(n5429), .A(n5430), .Z(n890) );
  XNOR U3974 ( .A(n5420), .B(n5431), .Z(SUM[1009]) );
  NANDN U3975 ( .A(n5418), .B(n5421), .Z(n5431) );
  OR U3976 ( .A(B[1009]), .B(A[1009]), .Z(n5421) );
  AND U3977 ( .A(B[1009]), .B(A[1009]), .Z(n5418) );
  NANDN U3978 ( .A(n5432), .B(n5433), .Z(n5420) );
  NAND U3979 ( .A(n5434), .B(n5435), .Z(n5433) );
  XNOR U3980 ( .A(n5434), .B(n5436), .Z(SUM[1008]) );
  NANDN U3981 ( .A(n5432), .B(n5435), .Z(n5436) );
  OR U3982 ( .A(B[1008]), .B(A[1008]), .Z(n5435) );
  AND U3983 ( .A(B[1008]), .B(A[1008]), .Z(n5432) );
  NANDN U3984 ( .A(n5437), .B(n5438), .Z(n5434) );
  NANDN U3985 ( .A(n5439), .B(n5440), .Z(n5438) );
  NANDN U3986 ( .A(n5441), .B(n5442), .Z(n5440) );
  NANDN U3987 ( .A(n5443), .B(n5444), .Z(n5442) );
  NANDN U3988 ( .A(n5445), .B(n5446), .Z(n5444) );
  NANDN U3989 ( .A(n5447), .B(n5448), .Z(n5446) );
  NANDN U3990 ( .A(n5449), .B(n5450), .Z(n5448) );
  NANDN U3991 ( .A(n5451), .B(n5452), .Z(n5450) );
  NANDN U3992 ( .A(n5453), .B(n5454), .Z(n5452) );
  NANDN U3993 ( .A(n5455), .B(n5456), .Z(n5454) );
  NANDN U3994 ( .A(n5457), .B(n5458), .Z(n5456) );
  AND U3995 ( .A(n5459), .B(n5460), .Z(n5458) );
  OR U3996 ( .A(n5461), .B(n5462), .Z(n5460) );
  OR U3997 ( .A(n5461), .B(n5463), .Z(n5459) );
  XOR U3998 ( .A(n5464), .B(n5465), .Z(SUM[1007]) );
  OR U3999 ( .A(n5439), .B(n5437), .Z(n5465) );
  AND U4000 ( .A(B[1007]), .B(A[1007]), .Z(n5437) );
  NOR U4001 ( .A(B[1007]), .B(A[1007]), .Z(n5439) );
  ANDN U4002 ( .B(n5466), .A(n5441), .Z(n5464) );
  NANDN U4003 ( .A(n5443), .B(n5467), .Z(n5466) );
  XNOR U4004 ( .A(n5467), .B(n5468), .Z(SUM[1006]) );
  OR U4005 ( .A(n5443), .B(n5441), .Z(n5468) );
  AND U4006 ( .A(B[1006]), .B(A[1006]), .Z(n5441) );
  NOR U4007 ( .A(B[1006]), .B(A[1006]), .Z(n5443) );
  NANDN U4008 ( .A(n5445), .B(n5469), .Z(n5467) );
  NANDN U4009 ( .A(n5447), .B(n5470), .Z(n5469) );
  XNOR U4010 ( .A(n5470), .B(n5471), .Z(SUM[1005]) );
  OR U4011 ( .A(n5447), .B(n5445), .Z(n5471) );
  AND U4012 ( .A(B[1005]), .B(A[1005]), .Z(n5445) );
  NOR U4013 ( .A(B[1005]), .B(A[1005]), .Z(n5447) );
  NANDN U4014 ( .A(n5449), .B(n5472), .Z(n5470) );
  NANDN U4015 ( .A(n5451), .B(n5473), .Z(n5472) );
  XNOR U4016 ( .A(n5473), .B(n5474), .Z(SUM[1004]) );
  OR U4017 ( .A(n5451), .B(n5449), .Z(n5474) );
  AND U4018 ( .A(B[1004]), .B(A[1004]), .Z(n5449) );
  NOR U4019 ( .A(B[1004]), .B(A[1004]), .Z(n5451) );
  NANDN U4020 ( .A(n5453), .B(n5475), .Z(n5473) );
  NANDN U4021 ( .A(n5455), .B(n5476), .Z(n5475) );
  NAND U4022 ( .A(n5477), .B(n5478), .Z(n5455) );
  AND U4023 ( .A(n5479), .B(n5480), .Z(n5478) );
  AND U4024 ( .A(n5481), .B(n5482), .Z(n5477) );
  NANDN U4025 ( .A(n5483), .B(n5484), .Z(n5453) );
  NAND U4026 ( .A(n5485), .B(n5482), .Z(n5484) );
  NANDN U4027 ( .A(n5486), .B(n5487), .Z(n5485) );
  NAND U4028 ( .A(n5488), .B(n5481), .Z(n5487) );
  NANDN U4029 ( .A(n5489), .B(n5490), .Z(n5488) );
  NAND U4030 ( .A(n5480), .B(n5491), .Z(n5490) );
  XOR U4031 ( .A(n5492), .B(n5493), .Z(SUM[1003]) );
  NANDN U4032 ( .A(n5483), .B(n5482), .Z(n5493) );
  OR U4033 ( .A(B[1003]), .B(A[1003]), .Z(n5482) );
  AND U4034 ( .A(B[1003]), .B(A[1003]), .Z(n5483) );
  ANDN U4035 ( .B(n5494), .A(n5486), .Z(n5492) );
  NAND U4036 ( .A(n5495), .B(n5481), .Z(n5494) );
  XNOR U4037 ( .A(n5495), .B(n5496), .Z(SUM[1002]) );
  NANDN U4038 ( .A(n5486), .B(n5481), .Z(n5496) );
  OR U4039 ( .A(B[1002]), .B(A[1002]), .Z(n5481) );
  AND U4040 ( .A(B[1002]), .B(A[1002]), .Z(n5486) );
  NANDN U4041 ( .A(n5489), .B(n5497), .Z(n5495) );
  NAND U4042 ( .A(n5498), .B(n5480), .Z(n5497) );
  XNOR U4043 ( .A(n5498), .B(n5499), .Z(SUM[1001]) );
  NANDN U4044 ( .A(n5489), .B(n5480), .Z(n5499) );
  OR U4045 ( .A(B[1001]), .B(A[1001]), .Z(n5480) );
  AND U4046 ( .A(B[1001]), .B(A[1001]), .Z(n5489) );
  NANDN U4047 ( .A(n5491), .B(n5500), .Z(n5498) );
  NAND U4048 ( .A(n5476), .B(n5479), .Z(n5500) );
  XNOR U4049 ( .A(n5476), .B(n5501), .Z(SUM[1000]) );
  NANDN U4050 ( .A(n5491), .B(n5479), .Z(n5501) );
  OR U4051 ( .A(B[1000]), .B(A[1000]), .Z(n5479) );
  AND U4052 ( .A(B[1000]), .B(A[1000]), .Z(n5491) );
  NANDN U4053 ( .A(n5457), .B(n5502), .Z(n5476) );
  OR U4054 ( .A(n5461), .B(n29), .Z(n5502) );
  AND U4055 ( .A(n5463), .B(n5462), .Z(n29) );
  ANDN U4056 ( .B(n5503), .A(n34), .Z(n5462) );
  AND U4057 ( .A(B[995]), .B(A[995]), .Z(n34) );
  NAND U4058 ( .A(n5504), .B(n35), .Z(n5503) );
  NANDN U4059 ( .A(n37), .B(n5505), .Z(n5504) );
  NAND U4060 ( .A(n5506), .B(n39), .Z(n5505) );
  NANDN U4061 ( .A(n41), .B(n5507), .Z(n5506) );
  NAND U4062 ( .A(n44), .B(n46), .Z(n5507) );
  AND U4063 ( .A(B[992]), .B(A[992]), .Z(n46) );
  AND U4064 ( .A(B[993]), .B(A[993]), .Z(n41) );
  AND U4065 ( .A(B[994]), .B(A[994]), .Z(n37) );
  NAND U4066 ( .A(n5508), .B(n5509), .Z(n5463) );
  AND U4067 ( .A(n44), .B(n5510), .Z(n5509) );
  AND U4068 ( .A(n35), .B(n39), .Z(n5510) );
  OR U4069 ( .A(B[994]), .B(A[994]), .Z(n39) );
  OR U4070 ( .A(B[995]), .B(A[995]), .Z(n35) );
  OR U4071 ( .A(B[993]), .B(A[993]), .Z(n44) );
  NOR U4072 ( .A(n48), .B(n49), .Z(n5508) );
  NOR U4073 ( .A(B[992]), .B(A[992]), .Z(n49) );
  ANDN U4074 ( .B(n5511), .A(n54), .Z(n48) );
  AND U4075 ( .A(B[991]), .B(A[991]), .Z(n54) );
  NANDN U4076 ( .A(n53), .B(n5512), .Z(n5511) );
  NANDN U4077 ( .A(n56), .B(n5513), .Z(n5512) );
  NANDN U4078 ( .A(n57), .B(n5514), .Z(n5513) );
  NANDN U4079 ( .A(n60), .B(n5515), .Z(n5514) );
  NANDN U4080 ( .A(n62), .B(n5516), .Z(n5515) );
  NANDN U4081 ( .A(n70), .B(n5517), .Z(n5516) );
  NANDN U4082 ( .A(n72), .B(n5518), .Z(n5517) );
  NANDN U4083 ( .A(n75), .B(n5519), .Z(n5518) );
  NANDN U4084 ( .A(n77), .B(n5520), .Z(n5519) );
  NANDN U4085 ( .A(n97), .B(n5521), .Z(n5520) );
  AND U4086 ( .A(n5522), .B(n5523), .Z(n5521) );
  NANDN U4087 ( .A(n99), .B(n119), .Z(n5523) );
  NANDN U4088 ( .A(n128), .B(n5524), .Z(n119) );
  NAND U4089 ( .A(n5525), .B(n129), .Z(n5524) );
  NANDN U4090 ( .A(n131), .B(n5526), .Z(n5525) );
  NAND U4091 ( .A(n5527), .B(n133), .Z(n5526) );
  NANDN U4092 ( .A(n135), .B(n5528), .Z(n5527) );
  NAND U4093 ( .A(n138), .B(n140), .Z(n5528) );
  AND U4094 ( .A(A[976]), .B(B[976]), .Z(n140) );
  AND U4095 ( .A(A[977]), .B(B[977]), .Z(n135) );
  AND U4096 ( .A(A[978]), .B(B[978]), .Z(n131) );
  AND U4097 ( .A(B[979]), .B(A[979]), .Z(n128) );
  NANDN U4098 ( .A(n99), .B(n120), .Z(n5522) );
  AND U4099 ( .A(n5529), .B(n5530), .Z(n120) );
  AND U4100 ( .A(n138), .B(n5531), .Z(n5530) );
  NOR U4101 ( .A(n142), .B(n143), .Z(n5531) );
  NOR U4102 ( .A(B[976]), .B(A[976]), .Z(n143) );
  ANDN U4103 ( .B(n5532), .A(n148), .Z(n142) );
  AND U4104 ( .A(B[975]), .B(A[975]), .Z(n148) );
  NANDN U4105 ( .A(n147), .B(n5533), .Z(n5532) );
  NANDN U4106 ( .A(n150), .B(n5534), .Z(n5533) );
  NANDN U4107 ( .A(n151), .B(n5535), .Z(n5534) );
  NANDN U4108 ( .A(n154), .B(n5536), .Z(n5535) );
  NANDN U4109 ( .A(n156), .B(n5537), .Z(n5536) );
  NANDN U4110 ( .A(n159), .B(n5538), .Z(n5537) );
  NANDN U4111 ( .A(n161), .B(n5539), .Z(n5538) );
  NANDN U4112 ( .A(n164), .B(n5540), .Z(n5539) );
  NANDN U4113 ( .A(n166), .B(n5541), .Z(n5540) );
  NANDN U4114 ( .A(n187), .B(n5542), .Z(n5541) );
  AND U4115 ( .A(n5543), .B(n5544), .Z(n5542) );
  NANDN U4116 ( .A(n189), .B(n209), .Z(n5544) );
  NANDN U4117 ( .A(n213), .B(n5545), .Z(n209) );
  NAND U4118 ( .A(n5546), .B(n214), .Z(n5545) );
  NANDN U4119 ( .A(n216), .B(n5547), .Z(n5546) );
  NAND U4120 ( .A(n5548), .B(n218), .Z(n5547) );
  NANDN U4121 ( .A(n220), .B(n5549), .Z(n5548) );
  NAND U4122 ( .A(n223), .B(n225), .Z(n5549) );
  AND U4123 ( .A(A[960]), .B(B[960]), .Z(n225) );
  AND U4124 ( .A(A[961]), .B(B[961]), .Z(n220) );
  AND U4125 ( .A(A[962]), .B(B[962]), .Z(n216) );
  AND U4126 ( .A(B[963]), .B(A[963]), .Z(n213) );
  NANDN U4127 ( .A(n189), .B(n210), .Z(n5543) );
  AND U4128 ( .A(n5550), .B(n5551), .Z(n210) );
  AND U4129 ( .A(n223), .B(n5552), .Z(n5551) );
  NOR U4130 ( .A(n227), .B(n228), .Z(n5552) );
  NOR U4131 ( .A(B[960]), .B(A[960]), .Z(n228) );
  ANDN U4132 ( .B(n5553), .A(n241), .Z(n227) );
  AND U4133 ( .A(B[959]), .B(A[959]), .Z(n241) );
  NANDN U4134 ( .A(n240), .B(n5554), .Z(n5553) );
  NANDN U4135 ( .A(n243), .B(n5555), .Z(n5554) );
  NANDN U4136 ( .A(n244), .B(n5556), .Z(n5555) );
  NANDN U4137 ( .A(n247), .B(n5557), .Z(n5556) );
  NANDN U4138 ( .A(n249), .B(n5558), .Z(n5557) );
  NAND U4139 ( .A(n5559), .B(n5560), .Z(n5558) );
  NAND U4140 ( .A(n5561), .B(n5562), .Z(n5560) );
  AND U4141 ( .A(n282), .B(n5563), .Z(n5562) );
  ANDN U4142 ( .B(n255), .A(n309), .Z(n5563) );
  ANDN U4143 ( .B(n5564), .A(n331), .Z(n309) );
  AND U4144 ( .A(B[943]), .B(A[943]), .Z(n331) );
  NANDN U4145 ( .A(n330), .B(n5565), .Z(n5564) );
  NANDN U4146 ( .A(n333), .B(n5566), .Z(n5565) );
  NANDN U4147 ( .A(n334), .B(n5567), .Z(n5566) );
  NANDN U4148 ( .A(n337), .B(n5568), .Z(n5567) );
  NANDN U4149 ( .A(n339), .B(n5569), .Z(n5568) );
  NAND U4150 ( .A(n5570), .B(n5571), .Z(n5569) );
  NAND U4151 ( .A(n5572), .B(n5573), .Z(n5571) );
  AND U4152 ( .A(n377), .B(n5574), .Z(n5573) );
  ANDN U4153 ( .B(n345), .A(n399), .Z(n5574) );
  ANDN U4154 ( .B(n5575), .A(n426), .Z(n399) );
  AND U4155 ( .A(B[927]), .B(A[927]), .Z(n426) );
  NANDN U4156 ( .A(n425), .B(n5576), .Z(n5575) );
  NANDN U4157 ( .A(n428), .B(n5577), .Z(n5576) );
  NANDN U4158 ( .A(n429), .B(n5578), .Z(n5577) );
  NANDN U4159 ( .A(n432), .B(n5579), .Z(n5578) );
  NANDN U4160 ( .A(n434), .B(n5580), .Z(n5579) );
  NAND U4161 ( .A(n5581), .B(n5582), .Z(n5580) );
  NAND U4162 ( .A(n5583), .B(n5584), .Z(n5582) );
  AND U4163 ( .A(n467), .B(n5585), .Z(n5584) );
  ANDN U4164 ( .B(n440), .A(n497), .Z(n5585) );
  ANDN U4165 ( .B(n5586), .A(n519), .Z(n497) );
  AND U4166 ( .A(B[911]), .B(A[911]), .Z(n519) );
  NANDN U4167 ( .A(n518), .B(n5587), .Z(n5586) );
  NANDN U4168 ( .A(n521), .B(n5588), .Z(n5587) );
  NANDN U4169 ( .A(n522), .B(n5589), .Z(n5588) );
  NANDN U4170 ( .A(n525), .B(n5590), .Z(n5589) );
  NANDN U4171 ( .A(n527), .B(n5591), .Z(n5590) );
  NAND U4172 ( .A(n5592), .B(n5593), .Z(n5591) );
  NAND U4173 ( .A(n5594), .B(n5595), .Z(n5593) );
  AND U4174 ( .A(n565), .B(n5596), .Z(n5595) );
  ANDN U4175 ( .B(n538), .A(n587), .Z(n5596) );
  ANDN U4176 ( .B(n5597), .A(n617), .Z(n587) );
  AND U4177 ( .A(B[895]), .B(A[895]), .Z(n617) );
  NANDN U4178 ( .A(n616), .B(n5598), .Z(n5597) );
  NANDN U4179 ( .A(n619), .B(n5599), .Z(n5598) );
  NANDN U4180 ( .A(n620), .B(n5600), .Z(n5599) );
  NANDN U4181 ( .A(n623), .B(n5601), .Z(n5600) );
  NANDN U4182 ( .A(n625), .B(n5602), .Z(n5601) );
  NAND U4183 ( .A(n5603), .B(n5604), .Z(n5602) );
  NAND U4184 ( .A(n5605), .B(n5606), .Z(n5604) );
  AND U4185 ( .A(n663), .B(n5607), .Z(n5606) );
  ANDN U4186 ( .B(n631), .A(n685), .Z(n5607) );
  ANDN U4187 ( .B(n5608), .A(n715), .Z(n685) );
  AND U4188 ( .A(B[879]), .B(A[879]), .Z(n715) );
  NANDN U4189 ( .A(n714), .B(n5609), .Z(n5608) );
  NANDN U4190 ( .A(n717), .B(n5610), .Z(n5609) );
  NANDN U4191 ( .A(n718), .B(n5611), .Z(n5610) );
  NANDN U4192 ( .A(n721), .B(n5612), .Z(n5611) );
  NANDN U4193 ( .A(n723), .B(n5613), .Z(n5612) );
  NAND U4194 ( .A(n5614), .B(n5615), .Z(n5613) );
  NAND U4195 ( .A(n5616), .B(n5617), .Z(n5615) );
  AND U4196 ( .A(n756), .B(n5618), .Z(n5617) );
  ANDN U4197 ( .B(n729), .A(n783), .Z(n5618) );
  ANDN U4198 ( .B(n5619), .A(n805), .Z(n783) );
  AND U4199 ( .A(B[863]), .B(A[863]), .Z(n805) );
  NANDN U4200 ( .A(n804), .B(n5620), .Z(n5619) );
  NANDN U4201 ( .A(n807), .B(n5621), .Z(n5620) );
  NANDN U4202 ( .A(n808), .B(n5622), .Z(n5621) );
  NANDN U4203 ( .A(n811), .B(n5623), .Z(n5622) );
  NANDN U4204 ( .A(n813), .B(n5624), .Z(n5623) );
  NAND U4205 ( .A(n5625), .B(n5626), .Z(n5624) );
  NAND U4206 ( .A(n5627), .B(n5628), .Z(n5626) );
  AND U4207 ( .A(n850), .B(n5629), .Z(n5628) );
  ANDN U4208 ( .B(n819), .A(n872), .Z(n5629) );
  ANDN U4209 ( .B(n5630), .A(n899), .Z(n872) );
  AND U4210 ( .A(B[847]), .B(A[847]), .Z(n899) );
  NANDN U4211 ( .A(n898), .B(n5631), .Z(n5630) );
  NANDN U4212 ( .A(n901), .B(n5632), .Z(n5631) );
  NANDN U4213 ( .A(n902), .B(n5633), .Z(n5632) );
  NANDN U4214 ( .A(n905), .B(n5634), .Z(n5633) );
  NANDN U4215 ( .A(n907), .B(n5635), .Z(n5634) );
  NAND U4216 ( .A(n5636), .B(n5637), .Z(n5635) );
  NAND U4217 ( .A(n5638), .B(n5639), .Z(n5637) );
  AND U4218 ( .A(n940), .B(n5640), .Z(n5639) );
  ANDN U4219 ( .B(n913), .A(n970), .Z(n5640) );
  ANDN U4220 ( .B(n5641), .A(n992), .Z(n970) );
  AND U4221 ( .A(B[831]), .B(A[831]), .Z(n992) );
  NANDN U4222 ( .A(n991), .B(n5642), .Z(n5641) );
  NANDN U4223 ( .A(n994), .B(n5643), .Z(n5642) );
  NANDN U4224 ( .A(n995), .B(n5644), .Z(n5643) );
  NANDN U4225 ( .A(n998), .B(n5645), .Z(n5644) );
  NANDN U4226 ( .A(n1000), .B(n5646), .Z(n5645) );
  NAND U4227 ( .A(n5647), .B(n5648), .Z(n5646) );
  NAND U4228 ( .A(n5649), .B(n5650), .Z(n5648) );
  AND U4229 ( .A(n1038), .B(n5651), .Z(n5650) );
  ANDN U4230 ( .B(n1011), .A(n1060), .Z(n5651) );
  ANDN U4231 ( .B(n5652), .A(n1086), .Z(n1060) );
  AND U4232 ( .A(B[815]), .B(A[815]), .Z(n1086) );
  NANDN U4233 ( .A(n1085), .B(n5653), .Z(n5652) );
  NANDN U4234 ( .A(n1088), .B(n5654), .Z(n5653) );
  NANDN U4235 ( .A(n1089), .B(n5655), .Z(n5654) );
  NANDN U4236 ( .A(n1092), .B(n5656), .Z(n5655) );
  NANDN U4237 ( .A(n1094), .B(n5657), .Z(n5656) );
  NAND U4238 ( .A(n5658), .B(n5659), .Z(n5657) );
  NAND U4239 ( .A(n5660), .B(n5661), .Z(n5659) );
  AND U4240 ( .A(n1128), .B(n5662), .Z(n5661) );
  ANDN U4241 ( .B(n1100), .A(n1150), .Z(n5662) );
  ANDN U4242 ( .B(n5663), .A(n1186), .Z(n1150) );
  AND U4243 ( .A(B[799]), .B(A[799]), .Z(n1186) );
  NANDN U4244 ( .A(n1185), .B(n5664), .Z(n5663) );
  NANDN U4245 ( .A(n1188), .B(n5665), .Z(n5664) );
  NANDN U4246 ( .A(n1189), .B(n5666), .Z(n5665) );
  NANDN U4247 ( .A(n1192), .B(n5667), .Z(n5666) );
  NANDN U4248 ( .A(n1194), .B(n5668), .Z(n5667) );
  NAND U4249 ( .A(n5669), .B(n5670), .Z(n5668) );
  NAND U4250 ( .A(n5671), .B(n5672), .Z(n5670) );
  AND U4251 ( .A(n1227), .B(n5673), .Z(n5672) );
  ANDN U4252 ( .B(n1200), .A(n1254), .Z(n5673) );
  ANDN U4253 ( .B(n5674), .A(n1276), .Z(n1254) );
  AND U4254 ( .A(B[783]), .B(A[783]), .Z(n1276) );
  NANDN U4255 ( .A(n1275), .B(n5675), .Z(n5674) );
  NANDN U4256 ( .A(n1278), .B(n5676), .Z(n5675) );
  NANDN U4257 ( .A(n1279), .B(n5677), .Z(n5676) );
  NANDN U4258 ( .A(n1282), .B(n5678), .Z(n5677) );
  NANDN U4259 ( .A(n1284), .B(n5679), .Z(n5678) );
  NAND U4260 ( .A(n5680), .B(n5681), .Z(n5679) );
  NAND U4261 ( .A(n5682), .B(n5683), .Z(n5681) );
  AND U4262 ( .A(n1322), .B(n5684), .Z(n5683) );
  ANDN U4263 ( .B(n1290), .A(n1344), .Z(n5684) );
  ANDN U4264 ( .B(n5685), .A(n1371), .Z(n1344) );
  AND U4265 ( .A(B[767]), .B(A[767]), .Z(n1371) );
  NANDN U4266 ( .A(n1370), .B(n5686), .Z(n5685) );
  NAND U4267 ( .A(n5687), .B(n5688), .Z(n5686) );
  NAND U4268 ( .A(n5689), .B(n5690), .Z(n5688) );
  AND U4269 ( .A(n5691), .B(n5692), .Z(n5690) );
  ANDN U4270 ( .B(n1380), .A(n1384), .Z(n5692) );
  AND U4271 ( .A(n1375), .B(n5693), .Z(n5691) );
  NANDN U4272 ( .A(n1461), .B(n5694), .Z(n5693) );
  NANDN U4273 ( .A(n1463), .B(n5695), .Z(n5694) );
  NANDN U4274 ( .A(n1558), .B(n5696), .Z(n5695) );
  NANDN U4275 ( .A(n1560), .B(n5697), .Z(n5696) );
  NANDN U4276 ( .A(n1651), .B(n5698), .Z(n5697) );
  NANDN U4277 ( .A(n1653), .B(n5699), .Z(n5698) );
  NANDN U4278 ( .A(n1752), .B(n5700), .Z(n5699) );
  NANDN U4279 ( .A(n1754), .B(n5701), .Z(n5700) );
  NANDN U4280 ( .A(n2134), .B(n5702), .Z(n5701) );
  AND U4281 ( .A(n5703), .B(n5704), .Z(n5702) );
  NANDN U4282 ( .A(n2136), .B(n2530), .Z(n5704) );
  NAND U4283 ( .A(n5705), .B(n5706), .Z(n2530) );
  NAND U4284 ( .A(n5707), .B(n2535), .Z(n5706) );
  NANDN U4285 ( .A(n2537), .B(n5708), .Z(n5707) );
  NAND U4286 ( .A(n5709), .B(n2539), .Z(n5708) );
  NANDN U4287 ( .A(n2541), .B(n5710), .Z(n5709) );
  NAND U4288 ( .A(n5711), .B(n2544), .Z(n5710) );
  NANDN U4289 ( .A(n2546), .B(n5712), .Z(n5711) );
  NAND U4290 ( .A(n5713), .B(n2549), .Z(n5712) );
  NANDN U4291 ( .A(n2551), .B(n5714), .Z(n5713) );
  NANDN U4292 ( .A(n2553), .B(n5715), .Z(n5714) );
  NANDN U4293 ( .A(n2578), .B(n5716), .Z(n5715) );
  NANDN U4294 ( .A(n2580), .B(n2601), .Z(n5716) );
  NANDN U4295 ( .A(n2606), .B(n5717), .Z(n2601) );
  NAND U4296 ( .A(n5718), .B(n2607), .Z(n5717) );
  NANDN U4297 ( .A(n2609), .B(n5719), .Z(n5718) );
  NAND U4298 ( .A(n5720), .B(n2611), .Z(n5719) );
  NANDN U4299 ( .A(n2613), .B(n5721), .Z(n5720) );
  NAND U4300 ( .A(n2616), .B(n2618), .Z(n5721) );
  AND U4301 ( .A(A[560]), .B(B[560]), .Z(n2618) );
  AND U4302 ( .A(A[561]), .B(B[561]), .Z(n2613) );
  AND U4303 ( .A(A[562]), .B(B[562]), .Z(n2609) );
  AND U4304 ( .A(B[563]), .B(A[563]), .Z(n2606) );
  NANDN U4305 ( .A(n2584), .B(n5722), .Z(n2578) );
  NAND U4306 ( .A(n5723), .B(n2585), .Z(n5722) );
  NANDN U4307 ( .A(n2587), .B(n5724), .Z(n5723) );
  NAND U4308 ( .A(n5725), .B(n2589), .Z(n5724) );
  NANDN U4309 ( .A(n2591), .B(n5726), .Z(n5725) );
  NAND U4310 ( .A(n2594), .B(n2596), .Z(n5726) );
  AND U4311 ( .A(A[564]), .B(B[564]), .Z(n2596) );
  AND U4312 ( .A(A[565]), .B(B[565]), .Z(n2591) );
  AND U4313 ( .A(A[566]), .B(B[566]), .Z(n2587) );
  AND U4314 ( .A(B[567]), .B(A[567]), .Z(n2584) );
  NANDN U4315 ( .A(n2557), .B(n5727), .Z(n2551) );
  NAND U4316 ( .A(n5728), .B(n2558), .Z(n5727) );
  NANDN U4317 ( .A(n2560), .B(n5729), .Z(n5728) );
  NAND U4318 ( .A(n5730), .B(n2562), .Z(n5729) );
  NANDN U4319 ( .A(n2564), .B(n5731), .Z(n5730) );
  NAND U4320 ( .A(n2567), .B(n2574), .Z(n5731) );
  AND U4321 ( .A(A[568]), .B(B[568]), .Z(n2574) );
  AND U4322 ( .A(A[569]), .B(B[569]), .Z(n2564) );
  AND U4323 ( .A(A[570]), .B(B[570]), .Z(n2560) );
  AND U4324 ( .A(B[571]), .B(A[571]), .Z(n2557) );
  AND U4325 ( .A(A[572]), .B(B[572]), .Z(n2546) );
  AND U4326 ( .A(A[573]), .B(B[573]), .Z(n2541) );
  AND U4327 ( .A(A[574]), .B(B[574]), .Z(n2537) );
  ANDN U4328 ( .B(n5732), .A(n2534), .Z(n5705) );
  AND U4329 ( .A(B[575]), .B(A[575]), .Z(n2534) );
  NANDN U4330 ( .A(n5733), .B(n5734), .Z(n5732) );
  NANDN U4331 ( .A(n2622), .B(n5735), .Z(n5734) );
  NANDN U4332 ( .A(n2624), .B(n5736), .Z(n5735) );
  NANDN U4333 ( .A(n2723), .B(n5737), .Z(n5736) );
  NANDN U4334 ( .A(n2725), .B(n2819), .Z(n5737) );
  NANDN U4335 ( .A(n2824), .B(n5738), .Z(n2819) );
  NAND U4336 ( .A(n5739), .B(n2825), .Z(n5738) );
  NANDN U4337 ( .A(n2827), .B(n5740), .Z(n5739) );
  NAND U4338 ( .A(n5741), .B(n2829), .Z(n5740) );
  NANDN U4339 ( .A(n2831), .B(n5742), .Z(n5741) );
  NAND U4340 ( .A(n5743), .B(n2834), .Z(n5742) );
  NANDN U4341 ( .A(n2836), .B(n5744), .Z(n5743) );
  NAND U4342 ( .A(n5745), .B(n2839), .Z(n5744) );
  NANDN U4343 ( .A(n2841), .B(n5746), .Z(n5745) );
  NANDN U4344 ( .A(n2843), .B(n5747), .Z(n5746) );
  NANDN U4345 ( .A(n2863), .B(n5748), .Z(n5747) );
  NANDN U4346 ( .A(n2865), .B(n2894), .Z(n5748) );
  NANDN U4347 ( .A(n2898), .B(n5749), .Z(n2894) );
  NAND U4348 ( .A(n5750), .B(n2899), .Z(n5749) );
  NANDN U4349 ( .A(n2901), .B(n5751), .Z(n5750) );
  NAND U4350 ( .A(n5752), .B(n2903), .Z(n5751) );
  NANDN U4351 ( .A(n2905), .B(n5753), .Z(n5752) );
  NAND U4352 ( .A(n2908), .B(n2910), .Z(n5753) );
  AND U4353 ( .A(A[512]), .B(B[512]), .Z(n2910) );
  AND U4354 ( .A(A[513]), .B(B[513]), .Z(n2905) );
  AND U4355 ( .A(A[514]), .B(B[514]), .Z(n2901) );
  AND U4356 ( .A(B[515]), .B(A[515]), .Z(n2898) );
  NANDN U4357 ( .A(n2877), .B(n5754), .Z(n2863) );
  NAND U4358 ( .A(n5755), .B(n2878), .Z(n5754) );
  NANDN U4359 ( .A(n2880), .B(n5756), .Z(n5755) );
  NAND U4360 ( .A(n5757), .B(n2882), .Z(n5756) );
  NANDN U4361 ( .A(n2884), .B(n5758), .Z(n5757) );
  NAND U4362 ( .A(n2887), .B(n2889), .Z(n5758) );
  AND U4363 ( .A(A[516]), .B(B[516]), .Z(n2889) );
  AND U4364 ( .A(A[517]), .B(B[517]), .Z(n2884) );
  AND U4365 ( .A(A[518]), .B(B[518]), .Z(n2880) );
  AND U4366 ( .A(B[519]), .B(A[519]), .Z(n2877) );
  NANDN U4367 ( .A(n2847), .B(n5759), .Z(n2841) );
  NAND U4368 ( .A(n5760), .B(n2848), .Z(n5759) );
  NANDN U4369 ( .A(n2850), .B(n5761), .Z(n5760) );
  NAND U4370 ( .A(n5762), .B(n2852), .Z(n5761) );
  NANDN U4371 ( .A(n2854), .B(n5763), .Z(n5762) );
  NAND U4372 ( .A(n2857), .B(n2859), .Z(n5763) );
  AND U4373 ( .A(A[520]), .B(B[520]), .Z(n2859) );
  AND U4374 ( .A(A[521]), .B(B[521]), .Z(n2854) );
  AND U4375 ( .A(A[522]), .B(B[522]), .Z(n2850) );
  AND U4376 ( .A(B[523]), .B(A[523]), .Z(n2847) );
  AND U4377 ( .A(A[524]), .B(B[524]), .Z(n2836) );
  AND U4378 ( .A(A[525]), .B(B[525]), .Z(n2831) );
  AND U4379 ( .A(A[526]), .B(B[526]), .Z(n2827) );
  AND U4380 ( .A(B[527]), .B(A[527]), .Z(n2824) );
  NANDN U4381 ( .A(n2729), .B(n5764), .Z(n2723) );
  NAND U4382 ( .A(n5765), .B(n2730), .Z(n5764) );
  NANDN U4383 ( .A(n2732), .B(n5766), .Z(n5765) );
  NAND U4384 ( .A(n5767), .B(n2734), .Z(n5766) );
  NANDN U4385 ( .A(n2736), .B(n5768), .Z(n5767) );
  NAND U4386 ( .A(n5769), .B(n2739), .Z(n5768) );
  NANDN U4387 ( .A(n2741), .B(n5770), .Z(n5769) );
  NAND U4388 ( .A(n5771), .B(n2744), .Z(n5770) );
  NANDN U4389 ( .A(n2746), .B(n5772), .Z(n5771) );
  NANDN U4390 ( .A(n2748), .B(n5773), .Z(n5772) );
  NANDN U4391 ( .A(n2772), .B(n5774), .Z(n5773) );
  NANDN U4392 ( .A(n2774), .B(n2795), .Z(n5774) );
  NANDN U4393 ( .A(n2799), .B(n5775), .Z(n2795) );
  NAND U4394 ( .A(n5776), .B(n2800), .Z(n5775) );
  NANDN U4395 ( .A(n2802), .B(n5777), .Z(n5776) );
  NAND U4396 ( .A(n5778), .B(n2804), .Z(n5777) );
  NANDN U4397 ( .A(n2806), .B(n5779), .Z(n5778) );
  NAND U4398 ( .A(n2809), .B(n2814), .Z(n5779) );
  AND U4399 ( .A(A[528]), .B(B[528]), .Z(n2814) );
  AND U4400 ( .A(A[529]), .B(B[529]), .Z(n2806) );
  AND U4401 ( .A(A[530]), .B(B[530]), .Z(n2802) );
  AND U4402 ( .A(B[531]), .B(A[531]), .Z(n2799) );
  NANDN U4403 ( .A(n2778), .B(n5780), .Z(n2772) );
  NAND U4404 ( .A(n5781), .B(n2779), .Z(n5780) );
  NANDN U4405 ( .A(n2781), .B(n5782), .Z(n5781) );
  NAND U4406 ( .A(n5783), .B(n2783), .Z(n5782) );
  NANDN U4407 ( .A(n2785), .B(n5784), .Z(n5783) );
  NAND U4408 ( .A(n2788), .B(n2790), .Z(n5784) );
  AND U4409 ( .A(A[532]), .B(B[532]), .Z(n2790) );
  AND U4410 ( .A(A[533]), .B(B[533]), .Z(n2785) );
  AND U4411 ( .A(A[534]), .B(B[534]), .Z(n2781) );
  AND U4412 ( .A(B[535]), .B(A[535]), .Z(n2778) );
  NANDN U4413 ( .A(n2756), .B(n5785), .Z(n2746) );
  NAND U4414 ( .A(n5786), .B(n2757), .Z(n5785) );
  NANDN U4415 ( .A(n2759), .B(n5787), .Z(n5786) );
  NAND U4416 ( .A(n5788), .B(n2761), .Z(n5787) );
  NANDN U4417 ( .A(n2763), .B(n5789), .Z(n5788) );
  NAND U4418 ( .A(n2766), .B(n2768), .Z(n5789) );
  AND U4419 ( .A(A[536]), .B(B[536]), .Z(n2768) );
  AND U4420 ( .A(A[537]), .B(B[537]), .Z(n2763) );
  AND U4421 ( .A(A[538]), .B(B[538]), .Z(n2759) );
  AND U4422 ( .A(B[539]), .B(A[539]), .Z(n2756) );
  AND U4423 ( .A(A[540]), .B(B[540]), .Z(n2741) );
  AND U4424 ( .A(A[541]), .B(B[541]), .Z(n2736) );
  AND U4425 ( .A(A[542]), .B(B[542]), .Z(n2732) );
  AND U4426 ( .A(B[543]), .B(A[543]), .Z(n2729) );
  NANDN U4427 ( .A(n2636), .B(n5790), .Z(n2622) );
  NAND U4428 ( .A(n5791), .B(n2637), .Z(n5790) );
  NANDN U4429 ( .A(n2639), .B(n5792), .Z(n5791) );
  NAND U4430 ( .A(n5793), .B(n2641), .Z(n5792) );
  NANDN U4431 ( .A(n2643), .B(n5794), .Z(n5793) );
  NAND U4432 ( .A(n5795), .B(n2646), .Z(n5794) );
  NANDN U4433 ( .A(n2648), .B(n5796), .Z(n5795) );
  NAND U4434 ( .A(n5797), .B(n2651), .Z(n5796) );
  NANDN U4435 ( .A(n2653), .B(n5798), .Z(n5797) );
  NANDN U4436 ( .A(n2655), .B(n5799), .Z(n5798) );
  NANDN U4437 ( .A(n2675), .B(n5800), .Z(n5799) );
  NANDN U4438 ( .A(n2677), .B(n2703), .Z(n5800) );
  NANDN U4439 ( .A(n2707), .B(n5801), .Z(n2703) );
  NAND U4440 ( .A(n5802), .B(n2708), .Z(n5801) );
  NANDN U4441 ( .A(n2710), .B(n5803), .Z(n5802) );
  NAND U4442 ( .A(n5804), .B(n2712), .Z(n5803) );
  NANDN U4443 ( .A(n2714), .B(n5805), .Z(n5804) );
  NAND U4444 ( .A(n2717), .B(n2719), .Z(n5805) );
  AND U4445 ( .A(A[544]), .B(B[544]), .Z(n2719) );
  AND U4446 ( .A(A[545]), .B(B[545]), .Z(n2714) );
  AND U4447 ( .A(A[546]), .B(B[546]), .Z(n2710) );
  AND U4448 ( .A(B[547]), .B(A[547]), .Z(n2707) );
  NANDN U4449 ( .A(n2681), .B(n5806), .Z(n2675) );
  NAND U4450 ( .A(n5807), .B(n2682), .Z(n5806) );
  NANDN U4451 ( .A(n2684), .B(n5808), .Z(n5807) );
  NAND U4452 ( .A(n5809), .B(n2686), .Z(n5808) );
  NANDN U4453 ( .A(n2688), .B(n5810), .Z(n5809) );
  NAND U4454 ( .A(n2691), .B(n2698), .Z(n5810) );
  AND U4455 ( .A(A[548]), .B(B[548]), .Z(n2698) );
  AND U4456 ( .A(A[549]), .B(B[549]), .Z(n2688) );
  AND U4457 ( .A(A[550]), .B(B[550]), .Z(n2684) );
  AND U4458 ( .A(B[551]), .B(A[551]), .Z(n2681) );
  NANDN U4459 ( .A(n2659), .B(n5811), .Z(n2653) );
  NAND U4460 ( .A(n5812), .B(n2660), .Z(n5811) );
  NANDN U4461 ( .A(n2662), .B(n5813), .Z(n5812) );
  NAND U4462 ( .A(n5814), .B(n2664), .Z(n5813) );
  NANDN U4463 ( .A(n2666), .B(n5815), .Z(n5814) );
  NAND U4464 ( .A(n2669), .B(n2671), .Z(n5815) );
  AND U4465 ( .A(A[552]), .B(B[552]), .Z(n2671) );
  AND U4466 ( .A(A[553]), .B(B[553]), .Z(n2666) );
  AND U4467 ( .A(A[554]), .B(B[554]), .Z(n2662) );
  AND U4468 ( .A(B[555]), .B(A[555]), .Z(n2659) );
  AND U4469 ( .A(A[556]), .B(B[556]), .Z(n2648) );
  AND U4470 ( .A(A[557]), .B(B[557]), .Z(n2643) );
  AND U4471 ( .A(A[558]), .B(B[558]), .Z(n2639) );
  AND U4472 ( .A(B[559]), .B(A[559]), .Z(n2636) );
  NANDN U4473 ( .A(n2136), .B(n2531), .Z(n5703) );
  AND U4474 ( .A(n5816), .B(n5817), .Z(n2531) );
  ANDN U4475 ( .B(n5818), .A(n2624), .Z(n5817) );
  NAND U4476 ( .A(n5819), .B(n5820), .Z(n2624) );
  AND U4477 ( .A(n5821), .B(n5822), .Z(n5820) );
  AND U4478 ( .A(n2651), .B(n2646), .Z(n5822) );
  OR U4479 ( .A(A[557]), .B(B[557]), .Z(n2646) );
  OR U4480 ( .A(A[556]), .B(B[556]), .Z(n2651) );
  AND U4481 ( .A(n2641), .B(n2637), .Z(n5821) );
  OR U4482 ( .A(B[559]), .B(A[559]), .Z(n2637) );
  OR U4483 ( .A(A[558]), .B(B[558]), .Z(n2641) );
  ANDN U4484 ( .B(n5823), .A(n2704), .Z(n5819) );
  NAND U4485 ( .A(n5824), .B(n5825), .Z(n2704) );
  AND U4486 ( .A(n2721), .B(n2717), .Z(n5825) );
  OR U4487 ( .A(A[545]), .B(B[545]), .Z(n2717) );
  OR U4488 ( .A(A[544]), .B(B[544]), .Z(n2721) );
  AND U4489 ( .A(n2712), .B(n2708), .Z(n5824) );
  OR U4490 ( .A(B[547]), .B(A[547]), .Z(n2708) );
  OR U4491 ( .A(A[546]), .B(B[546]), .Z(n2712) );
  NOR U4492 ( .A(n2677), .B(n2655), .Z(n5823) );
  NAND U4493 ( .A(n5826), .B(n5827), .Z(n2655) );
  AND U4494 ( .A(n2673), .B(n2669), .Z(n5827) );
  OR U4495 ( .A(A[553]), .B(B[553]), .Z(n2669) );
  OR U4496 ( .A(A[552]), .B(B[552]), .Z(n2673) );
  AND U4497 ( .A(n2664), .B(n2660), .Z(n5826) );
  OR U4498 ( .A(B[555]), .B(A[555]), .Z(n2660) );
  OR U4499 ( .A(A[554]), .B(B[554]), .Z(n2664) );
  NAND U4500 ( .A(n5828), .B(n5829), .Z(n2677) );
  AND U4501 ( .A(n2700), .B(n2691), .Z(n5829) );
  OR U4502 ( .A(A[549]), .B(B[549]), .Z(n2691) );
  OR U4503 ( .A(A[548]), .B(B[548]), .Z(n2700) );
  AND U4504 ( .A(n2686), .B(n2682), .Z(n5828) );
  OR U4505 ( .A(B[551]), .B(A[551]), .Z(n2682) );
  OR U4506 ( .A(A[550]), .B(B[550]), .Z(n2686) );
  NOR U4507 ( .A(n2821), .B(n2725), .Z(n5818) );
  NAND U4508 ( .A(n5830), .B(n5831), .Z(n2725) );
  AND U4509 ( .A(n5832), .B(n5833), .Z(n5831) );
  AND U4510 ( .A(n2744), .B(n2739), .Z(n5833) );
  OR U4511 ( .A(A[541]), .B(B[541]), .Z(n2739) );
  OR U4512 ( .A(A[540]), .B(B[540]), .Z(n2744) );
  AND U4513 ( .A(n2734), .B(n2730), .Z(n5832) );
  OR U4514 ( .A(B[543]), .B(A[543]), .Z(n2730) );
  OR U4515 ( .A(A[542]), .B(B[542]), .Z(n2734) );
  ANDN U4516 ( .B(n5834), .A(n2796), .Z(n5830) );
  NAND U4517 ( .A(n5835), .B(n5836), .Z(n2796) );
  AND U4518 ( .A(n2816), .B(n2809), .Z(n5836) );
  OR U4519 ( .A(A[529]), .B(B[529]), .Z(n2809) );
  OR U4520 ( .A(A[528]), .B(B[528]), .Z(n2816) );
  AND U4521 ( .A(n2804), .B(n2800), .Z(n5835) );
  OR U4522 ( .A(B[531]), .B(A[531]), .Z(n2800) );
  OR U4523 ( .A(A[530]), .B(B[530]), .Z(n2804) );
  NOR U4524 ( .A(n2774), .B(n2748), .Z(n5834) );
  NAND U4525 ( .A(n5837), .B(n5838), .Z(n2748) );
  AND U4526 ( .A(n2770), .B(n2766), .Z(n5838) );
  OR U4527 ( .A(A[537]), .B(B[537]), .Z(n2766) );
  OR U4528 ( .A(A[536]), .B(B[536]), .Z(n2770) );
  AND U4529 ( .A(n2761), .B(n2757), .Z(n5837) );
  OR U4530 ( .A(B[539]), .B(A[539]), .Z(n2757) );
  OR U4531 ( .A(A[538]), .B(B[538]), .Z(n2761) );
  NAND U4532 ( .A(n5839), .B(n5840), .Z(n2774) );
  AND U4533 ( .A(n2792), .B(n2788), .Z(n5840) );
  OR U4534 ( .A(A[533]), .B(B[533]), .Z(n2788) );
  OR U4535 ( .A(A[532]), .B(B[532]), .Z(n2792) );
  AND U4536 ( .A(n2783), .B(n2779), .Z(n5839) );
  OR U4537 ( .A(B[535]), .B(A[535]), .Z(n2779) );
  OR U4538 ( .A(A[534]), .B(B[534]), .Z(n2783) );
  ANDN U4539 ( .B(n5841), .A(n2917), .Z(n2821) );
  AND U4540 ( .A(B[511]), .B(A[511]), .Z(n2917) );
  NANDN U4541 ( .A(n2916), .B(n5842), .Z(n5841) );
  NAND U4542 ( .A(n5843), .B(n5844), .Z(n5842) );
  NAND U4543 ( .A(n5845), .B(n5846), .Z(n5844) );
  AND U4544 ( .A(n5847), .B(n5848), .Z(n5846) );
  ANDN U4545 ( .B(n2926), .A(n2935), .Z(n5848) );
  AND U4546 ( .A(n2921), .B(n5849), .Z(n5847) );
  NANDN U4547 ( .A(n3013), .B(n5850), .Z(n5849) );
  NANDN U4548 ( .A(n3015), .B(n5851), .Z(n5850) );
  NANDN U4549 ( .A(n3102), .B(n5852), .Z(n5851) );
  NANDN U4550 ( .A(n3104), .B(n5853), .Z(n5852) );
  NANDN U4551 ( .A(n3203), .B(n5854), .Z(n5853) );
  NANDN U4552 ( .A(n3205), .B(n5855), .Z(n5854) );
  NANDN U4553 ( .A(n3301), .B(n5856), .Z(n5855) );
  NANDN U4554 ( .A(n3303), .B(n5857), .Z(n5856) );
  NANDN U4555 ( .A(n3689), .B(n5858), .Z(n5857) );
  AND U4556 ( .A(n5859), .B(n5860), .Z(n5858) );
  NANDN U4557 ( .A(n3691), .B(n4068), .Z(n5860) );
  NAND U4558 ( .A(n5861), .B(n5862), .Z(n4068) );
  NAND U4559 ( .A(n5863), .B(n4081), .Z(n5862) );
  NANDN U4560 ( .A(n4083), .B(n5864), .Z(n5863) );
  NAND U4561 ( .A(n5865), .B(n4085), .Z(n5864) );
  NANDN U4562 ( .A(n4087), .B(n5866), .Z(n5865) );
  NAND U4563 ( .A(n5867), .B(n4090), .Z(n5866) );
  NANDN U4564 ( .A(n4092), .B(n5868), .Z(n5867) );
  NAND U4565 ( .A(n5869), .B(n4095), .Z(n5868) );
  NANDN U4566 ( .A(n4097), .B(n5870), .Z(n5869) );
  NANDN U4567 ( .A(n4099), .B(n5871), .Z(n5870) );
  NANDN U4568 ( .A(n4119), .B(n5872), .Z(n5871) );
  NANDN U4569 ( .A(n4121), .B(n4147), .Z(n5872) );
  NANDN U4570 ( .A(n4152), .B(n5873), .Z(n4147) );
  NAND U4571 ( .A(n5874), .B(n4153), .Z(n5873) );
  NANDN U4572 ( .A(n4155), .B(n5875), .Z(n5874) );
  NAND U4573 ( .A(n5876), .B(n4157), .Z(n5875) );
  NANDN U4574 ( .A(n4159), .B(n5877), .Z(n5876) );
  NAND U4575 ( .A(n4162), .B(n4164), .Z(n5877) );
  AND U4576 ( .A(A[304]), .B(B[304]), .Z(n4164) );
  AND U4577 ( .A(A[305]), .B(B[305]), .Z(n4159) );
  AND U4578 ( .A(A[306]), .B(B[306]), .Z(n4155) );
  AND U4579 ( .A(B[307]), .B(A[307]), .Z(n4152) );
  NANDN U4580 ( .A(n4125), .B(n5878), .Z(n4119) );
  NAND U4581 ( .A(n5879), .B(n4126), .Z(n5878) );
  NANDN U4582 ( .A(n4128), .B(n5880), .Z(n5879) );
  NAND U4583 ( .A(n5881), .B(n4130), .Z(n5880) );
  NANDN U4584 ( .A(n4132), .B(n5882), .Z(n5881) );
  NAND U4585 ( .A(n4135), .B(n4142), .Z(n5882) );
  AND U4586 ( .A(A[308]), .B(B[308]), .Z(n4142) );
  AND U4587 ( .A(A[309]), .B(B[309]), .Z(n4132) );
  AND U4588 ( .A(A[310]), .B(B[310]), .Z(n4128) );
  AND U4589 ( .A(B[311]), .B(A[311]), .Z(n4125) );
  NANDN U4590 ( .A(n4103), .B(n5883), .Z(n4097) );
  NAND U4591 ( .A(n5884), .B(n4104), .Z(n5883) );
  NANDN U4592 ( .A(n4106), .B(n5885), .Z(n5884) );
  NAND U4593 ( .A(n5886), .B(n4108), .Z(n5885) );
  NANDN U4594 ( .A(n4110), .B(n5887), .Z(n5886) );
  NAND U4595 ( .A(n4113), .B(n4115), .Z(n5887) );
  AND U4596 ( .A(A[312]), .B(B[312]), .Z(n4115) );
  AND U4597 ( .A(A[313]), .B(B[313]), .Z(n4110) );
  AND U4598 ( .A(A[314]), .B(B[314]), .Z(n4106) );
  AND U4599 ( .A(B[315]), .B(A[315]), .Z(n4103) );
  AND U4600 ( .A(A[316]), .B(B[316]), .Z(n4092) );
  AND U4601 ( .A(A[317]), .B(B[317]), .Z(n4087) );
  AND U4602 ( .A(A[318]), .B(B[318]), .Z(n4083) );
  ANDN U4603 ( .B(n5888), .A(n4080), .Z(n5861) );
  AND U4604 ( .A(B[319]), .B(A[319]), .Z(n4080) );
  NANDN U4605 ( .A(n5889), .B(n5890), .Z(n5888) );
  NANDN U4606 ( .A(n4168), .B(n5891), .Z(n5890) );
  NANDN U4607 ( .A(n4170), .B(n5892), .Z(n5891) );
  NANDN U4608 ( .A(n4266), .B(n5893), .Z(n5892) );
  NANDN U4609 ( .A(n4268), .B(n4363), .Z(n5893) );
  NANDN U4610 ( .A(n4368), .B(n5894), .Z(n4363) );
  NAND U4611 ( .A(n5895), .B(n4369), .Z(n5894) );
  NANDN U4612 ( .A(n4371), .B(n5896), .Z(n5895) );
  NAND U4613 ( .A(n5897), .B(n4373), .Z(n5896) );
  NANDN U4614 ( .A(n4375), .B(n5898), .Z(n5897) );
  NAND U4615 ( .A(n5899), .B(n4378), .Z(n5898) );
  NANDN U4616 ( .A(n4385), .B(n5900), .Z(n5899) );
  NAND U4617 ( .A(n5901), .B(n4388), .Z(n5900) );
  NANDN U4618 ( .A(n4390), .B(n5902), .Z(n5901) );
  NANDN U4619 ( .A(n4392), .B(n5903), .Z(n5902) );
  NANDN U4620 ( .A(n4412), .B(n5904), .Z(n5903) );
  NANDN U4621 ( .A(n4414), .B(n4435), .Z(n5904) );
  NANDN U4622 ( .A(n4443), .B(n5905), .Z(n4435) );
  NAND U4623 ( .A(n5906), .B(n4444), .Z(n5905) );
  NANDN U4624 ( .A(n4446), .B(n5907), .Z(n5906) );
  NAND U4625 ( .A(n5908), .B(n4448), .Z(n5907) );
  NANDN U4626 ( .A(n4450), .B(n5909), .Z(n5908) );
  NAND U4627 ( .A(n4453), .B(n4455), .Z(n5909) );
  AND U4628 ( .A(A[256]), .B(B[256]), .Z(n4455) );
  AND U4629 ( .A(A[257]), .B(B[257]), .Z(n4450) );
  AND U4630 ( .A(A[258]), .B(B[258]), .Z(n4446) );
  AND U4631 ( .A(B[259]), .B(A[259]), .Z(n4443) );
  NANDN U4632 ( .A(n4418), .B(n5910), .Z(n4412) );
  NAND U4633 ( .A(n5911), .B(n4419), .Z(n5910) );
  NANDN U4634 ( .A(n4421), .B(n5912), .Z(n5911) );
  NAND U4635 ( .A(n5913), .B(n4423), .Z(n5912) );
  NANDN U4636 ( .A(n4425), .B(n5914), .Z(n5913) );
  NAND U4637 ( .A(n4428), .B(n4430), .Z(n5914) );
  AND U4638 ( .A(A[260]), .B(B[260]), .Z(n4430) );
  AND U4639 ( .A(A[261]), .B(B[261]), .Z(n4425) );
  AND U4640 ( .A(A[262]), .B(B[262]), .Z(n4421) );
  AND U4641 ( .A(B[263]), .B(A[263]), .Z(n4418) );
  NANDN U4642 ( .A(n4396), .B(n5915), .Z(n4390) );
  NAND U4643 ( .A(n5916), .B(n4397), .Z(n5915) );
  NANDN U4644 ( .A(n4399), .B(n5917), .Z(n5916) );
  NAND U4645 ( .A(n5918), .B(n4401), .Z(n5917) );
  NANDN U4646 ( .A(n4403), .B(n5919), .Z(n5918) );
  NAND U4647 ( .A(n4406), .B(n4408), .Z(n5919) );
  AND U4648 ( .A(A[264]), .B(B[264]), .Z(n4408) );
  AND U4649 ( .A(A[265]), .B(B[265]), .Z(n4403) );
  AND U4650 ( .A(A[266]), .B(B[266]), .Z(n4399) );
  AND U4651 ( .A(B[267]), .B(A[267]), .Z(n4396) );
  AND U4652 ( .A(A[268]), .B(B[268]), .Z(n4385) );
  AND U4653 ( .A(A[269]), .B(B[269]), .Z(n4375) );
  AND U4654 ( .A(A[270]), .B(B[270]), .Z(n4371) );
  AND U4655 ( .A(B[271]), .B(A[271]), .Z(n4368) );
  NANDN U4656 ( .A(n4272), .B(n5920), .Z(n4266) );
  NAND U4657 ( .A(n5921), .B(n4273), .Z(n5920) );
  NANDN U4658 ( .A(n4275), .B(n5922), .Z(n5921) );
  NAND U4659 ( .A(n5923), .B(n4277), .Z(n5922) );
  NANDN U4660 ( .A(n4279), .B(n5924), .Z(n5923) );
  NAND U4661 ( .A(n5925), .B(n4282), .Z(n5924) );
  NANDN U4662 ( .A(n4284), .B(n5926), .Z(n5925) );
  NAND U4663 ( .A(n5927), .B(n4287), .Z(n5926) );
  NANDN U4664 ( .A(n4289), .B(n5928), .Z(n5927) );
  NANDN U4665 ( .A(n4291), .B(n5929), .Z(n5928) );
  NANDN U4666 ( .A(n4311), .B(n5930), .Z(n5929) );
  NANDN U4667 ( .A(n4313), .B(n4342), .Z(n5930) );
  NANDN U4668 ( .A(n4346), .B(n5931), .Z(n4342) );
  NAND U4669 ( .A(n5932), .B(n4347), .Z(n5931) );
  NANDN U4670 ( .A(n4349), .B(n5933), .Z(n5932) );
  NAND U4671 ( .A(n5934), .B(n4351), .Z(n5933) );
  NANDN U4672 ( .A(n4353), .B(n5935), .Z(n5934) );
  NAND U4673 ( .A(n4356), .B(n4358), .Z(n5935) );
  AND U4674 ( .A(A[272]), .B(B[272]), .Z(n4358) );
  AND U4675 ( .A(A[273]), .B(B[273]), .Z(n4353) );
  AND U4676 ( .A(A[274]), .B(B[274]), .Z(n4349) );
  AND U4677 ( .A(B[275]), .B(A[275]), .Z(n4346) );
  NANDN U4678 ( .A(n4325), .B(n5936), .Z(n4311) );
  NAND U4679 ( .A(n5937), .B(n4326), .Z(n5936) );
  NANDN U4680 ( .A(n4328), .B(n5938), .Z(n5937) );
  NAND U4681 ( .A(n5939), .B(n4330), .Z(n5938) );
  NANDN U4682 ( .A(n4332), .B(n5940), .Z(n5939) );
  NAND U4683 ( .A(n4335), .B(n4337), .Z(n5940) );
  AND U4684 ( .A(A[276]), .B(B[276]), .Z(n4337) );
  AND U4685 ( .A(A[277]), .B(B[277]), .Z(n4332) );
  AND U4686 ( .A(A[278]), .B(B[278]), .Z(n4328) );
  AND U4687 ( .A(B[279]), .B(A[279]), .Z(n4325) );
  NANDN U4688 ( .A(n4295), .B(n5941), .Z(n4289) );
  NAND U4689 ( .A(n5942), .B(n4296), .Z(n5941) );
  NANDN U4690 ( .A(n4298), .B(n5943), .Z(n5942) );
  NAND U4691 ( .A(n5944), .B(n4300), .Z(n5943) );
  NANDN U4692 ( .A(n4302), .B(n5945), .Z(n5944) );
  NAND U4693 ( .A(n4305), .B(n4307), .Z(n5945) );
  AND U4694 ( .A(A[280]), .B(B[280]), .Z(n4307) );
  AND U4695 ( .A(A[281]), .B(B[281]), .Z(n4302) );
  AND U4696 ( .A(A[282]), .B(B[282]), .Z(n4298) );
  AND U4697 ( .A(B[283]), .B(A[283]), .Z(n4295) );
  AND U4698 ( .A(A[284]), .B(B[284]), .Z(n4284) );
  AND U4699 ( .A(A[285]), .B(B[285]), .Z(n4279) );
  AND U4700 ( .A(A[286]), .B(B[286]), .Z(n4275) );
  AND U4701 ( .A(B[287]), .B(A[287]), .Z(n4272) );
  NANDN U4702 ( .A(n4174), .B(n5946), .Z(n4168) );
  NAND U4703 ( .A(n5947), .B(n4175), .Z(n5946) );
  NANDN U4704 ( .A(n4177), .B(n5948), .Z(n5947) );
  NAND U4705 ( .A(n5949), .B(n4179), .Z(n5948) );
  NANDN U4706 ( .A(n4181), .B(n5950), .Z(n5949) );
  NAND U4707 ( .A(n5951), .B(n4184), .Z(n5950) );
  NANDN U4708 ( .A(n4186), .B(n5952), .Z(n5951) );
  NAND U4709 ( .A(n5953), .B(n4189), .Z(n5952) );
  NANDN U4710 ( .A(n4191), .B(n5954), .Z(n5953) );
  NANDN U4711 ( .A(n4193), .B(n5955), .Z(n5954) );
  NANDN U4712 ( .A(n4218), .B(n5956), .Z(n5955) );
  NANDN U4713 ( .A(n4220), .B(n4241), .Z(n5956) );
  NANDN U4714 ( .A(n4245), .B(n5957), .Z(n4241) );
  NAND U4715 ( .A(n5958), .B(n4246), .Z(n5957) );
  NANDN U4716 ( .A(n4248), .B(n5959), .Z(n5958) );
  NAND U4717 ( .A(n5960), .B(n4250), .Z(n5959) );
  NANDN U4718 ( .A(n4252), .B(n5961), .Z(n5960) );
  NAND U4719 ( .A(n4255), .B(n4262), .Z(n5961) );
  AND U4720 ( .A(A[288]), .B(B[288]), .Z(n4262) );
  AND U4721 ( .A(A[289]), .B(B[289]), .Z(n4252) );
  AND U4722 ( .A(A[290]), .B(B[290]), .Z(n4248) );
  AND U4723 ( .A(B[291]), .B(A[291]), .Z(n4245) );
  NANDN U4724 ( .A(n4224), .B(n5962), .Z(n4218) );
  NAND U4725 ( .A(n5963), .B(n4225), .Z(n5962) );
  NANDN U4726 ( .A(n4227), .B(n5964), .Z(n5963) );
  NAND U4727 ( .A(n5965), .B(n4229), .Z(n5964) );
  NANDN U4728 ( .A(n4231), .B(n5966), .Z(n5965) );
  NAND U4729 ( .A(n4234), .B(n4236), .Z(n5966) );
  AND U4730 ( .A(A[292]), .B(B[292]), .Z(n4236) );
  AND U4731 ( .A(A[293]), .B(B[293]), .Z(n4231) );
  AND U4732 ( .A(A[294]), .B(B[294]), .Z(n4227) );
  AND U4733 ( .A(B[295]), .B(A[295]), .Z(n4224) );
  NANDN U4734 ( .A(n4202), .B(n5967), .Z(n4191) );
  NAND U4735 ( .A(n5968), .B(n4203), .Z(n5967) );
  NANDN U4736 ( .A(n4205), .B(n5969), .Z(n5968) );
  NAND U4737 ( .A(n5970), .B(n4207), .Z(n5969) );
  NANDN U4738 ( .A(n4209), .B(n5971), .Z(n5970) );
  NAND U4739 ( .A(n4212), .B(n4214), .Z(n5971) );
  AND U4740 ( .A(A[296]), .B(B[296]), .Z(n4214) );
  AND U4741 ( .A(A[297]), .B(B[297]), .Z(n4209) );
  AND U4742 ( .A(A[298]), .B(B[298]), .Z(n4205) );
  AND U4743 ( .A(B[299]), .B(A[299]), .Z(n4202) );
  AND U4744 ( .A(A[300]), .B(B[300]), .Z(n4186) );
  AND U4745 ( .A(A[301]), .B(B[301]), .Z(n4181) );
  AND U4746 ( .A(A[302]), .B(B[302]), .Z(n4177) );
  AND U4747 ( .A(B[303]), .B(A[303]), .Z(n4174) );
  NANDN U4748 ( .A(n3691), .B(n4069), .Z(n5859) );
  AND U4749 ( .A(n5972), .B(n5973), .Z(n4069) );
  ANDN U4750 ( .B(n5974), .A(n4170), .Z(n5973) );
  NAND U4751 ( .A(n5975), .B(n5976), .Z(n4170) );
  AND U4752 ( .A(n5977), .B(n5978), .Z(n5976) );
  AND U4753 ( .A(n4189), .B(n4184), .Z(n5978) );
  OR U4754 ( .A(A[301]), .B(B[301]), .Z(n4184) );
  OR U4755 ( .A(A[300]), .B(B[300]), .Z(n4189) );
  AND U4756 ( .A(n4179), .B(n4175), .Z(n5977) );
  OR U4757 ( .A(B[303]), .B(A[303]), .Z(n4175) );
  OR U4758 ( .A(A[302]), .B(B[302]), .Z(n4179) );
  ANDN U4759 ( .B(n5979), .A(n4242), .Z(n5975) );
  NAND U4760 ( .A(n5980), .B(n5981), .Z(n4242) );
  AND U4761 ( .A(n4264), .B(n4255), .Z(n5981) );
  OR U4762 ( .A(A[289]), .B(B[289]), .Z(n4255) );
  OR U4763 ( .A(A[288]), .B(B[288]), .Z(n4264) );
  AND U4764 ( .A(n4250), .B(n4246), .Z(n5980) );
  OR U4765 ( .A(B[291]), .B(A[291]), .Z(n4246) );
  OR U4766 ( .A(A[290]), .B(B[290]), .Z(n4250) );
  NOR U4767 ( .A(n4220), .B(n4193), .Z(n5979) );
  NAND U4768 ( .A(n5982), .B(n5983), .Z(n4193) );
  AND U4769 ( .A(n4216), .B(n4212), .Z(n5983) );
  OR U4770 ( .A(A[297]), .B(B[297]), .Z(n4212) );
  OR U4771 ( .A(A[296]), .B(B[296]), .Z(n4216) );
  AND U4772 ( .A(n4207), .B(n4203), .Z(n5982) );
  OR U4773 ( .A(B[299]), .B(A[299]), .Z(n4203) );
  OR U4774 ( .A(A[298]), .B(B[298]), .Z(n4207) );
  NAND U4775 ( .A(n5984), .B(n5985), .Z(n4220) );
  AND U4776 ( .A(n4238), .B(n4234), .Z(n5985) );
  OR U4777 ( .A(A[293]), .B(B[293]), .Z(n4234) );
  OR U4778 ( .A(A[292]), .B(B[292]), .Z(n4238) );
  AND U4779 ( .A(n4229), .B(n4225), .Z(n5984) );
  OR U4780 ( .A(B[295]), .B(A[295]), .Z(n4225) );
  OR U4781 ( .A(A[294]), .B(B[294]), .Z(n4229) );
  NOR U4782 ( .A(n4365), .B(n4268), .Z(n5974) );
  NAND U4783 ( .A(n5986), .B(n5987), .Z(n4268) );
  AND U4784 ( .A(n5988), .B(n5989), .Z(n5987) );
  AND U4785 ( .A(n4287), .B(n4282), .Z(n5989) );
  OR U4786 ( .A(A[285]), .B(B[285]), .Z(n4282) );
  OR U4787 ( .A(A[284]), .B(B[284]), .Z(n4287) );
  AND U4788 ( .A(n4277), .B(n4273), .Z(n5988) );
  OR U4789 ( .A(B[287]), .B(A[287]), .Z(n4273) );
  OR U4790 ( .A(A[286]), .B(B[286]), .Z(n4277) );
  ANDN U4791 ( .B(n5990), .A(n4343), .Z(n5986) );
  NAND U4792 ( .A(n5991), .B(n5992), .Z(n4343) );
  AND U4793 ( .A(n4360), .B(n4356), .Z(n5992) );
  OR U4794 ( .A(A[273]), .B(B[273]), .Z(n4356) );
  OR U4795 ( .A(A[272]), .B(B[272]), .Z(n4360) );
  AND U4796 ( .A(n4351), .B(n4347), .Z(n5991) );
  OR U4797 ( .A(B[275]), .B(A[275]), .Z(n4347) );
  OR U4798 ( .A(A[274]), .B(B[274]), .Z(n4351) );
  NOR U4799 ( .A(n4313), .B(n4291), .Z(n5990) );
  NAND U4800 ( .A(n5993), .B(n5994), .Z(n4291) );
  AND U4801 ( .A(n4309), .B(n4305), .Z(n5994) );
  OR U4802 ( .A(A[281]), .B(B[281]), .Z(n4305) );
  OR U4803 ( .A(A[280]), .B(B[280]), .Z(n4309) );
  AND U4804 ( .A(n4300), .B(n4296), .Z(n5993) );
  OR U4805 ( .A(B[283]), .B(A[283]), .Z(n4296) );
  OR U4806 ( .A(A[282]), .B(B[282]), .Z(n4300) );
  NAND U4807 ( .A(n5995), .B(n5996), .Z(n4313) );
  AND U4808 ( .A(n4339), .B(n4335), .Z(n5996) );
  OR U4809 ( .A(A[277]), .B(B[277]), .Z(n4335) );
  OR U4810 ( .A(A[276]), .B(B[276]), .Z(n4339) );
  AND U4811 ( .A(n4330), .B(n4326), .Z(n5995) );
  OR U4812 ( .A(B[279]), .B(A[279]), .Z(n4326) );
  OR U4813 ( .A(A[278]), .B(B[278]), .Z(n4330) );
  ANDN U4814 ( .B(n5997), .A(n4462), .Z(n4365) );
  AND U4815 ( .A(B[255]), .B(A[255]), .Z(n4462) );
  NANDN U4816 ( .A(n4461), .B(n5998), .Z(n5997) );
  NANDN U4817 ( .A(n4464), .B(n5999), .Z(n5998) );
  NANDN U4818 ( .A(n4465), .B(n6000), .Z(n5999) );
  NANDN U4819 ( .A(n4468), .B(n6001), .Z(n6000) );
  NANDN U4820 ( .A(n4470), .B(n6002), .Z(n6001) );
  NAND U4821 ( .A(n6003), .B(n6004), .Z(n6002) );
  NAND U4822 ( .A(n6005), .B(n6006), .Z(n6004) );
  AND U4823 ( .A(n4508), .B(n6007), .Z(n6006) );
  ANDN U4824 ( .B(n4476), .A(n4530), .Z(n6007) );
  ANDN U4825 ( .B(n6008), .A(n4560), .Z(n4530) );
  AND U4826 ( .A(B[239]), .B(A[239]), .Z(n4560) );
  NANDN U4827 ( .A(n4559), .B(n6009), .Z(n6008) );
  NANDN U4828 ( .A(n4562), .B(n6010), .Z(n6009) );
  NANDN U4829 ( .A(n4563), .B(n6011), .Z(n6010) );
  NANDN U4830 ( .A(n4566), .B(n6012), .Z(n6011) );
  NANDN U4831 ( .A(n4568), .B(n6013), .Z(n6012) );
  NAND U4832 ( .A(n6014), .B(n6015), .Z(n6013) );
  NAND U4833 ( .A(n6016), .B(n6017), .Z(n6015) );
  AND U4834 ( .A(n4601), .B(n6018), .Z(n6017) );
  ANDN U4835 ( .B(n4574), .A(n4628), .Z(n6018) );
  ANDN U4836 ( .B(n6019), .A(n4650), .Z(n4628) );
  AND U4837 ( .A(B[223]), .B(A[223]), .Z(n4650) );
  NANDN U4838 ( .A(n4649), .B(n6020), .Z(n6019) );
  NANDN U4839 ( .A(n4652), .B(n6021), .Z(n6020) );
  NANDN U4840 ( .A(n4653), .B(n6022), .Z(n6021) );
  NANDN U4841 ( .A(n4656), .B(n6023), .Z(n6022) );
  NANDN U4842 ( .A(n4658), .B(n6024), .Z(n6023) );
  NAND U4843 ( .A(n6025), .B(n6026), .Z(n6024) );
  NAND U4844 ( .A(n6027), .B(n6028), .Z(n6026) );
  AND U4845 ( .A(n4695), .B(n6029), .Z(n6028) );
  ANDN U4846 ( .B(n4664), .A(n4717), .Z(n6029) );
  ANDN U4847 ( .B(n6030), .A(n4744), .Z(n4717) );
  AND U4848 ( .A(B[207]), .B(A[207]), .Z(n4744) );
  NANDN U4849 ( .A(n4743), .B(n6031), .Z(n6030) );
  NANDN U4850 ( .A(n4746), .B(n6032), .Z(n6031) );
  NANDN U4851 ( .A(n4747), .B(n6033), .Z(n6032) );
  NANDN U4852 ( .A(n4750), .B(n6034), .Z(n6033) );
  NANDN U4853 ( .A(n4752), .B(n6035), .Z(n6034) );
  NAND U4854 ( .A(n6036), .B(n6037), .Z(n6035) );
  NAND U4855 ( .A(n6038), .B(n6039), .Z(n6037) );
  AND U4856 ( .A(n4785), .B(n6040), .Z(n6039) );
  ANDN U4857 ( .B(n4758), .A(n4815), .Z(n6040) );
  ANDN U4858 ( .B(n6041), .A(n4837), .Z(n4815) );
  AND U4859 ( .A(B[191]), .B(A[191]), .Z(n4837) );
  NANDN U4860 ( .A(n4836), .B(n6042), .Z(n6041) );
  NAND U4861 ( .A(n6043), .B(n6044), .Z(n6042) );
  NAND U4862 ( .A(n6045), .B(n6046), .Z(n6044) );
  AND U4863 ( .A(n6047), .B(n6048), .Z(n6046) );
  ANDN U4864 ( .B(n4846), .A(n4855), .Z(n6048) );
  AND U4865 ( .A(n4841), .B(n4905), .Z(n6047) );
  NANDN U4866 ( .A(n6049), .B(n6050), .Z(n4905) );
  NANDN U4867 ( .A(n6051), .B(n4995), .Z(n6050) );
  NANDN U4868 ( .A(n6052), .B(n6053), .Z(n4995) );
  NANDN U4869 ( .A(n6054), .B(n5088), .Z(n6053) );
  NANDN U4870 ( .A(n6055), .B(n6056), .Z(n5088) );
  OR U4871 ( .A(n6057), .B(n5177), .Z(n6056) );
  ANDN U4872 ( .B(n6058), .A(n5203), .Z(n5177) );
  AND U4873 ( .A(B[127]), .B(A[127]), .Z(n5203) );
  NANDN U4874 ( .A(n5202), .B(n6059), .Z(n6058) );
  NAND U4875 ( .A(n6060), .B(n6061), .Z(n6059) );
  NAND U4876 ( .A(n6062), .B(n6063), .Z(n6061) );
  AND U4877 ( .A(n6064), .B(n6065), .Z(n6063) );
  ANDN U4878 ( .B(n5212), .A(n5216), .Z(n6065) );
  AND U4879 ( .A(n5207), .B(n6066), .Z(n6064) );
  NANDN U4880 ( .A(n5293), .B(n6067), .Z(n6066) );
  NANDN U4881 ( .A(n5295), .B(n6068), .Z(n6067) );
  NANDN U4882 ( .A(n5427), .B(n6069), .Z(n6068) );
  NANDN U4883 ( .A(n5428), .B(n6070), .Z(n6069) );
  NANDN U4884 ( .A(n5430), .B(n5429), .Z(n6070) );
  OR U4885 ( .A(n6071), .B(n1847), .Z(n5429) );
  ANDN U4886 ( .B(n6072), .A(n2141), .Z(n1847) );
  AND U4887 ( .A(B[63]), .B(A[63]), .Z(n2141) );
  NANDN U4888 ( .A(n2140), .B(n6073), .Z(n6072) );
  NANDN U4889 ( .A(n2143), .B(n6074), .Z(n6073) );
  NANDN U4890 ( .A(n2144), .B(n6075), .Z(n6074) );
  NANDN U4891 ( .A(n2205), .B(n6076), .Z(n6075) );
  NANDN U4892 ( .A(n2207), .B(n6077), .Z(n6076) );
  NANDN U4893 ( .A(n2264), .B(n6078), .Z(n6077) );
  NANDN U4894 ( .A(n2266), .B(n6079), .Z(n6078) );
  NANDN U4895 ( .A(n2325), .B(n6080), .Z(n6079) );
  NANDN U4896 ( .A(n2327), .B(n6081), .Z(n6080) );
  NANDN U4897 ( .A(n2569), .B(n6082), .Z(n6081) );
  AND U4898 ( .A(n6083), .B(n6084), .Z(n6082) );
  NANDN U4899 ( .A(n2571), .B(n2811), .Z(n6084) );
  NANDN U4900 ( .A(n2869), .B(n6085), .Z(n2811) );
  NAND U4901 ( .A(n6086), .B(n2870), .Z(n6085) );
  NANDN U4902 ( .A(n2872), .B(n6087), .Z(n6086) );
  NAND U4903 ( .A(n6088), .B(n2874), .Z(n6087) );
  NANDN U4904 ( .A(n2928), .B(n6089), .Z(n6088) );
  NAND U4905 ( .A(n2931), .B(n2991), .Z(n6089) );
  AND U4906 ( .A(A[48]), .B(B[48]), .Z(n2991) );
  AND U4907 ( .A(A[49]), .B(B[49]), .Z(n2928) );
  AND U4908 ( .A(A[50]), .B(B[50]), .Z(n2872) );
  AND U4909 ( .A(B[51]), .B(A[51]), .Z(n2869) );
  NANDN U4910 ( .A(n2571), .B(n2812), .Z(n6083) );
  AND U4911 ( .A(n6090), .B(n6091), .Z(n2812) );
  AND U4912 ( .A(n2874), .B(n6092), .Z(n6091) );
  AND U4913 ( .A(n2994), .B(n2931), .Z(n6092) );
  OR U4914 ( .A(A[49]), .B(B[49]), .Z(n2931) );
  OR U4915 ( .A(A[48]), .B(B[48]), .Z(n2994) );
  OR U4916 ( .A(A[50]), .B(B[50]), .Z(n2874) );
  ANDN U4917 ( .B(n2870), .A(n2993), .Z(n6090) );
  ANDN U4918 ( .B(n6093), .A(n3109), .Z(n2993) );
  AND U4919 ( .A(B[47]), .B(A[47]), .Z(n3109) );
  NANDN U4920 ( .A(n3108), .B(n6094), .Z(n6093) );
  NANDN U4921 ( .A(n3111), .B(n6095), .Z(n6094) );
  NANDN U4922 ( .A(n3112), .B(n6096), .Z(n6095) );
  NANDN U4923 ( .A(n3173), .B(n6097), .Z(n6096) );
  NANDN U4924 ( .A(n3175), .B(n6098), .Z(n6097) );
  NAND U4925 ( .A(n6099), .B(n6100), .Z(n6098) );
  NAND U4926 ( .A(n6101), .B(n6102), .Z(n6100) );
  AND U4927 ( .A(n3539), .B(n6103), .Z(n6102) );
  ANDN U4928 ( .B(n3234), .A(n3781), .Z(n6103) );
  ANDN U4929 ( .B(n6104), .A(n4073), .Z(n3781) );
  AND U4930 ( .A(B[31]), .B(A[31]), .Z(n4073) );
  NANDN U4931 ( .A(n4072), .B(n6105), .Z(n6104) );
  NANDN U4932 ( .A(n4075), .B(n6106), .Z(n6105) );
  NANDN U4933 ( .A(n4076), .B(n6107), .Z(n6106) );
  NANDN U4934 ( .A(n4137), .B(n6108), .Z(n6107) );
  NANDN U4935 ( .A(n4139), .B(n6109), .Z(n6108) );
  NAND U4936 ( .A(n6110), .B(n6111), .Z(n6109) );
  NAND U4937 ( .A(n6112), .B(n6113), .Z(n6111) );
  AND U4938 ( .A(n4499), .B(n6114), .Z(n6113) );
  ANDN U4939 ( .B(n4199), .A(n4735), .Z(n6114) );
  ANDN U4940 ( .B(n6115), .A(n5016), .Z(n4735) );
  AND U4941 ( .A(B[15]), .B(A[15]), .Z(n5016) );
  NAND U4942 ( .A(n5014), .B(n5017), .Z(n6115) );
  OR U4943 ( .A(B[15]), .B(A[15]), .Z(n5017) );
  NANDN U4944 ( .A(n5078), .B(n6116), .Z(n5014) );
  NAND U4945 ( .A(n5076), .B(n5079), .Z(n6116) );
  OR U4946 ( .A(B[14]), .B(A[14]), .Z(n5079) );
  NANDN U4947 ( .A(n5132), .B(n6117), .Z(n5076) );
  NAND U4948 ( .A(n5130), .B(n5133), .Z(n6117) );
  OR U4949 ( .A(B[13]), .B(A[13]), .Z(n5133) );
  NANDN U4950 ( .A(n5193), .B(n6118), .Z(n5130) );
  NAND U4951 ( .A(n5191), .B(n5194), .Z(n6118) );
  OR U4952 ( .A(B[12]), .B(A[12]), .Z(n5194) );
  NANDN U4953 ( .A(n5248), .B(n6119), .Z(n5191) );
  NANDN U4954 ( .A(n5247), .B(n6120), .Z(n6119) );
  NANDN U4955 ( .A(n5250), .B(n6121), .Z(n6120) );
  NANDN U4956 ( .A(n5251), .B(n6122), .Z(n6121) );
  NANDN U4957 ( .A(n3), .B(n6123), .Z(n6122) );
  NAND U4958 ( .A(n6124), .B(n4), .Z(n6123) );
  OR U4959 ( .A(A[9]), .B(B[9]), .Z(n4) );
  NANDN U4960 ( .A(n591), .B(n5311), .Z(n6124) );
  OR U4961 ( .A(n588), .B(n590), .Z(n5311) );
  NOR U4962 ( .A(B[8]), .B(A[8]), .Z(n590) );
  ANDN U4963 ( .B(n6125), .A(n1172), .Z(n588) );
  AND U4964 ( .A(B[7]), .B(A[7]), .Z(n1172) );
  NANDN U4965 ( .A(n1171), .B(n6126), .Z(n6125) );
  NANDN U4966 ( .A(n1174), .B(n1173), .Z(n6126) );
  NANDN U4967 ( .A(n1781), .B(n1779), .Z(n1173) );
  NANDN U4968 ( .A(n2386), .B(n6127), .Z(n1779) );
  NANDN U4969 ( .A(n2385), .B(n2383), .Z(n6127) );
  NANDN U4970 ( .A(n2989), .B(n6128), .Z(n2383) );
  NAND U4971 ( .A(n2988), .B(n2986), .Z(n6128) );
  AND U4972 ( .A(A[3]), .B(B[3]), .Z(n2986) );
  OR U4973 ( .A(B[4]), .B(A[4]), .Z(n2988) );
  AND U4974 ( .A(B[4]), .B(A[4]), .Z(n2989) );
  NOR U4975 ( .A(B[5]), .B(A[5]), .Z(n2385) );
  AND U4976 ( .A(B[5]), .B(A[5]), .Z(n2386) );
  NOR U4977 ( .A(B[6]), .B(A[6]), .Z(n1781) );
  AND U4978 ( .A(B[6]), .B(A[6]), .Z(n1174) );
  NOR U4979 ( .A(B[7]), .B(A[7]), .Z(n1171) );
  AND U4980 ( .A(B[8]), .B(A[8]), .Z(n591) );
  AND U4981 ( .A(B[9]), .B(A[9]), .Z(n3) );
  NOR U4982 ( .A(B[10]), .B(A[10]), .Z(n5251) );
  AND U4983 ( .A(B[10]), .B(A[10]), .Z(n5250) );
  NOR U4984 ( .A(B[11]), .B(A[11]), .Z(n5247) );
  AND U4985 ( .A(B[11]), .B(A[11]), .Z(n5248) );
  AND U4986 ( .A(B[12]), .B(A[12]), .Z(n5193) );
  AND U4987 ( .A(B[13]), .B(A[13]), .Z(n5132) );
  AND U4988 ( .A(B[14]), .B(A[14]), .Z(n5078) );
  NOR U4989 ( .A(n4734), .B(n4259), .Z(n6112) );
  NAND U4990 ( .A(n6129), .B(n6130), .Z(n4734) );
  AND U4991 ( .A(n4909), .B(n4851), .Z(n6130) );
  OR U4992 ( .A(B[16]), .B(A[16]), .Z(n4909) );
  ANDN U4993 ( .B(n4789), .A(n4792), .Z(n6129) );
  ANDN U4994 ( .B(n6131), .A(n4196), .Z(n6110) );
  AND U4995 ( .A(B[28]), .B(A[28]), .Z(n4196) );
  NAND U4996 ( .A(n6132), .B(n4199), .Z(n6131) );
  OR U4997 ( .A(A[28]), .B(B[28]), .Z(n4199) );
  NANDN U4998 ( .A(n4257), .B(n6133), .Z(n6132) );
  NANDN U4999 ( .A(n4259), .B(n6134), .Z(n6133) );
  NANDN U5000 ( .A(n4496), .B(n6135), .Z(n6134) );
  NAND U5001 ( .A(n4733), .B(n4499), .Z(n6135) );
  AND U5002 ( .A(n6136), .B(n6137), .Z(n4499) );
  AND U5003 ( .A(n4673), .B(n4619), .Z(n6137) );
  OR U5004 ( .A(B[20]), .B(A[20]), .Z(n4673) );
  AND U5005 ( .A(n4556), .B(n4552), .Z(n6136) );
  NANDN U5006 ( .A(n4788), .B(n6138), .Z(n4733) );
  NAND U5007 ( .A(n6139), .B(n4789), .Z(n6138) );
  OR U5008 ( .A(B[19]), .B(A[19]), .Z(n4789) );
  NANDN U5009 ( .A(n4791), .B(n6140), .Z(n6139) );
  NANDN U5010 ( .A(n4792), .B(n6141), .Z(n6140) );
  NANDN U5011 ( .A(n4848), .B(n6142), .Z(n6141) );
  NAND U5012 ( .A(n4851), .B(n4907), .Z(n6142) );
  AND U5013 ( .A(A[16]), .B(B[16]), .Z(n4907) );
  OR U5014 ( .A(B[17]), .B(A[17]), .Z(n4851) );
  AND U5015 ( .A(B[17]), .B(A[17]), .Z(n4848) );
  NOR U5016 ( .A(B[18]), .B(A[18]), .Z(n4792) );
  AND U5017 ( .A(B[18]), .B(A[18]), .Z(n4791) );
  AND U5018 ( .A(B[19]), .B(A[19]), .Z(n4788) );
  NANDN U5019 ( .A(n4551), .B(n6143), .Z(n4496) );
  NAND U5020 ( .A(n6144), .B(n4552), .Z(n6143) );
  OR U5021 ( .A(B[23]), .B(A[23]), .Z(n4552) );
  NANDN U5022 ( .A(n4554), .B(n6145), .Z(n6144) );
  NAND U5023 ( .A(n6146), .B(n4556), .Z(n6145) );
  OR U5024 ( .A(B[22]), .B(A[22]), .Z(n4556) );
  NANDN U5025 ( .A(n4616), .B(n6147), .Z(n6146) );
  NAND U5026 ( .A(n4619), .B(n4671), .Z(n6147) );
  AND U5027 ( .A(B[20]), .B(A[20]), .Z(n4671) );
  OR U5028 ( .A(B[21]), .B(A[21]), .Z(n4619) );
  AND U5029 ( .A(B[21]), .B(A[21]), .Z(n4616) );
  AND U5030 ( .A(B[22]), .B(A[22]), .Z(n4554) );
  AND U5031 ( .A(B[23]), .B(A[23]), .Z(n4551) );
  NAND U5032 ( .A(n6148), .B(n6149), .Z(n4259) );
  AND U5033 ( .A(n4440), .B(n4383), .Z(n6149) );
  OR U5034 ( .A(B[24]), .B(A[24]), .Z(n4440) );
  AND U5035 ( .A(n4322), .B(n4318), .Z(n6148) );
  NANDN U5036 ( .A(n4317), .B(n6150), .Z(n4257) );
  NAND U5037 ( .A(n6151), .B(n4318), .Z(n6150) );
  OR U5038 ( .A(B[27]), .B(A[27]), .Z(n4318) );
  NANDN U5039 ( .A(n4320), .B(n6152), .Z(n6151) );
  NAND U5040 ( .A(n6153), .B(n4322), .Z(n6152) );
  OR U5041 ( .A(B[26]), .B(A[26]), .Z(n4322) );
  NANDN U5042 ( .A(n4380), .B(n6154), .Z(n6153) );
  NAND U5043 ( .A(n4383), .B(n4438), .Z(n6154) );
  AND U5044 ( .A(B[24]), .B(A[24]), .Z(n4438) );
  OR U5045 ( .A(B[25]), .B(A[25]), .Z(n4383) );
  AND U5046 ( .A(B[25]), .B(A[25]), .Z(n4380) );
  AND U5047 ( .A(B[26]), .B(A[26]), .Z(n4320) );
  AND U5048 ( .A(B[27]), .B(A[27]), .Z(n4317) );
  NOR U5049 ( .A(B[29]), .B(A[29]), .Z(n4139) );
  AND U5050 ( .A(B[29]), .B(A[29]), .Z(n4137) );
  NOR U5051 ( .A(B[30]), .B(A[30]), .Z(n4076) );
  AND U5052 ( .A(B[30]), .B(A[30]), .Z(n4075) );
  NOR U5053 ( .A(B[31]), .B(A[31]), .Z(n4072) );
  NOR U5054 ( .A(n3780), .B(n3294), .Z(n6101) );
  NAND U5055 ( .A(n6155), .B(n6156), .Z(n3780) );
  AND U5056 ( .A(n3961), .B(n3904), .Z(n6156) );
  OR U5057 ( .A(B[32]), .B(A[32]), .Z(n3961) );
  ANDN U5058 ( .B(n3839), .A(n3842), .Z(n6155) );
  ANDN U5059 ( .B(n6157), .A(n3231), .Z(n6099) );
  AND U5060 ( .A(B[44]), .B(A[44]), .Z(n3231) );
  NAND U5061 ( .A(n6158), .B(n3234), .Z(n6157) );
  OR U5062 ( .A(A[44]), .B(B[44]), .Z(n3234) );
  NANDN U5063 ( .A(n3292), .B(n6159), .Z(n6158) );
  NANDN U5064 ( .A(n3294), .B(n6160), .Z(n6159) );
  NANDN U5065 ( .A(n3536), .B(n6161), .Z(n6160) );
  NAND U5066 ( .A(n3779), .B(n3539), .Z(n6161) );
  AND U5067 ( .A(n6162), .B(n6163), .Z(n3539) );
  AND U5068 ( .A(n3719), .B(n3662), .Z(n6163) );
  OR U5069 ( .A(B[36]), .B(A[36]), .Z(n3719) );
  AND U5070 ( .A(n3599), .B(n3595), .Z(n6162) );
  NANDN U5071 ( .A(n3838), .B(n6164), .Z(n3779) );
  NAND U5072 ( .A(n6165), .B(n3839), .Z(n6164) );
  OR U5073 ( .A(B[35]), .B(A[35]), .Z(n3839) );
  NANDN U5074 ( .A(n3841), .B(n6166), .Z(n6165) );
  NANDN U5075 ( .A(n3842), .B(n6167), .Z(n6166) );
  NANDN U5076 ( .A(n3901), .B(n6168), .Z(n6167) );
  NAND U5077 ( .A(n3904), .B(n3959), .Z(n6168) );
  AND U5078 ( .A(A[32]), .B(B[32]), .Z(n3959) );
  OR U5079 ( .A(B[33]), .B(A[33]), .Z(n3904) );
  AND U5080 ( .A(B[33]), .B(A[33]), .Z(n3901) );
  NOR U5081 ( .A(B[34]), .B(A[34]), .Z(n3842) );
  AND U5082 ( .A(B[34]), .B(A[34]), .Z(n3841) );
  AND U5083 ( .A(B[35]), .B(A[35]), .Z(n3838) );
  NANDN U5084 ( .A(n3594), .B(n6169), .Z(n3536) );
  NAND U5085 ( .A(n6170), .B(n3595), .Z(n6169) );
  OR U5086 ( .A(B[39]), .B(A[39]), .Z(n3595) );
  NANDN U5087 ( .A(n3597), .B(n6171), .Z(n6170) );
  NAND U5088 ( .A(n6172), .B(n3599), .Z(n6171) );
  OR U5089 ( .A(B[38]), .B(A[38]), .Z(n3599) );
  NANDN U5090 ( .A(n3659), .B(n6173), .Z(n6172) );
  NAND U5091 ( .A(n3662), .B(n3717), .Z(n6173) );
  AND U5092 ( .A(B[36]), .B(A[36]), .Z(n3717) );
  OR U5093 ( .A(B[37]), .B(A[37]), .Z(n3662) );
  AND U5094 ( .A(B[37]), .B(A[37]), .Z(n3659) );
  AND U5095 ( .A(B[38]), .B(A[38]), .Z(n3597) );
  AND U5096 ( .A(B[39]), .B(A[39]), .Z(n3594) );
  NAND U5097 ( .A(n6174), .B(n6175), .Z(n3294) );
  AND U5098 ( .A(n3476), .B(n3419), .Z(n6175) );
  OR U5099 ( .A(B[40]), .B(A[40]), .Z(n3476) );
  AND U5100 ( .A(n3357), .B(n3353), .Z(n6174) );
  NANDN U5101 ( .A(n3352), .B(n6176), .Z(n3292) );
  NAND U5102 ( .A(n6177), .B(n3353), .Z(n6176) );
  OR U5103 ( .A(B[43]), .B(A[43]), .Z(n3353) );
  NANDN U5104 ( .A(n3355), .B(n6178), .Z(n6177) );
  NAND U5105 ( .A(n6179), .B(n3357), .Z(n6178) );
  OR U5106 ( .A(B[42]), .B(A[42]), .Z(n3357) );
  NANDN U5107 ( .A(n3416), .B(n6180), .Z(n6179) );
  NAND U5108 ( .A(n3419), .B(n3474), .Z(n6180) );
  AND U5109 ( .A(B[40]), .B(A[40]), .Z(n3474) );
  OR U5110 ( .A(B[41]), .B(A[41]), .Z(n3419) );
  AND U5111 ( .A(B[41]), .B(A[41]), .Z(n3416) );
  AND U5112 ( .A(B[42]), .B(A[42]), .Z(n3355) );
  AND U5113 ( .A(B[43]), .B(A[43]), .Z(n3352) );
  NOR U5114 ( .A(B[45]), .B(A[45]), .Z(n3175) );
  AND U5115 ( .A(B[45]), .B(A[45]), .Z(n3173) );
  NOR U5116 ( .A(B[46]), .B(A[46]), .Z(n3112) );
  AND U5117 ( .A(B[46]), .B(A[46]), .Z(n3111) );
  NOR U5118 ( .A(B[47]), .B(A[47]), .Z(n3108) );
  OR U5119 ( .A(B[51]), .B(A[51]), .Z(n2870) );
  NAND U5120 ( .A(n6181), .B(n6182), .Z(n2571) );
  AND U5121 ( .A(n2753), .B(n2696), .Z(n6182) );
  OR U5122 ( .A(A[52]), .B(B[52]), .Z(n2753) );
  AND U5123 ( .A(n2633), .B(n2629), .Z(n6181) );
  NANDN U5124 ( .A(n2628), .B(n6183), .Z(n2569) );
  NAND U5125 ( .A(n6184), .B(n2629), .Z(n6183) );
  OR U5126 ( .A(B[55]), .B(A[55]), .Z(n2629) );
  NANDN U5127 ( .A(n2631), .B(n6185), .Z(n6184) );
  NAND U5128 ( .A(n6186), .B(n2633), .Z(n6185) );
  OR U5129 ( .A(A[54]), .B(B[54]), .Z(n2633) );
  NANDN U5130 ( .A(n2693), .B(n6187), .Z(n6186) );
  NAND U5131 ( .A(n2696), .B(n2751), .Z(n6187) );
  AND U5132 ( .A(A[52]), .B(B[52]), .Z(n2751) );
  OR U5133 ( .A(A[53]), .B(B[53]), .Z(n2696) );
  AND U5134 ( .A(A[53]), .B(B[53]), .Z(n2693) );
  AND U5135 ( .A(A[54]), .B(B[54]), .Z(n2631) );
  AND U5136 ( .A(B[55]), .B(A[55]), .Z(n2628) );
  NAND U5137 ( .A(n6188), .B(n6189), .Z(n2327) );
  AND U5138 ( .A(n2511), .B(n2454), .Z(n6189) );
  OR U5139 ( .A(B[56]), .B(A[56]), .Z(n2511) );
  AND U5140 ( .A(n2394), .B(n2390), .Z(n6188) );
  NANDN U5141 ( .A(n2389), .B(n6190), .Z(n2325) );
  NAND U5142 ( .A(n6191), .B(n2390), .Z(n6190) );
  OR U5143 ( .A(B[59]), .B(A[59]), .Z(n2390) );
  NANDN U5144 ( .A(n2392), .B(n6192), .Z(n6191) );
  NAND U5145 ( .A(n6193), .B(n2394), .Z(n6192) );
  OR U5146 ( .A(B[58]), .B(A[58]), .Z(n2394) );
  NANDN U5147 ( .A(n2451), .B(n6194), .Z(n6193) );
  NAND U5148 ( .A(n2454), .B(n2509), .Z(n6194) );
  AND U5149 ( .A(B[56]), .B(A[56]), .Z(n2509) );
  OR U5150 ( .A(B[57]), .B(A[57]), .Z(n2454) );
  AND U5151 ( .A(B[57]), .B(A[57]), .Z(n2451) );
  AND U5152 ( .A(B[58]), .B(A[58]), .Z(n2392) );
  AND U5153 ( .A(B[59]), .B(A[59]), .Z(n2389) );
  NOR U5154 ( .A(B[60]), .B(A[60]), .Z(n2266) );
  AND U5155 ( .A(B[60]), .B(A[60]), .Z(n2264) );
  NOR U5156 ( .A(B[61]), .B(A[61]), .Z(n2207) );
  AND U5157 ( .A(B[61]), .B(A[61]), .Z(n2205) );
  NOR U5158 ( .A(B[62]), .B(A[62]), .Z(n2144) );
  AND U5159 ( .A(B[62]), .B(A[62]), .Z(n2143) );
  NOR U5160 ( .A(B[63]), .B(A[63]), .Z(n2140) );
  NAND U5161 ( .A(n6195), .B(n6196), .Z(n6071) );
  AND U5162 ( .A(n6197), .B(n6198), .Z(n6196) );
  ANDN U5163 ( .B(n1245), .A(n1299), .Z(n6198) );
  ANDN U5164 ( .B(n1178), .A(n1181), .Z(n6197) );
  ANDN U5165 ( .B(n6199), .A(n1846), .Z(n6195) );
  NAND U5166 ( .A(n6200), .B(n6201), .Z(n1846) );
  AND U5167 ( .A(n2027), .B(n1970), .Z(n6201) );
  OR U5168 ( .A(B[64]), .B(A[64]), .Z(n2027) );
  ANDN U5169 ( .B(n1905), .A(n1908), .Z(n6200) );
  ANDN U5170 ( .B(n1602), .A(n1361), .Z(n6199) );
  NANDN U5171 ( .A(n1177), .B(n6202), .Z(n5430) );
  NAND U5172 ( .A(n6203), .B(n1178), .Z(n6202) );
  OR U5173 ( .A(B[79]), .B(A[79]), .Z(n1178) );
  NANDN U5174 ( .A(n1180), .B(n6204), .Z(n6203) );
  NANDN U5175 ( .A(n1181), .B(n6205), .Z(n6204) );
  NANDN U5176 ( .A(n1242), .B(n6206), .Z(n6205) );
  NAND U5177 ( .A(n6207), .B(n1245), .Z(n6206) );
  OR U5178 ( .A(B[77]), .B(A[77]), .Z(n1245) );
  NANDN U5179 ( .A(n1297), .B(n6208), .Z(n6207) );
  NANDN U5180 ( .A(n1299), .B(n6209), .Z(n6208) );
  NANDN U5181 ( .A(n1359), .B(n6210), .Z(n6209) );
  NANDN U5182 ( .A(n1361), .B(n6211), .Z(n6210) );
  NANDN U5183 ( .A(n1599), .B(n6212), .Z(n6211) );
  NAND U5184 ( .A(n1845), .B(n1602), .Z(n6212) );
  AND U5185 ( .A(n6213), .B(n6214), .Z(n1602) );
  AND U5186 ( .A(n1785), .B(n1725), .Z(n6214) );
  OR U5187 ( .A(B[68]), .B(A[68]), .Z(n1785) );
  AND U5188 ( .A(n1662), .B(n1658), .Z(n6213) );
  NANDN U5189 ( .A(n1904), .B(n6215), .Z(n1845) );
  NAND U5190 ( .A(n6216), .B(n1905), .Z(n6215) );
  OR U5191 ( .A(B[67]), .B(A[67]), .Z(n1905) );
  NANDN U5192 ( .A(n1907), .B(n6217), .Z(n6216) );
  NANDN U5193 ( .A(n1908), .B(n6218), .Z(n6217) );
  NANDN U5194 ( .A(n1967), .B(n6219), .Z(n6218) );
  NAND U5195 ( .A(n1970), .B(n2025), .Z(n6219) );
  AND U5196 ( .A(A[64]), .B(B[64]), .Z(n2025) );
  OR U5197 ( .A(B[65]), .B(A[65]), .Z(n1970) );
  AND U5198 ( .A(B[65]), .B(A[65]), .Z(n1967) );
  NOR U5199 ( .A(B[66]), .B(A[66]), .Z(n1908) );
  AND U5200 ( .A(B[66]), .B(A[66]), .Z(n1907) );
  AND U5201 ( .A(B[67]), .B(A[67]), .Z(n1904) );
  NANDN U5202 ( .A(n1657), .B(n6220), .Z(n1599) );
  NAND U5203 ( .A(n6221), .B(n1658), .Z(n6220) );
  OR U5204 ( .A(B[71]), .B(A[71]), .Z(n1658) );
  NANDN U5205 ( .A(n1660), .B(n6222), .Z(n6221) );
  NAND U5206 ( .A(n6223), .B(n1662), .Z(n6222) );
  OR U5207 ( .A(B[70]), .B(A[70]), .Z(n1662) );
  NANDN U5208 ( .A(n1722), .B(n6224), .Z(n6223) );
  NAND U5209 ( .A(n1725), .B(n1783), .Z(n6224) );
  AND U5210 ( .A(B[68]), .B(A[68]), .Z(n1783) );
  OR U5211 ( .A(B[69]), .B(A[69]), .Z(n1725) );
  AND U5212 ( .A(B[69]), .B(A[69]), .Z(n1722) );
  AND U5213 ( .A(B[70]), .B(A[70]), .Z(n1660) );
  AND U5214 ( .A(B[71]), .B(A[71]), .Z(n1657) );
  NAND U5215 ( .A(n6225), .B(n6226), .Z(n1361) );
  AND U5216 ( .A(n1539), .B(n1482), .Z(n6226) );
  OR U5217 ( .A(B[72]), .B(A[72]), .Z(n1539) );
  AND U5218 ( .A(n1420), .B(n1416), .Z(n6225) );
  NANDN U5219 ( .A(n1415), .B(n6227), .Z(n1359) );
  NAND U5220 ( .A(n6228), .B(n1416), .Z(n6227) );
  OR U5221 ( .A(B[75]), .B(A[75]), .Z(n1416) );
  NANDN U5222 ( .A(n1418), .B(n6229), .Z(n6228) );
  NAND U5223 ( .A(n6230), .B(n1420), .Z(n6229) );
  OR U5224 ( .A(B[74]), .B(A[74]), .Z(n1420) );
  NANDN U5225 ( .A(n1479), .B(n6231), .Z(n6230) );
  NAND U5226 ( .A(n1482), .B(n1537), .Z(n6231) );
  AND U5227 ( .A(B[72]), .B(A[72]), .Z(n1537) );
  OR U5228 ( .A(B[73]), .B(A[73]), .Z(n1482) );
  AND U5229 ( .A(B[73]), .B(A[73]), .Z(n1479) );
  AND U5230 ( .A(B[74]), .B(A[74]), .Z(n1418) );
  AND U5231 ( .A(B[75]), .B(A[75]), .Z(n1415) );
  NOR U5232 ( .A(B[76]), .B(A[76]), .Z(n1299) );
  AND U5233 ( .A(B[76]), .B(A[76]), .Z(n1297) );
  AND U5234 ( .A(B[77]), .B(A[77]), .Z(n1242) );
  NOR U5235 ( .A(B[78]), .B(A[78]), .Z(n1181) );
  AND U5236 ( .A(B[78]), .B(A[78]), .Z(n1180) );
  AND U5237 ( .A(B[79]), .B(A[79]), .Z(n1177) );
  NAND U5238 ( .A(n6232), .B(n6233), .Z(n5428) );
  AND U5239 ( .A(n6234), .B(n6235), .Z(n6233) );
  ANDN U5240 ( .B(n300), .A(n354), .Z(n6235) );
  ANDN U5241 ( .B(n233), .A(n236), .Z(n6234) );
  ANDN U5242 ( .B(n6236), .A(n889), .Z(n6232) );
  NAND U5243 ( .A(n6237), .B(n6238), .Z(n889) );
  AND U5244 ( .A(n1064), .B(n1006), .Z(n6238) );
  OR U5245 ( .A(B[80]), .B(A[80]), .Z(n1064) );
  ANDN U5246 ( .B(n944), .A(n947), .Z(n6237) );
  ANDN U5247 ( .B(n654), .A(n416), .Z(n6236) );
  NANDN U5248 ( .A(n232), .B(n6239), .Z(n5427) );
  NAND U5249 ( .A(n6240), .B(n233), .Z(n6239) );
  OR U5250 ( .A(B[95]), .B(A[95]), .Z(n233) );
  NANDN U5251 ( .A(n235), .B(n6241), .Z(n6240) );
  NANDN U5252 ( .A(n236), .B(n6242), .Z(n6241) );
  NANDN U5253 ( .A(n297), .B(n6243), .Z(n6242) );
  NAND U5254 ( .A(n6244), .B(n300), .Z(n6243) );
  OR U5255 ( .A(B[93]), .B(A[93]), .Z(n300) );
  NANDN U5256 ( .A(n352), .B(n6245), .Z(n6244) );
  NANDN U5257 ( .A(n354), .B(n6246), .Z(n6245) );
  NANDN U5258 ( .A(n414), .B(n6247), .Z(n6246) );
  NANDN U5259 ( .A(n416), .B(n6248), .Z(n6247) );
  NANDN U5260 ( .A(n651), .B(n6249), .Z(n6248) );
  NAND U5261 ( .A(n888), .B(n654), .Z(n6249) );
  AND U5262 ( .A(n6250), .B(n6251), .Z(n654) );
  AND U5263 ( .A(n828), .B(n774), .Z(n6251) );
  OR U5264 ( .A(B[84]), .B(A[84]), .Z(n828) );
  AND U5265 ( .A(n711), .B(n707), .Z(n6250) );
  NANDN U5266 ( .A(n943), .B(n6252), .Z(n888) );
  NAND U5267 ( .A(n6253), .B(n944), .Z(n6252) );
  OR U5268 ( .A(B[83]), .B(A[83]), .Z(n944) );
  NANDN U5269 ( .A(n946), .B(n6254), .Z(n6253) );
  NANDN U5270 ( .A(n947), .B(n6255), .Z(n6254) );
  NANDN U5271 ( .A(n1003), .B(n6256), .Z(n6255) );
  NAND U5272 ( .A(n1006), .B(n1062), .Z(n6256) );
  AND U5273 ( .A(A[80]), .B(B[80]), .Z(n1062) );
  OR U5274 ( .A(B[81]), .B(A[81]), .Z(n1006) );
  AND U5275 ( .A(B[81]), .B(A[81]), .Z(n1003) );
  NOR U5276 ( .A(B[82]), .B(A[82]), .Z(n947) );
  AND U5277 ( .A(B[82]), .B(A[82]), .Z(n946) );
  AND U5278 ( .A(B[83]), .B(A[83]), .Z(n943) );
  NANDN U5279 ( .A(n706), .B(n6257), .Z(n651) );
  NAND U5280 ( .A(n6258), .B(n707), .Z(n6257) );
  OR U5281 ( .A(B[87]), .B(A[87]), .Z(n707) );
  NANDN U5282 ( .A(n709), .B(n6259), .Z(n6258) );
  NAND U5283 ( .A(n6260), .B(n711), .Z(n6259) );
  OR U5284 ( .A(B[86]), .B(A[86]), .Z(n711) );
  NANDN U5285 ( .A(n771), .B(n6261), .Z(n6260) );
  NAND U5286 ( .A(n774), .B(n826), .Z(n6261) );
  AND U5287 ( .A(B[84]), .B(A[84]), .Z(n826) );
  OR U5288 ( .A(B[85]), .B(A[85]), .Z(n774) );
  AND U5289 ( .A(B[85]), .B(A[85]), .Z(n771) );
  AND U5290 ( .A(B[86]), .B(A[86]), .Z(n709) );
  AND U5291 ( .A(B[87]), .B(A[87]), .Z(n706) );
  NAND U5292 ( .A(n6262), .B(n6263), .Z(n416) );
  AND U5293 ( .A(n595), .B(n533), .Z(n6263) );
  OR U5294 ( .A(B[88]), .B(A[88]), .Z(n595) );
  AND U5295 ( .A(n475), .B(n471), .Z(n6262) );
  NANDN U5296 ( .A(n470), .B(n6264), .Z(n414) );
  NAND U5297 ( .A(n6265), .B(n471), .Z(n6264) );
  OR U5298 ( .A(B[91]), .B(A[91]), .Z(n471) );
  NANDN U5299 ( .A(n473), .B(n6266), .Z(n6265) );
  NAND U5300 ( .A(n6267), .B(n475), .Z(n6266) );
  OR U5301 ( .A(B[90]), .B(A[90]), .Z(n475) );
  NANDN U5302 ( .A(n530), .B(n6268), .Z(n6267) );
  NAND U5303 ( .A(n533), .B(n593), .Z(n6268) );
  AND U5304 ( .A(B[88]), .B(A[88]), .Z(n593) );
  OR U5305 ( .A(B[89]), .B(A[89]), .Z(n533) );
  AND U5306 ( .A(B[89]), .B(A[89]), .Z(n530) );
  AND U5307 ( .A(B[90]), .B(A[90]), .Z(n473) );
  AND U5308 ( .A(B[91]), .B(A[91]), .Z(n470) );
  NOR U5309 ( .A(B[92]), .B(A[92]), .Z(n354) );
  AND U5310 ( .A(B[92]), .B(A[92]), .Z(n352) );
  AND U5311 ( .A(B[93]), .B(A[93]), .Z(n297) );
  NOR U5312 ( .A(B[94]), .B(A[94]), .Z(n236) );
  AND U5313 ( .A(B[94]), .B(A[94]), .Z(n235) );
  AND U5314 ( .A(B[95]), .B(A[95]), .Z(n232) );
  NAND U5315 ( .A(n6269), .B(n6270), .Z(n5295) );
  AND U5316 ( .A(n6271), .B(n6272), .Z(n6270) );
  AND U5317 ( .A(n5316), .B(n5308), .Z(n6272) );
  AND U5318 ( .A(n5303), .B(n5299), .Z(n6271) );
  ANDN U5319 ( .B(n6273), .A(n5425), .Z(n6269) );
  NAND U5320 ( .A(n6274), .B(n6275), .Z(n5425) );
  AND U5321 ( .A(n12), .B(n68), .Z(n6275) );
  ANDN U5322 ( .B(n8), .A(n124), .Z(n6274) );
  NOR U5323 ( .A(B[96]), .B(A[96]), .Z(n124) );
  ANDN U5324 ( .B(n5320), .A(n5342), .Z(n6273) );
  NANDN U5325 ( .A(n5298), .B(n6276), .Z(n5293) );
  NAND U5326 ( .A(n6277), .B(n5299), .Z(n6276) );
  OR U5327 ( .A(B[111]), .B(A[111]), .Z(n5299) );
  NANDN U5328 ( .A(n5301), .B(n6278), .Z(n6277) );
  NAND U5329 ( .A(n6279), .B(n5303), .Z(n6278) );
  OR U5330 ( .A(B[110]), .B(A[110]), .Z(n5303) );
  NANDN U5331 ( .A(n5305), .B(n6280), .Z(n6279) );
  NAND U5332 ( .A(n6281), .B(n5308), .Z(n6280) );
  OR U5333 ( .A(B[109]), .B(A[109]), .Z(n5308) );
  NANDN U5334 ( .A(n5313), .B(n6282), .Z(n6281) );
  NAND U5335 ( .A(n6283), .B(n5316), .Z(n6282) );
  OR U5336 ( .A(B[108]), .B(A[108]), .Z(n5316) );
  NANDN U5337 ( .A(n5318), .B(n6284), .Z(n6283) );
  NAND U5338 ( .A(n6285), .B(n5320), .Z(n6284) );
  AND U5339 ( .A(n6286), .B(n6287), .Z(n5320) );
  AND U5340 ( .A(n5338), .B(n5334), .Z(n6287) );
  OR U5341 ( .A(B[104]), .B(A[104]), .Z(n5338) );
  AND U5342 ( .A(n5329), .B(n5325), .Z(n6286) );
  NANDN U5343 ( .A(n5340), .B(n6288), .Z(n6285) );
  NANDN U5344 ( .A(n5342), .B(n5424), .Z(n6288) );
  NANDN U5345 ( .A(n7), .B(n6289), .Z(n5424) );
  NAND U5346 ( .A(n6290), .B(n8), .Z(n6289) );
  OR U5347 ( .A(B[99]), .B(A[99]), .Z(n8) );
  NANDN U5348 ( .A(n10), .B(n6291), .Z(n6290) );
  NAND U5349 ( .A(n6292), .B(n12), .Z(n6291) );
  OR U5350 ( .A(B[98]), .B(A[98]), .Z(n12) );
  NANDN U5351 ( .A(n65), .B(n6293), .Z(n6292) );
  NAND U5352 ( .A(n68), .B(n122), .Z(n6293) );
  AND U5353 ( .A(B[96]), .B(A[96]), .Z(n122) );
  OR U5354 ( .A(B[97]), .B(A[97]), .Z(n68) );
  AND U5355 ( .A(B[97]), .B(A[97]), .Z(n65) );
  AND U5356 ( .A(A[98]), .B(B[98]), .Z(n10) );
  AND U5357 ( .A(B[99]), .B(A[99]), .Z(n7) );
  NAND U5358 ( .A(n6294), .B(n6295), .Z(n5342) );
  AND U5359 ( .A(n5371), .B(n5356), .Z(n6295) );
  OR U5360 ( .A(B[100]), .B(A[100]), .Z(n5371) );
  AND U5361 ( .A(n5351), .B(n5347), .Z(n6294) );
  NANDN U5362 ( .A(n5346), .B(n6296), .Z(n5340) );
  NAND U5363 ( .A(n6297), .B(n5347), .Z(n6296) );
  OR U5364 ( .A(B[103]), .B(A[103]), .Z(n5347) );
  NANDN U5365 ( .A(n5349), .B(n6298), .Z(n6297) );
  NAND U5366 ( .A(n6299), .B(n5351), .Z(n6298) );
  OR U5367 ( .A(B[102]), .B(A[102]), .Z(n5351) );
  NANDN U5368 ( .A(n5353), .B(n6300), .Z(n6299) );
  NAND U5369 ( .A(n5356), .B(n5369), .Z(n6300) );
  AND U5370 ( .A(B[100]), .B(A[100]), .Z(n5369) );
  OR U5371 ( .A(B[101]), .B(A[101]), .Z(n5356) );
  AND U5372 ( .A(B[101]), .B(A[101]), .Z(n5353) );
  AND U5373 ( .A(B[102]), .B(A[102]), .Z(n5349) );
  AND U5374 ( .A(B[103]), .B(A[103]), .Z(n5346) );
  NANDN U5375 ( .A(n5324), .B(n6301), .Z(n5318) );
  NAND U5376 ( .A(n6302), .B(n5325), .Z(n6301) );
  OR U5377 ( .A(B[107]), .B(A[107]), .Z(n5325) );
  NANDN U5378 ( .A(n5327), .B(n6303), .Z(n6302) );
  NAND U5379 ( .A(n6304), .B(n5329), .Z(n6303) );
  OR U5380 ( .A(B[106]), .B(A[106]), .Z(n5329) );
  NANDN U5381 ( .A(n5331), .B(n6305), .Z(n6304) );
  NAND U5382 ( .A(n5334), .B(n5336), .Z(n6305) );
  AND U5383 ( .A(B[104]), .B(A[104]), .Z(n5336) );
  OR U5384 ( .A(B[105]), .B(A[105]), .Z(n5334) );
  AND U5385 ( .A(B[105]), .B(A[105]), .Z(n5331) );
  AND U5386 ( .A(B[106]), .B(A[106]), .Z(n5327) );
  AND U5387 ( .A(B[107]), .B(A[107]), .Z(n5324) );
  AND U5388 ( .A(B[108]), .B(A[108]), .Z(n5313) );
  AND U5389 ( .A(B[109]), .B(A[109]), .Z(n5305) );
  AND U5390 ( .A(B[110]), .B(A[110]), .Z(n5301) );
  AND U5391 ( .A(B[111]), .B(A[111]), .Z(n5298) );
  ANDN U5392 ( .B(n6306), .A(n5273), .Z(n6062) );
  NAND U5393 ( .A(n6307), .B(n6308), .Z(n5273) );
  AND U5394 ( .A(n5291), .B(n5287), .Z(n6308) );
  OR U5395 ( .A(B[112]), .B(A[112]), .Z(n5291) );
  ANDN U5396 ( .B(n5278), .A(n5281), .Z(n6307) );
  ANDN U5397 ( .B(n5244), .A(n5221), .Z(n6306) );
  ANDN U5398 ( .B(n6309), .A(n5205), .Z(n6060) );
  AND U5399 ( .A(B[126]), .B(A[126]), .Z(n5205) );
  NAND U5400 ( .A(n6310), .B(n5207), .Z(n6309) );
  OR U5401 ( .A(A[126]), .B(B[126]), .Z(n5207) );
  NANDN U5402 ( .A(n5209), .B(n6311), .Z(n6310) );
  NAND U5403 ( .A(n6312), .B(n5212), .Z(n6311) );
  OR U5404 ( .A(B[125]), .B(A[125]), .Z(n5212) );
  NANDN U5405 ( .A(n5214), .B(n6313), .Z(n6312) );
  NANDN U5406 ( .A(n5216), .B(n6314), .Z(n6313) );
  NANDN U5407 ( .A(n5219), .B(n6315), .Z(n6314) );
  NANDN U5408 ( .A(n5221), .B(n6316), .Z(n6315) );
  NANDN U5409 ( .A(n5241), .B(n6317), .Z(n6316) );
  NAND U5410 ( .A(n5272), .B(n5244), .Z(n6317) );
  AND U5411 ( .A(n6318), .B(n6319), .Z(n5244) );
  AND U5412 ( .A(n5269), .B(n5265), .Z(n6319) );
  OR U5413 ( .A(B[116]), .B(A[116]), .Z(n5269) );
  AND U5414 ( .A(n5260), .B(n5256), .Z(n6318) );
  NANDN U5415 ( .A(n5277), .B(n6320), .Z(n5272) );
  NAND U5416 ( .A(n6321), .B(n5278), .Z(n6320) );
  OR U5417 ( .A(B[115]), .B(A[115]), .Z(n5278) );
  NANDN U5418 ( .A(n5280), .B(n6322), .Z(n6321) );
  NANDN U5419 ( .A(n5281), .B(n6323), .Z(n6322) );
  NANDN U5420 ( .A(n5284), .B(n6324), .Z(n6323) );
  NAND U5421 ( .A(n5287), .B(n5289), .Z(n6324) );
  AND U5422 ( .A(A[112]), .B(B[112]), .Z(n5289) );
  OR U5423 ( .A(B[113]), .B(A[113]), .Z(n5287) );
  AND U5424 ( .A(B[113]), .B(A[113]), .Z(n5284) );
  NOR U5425 ( .A(B[114]), .B(A[114]), .Z(n5281) );
  AND U5426 ( .A(B[114]), .B(A[114]), .Z(n5280) );
  AND U5427 ( .A(B[115]), .B(A[115]), .Z(n5277) );
  NANDN U5428 ( .A(n5255), .B(n6325), .Z(n5241) );
  NAND U5429 ( .A(n6326), .B(n5256), .Z(n6325) );
  OR U5430 ( .A(B[119]), .B(A[119]), .Z(n5256) );
  NANDN U5431 ( .A(n5258), .B(n6327), .Z(n6326) );
  NAND U5432 ( .A(n6328), .B(n5260), .Z(n6327) );
  OR U5433 ( .A(B[118]), .B(A[118]), .Z(n5260) );
  NANDN U5434 ( .A(n5262), .B(n6329), .Z(n6328) );
  NAND U5435 ( .A(n5265), .B(n5267), .Z(n6329) );
  AND U5436 ( .A(B[116]), .B(A[116]), .Z(n5267) );
  OR U5437 ( .A(B[117]), .B(A[117]), .Z(n5265) );
  AND U5438 ( .A(B[117]), .B(A[117]), .Z(n5262) );
  AND U5439 ( .A(B[118]), .B(A[118]), .Z(n5258) );
  AND U5440 ( .A(B[119]), .B(A[119]), .Z(n5255) );
  NAND U5441 ( .A(n6330), .B(n6331), .Z(n5221) );
  AND U5442 ( .A(n5239), .B(n5235), .Z(n6331) );
  OR U5443 ( .A(B[120]), .B(A[120]), .Z(n5239) );
  AND U5444 ( .A(n5230), .B(n5226), .Z(n6330) );
  NANDN U5445 ( .A(n5225), .B(n6332), .Z(n5219) );
  NAND U5446 ( .A(n6333), .B(n5226), .Z(n6332) );
  OR U5447 ( .A(B[123]), .B(A[123]), .Z(n5226) );
  NANDN U5448 ( .A(n5228), .B(n6334), .Z(n6333) );
  NAND U5449 ( .A(n6335), .B(n5230), .Z(n6334) );
  OR U5450 ( .A(B[122]), .B(A[122]), .Z(n5230) );
  NANDN U5451 ( .A(n5232), .B(n6336), .Z(n6335) );
  NAND U5452 ( .A(n5235), .B(n5237), .Z(n6336) );
  AND U5453 ( .A(B[120]), .B(A[120]), .Z(n5237) );
  OR U5454 ( .A(B[121]), .B(A[121]), .Z(n5235) );
  AND U5455 ( .A(B[121]), .B(A[121]), .Z(n5232) );
  AND U5456 ( .A(B[122]), .B(A[122]), .Z(n5228) );
  AND U5457 ( .A(B[123]), .B(A[123]), .Z(n5225) );
  NOR U5458 ( .A(B[124]), .B(A[124]), .Z(n5216) );
  AND U5459 ( .A(B[124]), .B(A[124]), .Z(n5214) );
  AND U5460 ( .A(B[125]), .B(A[125]), .Z(n5209) );
  NOR U5461 ( .A(B[127]), .B(A[127]), .Z(n5202) );
  NAND U5462 ( .A(n6337), .B(n6338), .Z(n6057) );
  AND U5463 ( .A(n6339), .B(n6340), .Z(n6338) );
  AND U5464 ( .A(n5124), .B(n5119), .Z(n6340) );
  AND U5465 ( .A(n5114), .B(n5110), .Z(n6339) );
  ANDN U5466 ( .B(n6341), .A(n5176), .Z(n6337) );
  NAND U5467 ( .A(n6342), .B(n6343), .Z(n5176) );
  AND U5468 ( .A(n5198), .B(n5190), .Z(n6343) );
  OR U5469 ( .A(B[128]), .B(A[128]), .Z(n5198) );
  AND U5470 ( .A(n5185), .B(n5181), .Z(n6342) );
  ANDN U5471 ( .B(n5128), .A(n5154), .Z(n6341) );
  NANDN U5472 ( .A(n5109), .B(n6344), .Z(n6055) );
  NAND U5473 ( .A(n6345), .B(n5110), .Z(n6344) );
  OR U5474 ( .A(B[143]), .B(A[143]), .Z(n5110) );
  NANDN U5475 ( .A(n5112), .B(n6346), .Z(n6345) );
  NAND U5476 ( .A(n6347), .B(n5114), .Z(n6346) );
  OR U5477 ( .A(B[142]), .B(A[142]), .Z(n5114) );
  NANDN U5478 ( .A(n5116), .B(n6348), .Z(n6347) );
  NAND U5479 ( .A(n6349), .B(n5119), .Z(n6348) );
  OR U5480 ( .A(B[141]), .B(A[141]), .Z(n5119) );
  NANDN U5481 ( .A(n5121), .B(n6350), .Z(n6349) );
  NAND U5482 ( .A(n6351), .B(n5124), .Z(n6350) );
  OR U5483 ( .A(B[140]), .B(A[140]), .Z(n5124) );
  NANDN U5484 ( .A(n5126), .B(n6352), .Z(n6351) );
  NAND U5485 ( .A(n6353), .B(n5128), .Z(n6352) );
  AND U5486 ( .A(n6354), .B(n6355), .Z(n5128) );
  AND U5487 ( .A(n5150), .B(n5146), .Z(n6355) );
  OR U5488 ( .A(B[136]), .B(A[136]), .Z(n5150) );
  AND U5489 ( .A(n5141), .B(n5137), .Z(n6354) );
  NANDN U5490 ( .A(n5152), .B(n6356), .Z(n6353) );
  NANDN U5491 ( .A(n5154), .B(n5175), .Z(n6356) );
  NANDN U5492 ( .A(n5180), .B(n6357), .Z(n5175) );
  NAND U5493 ( .A(n6358), .B(n5181), .Z(n6357) );
  OR U5494 ( .A(B[131]), .B(A[131]), .Z(n5181) );
  NANDN U5495 ( .A(n5183), .B(n6359), .Z(n6358) );
  NAND U5496 ( .A(n6360), .B(n5185), .Z(n6359) );
  OR U5497 ( .A(B[130]), .B(A[130]), .Z(n5185) );
  NANDN U5498 ( .A(n5187), .B(n6361), .Z(n6360) );
  NAND U5499 ( .A(n5190), .B(n5196), .Z(n6361) );
  AND U5500 ( .A(B[128]), .B(A[128]), .Z(n5196) );
  OR U5501 ( .A(B[129]), .B(A[129]), .Z(n5190) );
  AND U5502 ( .A(B[129]), .B(A[129]), .Z(n5187) );
  AND U5503 ( .A(B[130]), .B(A[130]), .Z(n5183) );
  AND U5504 ( .A(B[131]), .B(A[131]), .Z(n5180) );
  NAND U5505 ( .A(n6362), .B(n6363), .Z(n5154) );
  AND U5506 ( .A(n5172), .B(n5168), .Z(n6363) );
  OR U5507 ( .A(B[132]), .B(A[132]), .Z(n5172) );
  AND U5508 ( .A(n5163), .B(n5159), .Z(n6362) );
  NANDN U5509 ( .A(n5158), .B(n6364), .Z(n5152) );
  NAND U5510 ( .A(n6365), .B(n5159), .Z(n6364) );
  OR U5511 ( .A(B[135]), .B(A[135]), .Z(n5159) );
  NANDN U5512 ( .A(n5161), .B(n6366), .Z(n6365) );
  NAND U5513 ( .A(n6367), .B(n5163), .Z(n6366) );
  OR U5514 ( .A(B[134]), .B(A[134]), .Z(n5163) );
  NANDN U5515 ( .A(n5165), .B(n6368), .Z(n6367) );
  NAND U5516 ( .A(n5168), .B(n5170), .Z(n6368) );
  AND U5517 ( .A(B[132]), .B(A[132]), .Z(n5170) );
  OR U5518 ( .A(B[133]), .B(A[133]), .Z(n5168) );
  AND U5519 ( .A(B[133]), .B(A[133]), .Z(n5165) );
  AND U5520 ( .A(B[134]), .B(A[134]), .Z(n5161) );
  AND U5521 ( .A(B[135]), .B(A[135]), .Z(n5158) );
  NANDN U5522 ( .A(n5136), .B(n6369), .Z(n5126) );
  NAND U5523 ( .A(n6370), .B(n5137), .Z(n6369) );
  OR U5524 ( .A(B[139]), .B(A[139]), .Z(n5137) );
  NANDN U5525 ( .A(n5139), .B(n6371), .Z(n6370) );
  NAND U5526 ( .A(n6372), .B(n5141), .Z(n6371) );
  OR U5527 ( .A(B[138]), .B(A[138]), .Z(n5141) );
  NANDN U5528 ( .A(n5143), .B(n6373), .Z(n6372) );
  NAND U5529 ( .A(n5146), .B(n5148), .Z(n6373) );
  AND U5530 ( .A(B[136]), .B(A[136]), .Z(n5148) );
  OR U5531 ( .A(B[137]), .B(A[137]), .Z(n5146) );
  AND U5532 ( .A(B[137]), .B(A[137]), .Z(n5143) );
  AND U5533 ( .A(B[138]), .B(A[138]), .Z(n5139) );
  AND U5534 ( .A(B[139]), .B(A[139]), .Z(n5136) );
  AND U5535 ( .A(B[140]), .B(A[140]), .Z(n5121) );
  AND U5536 ( .A(B[141]), .B(A[141]), .Z(n5116) );
  AND U5537 ( .A(B[142]), .B(A[142]), .Z(n5112) );
  AND U5538 ( .A(B[143]), .B(A[143]), .Z(n5109) );
  NAND U5539 ( .A(n6374), .B(n6375), .Z(n6054) );
  AND U5540 ( .A(n6376), .B(n6377), .Z(n6375) );
  AND U5541 ( .A(n5035), .B(n5030), .Z(n6377) );
  AND U5542 ( .A(n5025), .B(n5021), .Z(n6376) );
  ANDN U5543 ( .B(n6378), .A(n5087), .Z(n6374) );
  NAND U5544 ( .A(n6379), .B(n6380), .Z(n5087) );
  AND U5545 ( .A(n5105), .B(n5101), .Z(n6380) );
  OR U5546 ( .A(B[144]), .B(A[144]), .Z(n5105) );
  AND U5547 ( .A(n5096), .B(n5092), .Z(n6379) );
  ANDN U5548 ( .B(n5039), .A(n5061), .Z(n6378) );
  NANDN U5549 ( .A(n5020), .B(n6381), .Z(n6052) );
  NAND U5550 ( .A(n6382), .B(n5021), .Z(n6381) );
  OR U5551 ( .A(B[159]), .B(A[159]), .Z(n5021) );
  NANDN U5552 ( .A(n5023), .B(n6383), .Z(n6382) );
  NAND U5553 ( .A(n6384), .B(n5025), .Z(n6383) );
  OR U5554 ( .A(B[158]), .B(A[158]), .Z(n5025) );
  NANDN U5555 ( .A(n5027), .B(n6385), .Z(n6384) );
  NAND U5556 ( .A(n6386), .B(n5030), .Z(n6385) );
  OR U5557 ( .A(B[157]), .B(A[157]), .Z(n5030) );
  NANDN U5558 ( .A(n5032), .B(n6387), .Z(n6386) );
  NAND U5559 ( .A(n6388), .B(n5035), .Z(n6387) );
  OR U5560 ( .A(B[156]), .B(A[156]), .Z(n5035) );
  NANDN U5561 ( .A(n5037), .B(n6389), .Z(n6388) );
  NAND U5562 ( .A(n6390), .B(n5039), .Z(n6389) );
  AND U5563 ( .A(n6391), .B(n6392), .Z(n5039) );
  AND U5564 ( .A(n5057), .B(n5053), .Z(n6392) );
  OR U5565 ( .A(B[152]), .B(A[152]), .Z(n5057) );
  AND U5566 ( .A(n5048), .B(n5044), .Z(n6391) );
  NANDN U5567 ( .A(n5059), .B(n6393), .Z(n6390) );
  NANDN U5568 ( .A(n5061), .B(n5086), .Z(n6393) );
  NANDN U5569 ( .A(n5091), .B(n6394), .Z(n5086) );
  NAND U5570 ( .A(n6395), .B(n5092), .Z(n6394) );
  OR U5571 ( .A(B[147]), .B(A[147]), .Z(n5092) );
  NANDN U5572 ( .A(n5094), .B(n6396), .Z(n6395) );
  NAND U5573 ( .A(n6397), .B(n5096), .Z(n6396) );
  OR U5574 ( .A(B[146]), .B(A[146]), .Z(n5096) );
  NANDN U5575 ( .A(n5098), .B(n6398), .Z(n6397) );
  NAND U5576 ( .A(n5101), .B(n5103), .Z(n6398) );
  AND U5577 ( .A(B[144]), .B(A[144]), .Z(n5103) );
  OR U5578 ( .A(B[145]), .B(A[145]), .Z(n5101) );
  AND U5579 ( .A(B[145]), .B(A[145]), .Z(n5098) );
  AND U5580 ( .A(B[146]), .B(A[146]), .Z(n5094) );
  AND U5581 ( .A(B[147]), .B(A[147]), .Z(n5091) );
  NAND U5582 ( .A(n6399), .B(n6400), .Z(n5061) );
  AND U5583 ( .A(n5083), .B(n5075), .Z(n6400) );
  OR U5584 ( .A(B[148]), .B(A[148]), .Z(n5083) );
  AND U5585 ( .A(n5070), .B(n5066), .Z(n6399) );
  NANDN U5586 ( .A(n5065), .B(n6401), .Z(n5059) );
  NAND U5587 ( .A(n6402), .B(n5066), .Z(n6401) );
  OR U5588 ( .A(B[151]), .B(A[151]), .Z(n5066) );
  NANDN U5589 ( .A(n5068), .B(n6403), .Z(n6402) );
  NAND U5590 ( .A(n6404), .B(n5070), .Z(n6403) );
  OR U5591 ( .A(B[150]), .B(A[150]), .Z(n5070) );
  NANDN U5592 ( .A(n5072), .B(n6405), .Z(n6404) );
  NAND U5593 ( .A(n5075), .B(n5081), .Z(n6405) );
  AND U5594 ( .A(B[148]), .B(A[148]), .Z(n5081) );
  OR U5595 ( .A(B[149]), .B(A[149]), .Z(n5075) );
  AND U5596 ( .A(B[149]), .B(A[149]), .Z(n5072) );
  AND U5597 ( .A(B[150]), .B(A[150]), .Z(n5068) );
  AND U5598 ( .A(B[151]), .B(A[151]), .Z(n5065) );
  NANDN U5599 ( .A(n5043), .B(n6406), .Z(n5037) );
  NAND U5600 ( .A(n6407), .B(n5044), .Z(n6406) );
  OR U5601 ( .A(B[155]), .B(A[155]), .Z(n5044) );
  NANDN U5602 ( .A(n5046), .B(n6408), .Z(n6407) );
  NAND U5603 ( .A(n6409), .B(n5048), .Z(n6408) );
  OR U5604 ( .A(B[154]), .B(A[154]), .Z(n5048) );
  NANDN U5605 ( .A(n5050), .B(n6410), .Z(n6409) );
  NAND U5606 ( .A(n5053), .B(n5055), .Z(n6410) );
  AND U5607 ( .A(B[152]), .B(A[152]), .Z(n5055) );
  OR U5608 ( .A(B[153]), .B(A[153]), .Z(n5053) );
  AND U5609 ( .A(B[153]), .B(A[153]), .Z(n5050) );
  AND U5610 ( .A(B[154]), .B(A[154]), .Z(n5046) );
  AND U5611 ( .A(B[155]), .B(A[155]), .Z(n5043) );
  AND U5612 ( .A(B[156]), .B(A[156]), .Z(n5032) );
  AND U5613 ( .A(B[157]), .B(A[157]), .Z(n5027) );
  AND U5614 ( .A(B[158]), .B(A[158]), .Z(n5023) );
  AND U5615 ( .A(B[159]), .B(A[159]), .Z(n5020) );
  NAND U5616 ( .A(n6411), .B(n6412), .Z(n6051) );
  AND U5617 ( .A(n6413), .B(n6414), .Z(n6412) );
  AND U5618 ( .A(n4945), .B(n4940), .Z(n6414) );
  AND U5619 ( .A(n4935), .B(n4931), .Z(n6413) );
  ANDN U5620 ( .B(n6415), .A(n4994), .Z(n6411) );
  NAND U5621 ( .A(n6416), .B(n6417), .Z(n4994) );
  AND U5622 ( .A(n5012), .B(n5008), .Z(n6417) );
  OR U5623 ( .A(B[160]), .B(A[160]), .Z(n5012) );
  AND U5624 ( .A(n5003), .B(n4999), .Z(n6416) );
  ANDN U5625 ( .B(n4949), .A(n4972), .Z(n6415) );
  NANDN U5626 ( .A(n4930), .B(n6418), .Z(n6049) );
  NAND U5627 ( .A(n6419), .B(n4931), .Z(n6418) );
  OR U5628 ( .A(B[175]), .B(A[175]), .Z(n4931) );
  NANDN U5629 ( .A(n4933), .B(n6420), .Z(n6419) );
  NAND U5630 ( .A(n6421), .B(n4935), .Z(n6420) );
  OR U5631 ( .A(B[174]), .B(A[174]), .Z(n4935) );
  NANDN U5632 ( .A(n4937), .B(n6422), .Z(n6421) );
  NAND U5633 ( .A(n6423), .B(n4940), .Z(n6422) );
  OR U5634 ( .A(B[173]), .B(A[173]), .Z(n4940) );
  NANDN U5635 ( .A(n4942), .B(n6424), .Z(n6423) );
  NAND U5636 ( .A(n6425), .B(n4945), .Z(n6424) );
  OR U5637 ( .A(B[172]), .B(A[172]), .Z(n4945) );
  NANDN U5638 ( .A(n4947), .B(n6426), .Z(n6425) );
  NAND U5639 ( .A(n6427), .B(n4949), .Z(n6426) );
  AND U5640 ( .A(n6428), .B(n6429), .Z(n4949) );
  AND U5641 ( .A(n4968), .B(n4963), .Z(n6429) );
  OR U5642 ( .A(B[168]), .B(A[168]), .Z(n4968) );
  AND U5643 ( .A(n4958), .B(n4954), .Z(n6428) );
  NANDN U5644 ( .A(n4970), .B(n6430), .Z(n6427) );
  NANDN U5645 ( .A(n4972), .B(n4993), .Z(n6430) );
  NANDN U5646 ( .A(n4998), .B(n6431), .Z(n4993) );
  NAND U5647 ( .A(n6432), .B(n4999), .Z(n6431) );
  OR U5648 ( .A(B[163]), .B(A[163]), .Z(n4999) );
  NANDN U5649 ( .A(n5001), .B(n6433), .Z(n6432) );
  NAND U5650 ( .A(n6434), .B(n5003), .Z(n6433) );
  OR U5651 ( .A(B[162]), .B(A[162]), .Z(n5003) );
  NANDN U5652 ( .A(n5005), .B(n6435), .Z(n6434) );
  NAND U5653 ( .A(n5008), .B(n5010), .Z(n6435) );
  AND U5654 ( .A(B[160]), .B(A[160]), .Z(n5010) );
  OR U5655 ( .A(B[161]), .B(A[161]), .Z(n5008) );
  AND U5656 ( .A(B[161]), .B(A[161]), .Z(n5005) );
  AND U5657 ( .A(B[162]), .B(A[162]), .Z(n5001) );
  AND U5658 ( .A(B[163]), .B(A[163]), .Z(n4998) );
  NAND U5659 ( .A(n6436), .B(n6437), .Z(n4972) );
  AND U5660 ( .A(n4990), .B(n4986), .Z(n6437) );
  OR U5661 ( .A(B[164]), .B(A[164]), .Z(n4990) );
  AND U5662 ( .A(n4981), .B(n4977), .Z(n6436) );
  NANDN U5663 ( .A(n4976), .B(n6438), .Z(n4970) );
  NAND U5664 ( .A(n6439), .B(n4977), .Z(n6438) );
  OR U5665 ( .A(B[167]), .B(A[167]), .Z(n4977) );
  NANDN U5666 ( .A(n4979), .B(n6440), .Z(n6439) );
  NAND U5667 ( .A(n6441), .B(n4981), .Z(n6440) );
  OR U5668 ( .A(B[166]), .B(A[166]), .Z(n4981) );
  NANDN U5669 ( .A(n4983), .B(n6442), .Z(n6441) );
  NAND U5670 ( .A(n4986), .B(n4988), .Z(n6442) );
  AND U5671 ( .A(B[164]), .B(A[164]), .Z(n4988) );
  OR U5672 ( .A(B[165]), .B(A[165]), .Z(n4986) );
  AND U5673 ( .A(B[165]), .B(A[165]), .Z(n4983) );
  AND U5674 ( .A(B[166]), .B(A[166]), .Z(n4979) );
  AND U5675 ( .A(B[167]), .B(A[167]), .Z(n4976) );
  NANDN U5676 ( .A(n4953), .B(n6443), .Z(n4947) );
  NAND U5677 ( .A(n6444), .B(n4954), .Z(n6443) );
  OR U5678 ( .A(B[171]), .B(A[171]), .Z(n4954) );
  NANDN U5679 ( .A(n4956), .B(n6445), .Z(n6444) );
  NAND U5680 ( .A(n6446), .B(n4958), .Z(n6445) );
  OR U5681 ( .A(B[170]), .B(A[170]), .Z(n4958) );
  NANDN U5682 ( .A(n4960), .B(n6447), .Z(n6446) );
  NAND U5683 ( .A(n4963), .B(n4966), .Z(n6447) );
  AND U5684 ( .A(B[168]), .B(A[168]), .Z(n4966) );
  OR U5685 ( .A(B[169]), .B(A[169]), .Z(n4963) );
  AND U5686 ( .A(B[169]), .B(A[169]), .Z(n4960) );
  AND U5687 ( .A(B[170]), .B(A[170]), .Z(n4956) );
  AND U5688 ( .A(B[171]), .B(A[171]), .Z(n4953) );
  AND U5689 ( .A(B[172]), .B(A[172]), .Z(n4942) );
  AND U5690 ( .A(B[173]), .B(A[173]), .Z(n4937) );
  AND U5691 ( .A(B[174]), .B(A[174]), .Z(n4933) );
  AND U5692 ( .A(B[175]), .B(A[175]), .Z(n4930) );
  ANDN U5693 ( .B(n6448), .A(n4904), .Z(n6045) );
  NAND U5694 ( .A(n6449), .B(n6450), .Z(n4904) );
  AND U5695 ( .A(n4926), .B(n4922), .Z(n6450) );
  OR U5696 ( .A(B[176]), .B(A[176]), .Z(n4926) );
  ANDN U5697 ( .B(n4913), .A(n4916), .Z(n6449) );
  ANDN U5698 ( .B(n4883), .A(n4860), .Z(n6448) );
  ANDN U5699 ( .B(n6451), .A(n4839), .Z(n6043) );
  AND U5700 ( .A(B[190]), .B(A[190]), .Z(n4839) );
  NAND U5701 ( .A(n6452), .B(n4841), .Z(n6451) );
  OR U5702 ( .A(A[190]), .B(B[190]), .Z(n4841) );
  NANDN U5703 ( .A(n4843), .B(n6453), .Z(n6452) );
  NAND U5704 ( .A(n6454), .B(n4846), .Z(n6453) );
  OR U5705 ( .A(B[189]), .B(A[189]), .Z(n4846) );
  NANDN U5706 ( .A(n4853), .B(n6455), .Z(n6454) );
  NANDN U5707 ( .A(n4855), .B(n6456), .Z(n6455) );
  NANDN U5708 ( .A(n4858), .B(n6457), .Z(n6456) );
  NANDN U5709 ( .A(n4860), .B(n6458), .Z(n6457) );
  NANDN U5710 ( .A(n4880), .B(n6459), .Z(n6458) );
  NAND U5711 ( .A(n4903), .B(n4883), .Z(n6459) );
  AND U5712 ( .A(n6460), .B(n6461), .Z(n4883) );
  AND U5713 ( .A(n4900), .B(n4896), .Z(n6461) );
  OR U5714 ( .A(B[180]), .B(A[180]), .Z(n4900) );
  AND U5715 ( .A(n4891), .B(n4887), .Z(n6460) );
  NANDN U5716 ( .A(n4912), .B(n6462), .Z(n4903) );
  NAND U5717 ( .A(n6463), .B(n4913), .Z(n6462) );
  OR U5718 ( .A(B[179]), .B(A[179]), .Z(n4913) );
  NANDN U5719 ( .A(n4915), .B(n6464), .Z(n6463) );
  NANDN U5720 ( .A(n4916), .B(n6465), .Z(n6464) );
  NANDN U5721 ( .A(n4919), .B(n6466), .Z(n6465) );
  NAND U5722 ( .A(n4922), .B(n4924), .Z(n6466) );
  AND U5723 ( .A(A[176]), .B(B[176]), .Z(n4924) );
  OR U5724 ( .A(B[177]), .B(A[177]), .Z(n4922) );
  AND U5725 ( .A(B[177]), .B(A[177]), .Z(n4919) );
  NOR U5726 ( .A(B[178]), .B(A[178]), .Z(n4916) );
  AND U5727 ( .A(B[178]), .B(A[178]), .Z(n4915) );
  AND U5728 ( .A(B[179]), .B(A[179]), .Z(n4912) );
  NANDN U5729 ( .A(n4886), .B(n6467), .Z(n4880) );
  NAND U5730 ( .A(n6468), .B(n4887), .Z(n6467) );
  OR U5731 ( .A(B[183]), .B(A[183]), .Z(n4887) );
  NANDN U5732 ( .A(n4889), .B(n6469), .Z(n6468) );
  NAND U5733 ( .A(n6470), .B(n4891), .Z(n6469) );
  OR U5734 ( .A(B[182]), .B(A[182]), .Z(n4891) );
  NANDN U5735 ( .A(n4893), .B(n6471), .Z(n6470) );
  NAND U5736 ( .A(n4896), .B(n4898), .Z(n6471) );
  AND U5737 ( .A(B[180]), .B(A[180]), .Z(n4898) );
  OR U5738 ( .A(B[181]), .B(A[181]), .Z(n4896) );
  AND U5739 ( .A(B[181]), .B(A[181]), .Z(n4893) );
  AND U5740 ( .A(B[182]), .B(A[182]), .Z(n4889) );
  AND U5741 ( .A(B[183]), .B(A[183]), .Z(n4886) );
  NAND U5742 ( .A(n6472), .B(n6473), .Z(n4860) );
  AND U5743 ( .A(n4878), .B(n4874), .Z(n6473) );
  OR U5744 ( .A(B[184]), .B(A[184]), .Z(n4878) );
  AND U5745 ( .A(n4869), .B(n4865), .Z(n6472) );
  NANDN U5746 ( .A(n4864), .B(n6474), .Z(n4858) );
  NAND U5747 ( .A(n6475), .B(n4865), .Z(n6474) );
  OR U5748 ( .A(B[187]), .B(A[187]), .Z(n4865) );
  NANDN U5749 ( .A(n4867), .B(n6476), .Z(n6475) );
  NAND U5750 ( .A(n6477), .B(n4869), .Z(n6476) );
  OR U5751 ( .A(B[186]), .B(A[186]), .Z(n4869) );
  NANDN U5752 ( .A(n4871), .B(n6478), .Z(n6477) );
  NAND U5753 ( .A(n4874), .B(n4876), .Z(n6478) );
  AND U5754 ( .A(B[184]), .B(A[184]), .Z(n4876) );
  OR U5755 ( .A(B[185]), .B(A[185]), .Z(n4874) );
  AND U5756 ( .A(B[185]), .B(A[185]), .Z(n4871) );
  AND U5757 ( .A(B[186]), .B(A[186]), .Z(n4867) );
  AND U5758 ( .A(B[187]), .B(A[187]), .Z(n4864) );
  NOR U5759 ( .A(B[188]), .B(A[188]), .Z(n4855) );
  AND U5760 ( .A(B[188]), .B(A[188]), .Z(n4853) );
  AND U5761 ( .A(B[189]), .B(A[189]), .Z(n4843) );
  NOR U5762 ( .A(B[191]), .B(A[191]), .Z(n4836) );
  NOR U5763 ( .A(n4814), .B(n4762), .Z(n6038) );
  NAND U5764 ( .A(n6479), .B(n6480), .Z(n4814) );
  AND U5765 ( .A(n4832), .B(n4828), .Z(n6480) );
  OR U5766 ( .A(B[192]), .B(A[192]), .Z(n4832) );
  ANDN U5767 ( .B(n4819), .A(n4822), .Z(n6479) );
  ANDN U5768 ( .B(n6481), .A(n4755), .Z(n6036) );
  AND U5769 ( .A(B[204]), .B(A[204]), .Z(n4755) );
  NAND U5770 ( .A(n6482), .B(n4758), .Z(n6481) );
  OR U5771 ( .A(A[204]), .B(B[204]), .Z(n4758) );
  NANDN U5772 ( .A(n4760), .B(n6483), .Z(n6482) );
  NANDN U5773 ( .A(n4762), .B(n6484), .Z(n6483) );
  NANDN U5774 ( .A(n4782), .B(n6485), .Z(n6484) );
  NAND U5775 ( .A(n4813), .B(n4785), .Z(n6485) );
  AND U5776 ( .A(n6486), .B(n6487), .Z(n4785) );
  AND U5777 ( .A(n4810), .B(n4806), .Z(n6487) );
  OR U5778 ( .A(B[196]), .B(A[196]), .Z(n4810) );
  AND U5779 ( .A(n4801), .B(n4797), .Z(n6486) );
  NANDN U5780 ( .A(n4818), .B(n6488), .Z(n4813) );
  NAND U5781 ( .A(n6489), .B(n4819), .Z(n6488) );
  OR U5782 ( .A(B[195]), .B(A[195]), .Z(n4819) );
  NANDN U5783 ( .A(n4821), .B(n6490), .Z(n6489) );
  NANDN U5784 ( .A(n4822), .B(n6491), .Z(n6490) );
  NANDN U5785 ( .A(n4825), .B(n6492), .Z(n6491) );
  NAND U5786 ( .A(n4828), .B(n4830), .Z(n6492) );
  AND U5787 ( .A(A[192]), .B(B[192]), .Z(n4830) );
  OR U5788 ( .A(B[193]), .B(A[193]), .Z(n4828) );
  AND U5789 ( .A(B[193]), .B(A[193]), .Z(n4825) );
  NOR U5790 ( .A(B[194]), .B(A[194]), .Z(n4822) );
  AND U5791 ( .A(B[194]), .B(A[194]), .Z(n4821) );
  AND U5792 ( .A(B[195]), .B(A[195]), .Z(n4818) );
  NANDN U5793 ( .A(n4796), .B(n6493), .Z(n4782) );
  NAND U5794 ( .A(n6494), .B(n4797), .Z(n6493) );
  OR U5795 ( .A(B[199]), .B(A[199]), .Z(n4797) );
  NANDN U5796 ( .A(n4799), .B(n6495), .Z(n6494) );
  NAND U5797 ( .A(n6496), .B(n4801), .Z(n6495) );
  OR U5798 ( .A(B[198]), .B(A[198]), .Z(n4801) );
  NANDN U5799 ( .A(n4803), .B(n6497), .Z(n6496) );
  NAND U5800 ( .A(n4806), .B(n4808), .Z(n6497) );
  AND U5801 ( .A(B[196]), .B(A[196]), .Z(n4808) );
  OR U5802 ( .A(B[197]), .B(A[197]), .Z(n4806) );
  AND U5803 ( .A(B[197]), .B(A[197]), .Z(n4803) );
  AND U5804 ( .A(B[198]), .B(A[198]), .Z(n4799) );
  AND U5805 ( .A(B[199]), .B(A[199]), .Z(n4796) );
  NAND U5806 ( .A(n6498), .B(n6499), .Z(n4762) );
  AND U5807 ( .A(n4780), .B(n4776), .Z(n6499) );
  OR U5808 ( .A(B[200]), .B(A[200]), .Z(n4780) );
  AND U5809 ( .A(n4771), .B(n4767), .Z(n6498) );
  NANDN U5810 ( .A(n4766), .B(n6500), .Z(n4760) );
  NAND U5811 ( .A(n6501), .B(n4767), .Z(n6500) );
  OR U5812 ( .A(B[203]), .B(A[203]), .Z(n4767) );
  NANDN U5813 ( .A(n4769), .B(n6502), .Z(n6501) );
  NAND U5814 ( .A(n6503), .B(n4771), .Z(n6502) );
  OR U5815 ( .A(B[202]), .B(A[202]), .Z(n4771) );
  NANDN U5816 ( .A(n4773), .B(n6504), .Z(n6503) );
  NAND U5817 ( .A(n4776), .B(n4778), .Z(n6504) );
  AND U5818 ( .A(B[200]), .B(A[200]), .Z(n4778) );
  OR U5819 ( .A(B[201]), .B(A[201]), .Z(n4776) );
  AND U5820 ( .A(B[201]), .B(A[201]), .Z(n4773) );
  AND U5821 ( .A(B[202]), .B(A[202]), .Z(n4769) );
  AND U5822 ( .A(B[203]), .B(A[203]), .Z(n4766) );
  NOR U5823 ( .A(B[205]), .B(A[205]), .Z(n4752) );
  AND U5824 ( .A(B[205]), .B(A[205]), .Z(n4750) );
  NOR U5825 ( .A(B[206]), .B(A[206]), .Z(n4747) );
  AND U5826 ( .A(B[206]), .B(A[206]), .Z(n4746) );
  NOR U5827 ( .A(B[207]), .B(A[207]), .Z(n4743) );
  NOR U5828 ( .A(n4716), .B(n4668), .Z(n6027) );
  NAND U5829 ( .A(n6505), .B(n6506), .Z(n4716) );
  AND U5830 ( .A(n4739), .B(n4730), .Z(n6506) );
  OR U5831 ( .A(B[208]), .B(A[208]), .Z(n4739) );
  ANDN U5832 ( .B(n4721), .A(n4724), .Z(n6505) );
  ANDN U5833 ( .B(n6507), .A(n4661), .Z(n6025) );
  AND U5834 ( .A(B[220]), .B(A[220]), .Z(n4661) );
  NAND U5835 ( .A(n6508), .B(n4664), .Z(n6507) );
  OR U5836 ( .A(A[220]), .B(B[220]), .Z(n4664) );
  NANDN U5837 ( .A(n4666), .B(n6509), .Z(n6508) );
  NANDN U5838 ( .A(n4668), .B(n6510), .Z(n6509) );
  NANDN U5839 ( .A(n4692), .B(n6511), .Z(n6510) );
  NAND U5840 ( .A(n4715), .B(n4695), .Z(n6511) );
  AND U5841 ( .A(n6512), .B(n6513), .Z(n4695) );
  AND U5842 ( .A(n4712), .B(n4708), .Z(n6513) );
  OR U5843 ( .A(B[212]), .B(A[212]), .Z(n4712) );
  AND U5844 ( .A(n4703), .B(n4699), .Z(n6512) );
  NANDN U5845 ( .A(n4720), .B(n6514), .Z(n4715) );
  NAND U5846 ( .A(n6515), .B(n4721), .Z(n6514) );
  OR U5847 ( .A(B[211]), .B(A[211]), .Z(n4721) );
  NANDN U5848 ( .A(n4723), .B(n6516), .Z(n6515) );
  NANDN U5849 ( .A(n4724), .B(n6517), .Z(n6516) );
  NANDN U5850 ( .A(n4727), .B(n6518), .Z(n6517) );
  NAND U5851 ( .A(n4730), .B(n4737), .Z(n6518) );
  AND U5852 ( .A(A[208]), .B(B[208]), .Z(n4737) );
  OR U5853 ( .A(B[209]), .B(A[209]), .Z(n4730) );
  AND U5854 ( .A(B[209]), .B(A[209]), .Z(n4727) );
  NOR U5855 ( .A(B[210]), .B(A[210]), .Z(n4724) );
  AND U5856 ( .A(B[210]), .B(A[210]), .Z(n4723) );
  AND U5857 ( .A(B[211]), .B(A[211]), .Z(n4720) );
  NANDN U5858 ( .A(n4698), .B(n6519), .Z(n4692) );
  NAND U5859 ( .A(n6520), .B(n4699), .Z(n6519) );
  OR U5860 ( .A(B[215]), .B(A[215]), .Z(n4699) );
  NANDN U5861 ( .A(n4701), .B(n6521), .Z(n6520) );
  NAND U5862 ( .A(n6522), .B(n4703), .Z(n6521) );
  OR U5863 ( .A(B[214]), .B(A[214]), .Z(n4703) );
  NANDN U5864 ( .A(n4705), .B(n6523), .Z(n6522) );
  NAND U5865 ( .A(n4708), .B(n4710), .Z(n6523) );
  AND U5866 ( .A(B[212]), .B(A[212]), .Z(n4710) );
  OR U5867 ( .A(B[213]), .B(A[213]), .Z(n4708) );
  AND U5868 ( .A(B[213]), .B(A[213]), .Z(n4705) );
  AND U5869 ( .A(B[214]), .B(A[214]), .Z(n4701) );
  AND U5870 ( .A(B[215]), .B(A[215]), .Z(n4698) );
  NAND U5871 ( .A(n6524), .B(n6525), .Z(n4668) );
  AND U5872 ( .A(n4690), .B(n4686), .Z(n6525) );
  OR U5873 ( .A(B[216]), .B(A[216]), .Z(n4690) );
  AND U5874 ( .A(n4681), .B(n4677), .Z(n6524) );
  NANDN U5875 ( .A(n4676), .B(n6526), .Z(n4666) );
  NAND U5876 ( .A(n6527), .B(n4677), .Z(n6526) );
  OR U5877 ( .A(B[219]), .B(A[219]), .Z(n4677) );
  NANDN U5878 ( .A(n4679), .B(n6528), .Z(n6527) );
  NAND U5879 ( .A(n6529), .B(n4681), .Z(n6528) );
  OR U5880 ( .A(B[218]), .B(A[218]), .Z(n4681) );
  NANDN U5881 ( .A(n4683), .B(n6530), .Z(n6529) );
  NAND U5882 ( .A(n4686), .B(n4688), .Z(n6530) );
  AND U5883 ( .A(B[216]), .B(A[216]), .Z(n4688) );
  OR U5884 ( .A(B[217]), .B(A[217]), .Z(n4686) );
  AND U5885 ( .A(B[217]), .B(A[217]), .Z(n4683) );
  AND U5886 ( .A(B[218]), .B(A[218]), .Z(n4679) );
  AND U5887 ( .A(B[219]), .B(A[219]), .Z(n4676) );
  NOR U5888 ( .A(B[221]), .B(A[221]), .Z(n4658) );
  AND U5889 ( .A(B[221]), .B(A[221]), .Z(n4656) );
  NOR U5890 ( .A(B[222]), .B(A[222]), .Z(n4653) );
  AND U5891 ( .A(B[222]), .B(A[222]), .Z(n4652) );
  NOR U5892 ( .A(B[223]), .B(A[223]), .Z(n4649) );
  NOR U5893 ( .A(n4627), .B(n4578), .Z(n6016) );
  NAND U5894 ( .A(n6531), .B(n6532), .Z(n4627) );
  AND U5895 ( .A(n4645), .B(n4641), .Z(n6532) );
  OR U5896 ( .A(B[224]), .B(A[224]), .Z(n4645) );
  ANDN U5897 ( .B(n4632), .A(n4635), .Z(n6531) );
  ANDN U5898 ( .B(n6533), .A(n4571), .Z(n6014) );
  AND U5899 ( .A(B[236]), .B(A[236]), .Z(n4571) );
  NAND U5900 ( .A(n6534), .B(n4574), .Z(n6533) );
  OR U5901 ( .A(A[236]), .B(B[236]), .Z(n4574) );
  NANDN U5902 ( .A(n4576), .B(n6535), .Z(n6534) );
  NANDN U5903 ( .A(n4578), .B(n6536), .Z(n6535) );
  NANDN U5904 ( .A(n4598), .B(n6537), .Z(n6536) );
  NAND U5905 ( .A(n4626), .B(n4601), .Z(n6537) );
  AND U5906 ( .A(n6538), .B(n6539), .Z(n4601) );
  AND U5907 ( .A(n4623), .B(n4614), .Z(n6539) );
  OR U5908 ( .A(B[228]), .B(A[228]), .Z(n4623) );
  AND U5909 ( .A(n4609), .B(n4605), .Z(n6538) );
  NANDN U5910 ( .A(n4631), .B(n6540), .Z(n4626) );
  NAND U5911 ( .A(n6541), .B(n4632), .Z(n6540) );
  OR U5912 ( .A(B[227]), .B(A[227]), .Z(n4632) );
  NANDN U5913 ( .A(n4634), .B(n6542), .Z(n6541) );
  NANDN U5914 ( .A(n4635), .B(n6543), .Z(n6542) );
  NANDN U5915 ( .A(n4638), .B(n6544), .Z(n6543) );
  NAND U5916 ( .A(n4641), .B(n4643), .Z(n6544) );
  AND U5917 ( .A(A[224]), .B(B[224]), .Z(n4643) );
  OR U5918 ( .A(B[225]), .B(A[225]), .Z(n4641) );
  AND U5919 ( .A(B[225]), .B(A[225]), .Z(n4638) );
  NOR U5920 ( .A(B[226]), .B(A[226]), .Z(n4635) );
  AND U5921 ( .A(B[226]), .B(A[226]), .Z(n4634) );
  AND U5922 ( .A(B[227]), .B(A[227]), .Z(n4631) );
  NANDN U5923 ( .A(n4604), .B(n6545), .Z(n4598) );
  NAND U5924 ( .A(n6546), .B(n4605), .Z(n6545) );
  OR U5925 ( .A(B[231]), .B(A[231]), .Z(n4605) );
  NANDN U5926 ( .A(n4607), .B(n6547), .Z(n6546) );
  NAND U5927 ( .A(n6548), .B(n4609), .Z(n6547) );
  OR U5928 ( .A(B[230]), .B(A[230]), .Z(n4609) );
  NANDN U5929 ( .A(n4611), .B(n6549), .Z(n6548) );
  NAND U5930 ( .A(n4614), .B(n4621), .Z(n6549) );
  AND U5931 ( .A(B[228]), .B(A[228]), .Z(n4621) );
  OR U5932 ( .A(B[229]), .B(A[229]), .Z(n4614) );
  AND U5933 ( .A(B[229]), .B(A[229]), .Z(n4611) );
  AND U5934 ( .A(B[230]), .B(A[230]), .Z(n4607) );
  AND U5935 ( .A(B[231]), .B(A[231]), .Z(n4604) );
  NAND U5936 ( .A(n6550), .B(n6551), .Z(n4578) );
  AND U5937 ( .A(n4596), .B(n4592), .Z(n6551) );
  OR U5938 ( .A(B[232]), .B(A[232]), .Z(n4596) );
  AND U5939 ( .A(n4587), .B(n4583), .Z(n6550) );
  NANDN U5940 ( .A(n4582), .B(n6552), .Z(n4576) );
  NAND U5941 ( .A(n6553), .B(n4583), .Z(n6552) );
  OR U5942 ( .A(B[235]), .B(A[235]), .Z(n4583) );
  NANDN U5943 ( .A(n4585), .B(n6554), .Z(n6553) );
  NAND U5944 ( .A(n6555), .B(n4587), .Z(n6554) );
  OR U5945 ( .A(B[234]), .B(A[234]), .Z(n4587) );
  NANDN U5946 ( .A(n4589), .B(n6556), .Z(n6555) );
  NAND U5947 ( .A(n4592), .B(n4594), .Z(n6556) );
  AND U5948 ( .A(B[232]), .B(A[232]), .Z(n4594) );
  OR U5949 ( .A(B[233]), .B(A[233]), .Z(n4592) );
  AND U5950 ( .A(B[233]), .B(A[233]), .Z(n4589) );
  AND U5951 ( .A(B[234]), .B(A[234]), .Z(n4585) );
  AND U5952 ( .A(B[235]), .B(A[235]), .Z(n4582) );
  NOR U5953 ( .A(B[237]), .B(A[237]), .Z(n4568) );
  AND U5954 ( .A(B[237]), .B(A[237]), .Z(n4566) );
  NOR U5955 ( .A(B[238]), .B(A[238]), .Z(n4563) );
  AND U5956 ( .A(B[238]), .B(A[238]), .Z(n4562) );
  NOR U5957 ( .A(B[239]), .B(A[239]), .Z(n4559) );
  NOR U5958 ( .A(n4529), .B(n4480), .Z(n6005) );
  NAND U5959 ( .A(n6557), .B(n6558), .Z(n4529) );
  AND U5960 ( .A(n4547), .B(n4543), .Z(n6558) );
  OR U5961 ( .A(B[240]), .B(A[240]), .Z(n4547) );
  ANDN U5962 ( .B(n4534), .A(n4537), .Z(n6557) );
  ANDN U5963 ( .B(n6559), .A(n4473), .Z(n6003) );
  AND U5964 ( .A(B[252]), .B(A[252]), .Z(n4473) );
  NAND U5965 ( .A(n6560), .B(n4476), .Z(n6559) );
  OR U5966 ( .A(A[252]), .B(B[252]), .Z(n4476) );
  NANDN U5967 ( .A(n4478), .B(n6561), .Z(n6560) );
  NANDN U5968 ( .A(n4480), .B(n6562), .Z(n6561) );
  NANDN U5969 ( .A(n4505), .B(n6563), .Z(n6562) );
  NAND U5970 ( .A(n4528), .B(n4508), .Z(n6563) );
  AND U5971 ( .A(n6564), .B(n6565), .Z(n4508) );
  AND U5972 ( .A(n4525), .B(n4521), .Z(n6565) );
  OR U5973 ( .A(B[244]), .B(A[244]), .Z(n4525) );
  AND U5974 ( .A(n4516), .B(n4512), .Z(n6564) );
  NANDN U5975 ( .A(n4533), .B(n6566), .Z(n4528) );
  NAND U5976 ( .A(n6567), .B(n4534), .Z(n6566) );
  OR U5977 ( .A(B[243]), .B(A[243]), .Z(n4534) );
  NANDN U5978 ( .A(n4536), .B(n6568), .Z(n6567) );
  NANDN U5979 ( .A(n4537), .B(n6569), .Z(n6568) );
  NANDN U5980 ( .A(n4540), .B(n6570), .Z(n6569) );
  NAND U5981 ( .A(n4543), .B(n4545), .Z(n6570) );
  AND U5982 ( .A(A[240]), .B(B[240]), .Z(n4545) );
  OR U5983 ( .A(B[241]), .B(A[241]), .Z(n4543) );
  AND U5984 ( .A(B[241]), .B(A[241]), .Z(n4540) );
  NOR U5985 ( .A(B[242]), .B(A[242]), .Z(n4537) );
  AND U5986 ( .A(B[242]), .B(A[242]), .Z(n4536) );
  AND U5987 ( .A(B[243]), .B(A[243]), .Z(n4533) );
  NANDN U5988 ( .A(n4511), .B(n6571), .Z(n4505) );
  NAND U5989 ( .A(n6572), .B(n4512), .Z(n6571) );
  OR U5990 ( .A(B[247]), .B(A[247]), .Z(n4512) );
  NANDN U5991 ( .A(n4514), .B(n6573), .Z(n6572) );
  NAND U5992 ( .A(n6574), .B(n4516), .Z(n6573) );
  OR U5993 ( .A(B[246]), .B(A[246]), .Z(n4516) );
  NANDN U5994 ( .A(n4518), .B(n6575), .Z(n6574) );
  NAND U5995 ( .A(n4521), .B(n4523), .Z(n6575) );
  AND U5996 ( .A(B[244]), .B(A[244]), .Z(n4523) );
  OR U5997 ( .A(B[245]), .B(A[245]), .Z(n4521) );
  AND U5998 ( .A(B[245]), .B(A[245]), .Z(n4518) );
  AND U5999 ( .A(B[246]), .B(A[246]), .Z(n4514) );
  AND U6000 ( .A(B[247]), .B(A[247]), .Z(n4511) );
  NAND U6001 ( .A(n6576), .B(n6577), .Z(n4480) );
  AND U6002 ( .A(n4503), .B(n4494), .Z(n6577) );
  OR U6003 ( .A(B[248]), .B(A[248]), .Z(n4503) );
  AND U6004 ( .A(n4489), .B(n4485), .Z(n6576) );
  NANDN U6005 ( .A(n4484), .B(n6578), .Z(n4478) );
  NAND U6006 ( .A(n6579), .B(n4485), .Z(n6578) );
  OR U6007 ( .A(B[251]), .B(A[251]), .Z(n4485) );
  NANDN U6008 ( .A(n4487), .B(n6580), .Z(n6579) );
  NAND U6009 ( .A(n6581), .B(n4489), .Z(n6580) );
  OR U6010 ( .A(B[250]), .B(A[250]), .Z(n4489) );
  NANDN U6011 ( .A(n4491), .B(n6582), .Z(n6581) );
  NAND U6012 ( .A(n4494), .B(n4501), .Z(n6582) );
  AND U6013 ( .A(B[248]), .B(A[248]), .Z(n4501) );
  OR U6014 ( .A(B[249]), .B(A[249]), .Z(n4494) );
  AND U6015 ( .A(B[249]), .B(A[249]), .Z(n4491) );
  AND U6016 ( .A(B[250]), .B(A[250]), .Z(n4487) );
  AND U6017 ( .A(B[251]), .B(A[251]), .Z(n4484) );
  NOR U6018 ( .A(B[253]), .B(A[253]), .Z(n4470) );
  AND U6019 ( .A(B[253]), .B(A[253]), .Z(n4468) );
  NOR U6020 ( .A(B[254]), .B(A[254]), .Z(n4465) );
  AND U6021 ( .A(B[254]), .B(A[254]), .Z(n4464) );
  NOR U6022 ( .A(B[255]), .B(A[255]), .Z(n4461) );
  NOR U6023 ( .A(n4364), .B(n5889), .Z(n5972) );
  NAND U6024 ( .A(n6583), .B(n6584), .Z(n5889) );
  AND U6025 ( .A(n6585), .B(n6586), .Z(n6584) );
  AND U6026 ( .A(n4095), .B(n4090), .Z(n6586) );
  OR U6027 ( .A(A[317]), .B(B[317]), .Z(n4090) );
  OR U6028 ( .A(A[316]), .B(B[316]), .Z(n4095) );
  AND U6029 ( .A(n4085), .B(n4081), .Z(n6585) );
  OR U6030 ( .A(B[319]), .B(A[319]), .Z(n4081) );
  OR U6031 ( .A(A[318]), .B(B[318]), .Z(n4085) );
  ANDN U6032 ( .B(n6587), .A(n4121), .Z(n6583) );
  NAND U6033 ( .A(n6588), .B(n6589), .Z(n4121) );
  AND U6034 ( .A(n4144), .B(n4135), .Z(n6589) );
  OR U6035 ( .A(A[309]), .B(B[309]), .Z(n4135) );
  OR U6036 ( .A(A[308]), .B(B[308]), .Z(n4144) );
  AND U6037 ( .A(n4130), .B(n4126), .Z(n6588) );
  OR U6038 ( .A(B[311]), .B(A[311]), .Z(n4126) );
  OR U6039 ( .A(A[310]), .B(B[310]), .Z(n4130) );
  NOR U6040 ( .A(n4148), .B(n4099), .Z(n6587) );
  NAND U6041 ( .A(n6590), .B(n6591), .Z(n4099) );
  AND U6042 ( .A(n4117), .B(n4113), .Z(n6591) );
  OR U6043 ( .A(A[313]), .B(B[313]), .Z(n4113) );
  OR U6044 ( .A(A[312]), .B(B[312]), .Z(n4117) );
  AND U6045 ( .A(n4108), .B(n4104), .Z(n6590) );
  OR U6046 ( .A(B[315]), .B(A[315]), .Z(n4104) );
  OR U6047 ( .A(A[314]), .B(B[314]), .Z(n4108) );
  NAND U6048 ( .A(n6592), .B(n6593), .Z(n4148) );
  AND U6049 ( .A(n4166), .B(n4162), .Z(n6593) );
  OR U6050 ( .A(A[305]), .B(B[305]), .Z(n4162) );
  OR U6051 ( .A(A[304]), .B(B[304]), .Z(n4166) );
  AND U6052 ( .A(n4157), .B(n4153), .Z(n6592) );
  OR U6053 ( .A(B[307]), .B(A[307]), .Z(n4153) );
  OR U6054 ( .A(A[306]), .B(B[306]), .Z(n4157) );
  NAND U6055 ( .A(n6594), .B(n6595), .Z(n4364) );
  AND U6056 ( .A(n6596), .B(n6597), .Z(n6595) );
  AND U6057 ( .A(n4388), .B(n4378), .Z(n6597) );
  OR U6058 ( .A(A[269]), .B(B[269]), .Z(n4378) );
  OR U6059 ( .A(A[268]), .B(B[268]), .Z(n4388) );
  AND U6060 ( .A(n4373), .B(n4369), .Z(n6596) );
  OR U6061 ( .A(B[271]), .B(A[271]), .Z(n4369) );
  OR U6062 ( .A(A[270]), .B(B[270]), .Z(n4373) );
  ANDN U6063 ( .B(n6598), .A(n4436), .Z(n6594) );
  NAND U6064 ( .A(n6599), .B(n6600), .Z(n4436) );
  AND U6065 ( .A(n4457), .B(n4453), .Z(n6600) );
  OR U6066 ( .A(A[257]), .B(B[257]), .Z(n4453) );
  OR U6067 ( .A(A[256]), .B(B[256]), .Z(n4457) );
  AND U6068 ( .A(n4448), .B(n4444), .Z(n6599) );
  OR U6069 ( .A(B[259]), .B(A[259]), .Z(n4444) );
  OR U6070 ( .A(A[258]), .B(B[258]), .Z(n4448) );
  NOR U6071 ( .A(n4414), .B(n4392), .Z(n6598) );
  NAND U6072 ( .A(n6601), .B(n6602), .Z(n4392) );
  AND U6073 ( .A(n4410), .B(n4406), .Z(n6602) );
  OR U6074 ( .A(A[265]), .B(B[265]), .Z(n4406) );
  OR U6075 ( .A(A[264]), .B(B[264]), .Z(n4410) );
  AND U6076 ( .A(n4401), .B(n4397), .Z(n6601) );
  OR U6077 ( .A(B[267]), .B(A[267]), .Z(n4397) );
  OR U6078 ( .A(A[266]), .B(B[266]), .Z(n4401) );
  NAND U6079 ( .A(n6603), .B(n6604), .Z(n4414) );
  AND U6080 ( .A(n4432), .B(n4428), .Z(n6604) );
  OR U6081 ( .A(A[261]), .B(B[261]), .Z(n4428) );
  OR U6082 ( .A(A[260]), .B(B[260]), .Z(n4432) );
  AND U6083 ( .A(n4423), .B(n4419), .Z(n6603) );
  OR U6084 ( .A(B[263]), .B(A[263]), .Z(n4419) );
  OR U6085 ( .A(A[262]), .B(B[262]), .Z(n4423) );
  NAND U6086 ( .A(n6605), .B(n6606), .Z(n3691) );
  NOR U6087 ( .A(n3885), .B(n3789), .Z(n6606) );
  NOR U6088 ( .A(n3982), .B(n6607), .Z(n6605) );
  NAND U6089 ( .A(n6608), .B(n6609), .Z(n3982) );
  AND U6090 ( .A(n6610), .B(n6611), .Z(n6609) );
  AND U6091 ( .A(n4000), .B(n3995), .Z(n6611) );
  AND U6092 ( .A(n3990), .B(n3986), .Z(n6610) );
  ANDN U6093 ( .B(n6612), .A(n4049), .Z(n6608) );
  NAND U6094 ( .A(n6613), .B(n6614), .Z(n4049) );
  AND U6095 ( .A(n4066), .B(n4062), .Z(n6614) );
  OR U6096 ( .A(A[320]), .B(B[320]), .Z(n4066) );
  AND U6097 ( .A(n4057), .B(n4053), .Z(n6613) );
  NOR U6098 ( .A(n4027), .B(n4004), .Z(n6612) );
  NAND U6099 ( .A(n6615), .B(n6616), .Z(n3689) );
  NAND U6100 ( .A(n6617), .B(n3696), .Z(n6616) );
  NANDN U6101 ( .A(n3698), .B(n6618), .Z(n6617) );
  NAND U6102 ( .A(n6619), .B(n3700), .Z(n6618) );
  NANDN U6103 ( .A(n3702), .B(n6620), .Z(n6619) );
  NAND U6104 ( .A(n6621), .B(n3705), .Z(n6620) );
  NANDN U6105 ( .A(n3707), .B(n6622), .Z(n6621) );
  NAND U6106 ( .A(n6623), .B(n3710), .Z(n6622) );
  NANDN U6107 ( .A(n3712), .B(n6624), .Z(n6623) );
  NANDN U6108 ( .A(n3714), .B(n6625), .Z(n6624) );
  NANDN U6109 ( .A(n3738), .B(n6626), .Z(n6625) );
  NANDN U6110 ( .A(n3740), .B(n3761), .Z(n6626) );
  NANDN U6111 ( .A(n3766), .B(n6627), .Z(n3761) );
  NAND U6112 ( .A(n6628), .B(n3767), .Z(n6627) );
  NANDN U6113 ( .A(n3769), .B(n6629), .Z(n6628) );
  NAND U6114 ( .A(n6630), .B(n3771), .Z(n6629) );
  NANDN U6115 ( .A(n3773), .B(n6631), .Z(n6630) );
  NAND U6116 ( .A(n3776), .B(n3783), .Z(n6631) );
  AND U6117 ( .A(A[368]), .B(B[368]), .Z(n3783) );
  AND U6118 ( .A(A[369]), .B(B[369]), .Z(n3773) );
  AND U6119 ( .A(A[370]), .B(B[370]), .Z(n3769) );
  AND U6120 ( .A(B[371]), .B(A[371]), .Z(n3766) );
  NANDN U6121 ( .A(n3744), .B(n6632), .Z(n3738) );
  NAND U6122 ( .A(n6633), .B(n3745), .Z(n6632) );
  NANDN U6123 ( .A(n3747), .B(n6634), .Z(n6633) );
  NAND U6124 ( .A(n6635), .B(n3749), .Z(n6634) );
  NANDN U6125 ( .A(n3751), .B(n6636), .Z(n6635) );
  NAND U6126 ( .A(n3754), .B(n3756), .Z(n6636) );
  AND U6127 ( .A(A[372]), .B(B[372]), .Z(n3756) );
  AND U6128 ( .A(A[373]), .B(B[373]), .Z(n3751) );
  AND U6129 ( .A(A[374]), .B(B[374]), .Z(n3747) );
  AND U6130 ( .A(B[375]), .B(A[375]), .Z(n3744) );
  NANDN U6131 ( .A(n3722), .B(n6637), .Z(n3712) );
  NAND U6132 ( .A(n6638), .B(n3723), .Z(n6637) );
  NANDN U6133 ( .A(n3725), .B(n6639), .Z(n6638) );
  NAND U6134 ( .A(n6640), .B(n3727), .Z(n6639) );
  NANDN U6135 ( .A(n3729), .B(n6641), .Z(n6640) );
  NAND U6136 ( .A(n3732), .B(n3734), .Z(n6641) );
  AND U6137 ( .A(A[376]), .B(B[376]), .Z(n3734) );
  AND U6138 ( .A(A[377]), .B(B[377]), .Z(n3729) );
  AND U6139 ( .A(A[378]), .B(B[378]), .Z(n3725) );
  AND U6140 ( .A(B[379]), .B(A[379]), .Z(n3722) );
  AND U6141 ( .A(A[380]), .B(B[380]), .Z(n3707) );
  AND U6142 ( .A(A[381]), .B(B[381]), .Z(n3702) );
  AND U6143 ( .A(A[382]), .B(B[382]), .Z(n3698) );
  ANDN U6144 ( .B(n6642), .A(n3695), .Z(n6615) );
  AND U6145 ( .A(B[383]), .B(A[383]), .Z(n3695) );
  NANDN U6146 ( .A(n6607), .B(n6643), .Z(n6642) );
  NANDN U6147 ( .A(n3787), .B(n6644), .Z(n6643) );
  NANDN U6148 ( .A(n3789), .B(n6645), .Z(n6644) );
  NANDN U6149 ( .A(n3883), .B(n6646), .Z(n6645) );
  NANDN U6150 ( .A(n3885), .B(n3981), .Z(n6646) );
  NANDN U6151 ( .A(n3985), .B(n6647), .Z(n3981) );
  NAND U6152 ( .A(n6648), .B(n3986), .Z(n6647) );
  OR U6153 ( .A(B[335]), .B(A[335]), .Z(n3986) );
  NANDN U6154 ( .A(n3988), .B(n6649), .Z(n6648) );
  NAND U6155 ( .A(n6650), .B(n3990), .Z(n6649) );
  OR U6156 ( .A(A[334]), .B(B[334]), .Z(n3990) );
  NANDN U6157 ( .A(n3992), .B(n6651), .Z(n6650) );
  NAND U6158 ( .A(n6652), .B(n3995), .Z(n6651) );
  OR U6159 ( .A(A[333]), .B(B[333]), .Z(n3995) );
  NANDN U6160 ( .A(n3997), .B(n6653), .Z(n6652) );
  NAND U6161 ( .A(n6654), .B(n4000), .Z(n6653) );
  OR U6162 ( .A(A[332]), .B(B[332]), .Z(n4000) );
  NANDN U6163 ( .A(n4002), .B(n6655), .Z(n6654) );
  NANDN U6164 ( .A(n4004), .B(n6656), .Z(n6655) );
  NANDN U6165 ( .A(n4025), .B(n6657), .Z(n6656) );
  NANDN U6166 ( .A(n4027), .B(n4048), .Z(n6657) );
  NANDN U6167 ( .A(n4052), .B(n6658), .Z(n4048) );
  NAND U6168 ( .A(n6659), .B(n4053), .Z(n6658) );
  OR U6169 ( .A(B[323]), .B(A[323]), .Z(n4053) );
  NANDN U6170 ( .A(n4055), .B(n6660), .Z(n6659) );
  NAND U6171 ( .A(n6661), .B(n4057), .Z(n6660) );
  OR U6172 ( .A(A[322]), .B(B[322]), .Z(n4057) );
  NANDN U6173 ( .A(n4059), .B(n6662), .Z(n6661) );
  NAND U6174 ( .A(n4062), .B(n4064), .Z(n6662) );
  AND U6175 ( .A(A[320]), .B(B[320]), .Z(n4064) );
  OR U6176 ( .A(A[321]), .B(B[321]), .Z(n4062) );
  AND U6177 ( .A(A[321]), .B(B[321]), .Z(n4059) );
  AND U6178 ( .A(A[322]), .B(B[322]), .Z(n4055) );
  AND U6179 ( .A(B[323]), .B(A[323]), .Z(n4052) );
  NAND U6180 ( .A(n6663), .B(n6664), .Z(n4027) );
  AND U6181 ( .A(n4045), .B(n4041), .Z(n6664) );
  OR U6182 ( .A(A[324]), .B(B[324]), .Z(n4045) );
  AND U6183 ( .A(n4036), .B(n4032), .Z(n6663) );
  NANDN U6184 ( .A(n4031), .B(n6665), .Z(n4025) );
  NAND U6185 ( .A(n6666), .B(n4032), .Z(n6665) );
  OR U6186 ( .A(B[327]), .B(A[327]), .Z(n4032) );
  NANDN U6187 ( .A(n4034), .B(n6667), .Z(n6666) );
  NAND U6188 ( .A(n6668), .B(n4036), .Z(n6667) );
  OR U6189 ( .A(A[326]), .B(B[326]), .Z(n4036) );
  NANDN U6190 ( .A(n4038), .B(n6669), .Z(n6668) );
  NAND U6191 ( .A(n4041), .B(n4043), .Z(n6669) );
  AND U6192 ( .A(A[324]), .B(B[324]), .Z(n4043) );
  OR U6193 ( .A(A[325]), .B(B[325]), .Z(n4041) );
  AND U6194 ( .A(A[325]), .B(B[325]), .Z(n4038) );
  AND U6195 ( .A(A[326]), .B(B[326]), .Z(n4034) );
  AND U6196 ( .A(B[327]), .B(A[327]), .Z(n4031) );
  NAND U6197 ( .A(n6670), .B(n6671), .Z(n4004) );
  AND U6198 ( .A(n4023), .B(n4018), .Z(n6671) );
  OR U6199 ( .A(A[328]), .B(B[328]), .Z(n4023) );
  AND U6200 ( .A(n4013), .B(n4009), .Z(n6670) );
  NANDN U6201 ( .A(n4008), .B(n6672), .Z(n4002) );
  NAND U6202 ( .A(n6673), .B(n4009), .Z(n6672) );
  OR U6203 ( .A(B[331]), .B(A[331]), .Z(n4009) );
  NANDN U6204 ( .A(n4011), .B(n6674), .Z(n6673) );
  NAND U6205 ( .A(n6675), .B(n4013), .Z(n6674) );
  OR U6206 ( .A(A[330]), .B(B[330]), .Z(n4013) );
  NANDN U6207 ( .A(n4015), .B(n6676), .Z(n6675) );
  NAND U6208 ( .A(n4018), .B(n4021), .Z(n6676) );
  AND U6209 ( .A(A[328]), .B(B[328]), .Z(n4021) );
  OR U6210 ( .A(A[329]), .B(B[329]), .Z(n4018) );
  AND U6211 ( .A(A[329]), .B(B[329]), .Z(n4015) );
  AND U6212 ( .A(A[330]), .B(B[330]), .Z(n4011) );
  AND U6213 ( .A(B[331]), .B(A[331]), .Z(n4008) );
  AND U6214 ( .A(A[332]), .B(B[332]), .Z(n3997) );
  AND U6215 ( .A(A[333]), .B(B[333]), .Z(n3992) );
  AND U6216 ( .A(A[334]), .B(B[334]), .Z(n3988) );
  AND U6217 ( .A(B[335]), .B(A[335]), .Z(n3985) );
  NAND U6218 ( .A(n6677), .B(n6678), .Z(n3885) );
  AND U6219 ( .A(n6679), .B(n6680), .Z(n6678) );
  AND U6220 ( .A(n3909), .B(n3899), .Z(n6680) );
  AND U6221 ( .A(n3894), .B(n3890), .Z(n6679) );
  ANDN U6222 ( .B(n6681), .A(n3957), .Z(n6677) );
  NAND U6223 ( .A(n6682), .B(n6683), .Z(n3957) );
  AND U6224 ( .A(n3978), .B(n3974), .Z(n6683) );
  OR U6225 ( .A(A[336]), .B(B[336]), .Z(n3978) );
  AND U6226 ( .A(n3969), .B(n3965), .Z(n6682) );
  NOR U6227 ( .A(n3935), .B(n3913), .Z(n6681) );
  NANDN U6228 ( .A(n3889), .B(n6684), .Z(n3883) );
  NAND U6229 ( .A(n6685), .B(n3890), .Z(n6684) );
  OR U6230 ( .A(B[351]), .B(A[351]), .Z(n3890) );
  NANDN U6231 ( .A(n3892), .B(n6686), .Z(n6685) );
  NAND U6232 ( .A(n6687), .B(n3894), .Z(n6686) );
  OR U6233 ( .A(A[350]), .B(B[350]), .Z(n3894) );
  NANDN U6234 ( .A(n3896), .B(n6688), .Z(n6687) );
  NAND U6235 ( .A(n6689), .B(n3899), .Z(n6688) );
  OR U6236 ( .A(A[349]), .B(B[349]), .Z(n3899) );
  NANDN U6237 ( .A(n3906), .B(n6690), .Z(n6689) );
  NAND U6238 ( .A(n6691), .B(n3909), .Z(n6690) );
  OR U6239 ( .A(A[348]), .B(B[348]), .Z(n3909) );
  NANDN U6240 ( .A(n3911), .B(n6692), .Z(n6691) );
  NANDN U6241 ( .A(n3913), .B(n6693), .Z(n6692) );
  NANDN U6242 ( .A(n3933), .B(n6694), .Z(n6693) );
  NANDN U6243 ( .A(n3935), .B(n3956), .Z(n6694) );
  NANDN U6244 ( .A(n3964), .B(n6695), .Z(n3956) );
  NAND U6245 ( .A(n6696), .B(n3965), .Z(n6695) );
  OR U6246 ( .A(B[339]), .B(A[339]), .Z(n3965) );
  NANDN U6247 ( .A(n3967), .B(n6697), .Z(n6696) );
  NAND U6248 ( .A(n6698), .B(n3969), .Z(n6697) );
  OR U6249 ( .A(A[338]), .B(B[338]), .Z(n3969) );
  NANDN U6250 ( .A(n3971), .B(n6699), .Z(n6698) );
  NAND U6251 ( .A(n3974), .B(n3976), .Z(n6699) );
  AND U6252 ( .A(A[336]), .B(B[336]), .Z(n3976) );
  OR U6253 ( .A(A[337]), .B(B[337]), .Z(n3974) );
  AND U6254 ( .A(A[337]), .B(B[337]), .Z(n3971) );
  AND U6255 ( .A(A[338]), .B(B[338]), .Z(n3967) );
  AND U6256 ( .A(B[339]), .B(A[339]), .Z(n3964) );
  NAND U6257 ( .A(n6700), .B(n6701), .Z(n3935) );
  AND U6258 ( .A(n3953), .B(n3949), .Z(n6701) );
  OR U6259 ( .A(A[340]), .B(B[340]), .Z(n3953) );
  AND U6260 ( .A(n3944), .B(n3940), .Z(n6700) );
  NANDN U6261 ( .A(n3939), .B(n6702), .Z(n3933) );
  NAND U6262 ( .A(n6703), .B(n3940), .Z(n6702) );
  OR U6263 ( .A(B[343]), .B(A[343]), .Z(n3940) );
  NANDN U6264 ( .A(n3942), .B(n6704), .Z(n6703) );
  NAND U6265 ( .A(n6705), .B(n3944), .Z(n6704) );
  OR U6266 ( .A(A[342]), .B(B[342]), .Z(n3944) );
  NANDN U6267 ( .A(n3946), .B(n6706), .Z(n6705) );
  NAND U6268 ( .A(n3949), .B(n3951), .Z(n6706) );
  AND U6269 ( .A(A[340]), .B(B[340]), .Z(n3951) );
  OR U6270 ( .A(A[341]), .B(B[341]), .Z(n3949) );
  AND U6271 ( .A(A[341]), .B(B[341]), .Z(n3946) );
  AND U6272 ( .A(A[342]), .B(B[342]), .Z(n3942) );
  AND U6273 ( .A(B[343]), .B(A[343]), .Z(n3939) );
  NAND U6274 ( .A(n6707), .B(n6708), .Z(n3913) );
  AND U6275 ( .A(n3931), .B(n3927), .Z(n6708) );
  OR U6276 ( .A(A[344]), .B(B[344]), .Z(n3931) );
  AND U6277 ( .A(n3922), .B(n3918), .Z(n6707) );
  NANDN U6278 ( .A(n3917), .B(n6709), .Z(n3911) );
  NAND U6279 ( .A(n6710), .B(n3918), .Z(n6709) );
  OR U6280 ( .A(B[347]), .B(A[347]), .Z(n3918) );
  NANDN U6281 ( .A(n3920), .B(n6711), .Z(n6710) );
  NAND U6282 ( .A(n6712), .B(n3922), .Z(n6711) );
  OR U6283 ( .A(A[346]), .B(B[346]), .Z(n3922) );
  NANDN U6284 ( .A(n3924), .B(n6713), .Z(n6712) );
  NAND U6285 ( .A(n3927), .B(n3929), .Z(n6713) );
  AND U6286 ( .A(A[344]), .B(B[344]), .Z(n3929) );
  OR U6287 ( .A(A[345]), .B(B[345]), .Z(n3927) );
  AND U6288 ( .A(A[345]), .B(B[345]), .Z(n3924) );
  AND U6289 ( .A(A[346]), .B(B[346]), .Z(n3920) );
  AND U6290 ( .A(B[347]), .B(A[347]), .Z(n3917) );
  AND U6291 ( .A(A[348]), .B(B[348]), .Z(n3906) );
  AND U6292 ( .A(A[349]), .B(B[349]), .Z(n3896) );
  AND U6293 ( .A(A[350]), .B(B[350]), .Z(n3892) );
  AND U6294 ( .A(B[351]), .B(A[351]), .Z(n3889) );
  NAND U6295 ( .A(n6714), .B(n6715), .Z(n3789) );
  AND U6296 ( .A(n6716), .B(n6717), .Z(n6715) );
  AND U6297 ( .A(n3808), .B(n3803), .Z(n6717) );
  AND U6298 ( .A(n3798), .B(n3794), .Z(n6716) );
  ANDN U6299 ( .B(n6718), .A(n3864), .Z(n6714) );
  NAND U6300 ( .A(n6719), .B(n6720), .Z(n3864) );
  AND U6301 ( .A(n3881), .B(n3877), .Z(n6720) );
  OR U6302 ( .A(A[352]), .B(B[352]), .Z(n3881) );
  AND U6303 ( .A(n3872), .B(n3868), .Z(n6719) );
  NOR U6304 ( .A(n3834), .B(n3812), .Z(n6718) );
  NANDN U6305 ( .A(n3793), .B(n6721), .Z(n3787) );
  NAND U6306 ( .A(n6722), .B(n3794), .Z(n6721) );
  OR U6307 ( .A(B[367]), .B(A[367]), .Z(n3794) );
  NANDN U6308 ( .A(n3796), .B(n6723), .Z(n6722) );
  NAND U6309 ( .A(n6724), .B(n3798), .Z(n6723) );
  OR U6310 ( .A(A[366]), .B(B[366]), .Z(n3798) );
  NANDN U6311 ( .A(n3800), .B(n6725), .Z(n6724) );
  NAND U6312 ( .A(n6726), .B(n3803), .Z(n6725) );
  OR U6313 ( .A(A[365]), .B(B[365]), .Z(n3803) );
  NANDN U6314 ( .A(n3805), .B(n6727), .Z(n6726) );
  NAND U6315 ( .A(n6728), .B(n3808), .Z(n6727) );
  OR U6316 ( .A(A[364]), .B(B[364]), .Z(n3808) );
  NANDN U6317 ( .A(n3810), .B(n6729), .Z(n6728) );
  NANDN U6318 ( .A(n3812), .B(n6730), .Z(n6729) );
  NANDN U6319 ( .A(n3832), .B(n6731), .Z(n6730) );
  NANDN U6320 ( .A(n3834), .B(n3863), .Z(n6731) );
  NANDN U6321 ( .A(n3867), .B(n6732), .Z(n3863) );
  NAND U6322 ( .A(n6733), .B(n3868), .Z(n6732) );
  OR U6323 ( .A(B[355]), .B(A[355]), .Z(n3868) );
  NANDN U6324 ( .A(n3870), .B(n6734), .Z(n6733) );
  NAND U6325 ( .A(n6735), .B(n3872), .Z(n6734) );
  OR U6326 ( .A(A[354]), .B(B[354]), .Z(n3872) );
  NANDN U6327 ( .A(n3874), .B(n6736), .Z(n6735) );
  NAND U6328 ( .A(n3877), .B(n3879), .Z(n6736) );
  AND U6329 ( .A(A[352]), .B(B[352]), .Z(n3879) );
  OR U6330 ( .A(A[353]), .B(B[353]), .Z(n3877) );
  AND U6331 ( .A(A[353]), .B(B[353]), .Z(n3874) );
  AND U6332 ( .A(A[354]), .B(B[354]), .Z(n3870) );
  AND U6333 ( .A(B[355]), .B(A[355]), .Z(n3867) );
  NAND U6334 ( .A(n6737), .B(n6738), .Z(n3834) );
  AND U6335 ( .A(n3860), .B(n3856), .Z(n6738) );
  OR U6336 ( .A(A[356]), .B(B[356]), .Z(n3860) );
  AND U6337 ( .A(n3851), .B(n3847), .Z(n6737) );
  NANDN U6338 ( .A(n3846), .B(n6739), .Z(n3832) );
  NAND U6339 ( .A(n6740), .B(n3847), .Z(n6739) );
  OR U6340 ( .A(B[359]), .B(A[359]), .Z(n3847) );
  NANDN U6341 ( .A(n3849), .B(n6741), .Z(n6740) );
  NAND U6342 ( .A(n6742), .B(n3851), .Z(n6741) );
  OR U6343 ( .A(A[358]), .B(B[358]), .Z(n3851) );
  NANDN U6344 ( .A(n3853), .B(n6743), .Z(n6742) );
  NAND U6345 ( .A(n3856), .B(n3858), .Z(n6743) );
  AND U6346 ( .A(A[356]), .B(B[356]), .Z(n3858) );
  OR U6347 ( .A(A[357]), .B(B[357]), .Z(n3856) );
  AND U6348 ( .A(A[357]), .B(B[357]), .Z(n3853) );
  AND U6349 ( .A(A[358]), .B(B[358]), .Z(n3849) );
  AND U6350 ( .A(B[359]), .B(A[359]), .Z(n3846) );
  NAND U6351 ( .A(n6744), .B(n6745), .Z(n3812) );
  AND U6352 ( .A(n3830), .B(n3826), .Z(n6745) );
  OR U6353 ( .A(A[360]), .B(B[360]), .Z(n3830) );
  AND U6354 ( .A(n3821), .B(n3817), .Z(n6744) );
  NANDN U6355 ( .A(n3816), .B(n6746), .Z(n3810) );
  NAND U6356 ( .A(n6747), .B(n3817), .Z(n6746) );
  OR U6357 ( .A(B[363]), .B(A[363]), .Z(n3817) );
  NANDN U6358 ( .A(n3819), .B(n6748), .Z(n6747) );
  NAND U6359 ( .A(n6749), .B(n3821), .Z(n6748) );
  OR U6360 ( .A(A[362]), .B(B[362]), .Z(n3821) );
  NANDN U6361 ( .A(n3823), .B(n6750), .Z(n6749) );
  NAND U6362 ( .A(n3826), .B(n3828), .Z(n6750) );
  AND U6363 ( .A(A[360]), .B(B[360]), .Z(n3828) );
  OR U6364 ( .A(A[361]), .B(B[361]), .Z(n3826) );
  AND U6365 ( .A(A[361]), .B(B[361]), .Z(n3823) );
  AND U6366 ( .A(A[362]), .B(B[362]), .Z(n3819) );
  AND U6367 ( .A(B[363]), .B(A[363]), .Z(n3816) );
  AND U6368 ( .A(A[364]), .B(B[364]), .Z(n3805) );
  AND U6369 ( .A(A[365]), .B(B[365]), .Z(n3800) );
  AND U6370 ( .A(A[366]), .B(B[366]), .Z(n3796) );
  AND U6371 ( .A(B[367]), .B(A[367]), .Z(n3793) );
  NAND U6372 ( .A(n6751), .B(n6752), .Z(n6607) );
  AND U6373 ( .A(n6753), .B(n6754), .Z(n6752) );
  AND U6374 ( .A(n3710), .B(n3705), .Z(n6754) );
  OR U6375 ( .A(A[381]), .B(B[381]), .Z(n3705) );
  OR U6376 ( .A(A[380]), .B(B[380]), .Z(n3710) );
  AND U6377 ( .A(n3700), .B(n3696), .Z(n6753) );
  OR U6378 ( .A(B[383]), .B(A[383]), .Z(n3696) );
  OR U6379 ( .A(A[382]), .B(B[382]), .Z(n3700) );
  ANDN U6380 ( .B(n6755), .A(n3740), .Z(n6751) );
  NAND U6381 ( .A(n6756), .B(n6757), .Z(n3740) );
  AND U6382 ( .A(n3758), .B(n3754), .Z(n6757) );
  OR U6383 ( .A(A[373]), .B(B[373]), .Z(n3754) );
  OR U6384 ( .A(A[372]), .B(B[372]), .Z(n3758) );
  AND U6385 ( .A(n3749), .B(n3745), .Z(n6756) );
  OR U6386 ( .A(B[375]), .B(A[375]), .Z(n3745) );
  OR U6387 ( .A(A[374]), .B(B[374]), .Z(n3749) );
  NOR U6388 ( .A(n3762), .B(n3714), .Z(n6755) );
  NAND U6389 ( .A(n6758), .B(n6759), .Z(n3714) );
  AND U6390 ( .A(n3736), .B(n3732), .Z(n6759) );
  OR U6391 ( .A(A[377]), .B(B[377]), .Z(n3732) );
  OR U6392 ( .A(A[376]), .B(B[376]), .Z(n3736) );
  AND U6393 ( .A(n3727), .B(n3723), .Z(n6758) );
  OR U6394 ( .A(B[379]), .B(A[379]), .Z(n3723) );
  OR U6395 ( .A(A[378]), .B(B[378]), .Z(n3727) );
  NAND U6396 ( .A(n6760), .B(n6761), .Z(n3762) );
  AND U6397 ( .A(n3785), .B(n3776), .Z(n6761) );
  OR U6398 ( .A(A[369]), .B(B[369]), .Z(n3776) );
  OR U6399 ( .A(A[368]), .B(B[368]), .Z(n3785) );
  AND U6400 ( .A(n3771), .B(n3767), .Z(n6760) );
  OR U6401 ( .A(B[371]), .B(A[371]), .Z(n3767) );
  OR U6402 ( .A(A[370]), .B(B[370]), .Z(n3771) );
  NAND U6403 ( .A(n6762), .B(n6763), .Z(n3303) );
  ANDN U6404 ( .B(n3400), .A(n3497), .Z(n6763) );
  NOR U6405 ( .A(n3590), .B(n6764), .Z(n6762) );
  NAND U6406 ( .A(n6765), .B(n6766), .Z(n3590) );
  AND U6407 ( .A(n6767), .B(n6768), .Z(n6766) );
  AND U6408 ( .A(n3617), .B(n3612), .Z(n6768) );
  AND U6409 ( .A(n3607), .B(n3603), .Z(n6767) );
  ANDN U6410 ( .B(n6769), .A(n3670), .Z(n6765) );
  NAND U6411 ( .A(n6770), .B(n6771), .Z(n3670) );
  AND U6412 ( .A(n3687), .B(n3683), .Z(n6771) );
  OR U6413 ( .A(B[384]), .B(A[384]), .Z(n3687) );
  AND U6414 ( .A(n3678), .B(n3674), .Z(n6770) );
  ANDN U6415 ( .B(n3621), .A(n3643), .Z(n6769) );
  NAND U6416 ( .A(n6772), .B(n6773), .Z(n3301) );
  NAND U6417 ( .A(n6774), .B(n3308), .Z(n6773) );
  NANDN U6418 ( .A(n3310), .B(n6775), .Z(n6774) );
  NAND U6419 ( .A(n6776), .B(n3312), .Z(n6775) );
  NANDN U6420 ( .A(n3314), .B(n6777), .Z(n6776) );
  NAND U6421 ( .A(n6778), .B(n3317), .Z(n6777) );
  NANDN U6422 ( .A(n3319), .B(n6779), .Z(n6778) );
  NAND U6423 ( .A(n6780), .B(n3322), .Z(n6779) );
  NANDN U6424 ( .A(n3324), .B(n6781), .Z(n6780) );
  NANDN U6425 ( .A(n3326), .B(n6782), .Z(n6781) );
  NANDN U6426 ( .A(n3346), .B(n6783), .Z(n6782) );
  NANDN U6427 ( .A(n3348), .B(n3377), .Z(n6783) );
  NANDN U6428 ( .A(n3382), .B(n6784), .Z(n3377) );
  NAND U6429 ( .A(n6785), .B(n3383), .Z(n6784) );
  NANDN U6430 ( .A(n3385), .B(n6786), .Z(n6785) );
  NAND U6431 ( .A(n6787), .B(n3387), .Z(n6786) );
  NANDN U6432 ( .A(n3389), .B(n6788), .Z(n6787) );
  NAND U6433 ( .A(n3392), .B(n3394), .Z(n6788) );
  AND U6434 ( .A(A[432]), .B(B[432]), .Z(n3394) );
  AND U6435 ( .A(A[433]), .B(B[433]), .Z(n3389) );
  AND U6436 ( .A(A[434]), .B(B[434]), .Z(n3385) );
  AND U6437 ( .A(B[435]), .B(A[435]), .Z(n3382) );
  NANDN U6438 ( .A(n3360), .B(n6789), .Z(n3346) );
  NAND U6439 ( .A(n6790), .B(n3361), .Z(n6789) );
  NANDN U6440 ( .A(n3363), .B(n6791), .Z(n6790) );
  NAND U6441 ( .A(n6792), .B(n3365), .Z(n6791) );
  NANDN U6442 ( .A(n3367), .B(n6793), .Z(n6792) );
  NAND U6443 ( .A(n3370), .B(n3372), .Z(n6793) );
  AND U6444 ( .A(A[436]), .B(B[436]), .Z(n3372) );
  AND U6445 ( .A(A[437]), .B(B[437]), .Z(n3367) );
  AND U6446 ( .A(A[438]), .B(B[438]), .Z(n3363) );
  AND U6447 ( .A(B[439]), .B(A[439]), .Z(n3360) );
  NANDN U6448 ( .A(n3330), .B(n6794), .Z(n3324) );
  NAND U6449 ( .A(n6795), .B(n3331), .Z(n6794) );
  NANDN U6450 ( .A(n3333), .B(n6796), .Z(n6795) );
  NAND U6451 ( .A(n6797), .B(n3335), .Z(n6796) );
  NANDN U6452 ( .A(n3337), .B(n6798), .Z(n6797) );
  NAND U6453 ( .A(n3340), .B(n3342), .Z(n6798) );
  AND U6454 ( .A(A[440]), .B(B[440]), .Z(n3342) );
  AND U6455 ( .A(A[441]), .B(B[441]), .Z(n3337) );
  AND U6456 ( .A(A[442]), .B(B[442]), .Z(n3333) );
  AND U6457 ( .A(B[443]), .B(A[443]), .Z(n3330) );
  AND U6458 ( .A(A[444]), .B(B[444]), .Z(n3319) );
  AND U6459 ( .A(A[445]), .B(B[445]), .Z(n3314) );
  AND U6460 ( .A(A[446]), .B(B[446]), .Z(n3310) );
  ANDN U6461 ( .B(n6799), .A(n3307), .Z(n6772) );
  AND U6462 ( .A(B[447]), .B(A[447]), .Z(n3307) );
  NANDN U6463 ( .A(n6764), .B(n6800), .Z(n6799) );
  NANDN U6464 ( .A(n3398), .B(n6801), .Z(n6800) );
  NAND U6465 ( .A(n6802), .B(n3400), .Z(n6801) );
  AND U6466 ( .A(n6803), .B(n6804), .Z(n3400) );
  AND U6467 ( .A(n6805), .B(n6806), .Z(n6804) );
  AND U6468 ( .A(n3424), .B(n3414), .Z(n6806) );
  AND U6469 ( .A(n3409), .B(n3405), .Z(n6805) );
  ANDN U6470 ( .B(n6807), .A(n3472), .Z(n6803) );
  NAND U6471 ( .A(n6808), .B(n6809), .Z(n3472) );
  AND U6472 ( .A(n3493), .B(n3489), .Z(n6809) );
  OR U6473 ( .A(B[416]), .B(A[416]), .Z(n3493) );
  AND U6474 ( .A(n3484), .B(n3480), .Z(n6808) );
  ANDN U6475 ( .B(n3428), .A(n3450), .Z(n6807) );
  NANDN U6476 ( .A(n3495), .B(n6810), .Z(n6802) );
  NANDN U6477 ( .A(n3497), .B(n3589), .Z(n6810) );
  NANDN U6478 ( .A(n3602), .B(n6811), .Z(n3589) );
  NAND U6479 ( .A(n6812), .B(n3603), .Z(n6811) );
  OR U6480 ( .A(B[399]), .B(A[399]), .Z(n3603) );
  NANDN U6481 ( .A(n3605), .B(n6813), .Z(n6812) );
  NAND U6482 ( .A(n6814), .B(n3607), .Z(n6813) );
  OR U6483 ( .A(B[398]), .B(A[398]), .Z(n3607) );
  NANDN U6484 ( .A(n3609), .B(n6815), .Z(n6814) );
  NAND U6485 ( .A(n6816), .B(n3612), .Z(n6815) );
  OR U6486 ( .A(B[397]), .B(A[397]), .Z(n3612) );
  NANDN U6487 ( .A(n3614), .B(n6817), .Z(n6816) );
  NAND U6488 ( .A(n6818), .B(n3617), .Z(n6817) );
  OR U6489 ( .A(B[396]), .B(A[396]), .Z(n3617) );
  NANDN U6490 ( .A(n3619), .B(n6819), .Z(n6818) );
  NAND U6491 ( .A(n6820), .B(n3621), .Z(n6819) );
  AND U6492 ( .A(n6821), .B(n6822), .Z(n3621) );
  AND U6493 ( .A(n3639), .B(n3635), .Z(n6822) );
  OR U6494 ( .A(B[392]), .B(A[392]), .Z(n3639) );
  AND U6495 ( .A(n3630), .B(n3626), .Z(n6821) );
  NANDN U6496 ( .A(n3641), .B(n6823), .Z(n6820) );
  NANDN U6497 ( .A(n3643), .B(n3669), .Z(n6823) );
  NANDN U6498 ( .A(n3673), .B(n6824), .Z(n3669) );
  NAND U6499 ( .A(n6825), .B(n3674), .Z(n6824) );
  OR U6500 ( .A(B[387]), .B(A[387]), .Z(n3674) );
  NANDN U6501 ( .A(n3676), .B(n6826), .Z(n6825) );
  NAND U6502 ( .A(n6827), .B(n3678), .Z(n6826) );
  OR U6503 ( .A(B[386]), .B(A[386]), .Z(n3678) );
  NANDN U6504 ( .A(n3680), .B(n6828), .Z(n6827) );
  NAND U6505 ( .A(n3683), .B(n3685), .Z(n6828) );
  AND U6506 ( .A(B[384]), .B(A[384]), .Z(n3685) );
  OR U6507 ( .A(B[385]), .B(A[385]), .Z(n3683) );
  AND U6508 ( .A(B[385]), .B(A[385]), .Z(n3680) );
  AND U6509 ( .A(B[386]), .B(A[386]), .Z(n3676) );
  AND U6510 ( .A(B[387]), .B(A[387]), .Z(n3673) );
  NAND U6511 ( .A(n6829), .B(n6830), .Z(n3643) );
  AND U6512 ( .A(n3666), .B(n3657), .Z(n6830) );
  OR U6513 ( .A(B[388]), .B(A[388]), .Z(n3666) );
  AND U6514 ( .A(n3652), .B(n3648), .Z(n6829) );
  NANDN U6515 ( .A(n3647), .B(n6831), .Z(n3641) );
  NAND U6516 ( .A(n6832), .B(n3648), .Z(n6831) );
  OR U6517 ( .A(B[391]), .B(A[391]), .Z(n3648) );
  NANDN U6518 ( .A(n3650), .B(n6833), .Z(n6832) );
  NAND U6519 ( .A(n6834), .B(n3652), .Z(n6833) );
  OR U6520 ( .A(B[390]), .B(A[390]), .Z(n3652) );
  NANDN U6521 ( .A(n3654), .B(n6835), .Z(n6834) );
  NAND U6522 ( .A(n3657), .B(n3664), .Z(n6835) );
  AND U6523 ( .A(B[388]), .B(A[388]), .Z(n3664) );
  OR U6524 ( .A(B[389]), .B(A[389]), .Z(n3657) );
  AND U6525 ( .A(B[389]), .B(A[389]), .Z(n3654) );
  AND U6526 ( .A(B[390]), .B(A[390]), .Z(n3650) );
  AND U6527 ( .A(B[391]), .B(A[391]), .Z(n3647) );
  NANDN U6528 ( .A(n3625), .B(n6836), .Z(n3619) );
  NAND U6529 ( .A(n6837), .B(n3626), .Z(n6836) );
  OR U6530 ( .A(B[395]), .B(A[395]), .Z(n3626) );
  NANDN U6531 ( .A(n3628), .B(n6838), .Z(n6837) );
  NAND U6532 ( .A(n6839), .B(n3630), .Z(n6838) );
  OR U6533 ( .A(B[394]), .B(A[394]), .Z(n3630) );
  NANDN U6534 ( .A(n3632), .B(n6840), .Z(n6839) );
  NAND U6535 ( .A(n3635), .B(n3637), .Z(n6840) );
  AND U6536 ( .A(B[392]), .B(A[392]), .Z(n3637) );
  OR U6537 ( .A(B[393]), .B(A[393]), .Z(n3635) );
  AND U6538 ( .A(B[393]), .B(A[393]), .Z(n3632) );
  AND U6539 ( .A(B[394]), .B(A[394]), .Z(n3628) );
  AND U6540 ( .A(B[395]), .B(A[395]), .Z(n3625) );
  AND U6541 ( .A(B[396]), .B(A[396]), .Z(n3614) );
  AND U6542 ( .A(B[397]), .B(A[397]), .Z(n3609) );
  AND U6543 ( .A(B[398]), .B(A[398]), .Z(n3605) );
  AND U6544 ( .A(B[399]), .B(A[399]), .Z(n3602) );
  NAND U6545 ( .A(n6841), .B(n6842), .Z(n3497) );
  AND U6546 ( .A(n6843), .B(n6844), .Z(n6842) );
  AND U6547 ( .A(n3516), .B(n3511), .Z(n6844) );
  AND U6548 ( .A(n3506), .B(n3502), .Z(n6843) );
  ANDN U6549 ( .B(n6845), .A(n3569), .Z(n6841) );
  NAND U6550 ( .A(n6846), .B(n6847), .Z(n3569) );
  AND U6551 ( .A(n3586), .B(n3582), .Z(n6847) );
  OR U6552 ( .A(B[400]), .B(A[400]), .Z(n3586) );
  AND U6553 ( .A(n3577), .B(n3573), .Z(n6846) );
  ANDN U6554 ( .B(n3520), .A(n3547), .Z(n6845) );
  NANDN U6555 ( .A(n3501), .B(n6848), .Z(n3495) );
  NAND U6556 ( .A(n6849), .B(n3502), .Z(n6848) );
  OR U6557 ( .A(B[415]), .B(A[415]), .Z(n3502) );
  NANDN U6558 ( .A(n3504), .B(n6850), .Z(n6849) );
  NAND U6559 ( .A(n6851), .B(n3506), .Z(n6850) );
  OR U6560 ( .A(B[414]), .B(A[414]), .Z(n3506) );
  NANDN U6561 ( .A(n3508), .B(n6852), .Z(n6851) );
  NAND U6562 ( .A(n6853), .B(n3511), .Z(n6852) );
  OR U6563 ( .A(B[413]), .B(A[413]), .Z(n3511) );
  NANDN U6564 ( .A(n3513), .B(n6854), .Z(n6853) );
  NAND U6565 ( .A(n6855), .B(n3516), .Z(n6854) );
  OR U6566 ( .A(B[412]), .B(A[412]), .Z(n3516) );
  NANDN U6567 ( .A(n3518), .B(n6856), .Z(n6855) );
  NAND U6568 ( .A(n6857), .B(n3520), .Z(n6856) );
  AND U6569 ( .A(n6858), .B(n6859), .Z(n3520) );
  AND U6570 ( .A(n3543), .B(n3534), .Z(n6859) );
  OR U6571 ( .A(B[408]), .B(A[408]), .Z(n3543) );
  AND U6572 ( .A(n3529), .B(n3525), .Z(n6858) );
  NANDN U6573 ( .A(n3545), .B(n6860), .Z(n6857) );
  NANDN U6574 ( .A(n3547), .B(n3568), .Z(n6860) );
  NANDN U6575 ( .A(n3572), .B(n6861), .Z(n3568) );
  NAND U6576 ( .A(n6862), .B(n3573), .Z(n6861) );
  OR U6577 ( .A(B[403]), .B(A[403]), .Z(n3573) );
  NANDN U6578 ( .A(n3575), .B(n6863), .Z(n6862) );
  NAND U6579 ( .A(n6864), .B(n3577), .Z(n6863) );
  OR U6580 ( .A(B[402]), .B(A[402]), .Z(n3577) );
  NANDN U6581 ( .A(n3579), .B(n6865), .Z(n6864) );
  NAND U6582 ( .A(n3582), .B(n3584), .Z(n6865) );
  AND U6583 ( .A(B[400]), .B(A[400]), .Z(n3584) );
  OR U6584 ( .A(B[401]), .B(A[401]), .Z(n3582) );
  AND U6585 ( .A(B[401]), .B(A[401]), .Z(n3579) );
  AND U6586 ( .A(B[402]), .B(A[402]), .Z(n3575) );
  AND U6587 ( .A(B[403]), .B(A[403]), .Z(n3572) );
  NAND U6588 ( .A(n6866), .B(n6867), .Z(n3547) );
  AND U6589 ( .A(n3565), .B(n3561), .Z(n6867) );
  OR U6590 ( .A(B[404]), .B(A[404]), .Z(n3565) );
  AND U6591 ( .A(n3556), .B(n3552), .Z(n6866) );
  NANDN U6592 ( .A(n3551), .B(n6868), .Z(n3545) );
  NAND U6593 ( .A(n6869), .B(n3552), .Z(n6868) );
  OR U6594 ( .A(B[407]), .B(A[407]), .Z(n3552) );
  NANDN U6595 ( .A(n3554), .B(n6870), .Z(n6869) );
  NAND U6596 ( .A(n6871), .B(n3556), .Z(n6870) );
  OR U6597 ( .A(B[406]), .B(A[406]), .Z(n3556) );
  NANDN U6598 ( .A(n3558), .B(n6872), .Z(n6871) );
  NAND U6599 ( .A(n3561), .B(n3563), .Z(n6872) );
  AND U6600 ( .A(B[404]), .B(A[404]), .Z(n3563) );
  OR U6601 ( .A(B[405]), .B(A[405]), .Z(n3561) );
  AND U6602 ( .A(B[405]), .B(A[405]), .Z(n3558) );
  AND U6603 ( .A(B[406]), .B(A[406]), .Z(n3554) );
  AND U6604 ( .A(B[407]), .B(A[407]), .Z(n3551) );
  NANDN U6605 ( .A(n3524), .B(n6873), .Z(n3518) );
  NAND U6606 ( .A(n6874), .B(n3525), .Z(n6873) );
  OR U6607 ( .A(B[411]), .B(A[411]), .Z(n3525) );
  NANDN U6608 ( .A(n3527), .B(n6875), .Z(n6874) );
  NAND U6609 ( .A(n6876), .B(n3529), .Z(n6875) );
  OR U6610 ( .A(B[410]), .B(A[410]), .Z(n3529) );
  NANDN U6611 ( .A(n3531), .B(n6877), .Z(n6876) );
  NAND U6612 ( .A(n3534), .B(n3541), .Z(n6877) );
  AND U6613 ( .A(B[408]), .B(A[408]), .Z(n3541) );
  OR U6614 ( .A(B[409]), .B(A[409]), .Z(n3534) );
  AND U6615 ( .A(B[409]), .B(A[409]), .Z(n3531) );
  AND U6616 ( .A(B[410]), .B(A[410]), .Z(n3527) );
  AND U6617 ( .A(B[411]), .B(A[411]), .Z(n3524) );
  AND U6618 ( .A(B[412]), .B(A[412]), .Z(n3513) );
  AND U6619 ( .A(B[413]), .B(A[413]), .Z(n3508) );
  AND U6620 ( .A(B[414]), .B(A[414]), .Z(n3504) );
  AND U6621 ( .A(B[415]), .B(A[415]), .Z(n3501) );
  NANDN U6622 ( .A(n3404), .B(n6878), .Z(n3398) );
  NAND U6623 ( .A(n6879), .B(n3405), .Z(n6878) );
  OR U6624 ( .A(B[431]), .B(A[431]), .Z(n3405) );
  NANDN U6625 ( .A(n3407), .B(n6880), .Z(n6879) );
  NAND U6626 ( .A(n6881), .B(n3409), .Z(n6880) );
  OR U6627 ( .A(B[430]), .B(A[430]), .Z(n3409) );
  NANDN U6628 ( .A(n3411), .B(n6882), .Z(n6881) );
  NAND U6629 ( .A(n6883), .B(n3414), .Z(n6882) );
  OR U6630 ( .A(B[429]), .B(A[429]), .Z(n3414) );
  NANDN U6631 ( .A(n3421), .B(n6884), .Z(n6883) );
  NAND U6632 ( .A(n6885), .B(n3424), .Z(n6884) );
  OR U6633 ( .A(B[428]), .B(A[428]), .Z(n3424) );
  NANDN U6634 ( .A(n3426), .B(n6886), .Z(n6885) );
  NAND U6635 ( .A(n6887), .B(n3428), .Z(n6886) );
  AND U6636 ( .A(n6888), .B(n6889), .Z(n3428) );
  AND U6637 ( .A(n3446), .B(n3442), .Z(n6889) );
  OR U6638 ( .A(B[424]), .B(A[424]), .Z(n3446) );
  AND U6639 ( .A(n3437), .B(n3433), .Z(n6888) );
  NANDN U6640 ( .A(n3448), .B(n6890), .Z(n6887) );
  NANDN U6641 ( .A(n3450), .B(n3471), .Z(n6890) );
  NANDN U6642 ( .A(n3479), .B(n6891), .Z(n3471) );
  NAND U6643 ( .A(n6892), .B(n3480), .Z(n6891) );
  OR U6644 ( .A(B[419]), .B(A[419]), .Z(n3480) );
  NANDN U6645 ( .A(n3482), .B(n6893), .Z(n6892) );
  NAND U6646 ( .A(n6894), .B(n3484), .Z(n6893) );
  OR U6647 ( .A(B[418]), .B(A[418]), .Z(n3484) );
  NANDN U6648 ( .A(n3486), .B(n6895), .Z(n6894) );
  NAND U6649 ( .A(n3489), .B(n3491), .Z(n6895) );
  AND U6650 ( .A(B[416]), .B(A[416]), .Z(n3491) );
  OR U6651 ( .A(B[417]), .B(A[417]), .Z(n3489) );
  AND U6652 ( .A(B[417]), .B(A[417]), .Z(n3486) );
  AND U6653 ( .A(B[418]), .B(A[418]), .Z(n3482) );
  AND U6654 ( .A(B[419]), .B(A[419]), .Z(n3479) );
  NAND U6655 ( .A(n6896), .B(n6897), .Z(n3450) );
  AND U6656 ( .A(n3468), .B(n3464), .Z(n6897) );
  OR U6657 ( .A(B[420]), .B(A[420]), .Z(n3468) );
  AND U6658 ( .A(n3459), .B(n3455), .Z(n6896) );
  NANDN U6659 ( .A(n3454), .B(n6898), .Z(n3448) );
  NAND U6660 ( .A(n6899), .B(n3455), .Z(n6898) );
  OR U6661 ( .A(B[423]), .B(A[423]), .Z(n3455) );
  NANDN U6662 ( .A(n3457), .B(n6900), .Z(n6899) );
  NAND U6663 ( .A(n6901), .B(n3459), .Z(n6900) );
  OR U6664 ( .A(B[422]), .B(A[422]), .Z(n3459) );
  NANDN U6665 ( .A(n3461), .B(n6902), .Z(n6901) );
  NAND U6666 ( .A(n3464), .B(n3466), .Z(n6902) );
  AND U6667 ( .A(B[420]), .B(A[420]), .Z(n3466) );
  OR U6668 ( .A(B[421]), .B(A[421]), .Z(n3464) );
  AND U6669 ( .A(B[421]), .B(A[421]), .Z(n3461) );
  AND U6670 ( .A(B[422]), .B(A[422]), .Z(n3457) );
  AND U6671 ( .A(B[423]), .B(A[423]), .Z(n3454) );
  NANDN U6672 ( .A(n3432), .B(n6903), .Z(n3426) );
  NAND U6673 ( .A(n6904), .B(n3433), .Z(n6903) );
  OR U6674 ( .A(B[427]), .B(A[427]), .Z(n3433) );
  NANDN U6675 ( .A(n3435), .B(n6905), .Z(n6904) );
  NAND U6676 ( .A(n6906), .B(n3437), .Z(n6905) );
  OR U6677 ( .A(B[426]), .B(A[426]), .Z(n3437) );
  NANDN U6678 ( .A(n3439), .B(n6907), .Z(n6906) );
  NAND U6679 ( .A(n3442), .B(n3444), .Z(n6907) );
  AND U6680 ( .A(B[424]), .B(A[424]), .Z(n3444) );
  OR U6681 ( .A(B[425]), .B(A[425]), .Z(n3442) );
  AND U6682 ( .A(B[425]), .B(A[425]), .Z(n3439) );
  AND U6683 ( .A(B[426]), .B(A[426]), .Z(n3435) );
  AND U6684 ( .A(B[427]), .B(A[427]), .Z(n3432) );
  AND U6685 ( .A(B[428]), .B(A[428]), .Z(n3421) );
  AND U6686 ( .A(B[429]), .B(A[429]), .Z(n3411) );
  AND U6687 ( .A(B[430]), .B(A[430]), .Z(n3407) );
  AND U6688 ( .A(B[431]), .B(A[431]), .Z(n3404) );
  NAND U6689 ( .A(n6908), .B(n6909), .Z(n6764) );
  AND U6690 ( .A(n6910), .B(n6911), .Z(n6909) );
  AND U6691 ( .A(n3322), .B(n3317), .Z(n6911) );
  OR U6692 ( .A(A[445]), .B(B[445]), .Z(n3317) );
  OR U6693 ( .A(A[444]), .B(B[444]), .Z(n3322) );
  AND U6694 ( .A(n3312), .B(n3308), .Z(n6910) );
  OR U6695 ( .A(B[447]), .B(A[447]), .Z(n3308) );
  OR U6696 ( .A(A[446]), .B(B[446]), .Z(n3312) );
  ANDN U6697 ( .B(n6912), .A(n3348), .Z(n6908) );
  NAND U6698 ( .A(n6913), .B(n6914), .Z(n3348) );
  AND U6699 ( .A(n3374), .B(n3370), .Z(n6914) );
  OR U6700 ( .A(A[437]), .B(B[437]), .Z(n3370) );
  OR U6701 ( .A(A[436]), .B(B[436]), .Z(n3374) );
  AND U6702 ( .A(n3365), .B(n3361), .Z(n6913) );
  OR U6703 ( .A(B[439]), .B(A[439]), .Z(n3361) );
  OR U6704 ( .A(A[438]), .B(B[438]), .Z(n3365) );
  NOR U6705 ( .A(n3378), .B(n3326), .Z(n6912) );
  NAND U6706 ( .A(n6915), .B(n6916), .Z(n3326) );
  AND U6707 ( .A(n3344), .B(n3340), .Z(n6916) );
  OR U6708 ( .A(A[441]), .B(B[441]), .Z(n3340) );
  OR U6709 ( .A(A[440]), .B(B[440]), .Z(n3344) );
  AND U6710 ( .A(n3335), .B(n3331), .Z(n6915) );
  OR U6711 ( .A(B[443]), .B(A[443]), .Z(n3331) );
  OR U6712 ( .A(A[442]), .B(B[442]), .Z(n3335) );
  NAND U6713 ( .A(n6917), .B(n6918), .Z(n3378) );
  AND U6714 ( .A(n3396), .B(n3392), .Z(n6918) );
  OR U6715 ( .A(A[433]), .B(B[433]), .Z(n3392) );
  OR U6716 ( .A(A[432]), .B(B[432]), .Z(n3396) );
  AND U6717 ( .A(n3387), .B(n3383), .Z(n6917) );
  OR U6718 ( .A(B[435]), .B(A[435]), .Z(n3383) );
  OR U6719 ( .A(A[434]), .B(B[434]), .Z(n3387) );
  NAND U6720 ( .A(n6919), .B(n6920), .Z(n3205) );
  AND U6721 ( .A(n6921), .B(n6922), .Z(n6920) );
  AND U6722 ( .A(n3224), .B(n3219), .Z(n6922) );
  AND U6723 ( .A(n3214), .B(n3210), .Z(n6921) );
  ANDN U6724 ( .B(n6923), .A(n3277), .Z(n6919) );
  NAND U6725 ( .A(n6924), .B(n6925), .Z(n3277) );
  AND U6726 ( .A(n3299), .B(n3290), .Z(n6925) );
  OR U6727 ( .A(B[448]), .B(A[448]), .Z(n3299) );
  AND U6728 ( .A(n3285), .B(n3281), .Z(n6924) );
  ANDN U6729 ( .B(n3228), .A(n3255), .Z(n6923) );
  NANDN U6730 ( .A(n3209), .B(n6926), .Z(n3203) );
  NAND U6731 ( .A(n6927), .B(n3210), .Z(n6926) );
  OR U6732 ( .A(B[463]), .B(A[463]), .Z(n3210) );
  NANDN U6733 ( .A(n3212), .B(n6928), .Z(n6927) );
  NAND U6734 ( .A(n6929), .B(n3214), .Z(n6928) );
  OR U6735 ( .A(B[462]), .B(A[462]), .Z(n3214) );
  NANDN U6736 ( .A(n3216), .B(n6930), .Z(n6929) );
  NAND U6737 ( .A(n6931), .B(n3219), .Z(n6930) );
  OR U6738 ( .A(B[461]), .B(A[461]), .Z(n3219) );
  NANDN U6739 ( .A(n3221), .B(n6932), .Z(n6931) );
  NAND U6740 ( .A(n6933), .B(n3224), .Z(n6932) );
  OR U6741 ( .A(B[460]), .B(A[460]), .Z(n3224) );
  NANDN U6742 ( .A(n3226), .B(n6934), .Z(n6933) );
  NAND U6743 ( .A(n6935), .B(n3228), .Z(n6934) );
  AND U6744 ( .A(n6936), .B(n6937), .Z(n3228) );
  AND U6745 ( .A(n3251), .B(n3247), .Z(n6937) );
  OR U6746 ( .A(B[456]), .B(A[456]), .Z(n3251) );
  AND U6747 ( .A(n3242), .B(n3238), .Z(n6936) );
  NANDN U6748 ( .A(n3253), .B(n6938), .Z(n6935) );
  NANDN U6749 ( .A(n3255), .B(n3276), .Z(n6938) );
  NANDN U6750 ( .A(n3280), .B(n6939), .Z(n3276) );
  NAND U6751 ( .A(n6940), .B(n3281), .Z(n6939) );
  OR U6752 ( .A(B[451]), .B(A[451]), .Z(n3281) );
  NANDN U6753 ( .A(n3283), .B(n6941), .Z(n6940) );
  NAND U6754 ( .A(n6942), .B(n3285), .Z(n6941) );
  OR U6755 ( .A(B[450]), .B(A[450]), .Z(n3285) );
  NANDN U6756 ( .A(n3287), .B(n6943), .Z(n6942) );
  NAND U6757 ( .A(n3290), .B(n3297), .Z(n6943) );
  AND U6758 ( .A(B[448]), .B(A[448]), .Z(n3297) );
  OR U6759 ( .A(B[449]), .B(A[449]), .Z(n3290) );
  AND U6760 ( .A(B[449]), .B(A[449]), .Z(n3287) );
  AND U6761 ( .A(B[450]), .B(A[450]), .Z(n3283) );
  AND U6762 ( .A(B[451]), .B(A[451]), .Z(n3280) );
  NAND U6763 ( .A(n6944), .B(n6945), .Z(n3255) );
  AND U6764 ( .A(n3273), .B(n3269), .Z(n6945) );
  OR U6765 ( .A(B[452]), .B(A[452]), .Z(n3273) );
  AND U6766 ( .A(n3264), .B(n3260), .Z(n6944) );
  NANDN U6767 ( .A(n3259), .B(n6946), .Z(n3253) );
  NAND U6768 ( .A(n6947), .B(n3260), .Z(n6946) );
  OR U6769 ( .A(B[455]), .B(A[455]), .Z(n3260) );
  NANDN U6770 ( .A(n3262), .B(n6948), .Z(n6947) );
  NAND U6771 ( .A(n6949), .B(n3264), .Z(n6948) );
  OR U6772 ( .A(B[454]), .B(A[454]), .Z(n3264) );
  NANDN U6773 ( .A(n3266), .B(n6950), .Z(n6949) );
  NAND U6774 ( .A(n3269), .B(n3271), .Z(n6950) );
  AND U6775 ( .A(B[452]), .B(A[452]), .Z(n3271) );
  OR U6776 ( .A(B[453]), .B(A[453]), .Z(n3269) );
  AND U6777 ( .A(B[453]), .B(A[453]), .Z(n3266) );
  AND U6778 ( .A(B[454]), .B(A[454]), .Z(n3262) );
  AND U6779 ( .A(B[455]), .B(A[455]), .Z(n3259) );
  NANDN U6780 ( .A(n3237), .B(n6951), .Z(n3226) );
  NAND U6781 ( .A(n6952), .B(n3238), .Z(n6951) );
  OR U6782 ( .A(B[459]), .B(A[459]), .Z(n3238) );
  NANDN U6783 ( .A(n3240), .B(n6953), .Z(n6952) );
  NAND U6784 ( .A(n6954), .B(n3242), .Z(n6953) );
  OR U6785 ( .A(B[458]), .B(A[458]), .Z(n3242) );
  NANDN U6786 ( .A(n3244), .B(n6955), .Z(n6954) );
  NAND U6787 ( .A(n3247), .B(n3249), .Z(n6955) );
  AND U6788 ( .A(B[456]), .B(A[456]), .Z(n3249) );
  OR U6789 ( .A(B[457]), .B(A[457]), .Z(n3247) );
  AND U6790 ( .A(B[457]), .B(A[457]), .Z(n3244) );
  AND U6791 ( .A(B[458]), .B(A[458]), .Z(n3240) );
  AND U6792 ( .A(B[459]), .B(A[459]), .Z(n3237) );
  AND U6793 ( .A(B[460]), .B(A[460]), .Z(n3221) );
  AND U6794 ( .A(B[461]), .B(A[461]), .Z(n3216) );
  AND U6795 ( .A(B[462]), .B(A[462]), .Z(n3212) );
  AND U6796 ( .A(B[463]), .B(A[463]), .Z(n3209) );
  NAND U6797 ( .A(n6956), .B(n6957), .Z(n3104) );
  AND U6798 ( .A(n6958), .B(n6959), .Z(n6957) );
  AND U6799 ( .A(n3131), .B(n3126), .Z(n6959) );
  AND U6800 ( .A(n3121), .B(n3117), .Z(n6958) );
  ANDN U6801 ( .B(n6960), .A(n3184), .Z(n6956) );
  NAND U6802 ( .A(n6961), .B(n6962), .Z(n3184) );
  AND U6803 ( .A(n3201), .B(n3197), .Z(n6962) );
  OR U6804 ( .A(B[464]), .B(A[464]), .Z(n3201) );
  AND U6805 ( .A(n3192), .B(n3188), .Z(n6961) );
  ANDN U6806 ( .B(n3135), .A(n3157), .Z(n6960) );
  NANDN U6807 ( .A(n3116), .B(n6963), .Z(n3102) );
  NAND U6808 ( .A(n6964), .B(n3117), .Z(n6963) );
  OR U6809 ( .A(B[479]), .B(A[479]), .Z(n3117) );
  NANDN U6810 ( .A(n3119), .B(n6965), .Z(n6964) );
  NAND U6811 ( .A(n6966), .B(n3121), .Z(n6965) );
  OR U6812 ( .A(B[478]), .B(A[478]), .Z(n3121) );
  NANDN U6813 ( .A(n3123), .B(n6967), .Z(n6966) );
  NAND U6814 ( .A(n6968), .B(n3126), .Z(n6967) );
  OR U6815 ( .A(B[477]), .B(A[477]), .Z(n3126) );
  NANDN U6816 ( .A(n3128), .B(n6969), .Z(n6968) );
  NAND U6817 ( .A(n6970), .B(n3131), .Z(n6969) );
  OR U6818 ( .A(B[476]), .B(A[476]), .Z(n3131) );
  NANDN U6819 ( .A(n3133), .B(n6971), .Z(n6970) );
  NAND U6820 ( .A(n6972), .B(n3135), .Z(n6971) );
  AND U6821 ( .A(n6973), .B(n6974), .Z(n3135) );
  AND U6822 ( .A(n3153), .B(n3149), .Z(n6974) );
  OR U6823 ( .A(B[472]), .B(A[472]), .Z(n3153) );
  AND U6824 ( .A(n3144), .B(n3140), .Z(n6973) );
  NANDN U6825 ( .A(n3155), .B(n6975), .Z(n6972) );
  NANDN U6826 ( .A(n3157), .B(n3183), .Z(n6975) );
  NANDN U6827 ( .A(n3187), .B(n6976), .Z(n3183) );
  NAND U6828 ( .A(n6977), .B(n3188), .Z(n6976) );
  OR U6829 ( .A(B[467]), .B(A[467]), .Z(n3188) );
  NANDN U6830 ( .A(n3190), .B(n6978), .Z(n6977) );
  NAND U6831 ( .A(n6979), .B(n3192), .Z(n6978) );
  OR U6832 ( .A(B[466]), .B(A[466]), .Z(n3192) );
  NANDN U6833 ( .A(n3194), .B(n6980), .Z(n6979) );
  NAND U6834 ( .A(n3197), .B(n3199), .Z(n6980) );
  AND U6835 ( .A(B[464]), .B(A[464]), .Z(n3199) );
  OR U6836 ( .A(B[465]), .B(A[465]), .Z(n3197) );
  AND U6837 ( .A(B[465]), .B(A[465]), .Z(n3194) );
  AND U6838 ( .A(B[466]), .B(A[466]), .Z(n3190) );
  AND U6839 ( .A(B[467]), .B(A[467]), .Z(n3187) );
  NAND U6840 ( .A(n6981), .B(n6982), .Z(n3157) );
  AND U6841 ( .A(n3180), .B(n3171), .Z(n6982) );
  OR U6842 ( .A(B[468]), .B(A[468]), .Z(n3180) );
  AND U6843 ( .A(n3166), .B(n3162), .Z(n6981) );
  NANDN U6844 ( .A(n3161), .B(n6983), .Z(n3155) );
  NAND U6845 ( .A(n6984), .B(n3162), .Z(n6983) );
  OR U6846 ( .A(B[471]), .B(A[471]), .Z(n3162) );
  NANDN U6847 ( .A(n3164), .B(n6985), .Z(n6984) );
  NAND U6848 ( .A(n6986), .B(n3166), .Z(n6985) );
  OR U6849 ( .A(B[470]), .B(A[470]), .Z(n3166) );
  NANDN U6850 ( .A(n3168), .B(n6987), .Z(n6986) );
  NAND U6851 ( .A(n3171), .B(n3178), .Z(n6987) );
  AND U6852 ( .A(B[468]), .B(A[468]), .Z(n3178) );
  OR U6853 ( .A(B[469]), .B(A[469]), .Z(n3171) );
  AND U6854 ( .A(B[469]), .B(A[469]), .Z(n3168) );
  AND U6855 ( .A(B[470]), .B(A[470]), .Z(n3164) );
  AND U6856 ( .A(B[471]), .B(A[471]), .Z(n3161) );
  NANDN U6857 ( .A(n3139), .B(n6988), .Z(n3133) );
  NAND U6858 ( .A(n6989), .B(n3140), .Z(n6988) );
  OR U6859 ( .A(B[475]), .B(A[475]), .Z(n3140) );
  NANDN U6860 ( .A(n3142), .B(n6990), .Z(n6989) );
  NAND U6861 ( .A(n6991), .B(n3144), .Z(n6990) );
  OR U6862 ( .A(B[474]), .B(A[474]), .Z(n3144) );
  NANDN U6863 ( .A(n3146), .B(n6992), .Z(n6991) );
  NAND U6864 ( .A(n3149), .B(n3151), .Z(n6992) );
  AND U6865 ( .A(B[472]), .B(A[472]), .Z(n3151) );
  OR U6866 ( .A(B[473]), .B(A[473]), .Z(n3149) );
  AND U6867 ( .A(B[473]), .B(A[473]), .Z(n3146) );
  AND U6868 ( .A(B[474]), .B(A[474]), .Z(n3142) );
  AND U6869 ( .A(B[475]), .B(A[475]), .Z(n3139) );
  AND U6870 ( .A(B[476]), .B(A[476]), .Z(n3128) );
  AND U6871 ( .A(B[477]), .B(A[477]), .Z(n3123) );
  AND U6872 ( .A(B[478]), .B(A[478]), .Z(n3119) );
  AND U6873 ( .A(B[479]), .B(A[479]), .Z(n3116) );
  NAND U6874 ( .A(n6993), .B(n6994), .Z(n3015) );
  AND U6875 ( .A(n6995), .B(n6996), .Z(n6994) );
  AND U6876 ( .A(n3034), .B(n3029), .Z(n6996) );
  AND U6877 ( .A(n3024), .B(n3020), .Z(n6995) );
  ANDN U6878 ( .B(n6997), .A(n3083), .Z(n6993) );
  NAND U6879 ( .A(n6998), .B(n6999), .Z(n3083) );
  AND U6880 ( .A(n3100), .B(n3096), .Z(n6999) );
  OR U6881 ( .A(B[480]), .B(A[480]), .Z(n3100) );
  AND U6882 ( .A(n3091), .B(n3087), .Z(n6998) );
  ANDN U6883 ( .B(n3038), .A(n3061), .Z(n6997) );
  NANDN U6884 ( .A(n3019), .B(n7000), .Z(n3013) );
  NAND U6885 ( .A(n7001), .B(n3020), .Z(n7000) );
  OR U6886 ( .A(B[495]), .B(A[495]), .Z(n3020) );
  NANDN U6887 ( .A(n3022), .B(n7002), .Z(n7001) );
  NAND U6888 ( .A(n7003), .B(n3024), .Z(n7002) );
  OR U6889 ( .A(B[494]), .B(A[494]), .Z(n3024) );
  NANDN U6890 ( .A(n3026), .B(n7004), .Z(n7003) );
  NAND U6891 ( .A(n7005), .B(n3029), .Z(n7004) );
  OR U6892 ( .A(B[493]), .B(A[493]), .Z(n3029) );
  NANDN U6893 ( .A(n3031), .B(n7006), .Z(n7005) );
  NAND U6894 ( .A(n7007), .B(n3034), .Z(n7006) );
  OR U6895 ( .A(B[492]), .B(A[492]), .Z(n3034) );
  NANDN U6896 ( .A(n3036), .B(n7008), .Z(n7007) );
  NAND U6897 ( .A(n7009), .B(n3038), .Z(n7008) );
  AND U6898 ( .A(n7010), .B(n7011), .Z(n3038) );
  AND U6899 ( .A(n3057), .B(n3052), .Z(n7011) );
  OR U6900 ( .A(B[488]), .B(A[488]), .Z(n3057) );
  AND U6901 ( .A(n3047), .B(n3043), .Z(n7010) );
  NANDN U6902 ( .A(n3059), .B(n7012), .Z(n7009) );
  NANDN U6903 ( .A(n3061), .B(n3082), .Z(n7012) );
  NANDN U6904 ( .A(n3086), .B(n7013), .Z(n3082) );
  NAND U6905 ( .A(n7014), .B(n3087), .Z(n7013) );
  OR U6906 ( .A(B[483]), .B(A[483]), .Z(n3087) );
  NANDN U6907 ( .A(n3089), .B(n7015), .Z(n7014) );
  NAND U6908 ( .A(n7016), .B(n3091), .Z(n7015) );
  OR U6909 ( .A(B[482]), .B(A[482]), .Z(n3091) );
  NANDN U6910 ( .A(n3093), .B(n7017), .Z(n7016) );
  NAND U6911 ( .A(n3096), .B(n3098), .Z(n7017) );
  AND U6912 ( .A(B[480]), .B(A[480]), .Z(n3098) );
  OR U6913 ( .A(B[481]), .B(A[481]), .Z(n3096) );
  AND U6914 ( .A(B[481]), .B(A[481]), .Z(n3093) );
  AND U6915 ( .A(B[482]), .B(A[482]), .Z(n3089) );
  AND U6916 ( .A(B[483]), .B(A[483]), .Z(n3086) );
  NAND U6917 ( .A(n7018), .B(n7019), .Z(n3061) );
  AND U6918 ( .A(n3079), .B(n3075), .Z(n7019) );
  OR U6919 ( .A(B[484]), .B(A[484]), .Z(n3079) );
  AND U6920 ( .A(n3070), .B(n3066), .Z(n7018) );
  NANDN U6921 ( .A(n3065), .B(n7020), .Z(n3059) );
  NAND U6922 ( .A(n7021), .B(n3066), .Z(n7020) );
  OR U6923 ( .A(B[487]), .B(A[487]), .Z(n3066) );
  NANDN U6924 ( .A(n3068), .B(n7022), .Z(n7021) );
  NAND U6925 ( .A(n7023), .B(n3070), .Z(n7022) );
  OR U6926 ( .A(B[486]), .B(A[486]), .Z(n3070) );
  NANDN U6927 ( .A(n3072), .B(n7024), .Z(n7023) );
  NAND U6928 ( .A(n3075), .B(n3077), .Z(n7024) );
  AND U6929 ( .A(B[484]), .B(A[484]), .Z(n3077) );
  OR U6930 ( .A(B[485]), .B(A[485]), .Z(n3075) );
  AND U6931 ( .A(B[485]), .B(A[485]), .Z(n3072) );
  AND U6932 ( .A(B[486]), .B(A[486]), .Z(n3068) );
  AND U6933 ( .A(B[487]), .B(A[487]), .Z(n3065) );
  NANDN U6934 ( .A(n3042), .B(n7025), .Z(n3036) );
  NAND U6935 ( .A(n7026), .B(n3043), .Z(n7025) );
  OR U6936 ( .A(B[491]), .B(A[491]), .Z(n3043) );
  NANDN U6937 ( .A(n3045), .B(n7027), .Z(n7026) );
  NAND U6938 ( .A(n7028), .B(n3047), .Z(n7027) );
  OR U6939 ( .A(B[490]), .B(A[490]), .Z(n3047) );
  NANDN U6940 ( .A(n3049), .B(n7029), .Z(n7028) );
  NAND U6941 ( .A(n3052), .B(n3055), .Z(n7029) );
  AND U6942 ( .A(B[488]), .B(A[488]), .Z(n3055) );
  OR U6943 ( .A(B[489]), .B(A[489]), .Z(n3052) );
  AND U6944 ( .A(B[489]), .B(A[489]), .Z(n3049) );
  AND U6945 ( .A(B[490]), .B(A[490]), .Z(n3045) );
  AND U6946 ( .A(B[491]), .B(A[491]), .Z(n3042) );
  AND U6947 ( .A(B[492]), .B(A[492]), .Z(n3031) );
  AND U6948 ( .A(B[493]), .B(A[493]), .Z(n3026) );
  AND U6949 ( .A(B[494]), .B(A[494]), .Z(n3022) );
  AND U6950 ( .A(B[495]), .B(A[495]), .Z(n3019) );
  ANDN U6951 ( .B(n7030), .A(n2984), .Z(n5845) );
  NAND U6952 ( .A(n7031), .B(n7032), .Z(n2984) );
  AND U6953 ( .A(n3011), .B(n3007), .Z(n7032) );
  OR U6954 ( .A(B[496]), .B(A[496]), .Z(n3011) );
  ANDN U6955 ( .B(n2998), .A(n3001), .Z(n7031) );
  ANDN U6956 ( .B(n2963), .A(n2940), .Z(n7030) );
  ANDN U6957 ( .B(n7033), .A(n2919), .Z(n5843) );
  AND U6958 ( .A(B[510]), .B(A[510]), .Z(n2919) );
  NAND U6959 ( .A(n7034), .B(n2921), .Z(n7033) );
  OR U6960 ( .A(A[510]), .B(B[510]), .Z(n2921) );
  NANDN U6961 ( .A(n2923), .B(n7035), .Z(n7034) );
  NAND U6962 ( .A(n7036), .B(n2926), .Z(n7035) );
  OR U6963 ( .A(B[509]), .B(A[509]), .Z(n2926) );
  NANDN U6964 ( .A(n2933), .B(n7037), .Z(n7036) );
  NANDN U6965 ( .A(n2935), .B(n7038), .Z(n7037) );
  NANDN U6966 ( .A(n2938), .B(n7039), .Z(n7038) );
  NANDN U6967 ( .A(n2940), .B(n7040), .Z(n7039) );
  NANDN U6968 ( .A(n2960), .B(n7041), .Z(n7040) );
  NAND U6969 ( .A(n2983), .B(n2963), .Z(n7041) );
  AND U6970 ( .A(n7042), .B(n7043), .Z(n2963) );
  AND U6971 ( .A(n2980), .B(n2976), .Z(n7043) );
  OR U6972 ( .A(B[500]), .B(A[500]), .Z(n2980) );
  AND U6973 ( .A(n2971), .B(n2967), .Z(n7042) );
  NANDN U6974 ( .A(n2997), .B(n7044), .Z(n2983) );
  NAND U6975 ( .A(n7045), .B(n2998), .Z(n7044) );
  OR U6976 ( .A(B[499]), .B(A[499]), .Z(n2998) );
  NANDN U6977 ( .A(n3000), .B(n7046), .Z(n7045) );
  NANDN U6978 ( .A(n3001), .B(n7047), .Z(n7046) );
  NANDN U6979 ( .A(n3004), .B(n7048), .Z(n7047) );
  NAND U6980 ( .A(n3007), .B(n3009), .Z(n7048) );
  AND U6981 ( .A(A[496]), .B(B[496]), .Z(n3009) );
  OR U6982 ( .A(B[497]), .B(A[497]), .Z(n3007) );
  AND U6983 ( .A(B[497]), .B(A[497]), .Z(n3004) );
  NOR U6984 ( .A(B[498]), .B(A[498]), .Z(n3001) );
  AND U6985 ( .A(B[498]), .B(A[498]), .Z(n3000) );
  AND U6986 ( .A(B[499]), .B(A[499]), .Z(n2997) );
  NANDN U6987 ( .A(n2966), .B(n7049), .Z(n2960) );
  NAND U6988 ( .A(n7050), .B(n2967), .Z(n7049) );
  OR U6989 ( .A(B[503]), .B(A[503]), .Z(n2967) );
  NANDN U6990 ( .A(n2969), .B(n7051), .Z(n7050) );
  NAND U6991 ( .A(n7052), .B(n2971), .Z(n7051) );
  OR U6992 ( .A(B[502]), .B(A[502]), .Z(n2971) );
  NANDN U6993 ( .A(n2973), .B(n7053), .Z(n7052) );
  NAND U6994 ( .A(n2976), .B(n2978), .Z(n7053) );
  AND U6995 ( .A(B[500]), .B(A[500]), .Z(n2978) );
  OR U6996 ( .A(B[501]), .B(A[501]), .Z(n2976) );
  AND U6997 ( .A(B[501]), .B(A[501]), .Z(n2973) );
  AND U6998 ( .A(B[502]), .B(A[502]), .Z(n2969) );
  AND U6999 ( .A(B[503]), .B(A[503]), .Z(n2966) );
  NAND U7000 ( .A(n7054), .B(n7055), .Z(n2940) );
  AND U7001 ( .A(n2958), .B(n2954), .Z(n7055) );
  OR U7002 ( .A(B[504]), .B(A[504]), .Z(n2958) );
  AND U7003 ( .A(n2949), .B(n2945), .Z(n7054) );
  NANDN U7004 ( .A(n2944), .B(n7056), .Z(n2938) );
  NAND U7005 ( .A(n7057), .B(n2945), .Z(n7056) );
  OR U7006 ( .A(B[507]), .B(A[507]), .Z(n2945) );
  NANDN U7007 ( .A(n2947), .B(n7058), .Z(n7057) );
  NAND U7008 ( .A(n7059), .B(n2949), .Z(n7058) );
  OR U7009 ( .A(B[506]), .B(A[506]), .Z(n2949) );
  NANDN U7010 ( .A(n2951), .B(n7060), .Z(n7059) );
  NAND U7011 ( .A(n2954), .B(n2956), .Z(n7060) );
  AND U7012 ( .A(B[504]), .B(A[504]), .Z(n2956) );
  OR U7013 ( .A(B[505]), .B(A[505]), .Z(n2954) );
  AND U7014 ( .A(B[505]), .B(A[505]), .Z(n2951) );
  AND U7015 ( .A(B[506]), .B(A[506]), .Z(n2947) );
  AND U7016 ( .A(B[507]), .B(A[507]), .Z(n2944) );
  NOR U7017 ( .A(B[508]), .B(A[508]), .Z(n2935) );
  AND U7018 ( .A(B[508]), .B(A[508]), .Z(n2933) );
  AND U7019 ( .A(B[509]), .B(A[509]), .Z(n2923) );
  NOR U7020 ( .A(B[511]), .B(A[511]), .Z(n2916) );
  NOR U7021 ( .A(n2820), .B(n5733), .Z(n5816) );
  NAND U7022 ( .A(n7061), .B(n7062), .Z(n5733) );
  AND U7023 ( .A(n7063), .B(n7064), .Z(n7062) );
  AND U7024 ( .A(n2549), .B(n2544), .Z(n7064) );
  OR U7025 ( .A(A[573]), .B(B[573]), .Z(n2544) );
  OR U7026 ( .A(A[572]), .B(B[572]), .Z(n2549) );
  AND U7027 ( .A(n2539), .B(n2535), .Z(n7063) );
  OR U7028 ( .A(B[575]), .B(A[575]), .Z(n2535) );
  OR U7029 ( .A(A[574]), .B(B[574]), .Z(n2539) );
  ANDN U7030 ( .B(n7065), .A(n2580), .Z(n7061) );
  NAND U7031 ( .A(n7066), .B(n7067), .Z(n2580) );
  AND U7032 ( .A(n2598), .B(n2594), .Z(n7067) );
  OR U7033 ( .A(A[565]), .B(B[565]), .Z(n2594) );
  OR U7034 ( .A(A[564]), .B(B[564]), .Z(n2598) );
  AND U7035 ( .A(n2589), .B(n2585), .Z(n7066) );
  OR U7036 ( .A(B[567]), .B(A[567]), .Z(n2585) );
  OR U7037 ( .A(A[566]), .B(B[566]), .Z(n2589) );
  NOR U7038 ( .A(n2602), .B(n2553), .Z(n7065) );
  NAND U7039 ( .A(n7068), .B(n7069), .Z(n2553) );
  AND U7040 ( .A(n2576), .B(n2567), .Z(n7069) );
  OR U7041 ( .A(A[569]), .B(B[569]), .Z(n2567) );
  OR U7042 ( .A(A[568]), .B(B[568]), .Z(n2576) );
  AND U7043 ( .A(n2562), .B(n2558), .Z(n7068) );
  OR U7044 ( .A(B[571]), .B(A[571]), .Z(n2558) );
  OR U7045 ( .A(A[570]), .B(B[570]), .Z(n2562) );
  NAND U7046 ( .A(n7070), .B(n7071), .Z(n2602) );
  AND U7047 ( .A(n2620), .B(n2616), .Z(n7071) );
  OR U7048 ( .A(A[561]), .B(B[561]), .Z(n2616) );
  OR U7049 ( .A(A[560]), .B(B[560]), .Z(n2620) );
  AND U7050 ( .A(n2611), .B(n2607), .Z(n7070) );
  OR U7051 ( .A(B[563]), .B(A[563]), .Z(n2607) );
  OR U7052 ( .A(A[562]), .B(B[562]), .Z(n2611) );
  NAND U7053 ( .A(n7072), .B(n7073), .Z(n2820) );
  AND U7054 ( .A(n7074), .B(n7075), .Z(n7073) );
  AND U7055 ( .A(n2839), .B(n2834), .Z(n7075) );
  OR U7056 ( .A(A[525]), .B(B[525]), .Z(n2834) );
  OR U7057 ( .A(A[524]), .B(B[524]), .Z(n2839) );
  AND U7058 ( .A(n2829), .B(n2825), .Z(n7074) );
  OR U7059 ( .A(B[527]), .B(A[527]), .Z(n2825) );
  OR U7060 ( .A(A[526]), .B(B[526]), .Z(n2829) );
  ANDN U7061 ( .B(n7076), .A(n2895), .Z(n7072) );
  NAND U7062 ( .A(n7077), .B(n7078), .Z(n2895) );
  AND U7063 ( .A(n2912), .B(n2908), .Z(n7078) );
  OR U7064 ( .A(A[513]), .B(B[513]), .Z(n2908) );
  OR U7065 ( .A(A[512]), .B(B[512]), .Z(n2912) );
  AND U7066 ( .A(n2903), .B(n2899), .Z(n7077) );
  OR U7067 ( .A(B[515]), .B(A[515]), .Z(n2899) );
  OR U7068 ( .A(A[514]), .B(B[514]), .Z(n2903) );
  NOR U7069 ( .A(n2865), .B(n2843), .Z(n7076) );
  NAND U7070 ( .A(n7079), .B(n7080), .Z(n2843) );
  AND U7071 ( .A(n2861), .B(n2857), .Z(n7080) );
  OR U7072 ( .A(A[521]), .B(B[521]), .Z(n2857) );
  OR U7073 ( .A(A[520]), .B(B[520]), .Z(n2861) );
  AND U7074 ( .A(n2852), .B(n2848), .Z(n7079) );
  OR U7075 ( .A(B[523]), .B(A[523]), .Z(n2848) );
  OR U7076 ( .A(A[522]), .B(B[522]), .Z(n2852) );
  NAND U7077 ( .A(n7081), .B(n7082), .Z(n2865) );
  AND U7078 ( .A(n2891), .B(n2887), .Z(n7082) );
  OR U7079 ( .A(A[517]), .B(B[517]), .Z(n2887) );
  OR U7080 ( .A(A[516]), .B(B[516]), .Z(n2891) );
  AND U7081 ( .A(n2882), .B(n2878), .Z(n7081) );
  OR U7082 ( .A(B[519]), .B(A[519]), .Z(n2878) );
  OR U7083 ( .A(A[518]), .B(B[518]), .Z(n2882) );
  NAND U7084 ( .A(n7083), .B(n7084), .Z(n2136) );
  NOR U7085 ( .A(n2336), .B(n2238), .Z(n7084) );
  NOR U7086 ( .A(n2436), .B(n7085), .Z(n7083) );
  NAND U7087 ( .A(n7086), .B(n7087), .Z(n2436) );
  AND U7088 ( .A(n7088), .B(n7089), .Z(n7087) );
  AND U7089 ( .A(n2459), .B(n2449), .Z(n7089) );
  AND U7090 ( .A(n2444), .B(n2440), .Z(n7088) );
  ANDN U7091 ( .B(n7090), .A(n2507), .Z(n7086) );
  NAND U7092 ( .A(n7091), .B(n7092), .Z(n2507) );
  AND U7093 ( .A(n2528), .B(n2524), .Z(n7092) );
  OR U7094 ( .A(A[576]), .B(B[576]), .Z(n2528) );
  AND U7095 ( .A(n2519), .B(n2515), .Z(n7091) );
  NOR U7096 ( .A(n2485), .B(n2463), .Z(n7090) );
  NAND U7097 ( .A(n7093), .B(n7094), .Z(n2134) );
  NAND U7098 ( .A(n7095), .B(n2149), .Z(n7094) );
  NANDN U7099 ( .A(n2151), .B(n7096), .Z(n7095) );
  NAND U7100 ( .A(n7097), .B(n2153), .Z(n7096) );
  NANDN U7101 ( .A(n2155), .B(n7098), .Z(n7097) );
  NAND U7102 ( .A(n7099), .B(n2158), .Z(n7098) );
  NANDN U7103 ( .A(n2160), .B(n7100), .Z(n7099) );
  NAND U7104 ( .A(n7101), .B(n2163), .Z(n7100) );
  NANDN U7105 ( .A(n2165), .B(n7102), .Z(n7101) );
  NANDN U7106 ( .A(n2167), .B(n7103), .Z(n7102) );
  NANDN U7107 ( .A(n2187), .B(n7104), .Z(n7103) );
  NANDN U7108 ( .A(n2189), .B(n2215), .Z(n7104) );
  NANDN U7109 ( .A(n2220), .B(n7105), .Z(n2215) );
  NAND U7110 ( .A(n7106), .B(n2221), .Z(n7105) );
  NANDN U7111 ( .A(n2223), .B(n7107), .Z(n7106) );
  NAND U7112 ( .A(n7108), .B(n2225), .Z(n7107) );
  NANDN U7113 ( .A(n2227), .B(n7109), .Z(n7108) );
  NAND U7114 ( .A(n2230), .B(n2232), .Z(n7109) );
  AND U7115 ( .A(A[624]), .B(B[624]), .Z(n2232) );
  AND U7116 ( .A(A[625]), .B(B[625]), .Z(n2227) );
  AND U7117 ( .A(A[626]), .B(B[626]), .Z(n2223) );
  AND U7118 ( .A(B[627]), .B(A[627]), .Z(n2220) );
  NANDN U7119 ( .A(n2193), .B(n7110), .Z(n2187) );
  NAND U7120 ( .A(n7111), .B(n2194), .Z(n7110) );
  NANDN U7121 ( .A(n2196), .B(n7112), .Z(n7111) );
  NAND U7122 ( .A(n7113), .B(n2198), .Z(n7112) );
  NANDN U7123 ( .A(n2200), .B(n7114), .Z(n7113) );
  NAND U7124 ( .A(n2203), .B(n2210), .Z(n7114) );
  AND U7125 ( .A(A[628]), .B(B[628]), .Z(n2210) );
  AND U7126 ( .A(A[629]), .B(B[629]), .Z(n2200) );
  AND U7127 ( .A(A[630]), .B(B[630]), .Z(n2196) );
  AND U7128 ( .A(B[631]), .B(A[631]), .Z(n2193) );
  NANDN U7129 ( .A(n2171), .B(n7115), .Z(n2165) );
  NAND U7130 ( .A(n7116), .B(n2172), .Z(n7115) );
  NANDN U7131 ( .A(n2174), .B(n7117), .Z(n7116) );
  NAND U7132 ( .A(n7118), .B(n2176), .Z(n7117) );
  NANDN U7133 ( .A(n2178), .B(n7119), .Z(n7118) );
  NAND U7134 ( .A(n2181), .B(n2183), .Z(n7119) );
  AND U7135 ( .A(A[632]), .B(B[632]), .Z(n2183) );
  AND U7136 ( .A(A[633]), .B(B[633]), .Z(n2178) );
  AND U7137 ( .A(A[634]), .B(B[634]), .Z(n2174) );
  AND U7138 ( .A(B[635]), .B(A[635]), .Z(n2171) );
  AND U7139 ( .A(A[636]), .B(B[636]), .Z(n2160) );
  AND U7140 ( .A(A[637]), .B(B[637]), .Z(n2155) );
  AND U7141 ( .A(A[638]), .B(B[638]), .Z(n2151) );
  ANDN U7142 ( .B(n7120), .A(n2148), .Z(n7093) );
  AND U7143 ( .A(B[639]), .B(A[639]), .Z(n2148) );
  NANDN U7144 ( .A(n7085), .B(n7121), .Z(n7120) );
  NANDN U7145 ( .A(n2236), .B(n7122), .Z(n7121) );
  NANDN U7146 ( .A(n2238), .B(n7123), .Z(n7122) );
  NANDN U7147 ( .A(n2334), .B(n7124), .Z(n7123) );
  NANDN U7148 ( .A(n2336), .B(n2435), .Z(n7124) );
  NANDN U7149 ( .A(n2439), .B(n7125), .Z(n2435) );
  NAND U7150 ( .A(n7126), .B(n2440), .Z(n7125) );
  OR U7151 ( .A(B[591]), .B(A[591]), .Z(n2440) );
  NANDN U7152 ( .A(n2442), .B(n7127), .Z(n7126) );
  NAND U7153 ( .A(n7128), .B(n2444), .Z(n7127) );
  OR U7154 ( .A(A[590]), .B(B[590]), .Z(n2444) );
  NANDN U7155 ( .A(n2446), .B(n7129), .Z(n7128) );
  NAND U7156 ( .A(n7130), .B(n2449), .Z(n7129) );
  OR U7157 ( .A(A[589]), .B(B[589]), .Z(n2449) );
  NANDN U7158 ( .A(n2456), .B(n7131), .Z(n7130) );
  NAND U7159 ( .A(n7132), .B(n2459), .Z(n7131) );
  OR U7160 ( .A(A[588]), .B(B[588]), .Z(n2459) );
  NANDN U7161 ( .A(n2461), .B(n7133), .Z(n7132) );
  NANDN U7162 ( .A(n2463), .B(n7134), .Z(n7133) );
  NANDN U7163 ( .A(n2483), .B(n7135), .Z(n7134) );
  NANDN U7164 ( .A(n2485), .B(n2506), .Z(n7135) );
  NANDN U7165 ( .A(n2514), .B(n7136), .Z(n2506) );
  NAND U7166 ( .A(n7137), .B(n2515), .Z(n7136) );
  OR U7167 ( .A(B[579]), .B(A[579]), .Z(n2515) );
  NANDN U7168 ( .A(n2517), .B(n7138), .Z(n7137) );
  NAND U7169 ( .A(n7139), .B(n2519), .Z(n7138) );
  OR U7170 ( .A(A[578]), .B(B[578]), .Z(n2519) );
  NANDN U7171 ( .A(n2521), .B(n7140), .Z(n7139) );
  NAND U7172 ( .A(n2524), .B(n2526), .Z(n7140) );
  AND U7173 ( .A(A[576]), .B(B[576]), .Z(n2526) );
  OR U7174 ( .A(A[577]), .B(B[577]), .Z(n2524) );
  AND U7175 ( .A(A[577]), .B(B[577]), .Z(n2521) );
  AND U7176 ( .A(A[578]), .B(B[578]), .Z(n2517) );
  AND U7177 ( .A(B[579]), .B(A[579]), .Z(n2514) );
  NAND U7178 ( .A(n7141), .B(n7142), .Z(n2485) );
  AND U7179 ( .A(n2503), .B(n2499), .Z(n7142) );
  OR U7180 ( .A(A[580]), .B(B[580]), .Z(n2503) );
  AND U7181 ( .A(n2494), .B(n2490), .Z(n7141) );
  NANDN U7182 ( .A(n2489), .B(n7143), .Z(n2483) );
  NAND U7183 ( .A(n7144), .B(n2490), .Z(n7143) );
  OR U7184 ( .A(B[583]), .B(A[583]), .Z(n2490) );
  NANDN U7185 ( .A(n2492), .B(n7145), .Z(n7144) );
  NAND U7186 ( .A(n7146), .B(n2494), .Z(n7145) );
  OR U7187 ( .A(A[582]), .B(B[582]), .Z(n2494) );
  NANDN U7188 ( .A(n2496), .B(n7147), .Z(n7146) );
  NAND U7189 ( .A(n2499), .B(n2501), .Z(n7147) );
  AND U7190 ( .A(A[580]), .B(B[580]), .Z(n2501) );
  OR U7191 ( .A(A[581]), .B(B[581]), .Z(n2499) );
  AND U7192 ( .A(A[581]), .B(B[581]), .Z(n2496) );
  AND U7193 ( .A(A[582]), .B(B[582]), .Z(n2492) );
  AND U7194 ( .A(B[583]), .B(A[583]), .Z(n2489) );
  NAND U7195 ( .A(n7148), .B(n7149), .Z(n2463) );
  AND U7196 ( .A(n2481), .B(n2477), .Z(n7149) );
  OR U7197 ( .A(A[584]), .B(B[584]), .Z(n2481) );
  AND U7198 ( .A(n2472), .B(n2468), .Z(n7148) );
  NANDN U7199 ( .A(n2467), .B(n7150), .Z(n2461) );
  NAND U7200 ( .A(n7151), .B(n2468), .Z(n7150) );
  OR U7201 ( .A(B[587]), .B(A[587]), .Z(n2468) );
  NANDN U7202 ( .A(n2470), .B(n7152), .Z(n7151) );
  NAND U7203 ( .A(n7153), .B(n2472), .Z(n7152) );
  OR U7204 ( .A(A[586]), .B(B[586]), .Z(n2472) );
  NANDN U7205 ( .A(n2474), .B(n7154), .Z(n7153) );
  NAND U7206 ( .A(n2477), .B(n2479), .Z(n7154) );
  AND U7207 ( .A(A[584]), .B(B[584]), .Z(n2479) );
  OR U7208 ( .A(A[585]), .B(B[585]), .Z(n2477) );
  AND U7209 ( .A(A[585]), .B(B[585]), .Z(n2474) );
  AND U7210 ( .A(A[586]), .B(B[586]), .Z(n2470) );
  AND U7211 ( .A(B[587]), .B(A[587]), .Z(n2467) );
  AND U7212 ( .A(A[588]), .B(B[588]), .Z(n2456) );
  AND U7213 ( .A(A[589]), .B(B[589]), .Z(n2446) );
  AND U7214 ( .A(A[590]), .B(B[590]), .Z(n2442) );
  AND U7215 ( .A(B[591]), .B(A[591]), .Z(n2439) );
  NAND U7216 ( .A(n7155), .B(n7156), .Z(n2336) );
  AND U7217 ( .A(n7157), .B(n7158), .Z(n7156) );
  AND U7218 ( .A(n2355), .B(n2350), .Z(n7158) );
  AND U7219 ( .A(n2345), .B(n2341), .Z(n7157) );
  ANDN U7220 ( .B(n7159), .A(n2415), .Z(n7155) );
  NAND U7221 ( .A(n7160), .B(n7161), .Z(n2415) );
  AND U7222 ( .A(n2432), .B(n2428), .Z(n7161) );
  OR U7223 ( .A(A[592]), .B(B[592]), .Z(n2432) );
  AND U7224 ( .A(n2423), .B(n2419), .Z(n7160) );
  NOR U7225 ( .A(n2381), .B(n2359), .Z(n7159) );
  NANDN U7226 ( .A(n2340), .B(n7162), .Z(n2334) );
  NAND U7227 ( .A(n7163), .B(n2341), .Z(n7162) );
  OR U7228 ( .A(B[607]), .B(A[607]), .Z(n2341) );
  NANDN U7229 ( .A(n2343), .B(n7164), .Z(n7163) );
  NAND U7230 ( .A(n7165), .B(n2345), .Z(n7164) );
  OR U7231 ( .A(A[606]), .B(B[606]), .Z(n2345) );
  NANDN U7232 ( .A(n2347), .B(n7166), .Z(n7165) );
  NAND U7233 ( .A(n7167), .B(n2350), .Z(n7166) );
  OR U7234 ( .A(A[605]), .B(B[605]), .Z(n2350) );
  NANDN U7235 ( .A(n2352), .B(n7168), .Z(n7167) );
  NAND U7236 ( .A(n7169), .B(n2355), .Z(n7168) );
  OR U7237 ( .A(A[604]), .B(B[604]), .Z(n2355) );
  NANDN U7238 ( .A(n2357), .B(n7170), .Z(n7169) );
  NANDN U7239 ( .A(n2359), .B(n7171), .Z(n7170) );
  NANDN U7240 ( .A(n2379), .B(n7172), .Z(n7171) );
  NANDN U7241 ( .A(n2381), .B(n2414), .Z(n7172) );
  NANDN U7242 ( .A(n2418), .B(n7173), .Z(n2414) );
  NAND U7243 ( .A(n7174), .B(n2419), .Z(n7173) );
  OR U7244 ( .A(B[595]), .B(A[595]), .Z(n2419) );
  NANDN U7245 ( .A(n2421), .B(n7175), .Z(n7174) );
  NAND U7246 ( .A(n7176), .B(n2423), .Z(n7175) );
  OR U7247 ( .A(A[594]), .B(B[594]), .Z(n2423) );
  NANDN U7248 ( .A(n2425), .B(n7177), .Z(n7176) );
  NAND U7249 ( .A(n2428), .B(n2430), .Z(n7177) );
  AND U7250 ( .A(A[592]), .B(B[592]), .Z(n2430) );
  OR U7251 ( .A(A[593]), .B(B[593]), .Z(n2428) );
  AND U7252 ( .A(A[593]), .B(B[593]), .Z(n2425) );
  AND U7253 ( .A(A[594]), .B(B[594]), .Z(n2421) );
  AND U7254 ( .A(B[595]), .B(A[595]), .Z(n2418) );
  NAND U7255 ( .A(n7178), .B(n7179), .Z(n2381) );
  AND U7256 ( .A(n2411), .B(n2407), .Z(n7179) );
  OR U7257 ( .A(A[596]), .B(B[596]), .Z(n2411) );
  AND U7258 ( .A(n2402), .B(n2398), .Z(n7178) );
  NANDN U7259 ( .A(n2397), .B(n7180), .Z(n2379) );
  NAND U7260 ( .A(n7181), .B(n2398), .Z(n7180) );
  OR U7261 ( .A(B[599]), .B(A[599]), .Z(n2398) );
  NANDN U7262 ( .A(n2400), .B(n7182), .Z(n7181) );
  NAND U7263 ( .A(n7183), .B(n2402), .Z(n7182) );
  OR U7264 ( .A(A[598]), .B(B[598]), .Z(n2402) );
  NANDN U7265 ( .A(n2404), .B(n7184), .Z(n7183) );
  NAND U7266 ( .A(n2407), .B(n2409), .Z(n7184) );
  AND U7267 ( .A(A[596]), .B(B[596]), .Z(n2409) );
  OR U7268 ( .A(A[597]), .B(B[597]), .Z(n2407) );
  AND U7269 ( .A(A[597]), .B(B[597]), .Z(n2404) );
  AND U7270 ( .A(A[598]), .B(B[598]), .Z(n2400) );
  AND U7271 ( .A(B[599]), .B(A[599]), .Z(n2397) );
  NAND U7272 ( .A(n7185), .B(n7186), .Z(n2359) );
  AND U7273 ( .A(n2377), .B(n2373), .Z(n7186) );
  OR U7274 ( .A(A[600]), .B(B[600]), .Z(n2377) );
  AND U7275 ( .A(n2368), .B(n2364), .Z(n7185) );
  NANDN U7276 ( .A(n2363), .B(n7187), .Z(n2357) );
  NAND U7277 ( .A(n7188), .B(n2364), .Z(n7187) );
  OR U7278 ( .A(B[603]), .B(A[603]), .Z(n2364) );
  NANDN U7279 ( .A(n2366), .B(n7189), .Z(n7188) );
  NAND U7280 ( .A(n7190), .B(n2368), .Z(n7189) );
  OR U7281 ( .A(A[602]), .B(B[602]), .Z(n2368) );
  NANDN U7282 ( .A(n2370), .B(n7191), .Z(n7190) );
  NAND U7283 ( .A(n2373), .B(n2375), .Z(n7191) );
  AND U7284 ( .A(A[600]), .B(B[600]), .Z(n2375) );
  OR U7285 ( .A(A[601]), .B(B[601]), .Z(n2373) );
  AND U7286 ( .A(A[601]), .B(B[601]), .Z(n2370) );
  AND U7287 ( .A(A[602]), .B(B[602]), .Z(n2366) );
  AND U7288 ( .A(B[603]), .B(A[603]), .Z(n2363) );
  AND U7289 ( .A(A[604]), .B(B[604]), .Z(n2352) );
  AND U7290 ( .A(A[605]), .B(B[605]), .Z(n2347) );
  AND U7291 ( .A(A[606]), .B(B[606]), .Z(n2343) );
  AND U7292 ( .A(B[607]), .B(A[607]), .Z(n2340) );
  NAND U7293 ( .A(n7192), .B(n7193), .Z(n2238) );
  AND U7294 ( .A(n7194), .B(n7195), .Z(n7193) );
  AND U7295 ( .A(n2257), .B(n2252), .Z(n7195) );
  AND U7296 ( .A(n2247), .B(n2243), .Z(n7194) );
  ANDN U7297 ( .B(n7196), .A(n2310), .Z(n7192) );
  NAND U7298 ( .A(n7197), .B(n7198), .Z(n2310) );
  AND U7299 ( .A(n2332), .B(n2323), .Z(n7198) );
  OR U7300 ( .A(A[608]), .B(B[608]), .Z(n2332) );
  AND U7301 ( .A(n2318), .B(n2314), .Z(n7197) );
  NOR U7302 ( .A(n2288), .B(n2261), .Z(n7196) );
  NANDN U7303 ( .A(n2242), .B(n7199), .Z(n2236) );
  NAND U7304 ( .A(n7200), .B(n2243), .Z(n7199) );
  OR U7305 ( .A(B[623]), .B(A[623]), .Z(n2243) );
  NANDN U7306 ( .A(n2245), .B(n7201), .Z(n7200) );
  NAND U7307 ( .A(n7202), .B(n2247), .Z(n7201) );
  OR U7308 ( .A(A[622]), .B(B[622]), .Z(n2247) );
  NANDN U7309 ( .A(n2249), .B(n7203), .Z(n7202) );
  NAND U7310 ( .A(n7204), .B(n2252), .Z(n7203) );
  OR U7311 ( .A(A[621]), .B(B[621]), .Z(n2252) );
  NANDN U7312 ( .A(n2254), .B(n7205), .Z(n7204) );
  NAND U7313 ( .A(n7206), .B(n2257), .Z(n7205) );
  OR U7314 ( .A(A[620]), .B(B[620]), .Z(n2257) );
  NANDN U7315 ( .A(n2259), .B(n7207), .Z(n7206) );
  NANDN U7316 ( .A(n2261), .B(n7208), .Z(n7207) );
  NANDN U7317 ( .A(n2286), .B(n7209), .Z(n7208) );
  NANDN U7318 ( .A(n2288), .B(n2309), .Z(n7209) );
  NANDN U7319 ( .A(n2313), .B(n7210), .Z(n2309) );
  NAND U7320 ( .A(n7211), .B(n2314), .Z(n7210) );
  OR U7321 ( .A(B[611]), .B(A[611]), .Z(n2314) );
  NANDN U7322 ( .A(n2316), .B(n7212), .Z(n7211) );
  NAND U7323 ( .A(n7213), .B(n2318), .Z(n7212) );
  OR U7324 ( .A(A[610]), .B(B[610]), .Z(n2318) );
  NANDN U7325 ( .A(n2320), .B(n7214), .Z(n7213) );
  NAND U7326 ( .A(n2323), .B(n2330), .Z(n7214) );
  AND U7327 ( .A(A[608]), .B(B[608]), .Z(n2330) );
  OR U7328 ( .A(A[609]), .B(B[609]), .Z(n2323) );
  AND U7329 ( .A(A[609]), .B(B[609]), .Z(n2320) );
  AND U7330 ( .A(A[610]), .B(B[610]), .Z(n2316) );
  AND U7331 ( .A(B[611]), .B(A[611]), .Z(n2313) );
  NAND U7332 ( .A(n7215), .B(n7216), .Z(n2288) );
  AND U7333 ( .A(n2306), .B(n2302), .Z(n7216) );
  OR U7334 ( .A(A[612]), .B(B[612]), .Z(n2306) );
  AND U7335 ( .A(n2297), .B(n2293), .Z(n7215) );
  NANDN U7336 ( .A(n2292), .B(n7217), .Z(n2286) );
  NAND U7337 ( .A(n7218), .B(n2293), .Z(n7217) );
  OR U7338 ( .A(B[615]), .B(A[615]), .Z(n2293) );
  NANDN U7339 ( .A(n2295), .B(n7219), .Z(n7218) );
  NAND U7340 ( .A(n7220), .B(n2297), .Z(n7219) );
  OR U7341 ( .A(A[614]), .B(B[614]), .Z(n2297) );
  NANDN U7342 ( .A(n2299), .B(n7221), .Z(n7220) );
  NAND U7343 ( .A(n2302), .B(n2304), .Z(n7221) );
  AND U7344 ( .A(A[612]), .B(B[612]), .Z(n2304) );
  OR U7345 ( .A(A[613]), .B(B[613]), .Z(n2302) );
  AND U7346 ( .A(A[613]), .B(B[613]), .Z(n2299) );
  AND U7347 ( .A(A[614]), .B(B[614]), .Z(n2295) );
  AND U7348 ( .A(B[615]), .B(A[615]), .Z(n2292) );
  NAND U7349 ( .A(n7222), .B(n7223), .Z(n2261) );
  AND U7350 ( .A(n2284), .B(n2280), .Z(n7223) );
  OR U7351 ( .A(A[616]), .B(B[616]), .Z(n2284) );
  AND U7352 ( .A(n2275), .B(n2271), .Z(n7222) );
  NANDN U7353 ( .A(n2270), .B(n7224), .Z(n2259) );
  NAND U7354 ( .A(n7225), .B(n2271), .Z(n7224) );
  OR U7355 ( .A(B[619]), .B(A[619]), .Z(n2271) );
  NANDN U7356 ( .A(n2273), .B(n7226), .Z(n7225) );
  NAND U7357 ( .A(n7227), .B(n2275), .Z(n7226) );
  OR U7358 ( .A(A[618]), .B(B[618]), .Z(n2275) );
  NANDN U7359 ( .A(n2277), .B(n7228), .Z(n7227) );
  NAND U7360 ( .A(n2280), .B(n2282), .Z(n7228) );
  AND U7361 ( .A(A[616]), .B(B[616]), .Z(n2282) );
  OR U7362 ( .A(A[617]), .B(B[617]), .Z(n2280) );
  AND U7363 ( .A(A[617]), .B(B[617]), .Z(n2277) );
  AND U7364 ( .A(A[618]), .B(B[618]), .Z(n2273) );
  AND U7365 ( .A(B[619]), .B(A[619]), .Z(n2270) );
  AND U7366 ( .A(A[620]), .B(B[620]), .Z(n2254) );
  AND U7367 ( .A(A[621]), .B(B[621]), .Z(n2249) );
  AND U7368 ( .A(A[622]), .B(B[622]), .Z(n2245) );
  AND U7369 ( .A(B[623]), .B(A[623]), .Z(n2242) );
  NAND U7370 ( .A(n7229), .B(n7230), .Z(n7085) );
  AND U7371 ( .A(n7231), .B(n7232), .Z(n7230) );
  AND U7372 ( .A(n2163), .B(n2158), .Z(n7232) );
  OR U7373 ( .A(A[637]), .B(B[637]), .Z(n2158) );
  OR U7374 ( .A(A[636]), .B(B[636]), .Z(n2163) );
  AND U7375 ( .A(n2153), .B(n2149), .Z(n7231) );
  OR U7376 ( .A(B[639]), .B(A[639]), .Z(n2149) );
  OR U7377 ( .A(A[638]), .B(B[638]), .Z(n2153) );
  ANDN U7378 ( .B(n7233), .A(n2189), .Z(n7229) );
  NAND U7379 ( .A(n7234), .B(n7235), .Z(n2189) );
  AND U7380 ( .A(n2212), .B(n2203), .Z(n7235) );
  OR U7381 ( .A(A[629]), .B(B[629]), .Z(n2203) );
  OR U7382 ( .A(A[628]), .B(B[628]), .Z(n2212) );
  AND U7383 ( .A(n2198), .B(n2194), .Z(n7234) );
  OR U7384 ( .A(B[631]), .B(A[631]), .Z(n2194) );
  OR U7385 ( .A(A[630]), .B(B[630]), .Z(n2198) );
  NOR U7386 ( .A(n2216), .B(n2167), .Z(n7233) );
  NAND U7387 ( .A(n7236), .B(n7237), .Z(n2167) );
  AND U7388 ( .A(n2185), .B(n2181), .Z(n7237) );
  OR U7389 ( .A(A[633]), .B(B[633]), .Z(n2181) );
  OR U7390 ( .A(A[632]), .B(B[632]), .Z(n2185) );
  AND U7391 ( .A(n2176), .B(n2172), .Z(n7236) );
  OR U7392 ( .A(B[635]), .B(A[635]), .Z(n2172) );
  OR U7393 ( .A(A[634]), .B(B[634]), .Z(n2176) );
  NAND U7394 ( .A(n7238), .B(n7239), .Z(n2216) );
  AND U7395 ( .A(n2234), .B(n2230), .Z(n7239) );
  OR U7396 ( .A(A[625]), .B(B[625]), .Z(n2230) );
  OR U7397 ( .A(A[624]), .B(B[624]), .Z(n2234) );
  AND U7398 ( .A(n2225), .B(n2221), .Z(n7238) );
  OR U7399 ( .A(B[627]), .B(A[627]), .Z(n2221) );
  OR U7400 ( .A(A[626]), .B(B[626]), .Z(n2225) );
  NAND U7401 ( .A(n7240), .B(n7241), .Z(n1754) );
  ANDN U7402 ( .B(n1855), .A(n1951), .Z(n7241) );
  NOR U7403 ( .A(n2048), .B(n7242), .Z(n7240) );
  NAND U7404 ( .A(n7243), .B(n7244), .Z(n2048) );
  AND U7405 ( .A(n7245), .B(n7246), .Z(n7244) );
  AND U7406 ( .A(n2066), .B(n2061), .Z(n7246) );
  AND U7407 ( .A(n2056), .B(n2052), .Z(n7245) );
  ANDN U7408 ( .B(n7247), .A(n2115), .Z(n7243) );
  NAND U7409 ( .A(n7248), .B(n7249), .Z(n2115) );
  AND U7410 ( .A(n2132), .B(n2128), .Z(n7249) );
  OR U7411 ( .A(B[640]), .B(A[640]), .Z(n2132) );
  AND U7412 ( .A(n2123), .B(n2119), .Z(n7248) );
  ANDN U7413 ( .B(n2070), .A(n2093), .Z(n7247) );
  NAND U7414 ( .A(n7250), .B(n7251), .Z(n1752) );
  NAND U7415 ( .A(n7252), .B(n1759), .Z(n7251) );
  NANDN U7416 ( .A(n1761), .B(n7253), .Z(n7252) );
  NAND U7417 ( .A(n7254), .B(n1763), .Z(n7253) );
  NANDN U7418 ( .A(n1765), .B(n7255), .Z(n7254) );
  NAND U7419 ( .A(n7256), .B(n1768), .Z(n7255) );
  NANDN U7420 ( .A(n1770), .B(n7257), .Z(n7256) );
  NAND U7421 ( .A(n7258), .B(n1773), .Z(n7257) );
  NANDN U7422 ( .A(n1775), .B(n7259), .Z(n7258) );
  NANDN U7423 ( .A(n1777), .B(n7260), .Z(n7259) );
  NANDN U7424 ( .A(n1804), .B(n7261), .Z(n7260) );
  NANDN U7425 ( .A(n1806), .B(n1827), .Z(n7261) );
  NANDN U7426 ( .A(n1832), .B(n7262), .Z(n1827) );
  NAND U7427 ( .A(n7263), .B(n1833), .Z(n7262) );
  NANDN U7428 ( .A(n1835), .B(n7264), .Z(n7263) );
  NAND U7429 ( .A(n7265), .B(n1837), .Z(n7264) );
  NANDN U7430 ( .A(n1839), .B(n7266), .Z(n7265) );
  NAND U7431 ( .A(n1842), .B(n1849), .Z(n7266) );
  AND U7432 ( .A(A[688]), .B(B[688]), .Z(n1849) );
  AND U7433 ( .A(A[689]), .B(B[689]), .Z(n1839) );
  AND U7434 ( .A(A[690]), .B(B[690]), .Z(n1835) );
  AND U7435 ( .A(B[691]), .B(A[691]), .Z(n1832) );
  NANDN U7436 ( .A(n1810), .B(n7267), .Z(n1804) );
  NAND U7437 ( .A(n7268), .B(n1811), .Z(n7267) );
  NANDN U7438 ( .A(n1813), .B(n7269), .Z(n7268) );
  NAND U7439 ( .A(n7270), .B(n1815), .Z(n7269) );
  NANDN U7440 ( .A(n1817), .B(n7271), .Z(n7270) );
  NAND U7441 ( .A(n1820), .B(n1822), .Z(n7271) );
  AND U7442 ( .A(A[692]), .B(B[692]), .Z(n1822) );
  AND U7443 ( .A(A[693]), .B(B[693]), .Z(n1817) );
  AND U7444 ( .A(A[694]), .B(B[694]), .Z(n1813) );
  AND U7445 ( .A(B[695]), .B(A[695]), .Z(n1810) );
  NANDN U7446 ( .A(n1788), .B(n7272), .Z(n1775) );
  NAND U7447 ( .A(n7273), .B(n1789), .Z(n7272) );
  NANDN U7448 ( .A(n1791), .B(n7274), .Z(n7273) );
  NAND U7449 ( .A(n7275), .B(n1793), .Z(n7274) );
  NANDN U7450 ( .A(n1795), .B(n7276), .Z(n7275) );
  NAND U7451 ( .A(n1798), .B(n1800), .Z(n7276) );
  AND U7452 ( .A(A[696]), .B(B[696]), .Z(n1800) );
  AND U7453 ( .A(A[697]), .B(B[697]), .Z(n1795) );
  AND U7454 ( .A(A[698]), .B(B[698]), .Z(n1791) );
  AND U7455 ( .A(B[699]), .B(A[699]), .Z(n1788) );
  AND U7456 ( .A(A[700]), .B(B[700]), .Z(n1770) );
  AND U7457 ( .A(A[701]), .B(B[701]), .Z(n1765) );
  AND U7458 ( .A(A[702]), .B(B[702]), .Z(n1761) );
  ANDN U7459 ( .B(n7277), .A(n1758), .Z(n7250) );
  AND U7460 ( .A(B[703]), .B(A[703]), .Z(n1758) );
  NANDN U7461 ( .A(n7242), .B(n7278), .Z(n7277) );
  NANDN U7462 ( .A(n1853), .B(n7279), .Z(n7278) );
  NAND U7463 ( .A(n7280), .B(n1855), .Z(n7279) );
  AND U7464 ( .A(n7281), .B(n7282), .Z(n1855) );
  AND U7465 ( .A(n7283), .B(n7284), .Z(n7282) );
  AND U7466 ( .A(n1874), .B(n1869), .Z(n7284) );
  AND U7467 ( .A(n1864), .B(n1860), .Z(n7283) );
  ANDN U7468 ( .B(n7285), .A(n1930), .Z(n7281) );
  NAND U7469 ( .A(n7286), .B(n7287), .Z(n1930) );
  AND U7470 ( .A(n1947), .B(n1943), .Z(n7287) );
  OR U7471 ( .A(B[672]), .B(A[672]), .Z(n1947) );
  AND U7472 ( .A(n1938), .B(n1934), .Z(n7286) );
  ANDN U7473 ( .B(n1878), .A(n1900), .Z(n7285) );
  NANDN U7474 ( .A(n1949), .B(n7288), .Z(n7280) );
  NANDN U7475 ( .A(n1951), .B(n2047), .Z(n7288) );
  NANDN U7476 ( .A(n2051), .B(n7289), .Z(n2047) );
  NAND U7477 ( .A(n7290), .B(n2052), .Z(n7289) );
  OR U7478 ( .A(B[655]), .B(A[655]), .Z(n2052) );
  NANDN U7479 ( .A(n2054), .B(n7291), .Z(n7290) );
  NAND U7480 ( .A(n7292), .B(n2056), .Z(n7291) );
  OR U7481 ( .A(B[654]), .B(A[654]), .Z(n2056) );
  NANDN U7482 ( .A(n2058), .B(n7293), .Z(n7292) );
  NAND U7483 ( .A(n7294), .B(n2061), .Z(n7293) );
  OR U7484 ( .A(B[653]), .B(A[653]), .Z(n2061) );
  NANDN U7485 ( .A(n2063), .B(n7295), .Z(n7294) );
  NAND U7486 ( .A(n7296), .B(n2066), .Z(n7295) );
  OR U7487 ( .A(B[652]), .B(A[652]), .Z(n2066) );
  NANDN U7488 ( .A(n2068), .B(n7297), .Z(n7296) );
  NAND U7489 ( .A(n7298), .B(n2070), .Z(n7297) );
  AND U7490 ( .A(n7299), .B(n7300), .Z(n2070) );
  AND U7491 ( .A(n2089), .B(n2084), .Z(n7300) );
  OR U7492 ( .A(B[648]), .B(A[648]), .Z(n2089) );
  AND U7493 ( .A(n2079), .B(n2075), .Z(n7299) );
  NANDN U7494 ( .A(n2091), .B(n7301), .Z(n7298) );
  NANDN U7495 ( .A(n2093), .B(n2114), .Z(n7301) );
  NANDN U7496 ( .A(n2118), .B(n7302), .Z(n2114) );
  NAND U7497 ( .A(n7303), .B(n2119), .Z(n7302) );
  OR U7498 ( .A(B[643]), .B(A[643]), .Z(n2119) );
  NANDN U7499 ( .A(n2121), .B(n7304), .Z(n7303) );
  NAND U7500 ( .A(n7305), .B(n2123), .Z(n7304) );
  OR U7501 ( .A(B[642]), .B(A[642]), .Z(n2123) );
  NANDN U7502 ( .A(n2125), .B(n7306), .Z(n7305) );
  NAND U7503 ( .A(n2128), .B(n2130), .Z(n7306) );
  AND U7504 ( .A(B[640]), .B(A[640]), .Z(n2130) );
  OR U7505 ( .A(B[641]), .B(A[641]), .Z(n2128) );
  AND U7506 ( .A(B[641]), .B(A[641]), .Z(n2125) );
  AND U7507 ( .A(B[642]), .B(A[642]), .Z(n2121) );
  AND U7508 ( .A(B[643]), .B(A[643]), .Z(n2118) );
  NAND U7509 ( .A(n7307), .B(n7308), .Z(n2093) );
  AND U7510 ( .A(n2111), .B(n2107), .Z(n7308) );
  OR U7511 ( .A(B[644]), .B(A[644]), .Z(n2111) );
  AND U7512 ( .A(n2102), .B(n2098), .Z(n7307) );
  NANDN U7513 ( .A(n2097), .B(n7309), .Z(n2091) );
  NAND U7514 ( .A(n7310), .B(n2098), .Z(n7309) );
  OR U7515 ( .A(B[647]), .B(A[647]), .Z(n2098) );
  NANDN U7516 ( .A(n2100), .B(n7311), .Z(n7310) );
  NAND U7517 ( .A(n7312), .B(n2102), .Z(n7311) );
  OR U7518 ( .A(B[646]), .B(A[646]), .Z(n2102) );
  NANDN U7519 ( .A(n2104), .B(n7313), .Z(n7312) );
  NAND U7520 ( .A(n2107), .B(n2109), .Z(n7313) );
  AND U7521 ( .A(B[644]), .B(A[644]), .Z(n2109) );
  OR U7522 ( .A(B[645]), .B(A[645]), .Z(n2107) );
  AND U7523 ( .A(B[645]), .B(A[645]), .Z(n2104) );
  AND U7524 ( .A(B[646]), .B(A[646]), .Z(n2100) );
  AND U7525 ( .A(B[647]), .B(A[647]), .Z(n2097) );
  NANDN U7526 ( .A(n2074), .B(n7314), .Z(n2068) );
  NAND U7527 ( .A(n7315), .B(n2075), .Z(n7314) );
  OR U7528 ( .A(B[651]), .B(A[651]), .Z(n2075) );
  NANDN U7529 ( .A(n2077), .B(n7316), .Z(n7315) );
  NAND U7530 ( .A(n7317), .B(n2079), .Z(n7316) );
  OR U7531 ( .A(B[650]), .B(A[650]), .Z(n2079) );
  NANDN U7532 ( .A(n2081), .B(n7318), .Z(n7317) );
  NAND U7533 ( .A(n2084), .B(n2087), .Z(n7318) );
  AND U7534 ( .A(B[648]), .B(A[648]), .Z(n2087) );
  OR U7535 ( .A(B[649]), .B(A[649]), .Z(n2084) );
  AND U7536 ( .A(B[649]), .B(A[649]), .Z(n2081) );
  AND U7537 ( .A(B[650]), .B(A[650]), .Z(n2077) );
  AND U7538 ( .A(B[651]), .B(A[651]), .Z(n2074) );
  AND U7539 ( .A(B[652]), .B(A[652]), .Z(n2063) );
  AND U7540 ( .A(B[653]), .B(A[653]), .Z(n2058) );
  AND U7541 ( .A(B[654]), .B(A[654]), .Z(n2054) );
  AND U7542 ( .A(B[655]), .B(A[655]), .Z(n2051) );
  NAND U7543 ( .A(n7319), .B(n7320), .Z(n1951) );
  AND U7544 ( .A(n7321), .B(n7322), .Z(n7320) );
  AND U7545 ( .A(n1975), .B(n1965), .Z(n7322) );
  AND U7546 ( .A(n1960), .B(n1956), .Z(n7321) );
  ANDN U7547 ( .B(n7323), .A(n2023), .Z(n7319) );
  NAND U7548 ( .A(n7324), .B(n7325), .Z(n2023) );
  AND U7549 ( .A(n2044), .B(n2040), .Z(n7325) );
  OR U7550 ( .A(B[656]), .B(A[656]), .Z(n2044) );
  AND U7551 ( .A(n2035), .B(n2031), .Z(n7324) );
  ANDN U7552 ( .B(n1979), .A(n2001), .Z(n7323) );
  NANDN U7553 ( .A(n1955), .B(n7326), .Z(n1949) );
  NAND U7554 ( .A(n7327), .B(n1956), .Z(n7326) );
  OR U7555 ( .A(B[671]), .B(A[671]), .Z(n1956) );
  NANDN U7556 ( .A(n1958), .B(n7328), .Z(n7327) );
  NAND U7557 ( .A(n7329), .B(n1960), .Z(n7328) );
  OR U7558 ( .A(B[670]), .B(A[670]), .Z(n1960) );
  NANDN U7559 ( .A(n1962), .B(n7330), .Z(n7329) );
  NAND U7560 ( .A(n7331), .B(n1965), .Z(n7330) );
  OR U7561 ( .A(B[669]), .B(A[669]), .Z(n1965) );
  NANDN U7562 ( .A(n1972), .B(n7332), .Z(n7331) );
  NAND U7563 ( .A(n7333), .B(n1975), .Z(n7332) );
  OR U7564 ( .A(B[668]), .B(A[668]), .Z(n1975) );
  NANDN U7565 ( .A(n1977), .B(n7334), .Z(n7333) );
  NAND U7566 ( .A(n7335), .B(n1979), .Z(n7334) );
  AND U7567 ( .A(n7336), .B(n7337), .Z(n1979) );
  AND U7568 ( .A(n1997), .B(n1993), .Z(n7337) );
  OR U7569 ( .A(B[664]), .B(A[664]), .Z(n1997) );
  AND U7570 ( .A(n1988), .B(n1984), .Z(n7336) );
  NANDN U7571 ( .A(n1999), .B(n7338), .Z(n7335) );
  NANDN U7572 ( .A(n2001), .B(n2022), .Z(n7338) );
  NANDN U7573 ( .A(n2030), .B(n7339), .Z(n2022) );
  NAND U7574 ( .A(n7340), .B(n2031), .Z(n7339) );
  OR U7575 ( .A(B[659]), .B(A[659]), .Z(n2031) );
  NANDN U7576 ( .A(n2033), .B(n7341), .Z(n7340) );
  NAND U7577 ( .A(n7342), .B(n2035), .Z(n7341) );
  OR U7578 ( .A(B[658]), .B(A[658]), .Z(n2035) );
  NANDN U7579 ( .A(n2037), .B(n7343), .Z(n7342) );
  NAND U7580 ( .A(n2040), .B(n2042), .Z(n7343) );
  AND U7581 ( .A(B[656]), .B(A[656]), .Z(n2042) );
  OR U7582 ( .A(B[657]), .B(A[657]), .Z(n2040) );
  AND U7583 ( .A(B[657]), .B(A[657]), .Z(n2037) );
  AND U7584 ( .A(B[658]), .B(A[658]), .Z(n2033) );
  AND U7585 ( .A(B[659]), .B(A[659]), .Z(n2030) );
  NAND U7586 ( .A(n7344), .B(n7345), .Z(n2001) );
  AND U7587 ( .A(n2019), .B(n2015), .Z(n7345) );
  OR U7588 ( .A(B[660]), .B(A[660]), .Z(n2019) );
  AND U7589 ( .A(n2010), .B(n2006), .Z(n7344) );
  NANDN U7590 ( .A(n2005), .B(n7346), .Z(n1999) );
  NAND U7591 ( .A(n7347), .B(n2006), .Z(n7346) );
  OR U7592 ( .A(B[663]), .B(A[663]), .Z(n2006) );
  NANDN U7593 ( .A(n2008), .B(n7348), .Z(n7347) );
  NAND U7594 ( .A(n7349), .B(n2010), .Z(n7348) );
  OR U7595 ( .A(B[662]), .B(A[662]), .Z(n2010) );
  NANDN U7596 ( .A(n2012), .B(n7350), .Z(n7349) );
  NAND U7597 ( .A(n2015), .B(n2017), .Z(n7350) );
  AND U7598 ( .A(B[660]), .B(A[660]), .Z(n2017) );
  OR U7599 ( .A(B[661]), .B(A[661]), .Z(n2015) );
  AND U7600 ( .A(B[661]), .B(A[661]), .Z(n2012) );
  AND U7601 ( .A(B[662]), .B(A[662]), .Z(n2008) );
  AND U7602 ( .A(B[663]), .B(A[663]), .Z(n2005) );
  NANDN U7603 ( .A(n1983), .B(n7351), .Z(n1977) );
  NAND U7604 ( .A(n7352), .B(n1984), .Z(n7351) );
  OR U7605 ( .A(B[667]), .B(A[667]), .Z(n1984) );
  NANDN U7606 ( .A(n1986), .B(n7353), .Z(n7352) );
  NAND U7607 ( .A(n7354), .B(n1988), .Z(n7353) );
  OR U7608 ( .A(B[666]), .B(A[666]), .Z(n1988) );
  NANDN U7609 ( .A(n1990), .B(n7355), .Z(n7354) );
  NAND U7610 ( .A(n1993), .B(n1995), .Z(n7355) );
  AND U7611 ( .A(B[664]), .B(A[664]), .Z(n1995) );
  OR U7612 ( .A(B[665]), .B(A[665]), .Z(n1993) );
  AND U7613 ( .A(B[665]), .B(A[665]), .Z(n1990) );
  AND U7614 ( .A(B[666]), .B(A[666]), .Z(n1986) );
  AND U7615 ( .A(B[667]), .B(A[667]), .Z(n1983) );
  AND U7616 ( .A(B[668]), .B(A[668]), .Z(n1972) );
  AND U7617 ( .A(B[669]), .B(A[669]), .Z(n1962) );
  AND U7618 ( .A(B[670]), .B(A[670]), .Z(n1958) );
  AND U7619 ( .A(B[671]), .B(A[671]), .Z(n1955) );
  NANDN U7620 ( .A(n1859), .B(n7356), .Z(n1853) );
  NAND U7621 ( .A(n7357), .B(n1860), .Z(n7356) );
  OR U7622 ( .A(B[687]), .B(A[687]), .Z(n1860) );
  NANDN U7623 ( .A(n1862), .B(n7358), .Z(n7357) );
  NAND U7624 ( .A(n7359), .B(n1864), .Z(n7358) );
  OR U7625 ( .A(B[686]), .B(A[686]), .Z(n1864) );
  NANDN U7626 ( .A(n1866), .B(n7360), .Z(n7359) );
  NAND U7627 ( .A(n7361), .B(n1869), .Z(n7360) );
  OR U7628 ( .A(B[685]), .B(A[685]), .Z(n1869) );
  NANDN U7629 ( .A(n1871), .B(n7362), .Z(n7361) );
  NAND U7630 ( .A(n7363), .B(n1874), .Z(n7362) );
  OR U7631 ( .A(B[684]), .B(A[684]), .Z(n1874) );
  NANDN U7632 ( .A(n1876), .B(n7364), .Z(n7363) );
  NAND U7633 ( .A(n7365), .B(n1878), .Z(n7364) );
  AND U7634 ( .A(n7366), .B(n7367), .Z(n1878) );
  AND U7635 ( .A(n1896), .B(n1892), .Z(n7367) );
  OR U7636 ( .A(B[680]), .B(A[680]), .Z(n1896) );
  AND U7637 ( .A(n1887), .B(n1883), .Z(n7366) );
  NANDN U7638 ( .A(n1898), .B(n7368), .Z(n7365) );
  NANDN U7639 ( .A(n1900), .B(n1929), .Z(n7368) );
  NANDN U7640 ( .A(n1933), .B(n7369), .Z(n1929) );
  NAND U7641 ( .A(n7370), .B(n1934), .Z(n7369) );
  OR U7642 ( .A(B[675]), .B(A[675]), .Z(n1934) );
  NANDN U7643 ( .A(n1936), .B(n7371), .Z(n7370) );
  NAND U7644 ( .A(n7372), .B(n1938), .Z(n7371) );
  OR U7645 ( .A(B[674]), .B(A[674]), .Z(n1938) );
  NANDN U7646 ( .A(n1940), .B(n7373), .Z(n7372) );
  NAND U7647 ( .A(n1943), .B(n1945), .Z(n7373) );
  AND U7648 ( .A(B[672]), .B(A[672]), .Z(n1945) );
  OR U7649 ( .A(B[673]), .B(A[673]), .Z(n1943) );
  AND U7650 ( .A(B[673]), .B(A[673]), .Z(n1940) );
  AND U7651 ( .A(B[674]), .B(A[674]), .Z(n1936) );
  AND U7652 ( .A(B[675]), .B(A[675]), .Z(n1933) );
  NAND U7653 ( .A(n7374), .B(n7375), .Z(n1900) );
  AND U7654 ( .A(n1926), .B(n1922), .Z(n7375) );
  OR U7655 ( .A(B[676]), .B(A[676]), .Z(n1926) );
  AND U7656 ( .A(n1917), .B(n1913), .Z(n7374) );
  NANDN U7657 ( .A(n1912), .B(n7376), .Z(n1898) );
  NAND U7658 ( .A(n7377), .B(n1913), .Z(n7376) );
  OR U7659 ( .A(B[679]), .B(A[679]), .Z(n1913) );
  NANDN U7660 ( .A(n1915), .B(n7378), .Z(n7377) );
  NAND U7661 ( .A(n7379), .B(n1917), .Z(n7378) );
  OR U7662 ( .A(B[678]), .B(A[678]), .Z(n1917) );
  NANDN U7663 ( .A(n1919), .B(n7380), .Z(n7379) );
  NAND U7664 ( .A(n1922), .B(n1924), .Z(n7380) );
  AND U7665 ( .A(B[676]), .B(A[676]), .Z(n1924) );
  OR U7666 ( .A(B[677]), .B(A[677]), .Z(n1922) );
  AND U7667 ( .A(B[677]), .B(A[677]), .Z(n1919) );
  AND U7668 ( .A(B[678]), .B(A[678]), .Z(n1915) );
  AND U7669 ( .A(B[679]), .B(A[679]), .Z(n1912) );
  NANDN U7670 ( .A(n1882), .B(n7381), .Z(n1876) );
  NAND U7671 ( .A(n7382), .B(n1883), .Z(n7381) );
  OR U7672 ( .A(B[683]), .B(A[683]), .Z(n1883) );
  NANDN U7673 ( .A(n1885), .B(n7383), .Z(n7382) );
  NAND U7674 ( .A(n7384), .B(n1887), .Z(n7383) );
  OR U7675 ( .A(B[682]), .B(A[682]), .Z(n1887) );
  NANDN U7676 ( .A(n1889), .B(n7385), .Z(n7384) );
  NAND U7677 ( .A(n1892), .B(n1894), .Z(n7385) );
  AND U7678 ( .A(B[680]), .B(A[680]), .Z(n1894) );
  OR U7679 ( .A(B[681]), .B(A[681]), .Z(n1892) );
  AND U7680 ( .A(B[681]), .B(A[681]), .Z(n1889) );
  AND U7681 ( .A(B[682]), .B(A[682]), .Z(n1885) );
  AND U7682 ( .A(B[683]), .B(A[683]), .Z(n1882) );
  AND U7683 ( .A(B[684]), .B(A[684]), .Z(n1871) );
  AND U7684 ( .A(B[685]), .B(A[685]), .Z(n1866) );
  AND U7685 ( .A(B[686]), .B(A[686]), .Z(n1862) );
  AND U7686 ( .A(B[687]), .B(A[687]), .Z(n1859) );
  NAND U7687 ( .A(n7386), .B(n7387), .Z(n7242) );
  AND U7688 ( .A(n7388), .B(n7389), .Z(n7387) );
  AND U7689 ( .A(n1773), .B(n1768), .Z(n7389) );
  OR U7690 ( .A(A[701]), .B(B[701]), .Z(n1768) );
  OR U7691 ( .A(A[700]), .B(B[700]), .Z(n1773) );
  AND U7692 ( .A(n1763), .B(n1759), .Z(n7388) );
  OR U7693 ( .A(B[703]), .B(A[703]), .Z(n1759) );
  OR U7694 ( .A(A[702]), .B(B[702]), .Z(n1763) );
  ANDN U7695 ( .B(n7390), .A(n1806), .Z(n7386) );
  NAND U7696 ( .A(n7391), .B(n7392), .Z(n1806) );
  AND U7697 ( .A(n1824), .B(n1820), .Z(n7392) );
  OR U7698 ( .A(A[693]), .B(B[693]), .Z(n1820) );
  OR U7699 ( .A(A[692]), .B(B[692]), .Z(n1824) );
  AND U7700 ( .A(n1815), .B(n1811), .Z(n7391) );
  OR U7701 ( .A(B[695]), .B(A[695]), .Z(n1811) );
  OR U7702 ( .A(A[694]), .B(B[694]), .Z(n1815) );
  NOR U7703 ( .A(n1828), .B(n1777), .Z(n7390) );
  NAND U7704 ( .A(n7393), .B(n7394), .Z(n1777) );
  AND U7705 ( .A(n1802), .B(n1798), .Z(n7394) );
  OR U7706 ( .A(A[697]), .B(B[697]), .Z(n1798) );
  OR U7707 ( .A(A[696]), .B(B[696]), .Z(n1802) );
  AND U7708 ( .A(n1793), .B(n1789), .Z(n7393) );
  OR U7709 ( .A(B[699]), .B(A[699]), .Z(n1789) );
  OR U7710 ( .A(A[698]), .B(B[698]), .Z(n1793) );
  NAND U7711 ( .A(n7395), .B(n7396), .Z(n1828) );
  AND U7712 ( .A(n1851), .B(n1842), .Z(n7396) );
  OR U7713 ( .A(A[689]), .B(B[689]), .Z(n1842) );
  OR U7714 ( .A(A[688]), .B(B[688]), .Z(n1851) );
  AND U7715 ( .A(n1837), .B(n1833), .Z(n7395) );
  OR U7716 ( .A(B[691]), .B(A[691]), .Z(n1833) );
  OR U7717 ( .A(A[690]), .B(B[690]), .Z(n1837) );
  NAND U7718 ( .A(n7397), .B(n7398), .Z(n1653) );
  AND U7719 ( .A(n7399), .B(n7400), .Z(n7398) );
  AND U7720 ( .A(n1680), .B(n1675), .Z(n7400) );
  AND U7721 ( .A(n1670), .B(n1666), .Z(n7399) );
  ANDN U7722 ( .B(n7401), .A(n1733), .Z(n7397) );
  NAND U7723 ( .A(n7402), .B(n7403), .Z(n1733) );
  AND U7724 ( .A(n1750), .B(n1746), .Z(n7403) );
  OR U7725 ( .A(B[704]), .B(A[704]), .Z(n1750) );
  AND U7726 ( .A(n1741), .B(n1737), .Z(n7402) );
  ANDN U7727 ( .B(n1684), .A(n1706), .Z(n7401) );
  NANDN U7728 ( .A(n1665), .B(n7404), .Z(n1651) );
  NAND U7729 ( .A(n7405), .B(n1666), .Z(n7404) );
  OR U7730 ( .A(B[719]), .B(A[719]), .Z(n1666) );
  NANDN U7731 ( .A(n1668), .B(n7406), .Z(n7405) );
  NAND U7732 ( .A(n7407), .B(n1670), .Z(n7406) );
  OR U7733 ( .A(B[718]), .B(A[718]), .Z(n1670) );
  NANDN U7734 ( .A(n1672), .B(n7408), .Z(n7407) );
  NAND U7735 ( .A(n7409), .B(n1675), .Z(n7408) );
  OR U7736 ( .A(B[717]), .B(A[717]), .Z(n1675) );
  NANDN U7737 ( .A(n1677), .B(n7410), .Z(n7409) );
  NAND U7738 ( .A(n7411), .B(n1680), .Z(n7410) );
  OR U7739 ( .A(B[716]), .B(A[716]), .Z(n1680) );
  NANDN U7740 ( .A(n1682), .B(n7412), .Z(n7411) );
  NAND U7741 ( .A(n7413), .B(n1684), .Z(n7412) );
  AND U7742 ( .A(n7414), .B(n7415), .Z(n1684) );
  AND U7743 ( .A(n1702), .B(n1698), .Z(n7415) );
  OR U7744 ( .A(B[712]), .B(A[712]), .Z(n1702) );
  AND U7745 ( .A(n1693), .B(n1689), .Z(n7414) );
  NANDN U7746 ( .A(n1704), .B(n7416), .Z(n7413) );
  NANDN U7747 ( .A(n1706), .B(n1732), .Z(n7416) );
  NANDN U7748 ( .A(n1736), .B(n7417), .Z(n1732) );
  NAND U7749 ( .A(n7418), .B(n1737), .Z(n7417) );
  OR U7750 ( .A(B[707]), .B(A[707]), .Z(n1737) );
  NANDN U7751 ( .A(n1739), .B(n7419), .Z(n7418) );
  NAND U7752 ( .A(n7420), .B(n1741), .Z(n7419) );
  OR U7753 ( .A(B[706]), .B(A[706]), .Z(n1741) );
  NANDN U7754 ( .A(n1743), .B(n7421), .Z(n7420) );
  NAND U7755 ( .A(n1746), .B(n1748), .Z(n7421) );
  AND U7756 ( .A(B[704]), .B(A[704]), .Z(n1748) );
  OR U7757 ( .A(B[705]), .B(A[705]), .Z(n1746) );
  AND U7758 ( .A(B[705]), .B(A[705]), .Z(n1743) );
  AND U7759 ( .A(B[706]), .B(A[706]), .Z(n1739) );
  AND U7760 ( .A(B[707]), .B(A[707]), .Z(n1736) );
  NAND U7761 ( .A(n7422), .B(n7423), .Z(n1706) );
  AND U7762 ( .A(n1729), .B(n1720), .Z(n7423) );
  OR U7763 ( .A(B[708]), .B(A[708]), .Z(n1729) );
  AND U7764 ( .A(n1715), .B(n1711), .Z(n7422) );
  NANDN U7765 ( .A(n1710), .B(n7424), .Z(n1704) );
  NAND U7766 ( .A(n7425), .B(n1711), .Z(n7424) );
  OR U7767 ( .A(B[711]), .B(A[711]), .Z(n1711) );
  NANDN U7768 ( .A(n1713), .B(n7426), .Z(n7425) );
  NAND U7769 ( .A(n7427), .B(n1715), .Z(n7426) );
  OR U7770 ( .A(B[710]), .B(A[710]), .Z(n1715) );
  NANDN U7771 ( .A(n1717), .B(n7428), .Z(n7427) );
  NAND U7772 ( .A(n1720), .B(n1727), .Z(n7428) );
  AND U7773 ( .A(B[708]), .B(A[708]), .Z(n1727) );
  OR U7774 ( .A(B[709]), .B(A[709]), .Z(n1720) );
  AND U7775 ( .A(B[709]), .B(A[709]), .Z(n1717) );
  AND U7776 ( .A(B[710]), .B(A[710]), .Z(n1713) );
  AND U7777 ( .A(B[711]), .B(A[711]), .Z(n1710) );
  NANDN U7778 ( .A(n1688), .B(n7429), .Z(n1682) );
  NAND U7779 ( .A(n7430), .B(n1689), .Z(n7429) );
  OR U7780 ( .A(B[715]), .B(A[715]), .Z(n1689) );
  NANDN U7781 ( .A(n1691), .B(n7431), .Z(n7430) );
  NAND U7782 ( .A(n7432), .B(n1693), .Z(n7431) );
  OR U7783 ( .A(B[714]), .B(A[714]), .Z(n1693) );
  NANDN U7784 ( .A(n1695), .B(n7433), .Z(n7432) );
  NAND U7785 ( .A(n1698), .B(n1700), .Z(n7433) );
  AND U7786 ( .A(B[712]), .B(A[712]), .Z(n1700) );
  OR U7787 ( .A(B[713]), .B(A[713]), .Z(n1698) );
  AND U7788 ( .A(B[713]), .B(A[713]), .Z(n1695) );
  AND U7789 ( .A(B[714]), .B(A[714]), .Z(n1691) );
  AND U7790 ( .A(B[715]), .B(A[715]), .Z(n1688) );
  AND U7791 ( .A(B[716]), .B(A[716]), .Z(n1677) );
  AND U7792 ( .A(B[717]), .B(A[717]), .Z(n1672) );
  AND U7793 ( .A(B[718]), .B(A[718]), .Z(n1668) );
  AND U7794 ( .A(B[719]), .B(A[719]), .Z(n1665) );
  NAND U7795 ( .A(n7434), .B(n7435), .Z(n1560) );
  AND U7796 ( .A(n7436), .B(n7437), .Z(n7435) );
  AND U7797 ( .A(n1579), .B(n1574), .Z(n7437) );
  AND U7798 ( .A(n1569), .B(n1565), .Z(n7436) );
  ANDN U7799 ( .B(n7438), .A(n1632), .Z(n7434) );
  NAND U7800 ( .A(n7439), .B(n7440), .Z(n1632) );
  AND U7801 ( .A(n1649), .B(n1645), .Z(n7440) );
  OR U7802 ( .A(B[720]), .B(A[720]), .Z(n1649) );
  AND U7803 ( .A(n1640), .B(n1636), .Z(n7439) );
  ANDN U7804 ( .B(n1583), .A(n1610), .Z(n7438) );
  NANDN U7805 ( .A(n1564), .B(n7441), .Z(n1558) );
  NAND U7806 ( .A(n7442), .B(n1565), .Z(n7441) );
  OR U7807 ( .A(B[735]), .B(A[735]), .Z(n1565) );
  NANDN U7808 ( .A(n1567), .B(n7443), .Z(n7442) );
  NAND U7809 ( .A(n7444), .B(n1569), .Z(n7443) );
  OR U7810 ( .A(B[734]), .B(A[734]), .Z(n1569) );
  NANDN U7811 ( .A(n1571), .B(n7445), .Z(n7444) );
  NAND U7812 ( .A(n7446), .B(n1574), .Z(n7445) );
  OR U7813 ( .A(B[733]), .B(A[733]), .Z(n1574) );
  NANDN U7814 ( .A(n1576), .B(n7447), .Z(n7446) );
  NAND U7815 ( .A(n7448), .B(n1579), .Z(n7447) );
  OR U7816 ( .A(B[732]), .B(A[732]), .Z(n1579) );
  NANDN U7817 ( .A(n1581), .B(n7449), .Z(n7448) );
  NAND U7818 ( .A(n7450), .B(n1583), .Z(n7449) );
  AND U7819 ( .A(n7451), .B(n7452), .Z(n1583) );
  AND U7820 ( .A(n1606), .B(n1597), .Z(n7452) );
  OR U7821 ( .A(B[728]), .B(A[728]), .Z(n1606) );
  AND U7822 ( .A(n1592), .B(n1588), .Z(n7451) );
  NANDN U7823 ( .A(n1608), .B(n7453), .Z(n7450) );
  NANDN U7824 ( .A(n1610), .B(n1631), .Z(n7453) );
  NANDN U7825 ( .A(n1635), .B(n7454), .Z(n1631) );
  NAND U7826 ( .A(n7455), .B(n1636), .Z(n7454) );
  OR U7827 ( .A(B[723]), .B(A[723]), .Z(n1636) );
  NANDN U7828 ( .A(n1638), .B(n7456), .Z(n7455) );
  NAND U7829 ( .A(n7457), .B(n1640), .Z(n7456) );
  OR U7830 ( .A(B[722]), .B(A[722]), .Z(n1640) );
  NANDN U7831 ( .A(n1642), .B(n7458), .Z(n7457) );
  NAND U7832 ( .A(n1645), .B(n1647), .Z(n7458) );
  AND U7833 ( .A(B[720]), .B(A[720]), .Z(n1647) );
  OR U7834 ( .A(B[721]), .B(A[721]), .Z(n1645) );
  AND U7835 ( .A(B[721]), .B(A[721]), .Z(n1642) );
  AND U7836 ( .A(B[722]), .B(A[722]), .Z(n1638) );
  AND U7837 ( .A(B[723]), .B(A[723]), .Z(n1635) );
  NAND U7838 ( .A(n7459), .B(n7460), .Z(n1610) );
  AND U7839 ( .A(n1628), .B(n1624), .Z(n7460) );
  OR U7840 ( .A(B[724]), .B(A[724]), .Z(n1628) );
  AND U7841 ( .A(n1619), .B(n1615), .Z(n7459) );
  NANDN U7842 ( .A(n1614), .B(n7461), .Z(n1608) );
  NAND U7843 ( .A(n7462), .B(n1615), .Z(n7461) );
  OR U7844 ( .A(B[727]), .B(A[727]), .Z(n1615) );
  NANDN U7845 ( .A(n1617), .B(n7463), .Z(n7462) );
  NAND U7846 ( .A(n7464), .B(n1619), .Z(n7463) );
  OR U7847 ( .A(B[726]), .B(A[726]), .Z(n1619) );
  NANDN U7848 ( .A(n1621), .B(n7465), .Z(n7464) );
  NAND U7849 ( .A(n1624), .B(n1626), .Z(n7465) );
  AND U7850 ( .A(B[724]), .B(A[724]), .Z(n1626) );
  OR U7851 ( .A(B[725]), .B(A[725]), .Z(n1624) );
  AND U7852 ( .A(B[725]), .B(A[725]), .Z(n1621) );
  AND U7853 ( .A(B[726]), .B(A[726]), .Z(n1617) );
  AND U7854 ( .A(B[727]), .B(A[727]), .Z(n1614) );
  NANDN U7855 ( .A(n1587), .B(n7466), .Z(n1581) );
  NAND U7856 ( .A(n7467), .B(n1588), .Z(n7466) );
  OR U7857 ( .A(B[731]), .B(A[731]), .Z(n1588) );
  NANDN U7858 ( .A(n1590), .B(n7468), .Z(n7467) );
  NAND U7859 ( .A(n7469), .B(n1592), .Z(n7468) );
  OR U7860 ( .A(B[730]), .B(A[730]), .Z(n1592) );
  NANDN U7861 ( .A(n1594), .B(n7470), .Z(n7469) );
  NAND U7862 ( .A(n1597), .B(n1604), .Z(n7470) );
  AND U7863 ( .A(B[728]), .B(A[728]), .Z(n1604) );
  OR U7864 ( .A(B[729]), .B(A[729]), .Z(n1597) );
  AND U7865 ( .A(B[729]), .B(A[729]), .Z(n1594) );
  AND U7866 ( .A(B[730]), .B(A[730]), .Z(n1590) );
  AND U7867 ( .A(B[731]), .B(A[731]), .Z(n1587) );
  AND U7868 ( .A(B[732]), .B(A[732]), .Z(n1576) );
  AND U7869 ( .A(B[733]), .B(A[733]), .Z(n1571) );
  AND U7870 ( .A(B[734]), .B(A[734]), .Z(n1567) );
  AND U7871 ( .A(B[735]), .B(A[735]), .Z(n1564) );
  NAND U7872 ( .A(n7471), .B(n7472), .Z(n1463) );
  AND U7873 ( .A(n7473), .B(n7474), .Z(n7472) );
  AND U7874 ( .A(n1487), .B(n1477), .Z(n7474) );
  AND U7875 ( .A(n1472), .B(n1468), .Z(n7473) );
  ANDN U7876 ( .B(n7475), .A(n1535), .Z(n7471) );
  NAND U7877 ( .A(n7476), .B(n7477), .Z(n1535) );
  AND U7878 ( .A(n1556), .B(n1552), .Z(n7477) );
  OR U7879 ( .A(B[736]), .B(A[736]), .Z(n1556) );
  AND U7880 ( .A(n1547), .B(n1543), .Z(n7476) );
  ANDN U7881 ( .B(n1491), .A(n1513), .Z(n7475) );
  NANDN U7882 ( .A(n1467), .B(n7478), .Z(n1461) );
  NAND U7883 ( .A(n7479), .B(n1468), .Z(n7478) );
  OR U7884 ( .A(B[751]), .B(A[751]), .Z(n1468) );
  NANDN U7885 ( .A(n1470), .B(n7480), .Z(n7479) );
  NAND U7886 ( .A(n7481), .B(n1472), .Z(n7480) );
  OR U7887 ( .A(B[750]), .B(A[750]), .Z(n1472) );
  NANDN U7888 ( .A(n1474), .B(n7482), .Z(n7481) );
  NAND U7889 ( .A(n7483), .B(n1477), .Z(n7482) );
  OR U7890 ( .A(B[749]), .B(A[749]), .Z(n1477) );
  NANDN U7891 ( .A(n1484), .B(n7484), .Z(n7483) );
  NAND U7892 ( .A(n7485), .B(n1487), .Z(n7484) );
  OR U7893 ( .A(B[748]), .B(A[748]), .Z(n1487) );
  NANDN U7894 ( .A(n1489), .B(n7486), .Z(n7485) );
  NAND U7895 ( .A(n7487), .B(n1491), .Z(n7486) );
  AND U7896 ( .A(n7488), .B(n7489), .Z(n1491) );
  AND U7897 ( .A(n1509), .B(n1505), .Z(n7489) );
  OR U7898 ( .A(B[744]), .B(A[744]), .Z(n1509) );
  AND U7899 ( .A(n1500), .B(n1496), .Z(n7488) );
  NANDN U7900 ( .A(n1511), .B(n7490), .Z(n7487) );
  NANDN U7901 ( .A(n1513), .B(n1534), .Z(n7490) );
  NANDN U7902 ( .A(n1542), .B(n7491), .Z(n1534) );
  NAND U7903 ( .A(n7492), .B(n1543), .Z(n7491) );
  OR U7904 ( .A(B[739]), .B(A[739]), .Z(n1543) );
  NANDN U7905 ( .A(n1545), .B(n7493), .Z(n7492) );
  NAND U7906 ( .A(n7494), .B(n1547), .Z(n7493) );
  OR U7907 ( .A(B[738]), .B(A[738]), .Z(n1547) );
  NANDN U7908 ( .A(n1549), .B(n7495), .Z(n7494) );
  NAND U7909 ( .A(n1552), .B(n1554), .Z(n7495) );
  AND U7910 ( .A(B[736]), .B(A[736]), .Z(n1554) );
  OR U7911 ( .A(B[737]), .B(A[737]), .Z(n1552) );
  AND U7912 ( .A(B[737]), .B(A[737]), .Z(n1549) );
  AND U7913 ( .A(B[738]), .B(A[738]), .Z(n1545) );
  AND U7914 ( .A(B[739]), .B(A[739]), .Z(n1542) );
  NAND U7915 ( .A(n7496), .B(n7497), .Z(n1513) );
  AND U7916 ( .A(n1531), .B(n1527), .Z(n7497) );
  OR U7917 ( .A(B[740]), .B(A[740]), .Z(n1531) );
  AND U7918 ( .A(n1522), .B(n1518), .Z(n7496) );
  NANDN U7919 ( .A(n1517), .B(n7498), .Z(n1511) );
  NAND U7920 ( .A(n7499), .B(n1518), .Z(n7498) );
  OR U7921 ( .A(B[743]), .B(A[743]), .Z(n1518) );
  NANDN U7922 ( .A(n1520), .B(n7500), .Z(n7499) );
  NAND U7923 ( .A(n7501), .B(n1522), .Z(n7500) );
  OR U7924 ( .A(B[742]), .B(A[742]), .Z(n1522) );
  NANDN U7925 ( .A(n1524), .B(n7502), .Z(n7501) );
  NAND U7926 ( .A(n1527), .B(n1529), .Z(n7502) );
  AND U7927 ( .A(B[740]), .B(A[740]), .Z(n1529) );
  OR U7928 ( .A(B[741]), .B(A[741]), .Z(n1527) );
  AND U7929 ( .A(B[741]), .B(A[741]), .Z(n1524) );
  AND U7930 ( .A(B[742]), .B(A[742]), .Z(n1520) );
  AND U7931 ( .A(B[743]), .B(A[743]), .Z(n1517) );
  NANDN U7932 ( .A(n1495), .B(n7503), .Z(n1489) );
  NAND U7933 ( .A(n7504), .B(n1496), .Z(n7503) );
  OR U7934 ( .A(B[747]), .B(A[747]), .Z(n1496) );
  NANDN U7935 ( .A(n1498), .B(n7505), .Z(n7504) );
  NAND U7936 ( .A(n7506), .B(n1500), .Z(n7505) );
  OR U7937 ( .A(B[746]), .B(A[746]), .Z(n1500) );
  NANDN U7938 ( .A(n1502), .B(n7507), .Z(n7506) );
  NAND U7939 ( .A(n1505), .B(n1507), .Z(n7507) );
  AND U7940 ( .A(B[744]), .B(A[744]), .Z(n1507) );
  OR U7941 ( .A(B[745]), .B(A[745]), .Z(n1505) );
  AND U7942 ( .A(B[745]), .B(A[745]), .Z(n1502) );
  AND U7943 ( .A(B[746]), .B(A[746]), .Z(n1498) );
  AND U7944 ( .A(B[747]), .B(A[747]), .Z(n1495) );
  AND U7945 ( .A(B[748]), .B(A[748]), .Z(n1484) );
  AND U7946 ( .A(B[749]), .B(A[749]), .Z(n1474) );
  AND U7947 ( .A(B[750]), .B(A[750]), .Z(n1470) );
  AND U7948 ( .A(B[751]), .B(A[751]), .Z(n1467) );
  ANDN U7949 ( .B(n7508), .A(n1441), .Z(n5689) );
  NAND U7950 ( .A(n7509), .B(n7510), .Z(n1441) );
  AND U7951 ( .A(n1459), .B(n1455), .Z(n7510) );
  OR U7952 ( .A(B[752]), .B(A[752]), .Z(n1459) );
  ANDN U7953 ( .B(n1446), .A(n1449), .Z(n7509) );
  ANDN U7954 ( .B(n1412), .A(n1389), .Z(n7508) );
  ANDN U7955 ( .B(n7511), .A(n1373), .Z(n5687) );
  AND U7956 ( .A(B[766]), .B(A[766]), .Z(n1373) );
  NAND U7957 ( .A(n7512), .B(n1375), .Z(n7511) );
  OR U7958 ( .A(A[766]), .B(B[766]), .Z(n1375) );
  NANDN U7959 ( .A(n1377), .B(n7513), .Z(n7512) );
  NAND U7960 ( .A(n7514), .B(n1380), .Z(n7513) );
  OR U7961 ( .A(B[765]), .B(A[765]), .Z(n1380) );
  NANDN U7962 ( .A(n1382), .B(n7515), .Z(n7514) );
  NANDN U7963 ( .A(n1384), .B(n7516), .Z(n7515) );
  NANDN U7964 ( .A(n1387), .B(n7517), .Z(n7516) );
  NANDN U7965 ( .A(n1389), .B(n7518), .Z(n7517) );
  NANDN U7966 ( .A(n1409), .B(n7519), .Z(n7518) );
  NAND U7967 ( .A(n1440), .B(n1412), .Z(n7519) );
  AND U7968 ( .A(n7520), .B(n7521), .Z(n1412) );
  AND U7969 ( .A(n1437), .B(n1433), .Z(n7521) );
  OR U7970 ( .A(B[756]), .B(A[756]), .Z(n1437) );
  AND U7971 ( .A(n1428), .B(n1424), .Z(n7520) );
  NANDN U7972 ( .A(n1445), .B(n7522), .Z(n1440) );
  NAND U7973 ( .A(n7523), .B(n1446), .Z(n7522) );
  OR U7974 ( .A(B[755]), .B(A[755]), .Z(n1446) );
  NANDN U7975 ( .A(n1448), .B(n7524), .Z(n7523) );
  NANDN U7976 ( .A(n1449), .B(n7525), .Z(n7524) );
  NANDN U7977 ( .A(n1452), .B(n7526), .Z(n7525) );
  NAND U7978 ( .A(n1455), .B(n1457), .Z(n7526) );
  AND U7979 ( .A(A[752]), .B(B[752]), .Z(n1457) );
  OR U7980 ( .A(B[753]), .B(A[753]), .Z(n1455) );
  AND U7981 ( .A(B[753]), .B(A[753]), .Z(n1452) );
  NOR U7982 ( .A(B[754]), .B(A[754]), .Z(n1449) );
  AND U7983 ( .A(B[754]), .B(A[754]), .Z(n1448) );
  AND U7984 ( .A(B[755]), .B(A[755]), .Z(n1445) );
  NANDN U7985 ( .A(n1423), .B(n7527), .Z(n1409) );
  NAND U7986 ( .A(n7528), .B(n1424), .Z(n7527) );
  OR U7987 ( .A(B[759]), .B(A[759]), .Z(n1424) );
  NANDN U7988 ( .A(n1426), .B(n7529), .Z(n7528) );
  NAND U7989 ( .A(n7530), .B(n1428), .Z(n7529) );
  OR U7990 ( .A(B[758]), .B(A[758]), .Z(n1428) );
  NANDN U7991 ( .A(n1430), .B(n7531), .Z(n7530) );
  NAND U7992 ( .A(n1433), .B(n1435), .Z(n7531) );
  AND U7993 ( .A(B[756]), .B(A[756]), .Z(n1435) );
  OR U7994 ( .A(B[757]), .B(A[757]), .Z(n1433) );
  AND U7995 ( .A(B[757]), .B(A[757]), .Z(n1430) );
  AND U7996 ( .A(B[758]), .B(A[758]), .Z(n1426) );
  AND U7997 ( .A(B[759]), .B(A[759]), .Z(n1423) );
  NAND U7998 ( .A(n7532), .B(n7533), .Z(n1389) );
  AND U7999 ( .A(n1407), .B(n1403), .Z(n7533) );
  OR U8000 ( .A(B[760]), .B(A[760]), .Z(n1407) );
  AND U8001 ( .A(n1398), .B(n1394), .Z(n7532) );
  NANDN U8002 ( .A(n1393), .B(n7534), .Z(n1387) );
  NAND U8003 ( .A(n7535), .B(n1394), .Z(n7534) );
  OR U8004 ( .A(B[763]), .B(A[763]), .Z(n1394) );
  NANDN U8005 ( .A(n1396), .B(n7536), .Z(n7535) );
  NAND U8006 ( .A(n7537), .B(n1398), .Z(n7536) );
  OR U8007 ( .A(B[762]), .B(A[762]), .Z(n1398) );
  NANDN U8008 ( .A(n1400), .B(n7538), .Z(n7537) );
  NAND U8009 ( .A(n1403), .B(n1405), .Z(n7538) );
  AND U8010 ( .A(B[760]), .B(A[760]), .Z(n1405) );
  OR U8011 ( .A(B[761]), .B(A[761]), .Z(n1403) );
  AND U8012 ( .A(B[761]), .B(A[761]), .Z(n1400) );
  AND U8013 ( .A(B[762]), .B(A[762]), .Z(n1396) );
  AND U8014 ( .A(B[763]), .B(A[763]), .Z(n1393) );
  NOR U8015 ( .A(B[764]), .B(A[764]), .Z(n1384) );
  AND U8016 ( .A(B[764]), .B(A[764]), .Z(n1382) );
  AND U8017 ( .A(B[765]), .B(A[765]), .Z(n1377) );
  NOR U8018 ( .A(B[767]), .B(A[767]), .Z(n1370) );
  NOR U8019 ( .A(n1343), .B(n1294), .Z(n5682) );
  NAND U8020 ( .A(n7539), .B(n7540), .Z(n1343) );
  AND U8021 ( .A(n1366), .B(n1357), .Z(n7540) );
  OR U8022 ( .A(B[768]), .B(A[768]), .Z(n1366) );
  ANDN U8023 ( .B(n1348), .A(n1351), .Z(n7539) );
  ANDN U8024 ( .B(n7541), .A(n1287), .Z(n5680) );
  AND U8025 ( .A(B[780]), .B(A[780]), .Z(n1287) );
  NAND U8026 ( .A(n7542), .B(n1290), .Z(n7541) );
  OR U8027 ( .A(A[780]), .B(B[780]), .Z(n1290) );
  NANDN U8028 ( .A(n1292), .B(n7543), .Z(n7542) );
  NANDN U8029 ( .A(n1294), .B(n7544), .Z(n7543) );
  NANDN U8030 ( .A(n1319), .B(n7545), .Z(n7544) );
  NAND U8031 ( .A(n1342), .B(n1322), .Z(n7545) );
  AND U8032 ( .A(n7546), .B(n7547), .Z(n1322) );
  AND U8033 ( .A(n1339), .B(n1335), .Z(n7547) );
  OR U8034 ( .A(B[772]), .B(A[772]), .Z(n1339) );
  AND U8035 ( .A(n1330), .B(n1326), .Z(n7546) );
  NANDN U8036 ( .A(n1347), .B(n7548), .Z(n1342) );
  NAND U8037 ( .A(n7549), .B(n1348), .Z(n7548) );
  OR U8038 ( .A(B[771]), .B(A[771]), .Z(n1348) );
  NANDN U8039 ( .A(n1350), .B(n7550), .Z(n7549) );
  NANDN U8040 ( .A(n1351), .B(n7551), .Z(n7550) );
  NANDN U8041 ( .A(n1354), .B(n7552), .Z(n7551) );
  NAND U8042 ( .A(n1357), .B(n1364), .Z(n7552) );
  AND U8043 ( .A(A[768]), .B(B[768]), .Z(n1364) );
  OR U8044 ( .A(B[769]), .B(A[769]), .Z(n1357) );
  AND U8045 ( .A(B[769]), .B(A[769]), .Z(n1354) );
  NOR U8046 ( .A(B[770]), .B(A[770]), .Z(n1351) );
  AND U8047 ( .A(B[770]), .B(A[770]), .Z(n1350) );
  AND U8048 ( .A(B[771]), .B(A[771]), .Z(n1347) );
  NANDN U8049 ( .A(n1325), .B(n7553), .Z(n1319) );
  NAND U8050 ( .A(n7554), .B(n1326), .Z(n7553) );
  OR U8051 ( .A(B[775]), .B(A[775]), .Z(n1326) );
  NANDN U8052 ( .A(n1328), .B(n7555), .Z(n7554) );
  NAND U8053 ( .A(n7556), .B(n1330), .Z(n7555) );
  OR U8054 ( .A(B[774]), .B(A[774]), .Z(n1330) );
  NANDN U8055 ( .A(n1332), .B(n7557), .Z(n7556) );
  NAND U8056 ( .A(n1335), .B(n1337), .Z(n7557) );
  AND U8057 ( .A(B[772]), .B(A[772]), .Z(n1337) );
  OR U8058 ( .A(B[773]), .B(A[773]), .Z(n1335) );
  AND U8059 ( .A(B[773]), .B(A[773]), .Z(n1332) );
  AND U8060 ( .A(B[774]), .B(A[774]), .Z(n1328) );
  AND U8061 ( .A(B[775]), .B(A[775]), .Z(n1325) );
  NAND U8062 ( .A(n7558), .B(n7559), .Z(n1294) );
  AND U8063 ( .A(n1317), .B(n1313), .Z(n7559) );
  OR U8064 ( .A(B[776]), .B(A[776]), .Z(n1317) );
  AND U8065 ( .A(n1308), .B(n1304), .Z(n7558) );
  NANDN U8066 ( .A(n1303), .B(n7560), .Z(n1292) );
  NAND U8067 ( .A(n7561), .B(n1304), .Z(n7560) );
  OR U8068 ( .A(B[779]), .B(A[779]), .Z(n1304) );
  NANDN U8069 ( .A(n1306), .B(n7562), .Z(n7561) );
  NAND U8070 ( .A(n7563), .B(n1308), .Z(n7562) );
  OR U8071 ( .A(B[778]), .B(A[778]), .Z(n1308) );
  NANDN U8072 ( .A(n1310), .B(n7564), .Z(n7563) );
  NAND U8073 ( .A(n1313), .B(n1315), .Z(n7564) );
  AND U8074 ( .A(B[776]), .B(A[776]), .Z(n1315) );
  OR U8075 ( .A(B[777]), .B(A[777]), .Z(n1313) );
  AND U8076 ( .A(B[777]), .B(A[777]), .Z(n1310) );
  AND U8077 ( .A(B[778]), .B(A[778]), .Z(n1306) );
  AND U8078 ( .A(B[779]), .B(A[779]), .Z(n1303) );
  NOR U8079 ( .A(B[781]), .B(A[781]), .Z(n1284) );
  AND U8080 ( .A(B[781]), .B(A[781]), .Z(n1282) );
  NOR U8081 ( .A(B[782]), .B(A[782]), .Z(n1279) );
  AND U8082 ( .A(B[782]), .B(A[782]), .Z(n1278) );
  NOR U8083 ( .A(B[783]), .B(A[783]), .Z(n1275) );
  NOR U8084 ( .A(n1253), .B(n1204), .Z(n5671) );
  NAND U8085 ( .A(n7565), .B(n7566), .Z(n1253) );
  AND U8086 ( .A(n1271), .B(n1267), .Z(n7566) );
  OR U8087 ( .A(B[784]), .B(A[784]), .Z(n1271) );
  ANDN U8088 ( .B(n1258), .A(n1261), .Z(n7565) );
  ANDN U8089 ( .B(n7567), .A(n1197), .Z(n5669) );
  AND U8090 ( .A(B[796]), .B(A[796]), .Z(n1197) );
  NAND U8091 ( .A(n7568), .B(n1200), .Z(n7567) );
  OR U8092 ( .A(A[796]), .B(B[796]), .Z(n1200) );
  NANDN U8093 ( .A(n1202), .B(n7569), .Z(n7568) );
  NANDN U8094 ( .A(n1204), .B(n7570), .Z(n7569) );
  NANDN U8095 ( .A(n1224), .B(n7571), .Z(n7570) );
  NAND U8096 ( .A(n1252), .B(n1227), .Z(n7571) );
  AND U8097 ( .A(n7572), .B(n7573), .Z(n1227) );
  AND U8098 ( .A(n1249), .B(n1240), .Z(n7573) );
  OR U8099 ( .A(B[788]), .B(A[788]), .Z(n1249) );
  AND U8100 ( .A(n1235), .B(n1231), .Z(n7572) );
  NANDN U8101 ( .A(n1257), .B(n7574), .Z(n1252) );
  NAND U8102 ( .A(n7575), .B(n1258), .Z(n7574) );
  OR U8103 ( .A(B[787]), .B(A[787]), .Z(n1258) );
  NANDN U8104 ( .A(n1260), .B(n7576), .Z(n7575) );
  NANDN U8105 ( .A(n1261), .B(n7577), .Z(n7576) );
  NANDN U8106 ( .A(n1264), .B(n7578), .Z(n7577) );
  NAND U8107 ( .A(n1267), .B(n1269), .Z(n7578) );
  AND U8108 ( .A(A[784]), .B(B[784]), .Z(n1269) );
  OR U8109 ( .A(B[785]), .B(A[785]), .Z(n1267) );
  AND U8110 ( .A(B[785]), .B(A[785]), .Z(n1264) );
  NOR U8111 ( .A(B[786]), .B(A[786]), .Z(n1261) );
  AND U8112 ( .A(B[786]), .B(A[786]), .Z(n1260) );
  AND U8113 ( .A(B[787]), .B(A[787]), .Z(n1257) );
  NANDN U8114 ( .A(n1230), .B(n7579), .Z(n1224) );
  NAND U8115 ( .A(n7580), .B(n1231), .Z(n7579) );
  OR U8116 ( .A(B[791]), .B(A[791]), .Z(n1231) );
  NANDN U8117 ( .A(n1233), .B(n7581), .Z(n7580) );
  NAND U8118 ( .A(n7582), .B(n1235), .Z(n7581) );
  OR U8119 ( .A(B[790]), .B(A[790]), .Z(n1235) );
  NANDN U8120 ( .A(n1237), .B(n7583), .Z(n7582) );
  NAND U8121 ( .A(n1240), .B(n1247), .Z(n7583) );
  AND U8122 ( .A(B[788]), .B(A[788]), .Z(n1247) );
  OR U8123 ( .A(B[789]), .B(A[789]), .Z(n1240) );
  AND U8124 ( .A(B[789]), .B(A[789]), .Z(n1237) );
  AND U8125 ( .A(B[790]), .B(A[790]), .Z(n1233) );
  AND U8126 ( .A(B[791]), .B(A[791]), .Z(n1230) );
  NAND U8127 ( .A(n7584), .B(n7585), .Z(n1204) );
  AND U8128 ( .A(n1222), .B(n1218), .Z(n7585) );
  OR U8129 ( .A(B[792]), .B(A[792]), .Z(n1222) );
  AND U8130 ( .A(n1213), .B(n1209), .Z(n7584) );
  NANDN U8131 ( .A(n1208), .B(n7586), .Z(n1202) );
  NAND U8132 ( .A(n7587), .B(n1209), .Z(n7586) );
  OR U8133 ( .A(B[795]), .B(A[795]), .Z(n1209) );
  NANDN U8134 ( .A(n1211), .B(n7588), .Z(n7587) );
  NAND U8135 ( .A(n7589), .B(n1213), .Z(n7588) );
  OR U8136 ( .A(B[794]), .B(A[794]), .Z(n1213) );
  NANDN U8137 ( .A(n1215), .B(n7590), .Z(n7589) );
  NAND U8138 ( .A(n1218), .B(n1220), .Z(n7590) );
  AND U8139 ( .A(B[792]), .B(A[792]), .Z(n1220) );
  OR U8140 ( .A(B[793]), .B(A[793]), .Z(n1218) );
  AND U8141 ( .A(B[793]), .B(A[793]), .Z(n1215) );
  AND U8142 ( .A(B[794]), .B(A[794]), .Z(n1211) );
  AND U8143 ( .A(B[795]), .B(A[795]), .Z(n1208) );
  NOR U8144 ( .A(B[797]), .B(A[797]), .Z(n1194) );
  AND U8145 ( .A(B[797]), .B(A[797]), .Z(n1192) );
  NOR U8146 ( .A(B[798]), .B(A[798]), .Z(n1189) );
  AND U8147 ( .A(B[798]), .B(A[798]), .Z(n1188) );
  NOR U8148 ( .A(B[799]), .B(A[799]), .Z(n1185) );
  NOR U8149 ( .A(n1149), .B(n1104), .Z(n5660) );
  NAND U8150 ( .A(n7591), .B(n7592), .Z(n1149) );
  AND U8151 ( .A(n1167), .B(n1163), .Z(n7592) );
  OR U8152 ( .A(B[800]), .B(A[800]), .Z(n1167) );
  ANDN U8153 ( .B(n1154), .A(n1157), .Z(n7591) );
  ANDN U8154 ( .B(n7593), .A(n1097), .Z(n5658) );
  AND U8155 ( .A(B[812]), .B(A[812]), .Z(n1097) );
  NAND U8156 ( .A(n7594), .B(n1100), .Z(n7593) );
  OR U8157 ( .A(A[812]), .B(B[812]), .Z(n1100) );
  NANDN U8158 ( .A(n1102), .B(n7595), .Z(n7594) );
  NANDN U8159 ( .A(n1104), .B(n7596), .Z(n7595) );
  NANDN U8160 ( .A(n1125), .B(n7597), .Z(n7596) );
  NAND U8161 ( .A(n1148), .B(n1128), .Z(n7597) );
  AND U8162 ( .A(n7598), .B(n7599), .Z(n1128) );
  AND U8163 ( .A(n1145), .B(n1141), .Z(n7599) );
  OR U8164 ( .A(B[804]), .B(A[804]), .Z(n1145) );
  AND U8165 ( .A(n1136), .B(n1132), .Z(n7598) );
  NANDN U8166 ( .A(n1153), .B(n7600), .Z(n1148) );
  NAND U8167 ( .A(n7601), .B(n1154), .Z(n7600) );
  OR U8168 ( .A(B[803]), .B(A[803]), .Z(n1154) );
  NANDN U8169 ( .A(n1156), .B(n7602), .Z(n7601) );
  NANDN U8170 ( .A(n1157), .B(n7603), .Z(n7602) );
  NANDN U8171 ( .A(n1160), .B(n7604), .Z(n7603) );
  NAND U8172 ( .A(n1163), .B(n1165), .Z(n7604) );
  AND U8173 ( .A(A[800]), .B(B[800]), .Z(n1165) );
  OR U8174 ( .A(B[801]), .B(A[801]), .Z(n1163) );
  AND U8175 ( .A(B[801]), .B(A[801]), .Z(n1160) );
  NOR U8176 ( .A(B[802]), .B(A[802]), .Z(n1157) );
  AND U8177 ( .A(B[802]), .B(A[802]), .Z(n1156) );
  AND U8178 ( .A(B[803]), .B(A[803]), .Z(n1153) );
  NANDN U8179 ( .A(n1131), .B(n7605), .Z(n1125) );
  NAND U8180 ( .A(n7606), .B(n1132), .Z(n7605) );
  OR U8181 ( .A(B[807]), .B(A[807]), .Z(n1132) );
  NANDN U8182 ( .A(n1134), .B(n7607), .Z(n7606) );
  NAND U8183 ( .A(n7608), .B(n1136), .Z(n7607) );
  OR U8184 ( .A(B[806]), .B(A[806]), .Z(n1136) );
  NANDN U8185 ( .A(n1138), .B(n7609), .Z(n7608) );
  NAND U8186 ( .A(n1141), .B(n1143), .Z(n7609) );
  AND U8187 ( .A(B[804]), .B(A[804]), .Z(n1143) );
  OR U8188 ( .A(B[805]), .B(A[805]), .Z(n1141) );
  AND U8189 ( .A(B[805]), .B(A[805]), .Z(n1138) );
  AND U8190 ( .A(B[806]), .B(A[806]), .Z(n1134) );
  AND U8191 ( .A(B[807]), .B(A[807]), .Z(n1131) );
  NAND U8192 ( .A(n7610), .B(n7611), .Z(n1104) );
  AND U8193 ( .A(n1123), .B(n1118), .Z(n7611) );
  OR U8194 ( .A(B[808]), .B(A[808]), .Z(n1123) );
  AND U8195 ( .A(n1113), .B(n1109), .Z(n7610) );
  NANDN U8196 ( .A(n1108), .B(n7612), .Z(n1102) );
  NAND U8197 ( .A(n7613), .B(n1109), .Z(n7612) );
  OR U8198 ( .A(B[811]), .B(A[811]), .Z(n1109) );
  NANDN U8199 ( .A(n1111), .B(n7614), .Z(n7613) );
  NAND U8200 ( .A(n7615), .B(n1113), .Z(n7614) );
  OR U8201 ( .A(B[810]), .B(A[810]), .Z(n1113) );
  NANDN U8202 ( .A(n1115), .B(n7616), .Z(n7615) );
  NAND U8203 ( .A(n1118), .B(n1121), .Z(n7616) );
  AND U8204 ( .A(B[808]), .B(A[808]), .Z(n1121) );
  OR U8205 ( .A(B[809]), .B(A[809]), .Z(n1118) );
  AND U8206 ( .A(B[809]), .B(A[809]), .Z(n1115) );
  AND U8207 ( .A(B[810]), .B(A[810]), .Z(n1111) );
  AND U8208 ( .A(B[811]), .B(A[811]), .Z(n1108) );
  NOR U8209 ( .A(B[813]), .B(A[813]), .Z(n1094) );
  AND U8210 ( .A(B[813]), .B(A[813]), .Z(n1092) );
  NOR U8211 ( .A(B[814]), .B(A[814]), .Z(n1089) );
  AND U8212 ( .A(B[814]), .B(A[814]), .Z(n1088) );
  NOR U8213 ( .A(B[815]), .B(A[815]), .Z(n1085) );
  NOR U8214 ( .A(n1059), .B(n1015), .Z(n5649) );
  NAND U8215 ( .A(n7617), .B(n7618), .Z(n1059) );
  AND U8216 ( .A(n1081), .B(n1077), .Z(n7618) );
  OR U8217 ( .A(B[816]), .B(A[816]), .Z(n1081) );
  ANDN U8218 ( .B(n1068), .A(n1071), .Z(n7617) );
  ANDN U8219 ( .B(n7619), .A(n1008), .Z(n5647) );
  AND U8220 ( .A(B[828]), .B(A[828]), .Z(n1008) );
  NAND U8221 ( .A(n7620), .B(n1011), .Z(n7619) );
  OR U8222 ( .A(A[828]), .B(B[828]), .Z(n1011) );
  NANDN U8223 ( .A(n1013), .B(n7621), .Z(n7620) );
  NANDN U8224 ( .A(n1015), .B(n7622), .Z(n7621) );
  NANDN U8225 ( .A(n1035), .B(n7623), .Z(n7622) );
  NAND U8226 ( .A(n1058), .B(n1038), .Z(n7623) );
  AND U8227 ( .A(n7624), .B(n7625), .Z(n1038) );
  AND U8228 ( .A(n1055), .B(n1051), .Z(n7625) );
  OR U8229 ( .A(B[820]), .B(A[820]), .Z(n1055) );
  AND U8230 ( .A(n1046), .B(n1042), .Z(n7624) );
  NANDN U8231 ( .A(n1067), .B(n7626), .Z(n1058) );
  NAND U8232 ( .A(n7627), .B(n1068), .Z(n7626) );
  OR U8233 ( .A(B[819]), .B(A[819]), .Z(n1068) );
  NANDN U8234 ( .A(n1070), .B(n7628), .Z(n7627) );
  NANDN U8235 ( .A(n1071), .B(n7629), .Z(n7628) );
  NANDN U8236 ( .A(n1074), .B(n7630), .Z(n7629) );
  NAND U8237 ( .A(n1077), .B(n1079), .Z(n7630) );
  AND U8238 ( .A(A[816]), .B(B[816]), .Z(n1079) );
  OR U8239 ( .A(B[817]), .B(A[817]), .Z(n1077) );
  AND U8240 ( .A(B[817]), .B(A[817]), .Z(n1074) );
  NOR U8241 ( .A(B[818]), .B(A[818]), .Z(n1071) );
  AND U8242 ( .A(B[818]), .B(A[818]), .Z(n1070) );
  AND U8243 ( .A(B[819]), .B(A[819]), .Z(n1067) );
  NANDN U8244 ( .A(n1041), .B(n7631), .Z(n1035) );
  NAND U8245 ( .A(n7632), .B(n1042), .Z(n7631) );
  OR U8246 ( .A(B[823]), .B(A[823]), .Z(n1042) );
  NANDN U8247 ( .A(n1044), .B(n7633), .Z(n7632) );
  NAND U8248 ( .A(n7634), .B(n1046), .Z(n7633) );
  OR U8249 ( .A(B[822]), .B(A[822]), .Z(n1046) );
  NANDN U8250 ( .A(n1048), .B(n7635), .Z(n7634) );
  NAND U8251 ( .A(n1051), .B(n1053), .Z(n7635) );
  AND U8252 ( .A(B[820]), .B(A[820]), .Z(n1053) );
  OR U8253 ( .A(B[821]), .B(A[821]), .Z(n1051) );
  AND U8254 ( .A(B[821]), .B(A[821]), .Z(n1048) );
  AND U8255 ( .A(B[822]), .B(A[822]), .Z(n1044) );
  AND U8256 ( .A(B[823]), .B(A[823]), .Z(n1041) );
  NAND U8257 ( .A(n7636), .B(n7637), .Z(n1015) );
  AND U8258 ( .A(n1033), .B(n1029), .Z(n7637) );
  OR U8259 ( .A(B[824]), .B(A[824]), .Z(n1033) );
  AND U8260 ( .A(n1024), .B(n1020), .Z(n7636) );
  NANDN U8261 ( .A(n1019), .B(n7638), .Z(n1013) );
  NAND U8262 ( .A(n7639), .B(n1020), .Z(n7638) );
  OR U8263 ( .A(B[827]), .B(A[827]), .Z(n1020) );
  NANDN U8264 ( .A(n1022), .B(n7640), .Z(n7639) );
  NAND U8265 ( .A(n7641), .B(n1024), .Z(n7640) );
  OR U8266 ( .A(B[826]), .B(A[826]), .Z(n1024) );
  NANDN U8267 ( .A(n1026), .B(n7642), .Z(n7641) );
  NAND U8268 ( .A(n1029), .B(n1031), .Z(n7642) );
  AND U8269 ( .A(B[824]), .B(A[824]), .Z(n1031) );
  OR U8270 ( .A(B[825]), .B(A[825]), .Z(n1029) );
  AND U8271 ( .A(B[825]), .B(A[825]), .Z(n1026) );
  AND U8272 ( .A(B[826]), .B(A[826]), .Z(n1022) );
  AND U8273 ( .A(B[827]), .B(A[827]), .Z(n1019) );
  NOR U8274 ( .A(B[829]), .B(A[829]), .Z(n1000) );
  AND U8275 ( .A(B[829]), .B(A[829]), .Z(n998) );
  NOR U8276 ( .A(B[830]), .B(A[830]), .Z(n995) );
  AND U8277 ( .A(B[830]), .B(A[830]), .Z(n994) );
  NOR U8278 ( .A(B[831]), .B(A[831]), .Z(n991) );
  NOR U8279 ( .A(n969), .B(n917), .Z(n5638) );
  NAND U8280 ( .A(n7643), .B(n7644), .Z(n969) );
  AND U8281 ( .A(n987), .B(n983), .Z(n7644) );
  OR U8282 ( .A(B[832]), .B(A[832]), .Z(n987) );
  ANDN U8283 ( .B(n974), .A(n977), .Z(n7643) );
  ANDN U8284 ( .B(n7645), .A(n910), .Z(n5636) );
  AND U8285 ( .A(B[844]), .B(A[844]), .Z(n910) );
  NAND U8286 ( .A(n7646), .B(n913), .Z(n7645) );
  OR U8287 ( .A(A[844]), .B(B[844]), .Z(n913) );
  NANDN U8288 ( .A(n915), .B(n7647), .Z(n7646) );
  NANDN U8289 ( .A(n917), .B(n7648), .Z(n7647) );
  NANDN U8290 ( .A(n937), .B(n7649), .Z(n7648) );
  NAND U8291 ( .A(n968), .B(n940), .Z(n7649) );
  AND U8292 ( .A(n7650), .B(n7651), .Z(n940) );
  AND U8293 ( .A(n965), .B(n961), .Z(n7651) );
  OR U8294 ( .A(B[836]), .B(A[836]), .Z(n965) );
  AND U8295 ( .A(n956), .B(n952), .Z(n7650) );
  NANDN U8296 ( .A(n973), .B(n7652), .Z(n968) );
  NAND U8297 ( .A(n7653), .B(n974), .Z(n7652) );
  OR U8298 ( .A(B[835]), .B(A[835]), .Z(n974) );
  NANDN U8299 ( .A(n976), .B(n7654), .Z(n7653) );
  NANDN U8300 ( .A(n977), .B(n7655), .Z(n7654) );
  NANDN U8301 ( .A(n980), .B(n7656), .Z(n7655) );
  NAND U8302 ( .A(n983), .B(n985), .Z(n7656) );
  AND U8303 ( .A(A[832]), .B(B[832]), .Z(n985) );
  OR U8304 ( .A(B[833]), .B(A[833]), .Z(n983) );
  AND U8305 ( .A(B[833]), .B(A[833]), .Z(n980) );
  NOR U8306 ( .A(B[834]), .B(A[834]), .Z(n977) );
  AND U8307 ( .A(B[834]), .B(A[834]), .Z(n976) );
  AND U8308 ( .A(B[835]), .B(A[835]), .Z(n973) );
  NANDN U8309 ( .A(n951), .B(n7657), .Z(n937) );
  NAND U8310 ( .A(n7658), .B(n952), .Z(n7657) );
  OR U8311 ( .A(B[839]), .B(A[839]), .Z(n952) );
  NANDN U8312 ( .A(n954), .B(n7659), .Z(n7658) );
  NAND U8313 ( .A(n7660), .B(n956), .Z(n7659) );
  OR U8314 ( .A(B[838]), .B(A[838]), .Z(n956) );
  NANDN U8315 ( .A(n958), .B(n7661), .Z(n7660) );
  NAND U8316 ( .A(n961), .B(n963), .Z(n7661) );
  AND U8317 ( .A(B[836]), .B(A[836]), .Z(n963) );
  OR U8318 ( .A(B[837]), .B(A[837]), .Z(n961) );
  AND U8319 ( .A(B[837]), .B(A[837]), .Z(n958) );
  AND U8320 ( .A(B[838]), .B(A[838]), .Z(n954) );
  AND U8321 ( .A(B[839]), .B(A[839]), .Z(n951) );
  NAND U8322 ( .A(n7662), .B(n7663), .Z(n917) );
  AND U8323 ( .A(n935), .B(n931), .Z(n7663) );
  OR U8324 ( .A(B[840]), .B(A[840]), .Z(n935) );
  AND U8325 ( .A(n926), .B(n922), .Z(n7662) );
  NANDN U8326 ( .A(n921), .B(n7664), .Z(n915) );
  NAND U8327 ( .A(n7665), .B(n922), .Z(n7664) );
  OR U8328 ( .A(B[843]), .B(A[843]), .Z(n922) );
  NANDN U8329 ( .A(n924), .B(n7666), .Z(n7665) );
  NAND U8330 ( .A(n7667), .B(n926), .Z(n7666) );
  OR U8331 ( .A(B[842]), .B(A[842]), .Z(n926) );
  NANDN U8332 ( .A(n928), .B(n7668), .Z(n7667) );
  NAND U8333 ( .A(n931), .B(n933), .Z(n7668) );
  AND U8334 ( .A(B[840]), .B(A[840]), .Z(n933) );
  OR U8335 ( .A(B[841]), .B(A[841]), .Z(n931) );
  AND U8336 ( .A(B[841]), .B(A[841]), .Z(n928) );
  AND U8337 ( .A(B[842]), .B(A[842]), .Z(n924) );
  AND U8338 ( .A(B[843]), .B(A[843]), .Z(n921) );
  NOR U8339 ( .A(B[845]), .B(A[845]), .Z(n907) );
  AND U8340 ( .A(B[845]), .B(A[845]), .Z(n905) );
  NOR U8341 ( .A(B[846]), .B(A[846]), .Z(n902) );
  AND U8342 ( .A(B[846]), .B(A[846]), .Z(n901) );
  NOR U8343 ( .A(B[847]), .B(A[847]), .Z(n898) );
  NOR U8344 ( .A(n871), .B(n823), .Z(n5627) );
  NAND U8345 ( .A(n7669), .B(n7670), .Z(n871) );
  AND U8346 ( .A(n894), .B(n885), .Z(n7670) );
  OR U8347 ( .A(B[848]), .B(A[848]), .Z(n894) );
  ANDN U8348 ( .B(n876), .A(n879), .Z(n7669) );
  ANDN U8349 ( .B(n7671), .A(n816), .Z(n5625) );
  AND U8350 ( .A(B[860]), .B(A[860]), .Z(n816) );
  NAND U8351 ( .A(n7672), .B(n819), .Z(n7671) );
  OR U8352 ( .A(A[860]), .B(B[860]), .Z(n819) );
  NANDN U8353 ( .A(n821), .B(n7673), .Z(n7672) );
  NANDN U8354 ( .A(n823), .B(n7674), .Z(n7673) );
  NANDN U8355 ( .A(n847), .B(n7675), .Z(n7674) );
  NAND U8356 ( .A(n870), .B(n850), .Z(n7675) );
  AND U8357 ( .A(n7676), .B(n7677), .Z(n850) );
  AND U8358 ( .A(n867), .B(n863), .Z(n7677) );
  OR U8359 ( .A(B[852]), .B(A[852]), .Z(n867) );
  AND U8360 ( .A(n858), .B(n854), .Z(n7676) );
  NANDN U8361 ( .A(n875), .B(n7678), .Z(n870) );
  NAND U8362 ( .A(n7679), .B(n876), .Z(n7678) );
  OR U8363 ( .A(B[851]), .B(A[851]), .Z(n876) );
  NANDN U8364 ( .A(n878), .B(n7680), .Z(n7679) );
  NANDN U8365 ( .A(n879), .B(n7681), .Z(n7680) );
  NANDN U8366 ( .A(n882), .B(n7682), .Z(n7681) );
  NAND U8367 ( .A(n885), .B(n892), .Z(n7682) );
  AND U8368 ( .A(A[848]), .B(B[848]), .Z(n892) );
  OR U8369 ( .A(B[849]), .B(A[849]), .Z(n885) );
  AND U8370 ( .A(B[849]), .B(A[849]), .Z(n882) );
  NOR U8371 ( .A(B[850]), .B(A[850]), .Z(n879) );
  AND U8372 ( .A(B[850]), .B(A[850]), .Z(n878) );
  AND U8373 ( .A(B[851]), .B(A[851]), .Z(n875) );
  NANDN U8374 ( .A(n853), .B(n7683), .Z(n847) );
  NAND U8375 ( .A(n7684), .B(n854), .Z(n7683) );
  OR U8376 ( .A(B[855]), .B(A[855]), .Z(n854) );
  NANDN U8377 ( .A(n856), .B(n7685), .Z(n7684) );
  NAND U8378 ( .A(n7686), .B(n858), .Z(n7685) );
  OR U8379 ( .A(B[854]), .B(A[854]), .Z(n858) );
  NANDN U8380 ( .A(n860), .B(n7687), .Z(n7686) );
  NAND U8381 ( .A(n863), .B(n865), .Z(n7687) );
  AND U8382 ( .A(B[852]), .B(A[852]), .Z(n865) );
  OR U8383 ( .A(B[853]), .B(A[853]), .Z(n863) );
  AND U8384 ( .A(B[853]), .B(A[853]), .Z(n860) );
  AND U8385 ( .A(B[854]), .B(A[854]), .Z(n856) );
  AND U8386 ( .A(B[855]), .B(A[855]), .Z(n853) );
  NAND U8387 ( .A(n7688), .B(n7689), .Z(n823) );
  AND U8388 ( .A(n845), .B(n841), .Z(n7689) );
  OR U8389 ( .A(B[856]), .B(A[856]), .Z(n845) );
  AND U8390 ( .A(n836), .B(n832), .Z(n7688) );
  NANDN U8391 ( .A(n831), .B(n7690), .Z(n821) );
  NAND U8392 ( .A(n7691), .B(n832), .Z(n7690) );
  OR U8393 ( .A(B[859]), .B(A[859]), .Z(n832) );
  NANDN U8394 ( .A(n834), .B(n7692), .Z(n7691) );
  NAND U8395 ( .A(n7693), .B(n836), .Z(n7692) );
  OR U8396 ( .A(B[858]), .B(A[858]), .Z(n836) );
  NANDN U8397 ( .A(n838), .B(n7694), .Z(n7693) );
  NAND U8398 ( .A(n841), .B(n843), .Z(n7694) );
  AND U8399 ( .A(B[856]), .B(A[856]), .Z(n843) );
  OR U8400 ( .A(B[857]), .B(A[857]), .Z(n841) );
  AND U8401 ( .A(B[857]), .B(A[857]), .Z(n838) );
  AND U8402 ( .A(B[858]), .B(A[858]), .Z(n834) );
  AND U8403 ( .A(B[859]), .B(A[859]), .Z(n831) );
  NOR U8404 ( .A(B[861]), .B(A[861]), .Z(n813) );
  AND U8405 ( .A(B[861]), .B(A[861]), .Z(n811) );
  NOR U8406 ( .A(B[862]), .B(A[862]), .Z(n808) );
  AND U8407 ( .A(B[862]), .B(A[862]), .Z(n807) );
  NOR U8408 ( .A(B[863]), .B(A[863]), .Z(n804) );
  NOR U8409 ( .A(n782), .B(n733), .Z(n5616) );
  NAND U8410 ( .A(n7695), .B(n7696), .Z(n782) );
  AND U8411 ( .A(n800), .B(n796), .Z(n7696) );
  OR U8412 ( .A(B[864]), .B(A[864]), .Z(n800) );
  ANDN U8413 ( .B(n787), .A(n790), .Z(n7695) );
  ANDN U8414 ( .B(n7697), .A(n726), .Z(n5614) );
  AND U8415 ( .A(B[876]), .B(A[876]), .Z(n726) );
  NAND U8416 ( .A(n7698), .B(n729), .Z(n7697) );
  OR U8417 ( .A(A[876]), .B(B[876]), .Z(n729) );
  NANDN U8418 ( .A(n731), .B(n7699), .Z(n7698) );
  NANDN U8419 ( .A(n733), .B(n7700), .Z(n7699) );
  NANDN U8420 ( .A(n753), .B(n7701), .Z(n7700) );
  NAND U8421 ( .A(n781), .B(n756), .Z(n7701) );
  AND U8422 ( .A(n7702), .B(n7703), .Z(n756) );
  AND U8423 ( .A(n778), .B(n769), .Z(n7703) );
  OR U8424 ( .A(B[868]), .B(A[868]), .Z(n778) );
  AND U8425 ( .A(n764), .B(n760), .Z(n7702) );
  NANDN U8426 ( .A(n786), .B(n7704), .Z(n781) );
  NAND U8427 ( .A(n7705), .B(n787), .Z(n7704) );
  OR U8428 ( .A(B[867]), .B(A[867]), .Z(n787) );
  NANDN U8429 ( .A(n789), .B(n7706), .Z(n7705) );
  NANDN U8430 ( .A(n790), .B(n7707), .Z(n7706) );
  NANDN U8431 ( .A(n793), .B(n7708), .Z(n7707) );
  NAND U8432 ( .A(n796), .B(n798), .Z(n7708) );
  AND U8433 ( .A(A[864]), .B(B[864]), .Z(n798) );
  OR U8434 ( .A(B[865]), .B(A[865]), .Z(n796) );
  AND U8435 ( .A(B[865]), .B(A[865]), .Z(n793) );
  NOR U8436 ( .A(B[866]), .B(A[866]), .Z(n790) );
  AND U8437 ( .A(B[866]), .B(A[866]), .Z(n789) );
  AND U8438 ( .A(B[867]), .B(A[867]), .Z(n786) );
  NANDN U8439 ( .A(n759), .B(n7709), .Z(n753) );
  NAND U8440 ( .A(n7710), .B(n760), .Z(n7709) );
  OR U8441 ( .A(B[871]), .B(A[871]), .Z(n760) );
  NANDN U8442 ( .A(n762), .B(n7711), .Z(n7710) );
  NAND U8443 ( .A(n7712), .B(n764), .Z(n7711) );
  OR U8444 ( .A(B[870]), .B(A[870]), .Z(n764) );
  NANDN U8445 ( .A(n766), .B(n7713), .Z(n7712) );
  NAND U8446 ( .A(n769), .B(n776), .Z(n7713) );
  AND U8447 ( .A(B[868]), .B(A[868]), .Z(n776) );
  OR U8448 ( .A(B[869]), .B(A[869]), .Z(n769) );
  AND U8449 ( .A(B[869]), .B(A[869]), .Z(n766) );
  AND U8450 ( .A(B[870]), .B(A[870]), .Z(n762) );
  AND U8451 ( .A(B[871]), .B(A[871]), .Z(n759) );
  NAND U8452 ( .A(n7714), .B(n7715), .Z(n733) );
  AND U8453 ( .A(n751), .B(n747), .Z(n7715) );
  OR U8454 ( .A(B[872]), .B(A[872]), .Z(n751) );
  AND U8455 ( .A(n742), .B(n738), .Z(n7714) );
  NANDN U8456 ( .A(n737), .B(n7716), .Z(n731) );
  NAND U8457 ( .A(n7717), .B(n738), .Z(n7716) );
  OR U8458 ( .A(B[875]), .B(A[875]), .Z(n738) );
  NANDN U8459 ( .A(n740), .B(n7718), .Z(n7717) );
  NAND U8460 ( .A(n7719), .B(n742), .Z(n7718) );
  OR U8461 ( .A(B[874]), .B(A[874]), .Z(n742) );
  NANDN U8462 ( .A(n744), .B(n7720), .Z(n7719) );
  NAND U8463 ( .A(n747), .B(n749), .Z(n7720) );
  AND U8464 ( .A(B[872]), .B(A[872]), .Z(n749) );
  OR U8465 ( .A(B[873]), .B(A[873]), .Z(n747) );
  AND U8466 ( .A(B[873]), .B(A[873]), .Z(n744) );
  AND U8467 ( .A(B[874]), .B(A[874]), .Z(n740) );
  AND U8468 ( .A(B[875]), .B(A[875]), .Z(n737) );
  NOR U8469 ( .A(B[877]), .B(A[877]), .Z(n723) );
  AND U8470 ( .A(B[877]), .B(A[877]), .Z(n721) );
  NOR U8471 ( .A(B[878]), .B(A[878]), .Z(n718) );
  AND U8472 ( .A(B[878]), .B(A[878]), .Z(n717) );
  NOR U8473 ( .A(B[879]), .B(A[879]), .Z(n714) );
  NOR U8474 ( .A(n684), .B(n635), .Z(n5605) );
  NAND U8475 ( .A(n7721), .B(n7722), .Z(n684) );
  AND U8476 ( .A(n702), .B(n698), .Z(n7722) );
  OR U8477 ( .A(B[880]), .B(A[880]), .Z(n702) );
  ANDN U8478 ( .B(n689), .A(n692), .Z(n7721) );
  ANDN U8479 ( .B(n7723), .A(n628), .Z(n5603) );
  AND U8480 ( .A(B[892]), .B(A[892]), .Z(n628) );
  NAND U8481 ( .A(n7724), .B(n631), .Z(n7723) );
  OR U8482 ( .A(A[892]), .B(B[892]), .Z(n631) );
  NANDN U8483 ( .A(n633), .B(n7725), .Z(n7724) );
  NANDN U8484 ( .A(n635), .B(n7726), .Z(n7725) );
  NANDN U8485 ( .A(n660), .B(n7727), .Z(n7726) );
  NAND U8486 ( .A(n683), .B(n663), .Z(n7727) );
  AND U8487 ( .A(n7728), .B(n7729), .Z(n663) );
  AND U8488 ( .A(n680), .B(n676), .Z(n7729) );
  OR U8489 ( .A(B[884]), .B(A[884]), .Z(n680) );
  AND U8490 ( .A(n671), .B(n667), .Z(n7728) );
  NANDN U8491 ( .A(n688), .B(n7730), .Z(n683) );
  NAND U8492 ( .A(n7731), .B(n689), .Z(n7730) );
  OR U8493 ( .A(B[883]), .B(A[883]), .Z(n689) );
  NANDN U8494 ( .A(n691), .B(n7732), .Z(n7731) );
  NANDN U8495 ( .A(n692), .B(n7733), .Z(n7732) );
  NANDN U8496 ( .A(n695), .B(n7734), .Z(n7733) );
  NAND U8497 ( .A(n698), .B(n700), .Z(n7734) );
  AND U8498 ( .A(A[880]), .B(B[880]), .Z(n700) );
  OR U8499 ( .A(B[881]), .B(A[881]), .Z(n698) );
  AND U8500 ( .A(B[881]), .B(A[881]), .Z(n695) );
  NOR U8501 ( .A(B[882]), .B(A[882]), .Z(n692) );
  AND U8502 ( .A(B[882]), .B(A[882]), .Z(n691) );
  AND U8503 ( .A(B[883]), .B(A[883]), .Z(n688) );
  NANDN U8504 ( .A(n666), .B(n7735), .Z(n660) );
  NAND U8505 ( .A(n7736), .B(n667), .Z(n7735) );
  OR U8506 ( .A(B[887]), .B(A[887]), .Z(n667) );
  NANDN U8507 ( .A(n669), .B(n7737), .Z(n7736) );
  NAND U8508 ( .A(n7738), .B(n671), .Z(n7737) );
  OR U8509 ( .A(B[886]), .B(A[886]), .Z(n671) );
  NANDN U8510 ( .A(n673), .B(n7739), .Z(n7738) );
  NAND U8511 ( .A(n676), .B(n678), .Z(n7739) );
  AND U8512 ( .A(B[884]), .B(A[884]), .Z(n678) );
  OR U8513 ( .A(B[885]), .B(A[885]), .Z(n676) );
  AND U8514 ( .A(B[885]), .B(A[885]), .Z(n673) );
  AND U8515 ( .A(B[886]), .B(A[886]), .Z(n669) );
  AND U8516 ( .A(B[887]), .B(A[887]), .Z(n666) );
  NAND U8517 ( .A(n7740), .B(n7741), .Z(n635) );
  AND U8518 ( .A(n658), .B(n649), .Z(n7741) );
  OR U8519 ( .A(B[888]), .B(A[888]), .Z(n658) );
  AND U8520 ( .A(n644), .B(n640), .Z(n7740) );
  NANDN U8521 ( .A(n639), .B(n7742), .Z(n633) );
  NAND U8522 ( .A(n7743), .B(n640), .Z(n7742) );
  OR U8523 ( .A(B[891]), .B(A[891]), .Z(n640) );
  NANDN U8524 ( .A(n642), .B(n7744), .Z(n7743) );
  NAND U8525 ( .A(n7745), .B(n644), .Z(n7744) );
  OR U8526 ( .A(B[890]), .B(A[890]), .Z(n644) );
  NANDN U8527 ( .A(n646), .B(n7746), .Z(n7745) );
  NAND U8528 ( .A(n649), .B(n656), .Z(n7746) );
  AND U8529 ( .A(B[888]), .B(A[888]), .Z(n656) );
  OR U8530 ( .A(B[889]), .B(A[889]), .Z(n649) );
  AND U8531 ( .A(B[889]), .B(A[889]), .Z(n646) );
  AND U8532 ( .A(B[890]), .B(A[890]), .Z(n642) );
  AND U8533 ( .A(B[891]), .B(A[891]), .Z(n639) );
  NOR U8534 ( .A(B[893]), .B(A[893]), .Z(n625) );
  AND U8535 ( .A(B[893]), .B(A[893]), .Z(n623) );
  NOR U8536 ( .A(B[894]), .B(A[894]), .Z(n620) );
  AND U8537 ( .A(B[894]), .B(A[894]), .Z(n619) );
  NOR U8538 ( .A(B[895]), .B(A[895]), .Z(n616) );
  NOR U8539 ( .A(n586), .B(n542), .Z(n5594) );
  NAND U8540 ( .A(n7747), .B(n7748), .Z(n586) );
  AND U8541 ( .A(n612), .B(n608), .Z(n7748) );
  OR U8542 ( .A(B[896]), .B(A[896]), .Z(n612) );
  ANDN U8543 ( .B(n599), .A(n602), .Z(n7747) );
  ANDN U8544 ( .B(n7749), .A(n535), .Z(n5592) );
  AND U8545 ( .A(B[908]), .B(A[908]), .Z(n535) );
  NAND U8546 ( .A(n7750), .B(n538), .Z(n7749) );
  OR U8547 ( .A(A[908]), .B(B[908]), .Z(n538) );
  NANDN U8548 ( .A(n540), .B(n7751), .Z(n7750) );
  NANDN U8549 ( .A(n542), .B(n7752), .Z(n7751) );
  NANDN U8550 ( .A(n562), .B(n7753), .Z(n7752) );
  NAND U8551 ( .A(n585), .B(n565), .Z(n7753) );
  AND U8552 ( .A(n7754), .B(n7755), .Z(n565) );
  AND U8553 ( .A(n582), .B(n578), .Z(n7755) );
  OR U8554 ( .A(B[900]), .B(A[900]), .Z(n582) );
  AND U8555 ( .A(n573), .B(n569), .Z(n7754) );
  NANDN U8556 ( .A(n598), .B(n7756), .Z(n585) );
  NAND U8557 ( .A(n7757), .B(n599), .Z(n7756) );
  OR U8558 ( .A(B[899]), .B(A[899]), .Z(n599) );
  NANDN U8559 ( .A(n601), .B(n7758), .Z(n7757) );
  NANDN U8560 ( .A(n602), .B(n7759), .Z(n7758) );
  NANDN U8561 ( .A(n605), .B(n7760), .Z(n7759) );
  NAND U8562 ( .A(n608), .B(n610), .Z(n7760) );
  AND U8563 ( .A(A[896]), .B(B[896]), .Z(n610) );
  OR U8564 ( .A(B[897]), .B(A[897]), .Z(n608) );
  AND U8565 ( .A(B[897]), .B(A[897]), .Z(n605) );
  NOR U8566 ( .A(B[898]), .B(A[898]), .Z(n602) );
  AND U8567 ( .A(B[898]), .B(A[898]), .Z(n601) );
  AND U8568 ( .A(B[899]), .B(A[899]), .Z(n598) );
  NANDN U8569 ( .A(n568), .B(n7761), .Z(n562) );
  NAND U8570 ( .A(n7762), .B(n569), .Z(n7761) );
  OR U8571 ( .A(B[903]), .B(A[903]), .Z(n569) );
  NANDN U8572 ( .A(n571), .B(n7763), .Z(n7762) );
  NAND U8573 ( .A(n7764), .B(n573), .Z(n7763) );
  OR U8574 ( .A(B[902]), .B(A[902]), .Z(n573) );
  NANDN U8575 ( .A(n575), .B(n7765), .Z(n7764) );
  NAND U8576 ( .A(n578), .B(n580), .Z(n7765) );
  AND U8577 ( .A(B[900]), .B(A[900]), .Z(n580) );
  OR U8578 ( .A(B[901]), .B(A[901]), .Z(n578) );
  AND U8579 ( .A(B[901]), .B(A[901]), .Z(n575) );
  AND U8580 ( .A(B[902]), .B(A[902]), .Z(n571) );
  AND U8581 ( .A(B[903]), .B(A[903]), .Z(n568) );
  NAND U8582 ( .A(n7766), .B(n7767), .Z(n542) );
  AND U8583 ( .A(n560), .B(n556), .Z(n7767) );
  OR U8584 ( .A(B[904]), .B(A[904]), .Z(n560) );
  AND U8585 ( .A(n551), .B(n547), .Z(n7766) );
  NANDN U8586 ( .A(n546), .B(n7768), .Z(n540) );
  NAND U8587 ( .A(n7769), .B(n547), .Z(n7768) );
  OR U8588 ( .A(B[907]), .B(A[907]), .Z(n547) );
  NANDN U8589 ( .A(n549), .B(n7770), .Z(n7769) );
  NAND U8590 ( .A(n7771), .B(n551), .Z(n7770) );
  OR U8591 ( .A(B[906]), .B(A[906]), .Z(n551) );
  NANDN U8592 ( .A(n553), .B(n7772), .Z(n7771) );
  NAND U8593 ( .A(n556), .B(n558), .Z(n7772) );
  AND U8594 ( .A(B[904]), .B(A[904]), .Z(n558) );
  OR U8595 ( .A(B[905]), .B(A[905]), .Z(n556) );
  AND U8596 ( .A(B[905]), .B(A[905]), .Z(n553) );
  AND U8597 ( .A(B[906]), .B(A[906]), .Z(n549) );
  AND U8598 ( .A(B[907]), .B(A[907]), .Z(n546) );
  NOR U8599 ( .A(B[909]), .B(A[909]), .Z(n527) );
  AND U8600 ( .A(B[909]), .B(A[909]), .Z(n525) );
  NOR U8601 ( .A(B[910]), .B(A[910]), .Z(n522) );
  AND U8602 ( .A(B[910]), .B(A[910]), .Z(n521) );
  NOR U8603 ( .A(B[911]), .B(A[911]), .Z(n518) );
  NOR U8604 ( .A(n496), .B(n444), .Z(n5583) );
  NAND U8605 ( .A(n7773), .B(n7774), .Z(n496) );
  AND U8606 ( .A(n514), .B(n510), .Z(n7774) );
  OR U8607 ( .A(B[912]), .B(A[912]), .Z(n514) );
  ANDN U8608 ( .B(n501), .A(n504), .Z(n7773) );
  ANDN U8609 ( .B(n7775), .A(n437), .Z(n5581) );
  AND U8610 ( .A(B[924]), .B(A[924]), .Z(n437) );
  NAND U8611 ( .A(n7776), .B(n440), .Z(n7775) );
  OR U8612 ( .A(A[924]), .B(B[924]), .Z(n440) );
  NANDN U8613 ( .A(n442), .B(n7777), .Z(n7776) );
  NANDN U8614 ( .A(n444), .B(n7778), .Z(n7777) );
  NANDN U8615 ( .A(n464), .B(n7779), .Z(n7778) );
  NAND U8616 ( .A(n495), .B(n467), .Z(n7779) );
  AND U8617 ( .A(n7780), .B(n7781), .Z(n467) );
  AND U8618 ( .A(n492), .B(n488), .Z(n7781) );
  OR U8619 ( .A(B[916]), .B(A[916]), .Z(n492) );
  AND U8620 ( .A(n483), .B(n479), .Z(n7780) );
  NANDN U8621 ( .A(n500), .B(n7782), .Z(n495) );
  NAND U8622 ( .A(n7783), .B(n501), .Z(n7782) );
  OR U8623 ( .A(B[915]), .B(A[915]), .Z(n501) );
  NANDN U8624 ( .A(n503), .B(n7784), .Z(n7783) );
  NANDN U8625 ( .A(n504), .B(n7785), .Z(n7784) );
  NANDN U8626 ( .A(n507), .B(n7786), .Z(n7785) );
  NAND U8627 ( .A(n510), .B(n512), .Z(n7786) );
  AND U8628 ( .A(A[912]), .B(B[912]), .Z(n512) );
  OR U8629 ( .A(B[913]), .B(A[913]), .Z(n510) );
  AND U8630 ( .A(B[913]), .B(A[913]), .Z(n507) );
  NOR U8631 ( .A(B[914]), .B(A[914]), .Z(n504) );
  AND U8632 ( .A(B[914]), .B(A[914]), .Z(n503) );
  AND U8633 ( .A(B[915]), .B(A[915]), .Z(n500) );
  NANDN U8634 ( .A(n478), .B(n7787), .Z(n464) );
  NAND U8635 ( .A(n7788), .B(n479), .Z(n7787) );
  OR U8636 ( .A(B[919]), .B(A[919]), .Z(n479) );
  NANDN U8637 ( .A(n481), .B(n7789), .Z(n7788) );
  NAND U8638 ( .A(n7790), .B(n483), .Z(n7789) );
  OR U8639 ( .A(B[918]), .B(A[918]), .Z(n483) );
  NANDN U8640 ( .A(n485), .B(n7791), .Z(n7790) );
  NAND U8641 ( .A(n488), .B(n490), .Z(n7791) );
  AND U8642 ( .A(B[916]), .B(A[916]), .Z(n490) );
  OR U8643 ( .A(B[917]), .B(A[917]), .Z(n488) );
  AND U8644 ( .A(B[917]), .B(A[917]), .Z(n485) );
  AND U8645 ( .A(B[918]), .B(A[918]), .Z(n481) );
  AND U8646 ( .A(B[919]), .B(A[919]), .Z(n478) );
  NAND U8647 ( .A(n7792), .B(n7793), .Z(n444) );
  AND U8648 ( .A(n462), .B(n458), .Z(n7793) );
  OR U8649 ( .A(B[920]), .B(A[920]), .Z(n462) );
  AND U8650 ( .A(n453), .B(n449), .Z(n7792) );
  NANDN U8651 ( .A(n448), .B(n7794), .Z(n442) );
  NAND U8652 ( .A(n7795), .B(n449), .Z(n7794) );
  OR U8653 ( .A(B[923]), .B(A[923]), .Z(n449) );
  NANDN U8654 ( .A(n451), .B(n7796), .Z(n7795) );
  NAND U8655 ( .A(n7797), .B(n453), .Z(n7796) );
  OR U8656 ( .A(B[922]), .B(A[922]), .Z(n453) );
  NANDN U8657 ( .A(n455), .B(n7798), .Z(n7797) );
  NAND U8658 ( .A(n458), .B(n460), .Z(n7798) );
  AND U8659 ( .A(B[920]), .B(A[920]), .Z(n460) );
  OR U8660 ( .A(B[921]), .B(A[921]), .Z(n458) );
  AND U8661 ( .A(B[921]), .B(A[921]), .Z(n455) );
  AND U8662 ( .A(B[922]), .B(A[922]), .Z(n451) );
  AND U8663 ( .A(B[923]), .B(A[923]), .Z(n448) );
  NOR U8664 ( .A(B[925]), .B(A[925]), .Z(n434) );
  AND U8665 ( .A(B[925]), .B(A[925]), .Z(n432) );
  NOR U8666 ( .A(B[926]), .B(A[926]), .Z(n429) );
  AND U8667 ( .A(B[926]), .B(A[926]), .Z(n428) );
  NOR U8668 ( .A(B[927]), .B(A[927]), .Z(n425) );
  NOR U8669 ( .A(n398), .B(n349), .Z(n5572) );
  NAND U8670 ( .A(n7799), .B(n7800), .Z(n398) );
  AND U8671 ( .A(n421), .B(n412), .Z(n7800) );
  OR U8672 ( .A(B[928]), .B(A[928]), .Z(n421) );
  ANDN U8673 ( .B(n403), .A(n406), .Z(n7799) );
  ANDN U8674 ( .B(n7801), .A(n342), .Z(n5570) );
  AND U8675 ( .A(B[940]), .B(A[940]), .Z(n342) );
  NAND U8676 ( .A(n7802), .B(n345), .Z(n7801) );
  OR U8677 ( .A(A[940]), .B(B[940]), .Z(n345) );
  NANDN U8678 ( .A(n347), .B(n7803), .Z(n7802) );
  NANDN U8679 ( .A(n349), .B(n7804), .Z(n7803) );
  NANDN U8680 ( .A(n374), .B(n7805), .Z(n7804) );
  NAND U8681 ( .A(n397), .B(n377), .Z(n7805) );
  AND U8682 ( .A(n7806), .B(n7807), .Z(n377) );
  AND U8683 ( .A(n394), .B(n390), .Z(n7807) );
  OR U8684 ( .A(B[932]), .B(A[932]), .Z(n394) );
  AND U8685 ( .A(n385), .B(n381), .Z(n7806) );
  NANDN U8686 ( .A(n402), .B(n7808), .Z(n397) );
  NAND U8687 ( .A(n7809), .B(n403), .Z(n7808) );
  OR U8688 ( .A(B[931]), .B(A[931]), .Z(n403) );
  NANDN U8689 ( .A(n405), .B(n7810), .Z(n7809) );
  NANDN U8690 ( .A(n406), .B(n7811), .Z(n7810) );
  NANDN U8691 ( .A(n409), .B(n7812), .Z(n7811) );
  NAND U8692 ( .A(n412), .B(n419), .Z(n7812) );
  AND U8693 ( .A(A[928]), .B(B[928]), .Z(n419) );
  OR U8694 ( .A(B[929]), .B(A[929]), .Z(n412) );
  AND U8695 ( .A(B[929]), .B(A[929]), .Z(n409) );
  NOR U8696 ( .A(B[930]), .B(A[930]), .Z(n406) );
  AND U8697 ( .A(B[930]), .B(A[930]), .Z(n405) );
  AND U8698 ( .A(B[931]), .B(A[931]), .Z(n402) );
  NANDN U8699 ( .A(n380), .B(n7813), .Z(n374) );
  NAND U8700 ( .A(n7814), .B(n381), .Z(n7813) );
  OR U8701 ( .A(B[935]), .B(A[935]), .Z(n381) );
  NANDN U8702 ( .A(n383), .B(n7815), .Z(n7814) );
  NAND U8703 ( .A(n7816), .B(n385), .Z(n7815) );
  OR U8704 ( .A(B[934]), .B(A[934]), .Z(n385) );
  NANDN U8705 ( .A(n387), .B(n7817), .Z(n7816) );
  NAND U8706 ( .A(n390), .B(n392), .Z(n7817) );
  AND U8707 ( .A(B[932]), .B(A[932]), .Z(n392) );
  OR U8708 ( .A(B[933]), .B(A[933]), .Z(n390) );
  AND U8709 ( .A(B[933]), .B(A[933]), .Z(n387) );
  AND U8710 ( .A(B[934]), .B(A[934]), .Z(n383) );
  AND U8711 ( .A(B[935]), .B(A[935]), .Z(n380) );
  NAND U8712 ( .A(n7818), .B(n7819), .Z(n349) );
  AND U8713 ( .A(n372), .B(n368), .Z(n7819) );
  OR U8714 ( .A(B[936]), .B(A[936]), .Z(n372) );
  AND U8715 ( .A(n363), .B(n359), .Z(n7818) );
  NANDN U8716 ( .A(n358), .B(n7820), .Z(n347) );
  NAND U8717 ( .A(n7821), .B(n359), .Z(n7820) );
  OR U8718 ( .A(B[939]), .B(A[939]), .Z(n359) );
  NANDN U8719 ( .A(n361), .B(n7822), .Z(n7821) );
  NAND U8720 ( .A(n7823), .B(n363), .Z(n7822) );
  OR U8721 ( .A(B[938]), .B(A[938]), .Z(n363) );
  NANDN U8722 ( .A(n365), .B(n7824), .Z(n7823) );
  NAND U8723 ( .A(n368), .B(n370), .Z(n7824) );
  AND U8724 ( .A(B[936]), .B(A[936]), .Z(n370) );
  OR U8725 ( .A(B[937]), .B(A[937]), .Z(n368) );
  AND U8726 ( .A(B[937]), .B(A[937]), .Z(n365) );
  AND U8727 ( .A(B[938]), .B(A[938]), .Z(n361) );
  AND U8728 ( .A(B[939]), .B(A[939]), .Z(n358) );
  NOR U8729 ( .A(B[941]), .B(A[941]), .Z(n339) );
  AND U8730 ( .A(B[941]), .B(A[941]), .Z(n337) );
  NOR U8731 ( .A(B[942]), .B(A[942]), .Z(n334) );
  AND U8732 ( .A(B[942]), .B(A[942]), .Z(n333) );
  NOR U8733 ( .A(B[943]), .B(A[943]), .Z(n330) );
  NOR U8734 ( .A(n308), .B(n259), .Z(n5561) );
  NAND U8735 ( .A(n7825), .B(n7826), .Z(n308) );
  AND U8736 ( .A(n326), .B(n322), .Z(n7826) );
  OR U8737 ( .A(B[944]), .B(A[944]), .Z(n326) );
  ANDN U8738 ( .B(n313), .A(n316), .Z(n7825) );
  ANDN U8739 ( .B(n7827), .A(n252), .Z(n5559) );
  AND U8740 ( .A(B[956]), .B(A[956]), .Z(n252) );
  NAND U8741 ( .A(n7828), .B(n255), .Z(n7827) );
  OR U8742 ( .A(A[956]), .B(B[956]), .Z(n255) );
  NANDN U8743 ( .A(n257), .B(n7829), .Z(n7828) );
  NANDN U8744 ( .A(n259), .B(n7830), .Z(n7829) );
  NANDN U8745 ( .A(n279), .B(n7831), .Z(n7830) );
  NAND U8746 ( .A(n307), .B(n282), .Z(n7831) );
  AND U8747 ( .A(n7832), .B(n7833), .Z(n282) );
  AND U8748 ( .A(n304), .B(n295), .Z(n7833) );
  OR U8749 ( .A(B[948]), .B(A[948]), .Z(n304) );
  AND U8750 ( .A(n290), .B(n286), .Z(n7832) );
  NANDN U8751 ( .A(n312), .B(n7834), .Z(n307) );
  NAND U8752 ( .A(n7835), .B(n313), .Z(n7834) );
  OR U8753 ( .A(B[947]), .B(A[947]), .Z(n313) );
  NANDN U8754 ( .A(n315), .B(n7836), .Z(n7835) );
  NANDN U8755 ( .A(n316), .B(n7837), .Z(n7836) );
  NANDN U8756 ( .A(n319), .B(n7838), .Z(n7837) );
  NAND U8757 ( .A(n322), .B(n324), .Z(n7838) );
  AND U8758 ( .A(A[944]), .B(B[944]), .Z(n324) );
  OR U8759 ( .A(B[945]), .B(A[945]), .Z(n322) );
  AND U8760 ( .A(B[945]), .B(A[945]), .Z(n319) );
  NOR U8761 ( .A(B[946]), .B(A[946]), .Z(n316) );
  AND U8762 ( .A(B[946]), .B(A[946]), .Z(n315) );
  AND U8763 ( .A(B[947]), .B(A[947]), .Z(n312) );
  NANDN U8764 ( .A(n285), .B(n7839), .Z(n279) );
  NAND U8765 ( .A(n7840), .B(n286), .Z(n7839) );
  OR U8766 ( .A(B[951]), .B(A[951]), .Z(n286) );
  NANDN U8767 ( .A(n288), .B(n7841), .Z(n7840) );
  NAND U8768 ( .A(n7842), .B(n290), .Z(n7841) );
  OR U8769 ( .A(B[950]), .B(A[950]), .Z(n290) );
  NANDN U8770 ( .A(n292), .B(n7843), .Z(n7842) );
  NAND U8771 ( .A(n295), .B(n302), .Z(n7843) );
  AND U8772 ( .A(B[948]), .B(A[948]), .Z(n302) );
  OR U8773 ( .A(B[949]), .B(A[949]), .Z(n295) );
  AND U8774 ( .A(B[949]), .B(A[949]), .Z(n292) );
  AND U8775 ( .A(B[950]), .B(A[950]), .Z(n288) );
  AND U8776 ( .A(B[951]), .B(A[951]), .Z(n285) );
  NAND U8777 ( .A(n7844), .B(n7845), .Z(n259) );
  AND U8778 ( .A(n277), .B(n273), .Z(n7845) );
  OR U8779 ( .A(B[952]), .B(A[952]), .Z(n277) );
  AND U8780 ( .A(n268), .B(n264), .Z(n7844) );
  NANDN U8781 ( .A(n263), .B(n7846), .Z(n257) );
  NAND U8782 ( .A(n7847), .B(n264), .Z(n7846) );
  OR U8783 ( .A(B[955]), .B(A[955]), .Z(n264) );
  NANDN U8784 ( .A(n266), .B(n7848), .Z(n7847) );
  NAND U8785 ( .A(n7849), .B(n268), .Z(n7848) );
  OR U8786 ( .A(B[954]), .B(A[954]), .Z(n268) );
  NANDN U8787 ( .A(n270), .B(n7850), .Z(n7849) );
  NAND U8788 ( .A(n273), .B(n275), .Z(n7850) );
  AND U8789 ( .A(B[952]), .B(A[952]), .Z(n275) );
  OR U8790 ( .A(B[953]), .B(A[953]), .Z(n273) );
  AND U8791 ( .A(B[953]), .B(A[953]), .Z(n270) );
  AND U8792 ( .A(B[954]), .B(A[954]), .Z(n266) );
  AND U8793 ( .A(B[955]), .B(A[955]), .Z(n263) );
  NOR U8794 ( .A(B[957]), .B(A[957]), .Z(n249) );
  AND U8795 ( .A(B[957]), .B(A[957]), .Z(n247) );
  NOR U8796 ( .A(B[958]), .B(A[958]), .Z(n244) );
  AND U8797 ( .A(B[958]), .B(A[958]), .Z(n243) );
  NOR U8798 ( .A(B[959]), .B(A[959]), .Z(n240) );
  OR U8799 ( .A(A[961]), .B(B[961]), .Z(n223) );
  AND U8800 ( .A(n218), .B(n214), .Z(n5550) );
  OR U8801 ( .A(B[963]), .B(A[963]), .Z(n214) );
  OR U8802 ( .A(A[962]), .B(B[962]), .Z(n218) );
  NAND U8803 ( .A(n7851), .B(n7852), .Z(n189) );
  AND U8804 ( .A(n207), .B(n203), .Z(n7852) );
  OR U8805 ( .A(A[964]), .B(B[964]), .Z(n207) );
  AND U8806 ( .A(n198), .B(n194), .Z(n7851) );
  NANDN U8807 ( .A(n193), .B(n7853), .Z(n187) );
  NAND U8808 ( .A(n7854), .B(n194), .Z(n7853) );
  OR U8809 ( .A(B[967]), .B(A[967]), .Z(n194) );
  NANDN U8810 ( .A(n196), .B(n7855), .Z(n7854) );
  NAND U8811 ( .A(n7856), .B(n198), .Z(n7855) );
  OR U8812 ( .A(A[966]), .B(B[966]), .Z(n198) );
  NANDN U8813 ( .A(n200), .B(n7857), .Z(n7856) );
  NAND U8814 ( .A(n203), .B(n205), .Z(n7857) );
  AND U8815 ( .A(A[964]), .B(B[964]), .Z(n205) );
  OR U8816 ( .A(A[965]), .B(B[965]), .Z(n203) );
  AND U8817 ( .A(A[965]), .B(B[965]), .Z(n200) );
  AND U8818 ( .A(A[966]), .B(B[966]), .Z(n196) );
  AND U8819 ( .A(B[967]), .B(A[967]), .Z(n193) );
  NAND U8820 ( .A(n7858), .B(n7859), .Z(n166) );
  AND U8821 ( .A(n185), .B(n180), .Z(n7859) );
  OR U8822 ( .A(B[968]), .B(A[968]), .Z(n185) );
  AND U8823 ( .A(n175), .B(n171), .Z(n7858) );
  NANDN U8824 ( .A(n170), .B(n7860), .Z(n164) );
  NAND U8825 ( .A(n7861), .B(n171), .Z(n7860) );
  OR U8826 ( .A(B[971]), .B(A[971]), .Z(n171) );
  NANDN U8827 ( .A(n173), .B(n7862), .Z(n7861) );
  NAND U8828 ( .A(n7863), .B(n175), .Z(n7862) );
  OR U8829 ( .A(B[970]), .B(A[970]), .Z(n175) );
  NANDN U8830 ( .A(n177), .B(n7864), .Z(n7863) );
  NAND U8831 ( .A(n180), .B(n183), .Z(n7864) );
  AND U8832 ( .A(B[968]), .B(A[968]), .Z(n183) );
  OR U8833 ( .A(B[969]), .B(A[969]), .Z(n180) );
  AND U8834 ( .A(B[969]), .B(A[969]), .Z(n177) );
  AND U8835 ( .A(B[970]), .B(A[970]), .Z(n173) );
  AND U8836 ( .A(B[971]), .B(A[971]), .Z(n170) );
  NOR U8837 ( .A(B[972]), .B(A[972]), .Z(n161) );
  AND U8838 ( .A(B[972]), .B(A[972]), .Z(n159) );
  NOR U8839 ( .A(B[973]), .B(A[973]), .Z(n156) );
  AND U8840 ( .A(B[973]), .B(A[973]), .Z(n154) );
  NOR U8841 ( .A(B[974]), .B(A[974]), .Z(n151) );
  AND U8842 ( .A(B[974]), .B(A[974]), .Z(n150) );
  NOR U8843 ( .A(B[975]), .B(A[975]), .Z(n147) );
  OR U8844 ( .A(A[977]), .B(B[977]), .Z(n138) );
  AND U8845 ( .A(n133), .B(n129), .Z(n5529) );
  OR U8846 ( .A(B[979]), .B(A[979]), .Z(n129) );
  OR U8847 ( .A(A[978]), .B(B[978]), .Z(n133) );
  NAND U8848 ( .A(n7865), .B(n7866), .Z(n99) );
  AND U8849 ( .A(n117), .B(n113), .Z(n7866) );
  OR U8850 ( .A(A[980]), .B(B[980]), .Z(n117) );
  AND U8851 ( .A(n108), .B(n104), .Z(n7865) );
  NANDN U8852 ( .A(n103), .B(n7867), .Z(n97) );
  NAND U8853 ( .A(n7868), .B(n104), .Z(n7867) );
  OR U8854 ( .A(B[983]), .B(A[983]), .Z(n104) );
  NANDN U8855 ( .A(n106), .B(n7869), .Z(n7868) );
  NAND U8856 ( .A(n7870), .B(n108), .Z(n7869) );
  OR U8857 ( .A(A[982]), .B(B[982]), .Z(n108) );
  NANDN U8858 ( .A(n110), .B(n7871), .Z(n7870) );
  NAND U8859 ( .A(n113), .B(n115), .Z(n7871) );
  AND U8860 ( .A(A[980]), .B(B[980]), .Z(n115) );
  OR U8861 ( .A(A[981]), .B(B[981]), .Z(n113) );
  AND U8862 ( .A(A[981]), .B(B[981]), .Z(n110) );
  AND U8863 ( .A(A[982]), .B(B[982]), .Z(n106) );
  AND U8864 ( .A(B[983]), .B(A[983]), .Z(n103) );
  NAND U8865 ( .A(n7872), .B(n7873), .Z(n77) );
  AND U8866 ( .A(n95), .B(n91), .Z(n7873) );
  OR U8867 ( .A(B[984]), .B(A[984]), .Z(n95) );
  AND U8868 ( .A(n86), .B(n82), .Z(n7872) );
  NANDN U8869 ( .A(n81), .B(n7874), .Z(n75) );
  NAND U8870 ( .A(n7875), .B(n82), .Z(n7874) );
  OR U8871 ( .A(B[987]), .B(A[987]), .Z(n82) );
  NANDN U8872 ( .A(n84), .B(n7876), .Z(n7875) );
  NAND U8873 ( .A(n7877), .B(n86), .Z(n7876) );
  OR U8874 ( .A(B[986]), .B(A[986]), .Z(n86) );
  NANDN U8875 ( .A(n88), .B(n7878), .Z(n7877) );
  NAND U8876 ( .A(n91), .B(n93), .Z(n7878) );
  AND U8877 ( .A(B[984]), .B(A[984]), .Z(n93) );
  OR U8878 ( .A(B[985]), .B(A[985]), .Z(n91) );
  AND U8879 ( .A(B[985]), .B(A[985]), .Z(n88) );
  AND U8880 ( .A(B[986]), .B(A[986]), .Z(n84) );
  AND U8881 ( .A(B[987]), .B(A[987]), .Z(n81) );
  NOR U8882 ( .A(B[988]), .B(A[988]), .Z(n72) );
  AND U8883 ( .A(B[988]), .B(A[988]), .Z(n70) );
  NOR U8884 ( .A(B[989]), .B(A[989]), .Z(n62) );
  AND U8885 ( .A(B[989]), .B(A[989]), .Z(n60) );
  NOR U8886 ( .A(B[990]), .B(A[990]), .Z(n57) );
  AND U8887 ( .A(B[990]), .B(A[990]), .Z(n56) );
  NOR U8888 ( .A(B[991]), .B(A[991]), .Z(n53) );
  NAND U8889 ( .A(n7879), .B(n7880), .Z(n5461) );
  AND U8890 ( .A(n20), .B(n25), .Z(n7880) );
  AND U8891 ( .A(n16), .B(n30), .Z(n7879) );
  OR U8892 ( .A(B[996]), .B(A[996]), .Z(n30) );
  NANDN U8893 ( .A(n15), .B(n7881), .Z(n5457) );
  NAND U8894 ( .A(n7882), .B(n16), .Z(n7881) );
  OR U8895 ( .A(B[999]), .B(A[999]), .Z(n16) );
  NANDN U8896 ( .A(n18), .B(n7883), .Z(n7882) );
  NAND U8897 ( .A(n7884), .B(n20), .Z(n7883) );
  OR U8898 ( .A(B[998]), .B(A[998]), .Z(n20) );
  NANDN U8899 ( .A(n22), .B(n7885), .Z(n7884) );
  NANDN U8900 ( .A(n27), .B(n25), .Z(n7885) );
  OR U8901 ( .A(B[997]), .B(A[997]), .Z(n25) );
  NAND U8902 ( .A(B[996]), .B(A[996]), .Z(n27) );
  AND U8903 ( .A(B[997]), .B(A[997]), .Z(n22) );
  AND U8904 ( .A(A[998]), .B(B[998]), .Z(n18) );
  AND U8905 ( .A(B[999]), .B(A[999]), .Z(n15) );
endmodule


module mult_N1024_CC256_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [3:0] A;
  input [1023:0] B;
  output [1027:0] PRODUCT;
  input TC;
  wire   \A1[1024] , \A1[1023] , \A1[1022] , \A1[1021] , \A1[1020] ,
         \A1[1019] , \A1[1018] , \A1[1017] , \A1[1016] , \A1[1015] ,
         \A1[1014] , \A1[1013] , \A1[1012] , \A1[1011] , \A1[1010] ,
         \A1[1009] , \A1[1008] , \A1[1007] , \A1[1006] , \A1[1005] ,
         \A1[1004] , \A1[1003] , \A1[1002] , \A1[1001] , \A1[1000] , \A1[999] ,
         \A1[998] , \A1[997] , \A1[996] , \A1[995] , \A1[994] , \A1[993] ,
         \A1[992] , \A1[991] , \A1[990] , \A1[989] , \A1[988] , \A1[987] ,
         \A1[986] , \A1[985] , \A1[984] , \A1[983] , \A1[982] , \A1[981] ,
         \A1[980] , \A1[979] , \A1[978] , \A1[977] , \A1[976] , \A1[975] ,
         \A1[974] , \A1[973] , \A1[972] , \A1[971] , \A1[970] , \A1[969] ,
         \A1[968] , \A1[967] , \A1[966] , \A1[965] , \A1[964] , \A1[963] ,
         \A1[962] , \A1[961] , \A1[960] , \A1[959] , \A1[958] , \A1[957] ,
         \A1[956] , \A1[955] , \A1[954] , \A1[953] , \A1[952] , \A1[951] ,
         \A1[950] , \A1[949] , \A1[948] , \A1[947] , \A1[946] , \A1[945] ,
         \A1[944] , \A1[943] , \A1[942] , \A1[941] , \A1[940] , \A1[939] ,
         \A1[938] , \A1[937] , \A1[936] , \A1[935] , \A1[934] , \A1[933] ,
         \A1[932] , \A1[931] , \A1[930] , \A1[929] , \A1[928] , \A1[927] ,
         \A1[926] , \A1[925] , \A1[924] , \A1[923] , \A1[922] , \A1[921] ,
         \A1[920] , \A1[919] , \A1[918] , \A1[917] , \A1[916] , \A1[915] ,
         \A1[914] , \A1[913] , \A1[912] , \A1[911] , \A1[910] , \A1[909] ,
         \A1[908] , \A1[907] , \A1[906] , \A1[905] , \A1[904] , \A1[903] ,
         \A1[902] , \A1[901] , \A1[900] , \A1[899] , \A1[898] , \A1[897] ,
         \A1[896] , \A1[895] , \A1[894] , \A1[893] , \A1[892] , \A1[891] ,
         \A1[890] , \A1[889] , \A1[888] , \A1[887] , \A1[886] , \A1[885] ,
         \A1[884] , \A1[883] , \A1[882] , \A1[881] , \A1[880] , \A1[879] ,
         \A1[878] , \A1[877] , \A1[876] , \A1[875] , \A1[874] , \A1[873] ,
         \A1[872] , \A1[871] , \A1[870] , \A1[869] , \A1[868] , \A1[867] ,
         \A1[866] , \A1[865] , \A1[864] , \A1[863] , \A1[862] , \A1[861] ,
         \A1[860] , \A1[859] , \A1[858] , \A1[857] , \A1[856] , \A1[855] ,
         \A1[854] , \A1[853] , \A1[852] , \A1[851] , \A1[850] , \A1[849] ,
         \A1[848] , \A1[847] , \A1[846] , \A1[845] , \A1[844] , \A1[843] ,
         \A1[842] , \A1[841] , \A1[840] , \A1[839] , \A1[838] , \A1[837] ,
         \A1[836] , \A1[835] , \A1[834] , \A1[833] , \A1[832] , \A1[831] ,
         \A1[830] , \A1[829] , \A1[828] , \A1[827] , \A1[826] , \A1[825] ,
         \A1[824] , \A1[823] , \A1[822] , \A1[821] , \A1[820] , \A1[819] ,
         \A1[818] , \A1[817] , \A1[816] , \A1[815] , \A1[814] , \A1[813] ,
         \A1[812] , \A1[811] , \A1[810] , \A1[809] , \A1[808] , \A1[807] ,
         \A1[806] , \A1[805] , \A1[804] , \A1[803] , \A1[802] , \A1[801] ,
         \A1[800] , \A1[799] , \A1[798] , \A1[797] , \A1[796] , \A1[795] ,
         \A1[794] , \A1[793] , \A1[792] , \A1[791] , \A1[790] , \A1[789] ,
         \A1[788] , \A1[787] , \A1[786] , \A1[785] , \A1[784] , \A1[783] ,
         \A1[782] , \A1[781] , \A1[780] , \A1[779] , \A1[778] , \A1[777] ,
         \A1[776] , \A1[775] , \A1[774] , \A1[773] , \A1[772] , \A1[771] ,
         \A1[770] , \A1[769] , \A1[768] , \A1[767] , \A1[766] , \A1[765] ,
         \A1[764] , \A1[763] , \A1[762] , \A1[761] , \A1[760] , \A1[759] ,
         \A1[758] , \A1[757] , \A1[756] , \A1[755] , \A1[754] , \A1[753] ,
         \A1[752] , \A1[751] , \A1[750] , \A1[749] , \A1[748] , \A1[747] ,
         \A1[746] , \A1[745] , \A1[744] , \A1[743] , \A1[742] , \A1[741] ,
         \A1[740] , \A1[739] , \A1[738] , \A1[737] , \A1[736] , \A1[735] ,
         \A1[734] , \A1[733] , \A1[732] , \A1[731] , \A1[730] , \A1[729] ,
         \A1[728] , \A1[727] , \A1[726] , \A1[725] , \A1[724] , \A1[723] ,
         \A1[722] , \A1[721] , \A1[720] , \A1[719] , \A1[718] , \A1[717] ,
         \A1[716] , \A1[715] , \A1[714] , \A1[713] , \A1[712] , \A1[711] ,
         \A1[710] , \A1[709] , \A1[708] , \A1[707] , \A1[706] , \A1[705] ,
         \A1[704] , \A1[703] , \A1[702] , \A1[701] , \A1[700] , \A1[699] ,
         \A1[698] , \A1[697] , \A1[696] , \A1[695] , \A1[694] , \A1[693] ,
         \A1[692] , \A1[691] , \A1[690] , \A1[689] , \A1[688] , \A1[687] ,
         \A1[686] , \A1[685] , \A1[684] , \A1[683] , \A1[682] , \A1[681] ,
         \A1[680] , \A1[679] , \A1[678] , \A1[677] , \A1[676] , \A1[675] ,
         \A1[674] , \A1[673] , \A1[672] , \A1[671] , \A1[670] , \A1[669] ,
         \A1[668] , \A1[667] , \A1[666] , \A1[665] , \A1[664] , \A1[663] ,
         \A1[662] , \A1[661] , \A1[660] , \A1[659] , \A1[658] , \A1[657] ,
         \A1[656] , \A1[655] , \A1[654] , \A1[653] , \A1[652] , \A1[651] ,
         \A1[650] , \A1[649] , \A1[648] , \A1[647] , \A1[646] , \A1[645] ,
         \A1[644] , \A1[643] , \A1[642] , \A1[641] , \A1[640] , \A1[639] ,
         \A1[638] , \A1[637] , \A1[636] , \A1[635] , \A1[634] , \A1[633] ,
         \A1[632] , \A1[631] , \A1[630] , \A1[629] , \A1[628] , \A1[627] ,
         \A1[626] , \A1[625] , \A1[624] , \A1[623] , \A1[622] , \A1[621] ,
         \A1[620] , \A1[619] , \A1[618] , \A1[617] , \A1[616] , \A1[615] ,
         \A1[614] , \A1[613] , \A1[612] , \A1[611] , \A1[610] , \A1[609] ,
         \A1[608] , \A1[607] , \A1[606] , \A1[605] , \A1[604] , \A1[603] ,
         \A1[602] , \A1[601] , \A1[600] , \A1[599] , \A1[598] , \A1[597] ,
         \A1[596] , \A1[595] , \A1[594] , \A1[593] , \A1[592] , \A1[591] ,
         \A1[590] , \A1[589] , \A1[588] , \A1[587] , \A1[586] , \A1[585] ,
         \A1[584] , \A1[583] , \A1[582] , \A1[581] , \A1[580] , \A1[579] ,
         \A1[578] , \A1[577] , \A1[576] , \A1[575] , \A1[574] , \A1[573] ,
         \A1[572] , \A1[571] , \A1[570] , \A1[569] , \A1[568] , \A1[567] ,
         \A1[566] , \A1[565] , \A1[564] , \A1[563] , \A1[562] , \A1[561] ,
         \A1[560] , \A1[559] , \A1[558] , \A1[557] , \A1[556] , \A1[555] ,
         \A1[554] , \A1[553] , \A1[552] , \A1[551] , \A1[550] , \A1[549] ,
         \A1[548] , \A1[547] , \A1[546] , \A1[545] , \A1[544] , \A1[543] ,
         \A1[542] , \A1[541] , \A1[540] , \A1[539] , \A1[538] , \A1[537] ,
         \A1[536] , \A1[535] , \A1[534] , \A1[533] , \A1[532] , \A1[531] ,
         \A1[530] , \A1[529] , \A1[528] , \A1[527] , \A1[526] , \A1[525] ,
         \A1[524] , \A1[523] , \A1[522] , \A1[521] , \A1[520] , \A1[519] ,
         \A1[518] , \A1[517] , \A1[516] , \A1[515] , \A1[514] , \A1[513] ,
         \A1[512] , \A1[511] , \A1[510] , \A1[509] , \A1[508] , \A1[507] ,
         \A1[506] , \A1[505] , \A1[504] , \A1[503] , \A1[502] , \A1[501] ,
         \A1[500] , \A1[499] , \A1[498] , \A1[497] , \A1[496] , \A1[495] ,
         \A1[494] , \A1[493] , \A1[492] , \A1[491] , \A1[490] , \A1[489] ,
         \A1[488] , \A1[487] , \A1[486] , \A1[485] , \A1[484] , \A1[483] ,
         \A1[482] , \A1[481] , \A1[480] , \A1[479] , \A1[478] , \A1[477] ,
         \A1[476] , \A1[475] , \A1[474] , \A1[473] , \A1[472] , \A1[471] ,
         \A1[470] , \A1[469] , \A1[468] , \A1[467] , \A1[466] , \A1[465] ,
         \A1[464] , \A1[463] , \A1[462] , \A1[461] , \A1[460] , \A1[459] ,
         \A1[458] , \A1[457] , \A1[456] , \A1[455] , \A1[454] , \A1[453] ,
         \A1[452] , \A1[451] , \A1[450] , \A1[449] , \A1[448] , \A1[447] ,
         \A1[446] , \A1[445] , \A1[444] , \A1[443] , \A1[442] , \A1[441] ,
         \A1[440] , \A1[439] , \A1[438] , \A1[437] , \A1[436] , \A1[435] ,
         \A1[434] , \A1[433] , \A1[432] , \A1[431] , \A1[430] , \A1[429] ,
         \A1[428] , \A1[427] , \A1[426] , \A1[425] , \A1[424] , \A1[423] ,
         \A1[422] , \A1[421] , \A1[420] , \A1[419] , \A1[418] , \A1[417] ,
         \A1[416] , \A1[415] , \A1[414] , \A1[413] , \A1[412] , \A1[411] ,
         \A1[410] , \A1[409] , \A1[408] , \A1[407] , \A1[406] , \A1[405] ,
         \A1[404] , \A1[403] , \A1[402] , \A1[401] , \A1[400] , \A1[399] ,
         \A1[398] , \A1[397] , \A1[396] , \A1[395] , \A1[394] , \A1[393] ,
         \A1[392] , \A1[391] , \A1[390] , \A1[389] , \A1[388] , \A1[387] ,
         \A1[386] , \A1[385] , \A1[384] , \A1[383] , \A1[382] , \A1[381] ,
         \A1[380] , \A1[379] , \A1[378] , \A1[377] , \A1[376] , \A1[375] ,
         \A1[374] , \A1[373] , \A1[372] , \A1[371] , \A1[370] , \A1[369] ,
         \A1[368] , \A1[367] , \A1[366] , \A1[365] , \A1[364] , \A1[363] ,
         \A1[362] , \A1[361] , \A1[360] , \A1[359] , \A1[358] , \A1[357] ,
         \A1[356] , \A1[355] , \A1[354] , \A1[353] , \A1[352] , \A1[351] ,
         \A1[350] , \A1[349] , \A1[348] , \A1[347] , \A1[346] , \A1[345] ,
         \A1[344] , \A1[343] , \A1[342] , \A1[341] , \A1[340] , \A1[339] ,
         \A1[338] , \A1[337] , \A1[336] , \A1[335] , \A1[334] , \A1[333] ,
         \A1[332] , \A1[331] , \A1[330] , \A1[329] , \A1[328] , \A1[327] ,
         \A1[326] , \A1[325] , \A1[324] , \A1[323] , \A1[322] , \A1[321] ,
         \A1[320] , \A1[319] , \A1[318] , \A1[317] , \A1[316] , \A1[315] ,
         \A1[314] , \A1[313] , \A1[312] , \A1[311] , \A1[310] , \A1[309] ,
         \A1[308] , \A1[307] , \A1[306] , \A1[305] , \A1[304] , \A1[303] ,
         \A1[302] , \A1[301] , \A1[300] , \A1[299] , \A1[298] , \A1[297] ,
         \A1[296] , \A1[295] , \A1[294] , \A1[293] , \A1[292] , \A1[291] ,
         \A1[290] , \A1[289] , \A1[288] , \A1[287] , \A1[286] , \A1[285] ,
         \A1[284] , \A1[283] , \A1[282] , \A1[281] , \A1[280] , \A1[279] ,
         \A1[278] , \A1[277] , \A1[276] , \A1[275] , \A1[274] , \A1[273] ,
         \A1[272] , \A1[271] , \A1[270] , \A1[269] , \A1[268] , \A1[267] ,
         \A1[266] , \A1[265] , \A1[264] , \A1[263] , \A1[262] , \A1[261] ,
         \A1[260] , \A1[259] , \A1[258] , \A1[257] , \A1[256] , \A1[255] ,
         \A1[254] , \A1[253] , \A1[252] , \A1[251] , \A1[250] , \A1[249] ,
         \A1[248] , \A1[247] , \A1[246] , \A1[245] , \A1[244] , \A1[243] ,
         \A1[242] , \A1[241] , \A1[240] , \A1[239] , \A1[238] , \A1[237] ,
         \A1[236] , \A1[235] , \A1[234] , \A1[233] , \A1[232] , \A1[231] ,
         \A1[230] , \A1[229] , \A1[228] , \A1[227] , \A1[226] , \A1[225] ,
         \A1[224] , \A1[223] , \A1[222] , \A1[221] , \A1[220] , \A1[219] ,
         \A1[218] , \A1[217] , \A1[216] , \A1[215] , \A1[214] , \A1[213] ,
         \A1[212] , \A1[211] , \A1[210] , \A1[209] , \A1[208] , \A1[207] ,
         \A1[206] , \A1[205] , \A1[204] , \A1[203] , \A1[202] , \A1[201] ,
         \A1[200] , \A1[199] , \A1[198] , \A1[197] , \A1[196] , \A1[195] ,
         \A1[194] , \A1[193] , \A1[192] , \A1[191] , \A1[190] , \A1[189] ,
         \A1[188] , \A1[187] , \A1[186] , \A1[185] , \A1[184] , \A1[183] ,
         \A1[182] , \A1[181] , \A1[180] , \A1[179] , \A1[178] , \A1[177] ,
         \A1[176] , \A1[175] , \A1[174] , \A1[173] , \A1[172] , \A1[171] ,
         \A1[170] , \A1[169] , \A1[168] , \A1[167] , \A1[166] , \A1[165] ,
         \A1[164] , \A1[163] , \A1[162] , \A1[161] , \A1[160] , \A1[159] ,
         \A1[158] , \A1[157] , \A1[156] , \A1[155] , \A1[154] , \A1[153] ,
         \A1[152] , \A1[151] , \A1[150] , \A1[149] , \A1[148] , \A1[147] ,
         \A1[146] , \A1[145] , \A1[144] , \A1[143] , \A1[142] , \A1[141] ,
         \A1[140] , \A1[139] , \A1[138] , \A1[137] , \A1[136] , \A1[135] ,
         \A1[134] , \A1[133] , \A1[132] , \A1[131] , \A1[130] , \A1[129] ,
         \A1[128] , \A1[127] , \A1[126] , \A1[125] , \A1[124] , \A1[123] ,
         \A1[122] , \A1[121] , \A1[120] , \A1[119] , \A1[118] , \A1[117] ,
         \A1[116] , \A1[115] , \A1[114] , \A1[113] , \A1[112] , \A1[111] ,
         \A1[110] , \A1[109] , \A1[108] , \A1[107] , \A1[106] , \A1[105] ,
         \A1[104] , \A1[103] , \A1[102] , \A1[101] , \A1[100] , \A1[99] ,
         \A1[98] , \A1[97] , \A1[96] , \A1[95] , \A1[94] , \A1[93] , \A1[92] ,
         \A1[91] , \A1[90] , \A1[89] , \A1[88] , \A1[87] , \A1[86] , \A1[85] ,
         \A1[84] , \A1[83] , \A1[82] , \A1[81] , \A1[80] , \A1[79] , \A1[78] ,
         \A1[77] , \A1[76] , \A1[75] , \A1[74] , \A1[73] , \A1[72] , \A1[71] ,
         \A1[70] , \A1[69] , \A1[68] , \A1[67] , \A1[66] , \A1[65] , \A1[64] ,
         \A1[63] , \A1[62] , \A1[61] , \A1[60] , \A1[59] , \A1[58] , \A1[57] ,
         \A1[56] , \A1[55] , \A1[54] , \A1[53] , \A1[52] , \A1[51] , \A1[50] ,
         \A1[49] , \A1[48] , \A1[47] , \A1[46] , \A1[45] , \A1[44] , \A1[43] ,
         \A1[42] , \A1[41] , \A1[40] , \A1[39] , \A1[38] , \A1[37] , \A1[36] ,
         \A1[35] , \A1[34] , \A1[33] , \A1[32] , \A1[31] , \A1[30] , \A1[29] ,
         \A1[28] , \A1[27] , \A1[26] , \A1[25] , \A1[24] , \A1[23] , \A1[22] ,
         \A1[21] , \A1[20] , \A1[19] , \A1[18] , \A1[17] , \A1[16] , \A1[15] ,
         \A1[14] , \A1[13] , \A1[12] , \A1[11] , \A1[10] , \A1[9] , \A1[8] ,
         \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] , \A1[1] ,
         \A1[0] , \A2[1025] , \A2[1024] , \A2[1023] , \A2[1022] , \A2[1021] ,
         \A2[1020] , \A2[1019] , \A2[1018] , \A2[1017] , \A2[1016] ,
         \A2[1015] , \A2[1014] , \A2[1013] , \A2[1012] , \A2[1011] ,
         \A2[1010] , \A2[1009] , \A2[1008] , \A2[1007] , \A2[1006] ,
         \A2[1005] , \A2[1004] , \A2[1003] , \A2[1002] , \A2[1001] ,
         \A2[1000] , \A2[999] , \A2[998] , \A2[997] , \A2[996] , \A2[995] ,
         \A2[994] , \A2[993] , \A2[992] , \A2[991] , \A2[990] , \A2[989] ,
         \A2[988] , \A2[987] , \A2[986] , \A2[985] , \A2[984] , \A2[983] ,
         \A2[982] , \A2[981] , \A2[980] , \A2[979] , \A2[978] , \A2[977] ,
         \A2[976] , \A2[975] , \A2[974] , \A2[973] , \A2[972] , \A2[971] ,
         \A2[970] , \A2[969] , \A2[968] , \A2[967] , \A2[966] , \A2[965] ,
         \A2[964] , \A2[963] , \A2[962] , \A2[961] , \A2[960] , \A2[959] ,
         \A2[958] , \A2[957] , \A2[956] , \A2[955] , \A2[954] , \A2[953] ,
         \A2[952] , \A2[951] , \A2[950] , \A2[949] , \A2[948] , \A2[947] ,
         \A2[946] , \A2[945] , \A2[944] , \A2[943] , \A2[942] , \A2[941] ,
         \A2[940] , \A2[939] , \A2[938] , \A2[937] , \A2[936] , \A2[935] ,
         \A2[934] , \A2[933] , \A2[932] , \A2[931] , \A2[930] , \A2[929] ,
         \A2[928] , \A2[927] , \A2[926] , \A2[925] , \A2[924] , \A2[923] ,
         \A2[922] , \A2[921] , \A2[920] , \A2[919] , \A2[918] , \A2[917] ,
         \A2[916] , \A2[915] , \A2[914] , \A2[913] , \A2[912] , \A2[911] ,
         \A2[910] , \A2[909] , \A2[908] , \A2[907] , \A2[906] , \A2[905] ,
         \A2[904] , \A2[903] , \A2[902] , \A2[901] , \A2[900] , \A2[899] ,
         \A2[898] , \A2[897] , \A2[896] , \A2[895] , \A2[894] , \A2[893] ,
         \A2[892] , \A2[891] , \A2[890] , \A2[889] , \A2[888] , \A2[887] ,
         \A2[886] , \A2[885] , \A2[884] , \A2[883] , \A2[882] , \A2[881] ,
         \A2[880] , \A2[879] , \A2[878] , \A2[877] , \A2[876] , \A2[875] ,
         \A2[874] , \A2[873] , \A2[872] , \A2[871] , \A2[870] , \A2[869] ,
         \A2[868] , \A2[867] , \A2[866] , \A2[865] , \A2[864] , \A2[863] ,
         \A2[862] , \A2[861] , \A2[860] , \A2[859] , \A2[858] , \A2[857] ,
         \A2[856] , \A2[855] , \A2[854] , \A2[853] , \A2[852] , \A2[851] ,
         \A2[850] , \A2[849] , \A2[848] , \A2[847] , \A2[846] , \A2[845] ,
         \A2[844] , \A2[843] , \A2[842] , \A2[841] , \A2[840] , \A2[839] ,
         \A2[838] , \A2[837] , \A2[836] , \A2[835] , \A2[834] , \A2[833] ,
         \A2[832] , \A2[831] , \A2[830] , \A2[829] , \A2[828] , \A2[827] ,
         \A2[826] , \A2[825] , \A2[824] , \A2[823] , \A2[822] , \A2[821] ,
         \A2[820] , \A2[819] , \A2[818] , \A2[817] , \A2[816] , \A2[815] ,
         \A2[814] , \A2[813] , \A2[812] , \A2[811] , \A2[810] , \A2[809] ,
         \A2[808] , \A2[807] , \A2[806] , \A2[805] , \A2[804] , \A2[803] ,
         \A2[802] , \A2[801] , \A2[800] , \A2[799] , \A2[798] , \A2[797] ,
         \A2[796] , \A2[795] , \A2[794] , \A2[793] , \A2[792] , \A2[791] ,
         \A2[790] , \A2[789] , \A2[788] , \A2[787] , \A2[786] , \A2[785] ,
         \A2[784] , \A2[783] , \A2[782] , \A2[781] , \A2[780] , \A2[779] ,
         \A2[778] , \A2[777] , \A2[776] , \A2[775] , \A2[774] , \A2[773] ,
         \A2[772] , \A2[771] , \A2[770] , \A2[769] , \A2[768] , \A2[767] ,
         \A2[766] , \A2[765] , \A2[764] , \A2[763] , \A2[762] , \A2[761] ,
         \A2[760] , \A2[759] , \A2[758] , \A2[757] , \A2[756] , \A2[755] ,
         \A2[754] , \A2[753] , \A2[752] , \A2[751] , \A2[750] , \A2[749] ,
         \A2[748] , \A2[747] , \A2[746] , \A2[745] , \A2[744] , \A2[743] ,
         \A2[742] , \A2[741] , \A2[740] , \A2[739] , \A2[738] , \A2[737] ,
         \A2[736] , \A2[735] , \A2[734] , \A2[733] , \A2[732] , \A2[731] ,
         \A2[730] , \A2[729] , \A2[728] , \A2[727] , \A2[726] , \A2[725] ,
         \A2[724] , \A2[723] , \A2[722] , \A2[721] , \A2[720] , \A2[719] ,
         \A2[718] , \A2[717] , \A2[716] , \A2[715] , \A2[714] , \A2[713] ,
         \A2[712] , \A2[711] , \A2[710] , \A2[709] , \A2[708] , \A2[707] ,
         \A2[706] , \A2[705] , \A2[704] , \A2[703] , \A2[702] , \A2[701] ,
         \A2[700] , \A2[699] , \A2[698] , \A2[697] , \A2[696] , \A2[695] ,
         \A2[694] , \A2[693] , \A2[692] , \A2[691] , \A2[690] , \A2[689] ,
         \A2[688] , \A2[687] , \A2[686] , \A2[685] , \A2[684] , \A2[683] ,
         \A2[682] , \A2[681] , \A2[680] , \A2[679] , \A2[678] , \A2[677] ,
         \A2[676] , \A2[675] , \A2[674] , \A2[673] , \A2[672] , \A2[671] ,
         \A2[670] , \A2[669] , \A2[668] , \A2[667] , \A2[666] , \A2[665] ,
         \A2[664] , \A2[663] , \A2[662] , \A2[661] , \A2[660] , \A2[659] ,
         \A2[658] , \A2[657] , \A2[656] , \A2[655] , \A2[654] , \A2[653] ,
         \A2[652] , \A2[651] , \A2[650] , \A2[649] , \A2[648] , \A2[647] ,
         \A2[646] , \A2[645] , \A2[644] , \A2[643] , \A2[642] , \A2[641] ,
         \A2[640] , \A2[639] , \A2[638] , \A2[637] , \A2[636] , \A2[635] ,
         \A2[634] , \A2[633] , \A2[632] , \A2[631] , \A2[630] , \A2[629] ,
         \A2[628] , \A2[627] , \A2[626] , \A2[625] , \A2[624] , \A2[623] ,
         \A2[622] , \A2[621] , \A2[620] , \A2[619] , \A2[618] , \A2[617] ,
         \A2[616] , \A2[615] , \A2[614] , \A2[613] , \A2[612] , \A2[611] ,
         \A2[610] , \A2[609] , \A2[608] , \A2[607] , \A2[606] , \A2[605] ,
         \A2[604] , \A2[603] , \A2[602] , \A2[601] , \A2[600] , \A2[599] ,
         \A2[598] , \A2[597] , \A2[596] , \A2[595] , \A2[594] , \A2[593] ,
         \A2[592] , \A2[591] , \A2[590] , \A2[589] , \A2[588] , \A2[587] ,
         \A2[586] , \A2[585] , \A2[584] , \A2[583] , \A2[582] , \A2[581] ,
         \A2[580] , \A2[579] , \A2[578] , \A2[577] , \A2[576] , \A2[575] ,
         \A2[574] , \A2[573] , \A2[572] , \A2[571] , \A2[570] , \A2[569] ,
         \A2[568] , \A2[567] , \A2[566] , \A2[565] , \A2[564] , \A2[563] ,
         \A2[562] , \A2[561] , \A2[560] , \A2[559] , \A2[558] , \A2[557] ,
         \A2[556] , \A2[555] , \A2[554] , \A2[553] , \A2[552] , \A2[551] ,
         \A2[550] , \A2[549] , \A2[548] , \A2[547] , \A2[546] , \A2[545] ,
         \A2[544] , \A2[543] , \A2[542] , \A2[541] , \A2[540] , \A2[539] ,
         \A2[538] , \A2[537] , \A2[536] , \A2[535] , \A2[534] , \A2[533] ,
         \A2[532] , \A2[531] , \A2[530] , \A2[529] , \A2[528] , \A2[527] ,
         \A2[526] , \A2[525] , \A2[524] , \A2[523] , \A2[522] , \A2[521] ,
         \A2[520] , \A2[519] , \A2[518] , \A2[517] , \A2[516] , \A2[515] ,
         \A2[514] , \A2[513] , \A2[512] , \A2[511] , \A2[510] , \A2[509] ,
         \A2[508] , \A2[507] , \A2[506] , \A2[505] , \A2[504] , \A2[503] ,
         \A2[502] , \A2[501] , \A2[500] , \A2[499] , \A2[498] , \A2[497] ,
         \A2[496] , \A2[495] , \A2[494] , \A2[493] , \A2[492] , \A2[491] ,
         \A2[490] , \A2[489] , \A2[488] , \A2[487] , \A2[486] , \A2[485] ,
         \A2[484] , \A2[483] , \A2[482] , \A2[481] , \A2[480] , \A2[479] ,
         \A2[478] , \A2[477] , \A2[476] , \A2[475] , \A2[474] , \A2[473] ,
         \A2[472] , \A2[471] , \A2[470] , \A2[469] , \A2[468] , \A2[467] ,
         \A2[466] , \A2[465] , \A2[464] , \A2[463] , \A2[462] , \A2[461] ,
         \A2[460] , \A2[459] , \A2[458] , \A2[457] , \A2[456] , \A2[455] ,
         \A2[454] , \A2[453] , \A2[452] , \A2[451] , \A2[450] , \A2[449] ,
         \A2[448] , \A2[447] , \A2[446] , \A2[445] , \A2[444] , \A2[443] ,
         \A2[442] , \A2[441] , \A2[440] , \A2[439] , \A2[438] , \A2[437] ,
         \A2[436] , \A2[435] , \A2[434] , \A2[433] , \A2[432] , \A2[431] ,
         \A2[430] , \A2[429] , \A2[428] , \A2[427] , \A2[426] , \A2[425] ,
         \A2[424] , \A2[423] , \A2[422] , \A2[421] , \A2[420] , \A2[419] ,
         \A2[418] , \A2[417] , \A2[416] , \A2[415] , \A2[414] , \A2[413] ,
         \A2[412] , \A2[411] , \A2[410] , \A2[409] , \A2[408] , \A2[407] ,
         \A2[406] , \A2[405] , \A2[404] , \A2[403] , \A2[402] , \A2[401] ,
         \A2[400] , \A2[399] , \A2[398] , \A2[397] , \A2[396] , \A2[395] ,
         \A2[394] , \A2[393] , \A2[392] , \A2[391] , \A2[390] , \A2[389] ,
         \A2[388] , \A2[387] , \A2[386] , \A2[385] , \A2[384] , \A2[383] ,
         \A2[382] , \A2[381] , \A2[380] , \A2[379] , \A2[378] , \A2[377] ,
         \A2[376] , \A2[375] , \A2[374] , \A2[373] , \A2[372] , \A2[371] ,
         \A2[370] , \A2[369] , \A2[368] , \A2[367] , \A2[366] , \A2[365] ,
         \A2[364] , \A2[363] , \A2[362] , \A2[361] , \A2[360] , \A2[359] ,
         \A2[358] , \A2[357] , \A2[356] , \A2[355] , \A2[354] , \A2[353] ,
         \A2[352] , \A2[351] , \A2[350] , \A2[349] , \A2[348] , \A2[347] ,
         \A2[346] , \A2[345] , \A2[344] , \A2[343] , \A2[342] , \A2[341] ,
         \A2[340] , \A2[339] , \A2[338] , \A2[337] , \A2[336] , \A2[335] ,
         \A2[334] , \A2[333] , \A2[332] , \A2[331] , \A2[330] , \A2[329] ,
         \A2[328] , \A2[327] , \A2[326] , \A2[325] , \A2[324] , \A2[323] ,
         \A2[322] , \A2[321] , \A2[320] , \A2[319] , \A2[318] , \A2[317] ,
         \A2[316] , \A2[315] , \A2[314] , \A2[313] , \A2[312] , \A2[311] ,
         \A2[310] , \A2[309] , \A2[308] , \A2[307] , \A2[306] , \A2[305] ,
         \A2[304] , \A2[303] , \A2[302] , \A2[301] , \A2[300] , \A2[299] ,
         \A2[298] , \A2[297] , \A2[296] , \A2[295] , \A2[294] , \A2[293] ,
         \A2[292] , \A2[291] , \A2[290] , \A2[289] , \A2[288] , \A2[287] ,
         \A2[286] , \A2[285] , \A2[284] , \A2[283] , \A2[282] , \A2[281] ,
         \A2[280] , \A2[279] , \A2[278] , \A2[277] , \A2[276] , \A2[275] ,
         \A2[274] , \A2[273] , \A2[272] , \A2[271] , \A2[270] , \A2[269] ,
         \A2[268] , \A2[267] , \A2[266] , \A2[265] , \A2[264] , \A2[263] ,
         \A2[262] , \A2[261] , \A2[260] , \A2[259] , \A2[258] , \A2[257] ,
         \A2[256] , \A2[255] , \A2[254] , \A2[253] , \A2[252] , \A2[251] ,
         \A2[250] , \A2[249] , \A2[248] , \A2[247] , \A2[246] , \A2[245] ,
         \A2[244] , \A2[243] , \A2[242] , \A2[241] , \A2[240] , \A2[239] ,
         \A2[238] , \A2[237] , \A2[236] , \A2[235] , \A2[234] , \A2[233] ,
         \A2[232] , \A2[231] , \A2[230] , \A2[229] , \A2[228] , \A2[227] ,
         \A2[226] , \A2[225] , \A2[224] , \A2[223] , \A2[222] , \A2[221] ,
         \A2[220] , \A2[219] , \A2[218] , \A2[217] , \A2[216] , \A2[215] ,
         \A2[214] , \A2[213] , \A2[212] , \A2[211] , \A2[210] , \A2[209] ,
         \A2[208] , \A2[207] , \A2[206] , \A2[205] , \A2[204] , \A2[203] ,
         \A2[202] , \A2[201] , \A2[200] , \A2[199] , \A2[198] , \A2[197] ,
         \A2[196] , \A2[195] , \A2[194] , \A2[193] , \A2[192] , \A2[191] ,
         \A2[190] , \A2[189] , \A2[188] , \A2[187] , \A2[186] , \A2[185] ,
         \A2[184] , \A2[183] , \A2[182] , \A2[181] , \A2[180] , \A2[179] ,
         \A2[178] , \A2[177] , \A2[176] , \A2[175] , \A2[174] , \A2[173] ,
         \A2[172] , \A2[171] , \A2[170] , \A2[169] , \A2[168] , \A2[167] ,
         \A2[166] , \A2[165] , \A2[164] , \A2[163] , \A2[162] , \A2[161] ,
         \A2[160] , \A2[159] , \A2[158] , \A2[157] , \A2[156] , \A2[155] ,
         \A2[154] , \A2[153] , \A2[152] , \A2[151] , \A2[150] , \A2[149] ,
         \A2[148] , \A2[147] , \A2[146] , \A2[145] , \A2[144] , \A2[143] ,
         \A2[142] , \A2[141] , \A2[140] , \A2[139] , \A2[138] , \A2[137] ,
         \A2[136] , \A2[135] , \A2[134] , \A2[133] , \A2[132] , \A2[131] ,
         \A2[130] , \A2[129] , \A2[128] , \A2[127] , \A2[126] , \A2[125] ,
         \A2[124] , \A2[123] , \A2[122] , \A2[121] , \A2[120] , \A2[119] ,
         \A2[118] , \A2[117] , \A2[116] , \A2[115] , \A2[114] , \A2[113] ,
         \A2[112] , \A2[111] , \A2[110] , \A2[109] , \A2[108] , \A2[107] ,
         \A2[106] , \A2[105] , \A2[104] , \A2[103] , \A2[102] , \A2[101] ,
         \A2[100] , \A2[99] , \A2[98] , \A2[97] , \A2[96] , \A2[95] , \A2[94] ,
         \A2[93] , \A2[92] , \A2[91] , \A2[90] , \A2[89] , \A2[88] , \A2[87] ,
         \A2[86] , \A2[85] , \A2[84] , \A2[83] , \A2[82] , \A2[81] , \A2[80] ,
         \A2[79] , \A2[78] , \A2[77] , \A2[76] , \A2[75] , \A2[74] , \A2[73] ,
         \A2[72] , \A2[71] , \A2[70] , \A2[69] , \A2[68] , \A2[67] , \A2[66] ,
         \A2[65] , \A2[64] , \A2[63] , \A2[62] , \A2[61] , \A2[60] , \A2[59] ,
         \A2[58] , \A2[57] , \A2[56] , \A2[55] , \A2[54] , \A2[53] , \A2[52] ,
         \A2[51] , \A2[50] , \A2[49] , \A2[48] , \A2[47] , \A2[46] , \A2[45] ,
         \A2[44] , \A2[43] , \A2[42] , \A2[41] , \A2[40] , \A2[39] , \A2[38] ,
         \A2[37] , \A2[36] , \A2[35] , \A2[34] , \A2[33] , \A2[32] , \A2[31] ,
         \A2[30] , \A2[29] , \A2[28] , \A2[27] , \A2[26] , \A2[25] , \A2[24] ,
         \A2[23] , \A2[22] , \A2[21] , \A2[20] , \A2[19] , \A2[18] , \A2[17] ,
         \A2[16] , \A2[15] , \A2[14] , \A2[13] , \A2[12] , \A2[11] , \A2[10] ,
         \A2[9] , \A2[8] , \A2[7] , \A2[6] , \A2[5] , \A2[4] , \A2[3] , n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
         n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
         n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
         n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
         n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
         n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
         n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
         n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
         n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
         n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
         n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
         n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
         n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
         n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
         n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
         n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
         n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
         n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
         n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
         n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
         n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
         n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
         n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
         n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
         n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
         n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
         n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
         n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
         n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
         n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
         n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
         n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
         n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
         n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
         n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
         n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
         n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
         n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
         n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
         n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
         n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
         n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
         n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
         n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
         n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
         n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
         n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
         n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534,
         n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
         n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
         n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564,
         n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574,
         n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
         n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
         n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
         n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
         n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
         n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944,
         n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
         n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
         n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
         n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
         n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
         n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
         n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
         n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
         n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
         n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
         n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
         n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
         n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
         n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
         n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
         n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
         n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
         n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
         n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
         n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
         n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219,
         n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227,
         n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235,
         n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243,
         n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251,
         n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259,
         n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267,
         n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275,
         n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283,
         n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291,
         n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299,
         n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307,
         n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315,
         n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323,
         n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331,
         n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
         n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347,
         n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355,
         n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363,
         n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371,
         n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379,
         n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387,
         n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395,
         n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
         n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411,
         n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419,
         n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427,
         n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435,
         n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443,
         n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451,
         n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459,
         n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467,
         n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475,
         n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483,
         n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491,
         n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499,
         n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507,
         n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515,
         n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523,
         n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531,
         n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539,
         n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547,
         n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555,
         n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563,
         n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571,
         n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579,
         n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587,
         n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595,
         n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603,
         n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611,
         n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619,
         n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627,
         n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635,
         n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643,
         n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651,
         n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659,
         n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667,
         n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675,
         n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683,
         n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691,
         n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699,
         n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707,
         n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715,
         n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723,
         n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731,
         n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739,
         n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747,
         n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755,
         n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763,
         n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771,
         n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779,
         n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787,
         n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795,
         n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803,
         n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811,
         n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819,
         n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827,
         n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835,
         n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843,
         n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851,
         n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859,
         n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867,
         n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875,
         n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883,
         n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891,
         n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899,
         n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907,
         n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915,
         n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923,
         n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931,
         n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939,
         n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947,
         n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955,
         n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963,
         n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971,
         n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979,
         n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987,
         n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995,
         n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003,
         n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011,
         n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019,
         n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027,
         n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035,
         n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043,
         n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051,
         n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059,
         n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067,
         n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075,
         n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083,
         n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091,
         n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099,
         n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107,
         n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115,
         n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123,
         n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131,
         n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139,
         n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147,
         n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155,
         n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163,
         n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171,
         n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179,
         n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187,
         n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195,
         n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203,
         n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211,
         n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219,
         n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227,
         n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235,
         n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243,
         n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251,
         n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259,
         n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267,
         n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275,
         n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283,
         n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291,
         n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299,
         n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307,
         n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315,
         n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323,
         n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331,
         n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339,
         n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347,
         n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355,
         n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363,
         n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371,
         n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379,
         n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387,
         n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395,
         n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403,
         n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411,
         n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419,
         n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427,
         n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435,
         n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443,
         n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451,
         n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459,
         n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467,
         n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475,
         n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483,
         n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491,
         n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499,
         n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507,
         n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515,
         n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523,
         n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531,
         n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539,
         n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547,
         n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555,
         n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563,
         n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571,
         n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579,
         n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587,
         n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595,
         n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603,
         n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611,
         n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619,
         n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627,
         n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635,
         n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643,
         n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651,
         n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659,
         n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667,
         n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675,
         n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683,
         n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691,
         n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699,
         n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707,
         n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715,
         n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723,
         n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731,
         n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739,
         n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747,
         n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755,
         n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763,
         n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771,
         n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779,
         n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787,
         n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795,
         n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803,
         n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811,
         n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819,
         n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827,
         n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835,
         n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843,
         n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851,
         n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859,
         n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867,
         n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875,
         n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883,
         n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891,
         n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899,
         n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907,
         n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915,
         n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923,
         n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931,
         n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939,
         n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947,
         n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955,
         n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963,
         n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971,
         n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979,
         n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987,
         n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995,
         n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003,
         n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011,
         n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019,
         n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027,
         n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035,
         n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043,
         n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051,
         n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059,
         n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067,
         n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075,
         n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083,
         n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091,
         n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099,
         n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107,
         n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115,
         n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123,
         n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131,
         n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139,
         n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147,
         n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155,
         n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163,
         n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171,
         n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179,
         n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187,
         n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195,
         n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203,
         n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211,
         n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219,
         n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227,
         n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235,
         n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243,
         n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251,
         n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259,
         n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267,
         n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275,
         n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283,
         n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291,
         n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299,
         n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307,
         n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315,
         n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323,
         n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331,
         n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339,
         n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347,
         n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355,
         n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363,
         n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371,
         n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379,
         n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387,
         n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395,
         n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403,
         n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411,
         n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419,
         n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427,
         n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435,
         n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443,
         n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451,
         n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459,
         n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467,
         n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475,
         n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483,
         n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491,
         n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499,
         n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507,
         n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515,
         n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523,
         n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531,
         n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539,
         n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547,
         n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555,
         n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563,
         n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571,
         n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579,
         n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587,
         n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595,
         n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603,
         n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611,
         n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619,
         n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627,
         n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635,
         n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643,
         n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651,
         n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659,
         n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667,
         n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675,
         n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683,
         n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691,
         n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699,
         n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707,
         n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715,
         n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723,
         n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731,
         n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739,
         n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747,
         n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755,
         n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763,
         n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771,
         n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779,
         n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787,
         n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795,
         n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803,
         n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811,
         n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819,
         n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827,
         n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835,
         n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843,
         n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851,
         n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859,
         n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867,
         n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875,
         n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883,
         n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891,
         n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899,
         n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907,
         n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915,
         n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923,
         n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931,
         n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939,
         n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947,
         n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955,
         n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963,
         n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971,
         n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979,
         n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987,
         n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995,
         n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003,
         n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011,
         n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019,
         n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027,
         n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035,
         n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043,
         n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051,
         n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059,
         n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067,
         n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075,
         n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083,
         n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091,
         n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099,
         n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107,
         n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115,
         n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123,
         n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131,
         n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139,
         n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147,
         n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155,
         n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163,
         n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171,
         n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179,
         n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187,
         n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195,
         n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203,
         n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211,
         n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219,
         n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227,
         n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235,
         n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243,
         n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251,
         n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259,
         n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267,
         n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275,
         n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283,
         n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291,
         n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299,
         n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307,
         n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315,
         n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323,
         n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331,
         n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339,
         n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347,
         n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355,
         n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363,
         n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371,
         n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379,
         n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387,
         n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395,
         n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403,
         n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411,
         n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419,
         n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427,
         n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435,
         n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443,
         n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451,
         n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459,
         n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467,
         n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475,
         n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483,
         n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491,
         n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499,
         n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507,
         n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515,
         n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523,
         n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531,
         n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539,
         n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547,
         n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555,
         n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563,
         n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571,
         n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579,
         n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587,
         n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595,
         n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603,
         n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611,
         n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619,
         n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627,
         n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635,
         n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643,
         n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651,
         n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659,
         n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667,
         n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675,
         n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683,
         n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691,
         n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699,
         n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707,
         n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715,
         n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723,
         n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731,
         n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739,
         n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747,
         n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755,
         n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763,
         n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771,
         n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779,
         n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787,
         n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795,
         n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803,
         n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811,
         n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819,
         n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827,
         n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835,
         n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843,
         n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851,
         n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859,
         n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867,
         n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875,
         n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883,
         n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891,
         n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899,
         n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907,
         n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915,
         n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923,
         n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931,
         n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939,
         n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947,
         n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955,
         n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963,
         n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971,
         n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979,
         n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987,
         n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995,
         n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003,
         n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011,
         n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019,
         n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027,
         n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035,
         n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043,
         n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051,
         n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059,
         n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067,
         n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075,
         n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083,
         n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091,
         n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099,
         n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107,
         n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115,
         n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123,
         n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131,
         n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139,
         n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147,
         n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155,
         n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163,
         n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171,
         n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179,
         n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187,
         n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195,
         n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203,
         n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211,
         n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219,
         n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227,
         n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235,
         n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243,
         n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251,
         n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259,
         n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267,
         n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275,
         n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283,
         n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291,
         n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299,
         n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307,
         n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315,
         n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323,
         n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331,
         n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339,
         n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347,
         n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355,
         n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363,
         n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371,
         n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379,
         n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387,
         n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395,
         n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403,
         n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411,
         n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419,
         n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427,
         n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435,
         n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443,
         n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451,
         n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459,
         n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467,
         n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475,
         n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483,
         n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491,
         n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499,
         n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507,
         n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515,
         n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523,
         n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531,
         n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539,
         n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547,
         n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555,
         n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563,
         n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571,
         n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579,
         n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587,
         n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595,
         n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603,
         n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611,
         n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619,
         n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627,
         n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635,
         n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643,
         n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651,
         n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659,
         n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667,
         n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675,
         n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683,
         n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691,
         n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699,
         n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707,
         n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715,
         n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723,
         n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731,
         n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739,
         n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747,
         n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755,
         n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763,
         n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771,
         n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779,
         n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787,
         n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795,
         n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803,
         n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811,
         n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819,
         n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827,
         n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835,
         n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843,
         n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851,
         n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859,
         n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867,
         n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875,
         n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883,
         n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891,
         n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899,
         n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907,
         n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915,
         n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923,
         n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931,
         n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
         n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947,
         n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955,
         n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963,
         n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971,
         n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979,
         n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987,
         n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995,
         n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003,
         n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011,
         n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019,
         n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027,
         n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035,
         n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043,
         n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051,
         n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059,
         n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067,
         n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075,
         n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083,
         n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091,
         n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099,
         n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107,
         n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115,
         n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123,
         n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131,
         n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139,
         n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147,
         n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155,
         n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163,
         n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171,
         n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179,
         n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187,
         n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195,
         n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203,
         n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211,
         n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219,
         n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227,
         n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235,
         n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243,
         n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251,
         n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259,
         n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267,
         n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275,
         n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283,
         n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291,
         n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299,
         n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307,
         n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315,
         n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323,
         n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331,
         n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339,
         n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347,
         n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355,
         n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363,
         n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371,
         n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379,
         n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387,
         n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395,
         n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403,
         n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411,
         n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419,
         n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427,
         n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435,
         n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443,
         n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451,
         n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459,
         n15460, n15461, n15462, n15463, n15464, n15465, n15466, n15467,
         n15468, n15469, n15470, n15471, n15472, n15473, n15474, n15475,
         n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483,
         n15484, n15485, n15486, n15487, n15488, n15489, n15490, n15491,
         n15492, n15493, n15494, n15495, n15496, n15497, n15498, n15499,
         n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507,
         n15508, n15509, n15510, n15511, n15512, n15513, n15514, n15515,
         n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523,
         n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531,
         n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15539,
         n15540, n15541, n15542, n15543, n15544, n15545, n15546, n15547,
         n15548, n15549, n15550, n15551, n15552, n15553, n15554, n15555,
         n15556, n15557, n15558, n15559, n15560, n15561, n15562, n15563,
         n15564, n15565, n15566, n15567, n15568, n15569, n15570, n15571,
         n15572, n15573, n15574, n15575, n15576, n15577, n15578, n15579,
         n15580, n15581, n15582, n15583, n15584, n15585, n15586, n15587,
         n15588, n15589, n15590, n15591, n15592, n15593, n15594, n15595,
         n15596, n15597, n15598, n15599, n15600, n15601, n15602, n15603,
         n15604, n15605, n15606, n15607, n15608, n15609, n15610, n15611,
         n15612, n15613, n15614, n15615, n15616, n15617, n15618, n15619,
         n15620, n15621, n15622, n15623, n15624, n15625, n15626, n15627,
         n15628, n15629, n15630, n15631, n15632, n15633, n15634, n15635,
         n15636, n15637, n15638, n15639, n15640, n15641, n15642, n15643,
         n15644, n15645, n15646, n15647, n15648, n15649, n15650, n15651,
         n15652, n15653, n15654, n15655, n15656, n15657, n15658, n15659,
         n15660, n15661, n15662, n15663, n15664, n15665, n15666, n15667,
         n15668, n15669, n15670, n15671, n15672, n15673, n15674, n15675,
         n15676, n15677, n15678, n15679, n15680, n15681, n15682, n15683,
         n15684, n15685, n15686, n15687, n15688, n15689, n15690, n15691,
         n15692, n15693, n15694, n15695, n15696, n15697, n15698, n15699,
         n15700, n15701, n15702, n15703, n15704, n15705, n15706, n15707,
         n15708, n15709, n15710, n15711, n15712, n15713, n15714, n15715,
         n15716, n15717, n15718, n15719, n15720, n15721, n15722, n15723,
         n15724, n15725, n15726, n15727, n15728, n15729, n15730, n15731,
         n15732, n15733, n15734, n15735, n15736, n15737, n15738, n15739,
         n15740, n15741, n15742, n15743, n15744, n15745, n15746, n15747,
         n15748, n15749, n15750, n15751, n15752, n15753, n15754, n15755,
         n15756, n15757, n15758, n15759, n15760, n15761, n15762, n15763,
         n15764, n15765, n15766, n15767, n15768, n15769, n15770, n15771,
         n15772, n15773, n15774, n15775, n15776, n15777, n15778, n15779,
         n15780, n15781, n15782, n15783, n15784, n15785, n15786, n15787,
         n15788, n15789, n15790, n15791, n15792, n15793, n15794, n15795,
         n15796, n15797, n15798, n15799, n15800, n15801, n15802, n15803,
         n15804, n15805, n15806, n15807, n15808, n15809, n15810, n15811,
         n15812, n15813, n15814, n15815, n15816, n15817, n15818, n15819,
         n15820, n15821, n15822, n15823, n15824, n15825, n15826, n15827,
         n15828, n15829, n15830, n15831, n15832, n15833, n15834, n15835,
         n15836, n15837, n15838, n15839, n15840, n15841, n15842, n15843,
         n15844, n15845, n15846, n15847, n15848, n15849, n15850, n15851,
         n15852, n15853, n15854, n15855, n15856, n15857, n15858, n15859,
         n15860, n15861, n15862, n15863, n15864, n15865, n15866, n15867,
         n15868, n15869, n15870, n15871, n15872, n15873, n15874, n15875,
         n15876, n15877, n15878, n15879, n15880, n15881, n15882, n15883,
         n15884, n15885, n15886, n15887, n15888, n15889, n15890, n15891,
         n15892, n15893, n15894, n15895, n15896, n15897, n15898, n15899,
         n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907,
         n15908, n15909, n15910, n15911, n15912, n15913, n15914, n15915,
         n15916, n15917, n15918, n15919, n15920, n15921, n15922, n15923,
         n15924, n15925, n15926, n15927, n15928, n15929, n15930, n15931,
         n15932, n15933, n15934, n15935, n15936, n15937, n15938, n15939,
         n15940, n15941, n15942, n15943, n15944, n15945, n15946, n15947,
         n15948, n15949, n15950, n15951, n15952, n15953, n15954, n15955,
         n15956, n15957, n15958, n15959, n15960, n15961, n15962, n15963,
         n15964, n15965, n15966, n15967, n15968, n15969, n15970, n15971,
         n15972, n15973, n15974, n15975, n15976, n15977, n15978, n15979,
         n15980, n15981, n15982, n15983, n15984, n15985, n15986, n15987,
         n15988, n15989, n15990, n15991, n15992, n15993, n15994, n15995,
         n15996, n15997, n15998, n15999, n16000, n16001, n16002, n16003,
         n16004, n16005, n16006, n16007, n16008, n16009, n16010, n16011,
         n16012, n16013, n16014, n16015, n16016, n16017, n16018, n16019,
         n16020, n16021, n16022, n16023, n16024, n16025, n16026, n16027,
         n16028, n16029, n16030, n16031, n16032, n16033, n16034, n16035,
         n16036, n16037, n16038, n16039, n16040, n16041, n16042, n16043,
         n16044, n16045, n16046, n16047, n16048, n16049, n16050, n16051,
         n16052, n16053, n16054, n16055, n16056, n16057, n16058, n16059,
         n16060, n16061, n16062, n16063, n16064, n16065, n16066, n16067,
         n16068, n16069, n16070, n16071, n16072, n16073, n16074, n16075,
         n16076, n16077, n16078, n16079, n16080, n16081, n16082, n16083,
         n16084, n16085, n16086, n16087, n16088, n16089, n16090, n16091,
         n16092, n16093, n16094, n16095, n16096, n16097, n16098, n16099,
         n16100, n16101, n16102, n16103, n16104, n16105, n16106, n16107,
         n16108, n16109, n16110, n16111, n16112, n16113, n16114, n16115,
         n16116, n16117, n16118, n16119, n16120, n16121, n16122, n16123,
         n16124, n16125, n16126, n16127, n16128, n16129, n16130, n16131,
         n16132, n16133, n16134, n16135, n16136, n16137, n16138, n16139,
         n16140, n16141, n16142, n16143, n16144, n16145, n16146, n16147,
         n16148, n16149, n16150, n16151, n16152, n16153, n16154, n16155,
         n16156, n16157, n16158, n16159, n16160, n16161, n16162, n16163,
         n16164, n16165, n16166, n16167, n16168, n16169, n16170, n16171,
         n16172, n16173, n16174, n16175, n16176, n16177, n16178, n16179,
         n16180, n16181, n16182, n16183, n16184, n16185, n16186, n16187,
         n16188, n16189, n16190, n16191, n16192, n16193, n16194, n16195,
         n16196, n16197, n16198, n16199, n16200, n16201, n16202, n16203,
         n16204, n16205, n16206, n16207, n16208, n16209, n16210, n16211,
         n16212, n16213, n16214, n16215, n16216, n16217, n16218, n16219,
         n16220, n16221, n16222, n16223, n16224, n16225, n16226, n16227,
         n16228, n16229, n16230, n16231, n16232, n16233, n16234, n16235,
         n16236, n16237, n16238, n16239, n16240, n16241, n16242, n16243,
         n16244, n16245, n16246, n16247, n16248, n16249, n16250, n16251,
         n16252, n16253, n16254, n16255, n16256, n16257, n16258, n16259,
         n16260, n16261, n16262, n16263, n16264, n16265, n16266, n16267,
         n16268, n16269, n16270, n16271, n16272, n16273, n16274, n16275,
         n16276, n16277, n16278, n16279, n16280, n16281, n16282, n16283,
         n16284, n16285, n16286, n16287, n16288, n16289, n16290, n16291,
         n16292, n16293, n16294, n16295, n16296, n16297, n16298, n16299,
         n16300, n16301, n16302, n16303, n16304, n16305, n16306, n16307,
         n16308, n16309, n16310, n16311, n16312, n16313, n16314, n16315,
         n16316, n16317, n16318, n16319, n16320, n16321, n16322, n16323,
         n16324, n16325, n16326, n16327, n16328, n16329, n16330, n16331,
         n16332, n16333, n16334, n16335, n16336, n16337, n16338, n16339,
         n16340, n16341, n16342, n16343, n16344, n16345, n16346, n16347,
         n16348, n16349, n16350, n16351, n16352, n16353, n16354, n16355,
         n16356, n16357, n16358, n16359, n16360, n16361, n16362, n16363,
         n16364, n16365, n16366, n16367, n16368, n16369, n16370, n16371,
         n16372, n16373, n16374, n16375, n16376, n16377, n16378, n16379,
         n16380, n16381, n16382, n16383, n16384, n16385, n16386, n16387,
         n16388, n16389, n16390, n16391, n16392, n16393, n16394, n16395,
         n16396, n16397, n16398, n16399, n16400, n16401, n16402, n16403,
         n16404, n16405, n16406, n16407, n16408, n16409, n16410, n16411,
         n16412, n16413, n16414, n16415, n16416, n16417, n16418, n16419,
         n16420, n16421, n16422, n16423, n16424, n16425, n16426, n16427,
         n16428, n16429, n16430, n16431, n16432, n16433, n16434, n16435,
         n16436, n16437, n16438, n16439, n16440, n16441, n16442, n16443,
         n16444, n16445, n16446, n16447, n16448, n16449, n16450, n16451,
         n16452, n16453, n16454, n16455, n16456, n16457, n16458, n16459,
         n16460, n16461, n16462, n16463, n16464, n16465, n16466, n16467,
         n16468, n16469, n16470, n16471, n16472, n16473, n16474, n16475,
         n16476, n16477, n16478, n16479, n16480, n16481, n16482, n16483,
         n16484, n16485, n16486, n16487, n16488, n16489, n16490, n16491,
         n16492, n16493, n16494, n16495, n16496, n16497, n16498, n16499,
         n16500, n16501, n16502, n16503, n16504, n16505, n16506, n16507,
         n16508, n16509, n16510, n16511, n16512, n16513, n16514, n16515,
         n16516, n16517, n16518, n16519, n16520, n16521, n16522, n16523,
         n16524, n16525, n16526, n16527, n16528, n16529, n16530, n16531,
         n16532, n16533, n16534, n16535, n16536, n16537, n16538, n16539,
         n16540, n16541, n16542, n16543, n16544, n16545, n16546, n16547,
         n16548, n16549, n16550, n16551, n16552, n16553, n16554, n16555,
         n16556, n16557, n16558, n16559, n16560, n16561, n16562, n16563,
         n16564, n16565, n16566, n16567, n16568, n16569, n16570, n16571,
         n16572, n16573, n16574, n16575, n16576, n16577, n16578, n16579,
         n16580, n16581, n16582, n16583, n16584, n16585, n16586, n16587,
         n16588, n16589, n16590, n16591, n16592, n16593, n16594, n16595,
         n16596, n16597, n16598, n16599, n16600, n16601, n16602, n16603,
         n16604, n16605, n16606, n16607, n16608, n16609, n16610, n16611,
         n16612, n16613, n16614, n16615, n16616, n16617, n16618, n16619,
         n16620, n16621, n16622, n16623, n16624, n16625, n16626, n16627,
         n16628, n16629, n16630, n16631, n16632, n16633, n16634, n16635,
         n16636, n16637, n16638, n16639, n16640, n16641, n16642, n16643,
         n16644, n16645, n16646, n16647, n16648, n16649, n16650, n16651,
         n16652, n16653, n16654, n16655, n16656, n16657, n16658, n16659,
         n16660, n16661, n16662, n16663, n16664, n16665, n16666, n16667,
         n16668, n16669, n16670, n16671, n16672, n16673, n16674, n16675,
         n16676, n16677, n16678, n16679, n16680, n16681, n16682, n16683,
         n16684, n16685, n16686, n16687, n16688, n16689, n16690, n16691,
         n16692, n16693, n16694, n16695, n16696, n16697, n16698, n16699,
         n16700, n16701, n16702, n16703, n16704, n16705, n16706, n16707,
         n16708, n16709, n16710, n16711, n16712, n16713, n16714, n16715,
         n16716, n16717, n16718, n16719, n16720, n16721, n16722, n16723,
         n16724, n16725, n16726, n16727, n16728, n16729, n16730, n16731,
         n16732, n16733, n16734, n16735, n16736, n16737, n16738, n16739,
         n16740, n16741, n16742, n16743, n16744, n16745, n16746, n16747,
         n16748, n16749, n16750, n16751, n16752, n16753, n16754, n16755,
         n16756, n16757, n16758, n16759, n16760, n16761, n16762, n16763,
         n16764, n16765, n16766, n16767, n16768, n16769, n16770, n16771,
         n16772, n16773, n16774, n16775, n16776, n16777, n16778, n16779,
         n16780, n16781, n16782, n16783, n16784, n16785, n16786, n16787,
         n16788, n16789, n16790, n16791, n16792, n16793, n16794, n16795,
         n16796, n16797, n16798, n16799, n16800, n16801, n16802, n16803,
         n16804, n16805, n16806, n16807, n16808, n16809, n16810, n16811,
         n16812, n16813, n16814, n16815, n16816, n16817, n16818, n16819,
         n16820, n16821, n16822, n16823, n16824, n16825, n16826, n16827,
         n16828, n16829, n16830, n16831, n16832, n16833, n16834, n16835,
         n16836, n16837, n16838, n16839, n16840, n16841, n16842, n16843,
         n16844, n16845, n16846, n16847, n16848, n16849, n16850, n16851,
         n16852, n16853, n16854, n16855, n16856, n16857, n16858, n16859,
         n16860, n16861, n16862, n16863, n16864, n16865, n16866, n16867,
         n16868, n16869, n16870, n16871, n16872, n16873, n16874, n16875,
         n16876, n16877, n16878, n16879, n16880, n16881, n16882, n16883,
         n16884, n16885, n16886, n16887, n16888, n16889, n16890, n16891,
         n16892, n16893, n16894, n16895, n16896, n16897, n16898, n16899,
         n16900, n16901, n16902, n16903, n16904, n16905, n16906, n16907,
         n16908, n16909, n16910, n16911, n16912, n16913, n16914, n16915,
         n16916, n16917, n16918, n16919, n16920, n16921, n16922, n16923,
         n16924, n16925, n16926, n16927, n16928, n16929, n16930, n16931,
         n16932, n16933, n16934, n16935, n16936, n16937, n16938, n16939,
         n16940, n16941, n16942, n16943, n16944, n16945, n16946, n16947,
         n16948, n16949, n16950, n16951, n16952, n16953, n16954, n16955,
         n16956, n16957, n16958, n16959, n16960, n16961, n16962, n16963,
         n16964, n16965, n16966, n16967, n16968, n16969, n16970, n16971,
         n16972, n16973, n16974, n16975, n16976, n16977, n16978, n16979,
         n16980, n16981, n16982, n16983, n16984, n16985, n16986, n16987,
         n16988, n16989, n16990, n16991, n16992, n16993, n16994, n16995,
         n16996, n16997, n16998, n16999, n17000, n17001, n17002, n17003,
         n17004, n17005, n17006, n17007, n17008, n17009, n17010, n17011,
         n17012, n17013, n17014, n17015, n17016, n17017, n17018, n17019,
         n17020, n17021, n17022, n17023, n17024, n17025, n17026, n17027,
         n17028, n17029, n17030, n17031, n17032, n17033, n17034, n17035,
         n17036, n17037, n17038, n17039, n17040, n17041, n17042, n17043,
         n17044, n17045, n17046, n17047, n17048, n17049, n17050, n17051,
         n17052, n17053, n17054, n17055, n17056, n17057, n17058, n17059,
         n17060, n17061, n17062, n17063, n17064, n17065, n17066, n17067,
         n17068, n17069, n17070, n17071, n17072, n17073, n17074, n17075,
         n17076, n17077, n17078, n17079, n17080, n17081, n17082, n17083,
         n17084, n17085, n17086, n17087, n17088, n17089, n17090, n17091,
         n17092, n17093, n17094, n17095, n17096, n17097, n17098, n17099,
         n17100, n17101, n17102, n17103, n17104, n17105, n17106, n17107,
         n17108, n17109, n17110, n17111, n17112, n17113, n17114, n17115,
         n17116, n17117, n17118, n17119, n17120, n17121, n17122, n17123,
         n17124, n17125, n17126, n17127, n17128, n17129, n17130, n17131,
         n17132, n17133, n17134, n17135, n17136, n17137, n17138, n17139,
         n17140, n17141, n17142, n17143, n17144, n17145, n17146, n17147,
         n17148, n17149, n17150, n17151, n17152, n17153, n17154, n17155,
         n17156, n17157, n17158, n17159, n17160, n17161, n17162, n17163,
         n17164, n17165, n17166, n17167, n17168, n17169, n17170, n17171,
         n17172, n17173, n17174, n17175, n17176, n17177, n17178, n17179,
         n17180, n17181, n17182, n17183, n17184, n17185, n17186, n17187,
         n17188, n17189, n17190, n17191, n17192, n17193, n17194, n17195,
         n17196, n17197, n17198, n17199, n17200, n17201, n17202, n17203,
         n17204, n17205, n17206, n17207, n17208, n17209, n17210, n17211,
         n17212, n17213, n17214, n17215, n17216, n17217, n17218, n17219,
         n17220, n17221, n17222, n17223, n17224, n17225, n17226, n17227,
         n17228, n17229, n17230, n17231, n17232, n17233, n17234, n17235,
         n17236, n17237, n17238, n17239, n17240, n17241, n17242, n17243,
         n17244, n17245, n17246, n17247, n17248, n17249, n17250, n17251,
         n17252, n17253, n17254, n17255, n17256, n17257, n17258, n17259,
         n17260, n17261, n17262, n17263, n17264, n17265, n17266, n17267,
         n17268, n17269, n17270, n17271, n17272, n17273, n17274, n17275,
         n17276, n17277, n17278, n17279, n17280, n17281, n17282, n17283,
         n17284, n17285, n17286, n17287, n17288, n17289, n17290, n17291,
         n17292, n17293, n17294, n17295, n17296, n17297, n17298, n17299,
         n17300, n17301, n17302, n17303, n17304, n17305, n17306, n17307,
         n17308, n17309, n17310, n17311, n17312, n17313, n17314, n17315,
         n17316, n17317, n17318, n17319, n17320, n17321, n17322, n17323,
         n17324, n17325, n17326, n17327, n17328, n17329, n17330, n17331,
         n17332, n17333, n17334, n17335, n17336, n17337, n17338, n17339,
         n17340, n17341, n17342, n17343, n17344, n17345, n17346, n17347,
         n17348, n17349, n17350, n17351, n17352, n17353, n17354, n17355,
         n17356, n17357, n17358, n17359, n17360, n17361, n17362, n17363,
         n17364, n17365, n17366, n17367, n17368, n17369, n17370, n17371,
         n17372, n17373, n17374, n17375, n17376, n17377, n17378, n17379,
         n17380, n17381, n17382, n17383, n17384, n17385, n17386, n17387,
         n17388, n17389, n17390, n17391, n17392, n17393, n17394, n17395,
         n17396, n17397, n17398, n17399, n17400, n17401, n17402, n17403,
         n17404, n17405, n17406, n17407, n17408, n17409, n17410, n17411,
         n17412, n17413, n17414, n17415, n17416, n17417, n17418, n17419,
         n17420, n17421, n17422, n17423, n17424, n17425, n17426, n17427,
         n17428, n17429, n17430, n17431, n17432, n17433, n17434, n17435,
         n17436, n17437, n17438, n17439, n17440, n17441, n17442, n17443,
         n17444, n17445, n17446, n17447, n17448, n17449, n17450, n17451,
         n17452, n17453, n17454, n17455, n17456, n17457, n17458, n17459,
         n17460, n17461, n17462, n17463, n17464, n17465, n17466, n17467,
         n17468, n17469, n17470, n17471, n17472, n17473, n17474, n17475,
         n17476, n17477, n17478, n17479, n17480, n17481, n17482, n17483,
         n17484, n17485, n17486, n17487, n17488, n17489, n17490, n17491,
         n17492, n17493, n17494, n17495, n17496, n17497, n17498, n17499,
         n17500, n17501, n17502, n17503, n17504, n17505, n17506, n17507,
         n17508, n17509, n17510, n17511, n17512, n17513, n17514, n17515,
         n17516, n17517, n17518, n17519, n17520, n17521, n17522, n17523,
         n17524, n17525, n17526, n17527, n17528, n17529, n17530, n17531,
         n17532, n17533, n17534, n17535, n17536, n17537, n17538, n17539,
         n17540, n17541, n17542, n17543, n17544, n17545, n17546, n17547,
         n17548, n17549, n17550, n17551, n17552, n17553, n17554, n17555,
         n17556, n17557, n17558, n17559, n17560, n17561, n17562, n17563,
         n17564, n17565, n17566, n17567, n17568, n17569, n17570, n17571,
         n17572, n17573, n17574, n17575, n17576, n17577, n17578, n17579,
         n17580, n17581, n17582, n17583, n17584, n17585, n17586, n17587,
         n17588, n17589, n17590, n17591, n17592, n17593, n17594, n17595,
         n17596, n17597, n17598, n17599, n17600, n17601, n17602, n17603,
         n17604, n17605, n17606, n17607, n17608, n17609, n17610, n17611,
         n17612, n17613, n17614, n17615, n17616, n17617, n17618, n17619,
         n17620, n17621, n17622, n17623, n17624, n17625, n17626, n17627,
         n17628, n17629, n17630, n17631, n17632, n17633, n17634, n17635,
         n17636, n17637, n17638, n17639, n17640, n17641, n17642, n17643,
         n17644, n17645, n17646, n17647, n17648, n17649, n17650, n17651,
         n17652, n17653, n17654, n17655, n17656, n17657, n17658, n17659,
         n17660, n17661, n17662, n17663, n17664, n17665, n17666, n17667,
         n17668, n17669, n17670, n17671, n17672, n17673, n17674, n17675,
         n17676, n17677, n17678, n17679, n17680, n17681, n17682, n17683,
         n17684, n17685, n17686, n17687, n17688, n17689, n17690, n17691,
         n17692, n17693, n17694, n17695, n17696, n17697, n17698, n17699,
         n17700, n17701, n17702, n17703, n17704, n17705, n17706, n17707,
         n17708, n17709, n17710, n17711, n17712, n17713, n17714, n17715,
         n17716, n17717, n17718, n17719, n17720, n17721, n17722, n17723,
         n17724, n17725, n17726, n17727, n17728, n17729, n17730, n17731,
         n17732, n17733, n17734, n17735, n17736, n17737, n17738, n17739,
         n17740, n17741, n17742, n17743, n17744, n17745, n17746, n17747,
         n17748, n17749, n17750, n17751, n17752, n17753, n17754, n17755,
         n17756, n17757, n17758, n17759, n17760, n17761, n17762, n17763,
         n17764, n17765, n17766, n17767, n17768, n17769, n17770, n17771,
         n17772, n17773, n17774, n17775, n17776, n17777, n17778, n17779,
         n17780, n17781, n17782, n17783, n17784, n17785, n17786, n17787,
         n17788, n17789, n17790, n17791, n17792, n17793, n17794, n17795,
         n17796, n17797, n17798, n17799, n17800, n17801, n17802, n17803,
         n17804, n17805, n17806, n17807, n17808, n17809, n17810, n17811,
         n17812, n17813, n17814, n17815, n17816, n17817, n17818, n17819,
         n17820, n17821, n17822, n17823, n17824, n17825, n17826, n17827,
         n17828, n17829, n17830, n17831, n17832, n17833, n17834, n17835,
         n17836, n17837, n17838, n17839, n17840, n17841, n17842, n17843,
         n17844, n17845, n17846, n17847, n17848, n17849, n17850, n17851,
         n17852, n17853, n17854, n17855, n17856, n17857, n17858, n17859,
         n17860, n17861, n17862, n17863, n17864, n17865, n17866, n17867,
         n17868, n17869, n17870, n17871, n17872, n17873, n17874, n17875,
         n17876, n17877, n17878, n17879, n17880, n17881, n17882, n17883,
         n17884, n17885, n17886, n17887, n17888, n17889, n17890, n17891,
         n17892, n17893, n17894, n17895, n17896, n17897, n17898, n17899,
         n17900, n17901, n17902, n17903, n17904, n17905, n17906, n17907,
         n17908, n17909, n17910, n17911, n17912, n17913, n17914, n17915,
         n17916, n17917, n17918, n17919, n17920, n17921, n17922, n17923,
         n17924, n17925, n17926, n17927, n17928, n17929, n17930, n17931,
         n17932, n17933, n17934, n17935, n17936, n17937, n17938, n17939,
         n17940, n17941, n17942, n17943, n17944, n17945, n17946, n17947,
         n17948, n17949, n17950, n17951, n17952, n17953, n17954, n17955,
         n17956, n17957, n17958, n17959, n17960, n17961, n17962, n17963,
         n17964, n17965, n17966, n17967, n17968, n17969, n17970, n17971,
         n17972, n17973, n17974, n17975, n17976, n17977, n17978, n17979,
         n17980, n17981, n17982, n17983, n17984, n17985, n17986, n17987,
         n17988, n17989, n17990, n17991, n17992, n17993, n17994, n17995,
         n17996, n17997, n17998, n17999, n18000, n18001, n18002, n18003,
         n18004, n18005, n18006, n18007, n18008, n18009, n18010, n18011,
         n18012, n18013, n18014, n18015, n18016, n18017, n18018, n18019,
         n18020, n18021, n18022, n18023, n18024, n18025, n18026, n18027,
         n18028, n18029, n18030, n18031, n18032, n18033, n18034, n18035,
         n18036, n18037, n18038, n18039, n18040, n18041, n18042, n18043,
         n18044, n18045, n18046, n18047, n18048, n18049, n18050, n18051,
         n18052, n18053, n18054, n18055, n18056, n18057, n18058, n18059,
         n18060, n18061, n18062, n18063, n18064, n18065, n18066, n18067,
         n18068, n18069, n18070, n18071, n18072, n18073, n18074, n18075,
         n18076, n18077, n18078, n18079, n18080, n18081, n18082, n18083,
         n18084, n18085, n18086, n18087, n18088, n18089, n18090, n18091,
         n18092, n18093, n18094, n18095, n18096, n18097, n18098, n18099,
         n18100, n18101, n18102, n18103, n18104, n18105, n18106, n18107,
         n18108, n18109, n18110, n18111, n18112, n18113, n18114, n18115,
         n18116, n18117, n18118, n18119, n18120, n18121, n18122, n18123,
         n18124, n18125, n18126, n18127, n18128, n18129, n18130, n18131,
         n18132, n18133, n18134, n18135, n18136, n18137, n18138, n18139,
         n18140, n18141, n18142, n18143, n18144, n18145, n18146, n18147,
         n18148, n18149, n18150, n18151, n18152, n18153, n18154, n18155,
         n18156, n18157, n18158, n18159, n18160, n18161, n18162, n18163,
         n18164, n18165, n18166, n18167, n18168, n18169, n18170, n18171,
         n18172, n18173, n18174, n18175, n18176, n18177, n18178, n18179,
         n18180, n18181, n18182, n18183, n18184, n18185, n18186, n18187,
         n18188, n18189, n18190, n18191, n18192, n18193, n18194, n18195,
         n18196, n18197, n18198, n18199, n18200, n18201, n18202, n18203,
         n18204, n18205, n18206, n18207, n18208, n18209, n18210, n18211,
         n18212, n18213, n18214, n18215, n18216, n18217, n18218, n18219,
         n18220, n18221, n18222, n18223, n18224, n18225, n18226, n18227,
         n18228, n18229, n18230, n18231, n18232, n18233, n18234, n18235,
         n18236, n18237, n18238, n18239, n18240, n18241, n18242, n18243,
         n18244, n18245, n18246, n18247, n18248, n18249, n18250, n18251,
         n18252, n18253, n18254, n18255, n18256, n18257, n18258, n18259,
         n18260, n18261, n18262, n18263, n18264, n18265, n18266, n18267,
         n18268, n18269, n18270, n18271, n18272, n18273, n18274, n18275,
         n18276, n18277, n18278, n18279, n18280, n18281, n18282, n18283,
         n18284, n18285, n18286, n18287, n18288, n18289, n18290, n18291,
         n18292, n18293, n18294, n18295, n18296, n18297, n18298, n18299,
         n18300, n18301, n18302, n18303, n18304, n18305, n18306, n18307,
         n18308, n18309, n18310, n18311, n18312, n18313, n18314, n18315,
         n18316, n18317, n18318, n18319, n18320, n18321, n18322, n18323,
         n18324, n18325, n18326, n18327, n18328, n18329, n18330, n18331,
         n18332, n18333, n18334, n18335, n18336, n18337, n18338, n18339,
         n18340, n18341, n18342, n18343, n18344, n18345, n18346, n18347,
         n18348, n18349, n18350, n18351, n18352, n18353, n18354, n18355,
         n18356, n18357, n18358, n18359, n18360, n18361, n18362, n18363,
         n18364, n18365, n18366, n18367, n18368, n18369, n18370, n18371,
         n18372, n18373, n18374, n18375, n18376, n18377, n18378, n18379,
         n18380, n18381, n18382, n18383, n18384, n18385, n18386, n18387,
         n18388, n18389, n18390, n18391, n18392, n18393, n18394, n18395,
         n18396, n18397, n18398, n18399, n18400, n18401, n18402, n18403,
         n18404, n18405, n18406, n18407, n18408, n18409, n18410, n18411,
         n18412, n18413, n18414, n18415, n18416, n18417, n18418, n18419,
         n18420, n18421, n18422, n18423, n18424, n18425, n18426, n18427,
         n18428, n18429, n18430, n18431, n18432, n18433, n18434, n18435,
         n18436, n18437, n18438, n18439, n18440, n18441, n18442, n18443,
         n18444, n18445, n18446, n18447, n18448, n18449, n18450, n18451,
         n18452, n18453, n18454, n18455, n18456, n18457, n18458, n18459,
         n18460, n18461, n18462, n18463, n18464, n18465, n18466, n18467,
         n18468, n18469, n18470, n18471, n18472, n18473, n18474, n18475,
         n18476, n18477, n18478, n18479, n18480, n18481, n18482, n18483,
         n18484, n18485, n18486, n18487, n18488, n18489, n18490, n18491,
         n18492, n18493, n18494, n18495, n18496, n18497, n18498, n18499,
         n18500, n18501, n18502, n18503, n18504, n18505, n18506, n18507,
         n18508, n18509, n18510, n18511, n18512, n18513, n18514, n18515,
         n18516, n18517, n18518, n18519, n18520, n18521, n18522, n18523,
         n18524, n18525, n18526, n18527, n18528, n18529, n18530, n18531,
         n18532, n18533, n18534, n18535, n18536, n18537, n18538, n18539,
         n18540, n18541, n18542, n18543, n18544, n18545, n18546, n18547,
         n18548, n18549, n18550, n18551, n18552, n18553, n18554, n18555,
         n18556, n18557, n18558, n18559, n18560, n18561, n18562, n18563,
         n18564, n18565, n18566, n18567, n18568, n18569, n18570, n18571,
         n18572, n18573, n18574, n18575, n18576, n18577, n18578, n18579,
         n18580, n18581, n18582, n18583, n18584, n18585, n18586, n18587,
         n18588, n18589, n18590, n18591, n18592, n18593, n18594, n18595,
         n18596, n18597, n18598, n18599, n18600, n18601, n18602, n18603,
         n18604, n18605, n18606, n18607, n18608, n18609, n18610, n18611,
         n18612, n18613, n18614, n18615, n18616, n18617, n18618, n18619,
         n18620, n18621, n18622, n18623, n18624, n18625, n18626, n18627,
         n18628, n18629, n18630, n18631, n18632, n18633, n18634, n18635,
         n18636, n18637, n18638, n18639, n18640, n18641, n18642, n18643,
         n18644, n18645, n18646, n18647, n18648, n18649, n18650, n18651,
         n18652, n18653, n18654, n18655, n18656, n18657, n18658, n18659,
         n18660, n18661, n18662, n18663, n18664, n18665, n18666, n18667,
         n18668, n18669, n18670, n18671, n18672, n18673, n18674, n18675,
         n18676, n18677, n18678, n18679, n18680, n18681, n18682, n18683,
         n18684, n18685, n18686, n18687, n18688, n18689, n18690, n18691,
         n18692, n18693, n18694, n18695, n18696, n18697, n18698, n18699,
         n18700, n18701, n18702, n18703, n18704, n18705, n18706, n18707,
         n18708, n18709, n18710, n18711, n18712, n18713, n18714, n18715,
         n18716, n18717, n18718, n18719, n18720, n18721, n18722, n18723,
         n18724, n18725, n18726, n18727, n18728, n18729, n18730, n18731,
         n18732, n18733, n18734, n18735, n18736, n18737, n18738, n18739,
         n18740, n18741, n18742, n18743, n18744, n18745, n18746, n18747,
         n18748, n18749, n18750, n18751, n18752, n18753, n18754, n18755,
         n18756, n18757, n18758, n18759, n18760, n18761, n18762, n18763,
         n18764, n18765, n18766, n18767, n18768, n18769, n18770, n18771,
         n18772, n18773, n18774, n18775, n18776, n18777, n18778, n18779,
         n18780, n18781, n18782, n18783, n18784, n18785, n18786, n18787,
         n18788, n18789, n18790, n18791, n18792, n18793, n18794, n18795,
         n18796, n18797, n18798, n18799, n18800, n18801, n18802, n18803,
         n18804, n18805, n18806, n18807, n18808, n18809, n18810, n18811,
         n18812, n18813, n18814, n18815, n18816, n18817, n18818, n18819,
         n18820, n18821, n18822, n18823, n18824, n18825, n18826, n18827,
         n18828, n18829, n18830, n18831, n18832, n18833, n18834, n18835,
         n18836, n18837, n18838, n18839, n18840, n18841, n18842, n18843,
         n18844, n18845, n18846, n18847, n18848, n18849, n18850, n18851,
         n18852, n18853, n18854, n18855, n18856, n18857, n18858, n18859,
         n18860, n18861, n18862, n18863, n18864, n18865, n18866, n18867,
         n18868, n18869, n18870, n18871, n18872, n18873, n18874, n18875,
         n18876, n18877, n18878, n18879, n18880, n18881, n18882, n18883,
         n18884, n18885, n18886, n18887, n18888, n18889, n18890, n18891,
         n18892, n18893, n18894, n18895, n18896, n18897, n18898, n18899,
         n18900, n18901, n18902, n18903, n18904, n18905, n18906, n18907,
         n18908, n18909, n18910, n18911, n18912, n18913, n18914, n18915,
         n18916, n18917, n18918, n18919, n18920, n18921, n18922, n18923,
         n18924, n18925, n18926, n18927, n18928, n18929, n18930, n18931,
         n18932, n18933, n18934, n18935, n18936, n18937, n18938, n18939,
         n18940, n18941, n18942, n18943, n18944, n18945, n18946, n18947,
         n18948, n18949, n18950, n18951, n18952, n18953, n18954, n18955,
         n18956, n18957, n18958, n18959, n18960, n18961, n18962, n18963,
         n18964, n18965, n18966, n18967, n18968, n18969, n18970, n18971,
         n18972, n18973, n18974, n18975, n18976, n18977, n18978, n18979,
         n18980, n18981, n18982, n18983, n18984, n18985, n18986, n18987,
         n18988, n18989, n18990, n18991, n18992, n18993, n18994, n18995,
         n18996, n18997, n18998, n18999, n19000, n19001, n19002, n19003,
         n19004, n19005, n19006, n19007, n19008, n19009, n19010, n19011,
         n19012, n19013, n19014, n19015, n19016, n19017, n19018, n19019,
         n19020, n19021, n19022, n19023, n19024, n19025, n19026, n19027,
         n19028, n19029, n19030, n19031, n19032, n19033, n19034, n19035,
         n19036, n19037, n19038, n19039, n19040, n19041, n19042, n19043,
         n19044, n19045, n19046, n19047, n19048, n19049, n19050, n19051,
         n19052, n19053, n19054, n19055, n19056, n19057, n19058, n19059,
         n19060, n19061, n19062, n19063, n19064, n19065, n19066, n19067,
         n19068, n19069, n19070, n19071, n19072, n19073, n19074, n19075,
         n19076, n19077, n19078, n19079, n19080, n19081, n19082, n19083,
         n19084, n19085, n19086, n19087, n19088, n19089, n19090, n19091,
         n19092, n19093, n19094, n19095, n19096, n19097, n19098, n19099,
         n19100, n19101, n19102, n19103, n19104, n19105, n19106, n19107,
         n19108, n19109, n19110, n19111, n19112, n19113, n19114, n19115,
         n19116, n19117, n19118, n19119, n19120, n19121, n19122, n19123,
         n19124, n19125, n19126, n19127, n19128, n19129, n19130, n19131,
         n19132, n19133, n19134, n19135, n19136, n19137, n19138, n19139,
         n19140, n19141, n19142, n19143, n19144, n19145, n19146, n19147,
         n19148, n19149, n19150, n19151, n19152, n19153, n19154, n19155,
         n19156, n19157, n19158, n19159, n19160, n19161, n19162, n19163,
         n19164, n19165, n19166, n19167, n19168, n19169, n19170, n19171,
         n19172, n19173, n19174, n19175, n19176, n19177, n19178, n19179,
         n19180, n19181, n19182, n19183, n19184, n19185, n19186, n19187,
         n19188, n19189, n19190, n19191, n19192, n19193, n19194, n19195,
         n19196, n19197, n19198, n19199, n19200, n19201, n19202, n19203,
         n19204, n19205, n19206, n19207, n19208, n19209, n19210, n19211,
         n19212, n19213, n19214, n19215, n19216, n19217, n19218, n19219,
         n19220, n19221, n19222, n19223, n19224, n19225, n19226, n19227,
         n19228, n19229, n19230, n19231, n19232, n19233, n19234, n19235,
         n19236, n19237, n19238, n19239, n19240, n19241, n19242, n19243,
         n19244, n19245, n19246, n19247, n19248, n19249, n19250, n19251,
         n19252, n19253, n19254, n19255, n19256, n19257, n19258, n19259,
         n19260, n19261, n19262, n19263, n19264, n19265, n19266, n19267,
         n19268, n19269, n19270, n19271, n19272, n19273, n19274, n19275,
         n19276, n19277, n19278, n19279, n19280, n19281, n19282, n19283,
         n19284, n19285, n19286, n19287, n19288, n19289, n19290, n19291,
         n19292, n19293, n19294, n19295, n19296, n19297, n19298, n19299,
         n19300, n19301, n19302, n19303, n19304, n19305, n19306, n19307,
         n19308, n19309, n19310, n19311, n19312, n19313, n19314, n19315,
         n19316, n19317, n19318, n19319, n19320, n19321, n19322, n19323,
         n19324, n19325, n19326, n19327, n19328, n19329, n19330, n19331,
         n19332, n19333, n19334, n19335, n19336, n19337, n19338, n19339,
         n19340, n19341, n19342, n19343, n19344, n19345, n19346, n19347,
         n19348, n19349, n19350, n19351, n19352, n19353, n19354, n19355,
         n19356, n19357, n19358, n19359, n19360, n19361, n19362, n19363,
         n19364, n19365, n19366, n19367, n19368, n19369, n19370, n19371,
         n19372, n19373, n19374, n19375, n19376, n19377, n19378, n19379,
         n19380, n19381, n19382, n19383, n19384, n19385, n19386, n19387,
         n19388, n19389, n19390, n19391, n19392, n19393, n19394, n19395,
         n19396, n19397, n19398, n19399, n19400, n19401, n19402, n19403,
         n19404, n19405, n19406, n19407, n19408, n19409, n19410, n19411,
         n19412, n19413, n19414, n19415, n19416, n19417, n19418, n19419,
         n19420, n19421, n19422, n19423, n19424, n19425, n19426, n19427,
         n19428, n19429, n19430, n19431, n19432, n19433, n19434, n19435,
         n19436, n19437, n19438, n19439, n19440, n19441, n19442, n19443,
         n19444, n19445, n19446, n19447, n19448, n19449, n19450, n19451,
         n19452, n19453, n19454, n19455, n19456, n19457, n19458, n19459,
         n19460, n19461;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;

  mult_N1024_CC256_DW01_add_0 FS_1 ( .A({1'b0, \A1[1024] , \A1[1023] , 
        \A1[1022] , \A1[1021] , \A1[1020] , \A1[1019] , \A1[1018] , \A1[1017] , 
        \A1[1016] , \A1[1015] , \A1[1014] , \A1[1013] , \A1[1012] , \A1[1011] , 
        \A1[1010] , \A1[1009] , \A1[1008] , \A1[1007] , \A1[1006] , \A1[1005] , 
        \A1[1004] , \A1[1003] , \A1[1002] , \A1[1001] , \A1[1000] , \A1[999] , 
        \A1[998] , \A1[997] , \A1[996] , \A1[995] , \A1[994] , \A1[993] , 
        \A1[992] , \A1[991] , \A1[990] , \A1[989] , \A1[988] , \A1[987] , 
        \A1[986] , \A1[985] , \A1[984] , \A1[983] , \A1[982] , \A1[981] , 
        \A1[980] , \A1[979] , \A1[978] , \A1[977] , \A1[976] , \A1[975] , 
        \A1[974] , \A1[973] , \A1[972] , \A1[971] , \A1[970] , \A1[969] , 
        \A1[968] , \A1[967] , \A1[966] , \A1[965] , \A1[964] , \A1[963] , 
        \A1[962] , \A1[961] , \A1[960] , \A1[959] , \A1[958] , \A1[957] , 
        \A1[956] , \A1[955] , \A1[954] , \A1[953] , \A1[952] , \A1[951] , 
        \A1[950] , \A1[949] , \A1[948] , \A1[947] , \A1[946] , \A1[945] , 
        \A1[944] , \A1[943] , \A1[942] , \A1[941] , \A1[940] , \A1[939] , 
        \A1[938] , \A1[937] , \A1[936] , \A1[935] , \A1[934] , \A1[933] , 
        \A1[932] , \A1[931] , \A1[930] , \A1[929] , \A1[928] , \A1[927] , 
        \A1[926] , \A1[925] , \A1[924] , \A1[923] , \A1[922] , \A1[921] , 
        \A1[920] , \A1[919] , \A1[918] , \A1[917] , \A1[916] , \A1[915] , 
        \A1[914] , \A1[913] , \A1[912] , \A1[911] , \A1[910] , \A1[909] , 
        \A1[908] , \A1[907] , \A1[906] , \A1[905] , \A1[904] , \A1[903] , 
        \A1[902] , \A1[901] , \A1[900] , \A1[899] , \A1[898] , \A1[897] , 
        \A1[896] , \A1[895] , \A1[894] , \A1[893] , \A1[892] , \A1[891] , 
        \A1[890] , \A1[889] , \A1[888] , \A1[887] , \A1[886] , \A1[885] , 
        \A1[884] , \A1[883] , \A1[882] , \A1[881] , \A1[880] , \A1[879] , 
        \A1[878] , \A1[877] , \A1[876] , \A1[875] , \A1[874] , \A1[873] , 
        \A1[872] , \A1[871] , \A1[870] , \A1[869] , \A1[868] , \A1[867] , 
        \A1[866] , \A1[865] , \A1[864] , \A1[863] , \A1[862] , \A1[861] , 
        \A1[860] , \A1[859] , \A1[858] , \A1[857] , \A1[856] , \A1[855] , 
        \A1[854] , \A1[853] , \A1[852] , \A1[851] , \A1[850] , \A1[849] , 
        \A1[848] , \A1[847] , \A1[846] , \A1[845] , \A1[844] , \A1[843] , 
        \A1[842] , \A1[841] , \A1[840] , \A1[839] , \A1[838] , \A1[837] , 
        \A1[836] , \A1[835] , \A1[834] , \A1[833] , \A1[832] , \A1[831] , 
        \A1[830] , \A1[829] , \A1[828] , \A1[827] , \A1[826] , \A1[825] , 
        \A1[824] , \A1[823] , \A1[822] , \A1[821] , \A1[820] , \A1[819] , 
        \A1[818] , \A1[817] , \A1[816] , \A1[815] , \A1[814] , \A1[813] , 
        \A1[812] , \A1[811] , \A1[810] , \A1[809] , \A1[808] , \A1[807] , 
        \A1[806] , \A1[805] , \A1[804] , \A1[803] , \A1[802] , \A1[801] , 
        \A1[800] , \A1[799] , \A1[798] , \A1[797] , \A1[796] , \A1[795] , 
        \A1[794] , \A1[793] , \A1[792] , \A1[791] , \A1[790] , \A1[789] , 
        \A1[788] , \A1[787] , \A1[786] , \A1[785] , \A1[784] , \A1[783] , 
        \A1[782] , \A1[781] , \A1[780] , \A1[779] , \A1[778] , \A1[777] , 
        \A1[776] , \A1[775] , \A1[774] , \A1[773] , \A1[772] , \A1[771] , 
        \A1[770] , \A1[769] , \A1[768] , \A1[767] , \A1[766] , \A1[765] , 
        \A1[764] , \A1[763] , \A1[762] , \A1[761] , \A1[760] , \A1[759] , 
        \A1[758] , \A1[757] , \A1[756] , \A1[755] , \A1[754] , \A1[753] , 
        \A1[752] , \A1[751] , \A1[750] , \A1[749] , \A1[748] , \A1[747] , 
        \A1[746] , \A1[745] , \A1[744] , \A1[743] , \A1[742] , \A1[741] , 
        \A1[740] , \A1[739] , \A1[738] , \A1[737] , \A1[736] , \A1[735] , 
        \A1[734] , \A1[733] , \A1[732] , \A1[731] , \A1[730] , \A1[729] , 
        \A1[728] , \A1[727] , \A1[726] , \A1[725] , \A1[724] , \A1[723] , 
        \A1[722] , \A1[721] , \A1[720] , \A1[719] , \A1[718] , \A1[717] , 
        \A1[716] , \A1[715] , \A1[714] , \A1[713] , \A1[712] , \A1[711] , 
        \A1[710] , \A1[709] , \A1[708] , \A1[707] , \A1[706] , \A1[705] , 
        \A1[704] , \A1[703] , \A1[702] , \A1[701] , \A1[700] , \A1[699] , 
        \A1[698] , \A1[697] , \A1[696] , \A1[695] , \A1[694] , \A1[693] , 
        \A1[692] , \A1[691] , \A1[690] , \A1[689] , \A1[688] , \A1[687] , 
        \A1[686] , \A1[685] , \A1[684] , \A1[683] , \A1[682] , \A1[681] , 
        \A1[680] , \A1[679] , \A1[678] , \A1[677] , \A1[676] , \A1[675] , 
        \A1[674] , \A1[673] , \A1[672] , \A1[671] , \A1[670] , \A1[669] , 
        \A1[668] , \A1[667] , \A1[666] , \A1[665] , \A1[664] , \A1[663] , 
        \A1[662] , \A1[661] , \A1[660] , \A1[659] , \A1[658] , \A1[657] , 
        \A1[656] , \A1[655] , \A1[654] , \A1[653] , \A1[652] , \A1[651] , 
        \A1[650] , \A1[649] , \A1[648] , \A1[647] , \A1[646] , \A1[645] , 
        \A1[644] , \A1[643] , \A1[642] , \A1[641] , \A1[640] , \A1[639] , 
        \A1[638] , \A1[637] , \A1[636] , \A1[635] , \A1[634] , \A1[633] , 
        \A1[632] , \A1[631] , \A1[630] , \A1[629] , \A1[628] , \A1[627] , 
        \A1[626] , \A1[625] , \A1[624] , \A1[623] , \A1[622] , \A1[621] , 
        \A1[620] , \A1[619] , \A1[618] , \A1[617] , \A1[616] , \A1[615] , 
        \A1[614] , \A1[613] , \A1[612] , \A1[611] , \A1[610] , \A1[609] , 
        \A1[608] , \A1[607] , \A1[606] , \A1[605] , \A1[604] , \A1[603] , 
        \A1[602] , \A1[601] , \A1[600] , \A1[599] , \A1[598] , \A1[597] , 
        \A1[596] , \A1[595] , \A1[594] , \A1[593] , \A1[592] , \A1[591] , 
        \A1[590] , \A1[589] , \A1[588] , \A1[587] , \A1[586] , \A1[585] , 
        \A1[584] , \A1[583] , \A1[582] , \A1[581] , \A1[580] , \A1[579] , 
        \A1[578] , \A1[577] , \A1[576] , \A1[575] , \A1[574] , \A1[573] , 
        \A1[572] , \A1[571] , \A1[570] , \A1[569] , \A1[568] , \A1[567] , 
        \A1[566] , \A1[565] , \A1[564] , \A1[563] , \A1[562] , \A1[561] , 
        \A1[560] , \A1[559] , \A1[558] , \A1[557] , \A1[556] , \A1[555] , 
        \A1[554] , \A1[553] , \A1[552] , \A1[551] , \A1[550] , \A1[549] , 
        \A1[548] , \A1[547] , \A1[546] , \A1[545] , \A1[544] , \A1[543] , 
        \A1[542] , \A1[541] , \A1[540] , \A1[539] , \A1[538] , \A1[537] , 
        \A1[536] , \A1[535] , \A1[534] , \A1[533] , \A1[532] , \A1[531] , 
        \A1[530] , \A1[529] , \A1[528] , \A1[527] , \A1[526] , \A1[525] , 
        \A1[524] , \A1[523] , \A1[522] , \A1[521] , \A1[520] , \A1[519] , 
        \A1[518] , \A1[517] , \A1[516] , \A1[515] , \A1[514] , \A1[513] , 
        \A1[512] , \A1[511] , \A1[510] , \A1[509] , \A1[508] , \A1[507] , 
        \A1[506] , \A1[505] , \A1[504] , \A1[503] , \A1[502] , \A1[501] , 
        \A1[500] , \A1[499] , \A1[498] , \A1[497] , \A1[496] , \A1[495] , 
        \A1[494] , \A1[493] , \A1[492] , \A1[491] , \A1[490] , \A1[489] , 
        \A1[488] , \A1[487] , \A1[486] , \A1[485] , \A1[484] , \A1[483] , 
        \A1[482] , \A1[481] , \A1[480] , \A1[479] , \A1[478] , \A1[477] , 
        \A1[476] , \A1[475] , \A1[474] , \A1[473] , \A1[472] , \A1[471] , 
        \A1[470] , \A1[469] , \A1[468] , \A1[467] , \A1[466] , \A1[465] , 
        \A1[464] , \A1[463] , \A1[462] , \A1[461] , \A1[460] , \A1[459] , 
        \A1[458] , \A1[457] , \A1[456] , \A1[455] , \A1[454] , \A1[453] , 
        \A1[452] , \A1[451] , \A1[450] , \A1[449] , \A1[448] , \A1[447] , 
        \A1[446] , \A1[445] , \A1[444] , \A1[443] , \A1[442] , \A1[441] , 
        \A1[440] , \A1[439] , \A1[438] , \A1[437] , \A1[436] , \A1[435] , 
        \A1[434] , \A1[433] , \A1[432] , \A1[431] , \A1[430] , \A1[429] , 
        \A1[428] , \A1[427] , \A1[426] , \A1[425] , \A1[424] , \A1[423] , 
        \A1[422] , \A1[421] , \A1[420] , \A1[419] , \A1[418] , \A1[417] , 
        \A1[416] , \A1[415] , \A1[414] , \A1[413] , \A1[412] , \A1[411] , 
        \A1[410] , \A1[409] , \A1[408] , \A1[407] , \A1[406] , \A1[405] , 
        \A1[404] , \A1[403] , \A1[402] , \A1[401] , \A1[400] , \A1[399] , 
        \A1[398] , \A1[397] , \A1[396] , \A1[395] , \A1[394] , \A1[393] , 
        \A1[392] , \A1[391] , \A1[390] , \A1[389] , \A1[388] , \A1[387] , 
        \A1[386] , \A1[385] , \A1[384] , \A1[383] , \A1[382] , \A1[381] , 
        \A1[380] , \A1[379] , \A1[378] , \A1[377] , \A1[376] , \A1[375] , 
        \A1[374] , \A1[373] , \A1[372] , \A1[371] , \A1[370] , \A1[369] , 
        \A1[368] , \A1[367] , \A1[366] , \A1[365] , \A1[364] , \A1[363] , 
        \A1[362] , \A1[361] , \A1[360] , \A1[359] , \A1[358] , \A1[357] , 
        \A1[356] , \A1[355] , \A1[354] , \A1[353] , \A1[352] , \A1[351] , 
        \A1[350] , \A1[349] , \A1[348] , \A1[347] , \A1[346] , \A1[345] , 
        \A1[344] , \A1[343] , \A1[342] , \A1[341] , \A1[340] , \A1[339] , 
        \A1[338] , \A1[337] , \A1[336] , \A1[335] , \A1[334] , \A1[333] , 
        \A1[332] , \A1[331] , \A1[330] , \A1[329] , \A1[328] , \A1[327] , 
        \A1[326] , \A1[325] , \A1[324] , \A1[323] , \A1[322] , \A1[321] , 
        \A1[320] , \A1[319] , \A1[318] , \A1[317] , \A1[316] , \A1[315] , 
        \A1[314] , \A1[313] , \A1[312] , \A1[311] , \A1[310] , \A1[309] , 
        \A1[308] , \A1[307] , \A1[306] , \A1[305] , \A1[304] , \A1[303] , 
        \A1[302] , \A1[301] , \A1[300] , \A1[299] , \A1[298] , \A1[297] , 
        \A1[296] , \A1[295] , \A1[294] , \A1[293] , \A1[292] , \A1[291] , 
        \A1[290] , \A1[289] , \A1[288] , \A1[287] , \A1[286] , \A1[285] , 
        \A1[284] , \A1[283] , \A1[282] , \A1[281] , \A1[280] , \A1[279] , 
        \A1[278] , \A1[277] , \A1[276] , \A1[275] , \A1[274] , \A1[273] , 
        \A1[272] , \A1[271] , \A1[270] , \A1[269] , \A1[268] , \A1[267] , 
        \A1[266] , \A1[265] , \A1[264] , \A1[263] , \A1[262] , \A1[261] , 
        \A1[260] , \A1[259] , \A1[258] , \A1[257] , \A1[256] , \A1[255] , 
        \A1[254] , \A1[253] , \A1[252] , \A1[251] , \A1[250] , \A1[249] , 
        \A1[248] , \A1[247] , \A1[246] , \A1[245] , \A1[244] , \A1[243] , 
        \A1[242] , \A1[241] , \A1[240] , \A1[239] , \A1[238] , \A1[237] , 
        \A1[236] , \A1[235] , \A1[234] , \A1[233] , \A1[232] , \A1[231] , 
        \A1[230] , \A1[229] , \A1[228] , \A1[227] , \A1[226] , \A1[225] , 
        \A1[224] , \A1[223] , \A1[222] , \A1[221] , \A1[220] , \A1[219] , 
        \A1[218] , \A1[217] , \A1[216] , \A1[215] , \A1[214] , \A1[213] , 
        \A1[212] , \A1[211] , \A1[210] , \A1[209] , \A1[208] , \A1[207] , 
        \A1[206] , \A1[205] , \A1[204] , \A1[203] , \A1[202] , \A1[201] , 
        \A1[200] , \A1[199] , \A1[198] , \A1[197] , \A1[196] , \A1[195] , 
        \A1[194] , \A1[193] , \A1[192] , \A1[191] , \A1[190] , \A1[189] , 
        \A1[188] , \A1[187] , \A1[186] , \A1[185] , \A1[184] , \A1[183] , 
        \A1[182] , \A1[181] , \A1[180] , \A1[179] , \A1[178] , \A1[177] , 
        \A1[176] , \A1[175] , \A1[174] , \A1[173] , \A1[172] , \A1[171] , 
        \A1[170] , \A1[169] , \A1[168] , \A1[167] , \A1[166] , \A1[165] , 
        \A1[164] , \A1[163] , \A1[162] , \A1[161] , \A1[160] , \A1[159] , 
        \A1[158] , \A1[157] , \A1[156] , \A1[155] , \A1[154] , \A1[153] , 
        \A1[152] , \A1[151] , \A1[150] , \A1[149] , \A1[148] , \A1[147] , 
        \A1[146] , \A1[145] , \A1[144] , \A1[143] , \A1[142] , \A1[141] , 
        \A1[140] , \A1[139] , \A1[138] , \A1[137] , \A1[136] , \A1[135] , 
        \A1[134] , \A1[133] , \A1[132] , \A1[131] , \A1[130] , \A1[129] , 
        \A1[128] , \A1[127] , \A1[126] , \A1[125] , \A1[124] , \A1[123] , 
        \A1[122] , \A1[121] , \A1[120] , \A1[119] , \A1[118] , \A1[117] , 
        \A1[116] , \A1[115] , \A1[114] , \A1[113] , \A1[112] , \A1[111] , 
        \A1[110] , \A1[109] , \A1[108] , \A1[107] , \A1[106] , \A1[105] , 
        \A1[104] , \A1[103] , \A1[102] , \A1[101] , \A1[100] , \A1[99] , 
        \A1[98] , \A1[97] , \A1[96] , \A1[95] , \A1[94] , \A1[93] , \A1[92] , 
        \A1[91] , \A1[90] , \A1[89] , \A1[88] , \A1[87] , \A1[86] , \A1[85] , 
        \A1[84] , \A1[83] , \A1[82] , \A1[81] , \A1[80] , \A1[79] , \A1[78] , 
        \A1[77] , \A1[76] , \A1[75] , \A1[74] , \A1[73] , \A1[72] , \A1[71] , 
        \A1[70] , \A1[69] , \A1[68] , \A1[67] , \A1[66] , \A1[65] , \A1[64] , 
        \A1[63] , \A1[62] , \A1[61] , \A1[60] , \A1[59] , \A1[58] , \A1[57] , 
        \A1[56] , \A1[55] , \A1[54] , \A1[53] , \A1[52] , \A1[51] , \A1[50] , 
        \A1[49] , \A1[48] , \A1[47] , \A1[46] , \A1[45] , \A1[44] , \A1[43] , 
        \A1[42] , \A1[41] , \A1[40] , \A1[39] , \A1[38] , \A1[37] , \A1[36] , 
        \A1[35] , \A1[34] , \A1[33] , \A1[32] , \A1[31] , \A1[30] , \A1[29] , 
        \A1[28] , \A1[27] , \A1[26] , \A1[25] , \A1[24] , \A1[23] , \A1[22] , 
        \A1[21] , \A1[20] , \A1[19] , \A1[18] , \A1[17] , \A1[16] , \A1[15] , 
        \A1[14] , \A1[13] , \A1[12] , \A1[11] , \A1[10] , \A1[9] , \A1[8] , 
        \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] , \A1[1] , \A1[0] }), .B({\A2[1025] , \A2[1024] , \A2[1023] , \A2[1022] , \A2[1021] , \A2[1020] , 
        \A2[1019] , \A2[1018] , \A2[1017] , \A2[1016] , \A2[1015] , \A2[1014] , 
        \A2[1013] , \A2[1012] , \A2[1011] , \A2[1010] , \A2[1009] , \A2[1008] , 
        \A2[1007] , \A2[1006] , \A2[1005] , \A2[1004] , \A2[1003] , \A2[1002] , 
        \A2[1001] , \A2[1000] , \A2[999] , \A2[998] , \A2[997] , \A2[996] , 
        \A2[995] , \A2[994] , \A2[993] , \A2[992] , \A2[991] , \A2[990] , 
        \A2[989] , \A2[988] , \A2[987] , \A2[986] , \A2[985] , \A2[984] , 
        \A2[983] , \A2[982] , \A2[981] , \A2[980] , \A2[979] , \A2[978] , 
        \A2[977] , \A2[976] , \A2[975] , \A2[974] , \A2[973] , \A2[972] , 
        \A2[971] , \A2[970] , \A2[969] , \A2[968] , \A2[967] , \A2[966] , 
        \A2[965] , \A2[964] , \A2[963] , \A2[962] , \A2[961] , \A2[960] , 
        \A2[959] , \A2[958] , \A2[957] , \A2[956] , \A2[955] , \A2[954] , 
        \A2[953] , \A2[952] , \A2[951] , \A2[950] , \A2[949] , \A2[948] , 
        \A2[947] , \A2[946] , \A2[945] , \A2[944] , \A2[943] , \A2[942] , 
        \A2[941] , \A2[940] , \A2[939] , \A2[938] , \A2[937] , \A2[936] , 
        \A2[935] , \A2[934] , \A2[933] , \A2[932] , \A2[931] , \A2[930] , 
        \A2[929] , \A2[928] , \A2[927] , \A2[926] , \A2[925] , \A2[924] , 
        \A2[923] , \A2[922] , \A2[921] , \A2[920] , \A2[919] , \A2[918] , 
        \A2[917] , \A2[916] , \A2[915] , \A2[914] , \A2[913] , \A2[912] , 
        \A2[911] , \A2[910] , \A2[909] , \A2[908] , \A2[907] , \A2[906] , 
        \A2[905] , \A2[904] , \A2[903] , \A2[902] , \A2[901] , \A2[900] , 
        \A2[899] , \A2[898] , \A2[897] , \A2[896] , \A2[895] , \A2[894] , 
        \A2[893] , \A2[892] , \A2[891] , \A2[890] , \A2[889] , \A2[888] , 
        \A2[887] , \A2[886] , \A2[885] , \A2[884] , \A2[883] , \A2[882] , 
        \A2[881] , \A2[880] , \A2[879] , \A2[878] , \A2[877] , \A2[876] , 
        \A2[875] , \A2[874] , \A2[873] , \A2[872] , \A2[871] , \A2[870] , 
        \A2[869] , \A2[868] , \A2[867] , \A2[866] , \A2[865] , \A2[864] , 
        \A2[863] , \A2[862] , \A2[861] , \A2[860] , \A2[859] , \A2[858] , 
        \A2[857] , \A2[856] , \A2[855] , \A2[854] , \A2[853] , \A2[852] , 
        \A2[851] , \A2[850] , \A2[849] , \A2[848] , \A2[847] , \A2[846] , 
        \A2[845] , \A2[844] , \A2[843] , \A2[842] , \A2[841] , \A2[840] , 
        \A2[839] , \A2[838] , \A2[837] , \A2[836] , \A2[835] , \A2[834] , 
        \A2[833] , \A2[832] , \A2[831] , \A2[830] , \A2[829] , \A2[828] , 
        \A2[827] , \A2[826] , \A2[825] , \A2[824] , \A2[823] , \A2[822] , 
        \A2[821] , \A2[820] , \A2[819] , \A2[818] , \A2[817] , \A2[816] , 
        \A2[815] , \A2[814] , \A2[813] , \A2[812] , \A2[811] , \A2[810] , 
        \A2[809] , \A2[808] , \A2[807] , \A2[806] , \A2[805] , \A2[804] , 
        \A2[803] , \A2[802] , \A2[801] , \A2[800] , \A2[799] , \A2[798] , 
        \A2[797] , \A2[796] , \A2[795] , \A2[794] , \A2[793] , \A2[792] , 
        \A2[791] , \A2[790] , \A2[789] , \A2[788] , \A2[787] , \A2[786] , 
        \A2[785] , \A2[784] , \A2[783] , \A2[782] , \A2[781] , \A2[780] , 
        \A2[779] , \A2[778] , \A2[777] , \A2[776] , \A2[775] , \A2[774] , 
        \A2[773] , \A2[772] , \A2[771] , \A2[770] , \A2[769] , \A2[768] , 
        \A2[767] , \A2[766] , \A2[765] , \A2[764] , \A2[763] , \A2[762] , 
        \A2[761] , \A2[760] , \A2[759] , \A2[758] , \A2[757] , \A2[756] , 
        \A2[755] , \A2[754] , \A2[753] , \A2[752] , \A2[751] , \A2[750] , 
        \A2[749] , \A2[748] , \A2[747] , \A2[746] , \A2[745] , \A2[744] , 
        \A2[743] , \A2[742] , \A2[741] , \A2[740] , \A2[739] , \A2[738] , 
        \A2[737] , \A2[736] , \A2[735] , \A2[734] , \A2[733] , \A2[732] , 
        \A2[731] , \A2[730] , \A2[729] , \A2[728] , \A2[727] , \A2[726] , 
        \A2[725] , \A2[724] , \A2[723] , \A2[722] , \A2[721] , \A2[720] , 
        \A2[719] , \A2[718] , \A2[717] , \A2[716] , \A2[715] , \A2[714] , 
        \A2[713] , \A2[712] , \A2[711] , \A2[710] , \A2[709] , \A2[708] , 
        \A2[707] , \A2[706] , \A2[705] , \A2[704] , \A2[703] , \A2[702] , 
        \A2[701] , \A2[700] , \A2[699] , \A2[698] , \A2[697] , \A2[696] , 
        \A2[695] , \A2[694] , \A2[693] , \A2[692] , \A2[691] , \A2[690] , 
        \A2[689] , \A2[688] , \A2[687] , \A2[686] , \A2[685] , \A2[684] , 
        \A2[683] , \A2[682] , \A2[681] , \A2[680] , \A2[679] , \A2[678] , 
        \A2[677] , \A2[676] , \A2[675] , \A2[674] , \A2[673] , \A2[672] , 
        \A2[671] , \A2[670] , \A2[669] , \A2[668] , \A2[667] , \A2[666] , 
        \A2[665] , \A2[664] , \A2[663] , \A2[662] , \A2[661] , \A2[660] , 
        \A2[659] , \A2[658] , \A2[657] , \A2[656] , \A2[655] , \A2[654] , 
        \A2[653] , \A2[652] , \A2[651] , \A2[650] , \A2[649] , \A2[648] , 
        \A2[647] , \A2[646] , \A2[645] , \A2[644] , \A2[643] , \A2[642] , 
        \A2[641] , \A2[640] , \A2[639] , \A2[638] , \A2[637] , \A2[636] , 
        \A2[635] , \A2[634] , \A2[633] , \A2[632] , \A2[631] , \A2[630] , 
        \A2[629] , \A2[628] , \A2[627] , \A2[626] , \A2[625] , \A2[624] , 
        \A2[623] , \A2[622] , \A2[621] , \A2[620] , \A2[619] , \A2[618] , 
        \A2[617] , \A2[616] , \A2[615] , \A2[614] , \A2[613] , \A2[612] , 
        \A2[611] , \A2[610] , \A2[609] , \A2[608] , \A2[607] , \A2[606] , 
        \A2[605] , \A2[604] , \A2[603] , \A2[602] , \A2[601] , \A2[600] , 
        \A2[599] , \A2[598] , \A2[597] , \A2[596] , \A2[595] , \A2[594] , 
        \A2[593] , \A2[592] , \A2[591] , \A2[590] , \A2[589] , \A2[588] , 
        \A2[587] , \A2[586] , \A2[585] , \A2[584] , \A2[583] , \A2[582] , 
        \A2[581] , \A2[580] , \A2[579] , \A2[578] , \A2[577] , \A2[576] , 
        \A2[575] , \A2[574] , \A2[573] , \A2[572] , \A2[571] , \A2[570] , 
        \A2[569] , \A2[568] , \A2[567] , \A2[566] , \A2[565] , \A2[564] , 
        \A2[563] , \A2[562] , \A2[561] , \A2[560] , \A2[559] , \A2[558] , 
        \A2[557] , \A2[556] , \A2[555] , \A2[554] , \A2[553] , \A2[552] , 
        \A2[551] , \A2[550] , \A2[549] , \A2[548] , \A2[547] , \A2[546] , 
        \A2[545] , \A2[544] , \A2[543] , \A2[542] , \A2[541] , \A2[540] , 
        \A2[539] , \A2[538] , \A2[537] , \A2[536] , \A2[535] , \A2[534] , 
        \A2[533] , \A2[532] , \A2[531] , \A2[530] , \A2[529] , \A2[528] , 
        \A2[527] , \A2[526] , \A2[525] , \A2[524] , \A2[523] , \A2[522] , 
        \A2[521] , \A2[520] , \A2[519] , \A2[518] , \A2[517] , \A2[516] , 
        \A2[515] , \A2[514] , \A2[513] , \A2[512] , \A2[511] , \A2[510] , 
        \A2[509] , \A2[508] , \A2[507] , \A2[506] , \A2[505] , \A2[504] , 
        \A2[503] , \A2[502] , \A2[501] , \A2[500] , \A2[499] , \A2[498] , 
        \A2[497] , \A2[496] , \A2[495] , \A2[494] , \A2[493] , \A2[492] , 
        \A2[491] , \A2[490] , \A2[489] , \A2[488] , \A2[487] , \A2[486] , 
        \A2[485] , \A2[484] , \A2[483] , \A2[482] , \A2[481] , \A2[480] , 
        \A2[479] , \A2[478] , \A2[477] , \A2[476] , \A2[475] , \A2[474] , 
        \A2[473] , \A2[472] , \A2[471] , \A2[470] , \A2[469] , \A2[468] , 
        \A2[467] , \A2[466] , \A2[465] , \A2[464] , \A2[463] , \A2[462] , 
        \A2[461] , \A2[460] , \A2[459] , \A2[458] , \A2[457] , \A2[456] , 
        \A2[455] , \A2[454] , \A2[453] , \A2[452] , \A2[451] , \A2[450] , 
        \A2[449] , \A2[448] , \A2[447] , \A2[446] , \A2[445] , \A2[444] , 
        \A2[443] , \A2[442] , \A2[441] , \A2[440] , \A2[439] , \A2[438] , 
        \A2[437] , \A2[436] , \A2[435] , \A2[434] , \A2[433] , \A2[432] , 
        \A2[431] , \A2[430] , \A2[429] , \A2[428] , \A2[427] , \A2[426] , 
        \A2[425] , \A2[424] , \A2[423] , \A2[422] , \A2[421] , \A2[420] , 
        \A2[419] , \A2[418] , \A2[417] , \A2[416] , \A2[415] , \A2[414] , 
        \A2[413] , \A2[412] , \A2[411] , \A2[410] , \A2[409] , \A2[408] , 
        \A2[407] , \A2[406] , \A2[405] , \A2[404] , \A2[403] , \A2[402] , 
        \A2[401] , \A2[400] , \A2[399] , \A2[398] , \A2[397] , \A2[396] , 
        \A2[395] , \A2[394] , \A2[393] , \A2[392] , \A2[391] , \A2[390] , 
        \A2[389] , \A2[388] , \A2[387] , \A2[386] , \A2[385] , \A2[384] , 
        \A2[383] , \A2[382] , \A2[381] , \A2[380] , \A2[379] , \A2[378] , 
        \A2[377] , \A2[376] , \A2[375] , \A2[374] , \A2[373] , \A2[372] , 
        \A2[371] , \A2[370] , \A2[369] , \A2[368] , \A2[367] , \A2[366] , 
        \A2[365] , \A2[364] , \A2[363] , \A2[362] , \A2[361] , \A2[360] , 
        \A2[359] , \A2[358] , \A2[357] , \A2[356] , \A2[355] , \A2[354] , 
        \A2[353] , \A2[352] , \A2[351] , \A2[350] , \A2[349] , \A2[348] , 
        \A2[347] , \A2[346] , \A2[345] , \A2[344] , \A2[343] , \A2[342] , 
        \A2[341] , \A2[340] , \A2[339] , \A2[338] , \A2[337] , \A2[336] , 
        \A2[335] , \A2[334] , \A2[333] , \A2[332] , \A2[331] , \A2[330] , 
        \A2[329] , \A2[328] , \A2[327] , \A2[326] , \A2[325] , \A2[324] , 
        \A2[323] , \A2[322] , \A2[321] , \A2[320] , \A2[319] , \A2[318] , 
        \A2[317] , \A2[316] , \A2[315] , \A2[314] , \A2[313] , \A2[312] , 
        \A2[311] , \A2[310] , \A2[309] , \A2[308] , \A2[307] , \A2[306] , 
        \A2[305] , \A2[304] , \A2[303] , \A2[302] , \A2[301] , \A2[300] , 
        \A2[299] , \A2[298] , \A2[297] , \A2[296] , \A2[295] , \A2[294] , 
        \A2[293] , \A2[292] , \A2[291] , \A2[290] , \A2[289] , \A2[288] , 
        \A2[287] , \A2[286] , \A2[285] , \A2[284] , \A2[283] , \A2[282] , 
        \A2[281] , \A2[280] , \A2[279] , \A2[278] , \A2[277] , \A2[276] , 
        \A2[275] , \A2[274] , \A2[273] , \A2[272] , \A2[271] , \A2[270] , 
        \A2[269] , \A2[268] , \A2[267] , \A2[266] , \A2[265] , \A2[264] , 
        \A2[263] , \A2[262] , \A2[261] , \A2[260] , \A2[259] , \A2[258] , 
        \A2[257] , \A2[256] , \A2[255] , \A2[254] , \A2[253] , \A2[252] , 
        \A2[251] , \A2[250] , \A2[249] , \A2[248] , \A2[247] , \A2[246] , 
        \A2[245] , \A2[244] , \A2[243] , \A2[242] , \A2[241] , \A2[240] , 
        \A2[239] , \A2[238] , \A2[237] , \A2[236] , \A2[235] , \A2[234] , 
        \A2[233] , \A2[232] , \A2[231] , \A2[230] , \A2[229] , \A2[228] , 
        \A2[227] , \A2[226] , \A2[225] , \A2[224] , \A2[223] , \A2[222] , 
        \A2[221] , \A2[220] , \A2[219] , \A2[218] , \A2[217] , \A2[216] , 
        \A2[215] , \A2[214] , \A2[213] , \A2[212] , \A2[211] , \A2[210] , 
        \A2[209] , \A2[208] , \A2[207] , \A2[206] , \A2[205] , \A2[204] , 
        \A2[203] , \A2[202] , \A2[201] , \A2[200] , \A2[199] , \A2[198] , 
        \A2[197] , \A2[196] , \A2[195] , \A2[194] , \A2[193] , \A2[192] , 
        \A2[191] , \A2[190] , \A2[189] , \A2[188] , \A2[187] , \A2[186] , 
        \A2[185] , \A2[184] , \A2[183] , \A2[182] , \A2[181] , \A2[180] , 
        \A2[179] , \A2[178] , \A2[177] , \A2[176] , \A2[175] , \A2[174] , 
        \A2[173] , \A2[172] , \A2[171] , \A2[170] , \A2[169] , \A2[168] , 
        \A2[167] , \A2[166] , \A2[165] , \A2[164] , \A2[163] , \A2[162] , 
        \A2[161] , \A2[160] , \A2[159] , \A2[158] , \A2[157] , \A2[156] , 
        \A2[155] , \A2[154] , \A2[153] , \A2[152] , \A2[151] , \A2[150] , 
        \A2[149] , \A2[148] , \A2[147] , \A2[146] , \A2[145] , \A2[144] , 
        \A2[143] , \A2[142] , \A2[141] , \A2[140] , \A2[139] , \A2[138] , 
        \A2[137] , \A2[136] , \A2[135] , \A2[134] , \A2[133] , \A2[132] , 
        \A2[131] , \A2[130] , \A2[129] , \A2[128] , \A2[127] , \A2[126] , 
        \A2[125] , \A2[124] , \A2[123] , \A2[122] , \A2[121] , \A2[120] , 
        \A2[119] , \A2[118] , \A2[117] , \A2[116] , \A2[115] , \A2[114] , 
        \A2[113] , \A2[112] , \A2[111] , \A2[110] , \A2[109] , \A2[108] , 
        \A2[107] , \A2[106] , \A2[105] , \A2[104] , \A2[103] , \A2[102] , 
        \A2[101] , \A2[100] , \A2[99] , \A2[98] , \A2[97] , \A2[96] , \A2[95] , 
        \A2[94] , \A2[93] , \A2[92] , \A2[91] , \A2[90] , \A2[89] , \A2[88] , 
        \A2[87] , \A2[86] , \A2[85] , \A2[84] , \A2[83] , \A2[82] , \A2[81] , 
        \A2[80] , \A2[79] , \A2[78] , \A2[77] , \A2[76] , \A2[75] , \A2[74] , 
        \A2[73] , \A2[72] , \A2[71] , \A2[70] , \A2[69] , \A2[68] , \A2[67] , 
        \A2[66] , \A2[65] , \A2[64] , \A2[63] , \A2[62] , \A2[61] , \A2[60] , 
        \A2[59] , \A2[58] , \A2[57] , \A2[56] , \A2[55] , \A2[54] , \A2[53] , 
        \A2[52] , \A2[51] , \A2[50] , \A2[49] , \A2[48] , \A2[47] , \A2[46] , 
        \A2[45] , \A2[44] , \A2[43] , \A2[42] , \A2[41] , \A2[40] , \A2[39] , 
        \A2[38] , \A2[37] , \A2[36] , \A2[35] , \A2[34] , \A2[33] , \A2[32] , 
        \A2[31] , \A2[30] , \A2[29] , \A2[28] , \A2[27] , \A2[26] , \A2[25] , 
        \A2[24] , \A2[23] , \A2[22] , \A2[21] , \A2[20] , \A2[19] , \A2[18] , 
        \A2[17] , \A2[16] , \A2[15] , \A2[14] , \A2[13] , \A2[12] , \A2[11] , 
        \A2[10] , \A2[9] , \A2[8] , \A2[7] , \A2[6] , \A2[5] , \A2[4] , 
        \A2[3] , 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, PRODUCT[1023:2]}) );
  NANDN U2 ( .A(n19142), .B(n19141), .Z(n19137) );
  NANDN U3 ( .A(n19176), .B(n19175), .Z(n19171) );
  NANDN U4 ( .A(n19210), .B(n19209), .Z(n19205) );
  NANDN U5 ( .A(n19244), .B(n19243), .Z(n19239) );
  NANDN U6 ( .A(n19304), .B(n19303), .Z(n19299) );
  NANDN U7 ( .A(n19338), .B(n19337), .Z(n19333) );
  NANDN U8 ( .A(n19372), .B(n19371), .Z(n19367) );
  NANDN U9 ( .A(n19406), .B(n19405), .Z(n19401) );
  NANDN U10 ( .A(n2141), .B(n2140), .Z(n2136) );
  NANDN U11 ( .A(n2175), .B(n2174), .Z(n2170) );
  NANDN U12 ( .A(n2209), .B(n2208), .Z(n2204) );
  NANDN U13 ( .A(n2243), .B(n2242), .Z(n2238) );
  NANDN U14 ( .A(n2292), .B(n2291), .Z(n2287) );
  NANDN U15 ( .A(n2326), .B(n2325), .Z(n2321) );
  NANDN U16 ( .A(n2360), .B(n2359), .Z(n2355) );
  NANDN U17 ( .A(n2394), .B(n2393), .Z(n2389) );
  NANDN U18 ( .A(n2428), .B(n2427), .Z(n2423) );
  NANDN U19 ( .A(n2480), .B(n2479), .Z(n2475) );
  NANDN U20 ( .A(n2514), .B(n2513), .Z(n2509) );
  NANDN U21 ( .A(n2548), .B(n2547), .Z(n2543) );
  NANDN U22 ( .A(n2582), .B(n2581), .Z(n2577) );
  NANDN U23 ( .A(n2616), .B(n2615), .Z(n2611) );
  NANDN U24 ( .A(n2667), .B(n2666), .Z(n2662) );
  NANDN U25 ( .A(n2701), .B(n2700), .Z(n2696) );
  NANDN U26 ( .A(n2735), .B(n2734), .Z(n2730) );
  NANDN U27 ( .A(n2769), .B(n2768), .Z(n2764) );
  NANDN U28 ( .A(n2803), .B(n2802), .Z(n2798) );
  NANDN U29 ( .A(n2854), .B(n2853), .Z(n2849) );
  NANDN U30 ( .A(n2888), .B(n2887), .Z(n2883) );
  NANDN U31 ( .A(n2922), .B(n2921), .Z(n2917) );
  NANDN U32 ( .A(n2956), .B(n2955), .Z(n2951) );
  NANDN U33 ( .A(n2990), .B(n2989), .Z(n2985) );
  NANDN U34 ( .A(n3041), .B(n3040), .Z(n3036) );
  NANDN U35 ( .A(n3075), .B(n3074), .Z(n3070) );
  NANDN U36 ( .A(n3109), .B(n3108), .Z(n3104) );
  NANDN U37 ( .A(n3143), .B(n3142), .Z(n3138) );
  NANDN U38 ( .A(n3177), .B(n3176), .Z(n3172) );
  NANDN U39 ( .A(n3228), .B(n3227), .Z(n3223) );
  NANDN U40 ( .A(n3262), .B(n3261), .Z(n3257) );
  NANDN U41 ( .A(n3296), .B(n3295), .Z(n3291) );
  NANDN U42 ( .A(n3330), .B(n3329), .Z(n3325) );
  NANDN U43 ( .A(n3364), .B(n3363), .Z(n3359) );
  NANDN U44 ( .A(n3415), .B(n3414), .Z(n3410) );
  NANDN U45 ( .A(n3449), .B(n3448), .Z(n3444) );
  NANDN U46 ( .A(n3483), .B(n3482), .Z(n3478) );
  NANDN U47 ( .A(n3517), .B(n3516), .Z(n3512) );
  NANDN U48 ( .A(n3551), .B(n3550), .Z(n3546) );
  NANDN U49 ( .A(n3602), .B(n3601), .Z(n3597) );
  NANDN U50 ( .A(n3636), .B(n3635), .Z(n3631) );
  NANDN U51 ( .A(n3670), .B(n3669), .Z(n3665) );
  NANDN U52 ( .A(n3704), .B(n3703), .Z(n3699) );
  NANDN U53 ( .A(n3738), .B(n3737), .Z(n3733) );
  NANDN U54 ( .A(n3789), .B(n3788), .Z(n3784) );
  NANDN U55 ( .A(n3823), .B(n3822), .Z(n3818) );
  NANDN U56 ( .A(n3857), .B(n3856), .Z(n3852) );
  NANDN U57 ( .A(n3891), .B(n3890), .Z(n3886) );
  NANDN U58 ( .A(n3925), .B(n3924), .Z(n3920) );
  NANDN U59 ( .A(n3991), .B(n3990), .Z(n3986) );
  NANDN U60 ( .A(n4025), .B(n4024), .Z(n4020) );
  NANDN U61 ( .A(n4059), .B(n4058), .Z(n4054) );
  NANDN U62 ( .A(n4093), .B(n4092), .Z(n4088) );
  NANDN U63 ( .A(n4127), .B(n4126), .Z(n4122) );
  NANDN U64 ( .A(n4178), .B(n4177), .Z(n4173) );
  NANDN U65 ( .A(n4212), .B(n4211), .Z(n4207) );
  NANDN U66 ( .A(n4246), .B(n4245), .Z(n4241) );
  NANDN U67 ( .A(n4280), .B(n4279), .Z(n4275) );
  NANDN U68 ( .A(n4314), .B(n4313), .Z(n4309) );
  NANDN U69 ( .A(n4365), .B(n4364), .Z(n4360) );
  NANDN U70 ( .A(n4399), .B(n4398), .Z(n4394) );
  NANDN U71 ( .A(n4433), .B(n4432), .Z(n4428) );
  NANDN U72 ( .A(n4467), .B(n4466), .Z(n4462) );
  NANDN U73 ( .A(n4501), .B(n4500), .Z(n4496) );
  NANDN U74 ( .A(n4552), .B(n4551), .Z(n4547) );
  NANDN U75 ( .A(n4586), .B(n4585), .Z(n4581) );
  NANDN U76 ( .A(n4620), .B(n4619), .Z(n4615) );
  NANDN U77 ( .A(n4654), .B(n4653), .Z(n4649) );
  NANDN U78 ( .A(n4688), .B(n4687), .Z(n4683) );
  NANDN U79 ( .A(n4739), .B(n4738), .Z(n4734) );
  NANDN U80 ( .A(n4773), .B(n4772), .Z(n4768) );
  NANDN U81 ( .A(n4807), .B(n4806), .Z(n4802) );
  NANDN U82 ( .A(n4841), .B(n4840), .Z(n4836) );
  NANDN U83 ( .A(n4875), .B(n4874), .Z(n4870) );
  NANDN U84 ( .A(n4926), .B(n4925), .Z(n4921) );
  NANDN U85 ( .A(n4960), .B(n4959), .Z(n4955) );
  NANDN U86 ( .A(n4994), .B(n4993), .Z(n4989) );
  NANDN U87 ( .A(n5028), .B(n5027), .Z(n5023) );
  NANDN U88 ( .A(n5062), .B(n5061), .Z(n5057) );
  NANDN U89 ( .A(n5113), .B(n5112), .Z(n5108) );
  NANDN U90 ( .A(n5147), .B(n5146), .Z(n5142) );
  NANDN U91 ( .A(n5181), .B(n5180), .Z(n5176) );
  NANDN U92 ( .A(n5215), .B(n5214), .Z(n5210) );
  NANDN U93 ( .A(n5249), .B(n5248), .Z(n5244) );
  NANDN U94 ( .A(n5300), .B(n5299), .Z(n5295) );
  NANDN U95 ( .A(n5334), .B(n5333), .Z(n5329) );
  NANDN U96 ( .A(n5368), .B(n5367), .Z(n5363) );
  NANDN U97 ( .A(n5402), .B(n5401), .Z(n5397) );
  NANDN U98 ( .A(n5436), .B(n5435), .Z(n5431) );
  NANDN U99 ( .A(n5487), .B(n5486), .Z(n5482) );
  NANDN U100 ( .A(n5521), .B(n5520), .Z(n5516) );
  NANDN U101 ( .A(n5555), .B(n5554), .Z(n5550) );
  NANDN U102 ( .A(n5589), .B(n5588), .Z(n5584) );
  NANDN U103 ( .A(n5623), .B(n5622), .Z(n5618) );
  NANDN U104 ( .A(n5674), .B(n5673), .Z(n5669) );
  NANDN U105 ( .A(n5708), .B(n5707), .Z(n5703) );
  NANDN U106 ( .A(n5742), .B(n5741), .Z(n5737) );
  NANDN U107 ( .A(n5776), .B(n5775), .Z(n5771) );
  NANDN U108 ( .A(n5810), .B(n5809), .Z(n5805) );
  NANDN U109 ( .A(n5879), .B(n5878), .Z(n5874) );
  NANDN U110 ( .A(n5913), .B(n5912), .Z(n5908) );
  NANDN U111 ( .A(n5947), .B(n5946), .Z(n5942) );
  NANDN U112 ( .A(n5981), .B(n5980), .Z(n5976) );
  NANDN U113 ( .A(n6015), .B(n6014), .Z(n6010) );
  NANDN U114 ( .A(n6066), .B(n6065), .Z(n6061) );
  NANDN U115 ( .A(n6100), .B(n6099), .Z(n6095) );
  NANDN U116 ( .A(n6134), .B(n6133), .Z(n6129) );
  NANDN U117 ( .A(n6168), .B(n6167), .Z(n6163) );
  NANDN U118 ( .A(n6202), .B(n6201), .Z(n6197) );
  NANDN U119 ( .A(n6253), .B(n6252), .Z(n6248) );
  NANDN U120 ( .A(n6287), .B(n6286), .Z(n6282) );
  NANDN U121 ( .A(n6321), .B(n6320), .Z(n6316) );
  NANDN U122 ( .A(n6355), .B(n6354), .Z(n6350) );
  NANDN U123 ( .A(n6389), .B(n6388), .Z(n6384) );
  NANDN U124 ( .A(n6440), .B(n6439), .Z(n6435) );
  NANDN U125 ( .A(n6474), .B(n6473), .Z(n6469) );
  NANDN U126 ( .A(n6508), .B(n6507), .Z(n6503) );
  NANDN U127 ( .A(n6542), .B(n6541), .Z(n6537) );
  NANDN U128 ( .A(n6576), .B(n6575), .Z(n6571) );
  NANDN U129 ( .A(n6627), .B(n6626), .Z(n6622) );
  NANDN U130 ( .A(n6661), .B(n6660), .Z(n6656) );
  NANDN U131 ( .A(n6695), .B(n6694), .Z(n6690) );
  NANDN U132 ( .A(n6729), .B(n6728), .Z(n6724) );
  NANDN U133 ( .A(n6763), .B(n6762), .Z(n6758) );
  NANDN U134 ( .A(n6814), .B(n6813), .Z(n6809) );
  NANDN U135 ( .A(n6848), .B(n6847), .Z(n6843) );
  NANDN U136 ( .A(n6882), .B(n6881), .Z(n6877) );
  NANDN U137 ( .A(n6916), .B(n6915), .Z(n6911) );
  NANDN U138 ( .A(n6950), .B(n6949), .Z(n6945) );
  NANDN U139 ( .A(n7001), .B(n7000), .Z(n6996) );
  NANDN U140 ( .A(n7035), .B(n7034), .Z(n7030) );
  NANDN U141 ( .A(n7069), .B(n7068), .Z(n7064) );
  NANDN U142 ( .A(n7103), .B(n7102), .Z(n7098) );
  NANDN U143 ( .A(n7137), .B(n7136), .Z(n7132) );
  NANDN U144 ( .A(n7188), .B(n7187), .Z(n7183) );
  NANDN U145 ( .A(n7222), .B(n7221), .Z(n7217) );
  NANDN U146 ( .A(n7256), .B(n7255), .Z(n7251) );
  NANDN U147 ( .A(n7290), .B(n7289), .Z(n7285) );
  NANDN U148 ( .A(n7324), .B(n7323), .Z(n7319) );
  NANDN U149 ( .A(n7375), .B(n7374), .Z(n7370) );
  NANDN U150 ( .A(n7409), .B(n7408), .Z(n7404) );
  NANDN U151 ( .A(n7443), .B(n7442), .Z(n7438) );
  NANDN U152 ( .A(n7477), .B(n7476), .Z(n7472) );
  NANDN U153 ( .A(n7511), .B(n7510), .Z(n7506) );
  NANDN U154 ( .A(n7562), .B(n7561), .Z(n7557) );
  NANDN U155 ( .A(n7596), .B(n7595), .Z(n7591) );
  NANDN U156 ( .A(n7630), .B(n7629), .Z(n7625) );
  NANDN U157 ( .A(n7664), .B(n7663), .Z(n7659) );
  NANDN U158 ( .A(n7698), .B(n7697), .Z(n7693) );
  NANDN U159 ( .A(n7766), .B(n7765), .Z(n7761) );
  NANDN U160 ( .A(n7800), .B(n7799), .Z(n7795) );
  NANDN U161 ( .A(n7834), .B(n7833), .Z(n7829) );
  NANDN U162 ( .A(n7868), .B(n7867), .Z(n7863) );
  NANDN U163 ( .A(n7902), .B(n7901), .Z(n7897) );
  NANDN U164 ( .A(n7953), .B(n7952), .Z(n7948) );
  NANDN U165 ( .A(n7987), .B(n7986), .Z(n7982) );
  NANDN U166 ( .A(n8021), .B(n8020), .Z(n8016) );
  NANDN U167 ( .A(n8055), .B(n8054), .Z(n8050) );
  NANDN U168 ( .A(n8089), .B(n8088), .Z(n8084) );
  NANDN U169 ( .A(n8140), .B(n8139), .Z(n8135) );
  NANDN U170 ( .A(n8174), .B(n8173), .Z(n8169) );
  NANDN U171 ( .A(n8208), .B(n8207), .Z(n8203) );
  NANDN U172 ( .A(n8242), .B(n8241), .Z(n8237) );
  NANDN U173 ( .A(n8276), .B(n8275), .Z(n8271) );
  NANDN U174 ( .A(n8327), .B(n8326), .Z(n8322) );
  NANDN U175 ( .A(n8361), .B(n8360), .Z(n8356) );
  NANDN U176 ( .A(n8395), .B(n8394), .Z(n8390) );
  NANDN U177 ( .A(n8429), .B(n8428), .Z(n8424) );
  NANDN U178 ( .A(n8463), .B(n8462), .Z(n8458) );
  NANDN U179 ( .A(n8514), .B(n8513), .Z(n8509) );
  NANDN U180 ( .A(n8548), .B(n8547), .Z(n8543) );
  NANDN U181 ( .A(n8582), .B(n8581), .Z(n8577) );
  NANDN U182 ( .A(n8616), .B(n8615), .Z(n8611) );
  NANDN U183 ( .A(n8650), .B(n8649), .Z(n8645) );
  NANDN U184 ( .A(n8701), .B(n8700), .Z(n8696) );
  NANDN U185 ( .A(n8735), .B(n8734), .Z(n8730) );
  NANDN U186 ( .A(n8769), .B(n8768), .Z(n8764) );
  NANDN U187 ( .A(n8803), .B(n8802), .Z(n8798) );
  NANDN U188 ( .A(n8837), .B(n8836), .Z(n8832) );
  NANDN U189 ( .A(n8888), .B(n8887), .Z(n8883) );
  NANDN U190 ( .A(n8922), .B(n8921), .Z(n8917) );
  NANDN U191 ( .A(n8956), .B(n8955), .Z(n8951) );
  NANDN U192 ( .A(n8990), .B(n8989), .Z(n8985) );
  NANDN U193 ( .A(n9024), .B(n9023), .Z(n9019) );
  NANDN U194 ( .A(n9075), .B(n9074), .Z(n9070) );
  NANDN U195 ( .A(n9109), .B(n9108), .Z(n9104) );
  NANDN U196 ( .A(n9143), .B(n9142), .Z(n9138) );
  NANDN U197 ( .A(n9177), .B(n9176), .Z(n9172) );
  NANDN U198 ( .A(n9211), .B(n9210), .Z(n9206) );
  NANDN U199 ( .A(n9262), .B(n9261), .Z(n9257) );
  NANDN U200 ( .A(n9296), .B(n9295), .Z(n9291) );
  NANDN U201 ( .A(n9330), .B(n9329), .Z(n9325) );
  NANDN U202 ( .A(n9364), .B(n9363), .Z(n9359) );
  NANDN U203 ( .A(n9398), .B(n9397), .Z(n9393) );
  NANDN U204 ( .A(n9449), .B(n9448), .Z(n9444) );
  NANDN U205 ( .A(n9483), .B(n9482), .Z(n9478) );
  NANDN U206 ( .A(n9517), .B(n9516), .Z(n9512) );
  NANDN U207 ( .A(n9551), .B(n9550), .Z(n9546) );
  NANDN U208 ( .A(n9585), .B(n9584), .Z(n9580) );
  NANDN U209 ( .A(n9653), .B(n9652), .Z(n9648) );
  NANDN U210 ( .A(n9687), .B(n9686), .Z(n9682) );
  NANDN U211 ( .A(n9721), .B(n9720), .Z(n9716) );
  NANDN U212 ( .A(n9755), .B(n9754), .Z(n9750) );
  NANDN U213 ( .A(n9789), .B(n9788), .Z(n9784) );
  NANDN U214 ( .A(n9840), .B(n9839), .Z(n9835) );
  NANDN U215 ( .A(n9874), .B(n9873), .Z(n9869) );
  NANDN U216 ( .A(n9908), .B(n9907), .Z(n9903) );
  NANDN U217 ( .A(n9942), .B(n9941), .Z(n9937) );
  NANDN U218 ( .A(n9976), .B(n9975), .Z(n9971) );
  NANDN U219 ( .A(n10027), .B(n10026), .Z(n10022) );
  NANDN U220 ( .A(n10061), .B(n10060), .Z(n10056) );
  NANDN U221 ( .A(n10095), .B(n10094), .Z(n10090) );
  NANDN U222 ( .A(n10129), .B(n10128), .Z(n10124) );
  NANDN U223 ( .A(n10163), .B(n10162), .Z(n10158) );
  NANDN U224 ( .A(n10214), .B(n10213), .Z(n10209) );
  NANDN U225 ( .A(n10248), .B(n10247), .Z(n10243) );
  NANDN U226 ( .A(n10282), .B(n10281), .Z(n10277) );
  NANDN U227 ( .A(n10316), .B(n10315), .Z(n10311) );
  NANDN U228 ( .A(n10350), .B(n10349), .Z(n10345) );
  NANDN U229 ( .A(n10401), .B(n10400), .Z(n10396) );
  NANDN U230 ( .A(n10435), .B(n10434), .Z(n10430) );
  NANDN U231 ( .A(n10469), .B(n10468), .Z(n10464) );
  NANDN U232 ( .A(n10503), .B(n10502), .Z(n10498) );
  NANDN U233 ( .A(n10537), .B(n10536), .Z(n10532) );
  NANDN U234 ( .A(n10588), .B(n10587), .Z(n10583) );
  NANDN U235 ( .A(n10622), .B(n10621), .Z(n10617) );
  NANDN U236 ( .A(n10656), .B(n10655), .Z(n10651) );
  NANDN U237 ( .A(n10690), .B(n10689), .Z(n10685) );
  NANDN U238 ( .A(n10724), .B(n10723), .Z(n10719) );
  NANDN U239 ( .A(n10775), .B(n10774), .Z(n10770) );
  NANDN U240 ( .A(n10809), .B(n10808), .Z(n10804) );
  NANDN U241 ( .A(n10843), .B(n10842), .Z(n10838) );
  NANDN U242 ( .A(n10877), .B(n10876), .Z(n10872) );
  NANDN U243 ( .A(n10911), .B(n10910), .Z(n10906) );
  NANDN U244 ( .A(n10962), .B(n10961), .Z(n10957) );
  NANDN U245 ( .A(n10996), .B(n10995), .Z(n10991) );
  NANDN U246 ( .A(n11030), .B(n11029), .Z(n11025) );
  NANDN U247 ( .A(n11064), .B(n11063), .Z(n11059) );
  NANDN U248 ( .A(n11098), .B(n11097), .Z(n11093) );
  NANDN U249 ( .A(n11149), .B(n11148), .Z(n11144) );
  NANDN U250 ( .A(n11183), .B(n11182), .Z(n11178) );
  NANDN U251 ( .A(n11217), .B(n11216), .Z(n11212) );
  NANDN U252 ( .A(n11251), .B(n11250), .Z(n11246) );
  NANDN U253 ( .A(n11285), .B(n11284), .Z(n11280) );
  NANDN U254 ( .A(n11336), .B(n11335), .Z(n11331) );
  NANDN U255 ( .A(n11370), .B(n11369), .Z(n11365) );
  NANDN U256 ( .A(n11404), .B(n11403), .Z(n11399) );
  NANDN U257 ( .A(n11438), .B(n11437), .Z(n11433) );
  NANDN U258 ( .A(n11472), .B(n11471), .Z(n11467) );
  NANDN U259 ( .A(n11540), .B(n11539), .Z(n11535) );
  NANDN U260 ( .A(n11574), .B(n11573), .Z(n11569) );
  NANDN U261 ( .A(n11608), .B(n11607), .Z(n11603) );
  NANDN U262 ( .A(n11642), .B(n11641), .Z(n11637) );
  NANDN U263 ( .A(n11676), .B(n11675), .Z(n11671) );
  NANDN U264 ( .A(n11727), .B(n11726), .Z(n11722) );
  NANDN U265 ( .A(n11761), .B(n11760), .Z(n11756) );
  NANDN U266 ( .A(n11795), .B(n11794), .Z(n11790) );
  NANDN U267 ( .A(n11829), .B(n11828), .Z(n11824) );
  NANDN U268 ( .A(n11863), .B(n11862), .Z(n11858) );
  NANDN U269 ( .A(n11914), .B(n11913), .Z(n11909) );
  NANDN U270 ( .A(n11948), .B(n11947), .Z(n11943) );
  NANDN U271 ( .A(n11982), .B(n11981), .Z(n11977) );
  NANDN U272 ( .A(n12016), .B(n12015), .Z(n12011) );
  NANDN U273 ( .A(n12050), .B(n12049), .Z(n12045) );
  NANDN U274 ( .A(n12101), .B(n12100), .Z(n12096) );
  NANDN U275 ( .A(n12135), .B(n12134), .Z(n12130) );
  NANDN U276 ( .A(n12169), .B(n12168), .Z(n12164) );
  NANDN U277 ( .A(n12203), .B(n12202), .Z(n12198) );
  NANDN U278 ( .A(n12237), .B(n12236), .Z(n12232) );
  NANDN U279 ( .A(n12288), .B(n12287), .Z(n12283) );
  NANDN U280 ( .A(n12322), .B(n12321), .Z(n12317) );
  NANDN U281 ( .A(n12356), .B(n12355), .Z(n12351) );
  NANDN U282 ( .A(n12390), .B(n12389), .Z(n12385) );
  NANDN U283 ( .A(n12424), .B(n12423), .Z(n12419) );
  NANDN U284 ( .A(n12475), .B(n12474), .Z(n12470) );
  NANDN U285 ( .A(n12509), .B(n12508), .Z(n12504) );
  NANDN U286 ( .A(n12543), .B(n12542), .Z(n12538) );
  NANDN U287 ( .A(n12577), .B(n12576), .Z(n12572) );
  NANDN U288 ( .A(n12611), .B(n12610), .Z(n12606) );
  NANDN U289 ( .A(n12662), .B(n12661), .Z(n12657) );
  NANDN U290 ( .A(n12696), .B(n12695), .Z(n12691) );
  NANDN U291 ( .A(n12730), .B(n12729), .Z(n12725) );
  NANDN U292 ( .A(n12764), .B(n12763), .Z(n12759) );
  NANDN U293 ( .A(n12798), .B(n12797), .Z(n12793) );
  NANDN U294 ( .A(n12849), .B(n12848), .Z(n12844) );
  NANDN U295 ( .A(n12883), .B(n12882), .Z(n12878) );
  NANDN U296 ( .A(n12917), .B(n12916), .Z(n12912) );
  NANDN U297 ( .A(n12951), .B(n12950), .Z(n12946) );
  NANDN U298 ( .A(n12985), .B(n12984), .Z(n12980) );
  NANDN U299 ( .A(n13036), .B(n13035), .Z(n13031) );
  NANDN U300 ( .A(n13070), .B(n13069), .Z(n13065) );
  NANDN U301 ( .A(n13104), .B(n13103), .Z(n13099) );
  NANDN U302 ( .A(n13138), .B(n13137), .Z(n13133) );
  NANDN U303 ( .A(n13172), .B(n13171), .Z(n13167) );
  NANDN U304 ( .A(n13223), .B(n13222), .Z(n13218) );
  NANDN U305 ( .A(n13257), .B(n13256), .Z(n13252) );
  NANDN U306 ( .A(n13291), .B(n13290), .Z(n13286) );
  NANDN U307 ( .A(n13325), .B(n13324), .Z(n13320) );
  NANDN U308 ( .A(n13359), .B(n13358), .Z(n13354) );
  NANDN U309 ( .A(n13427), .B(n13426), .Z(n13422) );
  NANDN U310 ( .A(n13461), .B(n13460), .Z(n13456) );
  NANDN U311 ( .A(n13495), .B(n13494), .Z(n13490) );
  NANDN U312 ( .A(n13529), .B(n13528), .Z(n13524) );
  NANDN U313 ( .A(n13563), .B(n13562), .Z(n13558) );
  NANDN U314 ( .A(n13614), .B(n13613), .Z(n13609) );
  NANDN U315 ( .A(n13648), .B(n13647), .Z(n13643) );
  NANDN U316 ( .A(n13682), .B(n13681), .Z(n13677) );
  NANDN U317 ( .A(n13716), .B(n13715), .Z(n13711) );
  NANDN U318 ( .A(n13750), .B(n13749), .Z(n13745) );
  NANDN U319 ( .A(n13801), .B(n13800), .Z(n13796) );
  NANDN U320 ( .A(n13835), .B(n13834), .Z(n13830) );
  NANDN U321 ( .A(n13869), .B(n13868), .Z(n13864) );
  NANDN U322 ( .A(n13903), .B(n13902), .Z(n13898) );
  NANDN U323 ( .A(n13937), .B(n13936), .Z(n13932) );
  NANDN U324 ( .A(n13988), .B(n13987), .Z(n13983) );
  NANDN U325 ( .A(n14022), .B(n14021), .Z(n14017) );
  NANDN U326 ( .A(n14056), .B(n14055), .Z(n14051) );
  NANDN U327 ( .A(n14090), .B(n14089), .Z(n14085) );
  NANDN U328 ( .A(n14124), .B(n14123), .Z(n14119) );
  NANDN U329 ( .A(n14175), .B(n14174), .Z(n14170) );
  NANDN U330 ( .A(n14209), .B(n14208), .Z(n14204) );
  NANDN U331 ( .A(n14243), .B(n14242), .Z(n14238) );
  NANDN U332 ( .A(n14277), .B(n14276), .Z(n14272) );
  NANDN U333 ( .A(n14311), .B(n14310), .Z(n14306) );
  NANDN U334 ( .A(n14362), .B(n14361), .Z(n14357) );
  NANDN U335 ( .A(n14396), .B(n14395), .Z(n14391) );
  NANDN U336 ( .A(n14430), .B(n14429), .Z(n14425) );
  NANDN U337 ( .A(n14464), .B(n14463), .Z(n14459) );
  NANDN U338 ( .A(n14498), .B(n14497), .Z(n14493) );
  NANDN U339 ( .A(n14549), .B(n14548), .Z(n14544) );
  NANDN U340 ( .A(n14583), .B(n14582), .Z(n14578) );
  NANDN U341 ( .A(n14617), .B(n14616), .Z(n14612) );
  NANDN U342 ( .A(n14651), .B(n14650), .Z(n14646) );
  NANDN U343 ( .A(n14685), .B(n14684), .Z(n14680) );
  NANDN U344 ( .A(n14736), .B(n14735), .Z(n14731) );
  NANDN U345 ( .A(n14770), .B(n14769), .Z(n14765) );
  NANDN U346 ( .A(n14804), .B(n14803), .Z(n14799) );
  NANDN U347 ( .A(n14838), .B(n14837), .Z(n14833) );
  NANDN U348 ( .A(n14872), .B(n14871), .Z(n14867) );
  NANDN U349 ( .A(n14923), .B(n14922), .Z(n14918) );
  NANDN U350 ( .A(n14957), .B(n14956), .Z(n14952) );
  NANDN U351 ( .A(n14991), .B(n14990), .Z(n14986) );
  NANDN U352 ( .A(n15025), .B(n15024), .Z(n15020) );
  NANDN U353 ( .A(n15059), .B(n15058), .Z(n15054) );
  NANDN U354 ( .A(n15110), .B(n15109), .Z(n15105) );
  NANDN U355 ( .A(n15144), .B(n15143), .Z(n15139) );
  NANDN U356 ( .A(n15178), .B(n15177), .Z(n15173) );
  NANDN U357 ( .A(n15212), .B(n15211), .Z(n15207) );
  NANDN U358 ( .A(n15246), .B(n15245), .Z(n15241) );
  NANDN U359 ( .A(n15314), .B(n15313), .Z(n15309) );
  NANDN U360 ( .A(n15348), .B(n15347), .Z(n15343) );
  NANDN U361 ( .A(n15382), .B(n15381), .Z(n15377) );
  NANDN U362 ( .A(n15416), .B(n15415), .Z(n15411) );
  NANDN U363 ( .A(n15450), .B(n15449), .Z(n15445) );
  NANDN U364 ( .A(n15501), .B(n15500), .Z(n15496) );
  NANDN U365 ( .A(n15535), .B(n15534), .Z(n15530) );
  NANDN U366 ( .A(n15569), .B(n15568), .Z(n15564) );
  NANDN U367 ( .A(n15603), .B(n15602), .Z(n15598) );
  NANDN U368 ( .A(n15637), .B(n15636), .Z(n15632) );
  NANDN U369 ( .A(n15688), .B(n15687), .Z(n15683) );
  NANDN U370 ( .A(n15722), .B(n15721), .Z(n15717) );
  NANDN U371 ( .A(n15756), .B(n15755), .Z(n15751) );
  NANDN U372 ( .A(n15790), .B(n15789), .Z(n15785) );
  NANDN U373 ( .A(n15824), .B(n15823), .Z(n15819) );
  NANDN U374 ( .A(n15875), .B(n15874), .Z(n15870) );
  NANDN U375 ( .A(n15909), .B(n15908), .Z(n15904) );
  NANDN U376 ( .A(n15943), .B(n15942), .Z(n15938) );
  NANDN U377 ( .A(n15977), .B(n15976), .Z(n15972) );
  NANDN U378 ( .A(n16011), .B(n16010), .Z(n16006) );
  NANDN U379 ( .A(n16062), .B(n16061), .Z(n16057) );
  NANDN U380 ( .A(n16096), .B(n16095), .Z(n16091) );
  NANDN U381 ( .A(n16130), .B(n16129), .Z(n16125) );
  NANDN U382 ( .A(n16164), .B(n16163), .Z(n16159) );
  NANDN U383 ( .A(n16198), .B(n16197), .Z(n16193) );
  NANDN U384 ( .A(n16249), .B(n16248), .Z(n16244) );
  NANDN U385 ( .A(n16283), .B(n16282), .Z(n16278) );
  NANDN U386 ( .A(n16317), .B(n16316), .Z(n16312) );
  NANDN U387 ( .A(n16351), .B(n16350), .Z(n16346) );
  NANDN U388 ( .A(n16385), .B(n16384), .Z(n16380) );
  NANDN U389 ( .A(n16436), .B(n16435), .Z(n16431) );
  NANDN U390 ( .A(n16470), .B(n16469), .Z(n16465) );
  NANDN U391 ( .A(n16504), .B(n16503), .Z(n16499) );
  NANDN U392 ( .A(n16538), .B(n16537), .Z(n16533) );
  NANDN U393 ( .A(n16572), .B(n16571), .Z(n16567) );
  NANDN U394 ( .A(n16623), .B(n16622), .Z(n16618) );
  NANDN U395 ( .A(n16657), .B(n16656), .Z(n16652) );
  NANDN U396 ( .A(n16691), .B(n16690), .Z(n16686) );
  NANDN U397 ( .A(n16725), .B(n16724), .Z(n16720) );
  NANDN U398 ( .A(n16759), .B(n16758), .Z(n16754) );
  NANDN U399 ( .A(n16810), .B(n16809), .Z(n16805) );
  NANDN U400 ( .A(n16844), .B(n16843), .Z(n16839) );
  NANDN U401 ( .A(n16878), .B(n16877), .Z(n16873) );
  NANDN U402 ( .A(n16912), .B(n16911), .Z(n16907) );
  NANDN U403 ( .A(n16946), .B(n16945), .Z(n16941) );
  NANDN U404 ( .A(n16997), .B(n16996), .Z(n16992) );
  NANDN U405 ( .A(n17031), .B(n17030), .Z(n17026) );
  NANDN U406 ( .A(n17065), .B(n17064), .Z(n17060) );
  NANDN U407 ( .A(n17099), .B(n17098), .Z(n17094) );
  NANDN U408 ( .A(n17133), .B(n17132), .Z(n17128) );
  NANDN U409 ( .A(n17195), .B(n17194), .Z(n17190) );
  NANDN U410 ( .A(n17229), .B(n17228), .Z(n17224) );
  NANDN U411 ( .A(n17263), .B(n17262), .Z(n17258) );
  NANDN U412 ( .A(n17297), .B(n17296), .Z(n17292) );
  NANDN U413 ( .A(n17331), .B(n17330), .Z(n17326) );
  NANDN U414 ( .A(n17382), .B(n17381), .Z(n17377) );
  NANDN U415 ( .A(n17416), .B(n17415), .Z(n17411) );
  NANDN U416 ( .A(n17450), .B(n17449), .Z(n17445) );
  NANDN U417 ( .A(n17484), .B(n17483), .Z(n17479) );
  NANDN U418 ( .A(n17518), .B(n17517), .Z(n17513) );
  NANDN U419 ( .A(n17569), .B(n17568), .Z(n17564) );
  NANDN U420 ( .A(n17603), .B(n17602), .Z(n17598) );
  NANDN U421 ( .A(n17637), .B(n17636), .Z(n17632) );
  NANDN U422 ( .A(n17671), .B(n17670), .Z(n17666) );
  NANDN U423 ( .A(n17705), .B(n17704), .Z(n17700) );
  NANDN U424 ( .A(n17756), .B(n17755), .Z(n17751) );
  NANDN U425 ( .A(n17790), .B(n17789), .Z(n17785) );
  NANDN U426 ( .A(n17824), .B(n17823), .Z(n17819) );
  NANDN U427 ( .A(n17858), .B(n17857), .Z(n17853) );
  NANDN U428 ( .A(n17892), .B(n17891), .Z(n17887) );
  NANDN U429 ( .A(n17943), .B(n17942), .Z(n17938) );
  NANDN U430 ( .A(n17977), .B(n17976), .Z(n17972) );
  NANDN U431 ( .A(n18011), .B(n18010), .Z(n18006) );
  NANDN U432 ( .A(n18045), .B(n18044), .Z(n18040) );
  NANDN U433 ( .A(n18079), .B(n18078), .Z(n18074) );
  NANDN U434 ( .A(n18130), .B(n18129), .Z(n18125) );
  NANDN U435 ( .A(n18164), .B(n18163), .Z(n18159) );
  NANDN U436 ( .A(n18198), .B(n18197), .Z(n18193) );
  NANDN U437 ( .A(n18232), .B(n18231), .Z(n18227) );
  NANDN U438 ( .A(n18266), .B(n18265), .Z(n18261) );
  NANDN U439 ( .A(n18317), .B(n18316), .Z(n18312) );
  NANDN U440 ( .A(n18351), .B(n18350), .Z(n18346) );
  NANDN U441 ( .A(n18385), .B(n18384), .Z(n18380) );
  NANDN U442 ( .A(n18419), .B(n18418), .Z(n18414) );
  NANDN U443 ( .A(n18453), .B(n18452), .Z(n18448) );
  NANDN U444 ( .A(n18504), .B(n18503), .Z(n18499) );
  NANDN U445 ( .A(n18538), .B(n18537), .Z(n18533) );
  NANDN U446 ( .A(n18572), .B(n18571), .Z(n18567) );
  NANDN U447 ( .A(n18606), .B(n18605), .Z(n18601) );
  NANDN U448 ( .A(n18640), .B(n18639), .Z(n18635) );
  NANDN U449 ( .A(n18691), .B(n18690), .Z(n18686) );
  NANDN U450 ( .A(n18725), .B(n18724), .Z(n18720) );
  NANDN U451 ( .A(n18759), .B(n18758), .Z(n18754) );
  NANDN U452 ( .A(n18793), .B(n18792), .Z(n18788) );
  NANDN U453 ( .A(n18827), .B(n18826), .Z(n18822) );
  NANDN U454 ( .A(n18887), .B(n18886), .Z(n18882) );
  NANDN U455 ( .A(n18921), .B(n18920), .Z(n18916) );
  NANDN U456 ( .A(n18955), .B(n18954), .Z(n18950) );
  NANDN U457 ( .A(n18989), .B(n18988), .Z(n18984) );
  NANDN U458 ( .A(n2633), .B(n2632), .Z(n2628) );
  NANDN U459 ( .A(n3007), .B(n3006), .Z(n3002) );
  NANDN U460 ( .A(n3381), .B(n3380), .Z(n3376) );
  NANDN U461 ( .A(n3755), .B(n3754), .Z(n3750) );
  NANDN U462 ( .A(n4144), .B(n4143), .Z(n4139) );
  NANDN U463 ( .A(n4518), .B(n4517), .Z(n4513) );
  NANDN U464 ( .A(n4892), .B(n4891), .Z(n4887) );
  NANDN U465 ( .A(n5266), .B(n5265), .Z(n5261) );
  NANDN U466 ( .A(n5640), .B(n5639), .Z(n5635) );
  NANDN U467 ( .A(n6032), .B(n6031), .Z(n6027) );
  NANDN U468 ( .A(n6406), .B(n6405), .Z(n6401) );
  NANDN U469 ( .A(n6780), .B(n6779), .Z(n6775) );
  NANDN U470 ( .A(n7154), .B(n7153), .Z(n7149) );
  NANDN U471 ( .A(n7528), .B(n7527), .Z(n7523) );
  NANDN U472 ( .A(n7919), .B(n7918), .Z(n7914) );
  NANDN U473 ( .A(n8293), .B(n8292), .Z(n8288) );
  NANDN U474 ( .A(n8667), .B(n8666), .Z(n8662) );
  NANDN U475 ( .A(n9041), .B(n9040), .Z(n9036) );
  NANDN U476 ( .A(n9415), .B(n9414), .Z(n9410) );
  NANDN U477 ( .A(n9806), .B(n9805), .Z(n9801) );
  NANDN U478 ( .A(n10180), .B(n10179), .Z(n10175) );
  NANDN U479 ( .A(n10554), .B(n10553), .Z(n10549) );
  NANDN U480 ( .A(n10928), .B(n10927), .Z(n10923) );
  NANDN U481 ( .A(n11302), .B(n11301), .Z(n11297) );
  NANDN U482 ( .A(n11693), .B(n11692), .Z(n11688) );
  NANDN U483 ( .A(n12067), .B(n12066), .Z(n12062) );
  NANDN U484 ( .A(n12441), .B(n12440), .Z(n12436) );
  NANDN U485 ( .A(n12815), .B(n12814), .Z(n12810) );
  NANDN U486 ( .A(n13189), .B(n13188), .Z(n13184) );
  NANDN U487 ( .A(n13580), .B(n13579), .Z(n13575) );
  NANDN U488 ( .A(n13954), .B(n13953), .Z(n13949) );
  NANDN U489 ( .A(n14328), .B(n14327), .Z(n14323) );
  NANDN U490 ( .A(n14702), .B(n14701), .Z(n14697) );
  NANDN U491 ( .A(n15076), .B(n15075), .Z(n15071) );
  NANDN U492 ( .A(n15467), .B(n15466), .Z(n15462) );
  NANDN U493 ( .A(n15841), .B(n15840), .Z(n15836) );
  NANDN U494 ( .A(n16215), .B(n16214), .Z(n16210) );
  NANDN U495 ( .A(n16589), .B(n16588), .Z(n16584) );
  NANDN U496 ( .A(n16963), .B(n16962), .Z(n16958) );
  NANDN U497 ( .A(n17348), .B(n17347), .Z(n17343) );
  NANDN U498 ( .A(n17722), .B(n17721), .Z(n17717) );
  NANDN U499 ( .A(n18096), .B(n18095), .Z(n18091) );
  NANDN U500 ( .A(n18470), .B(n18469), .Z(n18465) );
  NANDN U501 ( .A(n9602), .B(n9601), .Z(n9597) );
  NANDN U502 ( .A(n19108), .B(n19107), .Z(n19103) );
  NANDN U503 ( .A(n13376), .B(n13375), .Z(n13371) );
  NANDN U504 ( .A(n19057), .B(n19056), .Z(n19052) );
  NANDN U505 ( .A(n19024), .B(n19023), .Z(n19019) );
  NANDN U506 ( .A(n19125), .B(n19124), .Z(n19120) );
  NANDN U507 ( .A(n19159), .B(n19158), .Z(n19154) );
  NANDN U508 ( .A(n19193), .B(n19192), .Z(n19188) );
  NANDN U509 ( .A(n19227), .B(n19226), .Z(n19222) );
  NANDN U510 ( .A(n19287), .B(n19286), .Z(n19282) );
  NANDN U511 ( .A(n19321), .B(n19320), .Z(n19316) );
  NANDN U512 ( .A(n19355), .B(n19354), .Z(n19350) );
  NANDN U513 ( .A(n19389), .B(n19388), .Z(n19384) );
  NANDN U514 ( .A(n19423), .B(n19422), .Z(n19418) );
  NANDN U515 ( .A(n2123), .B(n2122), .Z(n2118) );
  NANDN U516 ( .A(n2158), .B(n2157), .Z(n2153) );
  NANDN U517 ( .A(n2192), .B(n2191), .Z(n2187) );
  NANDN U518 ( .A(n2226), .B(n2225), .Z(n2221) );
  NANDN U519 ( .A(n2275), .B(n2274), .Z(n2270) );
  NANDN U520 ( .A(n2309), .B(n2308), .Z(n2304) );
  NANDN U521 ( .A(n2343), .B(n2342), .Z(n2338) );
  NANDN U522 ( .A(n2377), .B(n2376), .Z(n2372) );
  NANDN U523 ( .A(n2411), .B(n2410), .Z(n2406) );
  NANDN U524 ( .A(n2463), .B(n2462), .Z(n2458) );
  NANDN U525 ( .A(n2497), .B(n2496), .Z(n2492) );
  NANDN U526 ( .A(n2531), .B(n2530), .Z(n2526) );
  NANDN U527 ( .A(n2565), .B(n2564), .Z(n2560) );
  NANDN U528 ( .A(n2599), .B(n2598), .Z(n2594) );
  NANDN U529 ( .A(n2650), .B(n2649), .Z(n2645) );
  NANDN U530 ( .A(n2684), .B(n2683), .Z(n2679) );
  NANDN U531 ( .A(n2718), .B(n2717), .Z(n2713) );
  NANDN U532 ( .A(n2752), .B(n2751), .Z(n2747) );
  NANDN U533 ( .A(n2786), .B(n2785), .Z(n2781) );
  NANDN U534 ( .A(n2837), .B(n2836), .Z(n2832) );
  NANDN U535 ( .A(n2871), .B(n2870), .Z(n2866) );
  NANDN U536 ( .A(n2905), .B(n2904), .Z(n2900) );
  NANDN U537 ( .A(n2939), .B(n2938), .Z(n2934) );
  NANDN U538 ( .A(n2973), .B(n2972), .Z(n2968) );
  NANDN U539 ( .A(n3024), .B(n3023), .Z(n3019) );
  NANDN U540 ( .A(n3058), .B(n3057), .Z(n3053) );
  NANDN U541 ( .A(n3092), .B(n3091), .Z(n3087) );
  NANDN U542 ( .A(n3126), .B(n3125), .Z(n3121) );
  NANDN U543 ( .A(n3160), .B(n3159), .Z(n3155) );
  NANDN U544 ( .A(n3211), .B(n3210), .Z(n3206) );
  NANDN U545 ( .A(n3245), .B(n3244), .Z(n3240) );
  NANDN U546 ( .A(n3279), .B(n3278), .Z(n3274) );
  NANDN U547 ( .A(n3313), .B(n3312), .Z(n3308) );
  NANDN U548 ( .A(n3347), .B(n3346), .Z(n3342) );
  NANDN U549 ( .A(n3398), .B(n3397), .Z(n3393) );
  NANDN U550 ( .A(n3432), .B(n3431), .Z(n3427) );
  NANDN U551 ( .A(n3466), .B(n3465), .Z(n3461) );
  NANDN U552 ( .A(n3500), .B(n3499), .Z(n3495) );
  NANDN U553 ( .A(n3534), .B(n3533), .Z(n3529) );
  NANDN U554 ( .A(n3585), .B(n3584), .Z(n3580) );
  NANDN U555 ( .A(n3619), .B(n3618), .Z(n3614) );
  NANDN U556 ( .A(n3653), .B(n3652), .Z(n3648) );
  NANDN U557 ( .A(n3687), .B(n3686), .Z(n3682) );
  NANDN U558 ( .A(n3721), .B(n3720), .Z(n3716) );
  NANDN U559 ( .A(n3772), .B(n3771), .Z(n3767) );
  NANDN U560 ( .A(n3806), .B(n3805), .Z(n3801) );
  NANDN U561 ( .A(n3840), .B(n3839), .Z(n3835) );
  NANDN U562 ( .A(n3874), .B(n3873), .Z(n3869) );
  NANDN U563 ( .A(n3908), .B(n3907), .Z(n3903) );
  NANDN U564 ( .A(n3974), .B(n3973), .Z(n3969) );
  NANDN U565 ( .A(n4008), .B(n4007), .Z(n4003) );
  NANDN U566 ( .A(n4042), .B(n4041), .Z(n4037) );
  NANDN U567 ( .A(n4076), .B(n4075), .Z(n4071) );
  NANDN U568 ( .A(n4110), .B(n4109), .Z(n4105) );
  NANDN U569 ( .A(n4161), .B(n4160), .Z(n4156) );
  NANDN U570 ( .A(n4195), .B(n4194), .Z(n4190) );
  NANDN U571 ( .A(n4229), .B(n4228), .Z(n4224) );
  NANDN U572 ( .A(n4263), .B(n4262), .Z(n4258) );
  NANDN U573 ( .A(n4297), .B(n4296), .Z(n4292) );
  NANDN U574 ( .A(n4348), .B(n4347), .Z(n4343) );
  NANDN U575 ( .A(n4382), .B(n4381), .Z(n4377) );
  NANDN U576 ( .A(n4416), .B(n4415), .Z(n4411) );
  NANDN U577 ( .A(n4450), .B(n4449), .Z(n4445) );
  NANDN U578 ( .A(n4484), .B(n4483), .Z(n4479) );
  NANDN U579 ( .A(n4535), .B(n4534), .Z(n4530) );
  NANDN U580 ( .A(n4569), .B(n4568), .Z(n4564) );
  NANDN U581 ( .A(n4603), .B(n4602), .Z(n4598) );
  NANDN U582 ( .A(n4637), .B(n4636), .Z(n4632) );
  NANDN U583 ( .A(n4671), .B(n4670), .Z(n4666) );
  NANDN U584 ( .A(n4722), .B(n4721), .Z(n4717) );
  NANDN U585 ( .A(n4756), .B(n4755), .Z(n4751) );
  NANDN U586 ( .A(n4790), .B(n4789), .Z(n4785) );
  NANDN U587 ( .A(n4824), .B(n4823), .Z(n4819) );
  NANDN U588 ( .A(n4858), .B(n4857), .Z(n4853) );
  NANDN U589 ( .A(n4909), .B(n4908), .Z(n4904) );
  NANDN U590 ( .A(n4943), .B(n4942), .Z(n4938) );
  NANDN U591 ( .A(n4977), .B(n4976), .Z(n4972) );
  NANDN U592 ( .A(n5011), .B(n5010), .Z(n5006) );
  NANDN U593 ( .A(n5045), .B(n5044), .Z(n5040) );
  NANDN U594 ( .A(n5096), .B(n5095), .Z(n5091) );
  NANDN U595 ( .A(n5130), .B(n5129), .Z(n5125) );
  NANDN U596 ( .A(n5164), .B(n5163), .Z(n5159) );
  NANDN U597 ( .A(n5198), .B(n5197), .Z(n5193) );
  NANDN U598 ( .A(n5232), .B(n5231), .Z(n5227) );
  NANDN U599 ( .A(n5283), .B(n5282), .Z(n5278) );
  NANDN U600 ( .A(n5317), .B(n5316), .Z(n5312) );
  NANDN U601 ( .A(n5351), .B(n5350), .Z(n5346) );
  NANDN U602 ( .A(n5385), .B(n5384), .Z(n5380) );
  NANDN U603 ( .A(n5419), .B(n5418), .Z(n5414) );
  NANDN U604 ( .A(n5470), .B(n5469), .Z(n5465) );
  NANDN U605 ( .A(n5504), .B(n5503), .Z(n5499) );
  NANDN U606 ( .A(n5538), .B(n5537), .Z(n5533) );
  NANDN U607 ( .A(n5572), .B(n5571), .Z(n5567) );
  NANDN U608 ( .A(n5606), .B(n5605), .Z(n5601) );
  NANDN U609 ( .A(n5657), .B(n5656), .Z(n5652) );
  NANDN U610 ( .A(n5691), .B(n5690), .Z(n5686) );
  NANDN U611 ( .A(n5725), .B(n5724), .Z(n5720) );
  NANDN U612 ( .A(n5759), .B(n5758), .Z(n5754) );
  NANDN U613 ( .A(n5793), .B(n5792), .Z(n5788) );
  NANDN U614 ( .A(n5862), .B(n5861), .Z(n5857) );
  NANDN U615 ( .A(n5896), .B(n5895), .Z(n5891) );
  NANDN U616 ( .A(n5930), .B(n5929), .Z(n5925) );
  NANDN U617 ( .A(n5964), .B(n5963), .Z(n5959) );
  NANDN U618 ( .A(n5998), .B(n5997), .Z(n5993) );
  NANDN U619 ( .A(n6049), .B(n6048), .Z(n6044) );
  NANDN U620 ( .A(n6083), .B(n6082), .Z(n6078) );
  NANDN U621 ( .A(n6117), .B(n6116), .Z(n6112) );
  NANDN U622 ( .A(n6151), .B(n6150), .Z(n6146) );
  NANDN U623 ( .A(n6185), .B(n6184), .Z(n6180) );
  NANDN U624 ( .A(n6236), .B(n6235), .Z(n6231) );
  NANDN U625 ( .A(n6270), .B(n6269), .Z(n6265) );
  NANDN U626 ( .A(n6304), .B(n6303), .Z(n6299) );
  NANDN U627 ( .A(n6338), .B(n6337), .Z(n6333) );
  NANDN U628 ( .A(n6372), .B(n6371), .Z(n6367) );
  NANDN U629 ( .A(n6423), .B(n6422), .Z(n6418) );
  NANDN U630 ( .A(n6457), .B(n6456), .Z(n6452) );
  NANDN U631 ( .A(n6491), .B(n6490), .Z(n6486) );
  NANDN U632 ( .A(n6525), .B(n6524), .Z(n6520) );
  NANDN U633 ( .A(n6559), .B(n6558), .Z(n6554) );
  NANDN U634 ( .A(n6610), .B(n6609), .Z(n6605) );
  NANDN U635 ( .A(n6644), .B(n6643), .Z(n6639) );
  NANDN U636 ( .A(n6678), .B(n6677), .Z(n6673) );
  NANDN U637 ( .A(n6712), .B(n6711), .Z(n6707) );
  NANDN U638 ( .A(n6746), .B(n6745), .Z(n6741) );
  NANDN U639 ( .A(n6797), .B(n6796), .Z(n6792) );
  NANDN U640 ( .A(n6831), .B(n6830), .Z(n6826) );
  NANDN U641 ( .A(n6865), .B(n6864), .Z(n6860) );
  NANDN U642 ( .A(n6899), .B(n6898), .Z(n6894) );
  NANDN U643 ( .A(n6933), .B(n6932), .Z(n6928) );
  NANDN U644 ( .A(n6984), .B(n6983), .Z(n6979) );
  NANDN U645 ( .A(n7018), .B(n7017), .Z(n7013) );
  NANDN U646 ( .A(n7052), .B(n7051), .Z(n7047) );
  NANDN U647 ( .A(n7086), .B(n7085), .Z(n7081) );
  NANDN U648 ( .A(n7120), .B(n7119), .Z(n7115) );
  NANDN U649 ( .A(n7171), .B(n7170), .Z(n7166) );
  NANDN U650 ( .A(n7205), .B(n7204), .Z(n7200) );
  NANDN U651 ( .A(n7239), .B(n7238), .Z(n7234) );
  NANDN U652 ( .A(n7273), .B(n7272), .Z(n7268) );
  NANDN U653 ( .A(n7307), .B(n7306), .Z(n7302) );
  NANDN U654 ( .A(n7358), .B(n7357), .Z(n7353) );
  NANDN U655 ( .A(n7392), .B(n7391), .Z(n7387) );
  NANDN U656 ( .A(n7426), .B(n7425), .Z(n7421) );
  NANDN U657 ( .A(n7460), .B(n7459), .Z(n7455) );
  NANDN U658 ( .A(n7494), .B(n7493), .Z(n7489) );
  NANDN U659 ( .A(n7545), .B(n7544), .Z(n7540) );
  NANDN U660 ( .A(n7579), .B(n7578), .Z(n7574) );
  NANDN U661 ( .A(n7613), .B(n7612), .Z(n7608) );
  NANDN U662 ( .A(n7647), .B(n7646), .Z(n7642) );
  NANDN U663 ( .A(n7681), .B(n7680), .Z(n7676) );
  NANDN U664 ( .A(n7749), .B(n7748), .Z(n7744) );
  NANDN U665 ( .A(n7783), .B(n7782), .Z(n7778) );
  NANDN U666 ( .A(n7817), .B(n7816), .Z(n7812) );
  NANDN U667 ( .A(n7851), .B(n7850), .Z(n7846) );
  NANDN U668 ( .A(n7885), .B(n7884), .Z(n7880) );
  NANDN U669 ( .A(n7936), .B(n7935), .Z(n7931) );
  NANDN U670 ( .A(n7970), .B(n7969), .Z(n7965) );
  NANDN U671 ( .A(n8004), .B(n8003), .Z(n7999) );
  NANDN U672 ( .A(n8038), .B(n8037), .Z(n8033) );
  NANDN U673 ( .A(n8072), .B(n8071), .Z(n8067) );
  NANDN U674 ( .A(n8123), .B(n8122), .Z(n8118) );
  NANDN U675 ( .A(n8157), .B(n8156), .Z(n8152) );
  NANDN U676 ( .A(n8191), .B(n8190), .Z(n8186) );
  NANDN U677 ( .A(n8225), .B(n8224), .Z(n8220) );
  NANDN U678 ( .A(n8259), .B(n8258), .Z(n8254) );
  NANDN U679 ( .A(n8310), .B(n8309), .Z(n8305) );
  NANDN U680 ( .A(n8344), .B(n8343), .Z(n8339) );
  NANDN U681 ( .A(n8378), .B(n8377), .Z(n8373) );
  NANDN U682 ( .A(n8412), .B(n8411), .Z(n8407) );
  NANDN U683 ( .A(n8446), .B(n8445), .Z(n8441) );
  NANDN U684 ( .A(n8497), .B(n8496), .Z(n8492) );
  NANDN U685 ( .A(n8531), .B(n8530), .Z(n8526) );
  NANDN U686 ( .A(n8565), .B(n8564), .Z(n8560) );
  NANDN U687 ( .A(n8599), .B(n8598), .Z(n8594) );
  NANDN U688 ( .A(n8633), .B(n8632), .Z(n8628) );
  NANDN U689 ( .A(n8684), .B(n8683), .Z(n8679) );
  NANDN U690 ( .A(n8718), .B(n8717), .Z(n8713) );
  NANDN U691 ( .A(n8752), .B(n8751), .Z(n8747) );
  NANDN U692 ( .A(n8786), .B(n8785), .Z(n8781) );
  NANDN U693 ( .A(n8820), .B(n8819), .Z(n8815) );
  NANDN U694 ( .A(n8871), .B(n8870), .Z(n8866) );
  NANDN U695 ( .A(n8905), .B(n8904), .Z(n8900) );
  NANDN U696 ( .A(n8939), .B(n8938), .Z(n8934) );
  NANDN U697 ( .A(n8973), .B(n8972), .Z(n8968) );
  NANDN U698 ( .A(n9007), .B(n9006), .Z(n9002) );
  NANDN U699 ( .A(n9058), .B(n9057), .Z(n9053) );
  NANDN U700 ( .A(n9092), .B(n9091), .Z(n9087) );
  NANDN U701 ( .A(n9126), .B(n9125), .Z(n9121) );
  NANDN U702 ( .A(n9160), .B(n9159), .Z(n9155) );
  NANDN U703 ( .A(n9194), .B(n9193), .Z(n9189) );
  NANDN U704 ( .A(n9245), .B(n9244), .Z(n9240) );
  NANDN U705 ( .A(n9279), .B(n9278), .Z(n9274) );
  NANDN U706 ( .A(n9313), .B(n9312), .Z(n9308) );
  NANDN U707 ( .A(n9347), .B(n9346), .Z(n9342) );
  NANDN U708 ( .A(n9381), .B(n9380), .Z(n9376) );
  NANDN U709 ( .A(n9432), .B(n9431), .Z(n9427) );
  NANDN U710 ( .A(n9466), .B(n9465), .Z(n9461) );
  NANDN U711 ( .A(n9500), .B(n9499), .Z(n9495) );
  NANDN U712 ( .A(n9534), .B(n9533), .Z(n9529) );
  NANDN U713 ( .A(n9568), .B(n9567), .Z(n9563) );
  NANDN U714 ( .A(n9636), .B(n9635), .Z(n9631) );
  NANDN U715 ( .A(n9670), .B(n9669), .Z(n9665) );
  NANDN U716 ( .A(n9704), .B(n9703), .Z(n9699) );
  NANDN U717 ( .A(n9738), .B(n9737), .Z(n9733) );
  NANDN U718 ( .A(n9772), .B(n9771), .Z(n9767) );
  NANDN U719 ( .A(n9823), .B(n9822), .Z(n9818) );
  NANDN U720 ( .A(n9857), .B(n9856), .Z(n9852) );
  NANDN U721 ( .A(n9891), .B(n9890), .Z(n9886) );
  NANDN U722 ( .A(n9925), .B(n9924), .Z(n9920) );
  NANDN U723 ( .A(n9959), .B(n9958), .Z(n9954) );
  NANDN U724 ( .A(n10010), .B(n10009), .Z(n10005) );
  NANDN U725 ( .A(n10044), .B(n10043), .Z(n10039) );
  NANDN U726 ( .A(n10078), .B(n10077), .Z(n10073) );
  NANDN U727 ( .A(n10112), .B(n10111), .Z(n10107) );
  NANDN U728 ( .A(n10146), .B(n10145), .Z(n10141) );
  NANDN U729 ( .A(n10197), .B(n10196), .Z(n10192) );
  NANDN U730 ( .A(n10231), .B(n10230), .Z(n10226) );
  NANDN U731 ( .A(n10265), .B(n10264), .Z(n10260) );
  NANDN U732 ( .A(n10299), .B(n10298), .Z(n10294) );
  NANDN U733 ( .A(n10333), .B(n10332), .Z(n10328) );
  NANDN U734 ( .A(n10384), .B(n10383), .Z(n10379) );
  NANDN U735 ( .A(n10418), .B(n10417), .Z(n10413) );
  NANDN U736 ( .A(n10452), .B(n10451), .Z(n10447) );
  NANDN U737 ( .A(n10486), .B(n10485), .Z(n10481) );
  NANDN U738 ( .A(n10520), .B(n10519), .Z(n10515) );
  NANDN U739 ( .A(n10571), .B(n10570), .Z(n10566) );
  NANDN U740 ( .A(n10605), .B(n10604), .Z(n10600) );
  NANDN U741 ( .A(n10639), .B(n10638), .Z(n10634) );
  NANDN U742 ( .A(n10673), .B(n10672), .Z(n10668) );
  NANDN U743 ( .A(n10707), .B(n10706), .Z(n10702) );
  NANDN U744 ( .A(n10758), .B(n10757), .Z(n10753) );
  NANDN U745 ( .A(n10792), .B(n10791), .Z(n10787) );
  NANDN U746 ( .A(n10826), .B(n10825), .Z(n10821) );
  NANDN U747 ( .A(n10860), .B(n10859), .Z(n10855) );
  NANDN U748 ( .A(n10894), .B(n10893), .Z(n10889) );
  NANDN U749 ( .A(n10945), .B(n10944), .Z(n10940) );
  NANDN U750 ( .A(n10979), .B(n10978), .Z(n10974) );
  NANDN U751 ( .A(n11013), .B(n11012), .Z(n11008) );
  NANDN U752 ( .A(n11047), .B(n11046), .Z(n11042) );
  NANDN U753 ( .A(n11081), .B(n11080), .Z(n11076) );
  NANDN U754 ( .A(n11132), .B(n11131), .Z(n11127) );
  NANDN U755 ( .A(n11166), .B(n11165), .Z(n11161) );
  NANDN U756 ( .A(n11200), .B(n11199), .Z(n11195) );
  NANDN U757 ( .A(n11234), .B(n11233), .Z(n11229) );
  NANDN U758 ( .A(n11268), .B(n11267), .Z(n11263) );
  NANDN U759 ( .A(n11319), .B(n11318), .Z(n11314) );
  NANDN U760 ( .A(n11353), .B(n11352), .Z(n11348) );
  NANDN U761 ( .A(n11387), .B(n11386), .Z(n11382) );
  NANDN U762 ( .A(n11421), .B(n11420), .Z(n11416) );
  NANDN U763 ( .A(n11455), .B(n11454), .Z(n11450) );
  NANDN U764 ( .A(n11523), .B(n11522), .Z(n11518) );
  NANDN U765 ( .A(n11557), .B(n11556), .Z(n11552) );
  NANDN U766 ( .A(n11591), .B(n11590), .Z(n11586) );
  NANDN U767 ( .A(n11625), .B(n11624), .Z(n11620) );
  NANDN U768 ( .A(n11659), .B(n11658), .Z(n11654) );
  NANDN U769 ( .A(n11710), .B(n11709), .Z(n11705) );
  NANDN U770 ( .A(n11744), .B(n11743), .Z(n11739) );
  NANDN U771 ( .A(n11778), .B(n11777), .Z(n11773) );
  NANDN U772 ( .A(n11812), .B(n11811), .Z(n11807) );
  NANDN U773 ( .A(n11846), .B(n11845), .Z(n11841) );
  NANDN U774 ( .A(n11897), .B(n11896), .Z(n11892) );
  NANDN U775 ( .A(n11931), .B(n11930), .Z(n11926) );
  NANDN U776 ( .A(n11965), .B(n11964), .Z(n11960) );
  NANDN U777 ( .A(n11999), .B(n11998), .Z(n11994) );
  NANDN U778 ( .A(n12033), .B(n12032), .Z(n12028) );
  NANDN U779 ( .A(n12084), .B(n12083), .Z(n12079) );
  NANDN U780 ( .A(n12118), .B(n12117), .Z(n12113) );
  NANDN U781 ( .A(n12152), .B(n12151), .Z(n12147) );
  NANDN U782 ( .A(n12186), .B(n12185), .Z(n12181) );
  NANDN U783 ( .A(n12220), .B(n12219), .Z(n12215) );
  NANDN U784 ( .A(n12271), .B(n12270), .Z(n12266) );
  NANDN U785 ( .A(n12305), .B(n12304), .Z(n12300) );
  NANDN U786 ( .A(n12339), .B(n12338), .Z(n12334) );
  NANDN U787 ( .A(n12373), .B(n12372), .Z(n12368) );
  NANDN U788 ( .A(n12407), .B(n12406), .Z(n12402) );
  NANDN U789 ( .A(n12458), .B(n12457), .Z(n12453) );
  NANDN U790 ( .A(n12492), .B(n12491), .Z(n12487) );
  NANDN U791 ( .A(n12526), .B(n12525), .Z(n12521) );
  NANDN U792 ( .A(n12560), .B(n12559), .Z(n12555) );
  NANDN U793 ( .A(n12594), .B(n12593), .Z(n12589) );
  NANDN U794 ( .A(n12645), .B(n12644), .Z(n12640) );
  NANDN U795 ( .A(n12679), .B(n12678), .Z(n12674) );
  NANDN U796 ( .A(n12713), .B(n12712), .Z(n12708) );
  NANDN U797 ( .A(n12747), .B(n12746), .Z(n12742) );
  NANDN U798 ( .A(n12781), .B(n12780), .Z(n12776) );
  NANDN U799 ( .A(n12832), .B(n12831), .Z(n12827) );
  NANDN U800 ( .A(n12866), .B(n12865), .Z(n12861) );
  NANDN U801 ( .A(n12900), .B(n12899), .Z(n12895) );
  NANDN U802 ( .A(n12934), .B(n12933), .Z(n12929) );
  NANDN U803 ( .A(n12968), .B(n12967), .Z(n12963) );
  NANDN U804 ( .A(n13019), .B(n13018), .Z(n13014) );
  NANDN U805 ( .A(n13053), .B(n13052), .Z(n13048) );
  NANDN U806 ( .A(n13087), .B(n13086), .Z(n13082) );
  NANDN U807 ( .A(n13121), .B(n13120), .Z(n13116) );
  NANDN U808 ( .A(n13155), .B(n13154), .Z(n13150) );
  NANDN U809 ( .A(n13206), .B(n13205), .Z(n13201) );
  NANDN U810 ( .A(n13240), .B(n13239), .Z(n13235) );
  NANDN U811 ( .A(n13274), .B(n13273), .Z(n13269) );
  NANDN U812 ( .A(n13308), .B(n13307), .Z(n13303) );
  NANDN U813 ( .A(n13342), .B(n13341), .Z(n13337) );
  NANDN U814 ( .A(n13410), .B(n13409), .Z(n13405) );
  NANDN U815 ( .A(n13444), .B(n13443), .Z(n13439) );
  NANDN U816 ( .A(n13478), .B(n13477), .Z(n13473) );
  NANDN U817 ( .A(n13512), .B(n13511), .Z(n13507) );
  NANDN U818 ( .A(n13546), .B(n13545), .Z(n13541) );
  NANDN U819 ( .A(n13597), .B(n13596), .Z(n13592) );
  NANDN U820 ( .A(n13631), .B(n13630), .Z(n13626) );
  NANDN U821 ( .A(n13665), .B(n13664), .Z(n13660) );
  NANDN U822 ( .A(n13699), .B(n13698), .Z(n13694) );
  NANDN U823 ( .A(n13733), .B(n13732), .Z(n13728) );
  NANDN U824 ( .A(n13784), .B(n13783), .Z(n13779) );
  NANDN U825 ( .A(n13818), .B(n13817), .Z(n13813) );
  NANDN U826 ( .A(n13852), .B(n13851), .Z(n13847) );
  NANDN U827 ( .A(n13886), .B(n13885), .Z(n13881) );
  NANDN U828 ( .A(n13920), .B(n13919), .Z(n13915) );
  NANDN U829 ( .A(n13971), .B(n13970), .Z(n13966) );
  NANDN U830 ( .A(n14005), .B(n14004), .Z(n14000) );
  NANDN U831 ( .A(n14039), .B(n14038), .Z(n14034) );
  NANDN U832 ( .A(n14073), .B(n14072), .Z(n14068) );
  NANDN U833 ( .A(n14107), .B(n14106), .Z(n14102) );
  NANDN U834 ( .A(n14158), .B(n14157), .Z(n14153) );
  NANDN U835 ( .A(n14192), .B(n14191), .Z(n14187) );
  NANDN U836 ( .A(n14226), .B(n14225), .Z(n14221) );
  NANDN U837 ( .A(n14260), .B(n14259), .Z(n14255) );
  NANDN U838 ( .A(n14294), .B(n14293), .Z(n14289) );
  NANDN U839 ( .A(n14345), .B(n14344), .Z(n14340) );
  NANDN U840 ( .A(n14379), .B(n14378), .Z(n14374) );
  NANDN U841 ( .A(n14413), .B(n14412), .Z(n14408) );
  NANDN U842 ( .A(n14447), .B(n14446), .Z(n14442) );
  NANDN U843 ( .A(n14481), .B(n14480), .Z(n14476) );
  NANDN U844 ( .A(n14532), .B(n14531), .Z(n14527) );
  NANDN U845 ( .A(n14566), .B(n14565), .Z(n14561) );
  NANDN U846 ( .A(n14600), .B(n14599), .Z(n14595) );
  NANDN U847 ( .A(n14634), .B(n14633), .Z(n14629) );
  NANDN U848 ( .A(n14668), .B(n14667), .Z(n14663) );
  NANDN U849 ( .A(n14719), .B(n14718), .Z(n14714) );
  NANDN U850 ( .A(n14753), .B(n14752), .Z(n14748) );
  NANDN U851 ( .A(n14787), .B(n14786), .Z(n14782) );
  NANDN U852 ( .A(n14821), .B(n14820), .Z(n14816) );
  NANDN U853 ( .A(n14855), .B(n14854), .Z(n14850) );
  NANDN U854 ( .A(n14906), .B(n14905), .Z(n14901) );
  NANDN U855 ( .A(n14940), .B(n14939), .Z(n14935) );
  NANDN U856 ( .A(n14974), .B(n14973), .Z(n14969) );
  NANDN U857 ( .A(n15008), .B(n15007), .Z(n15003) );
  NANDN U858 ( .A(n15042), .B(n15041), .Z(n15037) );
  NANDN U859 ( .A(n15093), .B(n15092), .Z(n15088) );
  NANDN U860 ( .A(n15127), .B(n15126), .Z(n15122) );
  NANDN U861 ( .A(n15161), .B(n15160), .Z(n15156) );
  NANDN U862 ( .A(n15195), .B(n15194), .Z(n15190) );
  NANDN U863 ( .A(n15229), .B(n15228), .Z(n15224) );
  NANDN U864 ( .A(n15297), .B(n15296), .Z(n15292) );
  NANDN U865 ( .A(n15331), .B(n15330), .Z(n15326) );
  NANDN U866 ( .A(n15365), .B(n15364), .Z(n15360) );
  NANDN U867 ( .A(n15399), .B(n15398), .Z(n15394) );
  NANDN U868 ( .A(n15433), .B(n15432), .Z(n15428) );
  NANDN U869 ( .A(n15484), .B(n15483), .Z(n15479) );
  NANDN U870 ( .A(n15518), .B(n15517), .Z(n15513) );
  NANDN U871 ( .A(n15552), .B(n15551), .Z(n15547) );
  NANDN U872 ( .A(n15586), .B(n15585), .Z(n15581) );
  NANDN U873 ( .A(n15620), .B(n15619), .Z(n15615) );
  NANDN U874 ( .A(n15671), .B(n15670), .Z(n15666) );
  NANDN U875 ( .A(n15705), .B(n15704), .Z(n15700) );
  NANDN U876 ( .A(n15739), .B(n15738), .Z(n15734) );
  NANDN U877 ( .A(n15773), .B(n15772), .Z(n15768) );
  NANDN U878 ( .A(n15807), .B(n15806), .Z(n15802) );
  NANDN U879 ( .A(n15858), .B(n15857), .Z(n15853) );
  NANDN U880 ( .A(n15892), .B(n15891), .Z(n15887) );
  NANDN U881 ( .A(n15926), .B(n15925), .Z(n15921) );
  NANDN U882 ( .A(n15960), .B(n15959), .Z(n15955) );
  NANDN U883 ( .A(n15994), .B(n15993), .Z(n15989) );
  NANDN U884 ( .A(n16045), .B(n16044), .Z(n16040) );
  NANDN U885 ( .A(n16079), .B(n16078), .Z(n16074) );
  NANDN U886 ( .A(n16113), .B(n16112), .Z(n16108) );
  NANDN U887 ( .A(n16147), .B(n16146), .Z(n16142) );
  NANDN U888 ( .A(n16181), .B(n16180), .Z(n16176) );
  NANDN U889 ( .A(n16232), .B(n16231), .Z(n16227) );
  NANDN U890 ( .A(n16266), .B(n16265), .Z(n16261) );
  NANDN U891 ( .A(n16300), .B(n16299), .Z(n16295) );
  NANDN U892 ( .A(n16334), .B(n16333), .Z(n16329) );
  NANDN U893 ( .A(n16368), .B(n16367), .Z(n16363) );
  NANDN U894 ( .A(n16419), .B(n16418), .Z(n16414) );
  NANDN U895 ( .A(n16453), .B(n16452), .Z(n16448) );
  NANDN U896 ( .A(n16487), .B(n16486), .Z(n16482) );
  NANDN U897 ( .A(n16521), .B(n16520), .Z(n16516) );
  NANDN U898 ( .A(n16555), .B(n16554), .Z(n16550) );
  NANDN U899 ( .A(n16606), .B(n16605), .Z(n16601) );
  NANDN U900 ( .A(n16640), .B(n16639), .Z(n16635) );
  NANDN U901 ( .A(n16674), .B(n16673), .Z(n16669) );
  NANDN U902 ( .A(n16708), .B(n16707), .Z(n16703) );
  NANDN U903 ( .A(n16742), .B(n16741), .Z(n16737) );
  NANDN U904 ( .A(n16793), .B(n16792), .Z(n16788) );
  NANDN U905 ( .A(n16827), .B(n16826), .Z(n16822) );
  NANDN U906 ( .A(n16861), .B(n16860), .Z(n16856) );
  NANDN U907 ( .A(n16895), .B(n16894), .Z(n16890) );
  NANDN U908 ( .A(n16929), .B(n16928), .Z(n16924) );
  NANDN U909 ( .A(n16980), .B(n16979), .Z(n16975) );
  NANDN U910 ( .A(n17014), .B(n17013), .Z(n17009) );
  NANDN U911 ( .A(n17048), .B(n17047), .Z(n17043) );
  NANDN U912 ( .A(n17082), .B(n17081), .Z(n17077) );
  NANDN U913 ( .A(n17116), .B(n17115), .Z(n17111) );
  NANDN U914 ( .A(n17178), .B(n17177), .Z(n17173) );
  NANDN U915 ( .A(n17212), .B(n17211), .Z(n17207) );
  NANDN U916 ( .A(n17246), .B(n17245), .Z(n17241) );
  NANDN U917 ( .A(n17280), .B(n17279), .Z(n17275) );
  NANDN U918 ( .A(n17314), .B(n17313), .Z(n17309) );
  NANDN U919 ( .A(n17365), .B(n17364), .Z(n17360) );
  NANDN U920 ( .A(n17399), .B(n17398), .Z(n17394) );
  NANDN U921 ( .A(n17433), .B(n17432), .Z(n17428) );
  NANDN U922 ( .A(n17467), .B(n17466), .Z(n17462) );
  NANDN U923 ( .A(n17501), .B(n17500), .Z(n17496) );
  NANDN U924 ( .A(n17552), .B(n17551), .Z(n17547) );
  NANDN U925 ( .A(n17586), .B(n17585), .Z(n17581) );
  NANDN U926 ( .A(n17620), .B(n17619), .Z(n17615) );
  NANDN U927 ( .A(n17654), .B(n17653), .Z(n17649) );
  NANDN U928 ( .A(n17688), .B(n17687), .Z(n17683) );
  NANDN U929 ( .A(n17739), .B(n17738), .Z(n17734) );
  NANDN U930 ( .A(n17773), .B(n17772), .Z(n17768) );
  NANDN U931 ( .A(n17807), .B(n17806), .Z(n17802) );
  NANDN U932 ( .A(n17841), .B(n17840), .Z(n17836) );
  NANDN U933 ( .A(n17875), .B(n17874), .Z(n17870) );
  NANDN U934 ( .A(n17926), .B(n17925), .Z(n17921) );
  NANDN U935 ( .A(n17960), .B(n17959), .Z(n17955) );
  NANDN U936 ( .A(n17994), .B(n17993), .Z(n17989) );
  NANDN U937 ( .A(n18028), .B(n18027), .Z(n18023) );
  NANDN U938 ( .A(n18062), .B(n18061), .Z(n18057) );
  NANDN U939 ( .A(n18113), .B(n18112), .Z(n18108) );
  NANDN U940 ( .A(n18147), .B(n18146), .Z(n18142) );
  NANDN U941 ( .A(n18181), .B(n18180), .Z(n18176) );
  NANDN U942 ( .A(n18215), .B(n18214), .Z(n18210) );
  NANDN U943 ( .A(n18249), .B(n18248), .Z(n18244) );
  NANDN U944 ( .A(n18300), .B(n18299), .Z(n18295) );
  NANDN U945 ( .A(n18334), .B(n18333), .Z(n18329) );
  NANDN U946 ( .A(n18368), .B(n18367), .Z(n18363) );
  NANDN U947 ( .A(n18402), .B(n18401), .Z(n18397) );
  NANDN U948 ( .A(n18436), .B(n18435), .Z(n18431) );
  NANDN U949 ( .A(n18487), .B(n18486), .Z(n18482) );
  NANDN U950 ( .A(n18521), .B(n18520), .Z(n18516) );
  NANDN U951 ( .A(n18555), .B(n18554), .Z(n18550) );
  NANDN U952 ( .A(n18589), .B(n18588), .Z(n18584) );
  NANDN U953 ( .A(n18623), .B(n18622), .Z(n18618) );
  NANDN U954 ( .A(n18674), .B(n18673), .Z(n18669) );
  NANDN U955 ( .A(n18708), .B(n18707), .Z(n18703) );
  NANDN U956 ( .A(n18742), .B(n18741), .Z(n18737) );
  NANDN U957 ( .A(n18776), .B(n18775), .Z(n18771) );
  NANDN U958 ( .A(n18810), .B(n18809), .Z(n18805) );
  NANDN U959 ( .A(n18870), .B(n18869), .Z(n18865) );
  NANDN U960 ( .A(n18904), .B(n18903), .Z(n18899) );
  NANDN U961 ( .A(n18938), .B(n18937), .Z(n18933) );
  NANDN U962 ( .A(n18972), .B(n18971), .Z(n18967) );
  NANDN U963 ( .A(n19074), .B(n19073), .Z(n19069) );
  NANDN U964 ( .A(n2445), .B(n2444), .Z(n2440) );
  NANDN U965 ( .A(n2820), .B(n2819), .Z(n2815) );
  NANDN U966 ( .A(n3194), .B(n3193), .Z(n3189) );
  NANDN U967 ( .A(n3568), .B(n3567), .Z(n3563) );
  NANDN U968 ( .A(n3957), .B(n3956), .Z(n3952) );
  NANDN U969 ( .A(n4331), .B(n4330), .Z(n4326) );
  NANDN U970 ( .A(n4705), .B(n4704), .Z(n4700) );
  NANDN U971 ( .A(n5079), .B(n5078), .Z(n5074) );
  NANDN U972 ( .A(n5453), .B(n5452), .Z(n5448) );
  NANDN U973 ( .A(n5845), .B(n5844), .Z(n5840) );
  NANDN U974 ( .A(n6219), .B(n6218), .Z(n6214) );
  NANDN U975 ( .A(n6593), .B(n6592), .Z(n6588) );
  NANDN U976 ( .A(n6967), .B(n6966), .Z(n6962) );
  NANDN U977 ( .A(n7341), .B(n7340), .Z(n7336) );
  NANDN U978 ( .A(n7732), .B(n7731), .Z(n7727) );
  NANDN U979 ( .A(n8106), .B(n8105), .Z(n8101) );
  NANDN U980 ( .A(n8480), .B(n8479), .Z(n8475) );
  NANDN U981 ( .A(n8854), .B(n8853), .Z(n8849) );
  NANDN U982 ( .A(n9228), .B(n9227), .Z(n9223) );
  NANDN U983 ( .A(n9619), .B(n9618), .Z(n9614) );
  NANDN U984 ( .A(n9993), .B(n9992), .Z(n9988) );
  NANDN U985 ( .A(n10367), .B(n10366), .Z(n10362) );
  NANDN U986 ( .A(n10741), .B(n10740), .Z(n10736) );
  NANDN U987 ( .A(n11115), .B(n11114), .Z(n11110) );
  NANDN U988 ( .A(n11506), .B(n11505), .Z(n11501) );
  NANDN U989 ( .A(n11880), .B(n11879), .Z(n11875) );
  NANDN U990 ( .A(n12254), .B(n12253), .Z(n12249) );
  NANDN U991 ( .A(n12628), .B(n12627), .Z(n12623) );
  NANDN U992 ( .A(n13002), .B(n13001), .Z(n12997) );
  NANDN U993 ( .A(n13393), .B(n13392), .Z(n13388) );
  NANDN U994 ( .A(n13767), .B(n13766), .Z(n13762) );
  NANDN U995 ( .A(n14141), .B(n14140), .Z(n14136) );
  NANDN U996 ( .A(n14515), .B(n14514), .Z(n14510) );
  NANDN U997 ( .A(n14889), .B(n14888), .Z(n14884) );
  NANDN U998 ( .A(n15280), .B(n15279), .Z(n15275) );
  NANDN U999 ( .A(n15654), .B(n15653), .Z(n15649) );
  NANDN U1000 ( .A(n16028), .B(n16027), .Z(n16023) );
  NANDN U1001 ( .A(n16402), .B(n16401), .Z(n16397) );
  NANDN U1002 ( .A(n16776), .B(n16775), .Z(n16771) );
  NANDN U1003 ( .A(n17161), .B(n17160), .Z(n17156) );
  NANDN U1004 ( .A(n17535), .B(n17534), .Z(n17530) );
  NANDN U1005 ( .A(n17909), .B(n17908), .Z(n17904) );
  NANDN U1006 ( .A(n18283), .B(n18282), .Z(n18278) );
  NANDN U1007 ( .A(n18657), .B(n18656), .Z(n18652) );
  NANDN U1008 ( .A(n5827), .B(n5826), .Z(n5822) );
  NANDN U1009 ( .A(n7715), .B(n7714), .Z(n7710) );
  NANDN U1010 ( .A(n11489), .B(n11488), .Z(n11484) );
  NAND U1011 ( .A(n2101), .B(n2100), .Z(n2096) );
  NAND U1012 ( .A(n2092), .B(n2091), .Z(n2087) );
  NAND U1013 ( .A(n2083), .B(n2082), .Z(n2078) );
  NANDN U1014 ( .A(n19091), .B(n19090), .Z(n19086) );
  NANDN U1015 ( .A(n15263), .B(n15262), .Z(n15258) );
  NANDN U1016 ( .A(n19040), .B(n19039), .Z(n19035) );
  NAND U1017 ( .A(n19006), .B(n19003), .Z(n19002) );
  IV U1018 ( .A(n19017), .Z(n2) );
  IV U1019 ( .A(B[1023]), .Z(n3) );
  IV U1020 ( .A(n19439), .Z(n4) );
  IV U1021 ( .A(n19448), .Z(n5) );
  IV U1022 ( .A(n19453), .Z(n6) );
  IV U1023 ( .A(B[1000]), .Z(n7) );
  IV U1024 ( .A(n19452), .Z(n8) );
  IV U1025 ( .A(n2116), .Z(n9) );
  IV U1026 ( .A(B[999]), .Z(n10) );
  IV U1027 ( .A(n19260), .Z(n11) );
  IV U1028 ( .A(n19269), .Z(n12) );
  IV U1029 ( .A(n19274), .Z(n13) );
  IV U1030 ( .A(B[100]), .Z(n14) );
  IV U1031 ( .A(n19273), .Z(n15) );
  IV U1032 ( .A(n2268), .Z(n16) );
  IV U1033 ( .A(B[99]), .Z(n17) );
  IV U1034 ( .A(n18843), .Z(n18) );
  IV U1035 ( .A(n18852), .Z(n19) );
  IV U1036 ( .A(n18857), .Z(n20) );
  IV U1037 ( .A(B[10]), .Z(n21) );
  IV U1038 ( .A(n18856), .Z(n22) );
  IV U1039 ( .A(n3950), .Z(n23) );
  IV U1040 ( .A(B[9]), .Z(n24) );
  IV U1041 ( .A(n17150), .Z(n25) );
  IV U1042 ( .A(A[3]), .Z(n26) );
  XNOR U1043 ( .A(n28), .B(n29), .Z(PRODUCT[1]) );
  AND U1044 ( .A(A[0]), .B(B[0]), .Z(PRODUCT[0]) );
  AND U1045 ( .A(n30), .B(n31), .Z(\A2[9] ) );
  AND U1046 ( .A(n32), .B(n33), .Z(\A2[99] ) );
  AND U1047 ( .A(n34), .B(n35), .Z(\A2[999] ) );
  AND U1048 ( .A(n36), .B(n37), .Z(\A2[998] ) );
  AND U1049 ( .A(n38), .B(n39), .Z(\A2[997] ) );
  AND U1050 ( .A(n40), .B(n41), .Z(\A2[996] ) );
  AND U1051 ( .A(n42), .B(n43), .Z(\A2[995] ) );
  AND U1052 ( .A(n44), .B(n45), .Z(\A2[994] ) );
  AND U1053 ( .A(n46), .B(n47), .Z(\A2[993] ) );
  AND U1054 ( .A(n48), .B(n49), .Z(\A2[992] ) );
  AND U1055 ( .A(n50), .B(n51), .Z(\A2[991] ) );
  AND U1056 ( .A(n52), .B(n53), .Z(\A2[990] ) );
  AND U1057 ( .A(n54), .B(n55), .Z(\A2[98] ) );
  AND U1058 ( .A(n56), .B(n57), .Z(\A2[989] ) );
  AND U1059 ( .A(n58), .B(n59), .Z(\A2[988] ) );
  AND U1060 ( .A(n60), .B(n61), .Z(\A2[987] ) );
  AND U1061 ( .A(n62), .B(n63), .Z(\A2[986] ) );
  AND U1062 ( .A(n64), .B(n65), .Z(\A2[985] ) );
  AND U1063 ( .A(n66), .B(n67), .Z(\A2[984] ) );
  AND U1064 ( .A(n68), .B(n69), .Z(\A2[983] ) );
  AND U1065 ( .A(n70), .B(n71), .Z(\A2[982] ) );
  AND U1066 ( .A(n72), .B(n73), .Z(\A2[981] ) );
  AND U1067 ( .A(n74), .B(n75), .Z(\A2[980] ) );
  AND U1068 ( .A(n76), .B(n77), .Z(\A2[97] ) );
  AND U1069 ( .A(n78), .B(n79), .Z(\A2[979] ) );
  AND U1070 ( .A(n80), .B(n81), .Z(\A2[978] ) );
  AND U1071 ( .A(n82), .B(n83), .Z(\A2[977] ) );
  AND U1072 ( .A(n84), .B(n85), .Z(\A2[976] ) );
  AND U1073 ( .A(n86), .B(n87), .Z(\A2[975] ) );
  AND U1074 ( .A(n88), .B(n89), .Z(\A2[974] ) );
  AND U1075 ( .A(n90), .B(n91), .Z(\A2[973] ) );
  AND U1076 ( .A(n92), .B(n93), .Z(\A2[972] ) );
  AND U1077 ( .A(n94), .B(n95), .Z(\A2[971] ) );
  AND U1078 ( .A(n96), .B(n97), .Z(\A2[970] ) );
  AND U1079 ( .A(n98), .B(n99), .Z(\A2[96] ) );
  AND U1080 ( .A(n100), .B(n101), .Z(\A2[969] ) );
  AND U1081 ( .A(n102), .B(n103), .Z(\A2[968] ) );
  AND U1082 ( .A(n104), .B(n105), .Z(\A2[967] ) );
  AND U1083 ( .A(n106), .B(n107), .Z(\A2[966] ) );
  AND U1084 ( .A(n108), .B(n109), .Z(\A2[965] ) );
  AND U1085 ( .A(n110), .B(n111), .Z(\A2[964] ) );
  AND U1086 ( .A(n112), .B(n113), .Z(\A2[963] ) );
  AND U1087 ( .A(n114), .B(n115), .Z(\A2[962] ) );
  AND U1088 ( .A(n116), .B(n117), .Z(\A2[961] ) );
  AND U1089 ( .A(n118), .B(n119), .Z(\A2[960] ) );
  AND U1090 ( .A(n120), .B(n121), .Z(\A2[95] ) );
  AND U1091 ( .A(n122), .B(n123), .Z(\A2[959] ) );
  AND U1092 ( .A(n124), .B(n125), .Z(\A2[958] ) );
  AND U1093 ( .A(n126), .B(n127), .Z(\A2[957] ) );
  AND U1094 ( .A(n128), .B(n129), .Z(\A2[956] ) );
  AND U1095 ( .A(n130), .B(n131), .Z(\A2[955] ) );
  AND U1096 ( .A(n132), .B(n133), .Z(\A2[954] ) );
  AND U1097 ( .A(n134), .B(n135), .Z(\A2[953] ) );
  AND U1098 ( .A(n136), .B(n137), .Z(\A2[952] ) );
  AND U1099 ( .A(n138), .B(n139), .Z(\A2[951] ) );
  AND U1100 ( .A(n140), .B(n141), .Z(\A2[950] ) );
  AND U1101 ( .A(n142), .B(n143), .Z(\A2[94] ) );
  AND U1102 ( .A(n144), .B(n145), .Z(\A2[949] ) );
  AND U1103 ( .A(n146), .B(n147), .Z(\A2[948] ) );
  AND U1104 ( .A(n148), .B(n149), .Z(\A2[947] ) );
  AND U1105 ( .A(n150), .B(n151), .Z(\A2[946] ) );
  AND U1106 ( .A(n152), .B(n153), .Z(\A2[945] ) );
  AND U1107 ( .A(n154), .B(n155), .Z(\A2[944] ) );
  AND U1108 ( .A(n156), .B(n157), .Z(\A2[943] ) );
  AND U1109 ( .A(n158), .B(n159), .Z(\A2[942] ) );
  AND U1110 ( .A(n160), .B(n161), .Z(\A2[941] ) );
  AND U1111 ( .A(n162), .B(n163), .Z(\A2[940] ) );
  AND U1112 ( .A(n164), .B(n165), .Z(\A2[93] ) );
  AND U1113 ( .A(n166), .B(n167), .Z(\A2[939] ) );
  AND U1114 ( .A(n168), .B(n169), .Z(\A2[938] ) );
  AND U1115 ( .A(n170), .B(n171), .Z(\A2[937] ) );
  AND U1116 ( .A(n172), .B(n173), .Z(\A2[936] ) );
  AND U1117 ( .A(n174), .B(n175), .Z(\A2[935] ) );
  AND U1118 ( .A(n176), .B(n177), .Z(\A2[934] ) );
  AND U1119 ( .A(n178), .B(n179), .Z(\A2[933] ) );
  AND U1120 ( .A(n180), .B(n181), .Z(\A2[932] ) );
  AND U1121 ( .A(n182), .B(n183), .Z(\A2[931] ) );
  AND U1122 ( .A(n184), .B(n185), .Z(\A2[930] ) );
  AND U1123 ( .A(n186), .B(n187), .Z(\A2[92] ) );
  AND U1124 ( .A(n188), .B(n189), .Z(\A2[929] ) );
  AND U1125 ( .A(n190), .B(n191), .Z(\A2[928] ) );
  AND U1126 ( .A(n192), .B(n193), .Z(\A2[927] ) );
  AND U1127 ( .A(n194), .B(n195), .Z(\A2[926] ) );
  AND U1128 ( .A(n196), .B(n197), .Z(\A2[925] ) );
  AND U1129 ( .A(n198), .B(n199), .Z(\A2[924] ) );
  AND U1130 ( .A(n200), .B(n201), .Z(\A2[923] ) );
  AND U1131 ( .A(n202), .B(n203), .Z(\A2[922] ) );
  AND U1132 ( .A(n204), .B(n205), .Z(\A2[921] ) );
  AND U1133 ( .A(n206), .B(n207), .Z(\A2[920] ) );
  AND U1134 ( .A(n208), .B(n209), .Z(\A2[91] ) );
  AND U1135 ( .A(n210), .B(n211), .Z(\A2[919] ) );
  AND U1136 ( .A(n212), .B(n213), .Z(\A2[918] ) );
  AND U1137 ( .A(n214), .B(n215), .Z(\A2[917] ) );
  AND U1138 ( .A(n216), .B(n217), .Z(\A2[916] ) );
  AND U1139 ( .A(n218), .B(n219), .Z(\A2[915] ) );
  AND U1140 ( .A(n220), .B(n221), .Z(\A2[914] ) );
  AND U1141 ( .A(n222), .B(n223), .Z(\A2[913] ) );
  AND U1142 ( .A(n224), .B(n225), .Z(\A2[912] ) );
  AND U1143 ( .A(n226), .B(n227), .Z(\A2[911] ) );
  AND U1144 ( .A(n228), .B(n229), .Z(\A2[910] ) );
  AND U1145 ( .A(n230), .B(n231), .Z(\A2[90] ) );
  AND U1146 ( .A(n232), .B(n233), .Z(\A2[909] ) );
  AND U1147 ( .A(n234), .B(n235), .Z(\A2[908] ) );
  AND U1148 ( .A(n236), .B(n237), .Z(\A2[907] ) );
  AND U1149 ( .A(n238), .B(n239), .Z(\A2[906] ) );
  AND U1150 ( .A(n240), .B(n241), .Z(\A2[905] ) );
  AND U1151 ( .A(n242), .B(n243), .Z(\A2[904] ) );
  AND U1152 ( .A(n244), .B(n245), .Z(\A2[903] ) );
  AND U1153 ( .A(n246), .B(n247), .Z(\A2[902] ) );
  AND U1154 ( .A(n248), .B(n249), .Z(\A2[901] ) );
  AND U1155 ( .A(n250), .B(n251), .Z(\A2[900] ) );
  AND U1156 ( .A(n252), .B(n253), .Z(\A2[8] ) );
  AND U1157 ( .A(n254), .B(n255), .Z(\A2[89] ) );
  AND U1158 ( .A(n256), .B(n257), .Z(\A2[899] ) );
  AND U1159 ( .A(n258), .B(n259), .Z(\A2[898] ) );
  AND U1160 ( .A(n260), .B(n261), .Z(\A2[897] ) );
  AND U1161 ( .A(n262), .B(n263), .Z(\A2[896] ) );
  AND U1162 ( .A(n264), .B(n265), .Z(\A2[895] ) );
  AND U1163 ( .A(n266), .B(n267), .Z(\A2[894] ) );
  AND U1164 ( .A(n268), .B(n269), .Z(\A2[893] ) );
  AND U1165 ( .A(n270), .B(n271), .Z(\A2[892] ) );
  AND U1166 ( .A(n272), .B(n273), .Z(\A2[891] ) );
  AND U1167 ( .A(n274), .B(n275), .Z(\A2[890] ) );
  AND U1168 ( .A(n276), .B(n277), .Z(\A2[88] ) );
  AND U1169 ( .A(n278), .B(n279), .Z(\A2[889] ) );
  AND U1170 ( .A(n280), .B(n281), .Z(\A2[888] ) );
  AND U1171 ( .A(n282), .B(n283), .Z(\A2[887] ) );
  AND U1172 ( .A(n284), .B(n285), .Z(\A2[886] ) );
  AND U1173 ( .A(n286), .B(n287), .Z(\A2[885] ) );
  AND U1174 ( .A(n288), .B(n289), .Z(\A2[884] ) );
  AND U1175 ( .A(n290), .B(n291), .Z(\A2[883] ) );
  AND U1176 ( .A(n292), .B(n293), .Z(\A2[882] ) );
  AND U1177 ( .A(n294), .B(n295), .Z(\A2[881] ) );
  AND U1178 ( .A(n296), .B(n297), .Z(\A2[880] ) );
  AND U1179 ( .A(n298), .B(n299), .Z(\A2[87] ) );
  AND U1180 ( .A(n300), .B(n301), .Z(\A2[879] ) );
  AND U1181 ( .A(n302), .B(n303), .Z(\A2[878] ) );
  AND U1182 ( .A(n304), .B(n305), .Z(\A2[877] ) );
  AND U1183 ( .A(n306), .B(n307), .Z(\A2[876] ) );
  AND U1184 ( .A(n308), .B(n309), .Z(\A2[875] ) );
  AND U1185 ( .A(n310), .B(n311), .Z(\A2[874] ) );
  AND U1186 ( .A(n312), .B(n313), .Z(\A2[873] ) );
  AND U1187 ( .A(n314), .B(n315), .Z(\A2[872] ) );
  AND U1188 ( .A(n316), .B(n317), .Z(\A2[871] ) );
  AND U1189 ( .A(n318), .B(n319), .Z(\A2[870] ) );
  AND U1190 ( .A(n320), .B(n321), .Z(\A2[86] ) );
  AND U1191 ( .A(n322), .B(n323), .Z(\A2[869] ) );
  AND U1192 ( .A(n324), .B(n325), .Z(\A2[868] ) );
  AND U1193 ( .A(n326), .B(n327), .Z(\A2[867] ) );
  AND U1194 ( .A(n328), .B(n329), .Z(\A2[866] ) );
  AND U1195 ( .A(n330), .B(n331), .Z(\A2[865] ) );
  AND U1196 ( .A(n332), .B(n333), .Z(\A2[864] ) );
  AND U1197 ( .A(n334), .B(n335), .Z(\A2[863] ) );
  AND U1198 ( .A(n336), .B(n337), .Z(\A2[862] ) );
  AND U1199 ( .A(n338), .B(n339), .Z(\A2[861] ) );
  AND U1200 ( .A(n340), .B(n341), .Z(\A2[860] ) );
  AND U1201 ( .A(n342), .B(n343), .Z(\A2[85] ) );
  AND U1202 ( .A(n344), .B(n345), .Z(\A2[859] ) );
  AND U1203 ( .A(n346), .B(n347), .Z(\A2[858] ) );
  AND U1204 ( .A(n348), .B(n349), .Z(\A2[857] ) );
  AND U1205 ( .A(n350), .B(n351), .Z(\A2[856] ) );
  AND U1206 ( .A(n352), .B(n353), .Z(\A2[855] ) );
  AND U1207 ( .A(n354), .B(n355), .Z(\A2[854] ) );
  AND U1208 ( .A(n356), .B(n357), .Z(\A2[853] ) );
  AND U1209 ( .A(n358), .B(n359), .Z(\A2[852] ) );
  AND U1210 ( .A(n360), .B(n361), .Z(\A2[851] ) );
  AND U1211 ( .A(n362), .B(n363), .Z(\A2[850] ) );
  AND U1212 ( .A(n364), .B(n365), .Z(\A2[84] ) );
  AND U1213 ( .A(n366), .B(n367), .Z(\A2[849] ) );
  AND U1214 ( .A(n368), .B(n369), .Z(\A2[848] ) );
  AND U1215 ( .A(n370), .B(n371), .Z(\A2[847] ) );
  AND U1216 ( .A(n372), .B(n373), .Z(\A2[846] ) );
  AND U1217 ( .A(n374), .B(n375), .Z(\A2[845] ) );
  AND U1218 ( .A(n376), .B(n377), .Z(\A2[844] ) );
  AND U1219 ( .A(n378), .B(n379), .Z(\A2[843] ) );
  AND U1220 ( .A(n380), .B(n381), .Z(\A2[842] ) );
  AND U1221 ( .A(n382), .B(n383), .Z(\A2[841] ) );
  AND U1222 ( .A(n384), .B(n385), .Z(\A2[840] ) );
  AND U1223 ( .A(n386), .B(n387), .Z(\A2[83] ) );
  AND U1224 ( .A(n388), .B(n389), .Z(\A2[839] ) );
  AND U1225 ( .A(n390), .B(n391), .Z(\A2[838] ) );
  AND U1226 ( .A(n392), .B(n393), .Z(\A2[837] ) );
  AND U1227 ( .A(n394), .B(n395), .Z(\A2[836] ) );
  AND U1228 ( .A(n396), .B(n397), .Z(\A2[835] ) );
  AND U1229 ( .A(n398), .B(n399), .Z(\A2[834] ) );
  AND U1230 ( .A(n400), .B(n401), .Z(\A2[833] ) );
  AND U1231 ( .A(n402), .B(n403), .Z(\A2[832] ) );
  AND U1232 ( .A(n404), .B(n405), .Z(\A2[831] ) );
  AND U1233 ( .A(n406), .B(n407), .Z(\A2[830] ) );
  AND U1234 ( .A(n408), .B(n409), .Z(\A2[82] ) );
  AND U1235 ( .A(n410), .B(n411), .Z(\A2[829] ) );
  AND U1236 ( .A(n412), .B(n413), .Z(\A2[828] ) );
  AND U1237 ( .A(n414), .B(n415), .Z(\A2[827] ) );
  AND U1238 ( .A(n416), .B(n417), .Z(\A2[826] ) );
  AND U1239 ( .A(n418), .B(n419), .Z(\A2[825] ) );
  AND U1240 ( .A(n420), .B(n421), .Z(\A2[824] ) );
  AND U1241 ( .A(n422), .B(n423), .Z(\A2[823] ) );
  AND U1242 ( .A(n424), .B(n425), .Z(\A2[822] ) );
  AND U1243 ( .A(n426), .B(n427), .Z(\A2[821] ) );
  AND U1244 ( .A(n428), .B(n429), .Z(\A2[820] ) );
  AND U1245 ( .A(n430), .B(n431), .Z(\A2[81] ) );
  AND U1246 ( .A(n432), .B(n433), .Z(\A2[819] ) );
  AND U1247 ( .A(n434), .B(n435), .Z(\A2[818] ) );
  AND U1248 ( .A(n436), .B(n437), .Z(\A2[817] ) );
  AND U1249 ( .A(n438), .B(n439), .Z(\A2[816] ) );
  AND U1250 ( .A(n440), .B(n441), .Z(\A2[815] ) );
  AND U1251 ( .A(n442), .B(n443), .Z(\A2[814] ) );
  AND U1252 ( .A(n444), .B(n445), .Z(\A2[813] ) );
  AND U1253 ( .A(n446), .B(n447), .Z(\A2[812] ) );
  AND U1254 ( .A(n448), .B(n449), .Z(\A2[811] ) );
  AND U1255 ( .A(n450), .B(n451), .Z(\A2[810] ) );
  AND U1256 ( .A(n452), .B(n453), .Z(\A2[80] ) );
  AND U1257 ( .A(n454), .B(n455), .Z(\A2[809] ) );
  AND U1258 ( .A(n456), .B(n457), .Z(\A2[808] ) );
  AND U1259 ( .A(n458), .B(n459), .Z(\A2[807] ) );
  AND U1260 ( .A(n460), .B(n461), .Z(\A2[806] ) );
  AND U1261 ( .A(n462), .B(n463), .Z(\A2[805] ) );
  AND U1262 ( .A(n464), .B(n465), .Z(\A2[804] ) );
  AND U1263 ( .A(n466), .B(n467), .Z(\A2[803] ) );
  AND U1264 ( .A(n468), .B(n469), .Z(\A2[802] ) );
  AND U1265 ( .A(n470), .B(n471), .Z(\A2[801] ) );
  AND U1266 ( .A(n472), .B(n473), .Z(\A2[800] ) );
  AND U1267 ( .A(n474), .B(n475), .Z(\A2[7] ) );
  AND U1268 ( .A(n476), .B(n477), .Z(\A2[79] ) );
  AND U1269 ( .A(n478), .B(n479), .Z(\A2[799] ) );
  AND U1270 ( .A(n480), .B(n481), .Z(\A2[798] ) );
  AND U1271 ( .A(n482), .B(n483), .Z(\A2[797] ) );
  AND U1272 ( .A(n484), .B(n485), .Z(\A2[796] ) );
  AND U1273 ( .A(n486), .B(n487), .Z(\A2[795] ) );
  AND U1274 ( .A(n488), .B(n489), .Z(\A2[794] ) );
  AND U1275 ( .A(n490), .B(n491), .Z(\A2[793] ) );
  AND U1276 ( .A(n492), .B(n493), .Z(\A2[792] ) );
  AND U1277 ( .A(n494), .B(n495), .Z(\A2[791] ) );
  AND U1278 ( .A(n496), .B(n497), .Z(\A2[790] ) );
  AND U1279 ( .A(n498), .B(n499), .Z(\A2[78] ) );
  AND U1280 ( .A(n500), .B(n501), .Z(\A2[789] ) );
  AND U1281 ( .A(n502), .B(n503), .Z(\A2[788] ) );
  AND U1282 ( .A(n504), .B(n505), .Z(\A2[787] ) );
  AND U1283 ( .A(n506), .B(n507), .Z(\A2[786] ) );
  AND U1284 ( .A(n508), .B(n509), .Z(\A2[785] ) );
  AND U1285 ( .A(n510), .B(n511), .Z(\A2[784] ) );
  AND U1286 ( .A(n512), .B(n513), .Z(\A2[783] ) );
  AND U1287 ( .A(n514), .B(n515), .Z(\A2[782] ) );
  AND U1288 ( .A(n516), .B(n517), .Z(\A2[781] ) );
  AND U1289 ( .A(n518), .B(n519), .Z(\A2[780] ) );
  AND U1290 ( .A(n520), .B(n521), .Z(\A2[77] ) );
  AND U1291 ( .A(n522), .B(n523), .Z(\A2[779] ) );
  AND U1292 ( .A(n524), .B(n525), .Z(\A2[778] ) );
  AND U1293 ( .A(n526), .B(n527), .Z(\A2[777] ) );
  AND U1294 ( .A(n528), .B(n529), .Z(\A2[776] ) );
  AND U1295 ( .A(n530), .B(n531), .Z(\A2[775] ) );
  AND U1296 ( .A(n532), .B(n533), .Z(\A2[774] ) );
  AND U1297 ( .A(n534), .B(n535), .Z(\A2[773] ) );
  AND U1298 ( .A(n536), .B(n537), .Z(\A2[772] ) );
  AND U1299 ( .A(n538), .B(n539), .Z(\A2[771] ) );
  AND U1300 ( .A(n540), .B(n541), .Z(\A2[770] ) );
  AND U1301 ( .A(n542), .B(n543), .Z(\A2[76] ) );
  AND U1302 ( .A(n544), .B(n545), .Z(\A2[769] ) );
  AND U1303 ( .A(n546), .B(n547), .Z(\A2[768] ) );
  AND U1304 ( .A(n548), .B(n549), .Z(\A2[767] ) );
  AND U1305 ( .A(n550), .B(n551), .Z(\A2[766] ) );
  AND U1306 ( .A(n552), .B(n553), .Z(\A2[765] ) );
  AND U1307 ( .A(n554), .B(n555), .Z(\A2[764] ) );
  AND U1308 ( .A(n556), .B(n557), .Z(\A2[763] ) );
  AND U1309 ( .A(n558), .B(n559), .Z(\A2[762] ) );
  AND U1310 ( .A(n560), .B(n561), .Z(\A2[761] ) );
  AND U1311 ( .A(n562), .B(n563), .Z(\A2[760] ) );
  AND U1312 ( .A(n564), .B(n565), .Z(\A2[75] ) );
  AND U1313 ( .A(n566), .B(n567), .Z(\A2[759] ) );
  AND U1314 ( .A(n568), .B(n569), .Z(\A2[758] ) );
  AND U1315 ( .A(n570), .B(n571), .Z(\A2[757] ) );
  AND U1316 ( .A(n572), .B(n573), .Z(\A2[756] ) );
  AND U1317 ( .A(n574), .B(n575), .Z(\A2[755] ) );
  AND U1318 ( .A(n576), .B(n577), .Z(\A2[754] ) );
  AND U1319 ( .A(n578), .B(n579), .Z(\A2[753] ) );
  AND U1320 ( .A(n580), .B(n581), .Z(\A2[752] ) );
  AND U1321 ( .A(n582), .B(n583), .Z(\A2[751] ) );
  AND U1322 ( .A(n584), .B(n585), .Z(\A2[750] ) );
  AND U1323 ( .A(n586), .B(n587), .Z(\A2[74] ) );
  AND U1324 ( .A(n588), .B(n589), .Z(\A2[749] ) );
  AND U1325 ( .A(n590), .B(n591), .Z(\A2[748] ) );
  AND U1326 ( .A(n592), .B(n593), .Z(\A2[747] ) );
  AND U1327 ( .A(n594), .B(n595), .Z(\A2[746] ) );
  AND U1328 ( .A(n596), .B(n597), .Z(\A2[745] ) );
  AND U1329 ( .A(n598), .B(n599), .Z(\A2[744] ) );
  AND U1330 ( .A(n600), .B(n601), .Z(\A2[743] ) );
  AND U1331 ( .A(n602), .B(n603), .Z(\A2[742] ) );
  AND U1332 ( .A(n604), .B(n605), .Z(\A2[741] ) );
  AND U1333 ( .A(n606), .B(n607), .Z(\A2[740] ) );
  AND U1334 ( .A(n608), .B(n609), .Z(\A2[73] ) );
  AND U1335 ( .A(n610), .B(n611), .Z(\A2[739] ) );
  AND U1336 ( .A(n612), .B(n613), .Z(\A2[738] ) );
  AND U1337 ( .A(n614), .B(n615), .Z(\A2[737] ) );
  AND U1338 ( .A(n616), .B(n617), .Z(\A2[736] ) );
  AND U1339 ( .A(n618), .B(n619), .Z(\A2[735] ) );
  AND U1340 ( .A(n620), .B(n621), .Z(\A2[734] ) );
  AND U1341 ( .A(n622), .B(n623), .Z(\A2[733] ) );
  AND U1342 ( .A(n624), .B(n625), .Z(\A2[732] ) );
  AND U1343 ( .A(n626), .B(n627), .Z(\A2[731] ) );
  AND U1344 ( .A(n628), .B(n629), .Z(\A2[730] ) );
  AND U1345 ( .A(n630), .B(n631), .Z(\A2[72] ) );
  AND U1346 ( .A(n632), .B(n633), .Z(\A2[729] ) );
  AND U1347 ( .A(n634), .B(n635), .Z(\A2[728] ) );
  AND U1348 ( .A(n636), .B(n637), .Z(\A2[727] ) );
  AND U1349 ( .A(n638), .B(n639), .Z(\A2[726] ) );
  AND U1350 ( .A(n640), .B(n641), .Z(\A2[725] ) );
  AND U1351 ( .A(n642), .B(n643), .Z(\A2[724] ) );
  AND U1352 ( .A(n644), .B(n645), .Z(\A2[723] ) );
  AND U1353 ( .A(n646), .B(n647), .Z(\A2[722] ) );
  AND U1354 ( .A(n648), .B(n649), .Z(\A2[721] ) );
  AND U1355 ( .A(n650), .B(n651), .Z(\A2[720] ) );
  AND U1356 ( .A(n652), .B(n653), .Z(\A2[71] ) );
  AND U1357 ( .A(n654), .B(n655), .Z(\A2[719] ) );
  AND U1358 ( .A(n656), .B(n657), .Z(\A2[718] ) );
  AND U1359 ( .A(n658), .B(n659), .Z(\A2[717] ) );
  AND U1360 ( .A(n660), .B(n661), .Z(\A2[716] ) );
  AND U1361 ( .A(n662), .B(n663), .Z(\A2[715] ) );
  AND U1362 ( .A(n664), .B(n665), .Z(\A2[714] ) );
  AND U1363 ( .A(n666), .B(n667), .Z(\A2[713] ) );
  AND U1364 ( .A(n668), .B(n669), .Z(\A2[712] ) );
  AND U1365 ( .A(n670), .B(n671), .Z(\A2[711] ) );
  AND U1366 ( .A(n672), .B(n673), .Z(\A2[710] ) );
  AND U1367 ( .A(n674), .B(n675), .Z(\A2[70] ) );
  AND U1368 ( .A(n676), .B(n677), .Z(\A2[709] ) );
  AND U1369 ( .A(n678), .B(n679), .Z(\A2[708] ) );
  AND U1370 ( .A(n680), .B(n681), .Z(\A2[707] ) );
  AND U1371 ( .A(n682), .B(n683), .Z(\A2[706] ) );
  AND U1372 ( .A(n684), .B(n685), .Z(\A2[705] ) );
  AND U1373 ( .A(n686), .B(n687), .Z(\A2[704] ) );
  AND U1374 ( .A(n688), .B(n689), .Z(\A2[703] ) );
  AND U1375 ( .A(n690), .B(n691), .Z(\A2[702] ) );
  AND U1376 ( .A(n692), .B(n693), .Z(\A2[701] ) );
  AND U1377 ( .A(n694), .B(n695), .Z(\A2[700] ) );
  AND U1378 ( .A(n696), .B(n697), .Z(\A2[6] ) );
  AND U1379 ( .A(n698), .B(n699), .Z(\A2[69] ) );
  AND U1380 ( .A(n700), .B(n701), .Z(\A2[699] ) );
  AND U1381 ( .A(n702), .B(n703), .Z(\A2[698] ) );
  AND U1382 ( .A(n704), .B(n705), .Z(\A2[697] ) );
  AND U1383 ( .A(n706), .B(n707), .Z(\A2[696] ) );
  AND U1384 ( .A(n708), .B(n709), .Z(\A2[695] ) );
  AND U1385 ( .A(n710), .B(n711), .Z(\A2[694] ) );
  AND U1386 ( .A(n712), .B(n713), .Z(\A2[693] ) );
  AND U1387 ( .A(n714), .B(n715), .Z(\A2[692] ) );
  AND U1388 ( .A(n716), .B(n717), .Z(\A2[691] ) );
  AND U1389 ( .A(n718), .B(n719), .Z(\A2[690] ) );
  AND U1390 ( .A(n720), .B(n721), .Z(\A2[68] ) );
  AND U1391 ( .A(n722), .B(n723), .Z(\A2[689] ) );
  AND U1392 ( .A(n724), .B(n725), .Z(\A2[688] ) );
  AND U1393 ( .A(n726), .B(n727), .Z(\A2[687] ) );
  AND U1394 ( .A(n728), .B(n729), .Z(\A2[686] ) );
  AND U1395 ( .A(n730), .B(n731), .Z(\A2[685] ) );
  AND U1396 ( .A(n732), .B(n733), .Z(\A2[684] ) );
  AND U1397 ( .A(n734), .B(n735), .Z(\A2[683] ) );
  AND U1398 ( .A(n736), .B(n737), .Z(\A2[682] ) );
  AND U1399 ( .A(n738), .B(n739), .Z(\A2[681] ) );
  AND U1400 ( .A(n740), .B(n741), .Z(\A2[680] ) );
  AND U1401 ( .A(n742), .B(n743), .Z(\A2[67] ) );
  AND U1402 ( .A(n744), .B(n745), .Z(\A2[679] ) );
  AND U1403 ( .A(n746), .B(n747), .Z(\A2[678] ) );
  AND U1404 ( .A(n748), .B(n749), .Z(\A2[677] ) );
  AND U1405 ( .A(n750), .B(n751), .Z(\A2[676] ) );
  AND U1406 ( .A(n752), .B(n753), .Z(\A2[675] ) );
  AND U1407 ( .A(n754), .B(n755), .Z(\A2[674] ) );
  AND U1408 ( .A(n756), .B(n757), .Z(\A2[673] ) );
  AND U1409 ( .A(n758), .B(n759), .Z(\A2[672] ) );
  AND U1410 ( .A(n760), .B(n761), .Z(\A2[671] ) );
  AND U1411 ( .A(n762), .B(n763), .Z(\A2[670] ) );
  AND U1412 ( .A(n764), .B(n765), .Z(\A2[66] ) );
  AND U1413 ( .A(n766), .B(n767), .Z(\A2[669] ) );
  AND U1414 ( .A(n768), .B(n769), .Z(\A2[668] ) );
  AND U1415 ( .A(n770), .B(n771), .Z(\A2[667] ) );
  AND U1416 ( .A(n772), .B(n773), .Z(\A2[666] ) );
  AND U1417 ( .A(n774), .B(n775), .Z(\A2[665] ) );
  AND U1418 ( .A(n776), .B(n777), .Z(\A2[664] ) );
  AND U1419 ( .A(n778), .B(n779), .Z(\A2[663] ) );
  AND U1420 ( .A(n780), .B(n781), .Z(\A2[662] ) );
  AND U1421 ( .A(n782), .B(n783), .Z(\A2[661] ) );
  AND U1422 ( .A(n784), .B(n785), .Z(\A2[660] ) );
  AND U1423 ( .A(n786), .B(n787), .Z(\A2[65] ) );
  AND U1424 ( .A(n788), .B(n789), .Z(\A2[659] ) );
  AND U1425 ( .A(n790), .B(n791), .Z(\A2[658] ) );
  AND U1426 ( .A(n792), .B(n793), .Z(\A2[657] ) );
  AND U1427 ( .A(n794), .B(n795), .Z(\A2[656] ) );
  AND U1428 ( .A(n796), .B(n797), .Z(\A2[655] ) );
  AND U1429 ( .A(n798), .B(n799), .Z(\A2[654] ) );
  AND U1430 ( .A(n800), .B(n801), .Z(\A2[653] ) );
  AND U1431 ( .A(n802), .B(n803), .Z(\A2[652] ) );
  AND U1432 ( .A(n804), .B(n805), .Z(\A2[651] ) );
  AND U1433 ( .A(n806), .B(n807), .Z(\A2[650] ) );
  AND U1434 ( .A(n808), .B(n809), .Z(\A2[64] ) );
  AND U1435 ( .A(n810), .B(n811), .Z(\A2[649] ) );
  AND U1436 ( .A(n812), .B(n813), .Z(\A2[648] ) );
  AND U1437 ( .A(n814), .B(n815), .Z(\A2[647] ) );
  AND U1438 ( .A(n816), .B(n817), .Z(\A2[646] ) );
  AND U1439 ( .A(n818), .B(n819), .Z(\A2[645] ) );
  AND U1440 ( .A(n820), .B(n821), .Z(\A2[644] ) );
  AND U1441 ( .A(n822), .B(n823), .Z(\A2[643] ) );
  AND U1442 ( .A(n824), .B(n825), .Z(\A2[642] ) );
  AND U1443 ( .A(n826), .B(n827), .Z(\A2[641] ) );
  AND U1444 ( .A(n828), .B(n829), .Z(\A2[640] ) );
  AND U1445 ( .A(n830), .B(n831), .Z(\A2[63] ) );
  AND U1446 ( .A(n832), .B(n833), .Z(\A2[639] ) );
  AND U1447 ( .A(n834), .B(n835), .Z(\A2[638] ) );
  AND U1448 ( .A(n836), .B(n837), .Z(\A2[637] ) );
  AND U1449 ( .A(n838), .B(n839), .Z(\A2[636] ) );
  AND U1450 ( .A(n840), .B(n841), .Z(\A2[635] ) );
  AND U1451 ( .A(n842), .B(n843), .Z(\A2[634] ) );
  AND U1452 ( .A(n844), .B(n845), .Z(\A2[633] ) );
  AND U1453 ( .A(n846), .B(n847), .Z(\A2[632] ) );
  AND U1454 ( .A(n848), .B(n849), .Z(\A2[631] ) );
  AND U1455 ( .A(n850), .B(n851), .Z(\A2[630] ) );
  AND U1456 ( .A(n852), .B(n853), .Z(\A2[62] ) );
  AND U1457 ( .A(n854), .B(n855), .Z(\A2[629] ) );
  AND U1458 ( .A(n856), .B(n857), .Z(\A2[628] ) );
  AND U1459 ( .A(n858), .B(n859), .Z(\A2[627] ) );
  AND U1460 ( .A(n860), .B(n861), .Z(\A2[626] ) );
  AND U1461 ( .A(n862), .B(n863), .Z(\A2[625] ) );
  AND U1462 ( .A(n864), .B(n865), .Z(\A2[624] ) );
  AND U1463 ( .A(n866), .B(n867), .Z(\A2[623] ) );
  AND U1464 ( .A(n868), .B(n869), .Z(\A2[622] ) );
  AND U1465 ( .A(n870), .B(n871), .Z(\A2[621] ) );
  AND U1466 ( .A(n872), .B(n873), .Z(\A2[620] ) );
  AND U1467 ( .A(n874), .B(n875), .Z(\A2[61] ) );
  AND U1468 ( .A(n876), .B(n877), .Z(\A2[619] ) );
  AND U1469 ( .A(n878), .B(n879), .Z(\A2[618] ) );
  AND U1470 ( .A(n880), .B(n881), .Z(\A2[617] ) );
  AND U1471 ( .A(n882), .B(n883), .Z(\A2[616] ) );
  AND U1472 ( .A(n884), .B(n885), .Z(\A2[615] ) );
  AND U1473 ( .A(n886), .B(n887), .Z(\A2[614] ) );
  AND U1474 ( .A(n888), .B(n889), .Z(\A2[613] ) );
  AND U1475 ( .A(n890), .B(n891), .Z(\A2[612] ) );
  AND U1476 ( .A(n892), .B(n893), .Z(\A2[611] ) );
  AND U1477 ( .A(n894), .B(n895), .Z(\A2[610] ) );
  AND U1478 ( .A(n896), .B(n897), .Z(\A2[60] ) );
  AND U1479 ( .A(n898), .B(n899), .Z(\A2[609] ) );
  AND U1480 ( .A(n900), .B(n901), .Z(\A2[608] ) );
  AND U1481 ( .A(n902), .B(n903), .Z(\A2[607] ) );
  AND U1482 ( .A(n904), .B(n905), .Z(\A2[606] ) );
  AND U1483 ( .A(n906), .B(n907), .Z(\A2[605] ) );
  AND U1484 ( .A(n908), .B(n909), .Z(\A2[604] ) );
  AND U1485 ( .A(n910), .B(n911), .Z(\A2[603] ) );
  AND U1486 ( .A(n912), .B(n913), .Z(\A2[602] ) );
  AND U1487 ( .A(n914), .B(n915), .Z(\A2[601] ) );
  AND U1488 ( .A(n916), .B(n917), .Z(\A2[600] ) );
  AND U1489 ( .A(n918), .B(n919), .Z(\A2[5] ) );
  AND U1490 ( .A(n920), .B(n921), .Z(\A2[59] ) );
  AND U1491 ( .A(n922), .B(n923), .Z(\A2[599] ) );
  AND U1492 ( .A(n924), .B(n925), .Z(\A2[598] ) );
  AND U1493 ( .A(n926), .B(n927), .Z(\A2[597] ) );
  AND U1494 ( .A(n928), .B(n929), .Z(\A2[596] ) );
  AND U1495 ( .A(n930), .B(n931), .Z(\A2[595] ) );
  AND U1496 ( .A(n932), .B(n933), .Z(\A2[594] ) );
  AND U1497 ( .A(n934), .B(n935), .Z(\A2[593] ) );
  AND U1498 ( .A(n936), .B(n937), .Z(\A2[592] ) );
  AND U1499 ( .A(n938), .B(n939), .Z(\A2[591] ) );
  AND U1500 ( .A(n940), .B(n941), .Z(\A2[590] ) );
  AND U1501 ( .A(n942), .B(n943), .Z(\A2[58] ) );
  AND U1502 ( .A(n944), .B(n945), .Z(\A2[589] ) );
  AND U1503 ( .A(n946), .B(n947), .Z(\A2[588] ) );
  AND U1504 ( .A(n948), .B(n949), .Z(\A2[587] ) );
  AND U1505 ( .A(n950), .B(n951), .Z(\A2[586] ) );
  AND U1506 ( .A(n952), .B(n953), .Z(\A2[585] ) );
  AND U1507 ( .A(n954), .B(n955), .Z(\A2[584] ) );
  AND U1508 ( .A(n956), .B(n957), .Z(\A2[583] ) );
  AND U1509 ( .A(n958), .B(n959), .Z(\A2[582] ) );
  AND U1510 ( .A(n960), .B(n961), .Z(\A2[581] ) );
  AND U1511 ( .A(n962), .B(n963), .Z(\A2[580] ) );
  AND U1512 ( .A(n964), .B(n965), .Z(\A2[57] ) );
  AND U1513 ( .A(n966), .B(n967), .Z(\A2[579] ) );
  AND U1514 ( .A(n968), .B(n969), .Z(\A2[578] ) );
  AND U1515 ( .A(n970), .B(n971), .Z(\A2[577] ) );
  AND U1516 ( .A(n972), .B(n973), .Z(\A2[576] ) );
  AND U1517 ( .A(n974), .B(n975), .Z(\A2[575] ) );
  AND U1518 ( .A(n976), .B(n977), .Z(\A2[574] ) );
  AND U1519 ( .A(n978), .B(n979), .Z(\A2[573] ) );
  AND U1520 ( .A(n980), .B(n981), .Z(\A2[572] ) );
  AND U1521 ( .A(n982), .B(n983), .Z(\A2[571] ) );
  AND U1522 ( .A(n984), .B(n985), .Z(\A2[570] ) );
  AND U1523 ( .A(n986), .B(n987), .Z(\A2[56] ) );
  AND U1524 ( .A(n988), .B(n989), .Z(\A2[569] ) );
  AND U1525 ( .A(n990), .B(n991), .Z(\A2[568] ) );
  AND U1526 ( .A(n992), .B(n993), .Z(\A2[567] ) );
  AND U1527 ( .A(n994), .B(n995), .Z(\A2[566] ) );
  AND U1528 ( .A(n996), .B(n997), .Z(\A2[565] ) );
  AND U1529 ( .A(n998), .B(n999), .Z(\A2[564] ) );
  AND U1530 ( .A(n1000), .B(n1001), .Z(\A2[563] ) );
  AND U1531 ( .A(n1002), .B(n1003), .Z(\A2[562] ) );
  AND U1532 ( .A(n1004), .B(n1005), .Z(\A2[561] ) );
  AND U1533 ( .A(n1006), .B(n1007), .Z(\A2[560] ) );
  AND U1534 ( .A(n1008), .B(n1009), .Z(\A2[55] ) );
  AND U1535 ( .A(n1010), .B(n1011), .Z(\A2[559] ) );
  AND U1536 ( .A(n1012), .B(n1013), .Z(\A2[558] ) );
  AND U1537 ( .A(n1014), .B(n1015), .Z(\A2[557] ) );
  AND U1538 ( .A(n1016), .B(n1017), .Z(\A2[556] ) );
  AND U1539 ( .A(n1018), .B(n1019), .Z(\A2[555] ) );
  AND U1540 ( .A(n1020), .B(n1021), .Z(\A2[554] ) );
  AND U1541 ( .A(n1022), .B(n1023), .Z(\A2[553] ) );
  AND U1542 ( .A(n1024), .B(n1025), .Z(\A2[552] ) );
  AND U1543 ( .A(n1026), .B(n1027), .Z(\A2[551] ) );
  AND U1544 ( .A(n1028), .B(n1029), .Z(\A2[550] ) );
  AND U1545 ( .A(n1030), .B(n1031), .Z(\A2[54] ) );
  AND U1546 ( .A(n1032), .B(n1033), .Z(\A2[549] ) );
  AND U1547 ( .A(n1034), .B(n1035), .Z(\A2[548] ) );
  AND U1548 ( .A(n1036), .B(n1037), .Z(\A2[547] ) );
  AND U1549 ( .A(n1038), .B(n1039), .Z(\A2[546] ) );
  AND U1550 ( .A(n1040), .B(n1041), .Z(\A2[545] ) );
  AND U1551 ( .A(n1042), .B(n1043), .Z(\A2[544] ) );
  AND U1552 ( .A(n1044), .B(n1045), .Z(\A2[543] ) );
  AND U1553 ( .A(n1046), .B(n1047), .Z(\A2[542] ) );
  AND U1554 ( .A(n1048), .B(n1049), .Z(\A2[541] ) );
  AND U1555 ( .A(n1050), .B(n1051), .Z(\A2[540] ) );
  AND U1556 ( .A(n1052), .B(n1053), .Z(\A2[53] ) );
  AND U1557 ( .A(n1054), .B(n1055), .Z(\A2[539] ) );
  AND U1558 ( .A(n1056), .B(n1057), .Z(\A2[538] ) );
  AND U1559 ( .A(n1058), .B(n1059), .Z(\A2[537] ) );
  AND U1560 ( .A(n1060), .B(n1061), .Z(\A2[536] ) );
  AND U1561 ( .A(n1062), .B(n1063), .Z(\A2[535] ) );
  AND U1562 ( .A(n1064), .B(n1065), .Z(\A2[534] ) );
  AND U1563 ( .A(n1066), .B(n1067), .Z(\A2[533] ) );
  AND U1564 ( .A(n1068), .B(n1069), .Z(\A2[532] ) );
  AND U1565 ( .A(n1070), .B(n1071), .Z(\A2[531] ) );
  AND U1566 ( .A(n1072), .B(n1073), .Z(\A2[530] ) );
  AND U1567 ( .A(n1074), .B(n1075), .Z(\A2[52] ) );
  AND U1568 ( .A(n1076), .B(n1077), .Z(\A2[529] ) );
  AND U1569 ( .A(n1078), .B(n1079), .Z(\A2[528] ) );
  AND U1570 ( .A(n1080), .B(n1081), .Z(\A2[527] ) );
  AND U1571 ( .A(n1082), .B(n1083), .Z(\A2[526] ) );
  AND U1572 ( .A(n1084), .B(n1085), .Z(\A2[525] ) );
  AND U1573 ( .A(n1086), .B(n1087), .Z(\A2[524] ) );
  AND U1574 ( .A(n1088), .B(n1089), .Z(\A2[523] ) );
  AND U1575 ( .A(n1090), .B(n1091), .Z(\A2[522] ) );
  AND U1576 ( .A(n1092), .B(n1093), .Z(\A2[521] ) );
  AND U1577 ( .A(n1094), .B(n1095), .Z(\A2[520] ) );
  AND U1578 ( .A(n1096), .B(n1097), .Z(\A2[51] ) );
  AND U1579 ( .A(n1098), .B(n1099), .Z(\A2[519] ) );
  AND U1580 ( .A(n1100), .B(n1101), .Z(\A2[518] ) );
  AND U1581 ( .A(n1102), .B(n1103), .Z(\A2[517] ) );
  AND U1582 ( .A(n1104), .B(n1105), .Z(\A2[516] ) );
  AND U1583 ( .A(n1106), .B(n1107), .Z(\A2[515] ) );
  AND U1584 ( .A(n1108), .B(n1109), .Z(\A2[514] ) );
  AND U1585 ( .A(n1110), .B(n1111), .Z(\A2[513] ) );
  AND U1586 ( .A(n1112), .B(n1113), .Z(\A2[512] ) );
  AND U1587 ( .A(n1114), .B(n1115), .Z(\A2[511] ) );
  AND U1588 ( .A(n1116), .B(n1117), .Z(\A2[510] ) );
  AND U1589 ( .A(n1118), .B(n1119), .Z(\A2[50] ) );
  AND U1590 ( .A(n1120), .B(n1121), .Z(\A2[509] ) );
  AND U1591 ( .A(n1122), .B(n1123), .Z(\A2[508] ) );
  AND U1592 ( .A(n1124), .B(n1125), .Z(\A2[507] ) );
  AND U1593 ( .A(n1126), .B(n1127), .Z(\A2[506] ) );
  AND U1594 ( .A(n1128), .B(n1129), .Z(\A2[505] ) );
  AND U1595 ( .A(n1130), .B(n1131), .Z(\A2[504] ) );
  AND U1596 ( .A(n1132), .B(n1133), .Z(\A2[503] ) );
  AND U1597 ( .A(n1134), .B(n1135), .Z(\A2[502] ) );
  AND U1598 ( .A(n1136), .B(n1137), .Z(\A2[501] ) );
  AND U1599 ( .A(n1138), .B(n1139), .Z(\A2[500] ) );
  AND U1600 ( .A(n1140), .B(n1141), .Z(\A2[4] ) );
  AND U1601 ( .A(n1142), .B(n1143), .Z(\A2[49] ) );
  AND U1602 ( .A(n1144), .B(n1145), .Z(\A2[499] ) );
  AND U1603 ( .A(n1146), .B(n1147), .Z(\A2[498] ) );
  AND U1604 ( .A(n1148), .B(n1149), .Z(\A2[497] ) );
  AND U1605 ( .A(n1150), .B(n1151), .Z(\A2[496] ) );
  AND U1606 ( .A(n1152), .B(n1153), .Z(\A2[495] ) );
  AND U1607 ( .A(n1154), .B(n1155), .Z(\A2[494] ) );
  AND U1608 ( .A(n1156), .B(n1157), .Z(\A2[493] ) );
  AND U1609 ( .A(n1158), .B(n1159), .Z(\A2[492] ) );
  AND U1610 ( .A(n1160), .B(n1161), .Z(\A2[491] ) );
  AND U1611 ( .A(n1162), .B(n1163), .Z(\A2[490] ) );
  AND U1612 ( .A(n1164), .B(n1165), .Z(\A2[48] ) );
  AND U1613 ( .A(n1166), .B(n1167), .Z(\A2[489] ) );
  AND U1614 ( .A(n1168), .B(n1169), .Z(\A2[488] ) );
  AND U1615 ( .A(n1170), .B(n1171), .Z(\A2[487] ) );
  AND U1616 ( .A(n1172), .B(n1173), .Z(\A2[486] ) );
  AND U1617 ( .A(n1174), .B(n1175), .Z(\A2[485] ) );
  AND U1618 ( .A(n1176), .B(n1177), .Z(\A2[484] ) );
  AND U1619 ( .A(n1178), .B(n1179), .Z(\A2[483] ) );
  AND U1620 ( .A(n1180), .B(n1181), .Z(\A2[482] ) );
  AND U1621 ( .A(n1182), .B(n1183), .Z(\A2[481] ) );
  AND U1622 ( .A(n1184), .B(n1185), .Z(\A2[480] ) );
  AND U1623 ( .A(n1186), .B(n1187), .Z(\A2[47] ) );
  AND U1624 ( .A(n1188), .B(n1189), .Z(\A2[479] ) );
  AND U1625 ( .A(n1190), .B(n1191), .Z(\A2[478] ) );
  AND U1626 ( .A(n1192), .B(n1193), .Z(\A2[477] ) );
  AND U1627 ( .A(n1194), .B(n1195), .Z(\A2[476] ) );
  AND U1628 ( .A(n1196), .B(n1197), .Z(\A2[475] ) );
  AND U1629 ( .A(n1198), .B(n1199), .Z(\A2[474] ) );
  AND U1630 ( .A(n1200), .B(n1201), .Z(\A2[473] ) );
  AND U1631 ( .A(n1202), .B(n1203), .Z(\A2[472] ) );
  AND U1632 ( .A(n1204), .B(n1205), .Z(\A2[471] ) );
  AND U1633 ( .A(n1206), .B(n1207), .Z(\A2[470] ) );
  AND U1634 ( .A(n1208), .B(n1209), .Z(\A2[46] ) );
  AND U1635 ( .A(n1210), .B(n1211), .Z(\A2[469] ) );
  AND U1636 ( .A(n1212), .B(n1213), .Z(\A2[468] ) );
  AND U1637 ( .A(n1214), .B(n1215), .Z(\A2[467] ) );
  AND U1638 ( .A(n1216), .B(n1217), .Z(\A2[466] ) );
  AND U1639 ( .A(n1218), .B(n1219), .Z(\A2[465] ) );
  AND U1640 ( .A(n1220), .B(n1221), .Z(\A2[464] ) );
  AND U1641 ( .A(n1222), .B(n1223), .Z(\A2[463] ) );
  AND U1642 ( .A(n1224), .B(n1225), .Z(\A2[462] ) );
  AND U1643 ( .A(n1226), .B(n1227), .Z(\A2[461] ) );
  AND U1644 ( .A(n1228), .B(n1229), .Z(\A2[460] ) );
  AND U1645 ( .A(n1230), .B(n1231), .Z(\A2[45] ) );
  AND U1646 ( .A(n1232), .B(n1233), .Z(\A2[459] ) );
  AND U1647 ( .A(n1234), .B(n1235), .Z(\A2[458] ) );
  AND U1648 ( .A(n1236), .B(n1237), .Z(\A2[457] ) );
  AND U1649 ( .A(n1238), .B(n1239), .Z(\A2[456] ) );
  AND U1650 ( .A(n1240), .B(n1241), .Z(\A2[455] ) );
  AND U1651 ( .A(n1242), .B(n1243), .Z(\A2[454] ) );
  AND U1652 ( .A(n1244), .B(n1245), .Z(\A2[453] ) );
  AND U1653 ( .A(n1246), .B(n1247), .Z(\A2[452] ) );
  AND U1654 ( .A(n1248), .B(n1249), .Z(\A2[451] ) );
  AND U1655 ( .A(n1250), .B(n1251), .Z(\A2[450] ) );
  AND U1656 ( .A(n1252), .B(n1253), .Z(\A2[44] ) );
  AND U1657 ( .A(n1254), .B(n1255), .Z(\A2[449] ) );
  AND U1658 ( .A(n1256), .B(n1257), .Z(\A2[448] ) );
  AND U1659 ( .A(n1258), .B(n1259), .Z(\A2[447] ) );
  AND U1660 ( .A(n1260), .B(n1261), .Z(\A2[446] ) );
  AND U1661 ( .A(n1262), .B(n1263), .Z(\A2[445] ) );
  AND U1662 ( .A(n1264), .B(n1265), .Z(\A2[444] ) );
  AND U1663 ( .A(n1266), .B(n1267), .Z(\A2[443] ) );
  AND U1664 ( .A(n1268), .B(n1269), .Z(\A2[442] ) );
  AND U1665 ( .A(n1270), .B(n1271), .Z(\A2[441] ) );
  AND U1666 ( .A(n1272), .B(n1273), .Z(\A2[440] ) );
  AND U1667 ( .A(n1274), .B(n1275), .Z(\A2[43] ) );
  AND U1668 ( .A(n1276), .B(n1277), .Z(\A2[439] ) );
  AND U1669 ( .A(n1278), .B(n1279), .Z(\A2[438] ) );
  AND U1670 ( .A(n1280), .B(n1281), .Z(\A2[437] ) );
  AND U1671 ( .A(n1282), .B(n1283), .Z(\A2[436] ) );
  AND U1672 ( .A(n1284), .B(n1285), .Z(\A2[435] ) );
  AND U1673 ( .A(n1286), .B(n1287), .Z(\A2[434] ) );
  AND U1674 ( .A(n1288), .B(n1289), .Z(\A2[433] ) );
  AND U1675 ( .A(n1290), .B(n1291), .Z(\A2[432] ) );
  AND U1676 ( .A(n1292), .B(n1293), .Z(\A2[431] ) );
  AND U1677 ( .A(n1294), .B(n1295), .Z(\A2[430] ) );
  AND U1678 ( .A(n1296), .B(n1297), .Z(\A2[42] ) );
  AND U1679 ( .A(n1298), .B(n1299), .Z(\A2[429] ) );
  AND U1680 ( .A(n1300), .B(n1301), .Z(\A2[428] ) );
  AND U1681 ( .A(n1302), .B(n1303), .Z(\A2[427] ) );
  AND U1682 ( .A(n1304), .B(n1305), .Z(\A2[426] ) );
  AND U1683 ( .A(n1306), .B(n1307), .Z(\A2[425] ) );
  AND U1684 ( .A(n1308), .B(n1309), .Z(\A2[424] ) );
  AND U1685 ( .A(n1310), .B(n1311), .Z(\A2[423] ) );
  AND U1686 ( .A(n1312), .B(n1313), .Z(\A2[422] ) );
  AND U1687 ( .A(n1314), .B(n1315), .Z(\A2[421] ) );
  AND U1688 ( .A(n1316), .B(n1317), .Z(\A2[420] ) );
  AND U1689 ( .A(n1318), .B(n1319), .Z(\A2[41] ) );
  AND U1690 ( .A(n1320), .B(n1321), .Z(\A2[419] ) );
  AND U1691 ( .A(n1322), .B(n1323), .Z(\A2[418] ) );
  AND U1692 ( .A(n1324), .B(n1325), .Z(\A2[417] ) );
  AND U1693 ( .A(n1326), .B(n1327), .Z(\A2[416] ) );
  AND U1694 ( .A(n1328), .B(n1329), .Z(\A2[415] ) );
  AND U1695 ( .A(n1330), .B(n1331), .Z(\A2[414] ) );
  AND U1696 ( .A(n1332), .B(n1333), .Z(\A2[413] ) );
  AND U1697 ( .A(n1334), .B(n1335), .Z(\A2[412] ) );
  AND U1698 ( .A(n1336), .B(n1337), .Z(\A2[411] ) );
  AND U1699 ( .A(n1338), .B(n1339), .Z(\A2[410] ) );
  AND U1700 ( .A(n1340), .B(n1341), .Z(\A2[40] ) );
  AND U1701 ( .A(n1342), .B(n1343), .Z(\A2[409] ) );
  AND U1702 ( .A(n1344), .B(n1345), .Z(\A2[408] ) );
  AND U1703 ( .A(n1346), .B(n1347), .Z(\A2[407] ) );
  AND U1704 ( .A(n1348), .B(n1349), .Z(\A2[406] ) );
  AND U1705 ( .A(n1350), .B(n1351), .Z(\A2[405] ) );
  AND U1706 ( .A(n1352), .B(n1353), .Z(\A2[404] ) );
  AND U1707 ( .A(n1354), .B(n1355), .Z(\A2[403] ) );
  AND U1708 ( .A(n1356), .B(n1357), .Z(\A2[402] ) );
  AND U1709 ( .A(n1358), .B(n1359), .Z(\A2[401] ) );
  AND U1710 ( .A(n1360), .B(n1361), .Z(\A2[400] ) );
  AND U1711 ( .A(n1362), .B(n1363), .Z(\A2[3] ) );
  AND U1712 ( .A(n1364), .B(n1365), .Z(\A2[39] ) );
  AND U1713 ( .A(n1366), .B(n1367), .Z(\A2[399] ) );
  AND U1714 ( .A(n1368), .B(n1369), .Z(\A2[398] ) );
  AND U1715 ( .A(n1370), .B(n1371), .Z(\A2[397] ) );
  AND U1716 ( .A(n1372), .B(n1373), .Z(\A2[396] ) );
  AND U1717 ( .A(n1374), .B(n1375), .Z(\A2[395] ) );
  AND U1718 ( .A(n1376), .B(n1377), .Z(\A2[394] ) );
  AND U1719 ( .A(n1378), .B(n1379), .Z(\A2[393] ) );
  AND U1720 ( .A(n1380), .B(n1381), .Z(\A2[392] ) );
  AND U1721 ( .A(n1382), .B(n1383), .Z(\A2[391] ) );
  AND U1722 ( .A(n1384), .B(n1385), .Z(\A2[390] ) );
  AND U1723 ( .A(n1386), .B(n1387), .Z(\A2[38] ) );
  AND U1724 ( .A(n1388), .B(n1389), .Z(\A2[389] ) );
  AND U1725 ( .A(n1390), .B(n1391), .Z(\A2[388] ) );
  AND U1726 ( .A(n1392), .B(n1393), .Z(\A2[387] ) );
  AND U1727 ( .A(n1394), .B(n1395), .Z(\A2[386] ) );
  AND U1728 ( .A(n1396), .B(n1397), .Z(\A2[385] ) );
  AND U1729 ( .A(n1398), .B(n1399), .Z(\A2[384] ) );
  AND U1730 ( .A(n1400), .B(n1401), .Z(\A2[383] ) );
  AND U1731 ( .A(n1402), .B(n1403), .Z(\A2[382] ) );
  AND U1732 ( .A(n1404), .B(n1405), .Z(\A2[381] ) );
  AND U1733 ( .A(n1406), .B(n1407), .Z(\A2[380] ) );
  AND U1734 ( .A(n1408), .B(n1409), .Z(\A2[37] ) );
  AND U1735 ( .A(n1410), .B(n1411), .Z(\A2[379] ) );
  AND U1736 ( .A(n1412), .B(n1413), .Z(\A2[378] ) );
  AND U1737 ( .A(n1414), .B(n1415), .Z(\A2[377] ) );
  AND U1738 ( .A(n1416), .B(n1417), .Z(\A2[376] ) );
  AND U1739 ( .A(n1418), .B(n1419), .Z(\A2[375] ) );
  AND U1740 ( .A(n1420), .B(n1421), .Z(\A2[374] ) );
  AND U1741 ( .A(n1422), .B(n1423), .Z(\A2[373] ) );
  AND U1742 ( .A(n1424), .B(n1425), .Z(\A2[372] ) );
  AND U1743 ( .A(n1426), .B(n1427), .Z(\A2[371] ) );
  AND U1744 ( .A(n1428), .B(n1429), .Z(\A2[370] ) );
  AND U1745 ( .A(n1430), .B(n1431), .Z(\A2[36] ) );
  AND U1746 ( .A(n1432), .B(n1433), .Z(\A2[369] ) );
  AND U1747 ( .A(n1434), .B(n1435), .Z(\A2[368] ) );
  AND U1748 ( .A(n1436), .B(n1437), .Z(\A2[367] ) );
  AND U1749 ( .A(n1438), .B(n1439), .Z(\A2[366] ) );
  AND U1750 ( .A(n1440), .B(n1441), .Z(\A2[365] ) );
  AND U1751 ( .A(n1442), .B(n1443), .Z(\A2[364] ) );
  AND U1752 ( .A(n1444), .B(n1445), .Z(\A2[363] ) );
  AND U1753 ( .A(n1446), .B(n1447), .Z(\A2[362] ) );
  AND U1754 ( .A(n1448), .B(n1449), .Z(\A2[361] ) );
  AND U1755 ( .A(n1450), .B(n1451), .Z(\A2[360] ) );
  AND U1756 ( .A(n1452), .B(n1453), .Z(\A2[35] ) );
  AND U1757 ( .A(n1454), .B(n1455), .Z(\A2[359] ) );
  AND U1758 ( .A(n1456), .B(n1457), .Z(\A2[358] ) );
  AND U1759 ( .A(n1458), .B(n1459), .Z(\A2[357] ) );
  AND U1760 ( .A(n1460), .B(n1461), .Z(\A2[356] ) );
  AND U1761 ( .A(n1462), .B(n1463), .Z(\A2[355] ) );
  AND U1762 ( .A(n1464), .B(n1465), .Z(\A2[354] ) );
  AND U1763 ( .A(n1466), .B(n1467), .Z(\A2[353] ) );
  AND U1764 ( .A(n1468), .B(n1469), .Z(\A2[352] ) );
  AND U1765 ( .A(n1470), .B(n1471), .Z(\A2[351] ) );
  AND U1766 ( .A(n1472), .B(n1473), .Z(\A2[350] ) );
  AND U1767 ( .A(n1474), .B(n1475), .Z(\A2[34] ) );
  AND U1768 ( .A(n1476), .B(n1477), .Z(\A2[349] ) );
  AND U1769 ( .A(n1478), .B(n1479), .Z(\A2[348] ) );
  AND U1770 ( .A(n1480), .B(n1481), .Z(\A2[347] ) );
  AND U1771 ( .A(n1482), .B(n1483), .Z(\A2[346] ) );
  AND U1772 ( .A(n1484), .B(n1485), .Z(\A2[345] ) );
  AND U1773 ( .A(n1486), .B(n1487), .Z(\A2[344] ) );
  AND U1774 ( .A(n1488), .B(n1489), .Z(\A2[343] ) );
  AND U1775 ( .A(n1490), .B(n1491), .Z(\A2[342] ) );
  AND U1776 ( .A(n1492), .B(n1493), .Z(\A2[341] ) );
  AND U1777 ( .A(n1494), .B(n1495), .Z(\A2[340] ) );
  AND U1778 ( .A(n1496), .B(n1497), .Z(\A2[33] ) );
  AND U1779 ( .A(n1498), .B(n1499), .Z(\A2[339] ) );
  AND U1780 ( .A(n1500), .B(n1501), .Z(\A2[338] ) );
  AND U1781 ( .A(n1502), .B(n1503), .Z(\A2[337] ) );
  AND U1782 ( .A(n1504), .B(n1505), .Z(\A2[336] ) );
  AND U1783 ( .A(n1506), .B(n1507), .Z(\A2[335] ) );
  AND U1784 ( .A(n1508), .B(n1509), .Z(\A2[334] ) );
  AND U1785 ( .A(n1510), .B(n1511), .Z(\A2[333] ) );
  AND U1786 ( .A(n1512), .B(n1513), .Z(\A2[332] ) );
  AND U1787 ( .A(n1514), .B(n1515), .Z(\A2[331] ) );
  AND U1788 ( .A(n1516), .B(n1517), .Z(\A2[330] ) );
  AND U1789 ( .A(n1518), .B(n1519), .Z(\A2[32] ) );
  AND U1790 ( .A(n1520), .B(n1521), .Z(\A2[329] ) );
  AND U1791 ( .A(n1522), .B(n1523), .Z(\A2[328] ) );
  AND U1792 ( .A(n1524), .B(n1525), .Z(\A2[327] ) );
  AND U1793 ( .A(n1526), .B(n1527), .Z(\A2[326] ) );
  AND U1794 ( .A(n1528), .B(n1529), .Z(\A2[325] ) );
  AND U1795 ( .A(n1530), .B(n1531), .Z(\A2[324] ) );
  AND U1796 ( .A(n1532), .B(n1533), .Z(\A2[323] ) );
  AND U1797 ( .A(n1534), .B(n1535), .Z(\A2[322] ) );
  AND U1798 ( .A(n1536), .B(n1537), .Z(\A2[321] ) );
  AND U1799 ( .A(n1538), .B(n1539), .Z(\A2[320] ) );
  AND U1800 ( .A(n1540), .B(n1541), .Z(\A2[31] ) );
  AND U1801 ( .A(n1542), .B(n1543), .Z(\A2[319] ) );
  AND U1802 ( .A(n1544), .B(n1545), .Z(\A2[318] ) );
  AND U1803 ( .A(n1546), .B(n1547), .Z(\A2[317] ) );
  AND U1804 ( .A(n1548), .B(n1549), .Z(\A2[316] ) );
  AND U1805 ( .A(n1550), .B(n1551), .Z(\A2[315] ) );
  AND U1806 ( .A(n1552), .B(n1553), .Z(\A2[314] ) );
  AND U1807 ( .A(n1554), .B(n1555), .Z(\A2[313] ) );
  AND U1808 ( .A(n1556), .B(n1557), .Z(\A2[312] ) );
  AND U1809 ( .A(n1558), .B(n1559), .Z(\A2[311] ) );
  AND U1810 ( .A(n1560), .B(n1561), .Z(\A2[310] ) );
  AND U1811 ( .A(n1562), .B(n1563), .Z(\A2[30] ) );
  AND U1812 ( .A(n1564), .B(n1565), .Z(\A2[309] ) );
  AND U1813 ( .A(n1566), .B(n1567), .Z(\A2[308] ) );
  AND U1814 ( .A(n1568), .B(n1569), .Z(\A2[307] ) );
  AND U1815 ( .A(n1570), .B(n1571), .Z(\A2[306] ) );
  AND U1816 ( .A(n1572), .B(n1573), .Z(\A2[305] ) );
  AND U1817 ( .A(n1574), .B(n1575), .Z(\A2[304] ) );
  AND U1818 ( .A(n1576), .B(n1577), .Z(\A2[303] ) );
  AND U1819 ( .A(n1578), .B(n1579), .Z(\A2[302] ) );
  AND U1820 ( .A(n1580), .B(n1581), .Z(\A2[301] ) );
  AND U1821 ( .A(n1582), .B(n1583), .Z(\A2[300] ) );
  AND U1822 ( .A(n1584), .B(n1585), .Z(\A2[29] ) );
  AND U1823 ( .A(n1586), .B(n1587), .Z(\A2[299] ) );
  AND U1824 ( .A(n1588), .B(n1589), .Z(\A2[298] ) );
  AND U1825 ( .A(n1590), .B(n1591), .Z(\A2[297] ) );
  AND U1826 ( .A(n1592), .B(n1593), .Z(\A2[296] ) );
  AND U1827 ( .A(n1594), .B(n1595), .Z(\A2[295] ) );
  AND U1828 ( .A(n1596), .B(n1597), .Z(\A2[294] ) );
  AND U1829 ( .A(n1598), .B(n1599), .Z(\A2[293] ) );
  AND U1830 ( .A(n1600), .B(n1601), .Z(\A2[292] ) );
  AND U1831 ( .A(n1602), .B(n1603), .Z(\A2[291] ) );
  AND U1832 ( .A(n1604), .B(n1605), .Z(\A2[290] ) );
  AND U1833 ( .A(n1606), .B(n1607), .Z(\A2[28] ) );
  AND U1834 ( .A(n1608), .B(n1609), .Z(\A2[289] ) );
  AND U1835 ( .A(n1610), .B(n1611), .Z(\A2[288] ) );
  AND U1836 ( .A(n1612), .B(n1613), .Z(\A2[287] ) );
  AND U1837 ( .A(n1614), .B(n1615), .Z(\A2[286] ) );
  AND U1838 ( .A(n1616), .B(n1617), .Z(\A2[285] ) );
  AND U1839 ( .A(n1618), .B(n1619), .Z(\A2[284] ) );
  AND U1840 ( .A(n1620), .B(n1621), .Z(\A2[283] ) );
  AND U1841 ( .A(n1622), .B(n1623), .Z(\A2[282] ) );
  AND U1842 ( .A(n1624), .B(n1625), .Z(\A2[281] ) );
  AND U1843 ( .A(n1626), .B(n1627), .Z(\A2[280] ) );
  AND U1844 ( .A(n1628), .B(n1629), .Z(\A2[27] ) );
  AND U1845 ( .A(n1630), .B(n1631), .Z(\A2[279] ) );
  AND U1846 ( .A(n1632), .B(n1633), .Z(\A2[278] ) );
  AND U1847 ( .A(n1634), .B(n1635), .Z(\A2[277] ) );
  AND U1848 ( .A(n1636), .B(n1637), .Z(\A2[276] ) );
  AND U1849 ( .A(n1638), .B(n1639), .Z(\A2[275] ) );
  AND U1850 ( .A(n1640), .B(n1641), .Z(\A2[274] ) );
  AND U1851 ( .A(n1642), .B(n1643), .Z(\A2[273] ) );
  AND U1852 ( .A(n1644), .B(n1645), .Z(\A2[272] ) );
  AND U1853 ( .A(n1646), .B(n1647), .Z(\A2[271] ) );
  AND U1854 ( .A(n1648), .B(n1649), .Z(\A2[270] ) );
  AND U1855 ( .A(n1650), .B(n1651), .Z(\A2[26] ) );
  AND U1856 ( .A(n1652), .B(n1653), .Z(\A2[269] ) );
  AND U1857 ( .A(n1654), .B(n1655), .Z(\A2[268] ) );
  AND U1858 ( .A(n1656), .B(n1657), .Z(\A2[267] ) );
  AND U1859 ( .A(n1658), .B(n1659), .Z(\A2[266] ) );
  AND U1860 ( .A(n1660), .B(n1661), .Z(\A2[265] ) );
  AND U1861 ( .A(n1662), .B(n1663), .Z(\A2[264] ) );
  AND U1862 ( .A(n1664), .B(n1665), .Z(\A2[263] ) );
  AND U1863 ( .A(n1666), .B(n1667), .Z(\A2[262] ) );
  AND U1864 ( .A(n1668), .B(n1669), .Z(\A2[261] ) );
  AND U1865 ( .A(n1670), .B(n1671), .Z(\A2[260] ) );
  AND U1866 ( .A(n1672), .B(n1673), .Z(\A2[25] ) );
  AND U1867 ( .A(n1674), .B(n1675), .Z(\A2[259] ) );
  AND U1868 ( .A(n1676), .B(n1677), .Z(\A2[258] ) );
  AND U1869 ( .A(n1678), .B(n1679), .Z(\A2[257] ) );
  AND U1870 ( .A(n1680), .B(n1681), .Z(\A2[256] ) );
  AND U1871 ( .A(n1682), .B(n1683), .Z(\A2[255] ) );
  AND U1872 ( .A(n1684), .B(n1685), .Z(\A2[254] ) );
  AND U1873 ( .A(n1686), .B(n1687), .Z(\A2[253] ) );
  AND U1874 ( .A(n1688), .B(n1689), .Z(\A2[252] ) );
  AND U1875 ( .A(n1690), .B(n1691), .Z(\A2[251] ) );
  AND U1876 ( .A(n1692), .B(n1693), .Z(\A2[250] ) );
  AND U1877 ( .A(n1694), .B(n1695), .Z(\A2[24] ) );
  AND U1878 ( .A(n1696), .B(n1697), .Z(\A2[249] ) );
  AND U1879 ( .A(n1698), .B(n1699), .Z(\A2[248] ) );
  AND U1880 ( .A(n1700), .B(n1701), .Z(\A2[247] ) );
  AND U1881 ( .A(n1702), .B(n1703), .Z(\A2[246] ) );
  AND U1882 ( .A(n1704), .B(n1705), .Z(\A2[245] ) );
  AND U1883 ( .A(n1706), .B(n1707), .Z(\A2[244] ) );
  AND U1884 ( .A(n1708), .B(n1709), .Z(\A2[243] ) );
  AND U1885 ( .A(n1710), .B(n1711), .Z(\A2[242] ) );
  AND U1886 ( .A(n1712), .B(n1713), .Z(\A2[241] ) );
  AND U1887 ( .A(n1714), .B(n1715), .Z(\A2[240] ) );
  AND U1888 ( .A(n1716), .B(n1717), .Z(\A2[23] ) );
  AND U1889 ( .A(n1718), .B(n1719), .Z(\A2[239] ) );
  AND U1890 ( .A(n1720), .B(n1721), .Z(\A2[238] ) );
  AND U1891 ( .A(n1722), .B(n1723), .Z(\A2[237] ) );
  AND U1892 ( .A(n1724), .B(n1725), .Z(\A2[236] ) );
  AND U1893 ( .A(n1726), .B(n1727), .Z(\A2[235] ) );
  AND U1894 ( .A(n1728), .B(n1729), .Z(\A2[234] ) );
  AND U1895 ( .A(n1730), .B(n1731), .Z(\A2[233] ) );
  AND U1896 ( .A(n1732), .B(n1733), .Z(\A2[232] ) );
  AND U1897 ( .A(n1734), .B(n1735), .Z(\A2[231] ) );
  AND U1898 ( .A(n1736), .B(n1737), .Z(\A2[230] ) );
  AND U1899 ( .A(n1738), .B(n1739), .Z(\A2[22] ) );
  AND U1900 ( .A(n1740), .B(n1741), .Z(\A2[229] ) );
  AND U1901 ( .A(n1742), .B(n1743), .Z(\A2[228] ) );
  AND U1902 ( .A(n1744), .B(n1745), .Z(\A2[227] ) );
  AND U1903 ( .A(n1746), .B(n1747), .Z(\A2[226] ) );
  AND U1904 ( .A(n1748), .B(n1749), .Z(\A2[225] ) );
  AND U1905 ( .A(n1750), .B(n1751), .Z(\A2[224] ) );
  AND U1906 ( .A(n1752), .B(n1753), .Z(\A2[223] ) );
  AND U1907 ( .A(n1754), .B(n1755), .Z(\A2[222] ) );
  AND U1908 ( .A(n1756), .B(n1757), .Z(\A2[221] ) );
  AND U1909 ( .A(n1758), .B(n1759), .Z(\A2[220] ) );
  AND U1910 ( .A(n1760), .B(n1761), .Z(\A2[21] ) );
  AND U1911 ( .A(n1762), .B(n1763), .Z(\A2[219] ) );
  AND U1912 ( .A(n1764), .B(n1765), .Z(\A2[218] ) );
  AND U1913 ( .A(n1766), .B(n1767), .Z(\A2[217] ) );
  AND U1914 ( .A(n1768), .B(n1769), .Z(\A2[216] ) );
  AND U1915 ( .A(n1770), .B(n1771), .Z(\A2[215] ) );
  AND U1916 ( .A(n1772), .B(n1773), .Z(\A2[214] ) );
  AND U1917 ( .A(n1774), .B(n1775), .Z(\A2[213] ) );
  AND U1918 ( .A(n1776), .B(n1777), .Z(\A2[212] ) );
  AND U1919 ( .A(n1778), .B(n1779), .Z(\A2[211] ) );
  AND U1920 ( .A(n1780), .B(n1781), .Z(\A2[210] ) );
  AND U1921 ( .A(n1782), .B(n1783), .Z(\A2[20] ) );
  AND U1922 ( .A(n1784), .B(n1785), .Z(\A2[209] ) );
  AND U1923 ( .A(n1786), .B(n1787), .Z(\A2[208] ) );
  AND U1924 ( .A(n1788), .B(n1789), .Z(\A2[207] ) );
  AND U1925 ( .A(n1790), .B(n1791), .Z(\A2[206] ) );
  AND U1926 ( .A(n1792), .B(n1793), .Z(\A2[205] ) );
  AND U1927 ( .A(n1794), .B(n1795), .Z(\A2[204] ) );
  AND U1928 ( .A(n1796), .B(n1797), .Z(\A2[203] ) );
  AND U1929 ( .A(n1798), .B(n1799), .Z(\A2[202] ) );
  AND U1930 ( .A(n1800), .B(n1801), .Z(\A2[201] ) );
  AND U1931 ( .A(n1802), .B(n1803), .Z(\A2[200] ) );
  AND U1932 ( .A(n1804), .B(n1805), .Z(\A2[19] ) );
  AND U1933 ( .A(n1806), .B(n1807), .Z(\A2[199] ) );
  AND U1934 ( .A(n1808), .B(n1809), .Z(\A2[198] ) );
  AND U1935 ( .A(n1810), .B(n1811), .Z(\A2[197] ) );
  AND U1936 ( .A(n1812), .B(n1813), .Z(\A2[196] ) );
  AND U1937 ( .A(n1814), .B(n1815), .Z(\A2[195] ) );
  AND U1938 ( .A(n1816), .B(n1817), .Z(\A2[194] ) );
  AND U1939 ( .A(n1818), .B(n1819), .Z(\A2[193] ) );
  AND U1940 ( .A(n1820), .B(n1821), .Z(\A2[192] ) );
  AND U1941 ( .A(n1822), .B(n1823), .Z(\A2[191] ) );
  AND U1942 ( .A(n1824), .B(n1825), .Z(\A2[190] ) );
  AND U1943 ( .A(n1826), .B(n1827), .Z(\A2[18] ) );
  AND U1944 ( .A(n1828), .B(n1829), .Z(\A2[189] ) );
  AND U1945 ( .A(n1830), .B(n1831), .Z(\A2[188] ) );
  AND U1946 ( .A(n1832), .B(n1833), .Z(\A2[187] ) );
  AND U1947 ( .A(n1834), .B(n1835), .Z(\A2[186] ) );
  AND U1948 ( .A(n1836), .B(n1837), .Z(\A2[185] ) );
  AND U1949 ( .A(n1838), .B(n1839), .Z(\A2[184] ) );
  AND U1950 ( .A(n1840), .B(n1841), .Z(\A2[183] ) );
  AND U1951 ( .A(n1842), .B(n1843), .Z(\A2[182] ) );
  AND U1952 ( .A(n1844), .B(n1845), .Z(\A2[181] ) );
  AND U1953 ( .A(n1846), .B(n1847), .Z(\A2[180] ) );
  AND U1954 ( .A(n1848), .B(n1849), .Z(\A2[17] ) );
  AND U1955 ( .A(n1850), .B(n1851), .Z(\A2[179] ) );
  AND U1956 ( .A(n1852), .B(n1853), .Z(\A2[178] ) );
  AND U1957 ( .A(n1854), .B(n1855), .Z(\A2[177] ) );
  AND U1958 ( .A(n1856), .B(n1857), .Z(\A2[176] ) );
  AND U1959 ( .A(n1858), .B(n1859), .Z(\A2[175] ) );
  AND U1960 ( .A(n1860), .B(n1861), .Z(\A2[174] ) );
  AND U1961 ( .A(n1862), .B(n1863), .Z(\A2[173] ) );
  AND U1962 ( .A(n1864), .B(n1865), .Z(\A2[172] ) );
  AND U1963 ( .A(n1866), .B(n1867), .Z(\A2[171] ) );
  AND U1964 ( .A(n1868), .B(n1869), .Z(\A2[170] ) );
  AND U1965 ( .A(n1870), .B(n1871), .Z(\A2[16] ) );
  AND U1966 ( .A(n1872), .B(n1873), .Z(\A2[169] ) );
  AND U1967 ( .A(n1874), .B(n1875), .Z(\A2[168] ) );
  AND U1968 ( .A(n1876), .B(n1877), .Z(\A2[167] ) );
  AND U1969 ( .A(n1878), .B(n1879), .Z(\A2[166] ) );
  AND U1970 ( .A(n1880), .B(n1881), .Z(\A2[165] ) );
  AND U1971 ( .A(n1882), .B(n1883), .Z(\A2[164] ) );
  AND U1972 ( .A(n1884), .B(n1885), .Z(\A2[163] ) );
  AND U1973 ( .A(n1886), .B(n1887), .Z(\A2[162] ) );
  AND U1974 ( .A(n1888), .B(n1889), .Z(\A2[161] ) );
  AND U1975 ( .A(n1890), .B(n1891), .Z(\A2[160] ) );
  AND U1976 ( .A(n1892), .B(n1893), .Z(\A2[15] ) );
  AND U1977 ( .A(n1894), .B(n1895), .Z(\A2[159] ) );
  AND U1978 ( .A(n1896), .B(n1897), .Z(\A2[158] ) );
  AND U1979 ( .A(n1898), .B(n1899), .Z(\A2[157] ) );
  AND U1980 ( .A(n1900), .B(n1901), .Z(\A2[156] ) );
  AND U1981 ( .A(n1902), .B(n1903), .Z(\A2[155] ) );
  AND U1982 ( .A(n1904), .B(n1905), .Z(\A2[154] ) );
  AND U1983 ( .A(n1906), .B(n1907), .Z(\A2[153] ) );
  AND U1984 ( .A(n1908), .B(n1909), .Z(\A2[152] ) );
  AND U1985 ( .A(n1910), .B(n1911), .Z(\A2[151] ) );
  AND U1986 ( .A(n1912), .B(n1913), .Z(\A2[150] ) );
  AND U1987 ( .A(n1914), .B(n1915), .Z(\A2[14] ) );
  AND U1988 ( .A(n1916), .B(n1917), .Z(\A2[149] ) );
  AND U1989 ( .A(n1918), .B(n1919), .Z(\A2[148] ) );
  AND U1990 ( .A(n1920), .B(n1921), .Z(\A2[147] ) );
  AND U1991 ( .A(n1922), .B(n1923), .Z(\A2[146] ) );
  AND U1992 ( .A(n1924), .B(n1925), .Z(\A2[145] ) );
  AND U1993 ( .A(n1926), .B(n1927), .Z(\A2[144] ) );
  AND U1994 ( .A(n1928), .B(n1929), .Z(\A2[143] ) );
  AND U1995 ( .A(n1930), .B(n1931), .Z(\A2[142] ) );
  AND U1996 ( .A(n1932), .B(n1933), .Z(\A2[141] ) );
  AND U1997 ( .A(n1934), .B(n1935), .Z(\A2[140] ) );
  AND U1998 ( .A(n1936), .B(n1937), .Z(\A2[13] ) );
  AND U1999 ( .A(n1938), .B(n1939), .Z(\A2[139] ) );
  AND U2000 ( .A(n1940), .B(n1941), .Z(\A2[138] ) );
  AND U2001 ( .A(n1942), .B(n1943), .Z(\A2[137] ) );
  AND U2002 ( .A(n1944), .B(n1945), .Z(\A2[136] ) );
  AND U2003 ( .A(n1946), .B(n1947), .Z(\A2[135] ) );
  AND U2004 ( .A(n1948), .B(n1949), .Z(\A2[134] ) );
  AND U2005 ( .A(n1950), .B(n1951), .Z(\A2[133] ) );
  AND U2006 ( .A(n1952), .B(n1953), .Z(\A2[132] ) );
  AND U2007 ( .A(n1954), .B(n1955), .Z(\A2[131] ) );
  AND U2008 ( .A(n1956), .B(n1957), .Z(\A2[130] ) );
  AND U2009 ( .A(n1958), .B(n1959), .Z(\A2[12] ) );
  AND U2010 ( .A(n1960), .B(n1961), .Z(\A2[129] ) );
  AND U2011 ( .A(n1962), .B(n1963), .Z(\A2[128] ) );
  AND U2012 ( .A(n1964), .B(n1965), .Z(\A2[127] ) );
  AND U2013 ( .A(n1966), .B(n1967), .Z(\A2[126] ) );
  AND U2014 ( .A(n1968), .B(n1969), .Z(\A2[125] ) );
  AND U2015 ( .A(n1970), .B(n1971), .Z(\A2[124] ) );
  AND U2016 ( .A(n1972), .B(n1973), .Z(\A2[123] ) );
  AND U2017 ( .A(n1974), .B(n1975), .Z(\A2[122] ) );
  AND U2018 ( .A(n1976), .B(n1977), .Z(\A2[121] ) );
  AND U2019 ( .A(n1978), .B(n1979), .Z(\A2[120] ) );
  AND U2020 ( .A(n1980), .B(n1981), .Z(\A2[11] ) );
  AND U2021 ( .A(n1982), .B(n1983), .Z(\A2[119] ) );
  AND U2022 ( .A(n1984), .B(n1985), .Z(\A2[118] ) );
  AND U2023 ( .A(n1986), .B(n1987), .Z(\A2[117] ) );
  AND U2024 ( .A(n1988), .B(n1989), .Z(\A2[116] ) );
  AND U2025 ( .A(n1990), .B(n1991), .Z(\A2[115] ) );
  AND U2026 ( .A(n1992), .B(n1993), .Z(\A2[114] ) );
  AND U2027 ( .A(n1994), .B(n1995), .Z(\A2[113] ) );
  AND U2028 ( .A(n1996), .B(n1997), .Z(\A2[112] ) );
  AND U2029 ( .A(n1998), .B(n1999), .Z(\A2[111] ) );
  AND U2030 ( .A(n2000), .B(n2001), .Z(\A2[110] ) );
  AND U2031 ( .A(n2002), .B(n2003), .Z(\A2[10] ) );
  AND U2032 ( .A(n2004), .B(n2005), .Z(\A2[109] ) );
  AND U2033 ( .A(n2006), .B(n2007), .Z(\A2[108] ) );
  AND U2034 ( .A(n2008), .B(n2009), .Z(\A2[107] ) );
  AND U2035 ( .A(n2010), .B(n2011), .Z(\A2[106] ) );
  AND U2036 ( .A(n2012), .B(n2013), .Z(\A2[105] ) );
  AND U2037 ( .A(n2014), .B(n2015), .Z(\A2[104] ) );
  AND U2038 ( .A(n2016), .B(n2017), .Z(\A2[103] ) );
  AND U2039 ( .A(n2018), .B(n2019), .Z(\A2[102] ) );
  ANDN U2040 ( .B(n2020), .A(n26), .Z(\A2[1025] ) );
  AND U2041 ( .A(n2021), .B(n2022), .Z(\A2[1024] ) );
  AND U2042 ( .A(n2023), .B(n2024), .Z(\A2[1023] ) );
  AND U2043 ( .A(n2025), .B(n2026), .Z(\A2[1022] ) );
  AND U2044 ( .A(n2027), .B(n2028), .Z(\A2[1021] ) );
  AND U2045 ( .A(n2029), .B(n2030), .Z(\A2[1020] ) );
  AND U2046 ( .A(n2031), .B(n2032), .Z(\A2[101] ) );
  AND U2047 ( .A(n2033), .B(n2034), .Z(\A2[1019] ) );
  AND U2048 ( .A(n2035), .B(n2036), .Z(\A2[1018] ) );
  AND U2049 ( .A(n2037), .B(n2038), .Z(\A2[1017] ) );
  AND U2050 ( .A(n2039), .B(n2040), .Z(\A2[1016] ) );
  AND U2051 ( .A(n2041), .B(n2042), .Z(\A2[1015] ) );
  AND U2052 ( .A(n2043), .B(n2044), .Z(\A2[1014] ) );
  AND U2053 ( .A(n2045), .B(n2046), .Z(\A2[1013] ) );
  AND U2054 ( .A(n2047), .B(n2048), .Z(\A2[1012] ) );
  AND U2055 ( .A(n2049), .B(n2050), .Z(\A2[1011] ) );
  AND U2056 ( .A(n2051), .B(n2052), .Z(\A2[1010] ) );
  AND U2057 ( .A(n2053), .B(n2054), .Z(\A2[100] ) );
  AND U2058 ( .A(n2055), .B(n2056), .Z(\A2[1009] ) );
  AND U2059 ( .A(n2057), .B(n2058), .Z(\A2[1008] ) );
  AND U2060 ( .A(n2059), .B(n2060), .Z(\A2[1007] ) );
  AND U2061 ( .A(n2061), .B(n2062), .Z(\A2[1006] ) );
  AND U2062 ( .A(n2063), .B(n2064), .Z(\A2[1005] ) );
  AND U2063 ( .A(n2065), .B(n2066), .Z(\A2[1004] ) );
  AND U2064 ( .A(n2067), .B(n2068), .Z(\A2[1003] ) );
  AND U2065 ( .A(n2069), .B(n2070), .Z(\A2[1002] ) );
  AND U2066 ( .A(n2071), .B(n2072), .Z(\A2[1001] ) );
  AND U2067 ( .A(n2073), .B(n2074), .Z(\A2[1000] ) );
  XOR U2068 ( .A(n2003), .B(n2002), .Z(\A1[9] ) );
  XNOR U2069 ( .A(n2075), .B(n2076), .Z(n2002) );
  XOR U2070 ( .A(n2077), .B(n19), .Z(n2076) );
  NAND U2071 ( .A(n2078), .B(n2079), .Z(n2003) );
  NANDN U2072 ( .A(n2080), .B(n2081), .Z(n2079) );
  OR U2073 ( .A(n2082), .B(n2083), .Z(n2081) );
  XOR U2074 ( .A(n2054), .B(n2053), .Z(\A1[99] ) );
  XNOR U2075 ( .A(n2084), .B(n2085), .Z(n2053) );
  XOR U2076 ( .A(n2086), .B(n12), .Z(n2085) );
  NAND U2077 ( .A(n2087), .B(n2088), .Z(n2054) );
  NANDN U2078 ( .A(n2089), .B(n2090), .Z(n2088) );
  OR U2079 ( .A(n2091), .B(n2092), .Z(n2090) );
  XOR U2080 ( .A(n2074), .B(n2073), .Z(\A1[999] ) );
  XNOR U2081 ( .A(n2093), .B(n2094), .Z(n2073) );
  XOR U2082 ( .A(n2095), .B(n5), .Z(n2094) );
  NAND U2083 ( .A(n2096), .B(n2097), .Z(n2074) );
  NANDN U2084 ( .A(n2098), .B(n2099), .Z(n2097) );
  OR U2085 ( .A(n2100), .B(n2101), .Z(n2099) );
  XOR U2086 ( .A(n35), .B(n34), .Z(\A1[998] ) );
  XNOR U2087 ( .A(n2098), .B(n2102), .Z(n34) );
  XOR U2088 ( .A(n2100), .B(n2101), .Z(n2102) );
  NAND U2089 ( .A(n2103), .B(n2104), .Z(n2101) );
  NANDN U2090 ( .A(n2105), .B(n2106), .Z(n2104) );
  NANDN U2091 ( .A(n2107), .B(n2108), .Z(n2106) );
  NANDN U2092 ( .A(n2108), .B(n2107), .Z(n2103) );
  AND U2093 ( .A(B[997]), .B(A[3]), .Z(n2100) );
  XOR U2094 ( .A(n6), .B(n2109), .Z(n2098) );
  XOR U2095 ( .A(n2110), .B(n8), .Z(n2109) );
  NAND U2096 ( .A(n2111), .B(n2112), .Z(n35) );
  NANDN U2097 ( .A(n2113), .B(n2114), .Z(n2112) );
  OR U2098 ( .A(n2115), .B(n2116), .Z(n2114) );
  NANDN U2099 ( .A(n9), .B(n2115), .Z(n2111) );
  XOR U2100 ( .A(n37), .B(n36), .Z(\A1[997] ) );
  XNOR U2101 ( .A(n9), .B(n2117), .Z(n36) );
  XNOR U2102 ( .A(n2115), .B(n2113), .Z(n2117) );
  AND U2103 ( .A(n2118), .B(n2119), .Z(n2113) );
  NANDN U2104 ( .A(n2120), .B(n2121), .Z(n2119) );
  NANDN U2105 ( .A(n2122), .B(n2123), .Z(n2121) );
  AND U2106 ( .A(B[996]), .B(A[3]), .Z(n2115) );
  XOR U2107 ( .A(n2105), .B(n2124), .Z(n2116) );
  XOR U2108 ( .A(n2107), .B(n2108), .Z(n2124) );
  NAND U2109 ( .A(A[2]), .B(B[997]), .Z(n2108) );
  ANDN U2110 ( .B(n2125), .A(n2126), .Z(n2107) );
  AND U2111 ( .A(A[0]), .B(B[998]), .Z(n2125) );
  XNOR U2112 ( .A(n2127), .B(n2128), .Z(n2105) );
  NANDN U2113 ( .A(n10), .B(A[0]), .Z(n2128) );
  NAND U2114 ( .A(n2129), .B(n2130), .Z(n37) );
  NANDN U2115 ( .A(n2131), .B(n2132), .Z(n2130) );
  OR U2116 ( .A(n2133), .B(n2134), .Z(n2132) );
  NAND U2117 ( .A(n2134), .B(n2133), .Z(n2129) );
  XOR U2118 ( .A(n39), .B(n38), .Z(\A1[996] ) );
  XOR U2119 ( .A(n2134), .B(n2135), .Z(n38) );
  XNOR U2120 ( .A(n2133), .B(n2131), .Z(n2135) );
  AND U2121 ( .A(n2136), .B(n2137), .Z(n2131) );
  NANDN U2122 ( .A(n2138), .B(n2139), .Z(n2137) );
  NANDN U2123 ( .A(n2140), .B(n2141), .Z(n2139) );
  AND U2124 ( .A(B[995]), .B(A[3]), .Z(n2133) );
  XNOR U2125 ( .A(n2122), .B(n2142), .Z(n2134) );
  XNOR U2126 ( .A(n2120), .B(n2123), .Z(n2142) );
  NAND U2127 ( .A(A[2]), .B(B[996]), .Z(n2123) );
  NAND U2128 ( .A(n2143), .B(B[997]), .Z(n2120) );
  ANDN U2129 ( .B(A[0]), .A(n2144), .Z(n2143) );
  XOR U2130 ( .A(n2126), .B(n2145), .Z(n2122) );
  NAND U2131 ( .A(A[0]), .B(B[998]), .Z(n2145) );
  NAND U2132 ( .A(B[997]), .B(A[1]), .Z(n2126) );
  NAND U2133 ( .A(n2146), .B(n2147), .Z(n39) );
  NANDN U2134 ( .A(n2148), .B(n2149), .Z(n2147) );
  OR U2135 ( .A(n2150), .B(n2151), .Z(n2149) );
  NAND U2136 ( .A(n2151), .B(n2150), .Z(n2146) );
  XOR U2137 ( .A(n41), .B(n40), .Z(\A1[995] ) );
  XOR U2138 ( .A(n2151), .B(n2152), .Z(n40) );
  XNOR U2139 ( .A(n2150), .B(n2148), .Z(n2152) );
  AND U2140 ( .A(n2153), .B(n2154), .Z(n2148) );
  NANDN U2141 ( .A(n2155), .B(n2156), .Z(n2154) );
  NANDN U2142 ( .A(n2157), .B(n2158), .Z(n2156) );
  AND U2143 ( .A(B[994]), .B(A[3]), .Z(n2150) );
  XNOR U2144 ( .A(n2140), .B(n2159), .Z(n2151) );
  XNOR U2145 ( .A(n2138), .B(n2141), .Z(n2159) );
  NAND U2146 ( .A(A[2]), .B(B[995]), .Z(n2141) );
  NANDN U2147 ( .A(n2160), .B(n2161), .Z(n2138) );
  AND U2148 ( .A(A[0]), .B(B[996]), .Z(n2161) );
  XOR U2149 ( .A(n2144), .B(n2162), .Z(n2140) );
  NAND U2150 ( .A(A[0]), .B(B[997]), .Z(n2162) );
  NAND U2151 ( .A(B[996]), .B(A[1]), .Z(n2144) );
  NAND U2152 ( .A(n2163), .B(n2164), .Z(n41) );
  NANDN U2153 ( .A(n2165), .B(n2166), .Z(n2164) );
  OR U2154 ( .A(n2167), .B(n2168), .Z(n2166) );
  NAND U2155 ( .A(n2168), .B(n2167), .Z(n2163) );
  XOR U2156 ( .A(n43), .B(n42), .Z(\A1[994] ) );
  XOR U2157 ( .A(n2168), .B(n2169), .Z(n42) );
  XNOR U2158 ( .A(n2167), .B(n2165), .Z(n2169) );
  AND U2159 ( .A(n2170), .B(n2171), .Z(n2165) );
  NANDN U2160 ( .A(n2172), .B(n2173), .Z(n2171) );
  NANDN U2161 ( .A(n2174), .B(n2175), .Z(n2173) );
  AND U2162 ( .A(B[993]), .B(A[3]), .Z(n2167) );
  XNOR U2163 ( .A(n2157), .B(n2176), .Z(n2168) );
  XNOR U2164 ( .A(n2155), .B(n2158), .Z(n2176) );
  NAND U2165 ( .A(A[2]), .B(B[994]), .Z(n2158) );
  NANDN U2166 ( .A(n2177), .B(n2178), .Z(n2155) );
  AND U2167 ( .A(A[0]), .B(B[995]), .Z(n2178) );
  XOR U2168 ( .A(n2160), .B(n2179), .Z(n2157) );
  NAND U2169 ( .A(A[0]), .B(B[996]), .Z(n2179) );
  NAND U2170 ( .A(B[995]), .B(A[1]), .Z(n2160) );
  NAND U2171 ( .A(n2180), .B(n2181), .Z(n43) );
  NANDN U2172 ( .A(n2182), .B(n2183), .Z(n2181) );
  OR U2173 ( .A(n2184), .B(n2185), .Z(n2183) );
  NAND U2174 ( .A(n2185), .B(n2184), .Z(n2180) );
  XOR U2175 ( .A(n45), .B(n44), .Z(\A1[993] ) );
  XOR U2176 ( .A(n2185), .B(n2186), .Z(n44) );
  XNOR U2177 ( .A(n2184), .B(n2182), .Z(n2186) );
  AND U2178 ( .A(n2187), .B(n2188), .Z(n2182) );
  NANDN U2179 ( .A(n2189), .B(n2190), .Z(n2188) );
  NANDN U2180 ( .A(n2191), .B(n2192), .Z(n2190) );
  AND U2181 ( .A(B[992]), .B(A[3]), .Z(n2184) );
  XNOR U2182 ( .A(n2174), .B(n2193), .Z(n2185) );
  XNOR U2183 ( .A(n2172), .B(n2175), .Z(n2193) );
  NAND U2184 ( .A(A[2]), .B(B[993]), .Z(n2175) );
  NANDN U2185 ( .A(n2194), .B(n2195), .Z(n2172) );
  AND U2186 ( .A(A[0]), .B(B[994]), .Z(n2195) );
  XOR U2187 ( .A(n2177), .B(n2196), .Z(n2174) );
  NAND U2188 ( .A(A[0]), .B(B[995]), .Z(n2196) );
  NAND U2189 ( .A(B[994]), .B(A[1]), .Z(n2177) );
  NAND U2190 ( .A(n2197), .B(n2198), .Z(n45) );
  NANDN U2191 ( .A(n2199), .B(n2200), .Z(n2198) );
  OR U2192 ( .A(n2201), .B(n2202), .Z(n2200) );
  NAND U2193 ( .A(n2202), .B(n2201), .Z(n2197) );
  XOR U2194 ( .A(n47), .B(n46), .Z(\A1[992] ) );
  XOR U2195 ( .A(n2202), .B(n2203), .Z(n46) );
  XNOR U2196 ( .A(n2201), .B(n2199), .Z(n2203) );
  AND U2197 ( .A(n2204), .B(n2205), .Z(n2199) );
  NANDN U2198 ( .A(n2206), .B(n2207), .Z(n2205) );
  NANDN U2199 ( .A(n2208), .B(n2209), .Z(n2207) );
  AND U2200 ( .A(B[991]), .B(A[3]), .Z(n2201) );
  XNOR U2201 ( .A(n2191), .B(n2210), .Z(n2202) );
  XNOR U2202 ( .A(n2189), .B(n2192), .Z(n2210) );
  NAND U2203 ( .A(A[2]), .B(B[992]), .Z(n2192) );
  NANDN U2204 ( .A(n2211), .B(n2212), .Z(n2189) );
  AND U2205 ( .A(A[0]), .B(B[993]), .Z(n2212) );
  XOR U2206 ( .A(n2194), .B(n2213), .Z(n2191) );
  NAND U2207 ( .A(A[0]), .B(B[994]), .Z(n2213) );
  NAND U2208 ( .A(B[993]), .B(A[1]), .Z(n2194) );
  NAND U2209 ( .A(n2214), .B(n2215), .Z(n47) );
  NANDN U2210 ( .A(n2216), .B(n2217), .Z(n2215) );
  OR U2211 ( .A(n2218), .B(n2219), .Z(n2217) );
  NAND U2212 ( .A(n2219), .B(n2218), .Z(n2214) );
  XOR U2213 ( .A(n49), .B(n48), .Z(\A1[991] ) );
  XOR U2214 ( .A(n2219), .B(n2220), .Z(n48) );
  XNOR U2215 ( .A(n2218), .B(n2216), .Z(n2220) );
  AND U2216 ( .A(n2221), .B(n2222), .Z(n2216) );
  NANDN U2217 ( .A(n2223), .B(n2224), .Z(n2222) );
  NANDN U2218 ( .A(n2225), .B(n2226), .Z(n2224) );
  AND U2219 ( .A(B[990]), .B(A[3]), .Z(n2218) );
  XNOR U2220 ( .A(n2208), .B(n2227), .Z(n2219) );
  XNOR U2221 ( .A(n2206), .B(n2209), .Z(n2227) );
  NAND U2222 ( .A(A[2]), .B(B[991]), .Z(n2209) );
  NANDN U2223 ( .A(n2228), .B(n2229), .Z(n2206) );
  AND U2224 ( .A(A[0]), .B(B[992]), .Z(n2229) );
  XOR U2225 ( .A(n2211), .B(n2230), .Z(n2208) );
  NAND U2226 ( .A(A[0]), .B(B[993]), .Z(n2230) );
  NAND U2227 ( .A(B[992]), .B(A[1]), .Z(n2211) );
  NAND U2228 ( .A(n2231), .B(n2232), .Z(n49) );
  NANDN U2229 ( .A(n2233), .B(n2234), .Z(n2232) );
  OR U2230 ( .A(n2235), .B(n2236), .Z(n2234) );
  NAND U2231 ( .A(n2236), .B(n2235), .Z(n2231) );
  XOR U2232 ( .A(n51), .B(n50), .Z(\A1[990] ) );
  XOR U2233 ( .A(n2236), .B(n2237), .Z(n50) );
  XNOR U2234 ( .A(n2235), .B(n2233), .Z(n2237) );
  AND U2235 ( .A(n2238), .B(n2239), .Z(n2233) );
  NANDN U2236 ( .A(n2240), .B(n2241), .Z(n2239) );
  NANDN U2237 ( .A(n2242), .B(n2243), .Z(n2241) );
  AND U2238 ( .A(B[989]), .B(A[3]), .Z(n2235) );
  XNOR U2239 ( .A(n2225), .B(n2244), .Z(n2236) );
  XNOR U2240 ( .A(n2223), .B(n2226), .Z(n2244) );
  NAND U2241 ( .A(A[2]), .B(B[990]), .Z(n2226) );
  NANDN U2242 ( .A(n2245), .B(n2246), .Z(n2223) );
  AND U2243 ( .A(A[0]), .B(B[991]), .Z(n2246) );
  XOR U2244 ( .A(n2228), .B(n2247), .Z(n2225) );
  NAND U2245 ( .A(A[0]), .B(B[992]), .Z(n2247) );
  NAND U2246 ( .A(B[991]), .B(A[1]), .Z(n2228) );
  NAND U2247 ( .A(n2248), .B(n2249), .Z(n51) );
  NANDN U2248 ( .A(n2250), .B(n2251), .Z(n2249) );
  OR U2249 ( .A(n2252), .B(n2253), .Z(n2251) );
  NAND U2250 ( .A(n2253), .B(n2252), .Z(n2248) );
  XOR U2251 ( .A(n33), .B(n32), .Z(\A1[98] ) );
  XNOR U2252 ( .A(n2089), .B(n2254), .Z(n32) );
  XOR U2253 ( .A(n2091), .B(n2092), .Z(n2254) );
  NAND U2254 ( .A(n2255), .B(n2256), .Z(n2092) );
  NANDN U2255 ( .A(n2257), .B(n2258), .Z(n2256) );
  NANDN U2256 ( .A(n2259), .B(n2260), .Z(n2258) );
  NANDN U2257 ( .A(n2260), .B(n2259), .Z(n2255) );
  AND U2258 ( .A(B[97]), .B(A[3]), .Z(n2091) );
  XOR U2259 ( .A(n13), .B(n2261), .Z(n2089) );
  XOR U2260 ( .A(n2262), .B(n15), .Z(n2261) );
  NAND U2261 ( .A(n2263), .B(n2264), .Z(n33) );
  NANDN U2262 ( .A(n2265), .B(n2266), .Z(n2264) );
  OR U2263 ( .A(n2267), .B(n2268), .Z(n2266) );
  NANDN U2264 ( .A(n16), .B(n2267), .Z(n2263) );
  XOR U2265 ( .A(n53), .B(n52), .Z(\A1[989] ) );
  XOR U2266 ( .A(n2253), .B(n2269), .Z(n52) );
  XNOR U2267 ( .A(n2252), .B(n2250), .Z(n2269) );
  AND U2268 ( .A(n2270), .B(n2271), .Z(n2250) );
  NANDN U2269 ( .A(n2272), .B(n2273), .Z(n2271) );
  NANDN U2270 ( .A(n2274), .B(n2275), .Z(n2273) );
  AND U2271 ( .A(B[988]), .B(A[3]), .Z(n2252) );
  XNOR U2272 ( .A(n2242), .B(n2276), .Z(n2253) );
  XNOR U2273 ( .A(n2240), .B(n2243), .Z(n2276) );
  NAND U2274 ( .A(A[2]), .B(B[989]), .Z(n2243) );
  NANDN U2275 ( .A(n2277), .B(n2278), .Z(n2240) );
  AND U2276 ( .A(A[0]), .B(B[990]), .Z(n2278) );
  XOR U2277 ( .A(n2245), .B(n2279), .Z(n2242) );
  NAND U2278 ( .A(A[0]), .B(B[991]), .Z(n2279) );
  NAND U2279 ( .A(B[990]), .B(A[1]), .Z(n2245) );
  NAND U2280 ( .A(n2280), .B(n2281), .Z(n53) );
  NANDN U2281 ( .A(n2282), .B(n2283), .Z(n2281) );
  OR U2282 ( .A(n2284), .B(n2285), .Z(n2283) );
  NAND U2283 ( .A(n2285), .B(n2284), .Z(n2280) );
  XOR U2284 ( .A(n57), .B(n56), .Z(\A1[988] ) );
  XOR U2285 ( .A(n2285), .B(n2286), .Z(n56) );
  XNOR U2286 ( .A(n2284), .B(n2282), .Z(n2286) );
  AND U2287 ( .A(n2287), .B(n2288), .Z(n2282) );
  NANDN U2288 ( .A(n2289), .B(n2290), .Z(n2288) );
  NANDN U2289 ( .A(n2291), .B(n2292), .Z(n2290) );
  AND U2290 ( .A(B[987]), .B(A[3]), .Z(n2284) );
  XNOR U2291 ( .A(n2274), .B(n2293), .Z(n2285) );
  XNOR U2292 ( .A(n2272), .B(n2275), .Z(n2293) );
  NAND U2293 ( .A(A[2]), .B(B[988]), .Z(n2275) );
  NANDN U2294 ( .A(n2294), .B(n2295), .Z(n2272) );
  AND U2295 ( .A(A[0]), .B(B[989]), .Z(n2295) );
  XOR U2296 ( .A(n2277), .B(n2296), .Z(n2274) );
  NAND U2297 ( .A(A[0]), .B(B[990]), .Z(n2296) );
  NAND U2298 ( .A(B[989]), .B(A[1]), .Z(n2277) );
  NAND U2299 ( .A(n2297), .B(n2298), .Z(n57) );
  NANDN U2300 ( .A(n2299), .B(n2300), .Z(n2298) );
  OR U2301 ( .A(n2301), .B(n2302), .Z(n2300) );
  NAND U2302 ( .A(n2302), .B(n2301), .Z(n2297) );
  XOR U2303 ( .A(n59), .B(n58), .Z(\A1[987] ) );
  XOR U2304 ( .A(n2302), .B(n2303), .Z(n58) );
  XNOR U2305 ( .A(n2301), .B(n2299), .Z(n2303) );
  AND U2306 ( .A(n2304), .B(n2305), .Z(n2299) );
  NANDN U2307 ( .A(n2306), .B(n2307), .Z(n2305) );
  NANDN U2308 ( .A(n2308), .B(n2309), .Z(n2307) );
  AND U2309 ( .A(B[986]), .B(A[3]), .Z(n2301) );
  XNOR U2310 ( .A(n2291), .B(n2310), .Z(n2302) );
  XNOR U2311 ( .A(n2289), .B(n2292), .Z(n2310) );
  NAND U2312 ( .A(A[2]), .B(B[987]), .Z(n2292) );
  NANDN U2313 ( .A(n2311), .B(n2312), .Z(n2289) );
  AND U2314 ( .A(A[0]), .B(B[988]), .Z(n2312) );
  XOR U2315 ( .A(n2294), .B(n2313), .Z(n2291) );
  NAND U2316 ( .A(A[0]), .B(B[989]), .Z(n2313) );
  NAND U2317 ( .A(B[988]), .B(A[1]), .Z(n2294) );
  NAND U2318 ( .A(n2314), .B(n2315), .Z(n59) );
  NANDN U2319 ( .A(n2316), .B(n2317), .Z(n2315) );
  OR U2320 ( .A(n2318), .B(n2319), .Z(n2317) );
  NAND U2321 ( .A(n2319), .B(n2318), .Z(n2314) );
  XOR U2322 ( .A(n61), .B(n60), .Z(\A1[986] ) );
  XOR U2323 ( .A(n2319), .B(n2320), .Z(n60) );
  XNOR U2324 ( .A(n2318), .B(n2316), .Z(n2320) );
  AND U2325 ( .A(n2321), .B(n2322), .Z(n2316) );
  NANDN U2326 ( .A(n2323), .B(n2324), .Z(n2322) );
  NANDN U2327 ( .A(n2325), .B(n2326), .Z(n2324) );
  AND U2328 ( .A(B[985]), .B(A[3]), .Z(n2318) );
  XNOR U2329 ( .A(n2308), .B(n2327), .Z(n2319) );
  XNOR U2330 ( .A(n2306), .B(n2309), .Z(n2327) );
  NAND U2331 ( .A(A[2]), .B(B[986]), .Z(n2309) );
  NANDN U2332 ( .A(n2328), .B(n2329), .Z(n2306) );
  AND U2333 ( .A(A[0]), .B(B[987]), .Z(n2329) );
  XOR U2334 ( .A(n2311), .B(n2330), .Z(n2308) );
  NAND U2335 ( .A(A[0]), .B(B[988]), .Z(n2330) );
  NAND U2336 ( .A(B[987]), .B(A[1]), .Z(n2311) );
  NAND U2337 ( .A(n2331), .B(n2332), .Z(n61) );
  NANDN U2338 ( .A(n2333), .B(n2334), .Z(n2332) );
  OR U2339 ( .A(n2335), .B(n2336), .Z(n2334) );
  NAND U2340 ( .A(n2336), .B(n2335), .Z(n2331) );
  XOR U2341 ( .A(n63), .B(n62), .Z(\A1[985] ) );
  XOR U2342 ( .A(n2336), .B(n2337), .Z(n62) );
  XNOR U2343 ( .A(n2335), .B(n2333), .Z(n2337) );
  AND U2344 ( .A(n2338), .B(n2339), .Z(n2333) );
  NANDN U2345 ( .A(n2340), .B(n2341), .Z(n2339) );
  NANDN U2346 ( .A(n2342), .B(n2343), .Z(n2341) );
  AND U2347 ( .A(B[984]), .B(A[3]), .Z(n2335) );
  XNOR U2348 ( .A(n2325), .B(n2344), .Z(n2336) );
  XNOR U2349 ( .A(n2323), .B(n2326), .Z(n2344) );
  NAND U2350 ( .A(A[2]), .B(B[985]), .Z(n2326) );
  NANDN U2351 ( .A(n2345), .B(n2346), .Z(n2323) );
  AND U2352 ( .A(A[0]), .B(B[986]), .Z(n2346) );
  XOR U2353 ( .A(n2328), .B(n2347), .Z(n2325) );
  NAND U2354 ( .A(A[0]), .B(B[987]), .Z(n2347) );
  NAND U2355 ( .A(B[986]), .B(A[1]), .Z(n2328) );
  NAND U2356 ( .A(n2348), .B(n2349), .Z(n63) );
  NANDN U2357 ( .A(n2350), .B(n2351), .Z(n2349) );
  OR U2358 ( .A(n2352), .B(n2353), .Z(n2351) );
  NAND U2359 ( .A(n2353), .B(n2352), .Z(n2348) );
  XOR U2360 ( .A(n65), .B(n64), .Z(\A1[984] ) );
  XOR U2361 ( .A(n2353), .B(n2354), .Z(n64) );
  XNOR U2362 ( .A(n2352), .B(n2350), .Z(n2354) );
  AND U2363 ( .A(n2355), .B(n2356), .Z(n2350) );
  NANDN U2364 ( .A(n2357), .B(n2358), .Z(n2356) );
  NANDN U2365 ( .A(n2359), .B(n2360), .Z(n2358) );
  AND U2366 ( .A(B[983]), .B(A[3]), .Z(n2352) );
  XNOR U2367 ( .A(n2342), .B(n2361), .Z(n2353) );
  XNOR U2368 ( .A(n2340), .B(n2343), .Z(n2361) );
  NAND U2369 ( .A(A[2]), .B(B[984]), .Z(n2343) );
  NANDN U2370 ( .A(n2362), .B(n2363), .Z(n2340) );
  AND U2371 ( .A(A[0]), .B(B[985]), .Z(n2363) );
  XOR U2372 ( .A(n2345), .B(n2364), .Z(n2342) );
  NAND U2373 ( .A(A[0]), .B(B[986]), .Z(n2364) );
  NAND U2374 ( .A(B[985]), .B(A[1]), .Z(n2345) );
  NAND U2375 ( .A(n2365), .B(n2366), .Z(n65) );
  NANDN U2376 ( .A(n2367), .B(n2368), .Z(n2366) );
  OR U2377 ( .A(n2369), .B(n2370), .Z(n2368) );
  NAND U2378 ( .A(n2370), .B(n2369), .Z(n2365) );
  XOR U2379 ( .A(n67), .B(n66), .Z(\A1[983] ) );
  XOR U2380 ( .A(n2370), .B(n2371), .Z(n66) );
  XNOR U2381 ( .A(n2369), .B(n2367), .Z(n2371) );
  AND U2382 ( .A(n2372), .B(n2373), .Z(n2367) );
  NANDN U2383 ( .A(n2374), .B(n2375), .Z(n2373) );
  NANDN U2384 ( .A(n2376), .B(n2377), .Z(n2375) );
  AND U2385 ( .A(B[982]), .B(A[3]), .Z(n2369) );
  XNOR U2386 ( .A(n2359), .B(n2378), .Z(n2370) );
  XNOR U2387 ( .A(n2357), .B(n2360), .Z(n2378) );
  NAND U2388 ( .A(A[2]), .B(B[983]), .Z(n2360) );
  NANDN U2389 ( .A(n2379), .B(n2380), .Z(n2357) );
  AND U2390 ( .A(A[0]), .B(B[984]), .Z(n2380) );
  XOR U2391 ( .A(n2362), .B(n2381), .Z(n2359) );
  NAND U2392 ( .A(A[0]), .B(B[985]), .Z(n2381) );
  NAND U2393 ( .A(B[984]), .B(A[1]), .Z(n2362) );
  NAND U2394 ( .A(n2382), .B(n2383), .Z(n67) );
  NANDN U2395 ( .A(n2384), .B(n2385), .Z(n2383) );
  OR U2396 ( .A(n2386), .B(n2387), .Z(n2385) );
  NAND U2397 ( .A(n2387), .B(n2386), .Z(n2382) );
  XOR U2398 ( .A(n69), .B(n68), .Z(\A1[982] ) );
  XOR U2399 ( .A(n2387), .B(n2388), .Z(n68) );
  XNOR U2400 ( .A(n2386), .B(n2384), .Z(n2388) );
  AND U2401 ( .A(n2389), .B(n2390), .Z(n2384) );
  NANDN U2402 ( .A(n2391), .B(n2392), .Z(n2390) );
  NANDN U2403 ( .A(n2393), .B(n2394), .Z(n2392) );
  AND U2404 ( .A(B[981]), .B(A[3]), .Z(n2386) );
  XNOR U2405 ( .A(n2376), .B(n2395), .Z(n2387) );
  XNOR U2406 ( .A(n2374), .B(n2377), .Z(n2395) );
  NAND U2407 ( .A(A[2]), .B(B[982]), .Z(n2377) );
  NANDN U2408 ( .A(n2396), .B(n2397), .Z(n2374) );
  AND U2409 ( .A(A[0]), .B(B[983]), .Z(n2397) );
  XOR U2410 ( .A(n2379), .B(n2398), .Z(n2376) );
  NAND U2411 ( .A(A[0]), .B(B[984]), .Z(n2398) );
  NAND U2412 ( .A(B[983]), .B(A[1]), .Z(n2379) );
  NAND U2413 ( .A(n2399), .B(n2400), .Z(n69) );
  NANDN U2414 ( .A(n2401), .B(n2402), .Z(n2400) );
  OR U2415 ( .A(n2403), .B(n2404), .Z(n2402) );
  NAND U2416 ( .A(n2404), .B(n2403), .Z(n2399) );
  XOR U2417 ( .A(n71), .B(n70), .Z(\A1[981] ) );
  XOR U2418 ( .A(n2404), .B(n2405), .Z(n70) );
  XNOR U2419 ( .A(n2403), .B(n2401), .Z(n2405) );
  AND U2420 ( .A(n2406), .B(n2407), .Z(n2401) );
  NANDN U2421 ( .A(n2408), .B(n2409), .Z(n2407) );
  NANDN U2422 ( .A(n2410), .B(n2411), .Z(n2409) );
  AND U2423 ( .A(B[980]), .B(A[3]), .Z(n2403) );
  XNOR U2424 ( .A(n2393), .B(n2412), .Z(n2404) );
  XNOR U2425 ( .A(n2391), .B(n2394), .Z(n2412) );
  NAND U2426 ( .A(A[2]), .B(B[981]), .Z(n2394) );
  NANDN U2427 ( .A(n2413), .B(n2414), .Z(n2391) );
  AND U2428 ( .A(A[0]), .B(B[982]), .Z(n2414) );
  XOR U2429 ( .A(n2396), .B(n2415), .Z(n2393) );
  NAND U2430 ( .A(A[0]), .B(B[983]), .Z(n2415) );
  NAND U2431 ( .A(B[982]), .B(A[1]), .Z(n2396) );
  NAND U2432 ( .A(n2416), .B(n2417), .Z(n71) );
  NANDN U2433 ( .A(n2418), .B(n2419), .Z(n2417) );
  OR U2434 ( .A(n2420), .B(n2421), .Z(n2419) );
  NAND U2435 ( .A(n2421), .B(n2420), .Z(n2416) );
  XOR U2436 ( .A(n73), .B(n72), .Z(\A1[980] ) );
  XOR U2437 ( .A(n2421), .B(n2422), .Z(n72) );
  XNOR U2438 ( .A(n2420), .B(n2418), .Z(n2422) );
  AND U2439 ( .A(n2423), .B(n2424), .Z(n2418) );
  NANDN U2440 ( .A(n2425), .B(n2426), .Z(n2424) );
  NANDN U2441 ( .A(n2427), .B(n2428), .Z(n2426) );
  AND U2442 ( .A(B[979]), .B(A[3]), .Z(n2420) );
  XNOR U2443 ( .A(n2410), .B(n2429), .Z(n2421) );
  XNOR U2444 ( .A(n2408), .B(n2411), .Z(n2429) );
  NAND U2445 ( .A(A[2]), .B(B[980]), .Z(n2411) );
  NANDN U2446 ( .A(n2430), .B(n2431), .Z(n2408) );
  AND U2447 ( .A(A[0]), .B(B[981]), .Z(n2431) );
  XOR U2448 ( .A(n2413), .B(n2432), .Z(n2410) );
  NAND U2449 ( .A(A[0]), .B(B[982]), .Z(n2432) );
  NAND U2450 ( .A(B[981]), .B(A[1]), .Z(n2413) );
  NAND U2451 ( .A(n2433), .B(n2434), .Z(n73) );
  NANDN U2452 ( .A(n2435), .B(n2436), .Z(n2434) );
  OR U2453 ( .A(n2437), .B(n2438), .Z(n2436) );
  NAND U2454 ( .A(n2438), .B(n2437), .Z(n2433) );
  XOR U2455 ( .A(n55), .B(n54), .Z(\A1[97] ) );
  XNOR U2456 ( .A(n16), .B(n2439), .Z(n54) );
  XNOR U2457 ( .A(n2267), .B(n2265), .Z(n2439) );
  AND U2458 ( .A(n2440), .B(n2441), .Z(n2265) );
  NANDN U2459 ( .A(n2442), .B(n2443), .Z(n2441) );
  NANDN U2460 ( .A(n2444), .B(n2445), .Z(n2443) );
  AND U2461 ( .A(B[96]), .B(A[3]), .Z(n2267) );
  XOR U2462 ( .A(n2257), .B(n2446), .Z(n2268) );
  XOR U2463 ( .A(n2259), .B(n2260), .Z(n2446) );
  NAND U2464 ( .A(A[2]), .B(B[97]), .Z(n2260) );
  ANDN U2465 ( .B(n2447), .A(n2448), .Z(n2259) );
  AND U2466 ( .A(A[0]), .B(B[98]), .Z(n2447) );
  XNOR U2467 ( .A(n2449), .B(n2450), .Z(n2257) );
  NANDN U2468 ( .A(n17), .B(A[0]), .Z(n2450) );
  NAND U2469 ( .A(n2451), .B(n2452), .Z(n55) );
  NANDN U2470 ( .A(n2453), .B(n2454), .Z(n2452) );
  OR U2471 ( .A(n2455), .B(n2456), .Z(n2454) );
  NAND U2472 ( .A(n2456), .B(n2455), .Z(n2451) );
  XOR U2473 ( .A(n75), .B(n74), .Z(\A1[979] ) );
  XOR U2474 ( .A(n2438), .B(n2457), .Z(n74) );
  XNOR U2475 ( .A(n2437), .B(n2435), .Z(n2457) );
  AND U2476 ( .A(n2458), .B(n2459), .Z(n2435) );
  NANDN U2477 ( .A(n2460), .B(n2461), .Z(n2459) );
  NANDN U2478 ( .A(n2462), .B(n2463), .Z(n2461) );
  AND U2479 ( .A(B[978]), .B(A[3]), .Z(n2437) );
  XNOR U2480 ( .A(n2427), .B(n2464), .Z(n2438) );
  XNOR U2481 ( .A(n2425), .B(n2428), .Z(n2464) );
  NAND U2482 ( .A(A[2]), .B(B[979]), .Z(n2428) );
  NANDN U2483 ( .A(n2465), .B(n2466), .Z(n2425) );
  AND U2484 ( .A(A[0]), .B(B[980]), .Z(n2466) );
  XOR U2485 ( .A(n2430), .B(n2467), .Z(n2427) );
  NAND U2486 ( .A(A[0]), .B(B[981]), .Z(n2467) );
  NAND U2487 ( .A(B[980]), .B(A[1]), .Z(n2430) );
  NAND U2488 ( .A(n2468), .B(n2469), .Z(n75) );
  NANDN U2489 ( .A(n2470), .B(n2471), .Z(n2469) );
  OR U2490 ( .A(n2472), .B(n2473), .Z(n2471) );
  NAND U2491 ( .A(n2473), .B(n2472), .Z(n2468) );
  XOR U2492 ( .A(n79), .B(n78), .Z(\A1[978] ) );
  XOR U2493 ( .A(n2473), .B(n2474), .Z(n78) );
  XNOR U2494 ( .A(n2472), .B(n2470), .Z(n2474) );
  AND U2495 ( .A(n2475), .B(n2476), .Z(n2470) );
  NANDN U2496 ( .A(n2477), .B(n2478), .Z(n2476) );
  NANDN U2497 ( .A(n2479), .B(n2480), .Z(n2478) );
  AND U2498 ( .A(B[977]), .B(A[3]), .Z(n2472) );
  XNOR U2499 ( .A(n2462), .B(n2481), .Z(n2473) );
  XNOR U2500 ( .A(n2460), .B(n2463), .Z(n2481) );
  NAND U2501 ( .A(A[2]), .B(B[978]), .Z(n2463) );
  NANDN U2502 ( .A(n2482), .B(n2483), .Z(n2460) );
  AND U2503 ( .A(A[0]), .B(B[979]), .Z(n2483) );
  XOR U2504 ( .A(n2465), .B(n2484), .Z(n2462) );
  NAND U2505 ( .A(A[0]), .B(B[980]), .Z(n2484) );
  NAND U2506 ( .A(B[979]), .B(A[1]), .Z(n2465) );
  NAND U2507 ( .A(n2485), .B(n2486), .Z(n79) );
  NANDN U2508 ( .A(n2487), .B(n2488), .Z(n2486) );
  OR U2509 ( .A(n2489), .B(n2490), .Z(n2488) );
  NAND U2510 ( .A(n2490), .B(n2489), .Z(n2485) );
  XOR U2511 ( .A(n81), .B(n80), .Z(\A1[977] ) );
  XOR U2512 ( .A(n2490), .B(n2491), .Z(n80) );
  XNOR U2513 ( .A(n2489), .B(n2487), .Z(n2491) );
  AND U2514 ( .A(n2492), .B(n2493), .Z(n2487) );
  NANDN U2515 ( .A(n2494), .B(n2495), .Z(n2493) );
  NANDN U2516 ( .A(n2496), .B(n2497), .Z(n2495) );
  AND U2517 ( .A(B[976]), .B(A[3]), .Z(n2489) );
  XNOR U2518 ( .A(n2479), .B(n2498), .Z(n2490) );
  XNOR U2519 ( .A(n2477), .B(n2480), .Z(n2498) );
  NAND U2520 ( .A(A[2]), .B(B[977]), .Z(n2480) );
  NANDN U2521 ( .A(n2499), .B(n2500), .Z(n2477) );
  AND U2522 ( .A(A[0]), .B(B[978]), .Z(n2500) );
  XOR U2523 ( .A(n2482), .B(n2501), .Z(n2479) );
  NAND U2524 ( .A(A[0]), .B(B[979]), .Z(n2501) );
  NAND U2525 ( .A(B[978]), .B(A[1]), .Z(n2482) );
  NAND U2526 ( .A(n2502), .B(n2503), .Z(n81) );
  NANDN U2527 ( .A(n2504), .B(n2505), .Z(n2503) );
  OR U2528 ( .A(n2506), .B(n2507), .Z(n2505) );
  NAND U2529 ( .A(n2507), .B(n2506), .Z(n2502) );
  XOR U2530 ( .A(n83), .B(n82), .Z(\A1[976] ) );
  XOR U2531 ( .A(n2507), .B(n2508), .Z(n82) );
  XNOR U2532 ( .A(n2506), .B(n2504), .Z(n2508) );
  AND U2533 ( .A(n2509), .B(n2510), .Z(n2504) );
  NANDN U2534 ( .A(n2511), .B(n2512), .Z(n2510) );
  NANDN U2535 ( .A(n2513), .B(n2514), .Z(n2512) );
  AND U2536 ( .A(B[975]), .B(A[3]), .Z(n2506) );
  XNOR U2537 ( .A(n2496), .B(n2515), .Z(n2507) );
  XNOR U2538 ( .A(n2494), .B(n2497), .Z(n2515) );
  NAND U2539 ( .A(A[2]), .B(B[976]), .Z(n2497) );
  NANDN U2540 ( .A(n2516), .B(n2517), .Z(n2494) );
  AND U2541 ( .A(A[0]), .B(B[977]), .Z(n2517) );
  XOR U2542 ( .A(n2499), .B(n2518), .Z(n2496) );
  NAND U2543 ( .A(A[0]), .B(B[978]), .Z(n2518) );
  NAND U2544 ( .A(B[977]), .B(A[1]), .Z(n2499) );
  NAND U2545 ( .A(n2519), .B(n2520), .Z(n83) );
  NANDN U2546 ( .A(n2521), .B(n2522), .Z(n2520) );
  OR U2547 ( .A(n2523), .B(n2524), .Z(n2522) );
  NAND U2548 ( .A(n2524), .B(n2523), .Z(n2519) );
  XOR U2549 ( .A(n85), .B(n84), .Z(\A1[975] ) );
  XOR U2550 ( .A(n2524), .B(n2525), .Z(n84) );
  XNOR U2551 ( .A(n2523), .B(n2521), .Z(n2525) );
  AND U2552 ( .A(n2526), .B(n2527), .Z(n2521) );
  NANDN U2553 ( .A(n2528), .B(n2529), .Z(n2527) );
  NANDN U2554 ( .A(n2530), .B(n2531), .Z(n2529) );
  AND U2555 ( .A(B[974]), .B(A[3]), .Z(n2523) );
  XNOR U2556 ( .A(n2513), .B(n2532), .Z(n2524) );
  XNOR U2557 ( .A(n2511), .B(n2514), .Z(n2532) );
  NAND U2558 ( .A(A[2]), .B(B[975]), .Z(n2514) );
  NANDN U2559 ( .A(n2533), .B(n2534), .Z(n2511) );
  AND U2560 ( .A(A[0]), .B(B[976]), .Z(n2534) );
  XOR U2561 ( .A(n2516), .B(n2535), .Z(n2513) );
  NAND U2562 ( .A(A[0]), .B(B[977]), .Z(n2535) );
  NAND U2563 ( .A(B[976]), .B(A[1]), .Z(n2516) );
  NAND U2564 ( .A(n2536), .B(n2537), .Z(n85) );
  NANDN U2565 ( .A(n2538), .B(n2539), .Z(n2537) );
  OR U2566 ( .A(n2540), .B(n2541), .Z(n2539) );
  NAND U2567 ( .A(n2541), .B(n2540), .Z(n2536) );
  XOR U2568 ( .A(n87), .B(n86), .Z(\A1[974] ) );
  XOR U2569 ( .A(n2541), .B(n2542), .Z(n86) );
  XNOR U2570 ( .A(n2540), .B(n2538), .Z(n2542) );
  AND U2571 ( .A(n2543), .B(n2544), .Z(n2538) );
  NANDN U2572 ( .A(n2545), .B(n2546), .Z(n2544) );
  NANDN U2573 ( .A(n2547), .B(n2548), .Z(n2546) );
  AND U2574 ( .A(B[973]), .B(A[3]), .Z(n2540) );
  XNOR U2575 ( .A(n2530), .B(n2549), .Z(n2541) );
  XNOR U2576 ( .A(n2528), .B(n2531), .Z(n2549) );
  NAND U2577 ( .A(A[2]), .B(B[974]), .Z(n2531) );
  NANDN U2578 ( .A(n2550), .B(n2551), .Z(n2528) );
  AND U2579 ( .A(A[0]), .B(B[975]), .Z(n2551) );
  XOR U2580 ( .A(n2533), .B(n2552), .Z(n2530) );
  NAND U2581 ( .A(A[0]), .B(B[976]), .Z(n2552) );
  NAND U2582 ( .A(B[975]), .B(A[1]), .Z(n2533) );
  NAND U2583 ( .A(n2553), .B(n2554), .Z(n87) );
  NANDN U2584 ( .A(n2555), .B(n2556), .Z(n2554) );
  OR U2585 ( .A(n2557), .B(n2558), .Z(n2556) );
  NAND U2586 ( .A(n2558), .B(n2557), .Z(n2553) );
  XOR U2587 ( .A(n89), .B(n88), .Z(\A1[973] ) );
  XOR U2588 ( .A(n2558), .B(n2559), .Z(n88) );
  XNOR U2589 ( .A(n2557), .B(n2555), .Z(n2559) );
  AND U2590 ( .A(n2560), .B(n2561), .Z(n2555) );
  NANDN U2591 ( .A(n2562), .B(n2563), .Z(n2561) );
  NANDN U2592 ( .A(n2564), .B(n2565), .Z(n2563) );
  AND U2593 ( .A(B[972]), .B(A[3]), .Z(n2557) );
  XNOR U2594 ( .A(n2547), .B(n2566), .Z(n2558) );
  XNOR U2595 ( .A(n2545), .B(n2548), .Z(n2566) );
  NAND U2596 ( .A(A[2]), .B(B[973]), .Z(n2548) );
  NANDN U2597 ( .A(n2567), .B(n2568), .Z(n2545) );
  AND U2598 ( .A(A[0]), .B(B[974]), .Z(n2568) );
  XOR U2599 ( .A(n2550), .B(n2569), .Z(n2547) );
  NAND U2600 ( .A(A[0]), .B(B[975]), .Z(n2569) );
  NAND U2601 ( .A(B[974]), .B(A[1]), .Z(n2550) );
  NAND U2602 ( .A(n2570), .B(n2571), .Z(n89) );
  NANDN U2603 ( .A(n2572), .B(n2573), .Z(n2571) );
  OR U2604 ( .A(n2574), .B(n2575), .Z(n2573) );
  NAND U2605 ( .A(n2575), .B(n2574), .Z(n2570) );
  XOR U2606 ( .A(n91), .B(n90), .Z(\A1[972] ) );
  XOR U2607 ( .A(n2575), .B(n2576), .Z(n90) );
  XNOR U2608 ( .A(n2574), .B(n2572), .Z(n2576) );
  AND U2609 ( .A(n2577), .B(n2578), .Z(n2572) );
  NANDN U2610 ( .A(n2579), .B(n2580), .Z(n2578) );
  NANDN U2611 ( .A(n2581), .B(n2582), .Z(n2580) );
  AND U2612 ( .A(B[971]), .B(A[3]), .Z(n2574) );
  XNOR U2613 ( .A(n2564), .B(n2583), .Z(n2575) );
  XNOR U2614 ( .A(n2562), .B(n2565), .Z(n2583) );
  NAND U2615 ( .A(A[2]), .B(B[972]), .Z(n2565) );
  NANDN U2616 ( .A(n2584), .B(n2585), .Z(n2562) );
  AND U2617 ( .A(A[0]), .B(B[973]), .Z(n2585) );
  XOR U2618 ( .A(n2567), .B(n2586), .Z(n2564) );
  NAND U2619 ( .A(A[0]), .B(B[974]), .Z(n2586) );
  NAND U2620 ( .A(B[973]), .B(A[1]), .Z(n2567) );
  NAND U2621 ( .A(n2587), .B(n2588), .Z(n91) );
  NANDN U2622 ( .A(n2589), .B(n2590), .Z(n2588) );
  OR U2623 ( .A(n2591), .B(n2592), .Z(n2590) );
  NAND U2624 ( .A(n2592), .B(n2591), .Z(n2587) );
  XOR U2625 ( .A(n93), .B(n92), .Z(\A1[971] ) );
  XOR U2626 ( .A(n2592), .B(n2593), .Z(n92) );
  XNOR U2627 ( .A(n2591), .B(n2589), .Z(n2593) );
  AND U2628 ( .A(n2594), .B(n2595), .Z(n2589) );
  NANDN U2629 ( .A(n2596), .B(n2597), .Z(n2595) );
  NANDN U2630 ( .A(n2598), .B(n2599), .Z(n2597) );
  AND U2631 ( .A(B[970]), .B(A[3]), .Z(n2591) );
  XNOR U2632 ( .A(n2581), .B(n2600), .Z(n2592) );
  XNOR U2633 ( .A(n2579), .B(n2582), .Z(n2600) );
  NAND U2634 ( .A(A[2]), .B(B[971]), .Z(n2582) );
  NANDN U2635 ( .A(n2601), .B(n2602), .Z(n2579) );
  AND U2636 ( .A(A[0]), .B(B[972]), .Z(n2602) );
  XOR U2637 ( .A(n2584), .B(n2603), .Z(n2581) );
  NAND U2638 ( .A(A[0]), .B(B[973]), .Z(n2603) );
  NAND U2639 ( .A(B[972]), .B(A[1]), .Z(n2584) );
  NAND U2640 ( .A(n2604), .B(n2605), .Z(n93) );
  NANDN U2641 ( .A(n2606), .B(n2607), .Z(n2605) );
  OR U2642 ( .A(n2608), .B(n2609), .Z(n2607) );
  NAND U2643 ( .A(n2609), .B(n2608), .Z(n2604) );
  XOR U2644 ( .A(n95), .B(n94), .Z(\A1[970] ) );
  XOR U2645 ( .A(n2609), .B(n2610), .Z(n94) );
  XNOR U2646 ( .A(n2608), .B(n2606), .Z(n2610) );
  AND U2647 ( .A(n2611), .B(n2612), .Z(n2606) );
  NANDN U2648 ( .A(n2613), .B(n2614), .Z(n2612) );
  NANDN U2649 ( .A(n2615), .B(n2616), .Z(n2614) );
  AND U2650 ( .A(B[969]), .B(A[3]), .Z(n2608) );
  XNOR U2651 ( .A(n2598), .B(n2617), .Z(n2609) );
  XNOR U2652 ( .A(n2596), .B(n2599), .Z(n2617) );
  NAND U2653 ( .A(A[2]), .B(B[970]), .Z(n2599) );
  NANDN U2654 ( .A(n2618), .B(n2619), .Z(n2596) );
  AND U2655 ( .A(A[0]), .B(B[971]), .Z(n2619) );
  XOR U2656 ( .A(n2601), .B(n2620), .Z(n2598) );
  NAND U2657 ( .A(A[0]), .B(B[972]), .Z(n2620) );
  NAND U2658 ( .A(B[971]), .B(A[1]), .Z(n2601) );
  NAND U2659 ( .A(n2621), .B(n2622), .Z(n95) );
  NANDN U2660 ( .A(n2623), .B(n2624), .Z(n2622) );
  OR U2661 ( .A(n2625), .B(n2626), .Z(n2624) );
  NAND U2662 ( .A(n2626), .B(n2625), .Z(n2621) );
  XOR U2663 ( .A(n77), .B(n76), .Z(\A1[96] ) );
  XOR U2664 ( .A(n2456), .B(n2627), .Z(n76) );
  XNOR U2665 ( .A(n2455), .B(n2453), .Z(n2627) );
  AND U2666 ( .A(n2628), .B(n2629), .Z(n2453) );
  NANDN U2667 ( .A(n2630), .B(n2631), .Z(n2629) );
  NANDN U2668 ( .A(n2632), .B(n2633), .Z(n2631) );
  AND U2669 ( .A(B[95]), .B(A[3]), .Z(n2455) );
  XNOR U2670 ( .A(n2444), .B(n2634), .Z(n2456) );
  XNOR U2671 ( .A(n2442), .B(n2445), .Z(n2634) );
  NAND U2672 ( .A(A[2]), .B(B[96]), .Z(n2445) );
  NAND U2673 ( .A(n2635), .B(B[97]), .Z(n2442) );
  ANDN U2674 ( .B(A[0]), .A(n2636), .Z(n2635) );
  XOR U2675 ( .A(n2448), .B(n2637), .Z(n2444) );
  NAND U2676 ( .A(A[0]), .B(B[98]), .Z(n2637) );
  NAND U2677 ( .A(B[97]), .B(A[1]), .Z(n2448) );
  NAND U2678 ( .A(n2638), .B(n2639), .Z(n77) );
  NANDN U2679 ( .A(n2640), .B(n2641), .Z(n2639) );
  OR U2680 ( .A(n2642), .B(n2643), .Z(n2641) );
  NAND U2681 ( .A(n2643), .B(n2642), .Z(n2638) );
  XOR U2682 ( .A(n97), .B(n96), .Z(\A1[969] ) );
  XOR U2683 ( .A(n2626), .B(n2644), .Z(n96) );
  XNOR U2684 ( .A(n2625), .B(n2623), .Z(n2644) );
  AND U2685 ( .A(n2645), .B(n2646), .Z(n2623) );
  NANDN U2686 ( .A(n2647), .B(n2648), .Z(n2646) );
  NANDN U2687 ( .A(n2649), .B(n2650), .Z(n2648) );
  AND U2688 ( .A(B[968]), .B(A[3]), .Z(n2625) );
  XNOR U2689 ( .A(n2615), .B(n2651), .Z(n2626) );
  XNOR U2690 ( .A(n2613), .B(n2616), .Z(n2651) );
  NAND U2691 ( .A(A[2]), .B(B[969]), .Z(n2616) );
  NANDN U2692 ( .A(n2652), .B(n2653), .Z(n2613) );
  AND U2693 ( .A(A[0]), .B(B[970]), .Z(n2653) );
  XOR U2694 ( .A(n2618), .B(n2654), .Z(n2615) );
  NAND U2695 ( .A(A[0]), .B(B[971]), .Z(n2654) );
  NAND U2696 ( .A(B[970]), .B(A[1]), .Z(n2618) );
  NAND U2697 ( .A(n2655), .B(n2656), .Z(n97) );
  NANDN U2698 ( .A(n2657), .B(n2658), .Z(n2656) );
  OR U2699 ( .A(n2659), .B(n2660), .Z(n2658) );
  NAND U2700 ( .A(n2660), .B(n2659), .Z(n2655) );
  XOR U2701 ( .A(n101), .B(n100), .Z(\A1[968] ) );
  XOR U2702 ( .A(n2660), .B(n2661), .Z(n100) );
  XNOR U2703 ( .A(n2659), .B(n2657), .Z(n2661) );
  AND U2704 ( .A(n2662), .B(n2663), .Z(n2657) );
  NANDN U2705 ( .A(n2664), .B(n2665), .Z(n2663) );
  NANDN U2706 ( .A(n2666), .B(n2667), .Z(n2665) );
  AND U2707 ( .A(B[967]), .B(A[3]), .Z(n2659) );
  XNOR U2708 ( .A(n2649), .B(n2668), .Z(n2660) );
  XNOR U2709 ( .A(n2647), .B(n2650), .Z(n2668) );
  NAND U2710 ( .A(A[2]), .B(B[968]), .Z(n2650) );
  NANDN U2711 ( .A(n2669), .B(n2670), .Z(n2647) );
  AND U2712 ( .A(A[0]), .B(B[969]), .Z(n2670) );
  XOR U2713 ( .A(n2652), .B(n2671), .Z(n2649) );
  NAND U2714 ( .A(A[0]), .B(B[970]), .Z(n2671) );
  NAND U2715 ( .A(B[969]), .B(A[1]), .Z(n2652) );
  NAND U2716 ( .A(n2672), .B(n2673), .Z(n101) );
  NANDN U2717 ( .A(n2674), .B(n2675), .Z(n2673) );
  OR U2718 ( .A(n2676), .B(n2677), .Z(n2675) );
  NAND U2719 ( .A(n2677), .B(n2676), .Z(n2672) );
  XOR U2720 ( .A(n103), .B(n102), .Z(\A1[967] ) );
  XOR U2721 ( .A(n2677), .B(n2678), .Z(n102) );
  XNOR U2722 ( .A(n2676), .B(n2674), .Z(n2678) );
  AND U2723 ( .A(n2679), .B(n2680), .Z(n2674) );
  NANDN U2724 ( .A(n2681), .B(n2682), .Z(n2680) );
  NANDN U2725 ( .A(n2683), .B(n2684), .Z(n2682) );
  AND U2726 ( .A(B[966]), .B(A[3]), .Z(n2676) );
  XNOR U2727 ( .A(n2666), .B(n2685), .Z(n2677) );
  XNOR U2728 ( .A(n2664), .B(n2667), .Z(n2685) );
  NAND U2729 ( .A(A[2]), .B(B[967]), .Z(n2667) );
  NANDN U2730 ( .A(n2686), .B(n2687), .Z(n2664) );
  AND U2731 ( .A(A[0]), .B(B[968]), .Z(n2687) );
  XOR U2732 ( .A(n2669), .B(n2688), .Z(n2666) );
  NAND U2733 ( .A(A[0]), .B(B[969]), .Z(n2688) );
  NAND U2734 ( .A(B[968]), .B(A[1]), .Z(n2669) );
  NAND U2735 ( .A(n2689), .B(n2690), .Z(n103) );
  NANDN U2736 ( .A(n2691), .B(n2692), .Z(n2690) );
  OR U2737 ( .A(n2693), .B(n2694), .Z(n2692) );
  NAND U2738 ( .A(n2694), .B(n2693), .Z(n2689) );
  XOR U2739 ( .A(n105), .B(n104), .Z(\A1[966] ) );
  XOR U2740 ( .A(n2694), .B(n2695), .Z(n104) );
  XNOR U2741 ( .A(n2693), .B(n2691), .Z(n2695) );
  AND U2742 ( .A(n2696), .B(n2697), .Z(n2691) );
  NANDN U2743 ( .A(n2698), .B(n2699), .Z(n2697) );
  NANDN U2744 ( .A(n2700), .B(n2701), .Z(n2699) );
  AND U2745 ( .A(B[965]), .B(A[3]), .Z(n2693) );
  XNOR U2746 ( .A(n2683), .B(n2702), .Z(n2694) );
  XNOR U2747 ( .A(n2681), .B(n2684), .Z(n2702) );
  NAND U2748 ( .A(A[2]), .B(B[966]), .Z(n2684) );
  NANDN U2749 ( .A(n2703), .B(n2704), .Z(n2681) );
  AND U2750 ( .A(A[0]), .B(B[967]), .Z(n2704) );
  XOR U2751 ( .A(n2686), .B(n2705), .Z(n2683) );
  NAND U2752 ( .A(A[0]), .B(B[968]), .Z(n2705) );
  NAND U2753 ( .A(B[967]), .B(A[1]), .Z(n2686) );
  NAND U2754 ( .A(n2706), .B(n2707), .Z(n105) );
  NANDN U2755 ( .A(n2708), .B(n2709), .Z(n2707) );
  OR U2756 ( .A(n2710), .B(n2711), .Z(n2709) );
  NAND U2757 ( .A(n2711), .B(n2710), .Z(n2706) );
  XOR U2758 ( .A(n107), .B(n106), .Z(\A1[965] ) );
  XOR U2759 ( .A(n2711), .B(n2712), .Z(n106) );
  XNOR U2760 ( .A(n2710), .B(n2708), .Z(n2712) );
  AND U2761 ( .A(n2713), .B(n2714), .Z(n2708) );
  NANDN U2762 ( .A(n2715), .B(n2716), .Z(n2714) );
  NANDN U2763 ( .A(n2717), .B(n2718), .Z(n2716) );
  AND U2764 ( .A(B[964]), .B(A[3]), .Z(n2710) );
  XNOR U2765 ( .A(n2700), .B(n2719), .Z(n2711) );
  XNOR U2766 ( .A(n2698), .B(n2701), .Z(n2719) );
  NAND U2767 ( .A(A[2]), .B(B[965]), .Z(n2701) );
  NANDN U2768 ( .A(n2720), .B(n2721), .Z(n2698) );
  AND U2769 ( .A(A[0]), .B(B[966]), .Z(n2721) );
  XOR U2770 ( .A(n2703), .B(n2722), .Z(n2700) );
  NAND U2771 ( .A(A[0]), .B(B[967]), .Z(n2722) );
  NAND U2772 ( .A(B[966]), .B(A[1]), .Z(n2703) );
  NAND U2773 ( .A(n2723), .B(n2724), .Z(n107) );
  NANDN U2774 ( .A(n2725), .B(n2726), .Z(n2724) );
  OR U2775 ( .A(n2727), .B(n2728), .Z(n2726) );
  NAND U2776 ( .A(n2728), .B(n2727), .Z(n2723) );
  XOR U2777 ( .A(n109), .B(n108), .Z(\A1[964] ) );
  XOR U2778 ( .A(n2728), .B(n2729), .Z(n108) );
  XNOR U2779 ( .A(n2727), .B(n2725), .Z(n2729) );
  AND U2780 ( .A(n2730), .B(n2731), .Z(n2725) );
  NANDN U2781 ( .A(n2732), .B(n2733), .Z(n2731) );
  NANDN U2782 ( .A(n2734), .B(n2735), .Z(n2733) );
  AND U2783 ( .A(B[963]), .B(A[3]), .Z(n2727) );
  XNOR U2784 ( .A(n2717), .B(n2736), .Z(n2728) );
  XNOR U2785 ( .A(n2715), .B(n2718), .Z(n2736) );
  NAND U2786 ( .A(A[2]), .B(B[964]), .Z(n2718) );
  NANDN U2787 ( .A(n2737), .B(n2738), .Z(n2715) );
  AND U2788 ( .A(A[0]), .B(B[965]), .Z(n2738) );
  XOR U2789 ( .A(n2720), .B(n2739), .Z(n2717) );
  NAND U2790 ( .A(A[0]), .B(B[966]), .Z(n2739) );
  NAND U2791 ( .A(B[965]), .B(A[1]), .Z(n2720) );
  NAND U2792 ( .A(n2740), .B(n2741), .Z(n109) );
  NANDN U2793 ( .A(n2742), .B(n2743), .Z(n2741) );
  OR U2794 ( .A(n2744), .B(n2745), .Z(n2743) );
  NAND U2795 ( .A(n2745), .B(n2744), .Z(n2740) );
  XOR U2796 ( .A(n111), .B(n110), .Z(\A1[963] ) );
  XOR U2797 ( .A(n2745), .B(n2746), .Z(n110) );
  XNOR U2798 ( .A(n2744), .B(n2742), .Z(n2746) );
  AND U2799 ( .A(n2747), .B(n2748), .Z(n2742) );
  NANDN U2800 ( .A(n2749), .B(n2750), .Z(n2748) );
  NANDN U2801 ( .A(n2751), .B(n2752), .Z(n2750) );
  AND U2802 ( .A(B[962]), .B(A[3]), .Z(n2744) );
  XNOR U2803 ( .A(n2734), .B(n2753), .Z(n2745) );
  XNOR U2804 ( .A(n2732), .B(n2735), .Z(n2753) );
  NAND U2805 ( .A(A[2]), .B(B[963]), .Z(n2735) );
  NANDN U2806 ( .A(n2754), .B(n2755), .Z(n2732) );
  AND U2807 ( .A(A[0]), .B(B[964]), .Z(n2755) );
  XOR U2808 ( .A(n2737), .B(n2756), .Z(n2734) );
  NAND U2809 ( .A(A[0]), .B(B[965]), .Z(n2756) );
  NAND U2810 ( .A(B[964]), .B(A[1]), .Z(n2737) );
  NAND U2811 ( .A(n2757), .B(n2758), .Z(n111) );
  NANDN U2812 ( .A(n2759), .B(n2760), .Z(n2758) );
  OR U2813 ( .A(n2761), .B(n2762), .Z(n2760) );
  NAND U2814 ( .A(n2762), .B(n2761), .Z(n2757) );
  XOR U2815 ( .A(n113), .B(n112), .Z(\A1[962] ) );
  XOR U2816 ( .A(n2762), .B(n2763), .Z(n112) );
  XNOR U2817 ( .A(n2761), .B(n2759), .Z(n2763) );
  AND U2818 ( .A(n2764), .B(n2765), .Z(n2759) );
  NANDN U2819 ( .A(n2766), .B(n2767), .Z(n2765) );
  NANDN U2820 ( .A(n2768), .B(n2769), .Z(n2767) );
  AND U2821 ( .A(B[961]), .B(A[3]), .Z(n2761) );
  XNOR U2822 ( .A(n2751), .B(n2770), .Z(n2762) );
  XNOR U2823 ( .A(n2749), .B(n2752), .Z(n2770) );
  NAND U2824 ( .A(A[2]), .B(B[962]), .Z(n2752) );
  NANDN U2825 ( .A(n2771), .B(n2772), .Z(n2749) );
  AND U2826 ( .A(A[0]), .B(B[963]), .Z(n2772) );
  XOR U2827 ( .A(n2754), .B(n2773), .Z(n2751) );
  NAND U2828 ( .A(A[0]), .B(B[964]), .Z(n2773) );
  NAND U2829 ( .A(B[963]), .B(A[1]), .Z(n2754) );
  NAND U2830 ( .A(n2774), .B(n2775), .Z(n113) );
  NANDN U2831 ( .A(n2776), .B(n2777), .Z(n2775) );
  OR U2832 ( .A(n2778), .B(n2779), .Z(n2777) );
  NAND U2833 ( .A(n2779), .B(n2778), .Z(n2774) );
  XOR U2834 ( .A(n115), .B(n114), .Z(\A1[961] ) );
  XOR U2835 ( .A(n2779), .B(n2780), .Z(n114) );
  XNOR U2836 ( .A(n2778), .B(n2776), .Z(n2780) );
  AND U2837 ( .A(n2781), .B(n2782), .Z(n2776) );
  NANDN U2838 ( .A(n2783), .B(n2784), .Z(n2782) );
  NANDN U2839 ( .A(n2785), .B(n2786), .Z(n2784) );
  AND U2840 ( .A(B[960]), .B(A[3]), .Z(n2778) );
  XNOR U2841 ( .A(n2768), .B(n2787), .Z(n2779) );
  XNOR U2842 ( .A(n2766), .B(n2769), .Z(n2787) );
  NAND U2843 ( .A(A[2]), .B(B[961]), .Z(n2769) );
  NANDN U2844 ( .A(n2788), .B(n2789), .Z(n2766) );
  AND U2845 ( .A(A[0]), .B(B[962]), .Z(n2789) );
  XOR U2846 ( .A(n2771), .B(n2790), .Z(n2768) );
  NAND U2847 ( .A(A[0]), .B(B[963]), .Z(n2790) );
  NAND U2848 ( .A(B[962]), .B(A[1]), .Z(n2771) );
  NAND U2849 ( .A(n2791), .B(n2792), .Z(n115) );
  NANDN U2850 ( .A(n2793), .B(n2794), .Z(n2792) );
  OR U2851 ( .A(n2795), .B(n2796), .Z(n2794) );
  NAND U2852 ( .A(n2796), .B(n2795), .Z(n2791) );
  XOR U2853 ( .A(n117), .B(n116), .Z(\A1[960] ) );
  XOR U2854 ( .A(n2796), .B(n2797), .Z(n116) );
  XNOR U2855 ( .A(n2795), .B(n2793), .Z(n2797) );
  AND U2856 ( .A(n2798), .B(n2799), .Z(n2793) );
  NANDN U2857 ( .A(n2800), .B(n2801), .Z(n2799) );
  NANDN U2858 ( .A(n2802), .B(n2803), .Z(n2801) );
  AND U2859 ( .A(B[959]), .B(A[3]), .Z(n2795) );
  XNOR U2860 ( .A(n2785), .B(n2804), .Z(n2796) );
  XNOR U2861 ( .A(n2783), .B(n2786), .Z(n2804) );
  NAND U2862 ( .A(A[2]), .B(B[960]), .Z(n2786) );
  NANDN U2863 ( .A(n2805), .B(n2806), .Z(n2783) );
  AND U2864 ( .A(A[0]), .B(B[961]), .Z(n2806) );
  XOR U2865 ( .A(n2788), .B(n2807), .Z(n2785) );
  NAND U2866 ( .A(A[0]), .B(B[962]), .Z(n2807) );
  NAND U2867 ( .A(B[961]), .B(A[1]), .Z(n2788) );
  NAND U2868 ( .A(n2808), .B(n2809), .Z(n117) );
  NANDN U2869 ( .A(n2810), .B(n2811), .Z(n2809) );
  OR U2870 ( .A(n2812), .B(n2813), .Z(n2811) );
  NAND U2871 ( .A(n2813), .B(n2812), .Z(n2808) );
  XOR U2872 ( .A(n99), .B(n98), .Z(\A1[95] ) );
  XOR U2873 ( .A(n2643), .B(n2814), .Z(n98) );
  XNOR U2874 ( .A(n2642), .B(n2640), .Z(n2814) );
  AND U2875 ( .A(n2815), .B(n2816), .Z(n2640) );
  NANDN U2876 ( .A(n2817), .B(n2818), .Z(n2816) );
  NANDN U2877 ( .A(n2819), .B(n2820), .Z(n2818) );
  AND U2878 ( .A(B[94]), .B(A[3]), .Z(n2642) );
  XNOR U2879 ( .A(n2632), .B(n2821), .Z(n2643) );
  XNOR U2880 ( .A(n2630), .B(n2633), .Z(n2821) );
  NAND U2881 ( .A(A[2]), .B(B[95]), .Z(n2633) );
  NANDN U2882 ( .A(n2822), .B(n2823), .Z(n2630) );
  AND U2883 ( .A(A[0]), .B(B[96]), .Z(n2823) );
  XOR U2884 ( .A(n2636), .B(n2824), .Z(n2632) );
  NAND U2885 ( .A(A[0]), .B(B[97]), .Z(n2824) );
  NAND U2886 ( .A(B[96]), .B(A[1]), .Z(n2636) );
  NAND U2887 ( .A(n2825), .B(n2826), .Z(n99) );
  NANDN U2888 ( .A(n2827), .B(n2828), .Z(n2826) );
  OR U2889 ( .A(n2829), .B(n2830), .Z(n2828) );
  NAND U2890 ( .A(n2830), .B(n2829), .Z(n2825) );
  XOR U2891 ( .A(n119), .B(n118), .Z(\A1[959] ) );
  XOR U2892 ( .A(n2813), .B(n2831), .Z(n118) );
  XNOR U2893 ( .A(n2812), .B(n2810), .Z(n2831) );
  AND U2894 ( .A(n2832), .B(n2833), .Z(n2810) );
  NANDN U2895 ( .A(n2834), .B(n2835), .Z(n2833) );
  NANDN U2896 ( .A(n2836), .B(n2837), .Z(n2835) );
  AND U2897 ( .A(B[958]), .B(A[3]), .Z(n2812) );
  XNOR U2898 ( .A(n2802), .B(n2838), .Z(n2813) );
  XNOR U2899 ( .A(n2800), .B(n2803), .Z(n2838) );
  NAND U2900 ( .A(A[2]), .B(B[959]), .Z(n2803) );
  NANDN U2901 ( .A(n2839), .B(n2840), .Z(n2800) );
  AND U2902 ( .A(A[0]), .B(B[960]), .Z(n2840) );
  XOR U2903 ( .A(n2805), .B(n2841), .Z(n2802) );
  NAND U2904 ( .A(A[0]), .B(B[961]), .Z(n2841) );
  NAND U2905 ( .A(B[960]), .B(A[1]), .Z(n2805) );
  NAND U2906 ( .A(n2842), .B(n2843), .Z(n119) );
  NANDN U2907 ( .A(n2844), .B(n2845), .Z(n2843) );
  OR U2908 ( .A(n2846), .B(n2847), .Z(n2845) );
  NAND U2909 ( .A(n2847), .B(n2846), .Z(n2842) );
  XOR U2910 ( .A(n123), .B(n122), .Z(\A1[958] ) );
  XOR U2911 ( .A(n2847), .B(n2848), .Z(n122) );
  XNOR U2912 ( .A(n2846), .B(n2844), .Z(n2848) );
  AND U2913 ( .A(n2849), .B(n2850), .Z(n2844) );
  NANDN U2914 ( .A(n2851), .B(n2852), .Z(n2850) );
  NANDN U2915 ( .A(n2853), .B(n2854), .Z(n2852) );
  AND U2916 ( .A(B[957]), .B(A[3]), .Z(n2846) );
  XNOR U2917 ( .A(n2836), .B(n2855), .Z(n2847) );
  XNOR U2918 ( .A(n2834), .B(n2837), .Z(n2855) );
  NAND U2919 ( .A(A[2]), .B(B[958]), .Z(n2837) );
  NANDN U2920 ( .A(n2856), .B(n2857), .Z(n2834) );
  AND U2921 ( .A(A[0]), .B(B[959]), .Z(n2857) );
  XOR U2922 ( .A(n2839), .B(n2858), .Z(n2836) );
  NAND U2923 ( .A(A[0]), .B(B[960]), .Z(n2858) );
  NAND U2924 ( .A(B[959]), .B(A[1]), .Z(n2839) );
  NAND U2925 ( .A(n2859), .B(n2860), .Z(n123) );
  NANDN U2926 ( .A(n2861), .B(n2862), .Z(n2860) );
  OR U2927 ( .A(n2863), .B(n2864), .Z(n2862) );
  NAND U2928 ( .A(n2864), .B(n2863), .Z(n2859) );
  XOR U2929 ( .A(n125), .B(n124), .Z(\A1[957] ) );
  XOR U2930 ( .A(n2864), .B(n2865), .Z(n124) );
  XNOR U2931 ( .A(n2863), .B(n2861), .Z(n2865) );
  AND U2932 ( .A(n2866), .B(n2867), .Z(n2861) );
  NANDN U2933 ( .A(n2868), .B(n2869), .Z(n2867) );
  NANDN U2934 ( .A(n2870), .B(n2871), .Z(n2869) );
  AND U2935 ( .A(B[956]), .B(A[3]), .Z(n2863) );
  XNOR U2936 ( .A(n2853), .B(n2872), .Z(n2864) );
  XNOR U2937 ( .A(n2851), .B(n2854), .Z(n2872) );
  NAND U2938 ( .A(A[2]), .B(B[957]), .Z(n2854) );
  NANDN U2939 ( .A(n2873), .B(n2874), .Z(n2851) );
  AND U2940 ( .A(A[0]), .B(B[958]), .Z(n2874) );
  XOR U2941 ( .A(n2856), .B(n2875), .Z(n2853) );
  NAND U2942 ( .A(A[0]), .B(B[959]), .Z(n2875) );
  NAND U2943 ( .A(B[958]), .B(A[1]), .Z(n2856) );
  NAND U2944 ( .A(n2876), .B(n2877), .Z(n125) );
  NANDN U2945 ( .A(n2878), .B(n2879), .Z(n2877) );
  OR U2946 ( .A(n2880), .B(n2881), .Z(n2879) );
  NAND U2947 ( .A(n2881), .B(n2880), .Z(n2876) );
  XOR U2948 ( .A(n127), .B(n126), .Z(\A1[956] ) );
  XOR U2949 ( .A(n2881), .B(n2882), .Z(n126) );
  XNOR U2950 ( .A(n2880), .B(n2878), .Z(n2882) );
  AND U2951 ( .A(n2883), .B(n2884), .Z(n2878) );
  NANDN U2952 ( .A(n2885), .B(n2886), .Z(n2884) );
  NANDN U2953 ( .A(n2887), .B(n2888), .Z(n2886) );
  AND U2954 ( .A(B[955]), .B(A[3]), .Z(n2880) );
  XNOR U2955 ( .A(n2870), .B(n2889), .Z(n2881) );
  XNOR U2956 ( .A(n2868), .B(n2871), .Z(n2889) );
  NAND U2957 ( .A(A[2]), .B(B[956]), .Z(n2871) );
  NANDN U2958 ( .A(n2890), .B(n2891), .Z(n2868) );
  AND U2959 ( .A(A[0]), .B(B[957]), .Z(n2891) );
  XOR U2960 ( .A(n2873), .B(n2892), .Z(n2870) );
  NAND U2961 ( .A(A[0]), .B(B[958]), .Z(n2892) );
  NAND U2962 ( .A(B[957]), .B(A[1]), .Z(n2873) );
  NAND U2963 ( .A(n2893), .B(n2894), .Z(n127) );
  NANDN U2964 ( .A(n2895), .B(n2896), .Z(n2894) );
  OR U2965 ( .A(n2897), .B(n2898), .Z(n2896) );
  NAND U2966 ( .A(n2898), .B(n2897), .Z(n2893) );
  XOR U2967 ( .A(n129), .B(n128), .Z(\A1[955] ) );
  XOR U2968 ( .A(n2898), .B(n2899), .Z(n128) );
  XNOR U2969 ( .A(n2897), .B(n2895), .Z(n2899) );
  AND U2970 ( .A(n2900), .B(n2901), .Z(n2895) );
  NANDN U2971 ( .A(n2902), .B(n2903), .Z(n2901) );
  NANDN U2972 ( .A(n2904), .B(n2905), .Z(n2903) );
  AND U2973 ( .A(B[954]), .B(A[3]), .Z(n2897) );
  XNOR U2974 ( .A(n2887), .B(n2906), .Z(n2898) );
  XNOR U2975 ( .A(n2885), .B(n2888), .Z(n2906) );
  NAND U2976 ( .A(A[2]), .B(B[955]), .Z(n2888) );
  NANDN U2977 ( .A(n2907), .B(n2908), .Z(n2885) );
  AND U2978 ( .A(A[0]), .B(B[956]), .Z(n2908) );
  XOR U2979 ( .A(n2890), .B(n2909), .Z(n2887) );
  NAND U2980 ( .A(A[0]), .B(B[957]), .Z(n2909) );
  NAND U2981 ( .A(B[956]), .B(A[1]), .Z(n2890) );
  NAND U2982 ( .A(n2910), .B(n2911), .Z(n129) );
  NANDN U2983 ( .A(n2912), .B(n2913), .Z(n2911) );
  OR U2984 ( .A(n2914), .B(n2915), .Z(n2913) );
  NAND U2985 ( .A(n2915), .B(n2914), .Z(n2910) );
  XOR U2986 ( .A(n131), .B(n130), .Z(\A1[954] ) );
  XOR U2987 ( .A(n2915), .B(n2916), .Z(n130) );
  XNOR U2988 ( .A(n2914), .B(n2912), .Z(n2916) );
  AND U2989 ( .A(n2917), .B(n2918), .Z(n2912) );
  NANDN U2990 ( .A(n2919), .B(n2920), .Z(n2918) );
  NANDN U2991 ( .A(n2921), .B(n2922), .Z(n2920) );
  AND U2992 ( .A(B[953]), .B(A[3]), .Z(n2914) );
  XNOR U2993 ( .A(n2904), .B(n2923), .Z(n2915) );
  XNOR U2994 ( .A(n2902), .B(n2905), .Z(n2923) );
  NAND U2995 ( .A(A[2]), .B(B[954]), .Z(n2905) );
  NANDN U2996 ( .A(n2924), .B(n2925), .Z(n2902) );
  AND U2997 ( .A(A[0]), .B(B[955]), .Z(n2925) );
  XOR U2998 ( .A(n2907), .B(n2926), .Z(n2904) );
  NAND U2999 ( .A(A[0]), .B(B[956]), .Z(n2926) );
  NAND U3000 ( .A(B[955]), .B(A[1]), .Z(n2907) );
  NAND U3001 ( .A(n2927), .B(n2928), .Z(n131) );
  NANDN U3002 ( .A(n2929), .B(n2930), .Z(n2928) );
  OR U3003 ( .A(n2931), .B(n2932), .Z(n2930) );
  NAND U3004 ( .A(n2932), .B(n2931), .Z(n2927) );
  XOR U3005 ( .A(n133), .B(n132), .Z(\A1[953] ) );
  XOR U3006 ( .A(n2932), .B(n2933), .Z(n132) );
  XNOR U3007 ( .A(n2931), .B(n2929), .Z(n2933) );
  AND U3008 ( .A(n2934), .B(n2935), .Z(n2929) );
  NANDN U3009 ( .A(n2936), .B(n2937), .Z(n2935) );
  NANDN U3010 ( .A(n2938), .B(n2939), .Z(n2937) );
  AND U3011 ( .A(B[952]), .B(A[3]), .Z(n2931) );
  XNOR U3012 ( .A(n2921), .B(n2940), .Z(n2932) );
  XNOR U3013 ( .A(n2919), .B(n2922), .Z(n2940) );
  NAND U3014 ( .A(A[2]), .B(B[953]), .Z(n2922) );
  NANDN U3015 ( .A(n2941), .B(n2942), .Z(n2919) );
  AND U3016 ( .A(A[0]), .B(B[954]), .Z(n2942) );
  XOR U3017 ( .A(n2924), .B(n2943), .Z(n2921) );
  NAND U3018 ( .A(A[0]), .B(B[955]), .Z(n2943) );
  NAND U3019 ( .A(B[954]), .B(A[1]), .Z(n2924) );
  NAND U3020 ( .A(n2944), .B(n2945), .Z(n133) );
  NANDN U3021 ( .A(n2946), .B(n2947), .Z(n2945) );
  OR U3022 ( .A(n2948), .B(n2949), .Z(n2947) );
  NAND U3023 ( .A(n2949), .B(n2948), .Z(n2944) );
  XOR U3024 ( .A(n135), .B(n134), .Z(\A1[952] ) );
  XOR U3025 ( .A(n2949), .B(n2950), .Z(n134) );
  XNOR U3026 ( .A(n2948), .B(n2946), .Z(n2950) );
  AND U3027 ( .A(n2951), .B(n2952), .Z(n2946) );
  NANDN U3028 ( .A(n2953), .B(n2954), .Z(n2952) );
  NANDN U3029 ( .A(n2955), .B(n2956), .Z(n2954) );
  AND U3030 ( .A(B[951]), .B(A[3]), .Z(n2948) );
  XNOR U3031 ( .A(n2938), .B(n2957), .Z(n2949) );
  XNOR U3032 ( .A(n2936), .B(n2939), .Z(n2957) );
  NAND U3033 ( .A(A[2]), .B(B[952]), .Z(n2939) );
  NANDN U3034 ( .A(n2958), .B(n2959), .Z(n2936) );
  AND U3035 ( .A(A[0]), .B(B[953]), .Z(n2959) );
  XOR U3036 ( .A(n2941), .B(n2960), .Z(n2938) );
  NAND U3037 ( .A(A[0]), .B(B[954]), .Z(n2960) );
  NAND U3038 ( .A(B[953]), .B(A[1]), .Z(n2941) );
  NAND U3039 ( .A(n2961), .B(n2962), .Z(n135) );
  NANDN U3040 ( .A(n2963), .B(n2964), .Z(n2962) );
  OR U3041 ( .A(n2965), .B(n2966), .Z(n2964) );
  NAND U3042 ( .A(n2966), .B(n2965), .Z(n2961) );
  XOR U3043 ( .A(n137), .B(n136), .Z(\A1[951] ) );
  XOR U3044 ( .A(n2966), .B(n2967), .Z(n136) );
  XNOR U3045 ( .A(n2965), .B(n2963), .Z(n2967) );
  AND U3046 ( .A(n2968), .B(n2969), .Z(n2963) );
  NANDN U3047 ( .A(n2970), .B(n2971), .Z(n2969) );
  NANDN U3048 ( .A(n2972), .B(n2973), .Z(n2971) );
  AND U3049 ( .A(B[950]), .B(A[3]), .Z(n2965) );
  XNOR U3050 ( .A(n2955), .B(n2974), .Z(n2966) );
  XNOR U3051 ( .A(n2953), .B(n2956), .Z(n2974) );
  NAND U3052 ( .A(A[2]), .B(B[951]), .Z(n2956) );
  NANDN U3053 ( .A(n2975), .B(n2976), .Z(n2953) );
  AND U3054 ( .A(A[0]), .B(B[952]), .Z(n2976) );
  XOR U3055 ( .A(n2958), .B(n2977), .Z(n2955) );
  NAND U3056 ( .A(A[0]), .B(B[953]), .Z(n2977) );
  NAND U3057 ( .A(B[952]), .B(A[1]), .Z(n2958) );
  NAND U3058 ( .A(n2978), .B(n2979), .Z(n137) );
  NANDN U3059 ( .A(n2980), .B(n2981), .Z(n2979) );
  OR U3060 ( .A(n2982), .B(n2983), .Z(n2981) );
  NAND U3061 ( .A(n2983), .B(n2982), .Z(n2978) );
  XOR U3062 ( .A(n139), .B(n138), .Z(\A1[950] ) );
  XOR U3063 ( .A(n2983), .B(n2984), .Z(n138) );
  XNOR U3064 ( .A(n2982), .B(n2980), .Z(n2984) );
  AND U3065 ( .A(n2985), .B(n2986), .Z(n2980) );
  NANDN U3066 ( .A(n2987), .B(n2988), .Z(n2986) );
  NANDN U3067 ( .A(n2989), .B(n2990), .Z(n2988) );
  AND U3068 ( .A(B[949]), .B(A[3]), .Z(n2982) );
  XNOR U3069 ( .A(n2972), .B(n2991), .Z(n2983) );
  XNOR U3070 ( .A(n2970), .B(n2973), .Z(n2991) );
  NAND U3071 ( .A(A[2]), .B(B[950]), .Z(n2973) );
  NANDN U3072 ( .A(n2992), .B(n2993), .Z(n2970) );
  AND U3073 ( .A(A[0]), .B(B[951]), .Z(n2993) );
  XOR U3074 ( .A(n2975), .B(n2994), .Z(n2972) );
  NAND U3075 ( .A(A[0]), .B(B[952]), .Z(n2994) );
  NAND U3076 ( .A(B[951]), .B(A[1]), .Z(n2975) );
  NAND U3077 ( .A(n2995), .B(n2996), .Z(n139) );
  NANDN U3078 ( .A(n2997), .B(n2998), .Z(n2996) );
  OR U3079 ( .A(n2999), .B(n3000), .Z(n2998) );
  NAND U3080 ( .A(n3000), .B(n2999), .Z(n2995) );
  XOR U3081 ( .A(n121), .B(n120), .Z(\A1[94] ) );
  XOR U3082 ( .A(n2830), .B(n3001), .Z(n120) );
  XNOR U3083 ( .A(n2829), .B(n2827), .Z(n3001) );
  AND U3084 ( .A(n3002), .B(n3003), .Z(n2827) );
  NANDN U3085 ( .A(n3004), .B(n3005), .Z(n3003) );
  NANDN U3086 ( .A(n3006), .B(n3007), .Z(n3005) );
  AND U3087 ( .A(B[93]), .B(A[3]), .Z(n2829) );
  XNOR U3088 ( .A(n2819), .B(n3008), .Z(n2830) );
  XNOR U3089 ( .A(n2817), .B(n2820), .Z(n3008) );
  NAND U3090 ( .A(A[2]), .B(B[94]), .Z(n2820) );
  NANDN U3091 ( .A(n3009), .B(n3010), .Z(n2817) );
  AND U3092 ( .A(A[0]), .B(B[95]), .Z(n3010) );
  XOR U3093 ( .A(n2822), .B(n3011), .Z(n2819) );
  NAND U3094 ( .A(A[0]), .B(B[96]), .Z(n3011) );
  NAND U3095 ( .A(B[95]), .B(A[1]), .Z(n2822) );
  NAND U3096 ( .A(n3012), .B(n3013), .Z(n121) );
  NANDN U3097 ( .A(n3014), .B(n3015), .Z(n3013) );
  OR U3098 ( .A(n3016), .B(n3017), .Z(n3015) );
  NAND U3099 ( .A(n3017), .B(n3016), .Z(n3012) );
  XOR U3100 ( .A(n141), .B(n140), .Z(\A1[949] ) );
  XOR U3101 ( .A(n3000), .B(n3018), .Z(n140) );
  XNOR U3102 ( .A(n2999), .B(n2997), .Z(n3018) );
  AND U3103 ( .A(n3019), .B(n3020), .Z(n2997) );
  NANDN U3104 ( .A(n3021), .B(n3022), .Z(n3020) );
  NANDN U3105 ( .A(n3023), .B(n3024), .Z(n3022) );
  AND U3106 ( .A(B[948]), .B(A[3]), .Z(n2999) );
  XNOR U3107 ( .A(n2989), .B(n3025), .Z(n3000) );
  XNOR U3108 ( .A(n2987), .B(n2990), .Z(n3025) );
  NAND U3109 ( .A(A[2]), .B(B[949]), .Z(n2990) );
  NANDN U3110 ( .A(n3026), .B(n3027), .Z(n2987) );
  AND U3111 ( .A(A[0]), .B(B[950]), .Z(n3027) );
  XOR U3112 ( .A(n2992), .B(n3028), .Z(n2989) );
  NAND U3113 ( .A(A[0]), .B(B[951]), .Z(n3028) );
  NAND U3114 ( .A(B[950]), .B(A[1]), .Z(n2992) );
  NAND U3115 ( .A(n3029), .B(n3030), .Z(n141) );
  NANDN U3116 ( .A(n3031), .B(n3032), .Z(n3030) );
  OR U3117 ( .A(n3033), .B(n3034), .Z(n3032) );
  NAND U3118 ( .A(n3034), .B(n3033), .Z(n3029) );
  XOR U3119 ( .A(n145), .B(n144), .Z(\A1[948] ) );
  XOR U3120 ( .A(n3034), .B(n3035), .Z(n144) );
  XNOR U3121 ( .A(n3033), .B(n3031), .Z(n3035) );
  AND U3122 ( .A(n3036), .B(n3037), .Z(n3031) );
  NANDN U3123 ( .A(n3038), .B(n3039), .Z(n3037) );
  NANDN U3124 ( .A(n3040), .B(n3041), .Z(n3039) );
  AND U3125 ( .A(B[947]), .B(A[3]), .Z(n3033) );
  XNOR U3126 ( .A(n3023), .B(n3042), .Z(n3034) );
  XNOR U3127 ( .A(n3021), .B(n3024), .Z(n3042) );
  NAND U3128 ( .A(A[2]), .B(B[948]), .Z(n3024) );
  NANDN U3129 ( .A(n3043), .B(n3044), .Z(n3021) );
  AND U3130 ( .A(A[0]), .B(B[949]), .Z(n3044) );
  XOR U3131 ( .A(n3026), .B(n3045), .Z(n3023) );
  NAND U3132 ( .A(A[0]), .B(B[950]), .Z(n3045) );
  NAND U3133 ( .A(B[949]), .B(A[1]), .Z(n3026) );
  NAND U3134 ( .A(n3046), .B(n3047), .Z(n145) );
  NANDN U3135 ( .A(n3048), .B(n3049), .Z(n3047) );
  OR U3136 ( .A(n3050), .B(n3051), .Z(n3049) );
  NAND U3137 ( .A(n3051), .B(n3050), .Z(n3046) );
  XOR U3138 ( .A(n147), .B(n146), .Z(\A1[947] ) );
  XOR U3139 ( .A(n3051), .B(n3052), .Z(n146) );
  XNOR U3140 ( .A(n3050), .B(n3048), .Z(n3052) );
  AND U3141 ( .A(n3053), .B(n3054), .Z(n3048) );
  NANDN U3142 ( .A(n3055), .B(n3056), .Z(n3054) );
  NANDN U3143 ( .A(n3057), .B(n3058), .Z(n3056) );
  AND U3144 ( .A(B[946]), .B(A[3]), .Z(n3050) );
  XNOR U3145 ( .A(n3040), .B(n3059), .Z(n3051) );
  XNOR U3146 ( .A(n3038), .B(n3041), .Z(n3059) );
  NAND U3147 ( .A(A[2]), .B(B[947]), .Z(n3041) );
  NANDN U3148 ( .A(n3060), .B(n3061), .Z(n3038) );
  AND U3149 ( .A(A[0]), .B(B[948]), .Z(n3061) );
  XOR U3150 ( .A(n3043), .B(n3062), .Z(n3040) );
  NAND U3151 ( .A(A[0]), .B(B[949]), .Z(n3062) );
  NAND U3152 ( .A(B[948]), .B(A[1]), .Z(n3043) );
  NAND U3153 ( .A(n3063), .B(n3064), .Z(n147) );
  NANDN U3154 ( .A(n3065), .B(n3066), .Z(n3064) );
  OR U3155 ( .A(n3067), .B(n3068), .Z(n3066) );
  NAND U3156 ( .A(n3068), .B(n3067), .Z(n3063) );
  XOR U3157 ( .A(n149), .B(n148), .Z(\A1[946] ) );
  XOR U3158 ( .A(n3068), .B(n3069), .Z(n148) );
  XNOR U3159 ( .A(n3067), .B(n3065), .Z(n3069) );
  AND U3160 ( .A(n3070), .B(n3071), .Z(n3065) );
  NANDN U3161 ( .A(n3072), .B(n3073), .Z(n3071) );
  NANDN U3162 ( .A(n3074), .B(n3075), .Z(n3073) );
  AND U3163 ( .A(B[945]), .B(A[3]), .Z(n3067) );
  XNOR U3164 ( .A(n3057), .B(n3076), .Z(n3068) );
  XNOR U3165 ( .A(n3055), .B(n3058), .Z(n3076) );
  NAND U3166 ( .A(A[2]), .B(B[946]), .Z(n3058) );
  NANDN U3167 ( .A(n3077), .B(n3078), .Z(n3055) );
  AND U3168 ( .A(A[0]), .B(B[947]), .Z(n3078) );
  XOR U3169 ( .A(n3060), .B(n3079), .Z(n3057) );
  NAND U3170 ( .A(A[0]), .B(B[948]), .Z(n3079) );
  NAND U3171 ( .A(B[947]), .B(A[1]), .Z(n3060) );
  NAND U3172 ( .A(n3080), .B(n3081), .Z(n149) );
  NANDN U3173 ( .A(n3082), .B(n3083), .Z(n3081) );
  OR U3174 ( .A(n3084), .B(n3085), .Z(n3083) );
  NAND U3175 ( .A(n3085), .B(n3084), .Z(n3080) );
  XOR U3176 ( .A(n151), .B(n150), .Z(\A1[945] ) );
  XOR U3177 ( .A(n3085), .B(n3086), .Z(n150) );
  XNOR U3178 ( .A(n3084), .B(n3082), .Z(n3086) );
  AND U3179 ( .A(n3087), .B(n3088), .Z(n3082) );
  NANDN U3180 ( .A(n3089), .B(n3090), .Z(n3088) );
  NANDN U3181 ( .A(n3091), .B(n3092), .Z(n3090) );
  AND U3182 ( .A(B[944]), .B(A[3]), .Z(n3084) );
  XNOR U3183 ( .A(n3074), .B(n3093), .Z(n3085) );
  XNOR U3184 ( .A(n3072), .B(n3075), .Z(n3093) );
  NAND U3185 ( .A(A[2]), .B(B[945]), .Z(n3075) );
  NANDN U3186 ( .A(n3094), .B(n3095), .Z(n3072) );
  AND U3187 ( .A(A[0]), .B(B[946]), .Z(n3095) );
  XOR U3188 ( .A(n3077), .B(n3096), .Z(n3074) );
  NAND U3189 ( .A(A[0]), .B(B[947]), .Z(n3096) );
  NAND U3190 ( .A(B[946]), .B(A[1]), .Z(n3077) );
  NAND U3191 ( .A(n3097), .B(n3098), .Z(n151) );
  NANDN U3192 ( .A(n3099), .B(n3100), .Z(n3098) );
  OR U3193 ( .A(n3101), .B(n3102), .Z(n3100) );
  NAND U3194 ( .A(n3102), .B(n3101), .Z(n3097) );
  XOR U3195 ( .A(n153), .B(n152), .Z(\A1[944] ) );
  XOR U3196 ( .A(n3102), .B(n3103), .Z(n152) );
  XNOR U3197 ( .A(n3101), .B(n3099), .Z(n3103) );
  AND U3198 ( .A(n3104), .B(n3105), .Z(n3099) );
  NANDN U3199 ( .A(n3106), .B(n3107), .Z(n3105) );
  NANDN U3200 ( .A(n3108), .B(n3109), .Z(n3107) );
  AND U3201 ( .A(B[943]), .B(A[3]), .Z(n3101) );
  XNOR U3202 ( .A(n3091), .B(n3110), .Z(n3102) );
  XNOR U3203 ( .A(n3089), .B(n3092), .Z(n3110) );
  NAND U3204 ( .A(A[2]), .B(B[944]), .Z(n3092) );
  NANDN U3205 ( .A(n3111), .B(n3112), .Z(n3089) );
  AND U3206 ( .A(A[0]), .B(B[945]), .Z(n3112) );
  XOR U3207 ( .A(n3094), .B(n3113), .Z(n3091) );
  NAND U3208 ( .A(A[0]), .B(B[946]), .Z(n3113) );
  NAND U3209 ( .A(B[945]), .B(A[1]), .Z(n3094) );
  NAND U3210 ( .A(n3114), .B(n3115), .Z(n153) );
  NANDN U3211 ( .A(n3116), .B(n3117), .Z(n3115) );
  OR U3212 ( .A(n3118), .B(n3119), .Z(n3117) );
  NAND U3213 ( .A(n3119), .B(n3118), .Z(n3114) );
  XOR U3214 ( .A(n155), .B(n154), .Z(\A1[943] ) );
  XOR U3215 ( .A(n3119), .B(n3120), .Z(n154) );
  XNOR U3216 ( .A(n3118), .B(n3116), .Z(n3120) );
  AND U3217 ( .A(n3121), .B(n3122), .Z(n3116) );
  NANDN U3218 ( .A(n3123), .B(n3124), .Z(n3122) );
  NANDN U3219 ( .A(n3125), .B(n3126), .Z(n3124) );
  AND U3220 ( .A(B[942]), .B(A[3]), .Z(n3118) );
  XNOR U3221 ( .A(n3108), .B(n3127), .Z(n3119) );
  XNOR U3222 ( .A(n3106), .B(n3109), .Z(n3127) );
  NAND U3223 ( .A(A[2]), .B(B[943]), .Z(n3109) );
  NANDN U3224 ( .A(n3128), .B(n3129), .Z(n3106) );
  AND U3225 ( .A(A[0]), .B(B[944]), .Z(n3129) );
  XOR U3226 ( .A(n3111), .B(n3130), .Z(n3108) );
  NAND U3227 ( .A(A[0]), .B(B[945]), .Z(n3130) );
  NAND U3228 ( .A(B[944]), .B(A[1]), .Z(n3111) );
  NAND U3229 ( .A(n3131), .B(n3132), .Z(n155) );
  NANDN U3230 ( .A(n3133), .B(n3134), .Z(n3132) );
  OR U3231 ( .A(n3135), .B(n3136), .Z(n3134) );
  NAND U3232 ( .A(n3136), .B(n3135), .Z(n3131) );
  XOR U3233 ( .A(n157), .B(n156), .Z(\A1[942] ) );
  XOR U3234 ( .A(n3136), .B(n3137), .Z(n156) );
  XNOR U3235 ( .A(n3135), .B(n3133), .Z(n3137) );
  AND U3236 ( .A(n3138), .B(n3139), .Z(n3133) );
  NANDN U3237 ( .A(n3140), .B(n3141), .Z(n3139) );
  NANDN U3238 ( .A(n3142), .B(n3143), .Z(n3141) );
  AND U3239 ( .A(B[941]), .B(A[3]), .Z(n3135) );
  XNOR U3240 ( .A(n3125), .B(n3144), .Z(n3136) );
  XNOR U3241 ( .A(n3123), .B(n3126), .Z(n3144) );
  NAND U3242 ( .A(A[2]), .B(B[942]), .Z(n3126) );
  NANDN U3243 ( .A(n3145), .B(n3146), .Z(n3123) );
  AND U3244 ( .A(A[0]), .B(B[943]), .Z(n3146) );
  XOR U3245 ( .A(n3128), .B(n3147), .Z(n3125) );
  NAND U3246 ( .A(A[0]), .B(B[944]), .Z(n3147) );
  NAND U3247 ( .A(B[943]), .B(A[1]), .Z(n3128) );
  NAND U3248 ( .A(n3148), .B(n3149), .Z(n157) );
  NANDN U3249 ( .A(n3150), .B(n3151), .Z(n3149) );
  OR U3250 ( .A(n3152), .B(n3153), .Z(n3151) );
  NAND U3251 ( .A(n3153), .B(n3152), .Z(n3148) );
  XOR U3252 ( .A(n159), .B(n158), .Z(\A1[941] ) );
  XOR U3253 ( .A(n3153), .B(n3154), .Z(n158) );
  XNOR U3254 ( .A(n3152), .B(n3150), .Z(n3154) );
  AND U3255 ( .A(n3155), .B(n3156), .Z(n3150) );
  NANDN U3256 ( .A(n3157), .B(n3158), .Z(n3156) );
  NANDN U3257 ( .A(n3159), .B(n3160), .Z(n3158) );
  AND U3258 ( .A(B[940]), .B(A[3]), .Z(n3152) );
  XNOR U3259 ( .A(n3142), .B(n3161), .Z(n3153) );
  XNOR U3260 ( .A(n3140), .B(n3143), .Z(n3161) );
  NAND U3261 ( .A(A[2]), .B(B[941]), .Z(n3143) );
  NANDN U3262 ( .A(n3162), .B(n3163), .Z(n3140) );
  AND U3263 ( .A(A[0]), .B(B[942]), .Z(n3163) );
  XOR U3264 ( .A(n3145), .B(n3164), .Z(n3142) );
  NAND U3265 ( .A(A[0]), .B(B[943]), .Z(n3164) );
  NAND U3266 ( .A(B[942]), .B(A[1]), .Z(n3145) );
  NAND U3267 ( .A(n3165), .B(n3166), .Z(n159) );
  NANDN U3268 ( .A(n3167), .B(n3168), .Z(n3166) );
  OR U3269 ( .A(n3169), .B(n3170), .Z(n3168) );
  NAND U3270 ( .A(n3170), .B(n3169), .Z(n3165) );
  XOR U3271 ( .A(n161), .B(n160), .Z(\A1[940] ) );
  XOR U3272 ( .A(n3170), .B(n3171), .Z(n160) );
  XNOR U3273 ( .A(n3169), .B(n3167), .Z(n3171) );
  AND U3274 ( .A(n3172), .B(n3173), .Z(n3167) );
  NANDN U3275 ( .A(n3174), .B(n3175), .Z(n3173) );
  NANDN U3276 ( .A(n3176), .B(n3177), .Z(n3175) );
  AND U3277 ( .A(B[939]), .B(A[3]), .Z(n3169) );
  XNOR U3278 ( .A(n3159), .B(n3178), .Z(n3170) );
  XNOR U3279 ( .A(n3157), .B(n3160), .Z(n3178) );
  NAND U3280 ( .A(A[2]), .B(B[940]), .Z(n3160) );
  NANDN U3281 ( .A(n3179), .B(n3180), .Z(n3157) );
  AND U3282 ( .A(A[0]), .B(B[941]), .Z(n3180) );
  XOR U3283 ( .A(n3162), .B(n3181), .Z(n3159) );
  NAND U3284 ( .A(A[0]), .B(B[942]), .Z(n3181) );
  NAND U3285 ( .A(B[941]), .B(A[1]), .Z(n3162) );
  NAND U3286 ( .A(n3182), .B(n3183), .Z(n161) );
  NANDN U3287 ( .A(n3184), .B(n3185), .Z(n3183) );
  OR U3288 ( .A(n3186), .B(n3187), .Z(n3185) );
  NAND U3289 ( .A(n3187), .B(n3186), .Z(n3182) );
  XOR U3290 ( .A(n143), .B(n142), .Z(\A1[93] ) );
  XOR U3291 ( .A(n3017), .B(n3188), .Z(n142) );
  XNOR U3292 ( .A(n3016), .B(n3014), .Z(n3188) );
  AND U3293 ( .A(n3189), .B(n3190), .Z(n3014) );
  NANDN U3294 ( .A(n3191), .B(n3192), .Z(n3190) );
  NANDN U3295 ( .A(n3193), .B(n3194), .Z(n3192) );
  AND U3296 ( .A(B[92]), .B(A[3]), .Z(n3016) );
  XNOR U3297 ( .A(n3006), .B(n3195), .Z(n3017) );
  XNOR U3298 ( .A(n3004), .B(n3007), .Z(n3195) );
  NAND U3299 ( .A(A[2]), .B(B[93]), .Z(n3007) );
  NANDN U3300 ( .A(n3196), .B(n3197), .Z(n3004) );
  AND U3301 ( .A(A[0]), .B(B[94]), .Z(n3197) );
  XOR U3302 ( .A(n3009), .B(n3198), .Z(n3006) );
  NAND U3303 ( .A(A[0]), .B(B[95]), .Z(n3198) );
  NAND U3304 ( .A(B[94]), .B(A[1]), .Z(n3009) );
  NAND U3305 ( .A(n3199), .B(n3200), .Z(n143) );
  NANDN U3306 ( .A(n3201), .B(n3202), .Z(n3200) );
  OR U3307 ( .A(n3203), .B(n3204), .Z(n3202) );
  NAND U3308 ( .A(n3204), .B(n3203), .Z(n3199) );
  XOR U3309 ( .A(n163), .B(n162), .Z(\A1[939] ) );
  XOR U3310 ( .A(n3187), .B(n3205), .Z(n162) );
  XNOR U3311 ( .A(n3186), .B(n3184), .Z(n3205) );
  AND U3312 ( .A(n3206), .B(n3207), .Z(n3184) );
  NANDN U3313 ( .A(n3208), .B(n3209), .Z(n3207) );
  NANDN U3314 ( .A(n3210), .B(n3211), .Z(n3209) );
  AND U3315 ( .A(B[938]), .B(A[3]), .Z(n3186) );
  XNOR U3316 ( .A(n3176), .B(n3212), .Z(n3187) );
  XNOR U3317 ( .A(n3174), .B(n3177), .Z(n3212) );
  NAND U3318 ( .A(A[2]), .B(B[939]), .Z(n3177) );
  NANDN U3319 ( .A(n3213), .B(n3214), .Z(n3174) );
  AND U3320 ( .A(A[0]), .B(B[940]), .Z(n3214) );
  XOR U3321 ( .A(n3179), .B(n3215), .Z(n3176) );
  NAND U3322 ( .A(A[0]), .B(B[941]), .Z(n3215) );
  NAND U3323 ( .A(B[940]), .B(A[1]), .Z(n3179) );
  NAND U3324 ( .A(n3216), .B(n3217), .Z(n163) );
  NANDN U3325 ( .A(n3218), .B(n3219), .Z(n3217) );
  OR U3326 ( .A(n3220), .B(n3221), .Z(n3219) );
  NAND U3327 ( .A(n3221), .B(n3220), .Z(n3216) );
  XOR U3328 ( .A(n167), .B(n166), .Z(\A1[938] ) );
  XOR U3329 ( .A(n3221), .B(n3222), .Z(n166) );
  XNOR U3330 ( .A(n3220), .B(n3218), .Z(n3222) );
  AND U3331 ( .A(n3223), .B(n3224), .Z(n3218) );
  NANDN U3332 ( .A(n3225), .B(n3226), .Z(n3224) );
  NANDN U3333 ( .A(n3227), .B(n3228), .Z(n3226) );
  AND U3334 ( .A(B[937]), .B(A[3]), .Z(n3220) );
  XNOR U3335 ( .A(n3210), .B(n3229), .Z(n3221) );
  XNOR U3336 ( .A(n3208), .B(n3211), .Z(n3229) );
  NAND U3337 ( .A(A[2]), .B(B[938]), .Z(n3211) );
  NANDN U3338 ( .A(n3230), .B(n3231), .Z(n3208) );
  AND U3339 ( .A(A[0]), .B(B[939]), .Z(n3231) );
  XOR U3340 ( .A(n3213), .B(n3232), .Z(n3210) );
  NAND U3341 ( .A(A[0]), .B(B[940]), .Z(n3232) );
  NAND U3342 ( .A(B[939]), .B(A[1]), .Z(n3213) );
  NAND U3343 ( .A(n3233), .B(n3234), .Z(n167) );
  NANDN U3344 ( .A(n3235), .B(n3236), .Z(n3234) );
  OR U3345 ( .A(n3237), .B(n3238), .Z(n3236) );
  NAND U3346 ( .A(n3238), .B(n3237), .Z(n3233) );
  XOR U3347 ( .A(n169), .B(n168), .Z(\A1[937] ) );
  XOR U3348 ( .A(n3238), .B(n3239), .Z(n168) );
  XNOR U3349 ( .A(n3237), .B(n3235), .Z(n3239) );
  AND U3350 ( .A(n3240), .B(n3241), .Z(n3235) );
  NANDN U3351 ( .A(n3242), .B(n3243), .Z(n3241) );
  NANDN U3352 ( .A(n3244), .B(n3245), .Z(n3243) );
  AND U3353 ( .A(B[936]), .B(A[3]), .Z(n3237) );
  XNOR U3354 ( .A(n3227), .B(n3246), .Z(n3238) );
  XNOR U3355 ( .A(n3225), .B(n3228), .Z(n3246) );
  NAND U3356 ( .A(A[2]), .B(B[937]), .Z(n3228) );
  NANDN U3357 ( .A(n3247), .B(n3248), .Z(n3225) );
  AND U3358 ( .A(A[0]), .B(B[938]), .Z(n3248) );
  XOR U3359 ( .A(n3230), .B(n3249), .Z(n3227) );
  NAND U3360 ( .A(A[0]), .B(B[939]), .Z(n3249) );
  NAND U3361 ( .A(B[938]), .B(A[1]), .Z(n3230) );
  NAND U3362 ( .A(n3250), .B(n3251), .Z(n169) );
  NANDN U3363 ( .A(n3252), .B(n3253), .Z(n3251) );
  OR U3364 ( .A(n3254), .B(n3255), .Z(n3253) );
  NAND U3365 ( .A(n3255), .B(n3254), .Z(n3250) );
  XOR U3366 ( .A(n171), .B(n170), .Z(\A1[936] ) );
  XOR U3367 ( .A(n3255), .B(n3256), .Z(n170) );
  XNOR U3368 ( .A(n3254), .B(n3252), .Z(n3256) );
  AND U3369 ( .A(n3257), .B(n3258), .Z(n3252) );
  NANDN U3370 ( .A(n3259), .B(n3260), .Z(n3258) );
  NANDN U3371 ( .A(n3261), .B(n3262), .Z(n3260) );
  AND U3372 ( .A(B[935]), .B(A[3]), .Z(n3254) );
  XNOR U3373 ( .A(n3244), .B(n3263), .Z(n3255) );
  XNOR U3374 ( .A(n3242), .B(n3245), .Z(n3263) );
  NAND U3375 ( .A(A[2]), .B(B[936]), .Z(n3245) );
  NANDN U3376 ( .A(n3264), .B(n3265), .Z(n3242) );
  AND U3377 ( .A(A[0]), .B(B[937]), .Z(n3265) );
  XOR U3378 ( .A(n3247), .B(n3266), .Z(n3244) );
  NAND U3379 ( .A(A[0]), .B(B[938]), .Z(n3266) );
  NAND U3380 ( .A(B[937]), .B(A[1]), .Z(n3247) );
  NAND U3381 ( .A(n3267), .B(n3268), .Z(n171) );
  NANDN U3382 ( .A(n3269), .B(n3270), .Z(n3268) );
  OR U3383 ( .A(n3271), .B(n3272), .Z(n3270) );
  NAND U3384 ( .A(n3272), .B(n3271), .Z(n3267) );
  XOR U3385 ( .A(n173), .B(n172), .Z(\A1[935] ) );
  XOR U3386 ( .A(n3272), .B(n3273), .Z(n172) );
  XNOR U3387 ( .A(n3271), .B(n3269), .Z(n3273) );
  AND U3388 ( .A(n3274), .B(n3275), .Z(n3269) );
  NANDN U3389 ( .A(n3276), .B(n3277), .Z(n3275) );
  NANDN U3390 ( .A(n3278), .B(n3279), .Z(n3277) );
  AND U3391 ( .A(B[934]), .B(A[3]), .Z(n3271) );
  XNOR U3392 ( .A(n3261), .B(n3280), .Z(n3272) );
  XNOR U3393 ( .A(n3259), .B(n3262), .Z(n3280) );
  NAND U3394 ( .A(A[2]), .B(B[935]), .Z(n3262) );
  NANDN U3395 ( .A(n3281), .B(n3282), .Z(n3259) );
  AND U3396 ( .A(A[0]), .B(B[936]), .Z(n3282) );
  XOR U3397 ( .A(n3264), .B(n3283), .Z(n3261) );
  NAND U3398 ( .A(A[0]), .B(B[937]), .Z(n3283) );
  NAND U3399 ( .A(B[936]), .B(A[1]), .Z(n3264) );
  NAND U3400 ( .A(n3284), .B(n3285), .Z(n173) );
  NANDN U3401 ( .A(n3286), .B(n3287), .Z(n3285) );
  OR U3402 ( .A(n3288), .B(n3289), .Z(n3287) );
  NAND U3403 ( .A(n3289), .B(n3288), .Z(n3284) );
  XOR U3404 ( .A(n175), .B(n174), .Z(\A1[934] ) );
  XOR U3405 ( .A(n3289), .B(n3290), .Z(n174) );
  XNOR U3406 ( .A(n3288), .B(n3286), .Z(n3290) );
  AND U3407 ( .A(n3291), .B(n3292), .Z(n3286) );
  NANDN U3408 ( .A(n3293), .B(n3294), .Z(n3292) );
  NANDN U3409 ( .A(n3295), .B(n3296), .Z(n3294) );
  AND U3410 ( .A(B[933]), .B(A[3]), .Z(n3288) );
  XNOR U3411 ( .A(n3278), .B(n3297), .Z(n3289) );
  XNOR U3412 ( .A(n3276), .B(n3279), .Z(n3297) );
  NAND U3413 ( .A(A[2]), .B(B[934]), .Z(n3279) );
  NANDN U3414 ( .A(n3298), .B(n3299), .Z(n3276) );
  AND U3415 ( .A(A[0]), .B(B[935]), .Z(n3299) );
  XOR U3416 ( .A(n3281), .B(n3300), .Z(n3278) );
  NAND U3417 ( .A(A[0]), .B(B[936]), .Z(n3300) );
  NAND U3418 ( .A(B[935]), .B(A[1]), .Z(n3281) );
  NAND U3419 ( .A(n3301), .B(n3302), .Z(n175) );
  NANDN U3420 ( .A(n3303), .B(n3304), .Z(n3302) );
  OR U3421 ( .A(n3305), .B(n3306), .Z(n3304) );
  NAND U3422 ( .A(n3306), .B(n3305), .Z(n3301) );
  XOR U3423 ( .A(n177), .B(n176), .Z(\A1[933] ) );
  XOR U3424 ( .A(n3306), .B(n3307), .Z(n176) );
  XNOR U3425 ( .A(n3305), .B(n3303), .Z(n3307) );
  AND U3426 ( .A(n3308), .B(n3309), .Z(n3303) );
  NANDN U3427 ( .A(n3310), .B(n3311), .Z(n3309) );
  NANDN U3428 ( .A(n3312), .B(n3313), .Z(n3311) );
  AND U3429 ( .A(B[932]), .B(A[3]), .Z(n3305) );
  XNOR U3430 ( .A(n3295), .B(n3314), .Z(n3306) );
  XNOR U3431 ( .A(n3293), .B(n3296), .Z(n3314) );
  NAND U3432 ( .A(A[2]), .B(B[933]), .Z(n3296) );
  NANDN U3433 ( .A(n3315), .B(n3316), .Z(n3293) );
  AND U3434 ( .A(A[0]), .B(B[934]), .Z(n3316) );
  XOR U3435 ( .A(n3298), .B(n3317), .Z(n3295) );
  NAND U3436 ( .A(A[0]), .B(B[935]), .Z(n3317) );
  NAND U3437 ( .A(B[934]), .B(A[1]), .Z(n3298) );
  NAND U3438 ( .A(n3318), .B(n3319), .Z(n177) );
  NANDN U3439 ( .A(n3320), .B(n3321), .Z(n3319) );
  OR U3440 ( .A(n3322), .B(n3323), .Z(n3321) );
  NAND U3441 ( .A(n3323), .B(n3322), .Z(n3318) );
  XOR U3442 ( .A(n179), .B(n178), .Z(\A1[932] ) );
  XOR U3443 ( .A(n3323), .B(n3324), .Z(n178) );
  XNOR U3444 ( .A(n3322), .B(n3320), .Z(n3324) );
  AND U3445 ( .A(n3325), .B(n3326), .Z(n3320) );
  NANDN U3446 ( .A(n3327), .B(n3328), .Z(n3326) );
  NANDN U3447 ( .A(n3329), .B(n3330), .Z(n3328) );
  AND U3448 ( .A(B[931]), .B(A[3]), .Z(n3322) );
  XNOR U3449 ( .A(n3312), .B(n3331), .Z(n3323) );
  XNOR U3450 ( .A(n3310), .B(n3313), .Z(n3331) );
  NAND U3451 ( .A(A[2]), .B(B[932]), .Z(n3313) );
  NANDN U3452 ( .A(n3332), .B(n3333), .Z(n3310) );
  AND U3453 ( .A(A[0]), .B(B[933]), .Z(n3333) );
  XOR U3454 ( .A(n3315), .B(n3334), .Z(n3312) );
  NAND U3455 ( .A(A[0]), .B(B[934]), .Z(n3334) );
  NAND U3456 ( .A(B[933]), .B(A[1]), .Z(n3315) );
  NAND U3457 ( .A(n3335), .B(n3336), .Z(n179) );
  NANDN U3458 ( .A(n3337), .B(n3338), .Z(n3336) );
  OR U3459 ( .A(n3339), .B(n3340), .Z(n3338) );
  NAND U3460 ( .A(n3340), .B(n3339), .Z(n3335) );
  XOR U3461 ( .A(n181), .B(n180), .Z(\A1[931] ) );
  XOR U3462 ( .A(n3340), .B(n3341), .Z(n180) );
  XNOR U3463 ( .A(n3339), .B(n3337), .Z(n3341) );
  AND U3464 ( .A(n3342), .B(n3343), .Z(n3337) );
  NANDN U3465 ( .A(n3344), .B(n3345), .Z(n3343) );
  NANDN U3466 ( .A(n3346), .B(n3347), .Z(n3345) );
  AND U3467 ( .A(B[930]), .B(A[3]), .Z(n3339) );
  XNOR U3468 ( .A(n3329), .B(n3348), .Z(n3340) );
  XNOR U3469 ( .A(n3327), .B(n3330), .Z(n3348) );
  NAND U3470 ( .A(A[2]), .B(B[931]), .Z(n3330) );
  NANDN U3471 ( .A(n3349), .B(n3350), .Z(n3327) );
  AND U3472 ( .A(A[0]), .B(B[932]), .Z(n3350) );
  XOR U3473 ( .A(n3332), .B(n3351), .Z(n3329) );
  NAND U3474 ( .A(A[0]), .B(B[933]), .Z(n3351) );
  NAND U3475 ( .A(B[932]), .B(A[1]), .Z(n3332) );
  NAND U3476 ( .A(n3352), .B(n3353), .Z(n181) );
  NANDN U3477 ( .A(n3354), .B(n3355), .Z(n3353) );
  OR U3478 ( .A(n3356), .B(n3357), .Z(n3355) );
  NAND U3479 ( .A(n3357), .B(n3356), .Z(n3352) );
  XOR U3480 ( .A(n183), .B(n182), .Z(\A1[930] ) );
  XOR U3481 ( .A(n3357), .B(n3358), .Z(n182) );
  XNOR U3482 ( .A(n3356), .B(n3354), .Z(n3358) );
  AND U3483 ( .A(n3359), .B(n3360), .Z(n3354) );
  NANDN U3484 ( .A(n3361), .B(n3362), .Z(n3360) );
  NANDN U3485 ( .A(n3363), .B(n3364), .Z(n3362) );
  AND U3486 ( .A(B[929]), .B(A[3]), .Z(n3356) );
  XNOR U3487 ( .A(n3346), .B(n3365), .Z(n3357) );
  XNOR U3488 ( .A(n3344), .B(n3347), .Z(n3365) );
  NAND U3489 ( .A(A[2]), .B(B[930]), .Z(n3347) );
  NANDN U3490 ( .A(n3366), .B(n3367), .Z(n3344) );
  AND U3491 ( .A(A[0]), .B(B[931]), .Z(n3367) );
  XOR U3492 ( .A(n3349), .B(n3368), .Z(n3346) );
  NAND U3493 ( .A(A[0]), .B(B[932]), .Z(n3368) );
  NAND U3494 ( .A(B[931]), .B(A[1]), .Z(n3349) );
  NAND U3495 ( .A(n3369), .B(n3370), .Z(n183) );
  NANDN U3496 ( .A(n3371), .B(n3372), .Z(n3370) );
  OR U3497 ( .A(n3373), .B(n3374), .Z(n3372) );
  NAND U3498 ( .A(n3374), .B(n3373), .Z(n3369) );
  XOR U3499 ( .A(n165), .B(n164), .Z(\A1[92] ) );
  XOR U3500 ( .A(n3204), .B(n3375), .Z(n164) );
  XNOR U3501 ( .A(n3203), .B(n3201), .Z(n3375) );
  AND U3502 ( .A(n3376), .B(n3377), .Z(n3201) );
  NANDN U3503 ( .A(n3378), .B(n3379), .Z(n3377) );
  NANDN U3504 ( .A(n3380), .B(n3381), .Z(n3379) );
  AND U3505 ( .A(B[91]), .B(A[3]), .Z(n3203) );
  XNOR U3506 ( .A(n3193), .B(n3382), .Z(n3204) );
  XNOR U3507 ( .A(n3191), .B(n3194), .Z(n3382) );
  NAND U3508 ( .A(A[2]), .B(B[92]), .Z(n3194) );
  NANDN U3509 ( .A(n3383), .B(n3384), .Z(n3191) );
  AND U3510 ( .A(A[0]), .B(B[93]), .Z(n3384) );
  XOR U3511 ( .A(n3196), .B(n3385), .Z(n3193) );
  NAND U3512 ( .A(A[0]), .B(B[94]), .Z(n3385) );
  NAND U3513 ( .A(B[93]), .B(A[1]), .Z(n3196) );
  NAND U3514 ( .A(n3386), .B(n3387), .Z(n165) );
  NANDN U3515 ( .A(n3388), .B(n3389), .Z(n3387) );
  OR U3516 ( .A(n3390), .B(n3391), .Z(n3389) );
  NAND U3517 ( .A(n3391), .B(n3390), .Z(n3386) );
  XOR U3518 ( .A(n185), .B(n184), .Z(\A1[929] ) );
  XOR U3519 ( .A(n3374), .B(n3392), .Z(n184) );
  XNOR U3520 ( .A(n3373), .B(n3371), .Z(n3392) );
  AND U3521 ( .A(n3393), .B(n3394), .Z(n3371) );
  NANDN U3522 ( .A(n3395), .B(n3396), .Z(n3394) );
  NANDN U3523 ( .A(n3397), .B(n3398), .Z(n3396) );
  AND U3524 ( .A(B[928]), .B(A[3]), .Z(n3373) );
  XNOR U3525 ( .A(n3363), .B(n3399), .Z(n3374) );
  XNOR U3526 ( .A(n3361), .B(n3364), .Z(n3399) );
  NAND U3527 ( .A(A[2]), .B(B[929]), .Z(n3364) );
  NANDN U3528 ( .A(n3400), .B(n3401), .Z(n3361) );
  AND U3529 ( .A(A[0]), .B(B[930]), .Z(n3401) );
  XOR U3530 ( .A(n3366), .B(n3402), .Z(n3363) );
  NAND U3531 ( .A(A[0]), .B(B[931]), .Z(n3402) );
  NAND U3532 ( .A(B[930]), .B(A[1]), .Z(n3366) );
  NAND U3533 ( .A(n3403), .B(n3404), .Z(n185) );
  NANDN U3534 ( .A(n3405), .B(n3406), .Z(n3404) );
  OR U3535 ( .A(n3407), .B(n3408), .Z(n3406) );
  NAND U3536 ( .A(n3408), .B(n3407), .Z(n3403) );
  XOR U3537 ( .A(n189), .B(n188), .Z(\A1[928] ) );
  XOR U3538 ( .A(n3408), .B(n3409), .Z(n188) );
  XNOR U3539 ( .A(n3407), .B(n3405), .Z(n3409) );
  AND U3540 ( .A(n3410), .B(n3411), .Z(n3405) );
  NANDN U3541 ( .A(n3412), .B(n3413), .Z(n3411) );
  NANDN U3542 ( .A(n3414), .B(n3415), .Z(n3413) );
  AND U3543 ( .A(B[927]), .B(A[3]), .Z(n3407) );
  XNOR U3544 ( .A(n3397), .B(n3416), .Z(n3408) );
  XNOR U3545 ( .A(n3395), .B(n3398), .Z(n3416) );
  NAND U3546 ( .A(A[2]), .B(B[928]), .Z(n3398) );
  NANDN U3547 ( .A(n3417), .B(n3418), .Z(n3395) );
  AND U3548 ( .A(A[0]), .B(B[929]), .Z(n3418) );
  XOR U3549 ( .A(n3400), .B(n3419), .Z(n3397) );
  NAND U3550 ( .A(A[0]), .B(B[930]), .Z(n3419) );
  NAND U3551 ( .A(B[929]), .B(A[1]), .Z(n3400) );
  NAND U3552 ( .A(n3420), .B(n3421), .Z(n189) );
  NANDN U3553 ( .A(n3422), .B(n3423), .Z(n3421) );
  OR U3554 ( .A(n3424), .B(n3425), .Z(n3423) );
  NAND U3555 ( .A(n3425), .B(n3424), .Z(n3420) );
  XOR U3556 ( .A(n191), .B(n190), .Z(\A1[927] ) );
  XOR U3557 ( .A(n3425), .B(n3426), .Z(n190) );
  XNOR U3558 ( .A(n3424), .B(n3422), .Z(n3426) );
  AND U3559 ( .A(n3427), .B(n3428), .Z(n3422) );
  NANDN U3560 ( .A(n3429), .B(n3430), .Z(n3428) );
  NANDN U3561 ( .A(n3431), .B(n3432), .Z(n3430) );
  AND U3562 ( .A(B[926]), .B(A[3]), .Z(n3424) );
  XNOR U3563 ( .A(n3414), .B(n3433), .Z(n3425) );
  XNOR U3564 ( .A(n3412), .B(n3415), .Z(n3433) );
  NAND U3565 ( .A(A[2]), .B(B[927]), .Z(n3415) );
  NANDN U3566 ( .A(n3434), .B(n3435), .Z(n3412) );
  AND U3567 ( .A(A[0]), .B(B[928]), .Z(n3435) );
  XOR U3568 ( .A(n3417), .B(n3436), .Z(n3414) );
  NAND U3569 ( .A(A[0]), .B(B[929]), .Z(n3436) );
  NAND U3570 ( .A(B[928]), .B(A[1]), .Z(n3417) );
  NAND U3571 ( .A(n3437), .B(n3438), .Z(n191) );
  NANDN U3572 ( .A(n3439), .B(n3440), .Z(n3438) );
  OR U3573 ( .A(n3441), .B(n3442), .Z(n3440) );
  NAND U3574 ( .A(n3442), .B(n3441), .Z(n3437) );
  XOR U3575 ( .A(n193), .B(n192), .Z(\A1[926] ) );
  XOR U3576 ( .A(n3442), .B(n3443), .Z(n192) );
  XNOR U3577 ( .A(n3441), .B(n3439), .Z(n3443) );
  AND U3578 ( .A(n3444), .B(n3445), .Z(n3439) );
  NANDN U3579 ( .A(n3446), .B(n3447), .Z(n3445) );
  NANDN U3580 ( .A(n3448), .B(n3449), .Z(n3447) );
  AND U3581 ( .A(B[925]), .B(A[3]), .Z(n3441) );
  XNOR U3582 ( .A(n3431), .B(n3450), .Z(n3442) );
  XNOR U3583 ( .A(n3429), .B(n3432), .Z(n3450) );
  NAND U3584 ( .A(A[2]), .B(B[926]), .Z(n3432) );
  NANDN U3585 ( .A(n3451), .B(n3452), .Z(n3429) );
  AND U3586 ( .A(A[0]), .B(B[927]), .Z(n3452) );
  XOR U3587 ( .A(n3434), .B(n3453), .Z(n3431) );
  NAND U3588 ( .A(A[0]), .B(B[928]), .Z(n3453) );
  NAND U3589 ( .A(B[927]), .B(A[1]), .Z(n3434) );
  NAND U3590 ( .A(n3454), .B(n3455), .Z(n193) );
  NANDN U3591 ( .A(n3456), .B(n3457), .Z(n3455) );
  OR U3592 ( .A(n3458), .B(n3459), .Z(n3457) );
  NAND U3593 ( .A(n3459), .B(n3458), .Z(n3454) );
  XOR U3594 ( .A(n195), .B(n194), .Z(\A1[925] ) );
  XOR U3595 ( .A(n3459), .B(n3460), .Z(n194) );
  XNOR U3596 ( .A(n3458), .B(n3456), .Z(n3460) );
  AND U3597 ( .A(n3461), .B(n3462), .Z(n3456) );
  NANDN U3598 ( .A(n3463), .B(n3464), .Z(n3462) );
  NANDN U3599 ( .A(n3465), .B(n3466), .Z(n3464) );
  AND U3600 ( .A(B[924]), .B(A[3]), .Z(n3458) );
  XNOR U3601 ( .A(n3448), .B(n3467), .Z(n3459) );
  XNOR U3602 ( .A(n3446), .B(n3449), .Z(n3467) );
  NAND U3603 ( .A(A[2]), .B(B[925]), .Z(n3449) );
  NANDN U3604 ( .A(n3468), .B(n3469), .Z(n3446) );
  AND U3605 ( .A(A[0]), .B(B[926]), .Z(n3469) );
  XOR U3606 ( .A(n3451), .B(n3470), .Z(n3448) );
  NAND U3607 ( .A(A[0]), .B(B[927]), .Z(n3470) );
  NAND U3608 ( .A(B[926]), .B(A[1]), .Z(n3451) );
  NAND U3609 ( .A(n3471), .B(n3472), .Z(n195) );
  NANDN U3610 ( .A(n3473), .B(n3474), .Z(n3472) );
  OR U3611 ( .A(n3475), .B(n3476), .Z(n3474) );
  NAND U3612 ( .A(n3476), .B(n3475), .Z(n3471) );
  XOR U3613 ( .A(n197), .B(n196), .Z(\A1[924] ) );
  XOR U3614 ( .A(n3476), .B(n3477), .Z(n196) );
  XNOR U3615 ( .A(n3475), .B(n3473), .Z(n3477) );
  AND U3616 ( .A(n3478), .B(n3479), .Z(n3473) );
  NANDN U3617 ( .A(n3480), .B(n3481), .Z(n3479) );
  NANDN U3618 ( .A(n3482), .B(n3483), .Z(n3481) );
  AND U3619 ( .A(B[923]), .B(A[3]), .Z(n3475) );
  XNOR U3620 ( .A(n3465), .B(n3484), .Z(n3476) );
  XNOR U3621 ( .A(n3463), .B(n3466), .Z(n3484) );
  NAND U3622 ( .A(A[2]), .B(B[924]), .Z(n3466) );
  NANDN U3623 ( .A(n3485), .B(n3486), .Z(n3463) );
  AND U3624 ( .A(A[0]), .B(B[925]), .Z(n3486) );
  XOR U3625 ( .A(n3468), .B(n3487), .Z(n3465) );
  NAND U3626 ( .A(A[0]), .B(B[926]), .Z(n3487) );
  NAND U3627 ( .A(B[925]), .B(A[1]), .Z(n3468) );
  NAND U3628 ( .A(n3488), .B(n3489), .Z(n197) );
  NANDN U3629 ( .A(n3490), .B(n3491), .Z(n3489) );
  OR U3630 ( .A(n3492), .B(n3493), .Z(n3491) );
  NAND U3631 ( .A(n3493), .B(n3492), .Z(n3488) );
  XOR U3632 ( .A(n199), .B(n198), .Z(\A1[923] ) );
  XOR U3633 ( .A(n3493), .B(n3494), .Z(n198) );
  XNOR U3634 ( .A(n3492), .B(n3490), .Z(n3494) );
  AND U3635 ( .A(n3495), .B(n3496), .Z(n3490) );
  NANDN U3636 ( .A(n3497), .B(n3498), .Z(n3496) );
  NANDN U3637 ( .A(n3499), .B(n3500), .Z(n3498) );
  AND U3638 ( .A(B[922]), .B(A[3]), .Z(n3492) );
  XNOR U3639 ( .A(n3482), .B(n3501), .Z(n3493) );
  XNOR U3640 ( .A(n3480), .B(n3483), .Z(n3501) );
  NAND U3641 ( .A(A[2]), .B(B[923]), .Z(n3483) );
  NANDN U3642 ( .A(n3502), .B(n3503), .Z(n3480) );
  AND U3643 ( .A(A[0]), .B(B[924]), .Z(n3503) );
  XOR U3644 ( .A(n3485), .B(n3504), .Z(n3482) );
  NAND U3645 ( .A(A[0]), .B(B[925]), .Z(n3504) );
  NAND U3646 ( .A(B[924]), .B(A[1]), .Z(n3485) );
  NAND U3647 ( .A(n3505), .B(n3506), .Z(n199) );
  NANDN U3648 ( .A(n3507), .B(n3508), .Z(n3506) );
  OR U3649 ( .A(n3509), .B(n3510), .Z(n3508) );
  NAND U3650 ( .A(n3510), .B(n3509), .Z(n3505) );
  XOR U3651 ( .A(n201), .B(n200), .Z(\A1[922] ) );
  XOR U3652 ( .A(n3510), .B(n3511), .Z(n200) );
  XNOR U3653 ( .A(n3509), .B(n3507), .Z(n3511) );
  AND U3654 ( .A(n3512), .B(n3513), .Z(n3507) );
  NANDN U3655 ( .A(n3514), .B(n3515), .Z(n3513) );
  NANDN U3656 ( .A(n3516), .B(n3517), .Z(n3515) );
  AND U3657 ( .A(B[921]), .B(A[3]), .Z(n3509) );
  XNOR U3658 ( .A(n3499), .B(n3518), .Z(n3510) );
  XNOR U3659 ( .A(n3497), .B(n3500), .Z(n3518) );
  NAND U3660 ( .A(A[2]), .B(B[922]), .Z(n3500) );
  NANDN U3661 ( .A(n3519), .B(n3520), .Z(n3497) );
  AND U3662 ( .A(A[0]), .B(B[923]), .Z(n3520) );
  XOR U3663 ( .A(n3502), .B(n3521), .Z(n3499) );
  NAND U3664 ( .A(A[0]), .B(B[924]), .Z(n3521) );
  NAND U3665 ( .A(B[923]), .B(A[1]), .Z(n3502) );
  NAND U3666 ( .A(n3522), .B(n3523), .Z(n201) );
  NANDN U3667 ( .A(n3524), .B(n3525), .Z(n3523) );
  OR U3668 ( .A(n3526), .B(n3527), .Z(n3525) );
  NAND U3669 ( .A(n3527), .B(n3526), .Z(n3522) );
  XOR U3670 ( .A(n203), .B(n202), .Z(\A1[921] ) );
  XOR U3671 ( .A(n3527), .B(n3528), .Z(n202) );
  XNOR U3672 ( .A(n3526), .B(n3524), .Z(n3528) );
  AND U3673 ( .A(n3529), .B(n3530), .Z(n3524) );
  NANDN U3674 ( .A(n3531), .B(n3532), .Z(n3530) );
  NANDN U3675 ( .A(n3533), .B(n3534), .Z(n3532) );
  AND U3676 ( .A(B[920]), .B(A[3]), .Z(n3526) );
  XNOR U3677 ( .A(n3516), .B(n3535), .Z(n3527) );
  XNOR U3678 ( .A(n3514), .B(n3517), .Z(n3535) );
  NAND U3679 ( .A(A[2]), .B(B[921]), .Z(n3517) );
  NANDN U3680 ( .A(n3536), .B(n3537), .Z(n3514) );
  AND U3681 ( .A(A[0]), .B(B[922]), .Z(n3537) );
  XOR U3682 ( .A(n3519), .B(n3538), .Z(n3516) );
  NAND U3683 ( .A(A[0]), .B(B[923]), .Z(n3538) );
  NAND U3684 ( .A(B[922]), .B(A[1]), .Z(n3519) );
  NAND U3685 ( .A(n3539), .B(n3540), .Z(n203) );
  NANDN U3686 ( .A(n3541), .B(n3542), .Z(n3540) );
  OR U3687 ( .A(n3543), .B(n3544), .Z(n3542) );
  NAND U3688 ( .A(n3544), .B(n3543), .Z(n3539) );
  XOR U3689 ( .A(n205), .B(n204), .Z(\A1[920] ) );
  XOR U3690 ( .A(n3544), .B(n3545), .Z(n204) );
  XNOR U3691 ( .A(n3543), .B(n3541), .Z(n3545) );
  AND U3692 ( .A(n3546), .B(n3547), .Z(n3541) );
  NANDN U3693 ( .A(n3548), .B(n3549), .Z(n3547) );
  NANDN U3694 ( .A(n3550), .B(n3551), .Z(n3549) );
  AND U3695 ( .A(B[919]), .B(A[3]), .Z(n3543) );
  XNOR U3696 ( .A(n3533), .B(n3552), .Z(n3544) );
  XNOR U3697 ( .A(n3531), .B(n3534), .Z(n3552) );
  NAND U3698 ( .A(A[2]), .B(B[920]), .Z(n3534) );
  NANDN U3699 ( .A(n3553), .B(n3554), .Z(n3531) );
  AND U3700 ( .A(A[0]), .B(B[921]), .Z(n3554) );
  XOR U3701 ( .A(n3536), .B(n3555), .Z(n3533) );
  NAND U3702 ( .A(A[0]), .B(B[922]), .Z(n3555) );
  NAND U3703 ( .A(B[921]), .B(A[1]), .Z(n3536) );
  NAND U3704 ( .A(n3556), .B(n3557), .Z(n205) );
  NANDN U3705 ( .A(n3558), .B(n3559), .Z(n3557) );
  OR U3706 ( .A(n3560), .B(n3561), .Z(n3559) );
  NAND U3707 ( .A(n3561), .B(n3560), .Z(n3556) );
  XOR U3708 ( .A(n187), .B(n186), .Z(\A1[91] ) );
  XOR U3709 ( .A(n3391), .B(n3562), .Z(n186) );
  XNOR U3710 ( .A(n3390), .B(n3388), .Z(n3562) );
  AND U3711 ( .A(n3563), .B(n3564), .Z(n3388) );
  NANDN U3712 ( .A(n3565), .B(n3566), .Z(n3564) );
  NANDN U3713 ( .A(n3567), .B(n3568), .Z(n3566) );
  AND U3714 ( .A(B[90]), .B(A[3]), .Z(n3390) );
  XNOR U3715 ( .A(n3380), .B(n3569), .Z(n3391) );
  XNOR U3716 ( .A(n3378), .B(n3381), .Z(n3569) );
  NAND U3717 ( .A(A[2]), .B(B[91]), .Z(n3381) );
  NANDN U3718 ( .A(n3570), .B(n3571), .Z(n3378) );
  AND U3719 ( .A(A[0]), .B(B[92]), .Z(n3571) );
  XOR U3720 ( .A(n3383), .B(n3572), .Z(n3380) );
  NAND U3721 ( .A(A[0]), .B(B[93]), .Z(n3572) );
  NAND U3722 ( .A(B[92]), .B(A[1]), .Z(n3383) );
  NAND U3723 ( .A(n3573), .B(n3574), .Z(n187) );
  NANDN U3724 ( .A(n3575), .B(n3576), .Z(n3574) );
  OR U3725 ( .A(n3577), .B(n3578), .Z(n3576) );
  NAND U3726 ( .A(n3578), .B(n3577), .Z(n3573) );
  XOR U3727 ( .A(n207), .B(n206), .Z(\A1[919] ) );
  XOR U3728 ( .A(n3561), .B(n3579), .Z(n206) );
  XNOR U3729 ( .A(n3560), .B(n3558), .Z(n3579) );
  AND U3730 ( .A(n3580), .B(n3581), .Z(n3558) );
  NANDN U3731 ( .A(n3582), .B(n3583), .Z(n3581) );
  NANDN U3732 ( .A(n3584), .B(n3585), .Z(n3583) );
  AND U3733 ( .A(B[918]), .B(A[3]), .Z(n3560) );
  XNOR U3734 ( .A(n3550), .B(n3586), .Z(n3561) );
  XNOR U3735 ( .A(n3548), .B(n3551), .Z(n3586) );
  NAND U3736 ( .A(A[2]), .B(B[919]), .Z(n3551) );
  NANDN U3737 ( .A(n3587), .B(n3588), .Z(n3548) );
  AND U3738 ( .A(A[0]), .B(B[920]), .Z(n3588) );
  XOR U3739 ( .A(n3553), .B(n3589), .Z(n3550) );
  NAND U3740 ( .A(A[0]), .B(B[921]), .Z(n3589) );
  NAND U3741 ( .A(B[920]), .B(A[1]), .Z(n3553) );
  NAND U3742 ( .A(n3590), .B(n3591), .Z(n207) );
  NANDN U3743 ( .A(n3592), .B(n3593), .Z(n3591) );
  OR U3744 ( .A(n3594), .B(n3595), .Z(n3593) );
  NAND U3745 ( .A(n3595), .B(n3594), .Z(n3590) );
  XOR U3746 ( .A(n211), .B(n210), .Z(\A1[918] ) );
  XOR U3747 ( .A(n3595), .B(n3596), .Z(n210) );
  XNOR U3748 ( .A(n3594), .B(n3592), .Z(n3596) );
  AND U3749 ( .A(n3597), .B(n3598), .Z(n3592) );
  NANDN U3750 ( .A(n3599), .B(n3600), .Z(n3598) );
  NANDN U3751 ( .A(n3601), .B(n3602), .Z(n3600) );
  AND U3752 ( .A(B[917]), .B(A[3]), .Z(n3594) );
  XNOR U3753 ( .A(n3584), .B(n3603), .Z(n3595) );
  XNOR U3754 ( .A(n3582), .B(n3585), .Z(n3603) );
  NAND U3755 ( .A(A[2]), .B(B[918]), .Z(n3585) );
  NANDN U3756 ( .A(n3604), .B(n3605), .Z(n3582) );
  AND U3757 ( .A(A[0]), .B(B[919]), .Z(n3605) );
  XOR U3758 ( .A(n3587), .B(n3606), .Z(n3584) );
  NAND U3759 ( .A(A[0]), .B(B[920]), .Z(n3606) );
  NAND U3760 ( .A(B[919]), .B(A[1]), .Z(n3587) );
  NAND U3761 ( .A(n3607), .B(n3608), .Z(n211) );
  NANDN U3762 ( .A(n3609), .B(n3610), .Z(n3608) );
  OR U3763 ( .A(n3611), .B(n3612), .Z(n3610) );
  NAND U3764 ( .A(n3612), .B(n3611), .Z(n3607) );
  XOR U3765 ( .A(n213), .B(n212), .Z(\A1[917] ) );
  XOR U3766 ( .A(n3612), .B(n3613), .Z(n212) );
  XNOR U3767 ( .A(n3611), .B(n3609), .Z(n3613) );
  AND U3768 ( .A(n3614), .B(n3615), .Z(n3609) );
  NANDN U3769 ( .A(n3616), .B(n3617), .Z(n3615) );
  NANDN U3770 ( .A(n3618), .B(n3619), .Z(n3617) );
  AND U3771 ( .A(B[916]), .B(A[3]), .Z(n3611) );
  XNOR U3772 ( .A(n3601), .B(n3620), .Z(n3612) );
  XNOR U3773 ( .A(n3599), .B(n3602), .Z(n3620) );
  NAND U3774 ( .A(A[2]), .B(B[917]), .Z(n3602) );
  NANDN U3775 ( .A(n3621), .B(n3622), .Z(n3599) );
  AND U3776 ( .A(A[0]), .B(B[918]), .Z(n3622) );
  XOR U3777 ( .A(n3604), .B(n3623), .Z(n3601) );
  NAND U3778 ( .A(A[0]), .B(B[919]), .Z(n3623) );
  NAND U3779 ( .A(B[918]), .B(A[1]), .Z(n3604) );
  NAND U3780 ( .A(n3624), .B(n3625), .Z(n213) );
  NANDN U3781 ( .A(n3626), .B(n3627), .Z(n3625) );
  OR U3782 ( .A(n3628), .B(n3629), .Z(n3627) );
  NAND U3783 ( .A(n3629), .B(n3628), .Z(n3624) );
  XOR U3784 ( .A(n215), .B(n214), .Z(\A1[916] ) );
  XOR U3785 ( .A(n3629), .B(n3630), .Z(n214) );
  XNOR U3786 ( .A(n3628), .B(n3626), .Z(n3630) );
  AND U3787 ( .A(n3631), .B(n3632), .Z(n3626) );
  NANDN U3788 ( .A(n3633), .B(n3634), .Z(n3632) );
  NANDN U3789 ( .A(n3635), .B(n3636), .Z(n3634) );
  AND U3790 ( .A(B[915]), .B(A[3]), .Z(n3628) );
  XNOR U3791 ( .A(n3618), .B(n3637), .Z(n3629) );
  XNOR U3792 ( .A(n3616), .B(n3619), .Z(n3637) );
  NAND U3793 ( .A(A[2]), .B(B[916]), .Z(n3619) );
  NANDN U3794 ( .A(n3638), .B(n3639), .Z(n3616) );
  AND U3795 ( .A(A[0]), .B(B[917]), .Z(n3639) );
  XOR U3796 ( .A(n3621), .B(n3640), .Z(n3618) );
  NAND U3797 ( .A(A[0]), .B(B[918]), .Z(n3640) );
  NAND U3798 ( .A(B[917]), .B(A[1]), .Z(n3621) );
  NAND U3799 ( .A(n3641), .B(n3642), .Z(n215) );
  NANDN U3800 ( .A(n3643), .B(n3644), .Z(n3642) );
  OR U3801 ( .A(n3645), .B(n3646), .Z(n3644) );
  NAND U3802 ( .A(n3646), .B(n3645), .Z(n3641) );
  XOR U3803 ( .A(n217), .B(n216), .Z(\A1[915] ) );
  XOR U3804 ( .A(n3646), .B(n3647), .Z(n216) );
  XNOR U3805 ( .A(n3645), .B(n3643), .Z(n3647) );
  AND U3806 ( .A(n3648), .B(n3649), .Z(n3643) );
  NANDN U3807 ( .A(n3650), .B(n3651), .Z(n3649) );
  NANDN U3808 ( .A(n3652), .B(n3653), .Z(n3651) );
  AND U3809 ( .A(B[914]), .B(A[3]), .Z(n3645) );
  XNOR U3810 ( .A(n3635), .B(n3654), .Z(n3646) );
  XNOR U3811 ( .A(n3633), .B(n3636), .Z(n3654) );
  NAND U3812 ( .A(A[2]), .B(B[915]), .Z(n3636) );
  NANDN U3813 ( .A(n3655), .B(n3656), .Z(n3633) );
  AND U3814 ( .A(A[0]), .B(B[916]), .Z(n3656) );
  XOR U3815 ( .A(n3638), .B(n3657), .Z(n3635) );
  NAND U3816 ( .A(A[0]), .B(B[917]), .Z(n3657) );
  NAND U3817 ( .A(B[916]), .B(A[1]), .Z(n3638) );
  NAND U3818 ( .A(n3658), .B(n3659), .Z(n217) );
  NANDN U3819 ( .A(n3660), .B(n3661), .Z(n3659) );
  OR U3820 ( .A(n3662), .B(n3663), .Z(n3661) );
  NAND U3821 ( .A(n3663), .B(n3662), .Z(n3658) );
  XOR U3822 ( .A(n219), .B(n218), .Z(\A1[914] ) );
  XOR U3823 ( .A(n3663), .B(n3664), .Z(n218) );
  XNOR U3824 ( .A(n3662), .B(n3660), .Z(n3664) );
  AND U3825 ( .A(n3665), .B(n3666), .Z(n3660) );
  NANDN U3826 ( .A(n3667), .B(n3668), .Z(n3666) );
  NANDN U3827 ( .A(n3669), .B(n3670), .Z(n3668) );
  AND U3828 ( .A(B[913]), .B(A[3]), .Z(n3662) );
  XNOR U3829 ( .A(n3652), .B(n3671), .Z(n3663) );
  XNOR U3830 ( .A(n3650), .B(n3653), .Z(n3671) );
  NAND U3831 ( .A(A[2]), .B(B[914]), .Z(n3653) );
  NANDN U3832 ( .A(n3672), .B(n3673), .Z(n3650) );
  AND U3833 ( .A(A[0]), .B(B[915]), .Z(n3673) );
  XOR U3834 ( .A(n3655), .B(n3674), .Z(n3652) );
  NAND U3835 ( .A(A[0]), .B(B[916]), .Z(n3674) );
  NAND U3836 ( .A(B[915]), .B(A[1]), .Z(n3655) );
  NAND U3837 ( .A(n3675), .B(n3676), .Z(n219) );
  NANDN U3838 ( .A(n3677), .B(n3678), .Z(n3676) );
  OR U3839 ( .A(n3679), .B(n3680), .Z(n3678) );
  NAND U3840 ( .A(n3680), .B(n3679), .Z(n3675) );
  XOR U3841 ( .A(n221), .B(n220), .Z(\A1[913] ) );
  XOR U3842 ( .A(n3680), .B(n3681), .Z(n220) );
  XNOR U3843 ( .A(n3679), .B(n3677), .Z(n3681) );
  AND U3844 ( .A(n3682), .B(n3683), .Z(n3677) );
  NANDN U3845 ( .A(n3684), .B(n3685), .Z(n3683) );
  NANDN U3846 ( .A(n3686), .B(n3687), .Z(n3685) );
  AND U3847 ( .A(B[912]), .B(A[3]), .Z(n3679) );
  XNOR U3848 ( .A(n3669), .B(n3688), .Z(n3680) );
  XNOR U3849 ( .A(n3667), .B(n3670), .Z(n3688) );
  NAND U3850 ( .A(A[2]), .B(B[913]), .Z(n3670) );
  NANDN U3851 ( .A(n3689), .B(n3690), .Z(n3667) );
  AND U3852 ( .A(A[0]), .B(B[914]), .Z(n3690) );
  XOR U3853 ( .A(n3672), .B(n3691), .Z(n3669) );
  NAND U3854 ( .A(A[0]), .B(B[915]), .Z(n3691) );
  NAND U3855 ( .A(B[914]), .B(A[1]), .Z(n3672) );
  NAND U3856 ( .A(n3692), .B(n3693), .Z(n221) );
  NANDN U3857 ( .A(n3694), .B(n3695), .Z(n3693) );
  OR U3858 ( .A(n3696), .B(n3697), .Z(n3695) );
  NAND U3859 ( .A(n3697), .B(n3696), .Z(n3692) );
  XOR U3860 ( .A(n223), .B(n222), .Z(\A1[912] ) );
  XOR U3861 ( .A(n3697), .B(n3698), .Z(n222) );
  XNOR U3862 ( .A(n3696), .B(n3694), .Z(n3698) );
  AND U3863 ( .A(n3699), .B(n3700), .Z(n3694) );
  NANDN U3864 ( .A(n3701), .B(n3702), .Z(n3700) );
  NANDN U3865 ( .A(n3703), .B(n3704), .Z(n3702) );
  AND U3866 ( .A(B[911]), .B(A[3]), .Z(n3696) );
  XNOR U3867 ( .A(n3686), .B(n3705), .Z(n3697) );
  XNOR U3868 ( .A(n3684), .B(n3687), .Z(n3705) );
  NAND U3869 ( .A(A[2]), .B(B[912]), .Z(n3687) );
  NANDN U3870 ( .A(n3706), .B(n3707), .Z(n3684) );
  AND U3871 ( .A(A[0]), .B(B[913]), .Z(n3707) );
  XOR U3872 ( .A(n3689), .B(n3708), .Z(n3686) );
  NAND U3873 ( .A(A[0]), .B(B[914]), .Z(n3708) );
  NAND U3874 ( .A(B[913]), .B(A[1]), .Z(n3689) );
  NAND U3875 ( .A(n3709), .B(n3710), .Z(n223) );
  NANDN U3876 ( .A(n3711), .B(n3712), .Z(n3710) );
  OR U3877 ( .A(n3713), .B(n3714), .Z(n3712) );
  NAND U3878 ( .A(n3714), .B(n3713), .Z(n3709) );
  XOR U3879 ( .A(n225), .B(n224), .Z(\A1[911] ) );
  XOR U3880 ( .A(n3714), .B(n3715), .Z(n224) );
  XNOR U3881 ( .A(n3713), .B(n3711), .Z(n3715) );
  AND U3882 ( .A(n3716), .B(n3717), .Z(n3711) );
  NANDN U3883 ( .A(n3718), .B(n3719), .Z(n3717) );
  NANDN U3884 ( .A(n3720), .B(n3721), .Z(n3719) );
  AND U3885 ( .A(B[910]), .B(A[3]), .Z(n3713) );
  XNOR U3886 ( .A(n3703), .B(n3722), .Z(n3714) );
  XNOR U3887 ( .A(n3701), .B(n3704), .Z(n3722) );
  NAND U3888 ( .A(A[2]), .B(B[911]), .Z(n3704) );
  NANDN U3889 ( .A(n3723), .B(n3724), .Z(n3701) );
  AND U3890 ( .A(A[0]), .B(B[912]), .Z(n3724) );
  XOR U3891 ( .A(n3706), .B(n3725), .Z(n3703) );
  NAND U3892 ( .A(A[0]), .B(B[913]), .Z(n3725) );
  NAND U3893 ( .A(B[912]), .B(A[1]), .Z(n3706) );
  NAND U3894 ( .A(n3726), .B(n3727), .Z(n225) );
  NANDN U3895 ( .A(n3728), .B(n3729), .Z(n3727) );
  OR U3896 ( .A(n3730), .B(n3731), .Z(n3729) );
  NAND U3897 ( .A(n3731), .B(n3730), .Z(n3726) );
  XOR U3898 ( .A(n227), .B(n226), .Z(\A1[910] ) );
  XOR U3899 ( .A(n3731), .B(n3732), .Z(n226) );
  XNOR U3900 ( .A(n3730), .B(n3728), .Z(n3732) );
  AND U3901 ( .A(n3733), .B(n3734), .Z(n3728) );
  NANDN U3902 ( .A(n3735), .B(n3736), .Z(n3734) );
  NANDN U3903 ( .A(n3737), .B(n3738), .Z(n3736) );
  AND U3904 ( .A(B[909]), .B(A[3]), .Z(n3730) );
  XNOR U3905 ( .A(n3720), .B(n3739), .Z(n3731) );
  XNOR U3906 ( .A(n3718), .B(n3721), .Z(n3739) );
  NAND U3907 ( .A(A[2]), .B(B[910]), .Z(n3721) );
  NANDN U3908 ( .A(n3740), .B(n3741), .Z(n3718) );
  AND U3909 ( .A(A[0]), .B(B[911]), .Z(n3741) );
  XOR U3910 ( .A(n3723), .B(n3742), .Z(n3720) );
  NAND U3911 ( .A(A[0]), .B(B[912]), .Z(n3742) );
  NAND U3912 ( .A(B[911]), .B(A[1]), .Z(n3723) );
  NAND U3913 ( .A(n3743), .B(n3744), .Z(n227) );
  NANDN U3914 ( .A(n3745), .B(n3746), .Z(n3744) );
  OR U3915 ( .A(n3747), .B(n3748), .Z(n3746) );
  NAND U3916 ( .A(n3748), .B(n3747), .Z(n3743) );
  XOR U3917 ( .A(n209), .B(n208), .Z(\A1[90] ) );
  XOR U3918 ( .A(n3578), .B(n3749), .Z(n208) );
  XNOR U3919 ( .A(n3577), .B(n3575), .Z(n3749) );
  AND U3920 ( .A(n3750), .B(n3751), .Z(n3575) );
  NANDN U3921 ( .A(n3752), .B(n3753), .Z(n3751) );
  NANDN U3922 ( .A(n3754), .B(n3755), .Z(n3753) );
  AND U3923 ( .A(B[89]), .B(A[3]), .Z(n3577) );
  XNOR U3924 ( .A(n3567), .B(n3756), .Z(n3578) );
  XNOR U3925 ( .A(n3565), .B(n3568), .Z(n3756) );
  NAND U3926 ( .A(A[2]), .B(B[90]), .Z(n3568) );
  NANDN U3927 ( .A(n3757), .B(n3758), .Z(n3565) );
  AND U3928 ( .A(A[0]), .B(B[91]), .Z(n3758) );
  XOR U3929 ( .A(n3570), .B(n3759), .Z(n3567) );
  NAND U3930 ( .A(A[0]), .B(B[92]), .Z(n3759) );
  NAND U3931 ( .A(B[91]), .B(A[1]), .Z(n3570) );
  NAND U3932 ( .A(n3760), .B(n3761), .Z(n209) );
  NANDN U3933 ( .A(n3762), .B(n3763), .Z(n3761) );
  OR U3934 ( .A(n3764), .B(n3765), .Z(n3763) );
  NAND U3935 ( .A(n3765), .B(n3764), .Z(n3760) );
  XOR U3936 ( .A(n229), .B(n228), .Z(\A1[909] ) );
  XOR U3937 ( .A(n3748), .B(n3766), .Z(n228) );
  XNOR U3938 ( .A(n3747), .B(n3745), .Z(n3766) );
  AND U3939 ( .A(n3767), .B(n3768), .Z(n3745) );
  NANDN U3940 ( .A(n3769), .B(n3770), .Z(n3768) );
  NANDN U3941 ( .A(n3771), .B(n3772), .Z(n3770) );
  AND U3942 ( .A(B[908]), .B(A[3]), .Z(n3747) );
  XNOR U3943 ( .A(n3737), .B(n3773), .Z(n3748) );
  XNOR U3944 ( .A(n3735), .B(n3738), .Z(n3773) );
  NAND U3945 ( .A(A[2]), .B(B[909]), .Z(n3738) );
  NANDN U3946 ( .A(n3774), .B(n3775), .Z(n3735) );
  AND U3947 ( .A(A[0]), .B(B[910]), .Z(n3775) );
  XOR U3948 ( .A(n3740), .B(n3776), .Z(n3737) );
  NAND U3949 ( .A(A[0]), .B(B[911]), .Z(n3776) );
  NAND U3950 ( .A(B[910]), .B(A[1]), .Z(n3740) );
  NAND U3951 ( .A(n3777), .B(n3778), .Z(n229) );
  NANDN U3952 ( .A(n3779), .B(n3780), .Z(n3778) );
  OR U3953 ( .A(n3781), .B(n3782), .Z(n3780) );
  NAND U3954 ( .A(n3782), .B(n3781), .Z(n3777) );
  XOR U3955 ( .A(n233), .B(n232), .Z(\A1[908] ) );
  XOR U3956 ( .A(n3782), .B(n3783), .Z(n232) );
  XNOR U3957 ( .A(n3781), .B(n3779), .Z(n3783) );
  AND U3958 ( .A(n3784), .B(n3785), .Z(n3779) );
  NANDN U3959 ( .A(n3786), .B(n3787), .Z(n3785) );
  NANDN U3960 ( .A(n3788), .B(n3789), .Z(n3787) );
  AND U3961 ( .A(B[907]), .B(A[3]), .Z(n3781) );
  XNOR U3962 ( .A(n3771), .B(n3790), .Z(n3782) );
  XNOR U3963 ( .A(n3769), .B(n3772), .Z(n3790) );
  NAND U3964 ( .A(A[2]), .B(B[908]), .Z(n3772) );
  NANDN U3965 ( .A(n3791), .B(n3792), .Z(n3769) );
  AND U3966 ( .A(A[0]), .B(B[909]), .Z(n3792) );
  XOR U3967 ( .A(n3774), .B(n3793), .Z(n3771) );
  NAND U3968 ( .A(A[0]), .B(B[910]), .Z(n3793) );
  NAND U3969 ( .A(B[909]), .B(A[1]), .Z(n3774) );
  NAND U3970 ( .A(n3794), .B(n3795), .Z(n233) );
  NANDN U3971 ( .A(n3796), .B(n3797), .Z(n3795) );
  OR U3972 ( .A(n3798), .B(n3799), .Z(n3797) );
  NAND U3973 ( .A(n3799), .B(n3798), .Z(n3794) );
  XOR U3974 ( .A(n235), .B(n234), .Z(\A1[907] ) );
  XOR U3975 ( .A(n3799), .B(n3800), .Z(n234) );
  XNOR U3976 ( .A(n3798), .B(n3796), .Z(n3800) );
  AND U3977 ( .A(n3801), .B(n3802), .Z(n3796) );
  NANDN U3978 ( .A(n3803), .B(n3804), .Z(n3802) );
  NANDN U3979 ( .A(n3805), .B(n3806), .Z(n3804) );
  AND U3980 ( .A(B[906]), .B(A[3]), .Z(n3798) );
  XNOR U3981 ( .A(n3788), .B(n3807), .Z(n3799) );
  XNOR U3982 ( .A(n3786), .B(n3789), .Z(n3807) );
  NAND U3983 ( .A(A[2]), .B(B[907]), .Z(n3789) );
  NANDN U3984 ( .A(n3808), .B(n3809), .Z(n3786) );
  AND U3985 ( .A(A[0]), .B(B[908]), .Z(n3809) );
  XOR U3986 ( .A(n3791), .B(n3810), .Z(n3788) );
  NAND U3987 ( .A(A[0]), .B(B[909]), .Z(n3810) );
  NAND U3988 ( .A(B[908]), .B(A[1]), .Z(n3791) );
  NAND U3989 ( .A(n3811), .B(n3812), .Z(n235) );
  NANDN U3990 ( .A(n3813), .B(n3814), .Z(n3812) );
  OR U3991 ( .A(n3815), .B(n3816), .Z(n3814) );
  NAND U3992 ( .A(n3816), .B(n3815), .Z(n3811) );
  XOR U3993 ( .A(n237), .B(n236), .Z(\A1[906] ) );
  XOR U3994 ( .A(n3816), .B(n3817), .Z(n236) );
  XNOR U3995 ( .A(n3815), .B(n3813), .Z(n3817) );
  AND U3996 ( .A(n3818), .B(n3819), .Z(n3813) );
  NANDN U3997 ( .A(n3820), .B(n3821), .Z(n3819) );
  NANDN U3998 ( .A(n3822), .B(n3823), .Z(n3821) );
  AND U3999 ( .A(B[905]), .B(A[3]), .Z(n3815) );
  XNOR U4000 ( .A(n3805), .B(n3824), .Z(n3816) );
  XNOR U4001 ( .A(n3803), .B(n3806), .Z(n3824) );
  NAND U4002 ( .A(A[2]), .B(B[906]), .Z(n3806) );
  NANDN U4003 ( .A(n3825), .B(n3826), .Z(n3803) );
  AND U4004 ( .A(A[0]), .B(B[907]), .Z(n3826) );
  XOR U4005 ( .A(n3808), .B(n3827), .Z(n3805) );
  NAND U4006 ( .A(A[0]), .B(B[908]), .Z(n3827) );
  NAND U4007 ( .A(B[907]), .B(A[1]), .Z(n3808) );
  NAND U4008 ( .A(n3828), .B(n3829), .Z(n237) );
  NANDN U4009 ( .A(n3830), .B(n3831), .Z(n3829) );
  OR U4010 ( .A(n3832), .B(n3833), .Z(n3831) );
  NAND U4011 ( .A(n3833), .B(n3832), .Z(n3828) );
  XOR U4012 ( .A(n239), .B(n238), .Z(\A1[905] ) );
  XOR U4013 ( .A(n3833), .B(n3834), .Z(n238) );
  XNOR U4014 ( .A(n3832), .B(n3830), .Z(n3834) );
  AND U4015 ( .A(n3835), .B(n3836), .Z(n3830) );
  NANDN U4016 ( .A(n3837), .B(n3838), .Z(n3836) );
  NANDN U4017 ( .A(n3839), .B(n3840), .Z(n3838) );
  AND U4018 ( .A(B[904]), .B(A[3]), .Z(n3832) );
  XNOR U4019 ( .A(n3822), .B(n3841), .Z(n3833) );
  XNOR U4020 ( .A(n3820), .B(n3823), .Z(n3841) );
  NAND U4021 ( .A(A[2]), .B(B[905]), .Z(n3823) );
  NANDN U4022 ( .A(n3842), .B(n3843), .Z(n3820) );
  AND U4023 ( .A(A[0]), .B(B[906]), .Z(n3843) );
  XOR U4024 ( .A(n3825), .B(n3844), .Z(n3822) );
  NAND U4025 ( .A(A[0]), .B(B[907]), .Z(n3844) );
  NAND U4026 ( .A(B[906]), .B(A[1]), .Z(n3825) );
  NAND U4027 ( .A(n3845), .B(n3846), .Z(n239) );
  NANDN U4028 ( .A(n3847), .B(n3848), .Z(n3846) );
  OR U4029 ( .A(n3849), .B(n3850), .Z(n3848) );
  NAND U4030 ( .A(n3850), .B(n3849), .Z(n3845) );
  XOR U4031 ( .A(n241), .B(n240), .Z(\A1[904] ) );
  XOR U4032 ( .A(n3850), .B(n3851), .Z(n240) );
  XNOR U4033 ( .A(n3849), .B(n3847), .Z(n3851) );
  AND U4034 ( .A(n3852), .B(n3853), .Z(n3847) );
  NANDN U4035 ( .A(n3854), .B(n3855), .Z(n3853) );
  NANDN U4036 ( .A(n3856), .B(n3857), .Z(n3855) );
  AND U4037 ( .A(B[903]), .B(A[3]), .Z(n3849) );
  XNOR U4038 ( .A(n3839), .B(n3858), .Z(n3850) );
  XNOR U4039 ( .A(n3837), .B(n3840), .Z(n3858) );
  NAND U4040 ( .A(A[2]), .B(B[904]), .Z(n3840) );
  NANDN U4041 ( .A(n3859), .B(n3860), .Z(n3837) );
  AND U4042 ( .A(A[0]), .B(B[905]), .Z(n3860) );
  XOR U4043 ( .A(n3842), .B(n3861), .Z(n3839) );
  NAND U4044 ( .A(A[0]), .B(B[906]), .Z(n3861) );
  NAND U4045 ( .A(B[905]), .B(A[1]), .Z(n3842) );
  NAND U4046 ( .A(n3862), .B(n3863), .Z(n241) );
  NANDN U4047 ( .A(n3864), .B(n3865), .Z(n3863) );
  OR U4048 ( .A(n3866), .B(n3867), .Z(n3865) );
  NAND U4049 ( .A(n3867), .B(n3866), .Z(n3862) );
  XOR U4050 ( .A(n243), .B(n242), .Z(\A1[903] ) );
  XOR U4051 ( .A(n3867), .B(n3868), .Z(n242) );
  XNOR U4052 ( .A(n3866), .B(n3864), .Z(n3868) );
  AND U4053 ( .A(n3869), .B(n3870), .Z(n3864) );
  NANDN U4054 ( .A(n3871), .B(n3872), .Z(n3870) );
  NANDN U4055 ( .A(n3873), .B(n3874), .Z(n3872) );
  AND U4056 ( .A(B[902]), .B(A[3]), .Z(n3866) );
  XNOR U4057 ( .A(n3856), .B(n3875), .Z(n3867) );
  XNOR U4058 ( .A(n3854), .B(n3857), .Z(n3875) );
  NAND U4059 ( .A(A[2]), .B(B[903]), .Z(n3857) );
  NANDN U4060 ( .A(n3876), .B(n3877), .Z(n3854) );
  AND U4061 ( .A(A[0]), .B(B[904]), .Z(n3877) );
  XOR U4062 ( .A(n3859), .B(n3878), .Z(n3856) );
  NAND U4063 ( .A(A[0]), .B(B[905]), .Z(n3878) );
  NAND U4064 ( .A(B[904]), .B(A[1]), .Z(n3859) );
  NAND U4065 ( .A(n3879), .B(n3880), .Z(n243) );
  NANDN U4066 ( .A(n3881), .B(n3882), .Z(n3880) );
  OR U4067 ( .A(n3883), .B(n3884), .Z(n3882) );
  NAND U4068 ( .A(n3884), .B(n3883), .Z(n3879) );
  XOR U4069 ( .A(n245), .B(n244), .Z(\A1[902] ) );
  XOR U4070 ( .A(n3884), .B(n3885), .Z(n244) );
  XNOR U4071 ( .A(n3883), .B(n3881), .Z(n3885) );
  AND U4072 ( .A(n3886), .B(n3887), .Z(n3881) );
  NANDN U4073 ( .A(n3888), .B(n3889), .Z(n3887) );
  NANDN U4074 ( .A(n3890), .B(n3891), .Z(n3889) );
  AND U4075 ( .A(B[901]), .B(A[3]), .Z(n3883) );
  XNOR U4076 ( .A(n3873), .B(n3892), .Z(n3884) );
  XNOR U4077 ( .A(n3871), .B(n3874), .Z(n3892) );
  NAND U4078 ( .A(A[2]), .B(B[902]), .Z(n3874) );
  NANDN U4079 ( .A(n3893), .B(n3894), .Z(n3871) );
  AND U4080 ( .A(A[0]), .B(B[903]), .Z(n3894) );
  XOR U4081 ( .A(n3876), .B(n3895), .Z(n3873) );
  NAND U4082 ( .A(A[0]), .B(B[904]), .Z(n3895) );
  NAND U4083 ( .A(B[903]), .B(A[1]), .Z(n3876) );
  NAND U4084 ( .A(n3896), .B(n3897), .Z(n245) );
  NANDN U4085 ( .A(n3898), .B(n3899), .Z(n3897) );
  OR U4086 ( .A(n3900), .B(n3901), .Z(n3899) );
  NAND U4087 ( .A(n3901), .B(n3900), .Z(n3896) );
  XOR U4088 ( .A(n247), .B(n246), .Z(\A1[901] ) );
  XOR U4089 ( .A(n3901), .B(n3902), .Z(n246) );
  XNOR U4090 ( .A(n3900), .B(n3898), .Z(n3902) );
  AND U4091 ( .A(n3903), .B(n3904), .Z(n3898) );
  NANDN U4092 ( .A(n3905), .B(n3906), .Z(n3904) );
  NANDN U4093 ( .A(n3907), .B(n3908), .Z(n3906) );
  AND U4094 ( .A(B[900]), .B(A[3]), .Z(n3900) );
  XNOR U4095 ( .A(n3890), .B(n3909), .Z(n3901) );
  XNOR U4096 ( .A(n3888), .B(n3891), .Z(n3909) );
  NAND U4097 ( .A(A[2]), .B(B[901]), .Z(n3891) );
  NANDN U4098 ( .A(n3910), .B(n3911), .Z(n3888) );
  AND U4099 ( .A(A[0]), .B(B[902]), .Z(n3911) );
  XOR U4100 ( .A(n3893), .B(n3912), .Z(n3890) );
  NAND U4101 ( .A(A[0]), .B(B[903]), .Z(n3912) );
  NAND U4102 ( .A(B[902]), .B(A[1]), .Z(n3893) );
  NAND U4103 ( .A(n3913), .B(n3914), .Z(n247) );
  NANDN U4104 ( .A(n3915), .B(n3916), .Z(n3914) );
  OR U4105 ( .A(n3917), .B(n3918), .Z(n3916) );
  NAND U4106 ( .A(n3918), .B(n3917), .Z(n3913) );
  XOR U4107 ( .A(n249), .B(n248), .Z(\A1[900] ) );
  XOR U4108 ( .A(n3918), .B(n3919), .Z(n248) );
  XNOR U4109 ( .A(n3917), .B(n3915), .Z(n3919) );
  AND U4110 ( .A(n3920), .B(n3921), .Z(n3915) );
  NANDN U4111 ( .A(n3922), .B(n3923), .Z(n3921) );
  NANDN U4112 ( .A(n3924), .B(n3925), .Z(n3923) );
  AND U4113 ( .A(B[899]), .B(A[3]), .Z(n3917) );
  XNOR U4114 ( .A(n3907), .B(n3926), .Z(n3918) );
  XNOR U4115 ( .A(n3905), .B(n3908), .Z(n3926) );
  NAND U4116 ( .A(A[2]), .B(B[900]), .Z(n3908) );
  NANDN U4117 ( .A(n3927), .B(n3928), .Z(n3905) );
  AND U4118 ( .A(A[0]), .B(B[901]), .Z(n3928) );
  XOR U4119 ( .A(n3910), .B(n3929), .Z(n3907) );
  NAND U4120 ( .A(A[0]), .B(B[902]), .Z(n3929) );
  NAND U4121 ( .A(B[901]), .B(A[1]), .Z(n3910) );
  NAND U4122 ( .A(n3930), .B(n3931), .Z(n249) );
  NANDN U4123 ( .A(n3932), .B(n3933), .Z(n3931) );
  OR U4124 ( .A(n3934), .B(n3935), .Z(n3933) );
  NAND U4125 ( .A(n3935), .B(n3934), .Z(n3930) );
  XOR U4126 ( .A(n31), .B(n30), .Z(\A1[8] ) );
  XNOR U4127 ( .A(n2080), .B(n3936), .Z(n30) );
  XOR U4128 ( .A(n2082), .B(n2083), .Z(n3936) );
  NAND U4129 ( .A(n3937), .B(n3938), .Z(n2083) );
  NANDN U4130 ( .A(n3939), .B(n3940), .Z(n3938) );
  NANDN U4131 ( .A(n3941), .B(n3942), .Z(n3940) );
  NANDN U4132 ( .A(n3942), .B(n3941), .Z(n3937) );
  AND U4133 ( .A(B[7]), .B(A[3]), .Z(n2082) );
  XOR U4134 ( .A(n20), .B(n3943), .Z(n2080) );
  XOR U4135 ( .A(n3944), .B(n22), .Z(n3943) );
  NAND U4136 ( .A(n3945), .B(n3946), .Z(n31) );
  NANDN U4137 ( .A(n3947), .B(n3948), .Z(n3946) );
  OR U4138 ( .A(n3949), .B(n3950), .Z(n3948) );
  NANDN U4139 ( .A(n23), .B(n3949), .Z(n3945) );
  XOR U4140 ( .A(n231), .B(n230), .Z(\A1[89] ) );
  XOR U4141 ( .A(n3765), .B(n3951), .Z(n230) );
  XNOR U4142 ( .A(n3764), .B(n3762), .Z(n3951) );
  AND U4143 ( .A(n3952), .B(n3953), .Z(n3762) );
  NANDN U4144 ( .A(n3954), .B(n3955), .Z(n3953) );
  NANDN U4145 ( .A(n3956), .B(n3957), .Z(n3955) );
  AND U4146 ( .A(B[88]), .B(A[3]), .Z(n3764) );
  XNOR U4147 ( .A(n3754), .B(n3958), .Z(n3765) );
  XNOR U4148 ( .A(n3752), .B(n3755), .Z(n3958) );
  NAND U4149 ( .A(A[2]), .B(B[89]), .Z(n3755) );
  NANDN U4150 ( .A(n3959), .B(n3960), .Z(n3752) );
  AND U4151 ( .A(A[0]), .B(B[90]), .Z(n3960) );
  XOR U4152 ( .A(n3757), .B(n3961), .Z(n3754) );
  NAND U4153 ( .A(A[0]), .B(B[91]), .Z(n3961) );
  NAND U4154 ( .A(B[90]), .B(A[1]), .Z(n3757) );
  NAND U4155 ( .A(n3962), .B(n3963), .Z(n231) );
  NANDN U4156 ( .A(n3964), .B(n3965), .Z(n3963) );
  OR U4157 ( .A(n3966), .B(n3967), .Z(n3965) );
  NAND U4158 ( .A(n3967), .B(n3966), .Z(n3962) );
  XOR U4159 ( .A(n251), .B(n250), .Z(\A1[899] ) );
  XOR U4160 ( .A(n3935), .B(n3968), .Z(n250) );
  XNOR U4161 ( .A(n3934), .B(n3932), .Z(n3968) );
  AND U4162 ( .A(n3969), .B(n3970), .Z(n3932) );
  NANDN U4163 ( .A(n3971), .B(n3972), .Z(n3970) );
  NANDN U4164 ( .A(n3973), .B(n3974), .Z(n3972) );
  AND U4165 ( .A(B[898]), .B(A[3]), .Z(n3934) );
  XNOR U4166 ( .A(n3924), .B(n3975), .Z(n3935) );
  XNOR U4167 ( .A(n3922), .B(n3925), .Z(n3975) );
  NAND U4168 ( .A(A[2]), .B(B[899]), .Z(n3925) );
  NANDN U4169 ( .A(n3976), .B(n3977), .Z(n3922) );
  AND U4170 ( .A(A[0]), .B(B[900]), .Z(n3977) );
  XOR U4171 ( .A(n3927), .B(n3978), .Z(n3924) );
  NAND U4172 ( .A(A[0]), .B(B[901]), .Z(n3978) );
  NAND U4173 ( .A(B[900]), .B(A[1]), .Z(n3927) );
  NAND U4174 ( .A(n3979), .B(n3980), .Z(n251) );
  NANDN U4175 ( .A(n3981), .B(n3982), .Z(n3980) );
  OR U4176 ( .A(n3983), .B(n3984), .Z(n3982) );
  NAND U4177 ( .A(n3984), .B(n3983), .Z(n3979) );
  XOR U4178 ( .A(n257), .B(n256), .Z(\A1[898] ) );
  XOR U4179 ( .A(n3984), .B(n3985), .Z(n256) );
  XNOR U4180 ( .A(n3983), .B(n3981), .Z(n3985) );
  AND U4181 ( .A(n3986), .B(n3987), .Z(n3981) );
  NANDN U4182 ( .A(n3988), .B(n3989), .Z(n3987) );
  NANDN U4183 ( .A(n3990), .B(n3991), .Z(n3989) );
  AND U4184 ( .A(B[897]), .B(A[3]), .Z(n3983) );
  XNOR U4185 ( .A(n3973), .B(n3992), .Z(n3984) );
  XNOR U4186 ( .A(n3971), .B(n3974), .Z(n3992) );
  NAND U4187 ( .A(A[2]), .B(B[898]), .Z(n3974) );
  NANDN U4188 ( .A(n3993), .B(n3994), .Z(n3971) );
  AND U4189 ( .A(A[0]), .B(B[899]), .Z(n3994) );
  XOR U4190 ( .A(n3976), .B(n3995), .Z(n3973) );
  NAND U4191 ( .A(A[0]), .B(B[900]), .Z(n3995) );
  NAND U4192 ( .A(B[899]), .B(A[1]), .Z(n3976) );
  NAND U4193 ( .A(n3996), .B(n3997), .Z(n257) );
  NANDN U4194 ( .A(n3998), .B(n3999), .Z(n3997) );
  OR U4195 ( .A(n4000), .B(n4001), .Z(n3999) );
  NAND U4196 ( .A(n4001), .B(n4000), .Z(n3996) );
  XOR U4197 ( .A(n259), .B(n258), .Z(\A1[897] ) );
  XOR U4198 ( .A(n4001), .B(n4002), .Z(n258) );
  XNOR U4199 ( .A(n4000), .B(n3998), .Z(n4002) );
  AND U4200 ( .A(n4003), .B(n4004), .Z(n3998) );
  NANDN U4201 ( .A(n4005), .B(n4006), .Z(n4004) );
  NANDN U4202 ( .A(n4007), .B(n4008), .Z(n4006) );
  AND U4203 ( .A(B[896]), .B(A[3]), .Z(n4000) );
  XNOR U4204 ( .A(n3990), .B(n4009), .Z(n4001) );
  XNOR U4205 ( .A(n3988), .B(n3991), .Z(n4009) );
  NAND U4206 ( .A(A[2]), .B(B[897]), .Z(n3991) );
  NANDN U4207 ( .A(n4010), .B(n4011), .Z(n3988) );
  AND U4208 ( .A(A[0]), .B(B[898]), .Z(n4011) );
  XOR U4209 ( .A(n3993), .B(n4012), .Z(n3990) );
  NAND U4210 ( .A(A[0]), .B(B[899]), .Z(n4012) );
  NAND U4211 ( .A(B[898]), .B(A[1]), .Z(n3993) );
  NAND U4212 ( .A(n4013), .B(n4014), .Z(n259) );
  NANDN U4213 ( .A(n4015), .B(n4016), .Z(n4014) );
  OR U4214 ( .A(n4017), .B(n4018), .Z(n4016) );
  NAND U4215 ( .A(n4018), .B(n4017), .Z(n4013) );
  XOR U4216 ( .A(n261), .B(n260), .Z(\A1[896] ) );
  XOR U4217 ( .A(n4018), .B(n4019), .Z(n260) );
  XNOR U4218 ( .A(n4017), .B(n4015), .Z(n4019) );
  AND U4219 ( .A(n4020), .B(n4021), .Z(n4015) );
  NANDN U4220 ( .A(n4022), .B(n4023), .Z(n4021) );
  NANDN U4221 ( .A(n4024), .B(n4025), .Z(n4023) );
  AND U4222 ( .A(B[895]), .B(A[3]), .Z(n4017) );
  XNOR U4223 ( .A(n4007), .B(n4026), .Z(n4018) );
  XNOR U4224 ( .A(n4005), .B(n4008), .Z(n4026) );
  NAND U4225 ( .A(A[2]), .B(B[896]), .Z(n4008) );
  NANDN U4226 ( .A(n4027), .B(n4028), .Z(n4005) );
  AND U4227 ( .A(A[0]), .B(B[897]), .Z(n4028) );
  XOR U4228 ( .A(n4010), .B(n4029), .Z(n4007) );
  NAND U4229 ( .A(A[0]), .B(B[898]), .Z(n4029) );
  NAND U4230 ( .A(B[897]), .B(A[1]), .Z(n4010) );
  NAND U4231 ( .A(n4030), .B(n4031), .Z(n261) );
  NANDN U4232 ( .A(n4032), .B(n4033), .Z(n4031) );
  OR U4233 ( .A(n4034), .B(n4035), .Z(n4033) );
  NAND U4234 ( .A(n4035), .B(n4034), .Z(n4030) );
  XOR U4235 ( .A(n263), .B(n262), .Z(\A1[895] ) );
  XOR U4236 ( .A(n4035), .B(n4036), .Z(n262) );
  XNOR U4237 ( .A(n4034), .B(n4032), .Z(n4036) );
  AND U4238 ( .A(n4037), .B(n4038), .Z(n4032) );
  NANDN U4239 ( .A(n4039), .B(n4040), .Z(n4038) );
  NANDN U4240 ( .A(n4041), .B(n4042), .Z(n4040) );
  AND U4241 ( .A(B[894]), .B(A[3]), .Z(n4034) );
  XNOR U4242 ( .A(n4024), .B(n4043), .Z(n4035) );
  XNOR U4243 ( .A(n4022), .B(n4025), .Z(n4043) );
  NAND U4244 ( .A(A[2]), .B(B[895]), .Z(n4025) );
  NANDN U4245 ( .A(n4044), .B(n4045), .Z(n4022) );
  AND U4246 ( .A(A[0]), .B(B[896]), .Z(n4045) );
  XOR U4247 ( .A(n4027), .B(n4046), .Z(n4024) );
  NAND U4248 ( .A(A[0]), .B(B[897]), .Z(n4046) );
  NAND U4249 ( .A(B[896]), .B(A[1]), .Z(n4027) );
  NAND U4250 ( .A(n4047), .B(n4048), .Z(n263) );
  NANDN U4251 ( .A(n4049), .B(n4050), .Z(n4048) );
  OR U4252 ( .A(n4051), .B(n4052), .Z(n4050) );
  NAND U4253 ( .A(n4052), .B(n4051), .Z(n4047) );
  XOR U4254 ( .A(n265), .B(n264), .Z(\A1[894] ) );
  XOR U4255 ( .A(n4052), .B(n4053), .Z(n264) );
  XNOR U4256 ( .A(n4051), .B(n4049), .Z(n4053) );
  AND U4257 ( .A(n4054), .B(n4055), .Z(n4049) );
  NANDN U4258 ( .A(n4056), .B(n4057), .Z(n4055) );
  NANDN U4259 ( .A(n4058), .B(n4059), .Z(n4057) );
  AND U4260 ( .A(B[893]), .B(A[3]), .Z(n4051) );
  XNOR U4261 ( .A(n4041), .B(n4060), .Z(n4052) );
  XNOR U4262 ( .A(n4039), .B(n4042), .Z(n4060) );
  NAND U4263 ( .A(A[2]), .B(B[894]), .Z(n4042) );
  NANDN U4264 ( .A(n4061), .B(n4062), .Z(n4039) );
  AND U4265 ( .A(A[0]), .B(B[895]), .Z(n4062) );
  XOR U4266 ( .A(n4044), .B(n4063), .Z(n4041) );
  NAND U4267 ( .A(A[0]), .B(B[896]), .Z(n4063) );
  NAND U4268 ( .A(B[895]), .B(A[1]), .Z(n4044) );
  NAND U4269 ( .A(n4064), .B(n4065), .Z(n265) );
  NANDN U4270 ( .A(n4066), .B(n4067), .Z(n4065) );
  OR U4271 ( .A(n4068), .B(n4069), .Z(n4067) );
  NAND U4272 ( .A(n4069), .B(n4068), .Z(n4064) );
  XOR U4273 ( .A(n267), .B(n266), .Z(\A1[893] ) );
  XOR U4274 ( .A(n4069), .B(n4070), .Z(n266) );
  XNOR U4275 ( .A(n4068), .B(n4066), .Z(n4070) );
  AND U4276 ( .A(n4071), .B(n4072), .Z(n4066) );
  NANDN U4277 ( .A(n4073), .B(n4074), .Z(n4072) );
  NANDN U4278 ( .A(n4075), .B(n4076), .Z(n4074) );
  AND U4279 ( .A(B[892]), .B(A[3]), .Z(n4068) );
  XNOR U4280 ( .A(n4058), .B(n4077), .Z(n4069) );
  XNOR U4281 ( .A(n4056), .B(n4059), .Z(n4077) );
  NAND U4282 ( .A(A[2]), .B(B[893]), .Z(n4059) );
  NANDN U4283 ( .A(n4078), .B(n4079), .Z(n4056) );
  AND U4284 ( .A(A[0]), .B(B[894]), .Z(n4079) );
  XOR U4285 ( .A(n4061), .B(n4080), .Z(n4058) );
  NAND U4286 ( .A(A[0]), .B(B[895]), .Z(n4080) );
  NAND U4287 ( .A(B[894]), .B(A[1]), .Z(n4061) );
  NAND U4288 ( .A(n4081), .B(n4082), .Z(n267) );
  NANDN U4289 ( .A(n4083), .B(n4084), .Z(n4082) );
  OR U4290 ( .A(n4085), .B(n4086), .Z(n4084) );
  NAND U4291 ( .A(n4086), .B(n4085), .Z(n4081) );
  XOR U4292 ( .A(n269), .B(n268), .Z(\A1[892] ) );
  XOR U4293 ( .A(n4086), .B(n4087), .Z(n268) );
  XNOR U4294 ( .A(n4085), .B(n4083), .Z(n4087) );
  AND U4295 ( .A(n4088), .B(n4089), .Z(n4083) );
  NANDN U4296 ( .A(n4090), .B(n4091), .Z(n4089) );
  NANDN U4297 ( .A(n4092), .B(n4093), .Z(n4091) );
  AND U4298 ( .A(B[891]), .B(A[3]), .Z(n4085) );
  XNOR U4299 ( .A(n4075), .B(n4094), .Z(n4086) );
  XNOR U4300 ( .A(n4073), .B(n4076), .Z(n4094) );
  NAND U4301 ( .A(A[2]), .B(B[892]), .Z(n4076) );
  NANDN U4302 ( .A(n4095), .B(n4096), .Z(n4073) );
  AND U4303 ( .A(A[0]), .B(B[893]), .Z(n4096) );
  XOR U4304 ( .A(n4078), .B(n4097), .Z(n4075) );
  NAND U4305 ( .A(A[0]), .B(B[894]), .Z(n4097) );
  NAND U4306 ( .A(B[893]), .B(A[1]), .Z(n4078) );
  NAND U4307 ( .A(n4098), .B(n4099), .Z(n269) );
  NANDN U4308 ( .A(n4100), .B(n4101), .Z(n4099) );
  OR U4309 ( .A(n4102), .B(n4103), .Z(n4101) );
  NAND U4310 ( .A(n4103), .B(n4102), .Z(n4098) );
  XOR U4311 ( .A(n271), .B(n270), .Z(\A1[891] ) );
  XOR U4312 ( .A(n4103), .B(n4104), .Z(n270) );
  XNOR U4313 ( .A(n4102), .B(n4100), .Z(n4104) );
  AND U4314 ( .A(n4105), .B(n4106), .Z(n4100) );
  NANDN U4315 ( .A(n4107), .B(n4108), .Z(n4106) );
  NANDN U4316 ( .A(n4109), .B(n4110), .Z(n4108) );
  AND U4317 ( .A(B[890]), .B(A[3]), .Z(n4102) );
  XNOR U4318 ( .A(n4092), .B(n4111), .Z(n4103) );
  XNOR U4319 ( .A(n4090), .B(n4093), .Z(n4111) );
  NAND U4320 ( .A(A[2]), .B(B[891]), .Z(n4093) );
  NANDN U4321 ( .A(n4112), .B(n4113), .Z(n4090) );
  AND U4322 ( .A(A[0]), .B(B[892]), .Z(n4113) );
  XOR U4323 ( .A(n4095), .B(n4114), .Z(n4092) );
  NAND U4324 ( .A(A[0]), .B(B[893]), .Z(n4114) );
  NAND U4325 ( .A(B[892]), .B(A[1]), .Z(n4095) );
  NAND U4326 ( .A(n4115), .B(n4116), .Z(n271) );
  NANDN U4327 ( .A(n4117), .B(n4118), .Z(n4116) );
  OR U4328 ( .A(n4119), .B(n4120), .Z(n4118) );
  NAND U4329 ( .A(n4120), .B(n4119), .Z(n4115) );
  XOR U4330 ( .A(n273), .B(n272), .Z(\A1[890] ) );
  XOR U4331 ( .A(n4120), .B(n4121), .Z(n272) );
  XNOR U4332 ( .A(n4119), .B(n4117), .Z(n4121) );
  AND U4333 ( .A(n4122), .B(n4123), .Z(n4117) );
  NANDN U4334 ( .A(n4124), .B(n4125), .Z(n4123) );
  NANDN U4335 ( .A(n4126), .B(n4127), .Z(n4125) );
  AND U4336 ( .A(B[889]), .B(A[3]), .Z(n4119) );
  XNOR U4337 ( .A(n4109), .B(n4128), .Z(n4120) );
  XNOR U4338 ( .A(n4107), .B(n4110), .Z(n4128) );
  NAND U4339 ( .A(A[2]), .B(B[890]), .Z(n4110) );
  NANDN U4340 ( .A(n4129), .B(n4130), .Z(n4107) );
  AND U4341 ( .A(A[0]), .B(B[891]), .Z(n4130) );
  XOR U4342 ( .A(n4112), .B(n4131), .Z(n4109) );
  NAND U4343 ( .A(A[0]), .B(B[892]), .Z(n4131) );
  NAND U4344 ( .A(B[891]), .B(A[1]), .Z(n4112) );
  NAND U4345 ( .A(n4132), .B(n4133), .Z(n273) );
  NANDN U4346 ( .A(n4134), .B(n4135), .Z(n4133) );
  OR U4347 ( .A(n4136), .B(n4137), .Z(n4135) );
  NAND U4348 ( .A(n4137), .B(n4136), .Z(n4132) );
  XOR U4349 ( .A(n255), .B(n254), .Z(\A1[88] ) );
  XOR U4350 ( .A(n3967), .B(n4138), .Z(n254) );
  XNOR U4351 ( .A(n3966), .B(n3964), .Z(n4138) );
  AND U4352 ( .A(n4139), .B(n4140), .Z(n3964) );
  NANDN U4353 ( .A(n4141), .B(n4142), .Z(n4140) );
  NANDN U4354 ( .A(n4143), .B(n4144), .Z(n4142) );
  AND U4355 ( .A(B[87]), .B(A[3]), .Z(n3966) );
  XNOR U4356 ( .A(n3956), .B(n4145), .Z(n3967) );
  XNOR U4357 ( .A(n3954), .B(n3957), .Z(n4145) );
  NAND U4358 ( .A(A[2]), .B(B[88]), .Z(n3957) );
  NANDN U4359 ( .A(n4146), .B(n4147), .Z(n3954) );
  AND U4360 ( .A(A[0]), .B(B[89]), .Z(n4147) );
  XOR U4361 ( .A(n3959), .B(n4148), .Z(n3956) );
  NAND U4362 ( .A(A[0]), .B(B[90]), .Z(n4148) );
  NAND U4363 ( .A(B[89]), .B(A[1]), .Z(n3959) );
  NAND U4364 ( .A(n4149), .B(n4150), .Z(n255) );
  NANDN U4365 ( .A(n4151), .B(n4152), .Z(n4150) );
  OR U4366 ( .A(n4153), .B(n4154), .Z(n4152) );
  NAND U4367 ( .A(n4154), .B(n4153), .Z(n4149) );
  XOR U4368 ( .A(n275), .B(n274), .Z(\A1[889] ) );
  XOR U4369 ( .A(n4137), .B(n4155), .Z(n274) );
  XNOR U4370 ( .A(n4136), .B(n4134), .Z(n4155) );
  AND U4371 ( .A(n4156), .B(n4157), .Z(n4134) );
  NANDN U4372 ( .A(n4158), .B(n4159), .Z(n4157) );
  NANDN U4373 ( .A(n4160), .B(n4161), .Z(n4159) );
  AND U4374 ( .A(B[888]), .B(A[3]), .Z(n4136) );
  XNOR U4375 ( .A(n4126), .B(n4162), .Z(n4137) );
  XNOR U4376 ( .A(n4124), .B(n4127), .Z(n4162) );
  NAND U4377 ( .A(A[2]), .B(B[889]), .Z(n4127) );
  NANDN U4378 ( .A(n4163), .B(n4164), .Z(n4124) );
  AND U4379 ( .A(A[0]), .B(B[890]), .Z(n4164) );
  XOR U4380 ( .A(n4129), .B(n4165), .Z(n4126) );
  NAND U4381 ( .A(A[0]), .B(B[891]), .Z(n4165) );
  NAND U4382 ( .A(B[890]), .B(A[1]), .Z(n4129) );
  NAND U4383 ( .A(n4166), .B(n4167), .Z(n275) );
  NANDN U4384 ( .A(n4168), .B(n4169), .Z(n4167) );
  OR U4385 ( .A(n4170), .B(n4171), .Z(n4169) );
  NAND U4386 ( .A(n4171), .B(n4170), .Z(n4166) );
  XOR U4387 ( .A(n279), .B(n278), .Z(\A1[888] ) );
  XOR U4388 ( .A(n4171), .B(n4172), .Z(n278) );
  XNOR U4389 ( .A(n4170), .B(n4168), .Z(n4172) );
  AND U4390 ( .A(n4173), .B(n4174), .Z(n4168) );
  NANDN U4391 ( .A(n4175), .B(n4176), .Z(n4174) );
  NANDN U4392 ( .A(n4177), .B(n4178), .Z(n4176) );
  AND U4393 ( .A(B[887]), .B(A[3]), .Z(n4170) );
  XNOR U4394 ( .A(n4160), .B(n4179), .Z(n4171) );
  XNOR U4395 ( .A(n4158), .B(n4161), .Z(n4179) );
  NAND U4396 ( .A(A[2]), .B(B[888]), .Z(n4161) );
  NANDN U4397 ( .A(n4180), .B(n4181), .Z(n4158) );
  AND U4398 ( .A(A[0]), .B(B[889]), .Z(n4181) );
  XOR U4399 ( .A(n4163), .B(n4182), .Z(n4160) );
  NAND U4400 ( .A(A[0]), .B(B[890]), .Z(n4182) );
  NAND U4401 ( .A(B[889]), .B(A[1]), .Z(n4163) );
  NAND U4402 ( .A(n4183), .B(n4184), .Z(n279) );
  NANDN U4403 ( .A(n4185), .B(n4186), .Z(n4184) );
  OR U4404 ( .A(n4187), .B(n4188), .Z(n4186) );
  NAND U4405 ( .A(n4188), .B(n4187), .Z(n4183) );
  XOR U4406 ( .A(n281), .B(n280), .Z(\A1[887] ) );
  XOR U4407 ( .A(n4188), .B(n4189), .Z(n280) );
  XNOR U4408 ( .A(n4187), .B(n4185), .Z(n4189) );
  AND U4409 ( .A(n4190), .B(n4191), .Z(n4185) );
  NANDN U4410 ( .A(n4192), .B(n4193), .Z(n4191) );
  NANDN U4411 ( .A(n4194), .B(n4195), .Z(n4193) );
  AND U4412 ( .A(B[886]), .B(A[3]), .Z(n4187) );
  XNOR U4413 ( .A(n4177), .B(n4196), .Z(n4188) );
  XNOR U4414 ( .A(n4175), .B(n4178), .Z(n4196) );
  NAND U4415 ( .A(A[2]), .B(B[887]), .Z(n4178) );
  NANDN U4416 ( .A(n4197), .B(n4198), .Z(n4175) );
  AND U4417 ( .A(A[0]), .B(B[888]), .Z(n4198) );
  XOR U4418 ( .A(n4180), .B(n4199), .Z(n4177) );
  NAND U4419 ( .A(A[0]), .B(B[889]), .Z(n4199) );
  NAND U4420 ( .A(B[888]), .B(A[1]), .Z(n4180) );
  NAND U4421 ( .A(n4200), .B(n4201), .Z(n281) );
  NANDN U4422 ( .A(n4202), .B(n4203), .Z(n4201) );
  OR U4423 ( .A(n4204), .B(n4205), .Z(n4203) );
  NAND U4424 ( .A(n4205), .B(n4204), .Z(n4200) );
  XOR U4425 ( .A(n283), .B(n282), .Z(\A1[886] ) );
  XOR U4426 ( .A(n4205), .B(n4206), .Z(n282) );
  XNOR U4427 ( .A(n4204), .B(n4202), .Z(n4206) );
  AND U4428 ( .A(n4207), .B(n4208), .Z(n4202) );
  NANDN U4429 ( .A(n4209), .B(n4210), .Z(n4208) );
  NANDN U4430 ( .A(n4211), .B(n4212), .Z(n4210) );
  AND U4431 ( .A(B[885]), .B(A[3]), .Z(n4204) );
  XNOR U4432 ( .A(n4194), .B(n4213), .Z(n4205) );
  XNOR U4433 ( .A(n4192), .B(n4195), .Z(n4213) );
  NAND U4434 ( .A(A[2]), .B(B[886]), .Z(n4195) );
  NANDN U4435 ( .A(n4214), .B(n4215), .Z(n4192) );
  AND U4436 ( .A(A[0]), .B(B[887]), .Z(n4215) );
  XOR U4437 ( .A(n4197), .B(n4216), .Z(n4194) );
  NAND U4438 ( .A(A[0]), .B(B[888]), .Z(n4216) );
  NAND U4439 ( .A(B[887]), .B(A[1]), .Z(n4197) );
  NAND U4440 ( .A(n4217), .B(n4218), .Z(n283) );
  NANDN U4441 ( .A(n4219), .B(n4220), .Z(n4218) );
  OR U4442 ( .A(n4221), .B(n4222), .Z(n4220) );
  NAND U4443 ( .A(n4222), .B(n4221), .Z(n4217) );
  XOR U4444 ( .A(n285), .B(n284), .Z(\A1[885] ) );
  XOR U4445 ( .A(n4222), .B(n4223), .Z(n284) );
  XNOR U4446 ( .A(n4221), .B(n4219), .Z(n4223) );
  AND U4447 ( .A(n4224), .B(n4225), .Z(n4219) );
  NANDN U4448 ( .A(n4226), .B(n4227), .Z(n4225) );
  NANDN U4449 ( .A(n4228), .B(n4229), .Z(n4227) );
  AND U4450 ( .A(B[884]), .B(A[3]), .Z(n4221) );
  XNOR U4451 ( .A(n4211), .B(n4230), .Z(n4222) );
  XNOR U4452 ( .A(n4209), .B(n4212), .Z(n4230) );
  NAND U4453 ( .A(A[2]), .B(B[885]), .Z(n4212) );
  NANDN U4454 ( .A(n4231), .B(n4232), .Z(n4209) );
  AND U4455 ( .A(A[0]), .B(B[886]), .Z(n4232) );
  XOR U4456 ( .A(n4214), .B(n4233), .Z(n4211) );
  NAND U4457 ( .A(A[0]), .B(B[887]), .Z(n4233) );
  NAND U4458 ( .A(B[886]), .B(A[1]), .Z(n4214) );
  NAND U4459 ( .A(n4234), .B(n4235), .Z(n285) );
  NANDN U4460 ( .A(n4236), .B(n4237), .Z(n4235) );
  OR U4461 ( .A(n4238), .B(n4239), .Z(n4237) );
  NAND U4462 ( .A(n4239), .B(n4238), .Z(n4234) );
  XOR U4463 ( .A(n287), .B(n286), .Z(\A1[884] ) );
  XOR U4464 ( .A(n4239), .B(n4240), .Z(n286) );
  XNOR U4465 ( .A(n4238), .B(n4236), .Z(n4240) );
  AND U4466 ( .A(n4241), .B(n4242), .Z(n4236) );
  NANDN U4467 ( .A(n4243), .B(n4244), .Z(n4242) );
  NANDN U4468 ( .A(n4245), .B(n4246), .Z(n4244) );
  AND U4469 ( .A(B[883]), .B(A[3]), .Z(n4238) );
  XNOR U4470 ( .A(n4228), .B(n4247), .Z(n4239) );
  XNOR U4471 ( .A(n4226), .B(n4229), .Z(n4247) );
  NAND U4472 ( .A(A[2]), .B(B[884]), .Z(n4229) );
  NANDN U4473 ( .A(n4248), .B(n4249), .Z(n4226) );
  AND U4474 ( .A(A[0]), .B(B[885]), .Z(n4249) );
  XOR U4475 ( .A(n4231), .B(n4250), .Z(n4228) );
  NAND U4476 ( .A(A[0]), .B(B[886]), .Z(n4250) );
  NAND U4477 ( .A(B[885]), .B(A[1]), .Z(n4231) );
  NAND U4478 ( .A(n4251), .B(n4252), .Z(n287) );
  NANDN U4479 ( .A(n4253), .B(n4254), .Z(n4252) );
  OR U4480 ( .A(n4255), .B(n4256), .Z(n4254) );
  NAND U4481 ( .A(n4256), .B(n4255), .Z(n4251) );
  XOR U4482 ( .A(n289), .B(n288), .Z(\A1[883] ) );
  XOR U4483 ( .A(n4256), .B(n4257), .Z(n288) );
  XNOR U4484 ( .A(n4255), .B(n4253), .Z(n4257) );
  AND U4485 ( .A(n4258), .B(n4259), .Z(n4253) );
  NANDN U4486 ( .A(n4260), .B(n4261), .Z(n4259) );
  NANDN U4487 ( .A(n4262), .B(n4263), .Z(n4261) );
  AND U4488 ( .A(B[882]), .B(A[3]), .Z(n4255) );
  XNOR U4489 ( .A(n4245), .B(n4264), .Z(n4256) );
  XNOR U4490 ( .A(n4243), .B(n4246), .Z(n4264) );
  NAND U4491 ( .A(A[2]), .B(B[883]), .Z(n4246) );
  NANDN U4492 ( .A(n4265), .B(n4266), .Z(n4243) );
  AND U4493 ( .A(A[0]), .B(B[884]), .Z(n4266) );
  XOR U4494 ( .A(n4248), .B(n4267), .Z(n4245) );
  NAND U4495 ( .A(A[0]), .B(B[885]), .Z(n4267) );
  NAND U4496 ( .A(B[884]), .B(A[1]), .Z(n4248) );
  NAND U4497 ( .A(n4268), .B(n4269), .Z(n289) );
  NANDN U4498 ( .A(n4270), .B(n4271), .Z(n4269) );
  OR U4499 ( .A(n4272), .B(n4273), .Z(n4271) );
  NAND U4500 ( .A(n4273), .B(n4272), .Z(n4268) );
  XOR U4501 ( .A(n291), .B(n290), .Z(\A1[882] ) );
  XOR U4502 ( .A(n4273), .B(n4274), .Z(n290) );
  XNOR U4503 ( .A(n4272), .B(n4270), .Z(n4274) );
  AND U4504 ( .A(n4275), .B(n4276), .Z(n4270) );
  NANDN U4505 ( .A(n4277), .B(n4278), .Z(n4276) );
  NANDN U4506 ( .A(n4279), .B(n4280), .Z(n4278) );
  AND U4507 ( .A(B[881]), .B(A[3]), .Z(n4272) );
  XNOR U4508 ( .A(n4262), .B(n4281), .Z(n4273) );
  XNOR U4509 ( .A(n4260), .B(n4263), .Z(n4281) );
  NAND U4510 ( .A(A[2]), .B(B[882]), .Z(n4263) );
  NANDN U4511 ( .A(n4282), .B(n4283), .Z(n4260) );
  AND U4512 ( .A(A[0]), .B(B[883]), .Z(n4283) );
  XOR U4513 ( .A(n4265), .B(n4284), .Z(n4262) );
  NAND U4514 ( .A(A[0]), .B(B[884]), .Z(n4284) );
  NAND U4515 ( .A(B[883]), .B(A[1]), .Z(n4265) );
  NAND U4516 ( .A(n4285), .B(n4286), .Z(n291) );
  NANDN U4517 ( .A(n4287), .B(n4288), .Z(n4286) );
  OR U4518 ( .A(n4289), .B(n4290), .Z(n4288) );
  NAND U4519 ( .A(n4290), .B(n4289), .Z(n4285) );
  XOR U4520 ( .A(n293), .B(n292), .Z(\A1[881] ) );
  XOR U4521 ( .A(n4290), .B(n4291), .Z(n292) );
  XNOR U4522 ( .A(n4289), .B(n4287), .Z(n4291) );
  AND U4523 ( .A(n4292), .B(n4293), .Z(n4287) );
  NANDN U4524 ( .A(n4294), .B(n4295), .Z(n4293) );
  NANDN U4525 ( .A(n4296), .B(n4297), .Z(n4295) );
  AND U4526 ( .A(B[880]), .B(A[3]), .Z(n4289) );
  XNOR U4527 ( .A(n4279), .B(n4298), .Z(n4290) );
  XNOR U4528 ( .A(n4277), .B(n4280), .Z(n4298) );
  NAND U4529 ( .A(A[2]), .B(B[881]), .Z(n4280) );
  NANDN U4530 ( .A(n4299), .B(n4300), .Z(n4277) );
  AND U4531 ( .A(A[0]), .B(B[882]), .Z(n4300) );
  XOR U4532 ( .A(n4282), .B(n4301), .Z(n4279) );
  NAND U4533 ( .A(A[0]), .B(B[883]), .Z(n4301) );
  NAND U4534 ( .A(B[882]), .B(A[1]), .Z(n4282) );
  NAND U4535 ( .A(n4302), .B(n4303), .Z(n293) );
  NANDN U4536 ( .A(n4304), .B(n4305), .Z(n4303) );
  OR U4537 ( .A(n4306), .B(n4307), .Z(n4305) );
  NAND U4538 ( .A(n4307), .B(n4306), .Z(n4302) );
  XOR U4539 ( .A(n295), .B(n294), .Z(\A1[880] ) );
  XOR U4540 ( .A(n4307), .B(n4308), .Z(n294) );
  XNOR U4541 ( .A(n4306), .B(n4304), .Z(n4308) );
  AND U4542 ( .A(n4309), .B(n4310), .Z(n4304) );
  NANDN U4543 ( .A(n4311), .B(n4312), .Z(n4310) );
  NANDN U4544 ( .A(n4313), .B(n4314), .Z(n4312) );
  AND U4545 ( .A(B[879]), .B(A[3]), .Z(n4306) );
  XNOR U4546 ( .A(n4296), .B(n4315), .Z(n4307) );
  XNOR U4547 ( .A(n4294), .B(n4297), .Z(n4315) );
  NAND U4548 ( .A(A[2]), .B(B[880]), .Z(n4297) );
  NANDN U4549 ( .A(n4316), .B(n4317), .Z(n4294) );
  AND U4550 ( .A(A[0]), .B(B[881]), .Z(n4317) );
  XOR U4551 ( .A(n4299), .B(n4318), .Z(n4296) );
  NAND U4552 ( .A(A[0]), .B(B[882]), .Z(n4318) );
  NAND U4553 ( .A(B[881]), .B(A[1]), .Z(n4299) );
  NAND U4554 ( .A(n4319), .B(n4320), .Z(n295) );
  NANDN U4555 ( .A(n4321), .B(n4322), .Z(n4320) );
  OR U4556 ( .A(n4323), .B(n4324), .Z(n4322) );
  NAND U4557 ( .A(n4324), .B(n4323), .Z(n4319) );
  XOR U4558 ( .A(n277), .B(n276), .Z(\A1[87] ) );
  XOR U4559 ( .A(n4154), .B(n4325), .Z(n276) );
  XNOR U4560 ( .A(n4153), .B(n4151), .Z(n4325) );
  AND U4561 ( .A(n4326), .B(n4327), .Z(n4151) );
  NANDN U4562 ( .A(n4328), .B(n4329), .Z(n4327) );
  NANDN U4563 ( .A(n4330), .B(n4331), .Z(n4329) );
  AND U4564 ( .A(B[86]), .B(A[3]), .Z(n4153) );
  XNOR U4565 ( .A(n4143), .B(n4332), .Z(n4154) );
  XNOR U4566 ( .A(n4141), .B(n4144), .Z(n4332) );
  NAND U4567 ( .A(A[2]), .B(B[87]), .Z(n4144) );
  NANDN U4568 ( .A(n4333), .B(n4334), .Z(n4141) );
  AND U4569 ( .A(A[0]), .B(B[88]), .Z(n4334) );
  XOR U4570 ( .A(n4146), .B(n4335), .Z(n4143) );
  NAND U4571 ( .A(A[0]), .B(B[89]), .Z(n4335) );
  NAND U4572 ( .A(B[88]), .B(A[1]), .Z(n4146) );
  NAND U4573 ( .A(n4336), .B(n4337), .Z(n277) );
  NANDN U4574 ( .A(n4338), .B(n4339), .Z(n4337) );
  OR U4575 ( .A(n4340), .B(n4341), .Z(n4339) );
  NAND U4576 ( .A(n4341), .B(n4340), .Z(n4336) );
  XOR U4577 ( .A(n297), .B(n296), .Z(\A1[879] ) );
  XOR U4578 ( .A(n4324), .B(n4342), .Z(n296) );
  XNOR U4579 ( .A(n4323), .B(n4321), .Z(n4342) );
  AND U4580 ( .A(n4343), .B(n4344), .Z(n4321) );
  NANDN U4581 ( .A(n4345), .B(n4346), .Z(n4344) );
  NANDN U4582 ( .A(n4347), .B(n4348), .Z(n4346) );
  AND U4583 ( .A(B[878]), .B(A[3]), .Z(n4323) );
  XNOR U4584 ( .A(n4313), .B(n4349), .Z(n4324) );
  XNOR U4585 ( .A(n4311), .B(n4314), .Z(n4349) );
  NAND U4586 ( .A(A[2]), .B(B[879]), .Z(n4314) );
  NANDN U4587 ( .A(n4350), .B(n4351), .Z(n4311) );
  AND U4588 ( .A(A[0]), .B(B[880]), .Z(n4351) );
  XOR U4589 ( .A(n4316), .B(n4352), .Z(n4313) );
  NAND U4590 ( .A(A[0]), .B(B[881]), .Z(n4352) );
  NAND U4591 ( .A(B[880]), .B(A[1]), .Z(n4316) );
  NAND U4592 ( .A(n4353), .B(n4354), .Z(n297) );
  NANDN U4593 ( .A(n4355), .B(n4356), .Z(n4354) );
  OR U4594 ( .A(n4357), .B(n4358), .Z(n4356) );
  NAND U4595 ( .A(n4358), .B(n4357), .Z(n4353) );
  XOR U4596 ( .A(n301), .B(n300), .Z(\A1[878] ) );
  XOR U4597 ( .A(n4358), .B(n4359), .Z(n300) );
  XNOR U4598 ( .A(n4357), .B(n4355), .Z(n4359) );
  AND U4599 ( .A(n4360), .B(n4361), .Z(n4355) );
  NANDN U4600 ( .A(n4362), .B(n4363), .Z(n4361) );
  NANDN U4601 ( .A(n4364), .B(n4365), .Z(n4363) );
  AND U4602 ( .A(B[877]), .B(A[3]), .Z(n4357) );
  XNOR U4603 ( .A(n4347), .B(n4366), .Z(n4358) );
  XNOR U4604 ( .A(n4345), .B(n4348), .Z(n4366) );
  NAND U4605 ( .A(A[2]), .B(B[878]), .Z(n4348) );
  NANDN U4606 ( .A(n4367), .B(n4368), .Z(n4345) );
  AND U4607 ( .A(A[0]), .B(B[879]), .Z(n4368) );
  XOR U4608 ( .A(n4350), .B(n4369), .Z(n4347) );
  NAND U4609 ( .A(A[0]), .B(B[880]), .Z(n4369) );
  NAND U4610 ( .A(B[879]), .B(A[1]), .Z(n4350) );
  NAND U4611 ( .A(n4370), .B(n4371), .Z(n301) );
  NANDN U4612 ( .A(n4372), .B(n4373), .Z(n4371) );
  OR U4613 ( .A(n4374), .B(n4375), .Z(n4373) );
  NAND U4614 ( .A(n4375), .B(n4374), .Z(n4370) );
  XOR U4615 ( .A(n303), .B(n302), .Z(\A1[877] ) );
  XOR U4616 ( .A(n4375), .B(n4376), .Z(n302) );
  XNOR U4617 ( .A(n4374), .B(n4372), .Z(n4376) );
  AND U4618 ( .A(n4377), .B(n4378), .Z(n4372) );
  NANDN U4619 ( .A(n4379), .B(n4380), .Z(n4378) );
  NANDN U4620 ( .A(n4381), .B(n4382), .Z(n4380) );
  AND U4621 ( .A(B[876]), .B(A[3]), .Z(n4374) );
  XNOR U4622 ( .A(n4364), .B(n4383), .Z(n4375) );
  XNOR U4623 ( .A(n4362), .B(n4365), .Z(n4383) );
  NAND U4624 ( .A(A[2]), .B(B[877]), .Z(n4365) );
  NANDN U4625 ( .A(n4384), .B(n4385), .Z(n4362) );
  AND U4626 ( .A(A[0]), .B(B[878]), .Z(n4385) );
  XOR U4627 ( .A(n4367), .B(n4386), .Z(n4364) );
  NAND U4628 ( .A(A[0]), .B(B[879]), .Z(n4386) );
  NAND U4629 ( .A(B[878]), .B(A[1]), .Z(n4367) );
  NAND U4630 ( .A(n4387), .B(n4388), .Z(n303) );
  NANDN U4631 ( .A(n4389), .B(n4390), .Z(n4388) );
  OR U4632 ( .A(n4391), .B(n4392), .Z(n4390) );
  NAND U4633 ( .A(n4392), .B(n4391), .Z(n4387) );
  XOR U4634 ( .A(n305), .B(n304), .Z(\A1[876] ) );
  XOR U4635 ( .A(n4392), .B(n4393), .Z(n304) );
  XNOR U4636 ( .A(n4391), .B(n4389), .Z(n4393) );
  AND U4637 ( .A(n4394), .B(n4395), .Z(n4389) );
  NANDN U4638 ( .A(n4396), .B(n4397), .Z(n4395) );
  NANDN U4639 ( .A(n4398), .B(n4399), .Z(n4397) );
  AND U4640 ( .A(B[875]), .B(A[3]), .Z(n4391) );
  XNOR U4641 ( .A(n4381), .B(n4400), .Z(n4392) );
  XNOR U4642 ( .A(n4379), .B(n4382), .Z(n4400) );
  NAND U4643 ( .A(A[2]), .B(B[876]), .Z(n4382) );
  NANDN U4644 ( .A(n4401), .B(n4402), .Z(n4379) );
  AND U4645 ( .A(A[0]), .B(B[877]), .Z(n4402) );
  XOR U4646 ( .A(n4384), .B(n4403), .Z(n4381) );
  NAND U4647 ( .A(A[0]), .B(B[878]), .Z(n4403) );
  NAND U4648 ( .A(B[877]), .B(A[1]), .Z(n4384) );
  NAND U4649 ( .A(n4404), .B(n4405), .Z(n305) );
  NANDN U4650 ( .A(n4406), .B(n4407), .Z(n4405) );
  OR U4651 ( .A(n4408), .B(n4409), .Z(n4407) );
  NAND U4652 ( .A(n4409), .B(n4408), .Z(n4404) );
  XOR U4653 ( .A(n307), .B(n306), .Z(\A1[875] ) );
  XOR U4654 ( .A(n4409), .B(n4410), .Z(n306) );
  XNOR U4655 ( .A(n4408), .B(n4406), .Z(n4410) );
  AND U4656 ( .A(n4411), .B(n4412), .Z(n4406) );
  NANDN U4657 ( .A(n4413), .B(n4414), .Z(n4412) );
  NANDN U4658 ( .A(n4415), .B(n4416), .Z(n4414) );
  AND U4659 ( .A(B[874]), .B(A[3]), .Z(n4408) );
  XNOR U4660 ( .A(n4398), .B(n4417), .Z(n4409) );
  XNOR U4661 ( .A(n4396), .B(n4399), .Z(n4417) );
  NAND U4662 ( .A(A[2]), .B(B[875]), .Z(n4399) );
  NANDN U4663 ( .A(n4418), .B(n4419), .Z(n4396) );
  AND U4664 ( .A(A[0]), .B(B[876]), .Z(n4419) );
  XOR U4665 ( .A(n4401), .B(n4420), .Z(n4398) );
  NAND U4666 ( .A(A[0]), .B(B[877]), .Z(n4420) );
  NAND U4667 ( .A(B[876]), .B(A[1]), .Z(n4401) );
  NAND U4668 ( .A(n4421), .B(n4422), .Z(n307) );
  NANDN U4669 ( .A(n4423), .B(n4424), .Z(n4422) );
  OR U4670 ( .A(n4425), .B(n4426), .Z(n4424) );
  NAND U4671 ( .A(n4426), .B(n4425), .Z(n4421) );
  XOR U4672 ( .A(n309), .B(n308), .Z(\A1[874] ) );
  XOR U4673 ( .A(n4426), .B(n4427), .Z(n308) );
  XNOR U4674 ( .A(n4425), .B(n4423), .Z(n4427) );
  AND U4675 ( .A(n4428), .B(n4429), .Z(n4423) );
  NANDN U4676 ( .A(n4430), .B(n4431), .Z(n4429) );
  NANDN U4677 ( .A(n4432), .B(n4433), .Z(n4431) );
  AND U4678 ( .A(B[873]), .B(A[3]), .Z(n4425) );
  XNOR U4679 ( .A(n4415), .B(n4434), .Z(n4426) );
  XNOR U4680 ( .A(n4413), .B(n4416), .Z(n4434) );
  NAND U4681 ( .A(A[2]), .B(B[874]), .Z(n4416) );
  NANDN U4682 ( .A(n4435), .B(n4436), .Z(n4413) );
  AND U4683 ( .A(A[0]), .B(B[875]), .Z(n4436) );
  XOR U4684 ( .A(n4418), .B(n4437), .Z(n4415) );
  NAND U4685 ( .A(A[0]), .B(B[876]), .Z(n4437) );
  NAND U4686 ( .A(B[875]), .B(A[1]), .Z(n4418) );
  NAND U4687 ( .A(n4438), .B(n4439), .Z(n309) );
  NANDN U4688 ( .A(n4440), .B(n4441), .Z(n4439) );
  OR U4689 ( .A(n4442), .B(n4443), .Z(n4441) );
  NAND U4690 ( .A(n4443), .B(n4442), .Z(n4438) );
  XOR U4691 ( .A(n311), .B(n310), .Z(\A1[873] ) );
  XOR U4692 ( .A(n4443), .B(n4444), .Z(n310) );
  XNOR U4693 ( .A(n4442), .B(n4440), .Z(n4444) );
  AND U4694 ( .A(n4445), .B(n4446), .Z(n4440) );
  NANDN U4695 ( .A(n4447), .B(n4448), .Z(n4446) );
  NANDN U4696 ( .A(n4449), .B(n4450), .Z(n4448) );
  AND U4697 ( .A(B[872]), .B(A[3]), .Z(n4442) );
  XNOR U4698 ( .A(n4432), .B(n4451), .Z(n4443) );
  XNOR U4699 ( .A(n4430), .B(n4433), .Z(n4451) );
  NAND U4700 ( .A(A[2]), .B(B[873]), .Z(n4433) );
  NANDN U4701 ( .A(n4452), .B(n4453), .Z(n4430) );
  AND U4702 ( .A(A[0]), .B(B[874]), .Z(n4453) );
  XOR U4703 ( .A(n4435), .B(n4454), .Z(n4432) );
  NAND U4704 ( .A(A[0]), .B(B[875]), .Z(n4454) );
  NAND U4705 ( .A(B[874]), .B(A[1]), .Z(n4435) );
  NAND U4706 ( .A(n4455), .B(n4456), .Z(n311) );
  NANDN U4707 ( .A(n4457), .B(n4458), .Z(n4456) );
  OR U4708 ( .A(n4459), .B(n4460), .Z(n4458) );
  NAND U4709 ( .A(n4460), .B(n4459), .Z(n4455) );
  XOR U4710 ( .A(n313), .B(n312), .Z(\A1[872] ) );
  XOR U4711 ( .A(n4460), .B(n4461), .Z(n312) );
  XNOR U4712 ( .A(n4459), .B(n4457), .Z(n4461) );
  AND U4713 ( .A(n4462), .B(n4463), .Z(n4457) );
  NANDN U4714 ( .A(n4464), .B(n4465), .Z(n4463) );
  NANDN U4715 ( .A(n4466), .B(n4467), .Z(n4465) );
  AND U4716 ( .A(B[871]), .B(A[3]), .Z(n4459) );
  XNOR U4717 ( .A(n4449), .B(n4468), .Z(n4460) );
  XNOR U4718 ( .A(n4447), .B(n4450), .Z(n4468) );
  NAND U4719 ( .A(A[2]), .B(B[872]), .Z(n4450) );
  NANDN U4720 ( .A(n4469), .B(n4470), .Z(n4447) );
  AND U4721 ( .A(A[0]), .B(B[873]), .Z(n4470) );
  XOR U4722 ( .A(n4452), .B(n4471), .Z(n4449) );
  NAND U4723 ( .A(A[0]), .B(B[874]), .Z(n4471) );
  NAND U4724 ( .A(B[873]), .B(A[1]), .Z(n4452) );
  NAND U4725 ( .A(n4472), .B(n4473), .Z(n313) );
  NANDN U4726 ( .A(n4474), .B(n4475), .Z(n4473) );
  OR U4727 ( .A(n4476), .B(n4477), .Z(n4475) );
  NAND U4728 ( .A(n4477), .B(n4476), .Z(n4472) );
  XOR U4729 ( .A(n315), .B(n314), .Z(\A1[871] ) );
  XOR U4730 ( .A(n4477), .B(n4478), .Z(n314) );
  XNOR U4731 ( .A(n4476), .B(n4474), .Z(n4478) );
  AND U4732 ( .A(n4479), .B(n4480), .Z(n4474) );
  NANDN U4733 ( .A(n4481), .B(n4482), .Z(n4480) );
  NANDN U4734 ( .A(n4483), .B(n4484), .Z(n4482) );
  AND U4735 ( .A(B[870]), .B(A[3]), .Z(n4476) );
  XNOR U4736 ( .A(n4466), .B(n4485), .Z(n4477) );
  XNOR U4737 ( .A(n4464), .B(n4467), .Z(n4485) );
  NAND U4738 ( .A(A[2]), .B(B[871]), .Z(n4467) );
  NANDN U4739 ( .A(n4486), .B(n4487), .Z(n4464) );
  AND U4740 ( .A(A[0]), .B(B[872]), .Z(n4487) );
  XOR U4741 ( .A(n4469), .B(n4488), .Z(n4466) );
  NAND U4742 ( .A(A[0]), .B(B[873]), .Z(n4488) );
  NAND U4743 ( .A(B[872]), .B(A[1]), .Z(n4469) );
  NAND U4744 ( .A(n4489), .B(n4490), .Z(n315) );
  NANDN U4745 ( .A(n4491), .B(n4492), .Z(n4490) );
  OR U4746 ( .A(n4493), .B(n4494), .Z(n4492) );
  NAND U4747 ( .A(n4494), .B(n4493), .Z(n4489) );
  XOR U4748 ( .A(n317), .B(n316), .Z(\A1[870] ) );
  XOR U4749 ( .A(n4494), .B(n4495), .Z(n316) );
  XNOR U4750 ( .A(n4493), .B(n4491), .Z(n4495) );
  AND U4751 ( .A(n4496), .B(n4497), .Z(n4491) );
  NANDN U4752 ( .A(n4498), .B(n4499), .Z(n4497) );
  NANDN U4753 ( .A(n4500), .B(n4501), .Z(n4499) );
  AND U4754 ( .A(B[869]), .B(A[3]), .Z(n4493) );
  XNOR U4755 ( .A(n4483), .B(n4502), .Z(n4494) );
  XNOR U4756 ( .A(n4481), .B(n4484), .Z(n4502) );
  NAND U4757 ( .A(A[2]), .B(B[870]), .Z(n4484) );
  NANDN U4758 ( .A(n4503), .B(n4504), .Z(n4481) );
  AND U4759 ( .A(A[0]), .B(B[871]), .Z(n4504) );
  XOR U4760 ( .A(n4486), .B(n4505), .Z(n4483) );
  NAND U4761 ( .A(A[0]), .B(B[872]), .Z(n4505) );
  NAND U4762 ( .A(B[871]), .B(A[1]), .Z(n4486) );
  NAND U4763 ( .A(n4506), .B(n4507), .Z(n317) );
  NANDN U4764 ( .A(n4508), .B(n4509), .Z(n4507) );
  OR U4765 ( .A(n4510), .B(n4511), .Z(n4509) );
  NAND U4766 ( .A(n4511), .B(n4510), .Z(n4506) );
  XOR U4767 ( .A(n299), .B(n298), .Z(\A1[86] ) );
  XOR U4768 ( .A(n4341), .B(n4512), .Z(n298) );
  XNOR U4769 ( .A(n4340), .B(n4338), .Z(n4512) );
  AND U4770 ( .A(n4513), .B(n4514), .Z(n4338) );
  NANDN U4771 ( .A(n4515), .B(n4516), .Z(n4514) );
  NANDN U4772 ( .A(n4517), .B(n4518), .Z(n4516) );
  AND U4773 ( .A(B[85]), .B(A[3]), .Z(n4340) );
  XNOR U4774 ( .A(n4330), .B(n4519), .Z(n4341) );
  XNOR U4775 ( .A(n4328), .B(n4331), .Z(n4519) );
  NAND U4776 ( .A(A[2]), .B(B[86]), .Z(n4331) );
  NANDN U4777 ( .A(n4520), .B(n4521), .Z(n4328) );
  AND U4778 ( .A(A[0]), .B(B[87]), .Z(n4521) );
  XOR U4779 ( .A(n4333), .B(n4522), .Z(n4330) );
  NAND U4780 ( .A(A[0]), .B(B[88]), .Z(n4522) );
  NAND U4781 ( .A(B[87]), .B(A[1]), .Z(n4333) );
  NAND U4782 ( .A(n4523), .B(n4524), .Z(n299) );
  NANDN U4783 ( .A(n4525), .B(n4526), .Z(n4524) );
  OR U4784 ( .A(n4527), .B(n4528), .Z(n4526) );
  NAND U4785 ( .A(n4528), .B(n4527), .Z(n4523) );
  XOR U4786 ( .A(n319), .B(n318), .Z(\A1[869] ) );
  XOR U4787 ( .A(n4511), .B(n4529), .Z(n318) );
  XNOR U4788 ( .A(n4510), .B(n4508), .Z(n4529) );
  AND U4789 ( .A(n4530), .B(n4531), .Z(n4508) );
  NANDN U4790 ( .A(n4532), .B(n4533), .Z(n4531) );
  NANDN U4791 ( .A(n4534), .B(n4535), .Z(n4533) );
  AND U4792 ( .A(B[868]), .B(A[3]), .Z(n4510) );
  XNOR U4793 ( .A(n4500), .B(n4536), .Z(n4511) );
  XNOR U4794 ( .A(n4498), .B(n4501), .Z(n4536) );
  NAND U4795 ( .A(A[2]), .B(B[869]), .Z(n4501) );
  NANDN U4796 ( .A(n4537), .B(n4538), .Z(n4498) );
  AND U4797 ( .A(A[0]), .B(B[870]), .Z(n4538) );
  XOR U4798 ( .A(n4503), .B(n4539), .Z(n4500) );
  NAND U4799 ( .A(A[0]), .B(B[871]), .Z(n4539) );
  NAND U4800 ( .A(B[870]), .B(A[1]), .Z(n4503) );
  NAND U4801 ( .A(n4540), .B(n4541), .Z(n319) );
  NANDN U4802 ( .A(n4542), .B(n4543), .Z(n4541) );
  OR U4803 ( .A(n4544), .B(n4545), .Z(n4543) );
  NAND U4804 ( .A(n4545), .B(n4544), .Z(n4540) );
  XOR U4805 ( .A(n323), .B(n322), .Z(\A1[868] ) );
  XOR U4806 ( .A(n4545), .B(n4546), .Z(n322) );
  XNOR U4807 ( .A(n4544), .B(n4542), .Z(n4546) );
  AND U4808 ( .A(n4547), .B(n4548), .Z(n4542) );
  NANDN U4809 ( .A(n4549), .B(n4550), .Z(n4548) );
  NANDN U4810 ( .A(n4551), .B(n4552), .Z(n4550) );
  AND U4811 ( .A(B[867]), .B(A[3]), .Z(n4544) );
  XNOR U4812 ( .A(n4534), .B(n4553), .Z(n4545) );
  XNOR U4813 ( .A(n4532), .B(n4535), .Z(n4553) );
  NAND U4814 ( .A(A[2]), .B(B[868]), .Z(n4535) );
  NANDN U4815 ( .A(n4554), .B(n4555), .Z(n4532) );
  AND U4816 ( .A(A[0]), .B(B[869]), .Z(n4555) );
  XOR U4817 ( .A(n4537), .B(n4556), .Z(n4534) );
  NAND U4818 ( .A(A[0]), .B(B[870]), .Z(n4556) );
  NAND U4819 ( .A(B[869]), .B(A[1]), .Z(n4537) );
  NAND U4820 ( .A(n4557), .B(n4558), .Z(n323) );
  NANDN U4821 ( .A(n4559), .B(n4560), .Z(n4558) );
  OR U4822 ( .A(n4561), .B(n4562), .Z(n4560) );
  NAND U4823 ( .A(n4562), .B(n4561), .Z(n4557) );
  XOR U4824 ( .A(n325), .B(n324), .Z(\A1[867] ) );
  XOR U4825 ( .A(n4562), .B(n4563), .Z(n324) );
  XNOR U4826 ( .A(n4561), .B(n4559), .Z(n4563) );
  AND U4827 ( .A(n4564), .B(n4565), .Z(n4559) );
  NANDN U4828 ( .A(n4566), .B(n4567), .Z(n4565) );
  NANDN U4829 ( .A(n4568), .B(n4569), .Z(n4567) );
  AND U4830 ( .A(B[866]), .B(A[3]), .Z(n4561) );
  XNOR U4831 ( .A(n4551), .B(n4570), .Z(n4562) );
  XNOR U4832 ( .A(n4549), .B(n4552), .Z(n4570) );
  NAND U4833 ( .A(A[2]), .B(B[867]), .Z(n4552) );
  NANDN U4834 ( .A(n4571), .B(n4572), .Z(n4549) );
  AND U4835 ( .A(A[0]), .B(B[868]), .Z(n4572) );
  XOR U4836 ( .A(n4554), .B(n4573), .Z(n4551) );
  NAND U4837 ( .A(A[0]), .B(B[869]), .Z(n4573) );
  NAND U4838 ( .A(B[868]), .B(A[1]), .Z(n4554) );
  NAND U4839 ( .A(n4574), .B(n4575), .Z(n325) );
  NANDN U4840 ( .A(n4576), .B(n4577), .Z(n4575) );
  OR U4841 ( .A(n4578), .B(n4579), .Z(n4577) );
  NAND U4842 ( .A(n4579), .B(n4578), .Z(n4574) );
  XOR U4843 ( .A(n327), .B(n326), .Z(\A1[866] ) );
  XOR U4844 ( .A(n4579), .B(n4580), .Z(n326) );
  XNOR U4845 ( .A(n4578), .B(n4576), .Z(n4580) );
  AND U4846 ( .A(n4581), .B(n4582), .Z(n4576) );
  NANDN U4847 ( .A(n4583), .B(n4584), .Z(n4582) );
  NANDN U4848 ( .A(n4585), .B(n4586), .Z(n4584) );
  AND U4849 ( .A(B[865]), .B(A[3]), .Z(n4578) );
  XNOR U4850 ( .A(n4568), .B(n4587), .Z(n4579) );
  XNOR U4851 ( .A(n4566), .B(n4569), .Z(n4587) );
  NAND U4852 ( .A(A[2]), .B(B[866]), .Z(n4569) );
  NANDN U4853 ( .A(n4588), .B(n4589), .Z(n4566) );
  AND U4854 ( .A(A[0]), .B(B[867]), .Z(n4589) );
  XOR U4855 ( .A(n4571), .B(n4590), .Z(n4568) );
  NAND U4856 ( .A(A[0]), .B(B[868]), .Z(n4590) );
  NAND U4857 ( .A(B[867]), .B(A[1]), .Z(n4571) );
  NAND U4858 ( .A(n4591), .B(n4592), .Z(n327) );
  NANDN U4859 ( .A(n4593), .B(n4594), .Z(n4592) );
  OR U4860 ( .A(n4595), .B(n4596), .Z(n4594) );
  NAND U4861 ( .A(n4596), .B(n4595), .Z(n4591) );
  XOR U4862 ( .A(n329), .B(n328), .Z(\A1[865] ) );
  XOR U4863 ( .A(n4596), .B(n4597), .Z(n328) );
  XNOR U4864 ( .A(n4595), .B(n4593), .Z(n4597) );
  AND U4865 ( .A(n4598), .B(n4599), .Z(n4593) );
  NANDN U4866 ( .A(n4600), .B(n4601), .Z(n4599) );
  NANDN U4867 ( .A(n4602), .B(n4603), .Z(n4601) );
  AND U4868 ( .A(B[864]), .B(A[3]), .Z(n4595) );
  XNOR U4869 ( .A(n4585), .B(n4604), .Z(n4596) );
  XNOR U4870 ( .A(n4583), .B(n4586), .Z(n4604) );
  NAND U4871 ( .A(A[2]), .B(B[865]), .Z(n4586) );
  NANDN U4872 ( .A(n4605), .B(n4606), .Z(n4583) );
  AND U4873 ( .A(A[0]), .B(B[866]), .Z(n4606) );
  XOR U4874 ( .A(n4588), .B(n4607), .Z(n4585) );
  NAND U4875 ( .A(A[0]), .B(B[867]), .Z(n4607) );
  NAND U4876 ( .A(B[866]), .B(A[1]), .Z(n4588) );
  NAND U4877 ( .A(n4608), .B(n4609), .Z(n329) );
  NANDN U4878 ( .A(n4610), .B(n4611), .Z(n4609) );
  OR U4879 ( .A(n4612), .B(n4613), .Z(n4611) );
  NAND U4880 ( .A(n4613), .B(n4612), .Z(n4608) );
  XOR U4881 ( .A(n331), .B(n330), .Z(\A1[864] ) );
  XOR U4882 ( .A(n4613), .B(n4614), .Z(n330) );
  XNOR U4883 ( .A(n4612), .B(n4610), .Z(n4614) );
  AND U4884 ( .A(n4615), .B(n4616), .Z(n4610) );
  NANDN U4885 ( .A(n4617), .B(n4618), .Z(n4616) );
  NANDN U4886 ( .A(n4619), .B(n4620), .Z(n4618) );
  AND U4887 ( .A(B[863]), .B(A[3]), .Z(n4612) );
  XNOR U4888 ( .A(n4602), .B(n4621), .Z(n4613) );
  XNOR U4889 ( .A(n4600), .B(n4603), .Z(n4621) );
  NAND U4890 ( .A(A[2]), .B(B[864]), .Z(n4603) );
  NANDN U4891 ( .A(n4622), .B(n4623), .Z(n4600) );
  AND U4892 ( .A(A[0]), .B(B[865]), .Z(n4623) );
  XOR U4893 ( .A(n4605), .B(n4624), .Z(n4602) );
  NAND U4894 ( .A(A[0]), .B(B[866]), .Z(n4624) );
  NAND U4895 ( .A(B[865]), .B(A[1]), .Z(n4605) );
  NAND U4896 ( .A(n4625), .B(n4626), .Z(n331) );
  NANDN U4897 ( .A(n4627), .B(n4628), .Z(n4626) );
  OR U4898 ( .A(n4629), .B(n4630), .Z(n4628) );
  NAND U4899 ( .A(n4630), .B(n4629), .Z(n4625) );
  XOR U4900 ( .A(n333), .B(n332), .Z(\A1[863] ) );
  XOR U4901 ( .A(n4630), .B(n4631), .Z(n332) );
  XNOR U4902 ( .A(n4629), .B(n4627), .Z(n4631) );
  AND U4903 ( .A(n4632), .B(n4633), .Z(n4627) );
  NANDN U4904 ( .A(n4634), .B(n4635), .Z(n4633) );
  NANDN U4905 ( .A(n4636), .B(n4637), .Z(n4635) );
  AND U4906 ( .A(B[862]), .B(A[3]), .Z(n4629) );
  XNOR U4907 ( .A(n4619), .B(n4638), .Z(n4630) );
  XNOR U4908 ( .A(n4617), .B(n4620), .Z(n4638) );
  NAND U4909 ( .A(A[2]), .B(B[863]), .Z(n4620) );
  NANDN U4910 ( .A(n4639), .B(n4640), .Z(n4617) );
  AND U4911 ( .A(A[0]), .B(B[864]), .Z(n4640) );
  XOR U4912 ( .A(n4622), .B(n4641), .Z(n4619) );
  NAND U4913 ( .A(A[0]), .B(B[865]), .Z(n4641) );
  NAND U4914 ( .A(B[864]), .B(A[1]), .Z(n4622) );
  NAND U4915 ( .A(n4642), .B(n4643), .Z(n333) );
  NANDN U4916 ( .A(n4644), .B(n4645), .Z(n4643) );
  OR U4917 ( .A(n4646), .B(n4647), .Z(n4645) );
  NAND U4918 ( .A(n4647), .B(n4646), .Z(n4642) );
  XOR U4919 ( .A(n335), .B(n334), .Z(\A1[862] ) );
  XOR U4920 ( .A(n4647), .B(n4648), .Z(n334) );
  XNOR U4921 ( .A(n4646), .B(n4644), .Z(n4648) );
  AND U4922 ( .A(n4649), .B(n4650), .Z(n4644) );
  NANDN U4923 ( .A(n4651), .B(n4652), .Z(n4650) );
  NANDN U4924 ( .A(n4653), .B(n4654), .Z(n4652) );
  AND U4925 ( .A(B[861]), .B(A[3]), .Z(n4646) );
  XNOR U4926 ( .A(n4636), .B(n4655), .Z(n4647) );
  XNOR U4927 ( .A(n4634), .B(n4637), .Z(n4655) );
  NAND U4928 ( .A(A[2]), .B(B[862]), .Z(n4637) );
  NANDN U4929 ( .A(n4656), .B(n4657), .Z(n4634) );
  AND U4930 ( .A(A[0]), .B(B[863]), .Z(n4657) );
  XOR U4931 ( .A(n4639), .B(n4658), .Z(n4636) );
  NAND U4932 ( .A(A[0]), .B(B[864]), .Z(n4658) );
  NAND U4933 ( .A(B[863]), .B(A[1]), .Z(n4639) );
  NAND U4934 ( .A(n4659), .B(n4660), .Z(n335) );
  NANDN U4935 ( .A(n4661), .B(n4662), .Z(n4660) );
  OR U4936 ( .A(n4663), .B(n4664), .Z(n4662) );
  NAND U4937 ( .A(n4664), .B(n4663), .Z(n4659) );
  XOR U4938 ( .A(n337), .B(n336), .Z(\A1[861] ) );
  XOR U4939 ( .A(n4664), .B(n4665), .Z(n336) );
  XNOR U4940 ( .A(n4663), .B(n4661), .Z(n4665) );
  AND U4941 ( .A(n4666), .B(n4667), .Z(n4661) );
  NANDN U4942 ( .A(n4668), .B(n4669), .Z(n4667) );
  NANDN U4943 ( .A(n4670), .B(n4671), .Z(n4669) );
  AND U4944 ( .A(B[860]), .B(A[3]), .Z(n4663) );
  XNOR U4945 ( .A(n4653), .B(n4672), .Z(n4664) );
  XNOR U4946 ( .A(n4651), .B(n4654), .Z(n4672) );
  NAND U4947 ( .A(A[2]), .B(B[861]), .Z(n4654) );
  NANDN U4948 ( .A(n4673), .B(n4674), .Z(n4651) );
  AND U4949 ( .A(A[0]), .B(B[862]), .Z(n4674) );
  XOR U4950 ( .A(n4656), .B(n4675), .Z(n4653) );
  NAND U4951 ( .A(A[0]), .B(B[863]), .Z(n4675) );
  NAND U4952 ( .A(B[862]), .B(A[1]), .Z(n4656) );
  NAND U4953 ( .A(n4676), .B(n4677), .Z(n337) );
  NANDN U4954 ( .A(n4678), .B(n4679), .Z(n4677) );
  OR U4955 ( .A(n4680), .B(n4681), .Z(n4679) );
  NAND U4956 ( .A(n4681), .B(n4680), .Z(n4676) );
  XOR U4957 ( .A(n339), .B(n338), .Z(\A1[860] ) );
  XOR U4958 ( .A(n4681), .B(n4682), .Z(n338) );
  XNOR U4959 ( .A(n4680), .B(n4678), .Z(n4682) );
  AND U4960 ( .A(n4683), .B(n4684), .Z(n4678) );
  NANDN U4961 ( .A(n4685), .B(n4686), .Z(n4684) );
  NANDN U4962 ( .A(n4687), .B(n4688), .Z(n4686) );
  AND U4963 ( .A(B[859]), .B(A[3]), .Z(n4680) );
  XNOR U4964 ( .A(n4670), .B(n4689), .Z(n4681) );
  XNOR U4965 ( .A(n4668), .B(n4671), .Z(n4689) );
  NAND U4966 ( .A(A[2]), .B(B[860]), .Z(n4671) );
  NANDN U4967 ( .A(n4690), .B(n4691), .Z(n4668) );
  AND U4968 ( .A(A[0]), .B(B[861]), .Z(n4691) );
  XOR U4969 ( .A(n4673), .B(n4692), .Z(n4670) );
  NAND U4970 ( .A(A[0]), .B(B[862]), .Z(n4692) );
  NAND U4971 ( .A(B[861]), .B(A[1]), .Z(n4673) );
  NAND U4972 ( .A(n4693), .B(n4694), .Z(n339) );
  NANDN U4973 ( .A(n4695), .B(n4696), .Z(n4694) );
  OR U4974 ( .A(n4697), .B(n4698), .Z(n4696) );
  NAND U4975 ( .A(n4698), .B(n4697), .Z(n4693) );
  XOR U4976 ( .A(n321), .B(n320), .Z(\A1[85] ) );
  XOR U4977 ( .A(n4528), .B(n4699), .Z(n320) );
  XNOR U4978 ( .A(n4527), .B(n4525), .Z(n4699) );
  AND U4979 ( .A(n4700), .B(n4701), .Z(n4525) );
  NANDN U4980 ( .A(n4702), .B(n4703), .Z(n4701) );
  NANDN U4981 ( .A(n4704), .B(n4705), .Z(n4703) );
  AND U4982 ( .A(B[84]), .B(A[3]), .Z(n4527) );
  XNOR U4983 ( .A(n4517), .B(n4706), .Z(n4528) );
  XNOR U4984 ( .A(n4515), .B(n4518), .Z(n4706) );
  NAND U4985 ( .A(A[2]), .B(B[85]), .Z(n4518) );
  NANDN U4986 ( .A(n4707), .B(n4708), .Z(n4515) );
  AND U4987 ( .A(A[0]), .B(B[86]), .Z(n4708) );
  XOR U4988 ( .A(n4520), .B(n4709), .Z(n4517) );
  NAND U4989 ( .A(A[0]), .B(B[87]), .Z(n4709) );
  NAND U4990 ( .A(B[86]), .B(A[1]), .Z(n4520) );
  NAND U4991 ( .A(n4710), .B(n4711), .Z(n321) );
  NANDN U4992 ( .A(n4712), .B(n4713), .Z(n4711) );
  OR U4993 ( .A(n4714), .B(n4715), .Z(n4713) );
  NAND U4994 ( .A(n4715), .B(n4714), .Z(n4710) );
  XOR U4995 ( .A(n341), .B(n340), .Z(\A1[859] ) );
  XOR U4996 ( .A(n4698), .B(n4716), .Z(n340) );
  XNOR U4997 ( .A(n4697), .B(n4695), .Z(n4716) );
  AND U4998 ( .A(n4717), .B(n4718), .Z(n4695) );
  NANDN U4999 ( .A(n4719), .B(n4720), .Z(n4718) );
  NANDN U5000 ( .A(n4721), .B(n4722), .Z(n4720) );
  AND U5001 ( .A(B[858]), .B(A[3]), .Z(n4697) );
  XNOR U5002 ( .A(n4687), .B(n4723), .Z(n4698) );
  XNOR U5003 ( .A(n4685), .B(n4688), .Z(n4723) );
  NAND U5004 ( .A(A[2]), .B(B[859]), .Z(n4688) );
  NANDN U5005 ( .A(n4724), .B(n4725), .Z(n4685) );
  AND U5006 ( .A(A[0]), .B(B[860]), .Z(n4725) );
  XOR U5007 ( .A(n4690), .B(n4726), .Z(n4687) );
  NAND U5008 ( .A(A[0]), .B(B[861]), .Z(n4726) );
  NAND U5009 ( .A(B[860]), .B(A[1]), .Z(n4690) );
  NAND U5010 ( .A(n4727), .B(n4728), .Z(n341) );
  NANDN U5011 ( .A(n4729), .B(n4730), .Z(n4728) );
  OR U5012 ( .A(n4731), .B(n4732), .Z(n4730) );
  NAND U5013 ( .A(n4732), .B(n4731), .Z(n4727) );
  XOR U5014 ( .A(n345), .B(n344), .Z(\A1[858] ) );
  XOR U5015 ( .A(n4732), .B(n4733), .Z(n344) );
  XNOR U5016 ( .A(n4731), .B(n4729), .Z(n4733) );
  AND U5017 ( .A(n4734), .B(n4735), .Z(n4729) );
  NANDN U5018 ( .A(n4736), .B(n4737), .Z(n4735) );
  NANDN U5019 ( .A(n4738), .B(n4739), .Z(n4737) );
  AND U5020 ( .A(B[857]), .B(A[3]), .Z(n4731) );
  XNOR U5021 ( .A(n4721), .B(n4740), .Z(n4732) );
  XNOR U5022 ( .A(n4719), .B(n4722), .Z(n4740) );
  NAND U5023 ( .A(A[2]), .B(B[858]), .Z(n4722) );
  NANDN U5024 ( .A(n4741), .B(n4742), .Z(n4719) );
  AND U5025 ( .A(A[0]), .B(B[859]), .Z(n4742) );
  XOR U5026 ( .A(n4724), .B(n4743), .Z(n4721) );
  NAND U5027 ( .A(A[0]), .B(B[860]), .Z(n4743) );
  NAND U5028 ( .A(B[859]), .B(A[1]), .Z(n4724) );
  NAND U5029 ( .A(n4744), .B(n4745), .Z(n345) );
  NANDN U5030 ( .A(n4746), .B(n4747), .Z(n4745) );
  OR U5031 ( .A(n4748), .B(n4749), .Z(n4747) );
  NAND U5032 ( .A(n4749), .B(n4748), .Z(n4744) );
  XOR U5033 ( .A(n347), .B(n346), .Z(\A1[857] ) );
  XOR U5034 ( .A(n4749), .B(n4750), .Z(n346) );
  XNOR U5035 ( .A(n4748), .B(n4746), .Z(n4750) );
  AND U5036 ( .A(n4751), .B(n4752), .Z(n4746) );
  NANDN U5037 ( .A(n4753), .B(n4754), .Z(n4752) );
  NANDN U5038 ( .A(n4755), .B(n4756), .Z(n4754) );
  AND U5039 ( .A(B[856]), .B(A[3]), .Z(n4748) );
  XNOR U5040 ( .A(n4738), .B(n4757), .Z(n4749) );
  XNOR U5041 ( .A(n4736), .B(n4739), .Z(n4757) );
  NAND U5042 ( .A(A[2]), .B(B[857]), .Z(n4739) );
  NANDN U5043 ( .A(n4758), .B(n4759), .Z(n4736) );
  AND U5044 ( .A(A[0]), .B(B[858]), .Z(n4759) );
  XOR U5045 ( .A(n4741), .B(n4760), .Z(n4738) );
  NAND U5046 ( .A(A[0]), .B(B[859]), .Z(n4760) );
  NAND U5047 ( .A(B[858]), .B(A[1]), .Z(n4741) );
  NAND U5048 ( .A(n4761), .B(n4762), .Z(n347) );
  NANDN U5049 ( .A(n4763), .B(n4764), .Z(n4762) );
  OR U5050 ( .A(n4765), .B(n4766), .Z(n4764) );
  NAND U5051 ( .A(n4766), .B(n4765), .Z(n4761) );
  XOR U5052 ( .A(n349), .B(n348), .Z(\A1[856] ) );
  XOR U5053 ( .A(n4766), .B(n4767), .Z(n348) );
  XNOR U5054 ( .A(n4765), .B(n4763), .Z(n4767) );
  AND U5055 ( .A(n4768), .B(n4769), .Z(n4763) );
  NANDN U5056 ( .A(n4770), .B(n4771), .Z(n4769) );
  NANDN U5057 ( .A(n4772), .B(n4773), .Z(n4771) );
  AND U5058 ( .A(B[855]), .B(A[3]), .Z(n4765) );
  XNOR U5059 ( .A(n4755), .B(n4774), .Z(n4766) );
  XNOR U5060 ( .A(n4753), .B(n4756), .Z(n4774) );
  NAND U5061 ( .A(A[2]), .B(B[856]), .Z(n4756) );
  NANDN U5062 ( .A(n4775), .B(n4776), .Z(n4753) );
  AND U5063 ( .A(A[0]), .B(B[857]), .Z(n4776) );
  XOR U5064 ( .A(n4758), .B(n4777), .Z(n4755) );
  NAND U5065 ( .A(A[0]), .B(B[858]), .Z(n4777) );
  NAND U5066 ( .A(B[857]), .B(A[1]), .Z(n4758) );
  NAND U5067 ( .A(n4778), .B(n4779), .Z(n349) );
  NANDN U5068 ( .A(n4780), .B(n4781), .Z(n4779) );
  OR U5069 ( .A(n4782), .B(n4783), .Z(n4781) );
  NAND U5070 ( .A(n4783), .B(n4782), .Z(n4778) );
  XOR U5071 ( .A(n351), .B(n350), .Z(\A1[855] ) );
  XOR U5072 ( .A(n4783), .B(n4784), .Z(n350) );
  XNOR U5073 ( .A(n4782), .B(n4780), .Z(n4784) );
  AND U5074 ( .A(n4785), .B(n4786), .Z(n4780) );
  NANDN U5075 ( .A(n4787), .B(n4788), .Z(n4786) );
  NANDN U5076 ( .A(n4789), .B(n4790), .Z(n4788) );
  AND U5077 ( .A(B[854]), .B(A[3]), .Z(n4782) );
  XNOR U5078 ( .A(n4772), .B(n4791), .Z(n4783) );
  XNOR U5079 ( .A(n4770), .B(n4773), .Z(n4791) );
  NAND U5080 ( .A(A[2]), .B(B[855]), .Z(n4773) );
  NANDN U5081 ( .A(n4792), .B(n4793), .Z(n4770) );
  AND U5082 ( .A(A[0]), .B(B[856]), .Z(n4793) );
  XOR U5083 ( .A(n4775), .B(n4794), .Z(n4772) );
  NAND U5084 ( .A(A[0]), .B(B[857]), .Z(n4794) );
  NAND U5085 ( .A(B[856]), .B(A[1]), .Z(n4775) );
  NAND U5086 ( .A(n4795), .B(n4796), .Z(n351) );
  NANDN U5087 ( .A(n4797), .B(n4798), .Z(n4796) );
  OR U5088 ( .A(n4799), .B(n4800), .Z(n4798) );
  NAND U5089 ( .A(n4800), .B(n4799), .Z(n4795) );
  XOR U5090 ( .A(n353), .B(n352), .Z(\A1[854] ) );
  XOR U5091 ( .A(n4800), .B(n4801), .Z(n352) );
  XNOR U5092 ( .A(n4799), .B(n4797), .Z(n4801) );
  AND U5093 ( .A(n4802), .B(n4803), .Z(n4797) );
  NANDN U5094 ( .A(n4804), .B(n4805), .Z(n4803) );
  NANDN U5095 ( .A(n4806), .B(n4807), .Z(n4805) );
  AND U5096 ( .A(B[853]), .B(A[3]), .Z(n4799) );
  XNOR U5097 ( .A(n4789), .B(n4808), .Z(n4800) );
  XNOR U5098 ( .A(n4787), .B(n4790), .Z(n4808) );
  NAND U5099 ( .A(A[2]), .B(B[854]), .Z(n4790) );
  NANDN U5100 ( .A(n4809), .B(n4810), .Z(n4787) );
  AND U5101 ( .A(A[0]), .B(B[855]), .Z(n4810) );
  XOR U5102 ( .A(n4792), .B(n4811), .Z(n4789) );
  NAND U5103 ( .A(A[0]), .B(B[856]), .Z(n4811) );
  NAND U5104 ( .A(B[855]), .B(A[1]), .Z(n4792) );
  NAND U5105 ( .A(n4812), .B(n4813), .Z(n353) );
  NANDN U5106 ( .A(n4814), .B(n4815), .Z(n4813) );
  OR U5107 ( .A(n4816), .B(n4817), .Z(n4815) );
  NAND U5108 ( .A(n4817), .B(n4816), .Z(n4812) );
  XOR U5109 ( .A(n355), .B(n354), .Z(\A1[853] ) );
  XOR U5110 ( .A(n4817), .B(n4818), .Z(n354) );
  XNOR U5111 ( .A(n4816), .B(n4814), .Z(n4818) );
  AND U5112 ( .A(n4819), .B(n4820), .Z(n4814) );
  NANDN U5113 ( .A(n4821), .B(n4822), .Z(n4820) );
  NANDN U5114 ( .A(n4823), .B(n4824), .Z(n4822) );
  AND U5115 ( .A(B[852]), .B(A[3]), .Z(n4816) );
  XNOR U5116 ( .A(n4806), .B(n4825), .Z(n4817) );
  XNOR U5117 ( .A(n4804), .B(n4807), .Z(n4825) );
  NAND U5118 ( .A(A[2]), .B(B[853]), .Z(n4807) );
  NANDN U5119 ( .A(n4826), .B(n4827), .Z(n4804) );
  AND U5120 ( .A(A[0]), .B(B[854]), .Z(n4827) );
  XOR U5121 ( .A(n4809), .B(n4828), .Z(n4806) );
  NAND U5122 ( .A(A[0]), .B(B[855]), .Z(n4828) );
  NAND U5123 ( .A(B[854]), .B(A[1]), .Z(n4809) );
  NAND U5124 ( .A(n4829), .B(n4830), .Z(n355) );
  NANDN U5125 ( .A(n4831), .B(n4832), .Z(n4830) );
  OR U5126 ( .A(n4833), .B(n4834), .Z(n4832) );
  NAND U5127 ( .A(n4834), .B(n4833), .Z(n4829) );
  XOR U5128 ( .A(n357), .B(n356), .Z(\A1[852] ) );
  XOR U5129 ( .A(n4834), .B(n4835), .Z(n356) );
  XNOR U5130 ( .A(n4833), .B(n4831), .Z(n4835) );
  AND U5131 ( .A(n4836), .B(n4837), .Z(n4831) );
  NANDN U5132 ( .A(n4838), .B(n4839), .Z(n4837) );
  NANDN U5133 ( .A(n4840), .B(n4841), .Z(n4839) );
  AND U5134 ( .A(B[851]), .B(A[3]), .Z(n4833) );
  XNOR U5135 ( .A(n4823), .B(n4842), .Z(n4834) );
  XNOR U5136 ( .A(n4821), .B(n4824), .Z(n4842) );
  NAND U5137 ( .A(A[2]), .B(B[852]), .Z(n4824) );
  NANDN U5138 ( .A(n4843), .B(n4844), .Z(n4821) );
  AND U5139 ( .A(A[0]), .B(B[853]), .Z(n4844) );
  XOR U5140 ( .A(n4826), .B(n4845), .Z(n4823) );
  NAND U5141 ( .A(A[0]), .B(B[854]), .Z(n4845) );
  NAND U5142 ( .A(B[853]), .B(A[1]), .Z(n4826) );
  NAND U5143 ( .A(n4846), .B(n4847), .Z(n357) );
  NANDN U5144 ( .A(n4848), .B(n4849), .Z(n4847) );
  OR U5145 ( .A(n4850), .B(n4851), .Z(n4849) );
  NAND U5146 ( .A(n4851), .B(n4850), .Z(n4846) );
  XOR U5147 ( .A(n359), .B(n358), .Z(\A1[851] ) );
  XOR U5148 ( .A(n4851), .B(n4852), .Z(n358) );
  XNOR U5149 ( .A(n4850), .B(n4848), .Z(n4852) );
  AND U5150 ( .A(n4853), .B(n4854), .Z(n4848) );
  NANDN U5151 ( .A(n4855), .B(n4856), .Z(n4854) );
  NANDN U5152 ( .A(n4857), .B(n4858), .Z(n4856) );
  AND U5153 ( .A(B[850]), .B(A[3]), .Z(n4850) );
  XNOR U5154 ( .A(n4840), .B(n4859), .Z(n4851) );
  XNOR U5155 ( .A(n4838), .B(n4841), .Z(n4859) );
  NAND U5156 ( .A(A[2]), .B(B[851]), .Z(n4841) );
  NANDN U5157 ( .A(n4860), .B(n4861), .Z(n4838) );
  AND U5158 ( .A(A[0]), .B(B[852]), .Z(n4861) );
  XOR U5159 ( .A(n4843), .B(n4862), .Z(n4840) );
  NAND U5160 ( .A(A[0]), .B(B[853]), .Z(n4862) );
  NAND U5161 ( .A(B[852]), .B(A[1]), .Z(n4843) );
  NAND U5162 ( .A(n4863), .B(n4864), .Z(n359) );
  NANDN U5163 ( .A(n4865), .B(n4866), .Z(n4864) );
  OR U5164 ( .A(n4867), .B(n4868), .Z(n4866) );
  NAND U5165 ( .A(n4868), .B(n4867), .Z(n4863) );
  XOR U5166 ( .A(n361), .B(n360), .Z(\A1[850] ) );
  XOR U5167 ( .A(n4868), .B(n4869), .Z(n360) );
  XNOR U5168 ( .A(n4867), .B(n4865), .Z(n4869) );
  AND U5169 ( .A(n4870), .B(n4871), .Z(n4865) );
  NANDN U5170 ( .A(n4872), .B(n4873), .Z(n4871) );
  NANDN U5171 ( .A(n4874), .B(n4875), .Z(n4873) );
  AND U5172 ( .A(B[849]), .B(A[3]), .Z(n4867) );
  XNOR U5173 ( .A(n4857), .B(n4876), .Z(n4868) );
  XNOR U5174 ( .A(n4855), .B(n4858), .Z(n4876) );
  NAND U5175 ( .A(A[2]), .B(B[850]), .Z(n4858) );
  NANDN U5176 ( .A(n4877), .B(n4878), .Z(n4855) );
  AND U5177 ( .A(A[0]), .B(B[851]), .Z(n4878) );
  XOR U5178 ( .A(n4860), .B(n4879), .Z(n4857) );
  NAND U5179 ( .A(A[0]), .B(B[852]), .Z(n4879) );
  NAND U5180 ( .A(B[851]), .B(A[1]), .Z(n4860) );
  NAND U5181 ( .A(n4880), .B(n4881), .Z(n361) );
  NANDN U5182 ( .A(n4882), .B(n4883), .Z(n4881) );
  OR U5183 ( .A(n4884), .B(n4885), .Z(n4883) );
  NAND U5184 ( .A(n4885), .B(n4884), .Z(n4880) );
  XOR U5185 ( .A(n343), .B(n342), .Z(\A1[84] ) );
  XOR U5186 ( .A(n4715), .B(n4886), .Z(n342) );
  XNOR U5187 ( .A(n4714), .B(n4712), .Z(n4886) );
  AND U5188 ( .A(n4887), .B(n4888), .Z(n4712) );
  NANDN U5189 ( .A(n4889), .B(n4890), .Z(n4888) );
  NANDN U5190 ( .A(n4891), .B(n4892), .Z(n4890) );
  AND U5191 ( .A(B[83]), .B(A[3]), .Z(n4714) );
  XNOR U5192 ( .A(n4704), .B(n4893), .Z(n4715) );
  XNOR U5193 ( .A(n4702), .B(n4705), .Z(n4893) );
  NAND U5194 ( .A(A[2]), .B(B[84]), .Z(n4705) );
  NANDN U5195 ( .A(n4894), .B(n4895), .Z(n4702) );
  AND U5196 ( .A(A[0]), .B(B[85]), .Z(n4895) );
  XOR U5197 ( .A(n4707), .B(n4896), .Z(n4704) );
  NAND U5198 ( .A(A[0]), .B(B[86]), .Z(n4896) );
  NAND U5199 ( .A(B[85]), .B(A[1]), .Z(n4707) );
  NAND U5200 ( .A(n4897), .B(n4898), .Z(n343) );
  NANDN U5201 ( .A(n4899), .B(n4900), .Z(n4898) );
  OR U5202 ( .A(n4901), .B(n4902), .Z(n4900) );
  NAND U5203 ( .A(n4902), .B(n4901), .Z(n4897) );
  XOR U5204 ( .A(n363), .B(n362), .Z(\A1[849] ) );
  XOR U5205 ( .A(n4885), .B(n4903), .Z(n362) );
  XNOR U5206 ( .A(n4884), .B(n4882), .Z(n4903) );
  AND U5207 ( .A(n4904), .B(n4905), .Z(n4882) );
  NANDN U5208 ( .A(n4906), .B(n4907), .Z(n4905) );
  NANDN U5209 ( .A(n4908), .B(n4909), .Z(n4907) );
  AND U5210 ( .A(B[848]), .B(A[3]), .Z(n4884) );
  XNOR U5211 ( .A(n4874), .B(n4910), .Z(n4885) );
  XNOR U5212 ( .A(n4872), .B(n4875), .Z(n4910) );
  NAND U5213 ( .A(A[2]), .B(B[849]), .Z(n4875) );
  NANDN U5214 ( .A(n4911), .B(n4912), .Z(n4872) );
  AND U5215 ( .A(A[0]), .B(B[850]), .Z(n4912) );
  XOR U5216 ( .A(n4877), .B(n4913), .Z(n4874) );
  NAND U5217 ( .A(A[0]), .B(B[851]), .Z(n4913) );
  NAND U5218 ( .A(B[850]), .B(A[1]), .Z(n4877) );
  NAND U5219 ( .A(n4914), .B(n4915), .Z(n363) );
  NANDN U5220 ( .A(n4916), .B(n4917), .Z(n4915) );
  OR U5221 ( .A(n4918), .B(n4919), .Z(n4917) );
  NAND U5222 ( .A(n4919), .B(n4918), .Z(n4914) );
  XOR U5223 ( .A(n367), .B(n366), .Z(\A1[848] ) );
  XOR U5224 ( .A(n4919), .B(n4920), .Z(n366) );
  XNOR U5225 ( .A(n4918), .B(n4916), .Z(n4920) );
  AND U5226 ( .A(n4921), .B(n4922), .Z(n4916) );
  NANDN U5227 ( .A(n4923), .B(n4924), .Z(n4922) );
  NANDN U5228 ( .A(n4925), .B(n4926), .Z(n4924) );
  AND U5229 ( .A(B[847]), .B(A[3]), .Z(n4918) );
  XNOR U5230 ( .A(n4908), .B(n4927), .Z(n4919) );
  XNOR U5231 ( .A(n4906), .B(n4909), .Z(n4927) );
  NAND U5232 ( .A(A[2]), .B(B[848]), .Z(n4909) );
  NANDN U5233 ( .A(n4928), .B(n4929), .Z(n4906) );
  AND U5234 ( .A(A[0]), .B(B[849]), .Z(n4929) );
  XOR U5235 ( .A(n4911), .B(n4930), .Z(n4908) );
  NAND U5236 ( .A(A[0]), .B(B[850]), .Z(n4930) );
  NAND U5237 ( .A(B[849]), .B(A[1]), .Z(n4911) );
  NAND U5238 ( .A(n4931), .B(n4932), .Z(n367) );
  NANDN U5239 ( .A(n4933), .B(n4934), .Z(n4932) );
  OR U5240 ( .A(n4935), .B(n4936), .Z(n4934) );
  NAND U5241 ( .A(n4936), .B(n4935), .Z(n4931) );
  XOR U5242 ( .A(n369), .B(n368), .Z(\A1[847] ) );
  XOR U5243 ( .A(n4936), .B(n4937), .Z(n368) );
  XNOR U5244 ( .A(n4935), .B(n4933), .Z(n4937) );
  AND U5245 ( .A(n4938), .B(n4939), .Z(n4933) );
  NANDN U5246 ( .A(n4940), .B(n4941), .Z(n4939) );
  NANDN U5247 ( .A(n4942), .B(n4943), .Z(n4941) );
  AND U5248 ( .A(B[846]), .B(A[3]), .Z(n4935) );
  XNOR U5249 ( .A(n4925), .B(n4944), .Z(n4936) );
  XNOR U5250 ( .A(n4923), .B(n4926), .Z(n4944) );
  NAND U5251 ( .A(A[2]), .B(B[847]), .Z(n4926) );
  NANDN U5252 ( .A(n4945), .B(n4946), .Z(n4923) );
  AND U5253 ( .A(A[0]), .B(B[848]), .Z(n4946) );
  XOR U5254 ( .A(n4928), .B(n4947), .Z(n4925) );
  NAND U5255 ( .A(A[0]), .B(B[849]), .Z(n4947) );
  NAND U5256 ( .A(B[848]), .B(A[1]), .Z(n4928) );
  NAND U5257 ( .A(n4948), .B(n4949), .Z(n369) );
  NANDN U5258 ( .A(n4950), .B(n4951), .Z(n4949) );
  OR U5259 ( .A(n4952), .B(n4953), .Z(n4951) );
  NAND U5260 ( .A(n4953), .B(n4952), .Z(n4948) );
  XOR U5261 ( .A(n371), .B(n370), .Z(\A1[846] ) );
  XOR U5262 ( .A(n4953), .B(n4954), .Z(n370) );
  XNOR U5263 ( .A(n4952), .B(n4950), .Z(n4954) );
  AND U5264 ( .A(n4955), .B(n4956), .Z(n4950) );
  NANDN U5265 ( .A(n4957), .B(n4958), .Z(n4956) );
  NANDN U5266 ( .A(n4959), .B(n4960), .Z(n4958) );
  AND U5267 ( .A(B[845]), .B(A[3]), .Z(n4952) );
  XNOR U5268 ( .A(n4942), .B(n4961), .Z(n4953) );
  XNOR U5269 ( .A(n4940), .B(n4943), .Z(n4961) );
  NAND U5270 ( .A(A[2]), .B(B[846]), .Z(n4943) );
  NANDN U5271 ( .A(n4962), .B(n4963), .Z(n4940) );
  AND U5272 ( .A(A[0]), .B(B[847]), .Z(n4963) );
  XOR U5273 ( .A(n4945), .B(n4964), .Z(n4942) );
  NAND U5274 ( .A(A[0]), .B(B[848]), .Z(n4964) );
  NAND U5275 ( .A(B[847]), .B(A[1]), .Z(n4945) );
  NAND U5276 ( .A(n4965), .B(n4966), .Z(n371) );
  NANDN U5277 ( .A(n4967), .B(n4968), .Z(n4966) );
  OR U5278 ( .A(n4969), .B(n4970), .Z(n4968) );
  NAND U5279 ( .A(n4970), .B(n4969), .Z(n4965) );
  XOR U5280 ( .A(n373), .B(n372), .Z(\A1[845] ) );
  XOR U5281 ( .A(n4970), .B(n4971), .Z(n372) );
  XNOR U5282 ( .A(n4969), .B(n4967), .Z(n4971) );
  AND U5283 ( .A(n4972), .B(n4973), .Z(n4967) );
  NANDN U5284 ( .A(n4974), .B(n4975), .Z(n4973) );
  NANDN U5285 ( .A(n4976), .B(n4977), .Z(n4975) );
  AND U5286 ( .A(B[844]), .B(A[3]), .Z(n4969) );
  XNOR U5287 ( .A(n4959), .B(n4978), .Z(n4970) );
  XNOR U5288 ( .A(n4957), .B(n4960), .Z(n4978) );
  NAND U5289 ( .A(A[2]), .B(B[845]), .Z(n4960) );
  NANDN U5290 ( .A(n4979), .B(n4980), .Z(n4957) );
  AND U5291 ( .A(A[0]), .B(B[846]), .Z(n4980) );
  XOR U5292 ( .A(n4962), .B(n4981), .Z(n4959) );
  NAND U5293 ( .A(A[0]), .B(B[847]), .Z(n4981) );
  NAND U5294 ( .A(B[846]), .B(A[1]), .Z(n4962) );
  NAND U5295 ( .A(n4982), .B(n4983), .Z(n373) );
  NANDN U5296 ( .A(n4984), .B(n4985), .Z(n4983) );
  OR U5297 ( .A(n4986), .B(n4987), .Z(n4985) );
  NAND U5298 ( .A(n4987), .B(n4986), .Z(n4982) );
  XOR U5299 ( .A(n375), .B(n374), .Z(\A1[844] ) );
  XOR U5300 ( .A(n4987), .B(n4988), .Z(n374) );
  XNOR U5301 ( .A(n4986), .B(n4984), .Z(n4988) );
  AND U5302 ( .A(n4989), .B(n4990), .Z(n4984) );
  NANDN U5303 ( .A(n4991), .B(n4992), .Z(n4990) );
  NANDN U5304 ( .A(n4993), .B(n4994), .Z(n4992) );
  AND U5305 ( .A(B[843]), .B(A[3]), .Z(n4986) );
  XNOR U5306 ( .A(n4976), .B(n4995), .Z(n4987) );
  XNOR U5307 ( .A(n4974), .B(n4977), .Z(n4995) );
  NAND U5308 ( .A(A[2]), .B(B[844]), .Z(n4977) );
  NANDN U5309 ( .A(n4996), .B(n4997), .Z(n4974) );
  AND U5310 ( .A(A[0]), .B(B[845]), .Z(n4997) );
  XOR U5311 ( .A(n4979), .B(n4998), .Z(n4976) );
  NAND U5312 ( .A(A[0]), .B(B[846]), .Z(n4998) );
  NAND U5313 ( .A(B[845]), .B(A[1]), .Z(n4979) );
  NAND U5314 ( .A(n4999), .B(n5000), .Z(n375) );
  NANDN U5315 ( .A(n5001), .B(n5002), .Z(n5000) );
  OR U5316 ( .A(n5003), .B(n5004), .Z(n5002) );
  NAND U5317 ( .A(n5004), .B(n5003), .Z(n4999) );
  XOR U5318 ( .A(n377), .B(n376), .Z(\A1[843] ) );
  XOR U5319 ( .A(n5004), .B(n5005), .Z(n376) );
  XNOR U5320 ( .A(n5003), .B(n5001), .Z(n5005) );
  AND U5321 ( .A(n5006), .B(n5007), .Z(n5001) );
  NANDN U5322 ( .A(n5008), .B(n5009), .Z(n5007) );
  NANDN U5323 ( .A(n5010), .B(n5011), .Z(n5009) );
  AND U5324 ( .A(B[842]), .B(A[3]), .Z(n5003) );
  XNOR U5325 ( .A(n4993), .B(n5012), .Z(n5004) );
  XNOR U5326 ( .A(n4991), .B(n4994), .Z(n5012) );
  NAND U5327 ( .A(A[2]), .B(B[843]), .Z(n4994) );
  NANDN U5328 ( .A(n5013), .B(n5014), .Z(n4991) );
  AND U5329 ( .A(A[0]), .B(B[844]), .Z(n5014) );
  XOR U5330 ( .A(n4996), .B(n5015), .Z(n4993) );
  NAND U5331 ( .A(A[0]), .B(B[845]), .Z(n5015) );
  NAND U5332 ( .A(B[844]), .B(A[1]), .Z(n4996) );
  NAND U5333 ( .A(n5016), .B(n5017), .Z(n377) );
  NANDN U5334 ( .A(n5018), .B(n5019), .Z(n5017) );
  OR U5335 ( .A(n5020), .B(n5021), .Z(n5019) );
  NAND U5336 ( .A(n5021), .B(n5020), .Z(n5016) );
  XOR U5337 ( .A(n379), .B(n378), .Z(\A1[842] ) );
  XOR U5338 ( .A(n5021), .B(n5022), .Z(n378) );
  XNOR U5339 ( .A(n5020), .B(n5018), .Z(n5022) );
  AND U5340 ( .A(n5023), .B(n5024), .Z(n5018) );
  NANDN U5341 ( .A(n5025), .B(n5026), .Z(n5024) );
  NANDN U5342 ( .A(n5027), .B(n5028), .Z(n5026) );
  AND U5343 ( .A(B[841]), .B(A[3]), .Z(n5020) );
  XNOR U5344 ( .A(n5010), .B(n5029), .Z(n5021) );
  XNOR U5345 ( .A(n5008), .B(n5011), .Z(n5029) );
  NAND U5346 ( .A(A[2]), .B(B[842]), .Z(n5011) );
  NANDN U5347 ( .A(n5030), .B(n5031), .Z(n5008) );
  AND U5348 ( .A(A[0]), .B(B[843]), .Z(n5031) );
  XOR U5349 ( .A(n5013), .B(n5032), .Z(n5010) );
  NAND U5350 ( .A(A[0]), .B(B[844]), .Z(n5032) );
  NAND U5351 ( .A(B[843]), .B(A[1]), .Z(n5013) );
  NAND U5352 ( .A(n5033), .B(n5034), .Z(n379) );
  NANDN U5353 ( .A(n5035), .B(n5036), .Z(n5034) );
  OR U5354 ( .A(n5037), .B(n5038), .Z(n5036) );
  NAND U5355 ( .A(n5038), .B(n5037), .Z(n5033) );
  XOR U5356 ( .A(n381), .B(n380), .Z(\A1[841] ) );
  XOR U5357 ( .A(n5038), .B(n5039), .Z(n380) );
  XNOR U5358 ( .A(n5037), .B(n5035), .Z(n5039) );
  AND U5359 ( .A(n5040), .B(n5041), .Z(n5035) );
  NANDN U5360 ( .A(n5042), .B(n5043), .Z(n5041) );
  NANDN U5361 ( .A(n5044), .B(n5045), .Z(n5043) );
  AND U5362 ( .A(B[840]), .B(A[3]), .Z(n5037) );
  XNOR U5363 ( .A(n5027), .B(n5046), .Z(n5038) );
  XNOR U5364 ( .A(n5025), .B(n5028), .Z(n5046) );
  NAND U5365 ( .A(A[2]), .B(B[841]), .Z(n5028) );
  NANDN U5366 ( .A(n5047), .B(n5048), .Z(n5025) );
  AND U5367 ( .A(A[0]), .B(B[842]), .Z(n5048) );
  XOR U5368 ( .A(n5030), .B(n5049), .Z(n5027) );
  NAND U5369 ( .A(A[0]), .B(B[843]), .Z(n5049) );
  NAND U5370 ( .A(B[842]), .B(A[1]), .Z(n5030) );
  NAND U5371 ( .A(n5050), .B(n5051), .Z(n381) );
  NANDN U5372 ( .A(n5052), .B(n5053), .Z(n5051) );
  OR U5373 ( .A(n5054), .B(n5055), .Z(n5053) );
  NAND U5374 ( .A(n5055), .B(n5054), .Z(n5050) );
  XOR U5375 ( .A(n383), .B(n382), .Z(\A1[840] ) );
  XOR U5376 ( .A(n5055), .B(n5056), .Z(n382) );
  XNOR U5377 ( .A(n5054), .B(n5052), .Z(n5056) );
  AND U5378 ( .A(n5057), .B(n5058), .Z(n5052) );
  NANDN U5379 ( .A(n5059), .B(n5060), .Z(n5058) );
  NANDN U5380 ( .A(n5061), .B(n5062), .Z(n5060) );
  AND U5381 ( .A(B[839]), .B(A[3]), .Z(n5054) );
  XNOR U5382 ( .A(n5044), .B(n5063), .Z(n5055) );
  XNOR U5383 ( .A(n5042), .B(n5045), .Z(n5063) );
  NAND U5384 ( .A(A[2]), .B(B[840]), .Z(n5045) );
  NANDN U5385 ( .A(n5064), .B(n5065), .Z(n5042) );
  AND U5386 ( .A(A[0]), .B(B[841]), .Z(n5065) );
  XOR U5387 ( .A(n5047), .B(n5066), .Z(n5044) );
  NAND U5388 ( .A(A[0]), .B(B[842]), .Z(n5066) );
  NAND U5389 ( .A(B[841]), .B(A[1]), .Z(n5047) );
  NAND U5390 ( .A(n5067), .B(n5068), .Z(n383) );
  NANDN U5391 ( .A(n5069), .B(n5070), .Z(n5068) );
  OR U5392 ( .A(n5071), .B(n5072), .Z(n5070) );
  NAND U5393 ( .A(n5072), .B(n5071), .Z(n5067) );
  XOR U5394 ( .A(n365), .B(n364), .Z(\A1[83] ) );
  XOR U5395 ( .A(n4902), .B(n5073), .Z(n364) );
  XNOR U5396 ( .A(n4901), .B(n4899), .Z(n5073) );
  AND U5397 ( .A(n5074), .B(n5075), .Z(n4899) );
  NANDN U5398 ( .A(n5076), .B(n5077), .Z(n5075) );
  NANDN U5399 ( .A(n5078), .B(n5079), .Z(n5077) );
  AND U5400 ( .A(B[82]), .B(A[3]), .Z(n4901) );
  XNOR U5401 ( .A(n4891), .B(n5080), .Z(n4902) );
  XNOR U5402 ( .A(n4889), .B(n4892), .Z(n5080) );
  NAND U5403 ( .A(A[2]), .B(B[83]), .Z(n4892) );
  NANDN U5404 ( .A(n5081), .B(n5082), .Z(n4889) );
  AND U5405 ( .A(A[0]), .B(B[84]), .Z(n5082) );
  XOR U5406 ( .A(n4894), .B(n5083), .Z(n4891) );
  NAND U5407 ( .A(A[0]), .B(B[85]), .Z(n5083) );
  NAND U5408 ( .A(B[84]), .B(A[1]), .Z(n4894) );
  NAND U5409 ( .A(n5084), .B(n5085), .Z(n365) );
  NANDN U5410 ( .A(n5086), .B(n5087), .Z(n5085) );
  OR U5411 ( .A(n5088), .B(n5089), .Z(n5087) );
  NAND U5412 ( .A(n5089), .B(n5088), .Z(n5084) );
  XOR U5413 ( .A(n385), .B(n384), .Z(\A1[839] ) );
  XOR U5414 ( .A(n5072), .B(n5090), .Z(n384) );
  XNOR U5415 ( .A(n5071), .B(n5069), .Z(n5090) );
  AND U5416 ( .A(n5091), .B(n5092), .Z(n5069) );
  NANDN U5417 ( .A(n5093), .B(n5094), .Z(n5092) );
  NANDN U5418 ( .A(n5095), .B(n5096), .Z(n5094) );
  AND U5419 ( .A(B[838]), .B(A[3]), .Z(n5071) );
  XNOR U5420 ( .A(n5061), .B(n5097), .Z(n5072) );
  XNOR U5421 ( .A(n5059), .B(n5062), .Z(n5097) );
  NAND U5422 ( .A(A[2]), .B(B[839]), .Z(n5062) );
  NANDN U5423 ( .A(n5098), .B(n5099), .Z(n5059) );
  AND U5424 ( .A(A[0]), .B(B[840]), .Z(n5099) );
  XOR U5425 ( .A(n5064), .B(n5100), .Z(n5061) );
  NAND U5426 ( .A(A[0]), .B(B[841]), .Z(n5100) );
  NAND U5427 ( .A(B[840]), .B(A[1]), .Z(n5064) );
  NAND U5428 ( .A(n5101), .B(n5102), .Z(n385) );
  NANDN U5429 ( .A(n5103), .B(n5104), .Z(n5102) );
  OR U5430 ( .A(n5105), .B(n5106), .Z(n5104) );
  NAND U5431 ( .A(n5106), .B(n5105), .Z(n5101) );
  XOR U5432 ( .A(n389), .B(n388), .Z(\A1[838] ) );
  XOR U5433 ( .A(n5106), .B(n5107), .Z(n388) );
  XNOR U5434 ( .A(n5105), .B(n5103), .Z(n5107) );
  AND U5435 ( .A(n5108), .B(n5109), .Z(n5103) );
  NANDN U5436 ( .A(n5110), .B(n5111), .Z(n5109) );
  NANDN U5437 ( .A(n5112), .B(n5113), .Z(n5111) );
  AND U5438 ( .A(B[837]), .B(A[3]), .Z(n5105) );
  XNOR U5439 ( .A(n5095), .B(n5114), .Z(n5106) );
  XNOR U5440 ( .A(n5093), .B(n5096), .Z(n5114) );
  NAND U5441 ( .A(A[2]), .B(B[838]), .Z(n5096) );
  NANDN U5442 ( .A(n5115), .B(n5116), .Z(n5093) );
  AND U5443 ( .A(A[0]), .B(B[839]), .Z(n5116) );
  XOR U5444 ( .A(n5098), .B(n5117), .Z(n5095) );
  NAND U5445 ( .A(A[0]), .B(B[840]), .Z(n5117) );
  NAND U5446 ( .A(B[839]), .B(A[1]), .Z(n5098) );
  NAND U5447 ( .A(n5118), .B(n5119), .Z(n389) );
  NANDN U5448 ( .A(n5120), .B(n5121), .Z(n5119) );
  OR U5449 ( .A(n5122), .B(n5123), .Z(n5121) );
  NAND U5450 ( .A(n5123), .B(n5122), .Z(n5118) );
  XOR U5451 ( .A(n391), .B(n390), .Z(\A1[837] ) );
  XOR U5452 ( .A(n5123), .B(n5124), .Z(n390) );
  XNOR U5453 ( .A(n5122), .B(n5120), .Z(n5124) );
  AND U5454 ( .A(n5125), .B(n5126), .Z(n5120) );
  NANDN U5455 ( .A(n5127), .B(n5128), .Z(n5126) );
  NANDN U5456 ( .A(n5129), .B(n5130), .Z(n5128) );
  AND U5457 ( .A(B[836]), .B(A[3]), .Z(n5122) );
  XNOR U5458 ( .A(n5112), .B(n5131), .Z(n5123) );
  XNOR U5459 ( .A(n5110), .B(n5113), .Z(n5131) );
  NAND U5460 ( .A(A[2]), .B(B[837]), .Z(n5113) );
  NANDN U5461 ( .A(n5132), .B(n5133), .Z(n5110) );
  AND U5462 ( .A(A[0]), .B(B[838]), .Z(n5133) );
  XOR U5463 ( .A(n5115), .B(n5134), .Z(n5112) );
  NAND U5464 ( .A(A[0]), .B(B[839]), .Z(n5134) );
  NAND U5465 ( .A(B[838]), .B(A[1]), .Z(n5115) );
  NAND U5466 ( .A(n5135), .B(n5136), .Z(n391) );
  NANDN U5467 ( .A(n5137), .B(n5138), .Z(n5136) );
  OR U5468 ( .A(n5139), .B(n5140), .Z(n5138) );
  NAND U5469 ( .A(n5140), .B(n5139), .Z(n5135) );
  XOR U5470 ( .A(n393), .B(n392), .Z(\A1[836] ) );
  XOR U5471 ( .A(n5140), .B(n5141), .Z(n392) );
  XNOR U5472 ( .A(n5139), .B(n5137), .Z(n5141) );
  AND U5473 ( .A(n5142), .B(n5143), .Z(n5137) );
  NANDN U5474 ( .A(n5144), .B(n5145), .Z(n5143) );
  NANDN U5475 ( .A(n5146), .B(n5147), .Z(n5145) );
  AND U5476 ( .A(B[835]), .B(A[3]), .Z(n5139) );
  XNOR U5477 ( .A(n5129), .B(n5148), .Z(n5140) );
  XNOR U5478 ( .A(n5127), .B(n5130), .Z(n5148) );
  NAND U5479 ( .A(A[2]), .B(B[836]), .Z(n5130) );
  NANDN U5480 ( .A(n5149), .B(n5150), .Z(n5127) );
  AND U5481 ( .A(A[0]), .B(B[837]), .Z(n5150) );
  XOR U5482 ( .A(n5132), .B(n5151), .Z(n5129) );
  NAND U5483 ( .A(A[0]), .B(B[838]), .Z(n5151) );
  NAND U5484 ( .A(B[837]), .B(A[1]), .Z(n5132) );
  NAND U5485 ( .A(n5152), .B(n5153), .Z(n393) );
  NANDN U5486 ( .A(n5154), .B(n5155), .Z(n5153) );
  OR U5487 ( .A(n5156), .B(n5157), .Z(n5155) );
  NAND U5488 ( .A(n5157), .B(n5156), .Z(n5152) );
  XOR U5489 ( .A(n395), .B(n394), .Z(\A1[835] ) );
  XOR U5490 ( .A(n5157), .B(n5158), .Z(n394) );
  XNOR U5491 ( .A(n5156), .B(n5154), .Z(n5158) );
  AND U5492 ( .A(n5159), .B(n5160), .Z(n5154) );
  NANDN U5493 ( .A(n5161), .B(n5162), .Z(n5160) );
  NANDN U5494 ( .A(n5163), .B(n5164), .Z(n5162) );
  AND U5495 ( .A(B[834]), .B(A[3]), .Z(n5156) );
  XNOR U5496 ( .A(n5146), .B(n5165), .Z(n5157) );
  XNOR U5497 ( .A(n5144), .B(n5147), .Z(n5165) );
  NAND U5498 ( .A(A[2]), .B(B[835]), .Z(n5147) );
  NANDN U5499 ( .A(n5166), .B(n5167), .Z(n5144) );
  AND U5500 ( .A(A[0]), .B(B[836]), .Z(n5167) );
  XOR U5501 ( .A(n5149), .B(n5168), .Z(n5146) );
  NAND U5502 ( .A(A[0]), .B(B[837]), .Z(n5168) );
  NAND U5503 ( .A(B[836]), .B(A[1]), .Z(n5149) );
  NAND U5504 ( .A(n5169), .B(n5170), .Z(n395) );
  NANDN U5505 ( .A(n5171), .B(n5172), .Z(n5170) );
  OR U5506 ( .A(n5173), .B(n5174), .Z(n5172) );
  NAND U5507 ( .A(n5174), .B(n5173), .Z(n5169) );
  XOR U5508 ( .A(n397), .B(n396), .Z(\A1[834] ) );
  XOR U5509 ( .A(n5174), .B(n5175), .Z(n396) );
  XNOR U5510 ( .A(n5173), .B(n5171), .Z(n5175) );
  AND U5511 ( .A(n5176), .B(n5177), .Z(n5171) );
  NANDN U5512 ( .A(n5178), .B(n5179), .Z(n5177) );
  NANDN U5513 ( .A(n5180), .B(n5181), .Z(n5179) );
  AND U5514 ( .A(B[833]), .B(A[3]), .Z(n5173) );
  XNOR U5515 ( .A(n5163), .B(n5182), .Z(n5174) );
  XNOR U5516 ( .A(n5161), .B(n5164), .Z(n5182) );
  NAND U5517 ( .A(A[2]), .B(B[834]), .Z(n5164) );
  NANDN U5518 ( .A(n5183), .B(n5184), .Z(n5161) );
  AND U5519 ( .A(A[0]), .B(B[835]), .Z(n5184) );
  XOR U5520 ( .A(n5166), .B(n5185), .Z(n5163) );
  NAND U5521 ( .A(A[0]), .B(B[836]), .Z(n5185) );
  NAND U5522 ( .A(B[835]), .B(A[1]), .Z(n5166) );
  NAND U5523 ( .A(n5186), .B(n5187), .Z(n397) );
  NANDN U5524 ( .A(n5188), .B(n5189), .Z(n5187) );
  OR U5525 ( .A(n5190), .B(n5191), .Z(n5189) );
  NAND U5526 ( .A(n5191), .B(n5190), .Z(n5186) );
  XOR U5527 ( .A(n399), .B(n398), .Z(\A1[833] ) );
  XOR U5528 ( .A(n5191), .B(n5192), .Z(n398) );
  XNOR U5529 ( .A(n5190), .B(n5188), .Z(n5192) );
  AND U5530 ( .A(n5193), .B(n5194), .Z(n5188) );
  NANDN U5531 ( .A(n5195), .B(n5196), .Z(n5194) );
  NANDN U5532 ( .A(n5197), .B(n5198), .Z(n5196) );
  AND U5533 ( .A(B[832]), .B(A[3]), .Z(n5190) );
  XNOR U5534 ( .A(n5180), .B(n5199), .Z(n5191) );
  XNOR U5535 ( .A(n5178), .B(n5181), .Z(n5199) );
  NAND U5536 ( .A(A[2]), .B(B[833]), .Z(n5181) );
  NANDN U5537 ( .A(n5200), .B(n5201), .Z(n5178) );
  AND U5538 ( .A(A[0]), .B(B[834]), .Z(n5201) );
  XOR U5539 ( .A(n5183), .B(n5202), .Z(n5180) );
  NAND U5540 ( .A(A[0]), .B(B[835]), .Z(n5202) );
  NAND U5541 ( .A(B[834]), .B(A[1]), .Z(n5183) );
  NAND U5542 ( .A(n5203), .B(n5204), .Z(n399) );
  NANDN U5543 ( .A(n5205), .B(n5206), .Z(n5204) );
  OR U5544 ( .A(n5207), .B(n5208), .Z(n5206) );
  NAND U5545 ( .A(n5208), .B(n5207), .Z(n5203) );
  XOR U5546 ( .A(n401), .B(n400), .Z(\A1[832] ) );
  XOR U5547 ( .A(n5208), .B(n5209), .Z(n400) );
  XNOR U5548 ( .A(n5207), .B(n5205), .Z(n5209) );
  AND U5549 ( .A(n5210), .B(n5211), .Z(n5205) );
  NANDN U5550 ( .A(n5212), .B(n5213), .Z(n5211) );
  NANDN U5551 ( .A(n5214), .B(n5215), .Z(n5213) );
  AND U5552 ( .A(B[831]), .B(A[3]), .Z(n5207) );
  XNOR U5553 ( .A(n5197), .B(n5216), .Z(n5208) );
  XNOR U5554 ( .A(n5195), .B(n5198), .Z(n5216) );
  NAND U5555 ( .A(A[2]), .B(B[832]), .Z(n5198) );
  NANDN U5556 ( .A(n5217), .B(n5218), .Z(n5195) );
  AND U5557 ( .A(A[0]), .B(B[833]), .Z(n5218) );
  XOR U5558 ( .A(n5200), .B(n5219), .Z(n5197) );
  NAND U5559 ( .A(A[0]), .B(B[834]), .Z(n5219) );
  NAND U5560 ( .A(B[833]), .B(A[1]), .Z(n5200) );
  NAND U5561 ( .A(n5220), .B(n5221), .Z(n401) );
  NANDN U5562 ( .A(n5222), .B(n5223), .Z(n5221) );
  OR U5563 ( .A(n5224), .B(n5225), .Z(n5223) );
  NAND U5564 ( .A(n5225), .B(n5224), .Z(n5220) );
  XOR U5565 ( .A(n403), .B(n402), .Z(\A1[831] ) );
  XOR U5566 ( .A(n5225), .B(n5226), .Z(n402) );
  XNOR U5567 ( .A(n5224), .B(n5222), .Z(n5226) );
  AND U5568 ( .A(n5227), .B(n5228), .Z(n5222) );
  NANDN U5569 ( .A(n5229), .B(n5230), .Z(n5228) );
  NANDN U5570 ( .A(n5231), .B(n5232), .Z(n5230) );
  AND U5571 ( .A(B[830]), .B(A[3]), .Z(n5224) );
  XNOR U5572 ( .A(n5214), .B(n5233), .Z(n5225) );
  XNOR U5573 ( .A(n5212), .B(n5215), .Z(n5233) );
  NAND U5574 ( .A(A[2]), .B(B[831]), .Z(n5215) );
  NANDN U5575 ( .A(n5234), .B(n5235), .Z(n5212) );
  AND U5576 ( .A(A[0]), .B(B[832]), .Z(n5235) );
  XOR U5577 ( .A(n5217), .B(n5236), .Z(n5214) );
  NAND U5578 ( .A(A[0]), .B(B[833]), .Z(n5236) );
  NAND U5579 ( .A(B[832]), .B(A[1]), .Z(n5217) );
  NAND U5580 ( .A(n5237), .B(n5238), .Z(n403) );
  NANDN U5581 ( .A(n5239), .B(n5240), .Z(n5238) );
  OR U5582 ( .A(n5241), .B(n5242), .Z(n5240) );
  NAND U5583 ( .A(n5242), .B(n5241), .Z(n5237) );
  XOR U5584 ( .A(n405), .B(n404), .Z(\A1[830] ) );
  XOR U5585 ( .A(n5242), .B(n5243), .Z(n404) );
  XNOR U5586 ( .A(n5241), .B(n5239), .Z(n5243) );
  AND U5587 ( .A(n5244), .B(n5245), .Z(n5239) );
  NANDN U5588 ( .A(n5246), .B(n5247), .Z(n5245) );
  NANDN U5589 ( .A(n5248), .B(n5249), .Z(n5247) );
  AND U5590 ( .A(B[829]), .B(A[3]), .Z(n5241) );
  XNOR U5591 ( .A(n5231), .B(n5250), .Z(n5242) );
  XNOR U5592 ( .A(n5229), .B(n5232), .Z(n5250) );
  NAND U5593 ( .A(A[2]), .B(B[830]), .Z(n5232) );
  NANDN U5594 ( .A(n5251), .B(n5252), .Z(n5229) );
  AND U5595 ( .A(A[0]), .B(B[831]), .Z(n5252) );
  XOR U5596 ( .A(n5234), .B(n5253), .Z(n5231) );
  NAND U5597 ( .A(A[0]), .B(B[832]), .Z(n5253) );
  NAND U5598 ( .A(B[831]), .B(A[1]), .Z(n5234) );
  NAND U5599 ( .A(n5254), .B(n5255), .Z(n405) );
  NANDN U5600 ( .A(n5256), .B(n5257), .Z(n5255) );
  OR U5601 ( .A(n5258), .B(n5259), .Z(n5257) );
  NAND U5602 ( .A(n5259), .B(n5258), .Z(n5254) );
  XOR U5603 ( .A(n387), .B(n386), .Z(\A1[82] ) );
  XOR U5604 ( .A(n5089), .B(n5260), .Z(n386) );
  XNOR U5605 ( .A(n5088), .B(n5086), .Z(n5260) );
  AND U5606 ( .A(n5261), .B(n5262), .Z(n5086) );
  NANDN U5607 ( .A(n5263), .B(n5264), .Z(n5262) );
  NANDN U5608 ( .A(n5265), .B(n5266), .Z(n5264) );
  AND U5609 ( .A(B[81]), .B(A[3]), .Z(n5088) );
  XNOR U5610 ( .A(n5078), .B(n5267), .Z(n5089) );
  XNOR U5611 ( .A(n5076), .B(n5079), .Z(n5267) );
  NAND U5612 ( .A(A[2]), .B(B[82]), .Z(n5079) );
  NANDN U5613 ( .A(n5268), .B(n5269), .Z(n5076) );
  AND U5614 ( .A(A[0]), .B(B[83]), .Z(n5269) );
  XOR U5615 ( .A(n5081), .B(n5270), .Z(n5078) );
  NAND U5616 ( .A(A[0]), .B(B[84]), .Z(n5270) );
  NAND U5617 ( .A(B[83]), .B(A[1]), .Z(n5081) );
  NAND U5618 ( .A(n5271), .B(n5272), .Z(n387) );
  NANDN U5619 ( .A(n5273), .B(n5274), .Z(n5272) );
  OR U5620 ( .A(n5275), .B(n5276), .Z(n5274) );
  NAND U5621 ( .A(n5276), .B(n5275), .Z(n5271) );
  XOR U5622 ( .A(n407), .B(n406), .Z(\A1[829] ) );
  XOR U5623 ( .A(n5259), .B(n5277), .Z(n406) );
  XNOR U5624 ( .A(n5258), .B(n5256), .Z(n5277) );
  AND U5625 ( .A(n5278), .B(n5279), .Z(n5256) );
  NANDN U5626 ( .A(n5280), .B(n5281), .Z(n5279) );
  NANDN U5627 ( .A(n5282), .B(n5283), .Z(n5281) );
  AND U5628 ( .A(B[828]), .B(A[3]), .Z(n5258) );
  XNOR U5629 ( .A(n5248), .B(n5284), .Z(n5259) );
  XNOR U5630 ( .A(n5246), .B(n5249), .Z(n5284) );
  NAND U5631 ( .A(A[2]), .B(B[829]), .Z(n5249) );
  NANDN U5632 ( .A(n5285), .B(n5286), .Z(n5246) );
  AND U5633 ( .A(A[0]), .B(B[830]), .Z(n5286) );
  XOR U5634 ( .A(n5251), .B(n5287), .Z(n5248) );
  NAND U5635 ( .A(A[0]), .B(B[831]), .Z(n5287) );
  NAND U5636 ( .A(B[830]), .B(A[1]), .Z(n5251) );
  NAND U5637 ( .A(n5288), .B(n5289), .Z(n407) );
  NANDN U5638 ( .A(n5290), .B(n5291), .Z(n5289) );
  OR U5639 ( .A(n5292), .B(n5293), .Z(n5291) );
  NAND U5640 ( .A(n5293), .B(n5292), .Z(n5288) );
  XOR U5641 ( .A(n411), .B(n410), .Z(\A1[828] ) );
  XOR U5642 ( .A(n5293), .B(n5294), .Z(n410) );
  XNOR U5643 ( .A(n5292), .B(n5290), .Z(n5294) );
  AND U5644 ( .A(n5295), .B(n5296), .Z(n5290) );
  NANDN U5645 ( .A(n5297), .B(n5298), .Z(n5296) );
  NANDN U5646 ( .A(n5299), .B(n5300), .Z(n5298) );
  AND U5647 ( .A(B[827]), .B(A[3]), .Z(n5292) );
  XNOR U5648 ( .A(n5282), .B(n5301), .Z(n5293) );
  XNOR U5649 ( .A(n5280), .B(n5283), .Z(n5301) );
  NAND U5650 ( .A(A[2]), .B(B[828]), .Z(n5283) );
  NANDN U5651 ( .A(n5302), .B(n5303), .Z(n5280) );
  AND U5652 ( .A(A[0]), .B(B[829]), .Z(n5303) );
  XOR U5653 ( .A(n5285), .B(n5304), .Z(n5282) );
  NAND U5654 ( .A(A[0]), .B(B[830]), .Z(n5304) );
  NAND U5655 ( .A(B[829]), .B(A[1]), .Z(n5285) );
  NAND U5656 ( .A(n5305), .B(n5306), .Z(n411) );
  NANDN U5657 ( .A(n5307), .B(n5308), .Z(n5306) );
  OR U5658 ( .A(n5309), .B(n5310), .Z(n5308) );
  NAND U5659 ( .A(n5310), .B(n5309), .Z(n5305) );
  XOR U5660 ( .A(n413), .B(n412), .Z(\A1[827] ) );
  XOR U5661 ( .A(n5310), .B(n5311), .Z(n412) );
  XNOR U5662 ( .A(n5309), .B(n5307), .Z(n5311) );
  AND U5663 ( .A(n5312), .B(n5313), .Z(n5307) );
  NANDN U5664 ( .A(n5314), .B(n5315), .Z(n5313) );
  NANDN U5665 ( .A(n5316), .B(n5317), .Z(n5315) );
  AND U5666 ( .A(B[826]), .B(A[3]), .Z(n5309) );
  XNOR U5667 ( .A(n5299), .B(n5318), .Z(n5310) );
  XNOR U5668 ( .A(n5297), .B(n5300), .Z(n5318) );
  NAND U5669 ( .A(A[2]), .B(B[827]), .Z(n5300) );
  NANDN U5670 ( .A(n5319), .B(n5320), .Z(n5297) );
  AND U5671 ( .A(A[0]), .B(B[828]), .Z(n5320) );
  XOR U5672 ( .A(n5302), .B(n5321), .Z(n5299) );
  NAND U5673 ( .A(A[0]), .B(B[829]), .Z(n5321) );
  NAND U5674 ( .A(B[828]), .B(A[1]), .Z(n5302) );
  NAND U5675 ( .A(n5322), .B(n5323), .Z(n413) );
  NANDN U5676 ( .A(n5324), .B(n5325), .Z(n5323) );
  OR U5677 ( .A(n5326), .B(n5327), .Z(n5325) );
  NAND U5678 ( .A(n5327), .B(n5326), .Z(n5322) );
  XOR U5679 ( .A(n415), .B(n414), .Z(\A1[826] ) );
  XOR U5680 ( .A(n5327), .B(n5328), .Z(n414) );
  XNOR U5681 ( .A(n5326), .B(n5324), .Z(n5328) );
  AND U5682 ( .A(n5329), .B(n5330), .Z(n5324) );
  NANDN U5683 ( .A(n5331), .B(n5332), .Z(n5330) );
  NANDN U5684 ( .A(n5333), .B(n5334), .Z(n5332) );
  AND U5685 ( .A(B[825]), .B(A[3]), .Z(n5326) );
  XNOR U5686 ( .A(n5316), .B(n5335), .Z(n5327) );
  XNOR U5687 ( .A(n5314), .B(n5317), .Z(n5335) );
  NAND U5688 ( .A(A[2]), .B(B[826]), .Z(n5317) );
  NANDN U5689 ( .A(n5336), .B(n5337), .Z(n5314) );
  AND U5690 ( .A(A[0]), .B(B[827]), .Z(n5337) );
  XOR U5691 ( .A(n5319), .B(n5338), .Z(n5316) );
  NAND U5692 ( .A(A[0]), .B(B[828]), .Z(n5338) );
  NAND U5693 ( .A(B[827]), .B(A[1]), .Z(n5319) );
  NAND U5694 ( .A(n5339), .B(n5340), .Z(n415) );
  NANDN U5695 ( .A(n5341), .B(n5342), .Z(n5340) );
  OR U5696 ( .A(n5343), .B(n5344), .Z(n5342) );
  NAND U5697 ( .A(n5344), .B(n5343), .Z(n5339) );
  XOR U5698 ( .A(n417), .B(n416), .Z(\A1[825] ) );
  XOR U5699 ( .A(n5344), .B(n5345), .Z(n416) );
  XNOR U5700 ( .A(n5343), .B(n5341), .Z(n5345) );
  AND U5701 ( .A(n5346), .B(n5347), .Z(n5341) );
  NANDN U5702 ( .A(n5348), .B(n5349), .Z(n5347) );
  NANDN U5703 ( .A(n5350), .B(n5351), .Z(n5349) );
  AND U5704 ( .A(B[824]), .B(A[3]), .Z(n5343) );
  XNOR U5705 ( .A(n5333), .B(n5352), .Z(n5344) );
  XNOR U5706 ( .A(n5331), .B(n5334), .Z(n5352) );
  NAND U5707 ( .A(A[2]), .B(B[825]), .Z(n5334) );
  NANDN U5708 ( .A(n5353), .B(n5354), .Z(n5331) );
  AND U5709 ( .A(A[0]), .B(B[826]), .Z(n5354) );
  XOR U5710 ( .A(n5336), .B(n5355), .Z(n5333) );
  NAND U5711 ( .A(A[0]), .B(B[827]), .Z(n5355) );
  NAND U5712 ( .A(B[826]), .B(A[1]), .Z(n5336) );
  NAND U5713 ( .A(n5356), .B(n5357), .Z(n417) );
  NANDN U5714 ( .A(n5358), .B(n5359), .Z(n5357) );
  OR U5715 ( .A(n5360), .B(n5361), .Z(n5359) );
  NAND U5716 ( .A(n5361), .B(n5360), .Z(n5356) );
  XOR U5717 ( .A(n419), .B(n418), .Z(\A1[824] ) );
  XOR U5718 ( .A(n5361), .B(n5362), .Z(n418) );
  XNOR U5719 ( .A(n5360), .B(n5358), .Z(n5362) );
  AND U5720 ( .A(n5363), .B(n5364), .Z(n5358) );
  NANDN U5721 ( .A(n5365), .B(n5366), .Z(n5364) );
  NANDN U5722 ( .A(n5367), .B(n5368), .Z(n5366) );
  AND U5723 ( .A(B[823]), .B(A[3]), .Z(n5360) );
  XNOR U5724 ( .A(n5350), .B(n5369), .Z(n5361) );
  XNOR U5725 ( .A(n5348), .B(n5351), .Z(n5369) );
  NAND U5726 ( .A(A[2]), .B(B[824]), .Z(n5351) );
  NANDN U5727 ( .A(n5370), .B(n5371), .Z(n5348) );
  AND U5728 ( .A(A[0]), .B(B[825]), .Z(n5371) );
  XOR U5729 ( .A(n5353), .B(n5372), .Z(n5350) );
  NAND U5730 ( .A(A[0]), .B(B[826]), .Z(n5372) );
  NAND U5731 ( .A(B[825]), .B(A[1]), .Z(n5353) );
  NAND U5732 ( .A(n5373), .B(n5374), .Z(n419) );
  NANDN U5733 ( .A(n5375), .B(n5376), .Z(n5374) );
  OR U5734 ( .A(n5377), .B(n5378), .Z(n5376) );
  NAND U5735 ( .A(n5378), .B(n5377), .Z(n5373) );
  XOR U5736 ( .A(n421), .B(n420), .Z(\A1[823] ) );
  XOR U5737 ( .A(n5378), .B(n5379), .Z(n420) );
  XNOR U5738 ( .A(n5377), .B(n5375), .Z(n5379) );
  AND U5739 ( .A(n5380), .B(n5381), .Z(n5375) );
  NANDN U5740 ( .A(n5382), .B(n5383), .Z(n5381) );
  NANDN U5741 ( .A(n5384), .B(n5385), .Z(n5383) );
  AND U5742 ( .A(B[822]), .B(A[3]), .Z(n5377) );
  XNOR U5743 ( .A(n5367), .B(n5386), .Z(n5378) );
  XNOR U5744 ( .A(n5365), .B(n5368), .Z(n5386) );
  NAND U5745 ( .A(A[2]), .B(B[823]), .Z(n5368) );
  NANDN U5746 ( .A(n5387), .B(n5388), .Z(n5365) );
  AND U5747 ( .A(A[0]), .B(B[824]), .Z(n5388) );
  XOR U5748 ( .A(n5370), .B(n5389), .Z(n5367) );
  NAND U5749 ( .A(A[0]), .B(B[825]), .Z(n5389) );
  NAND U5750 ( .A(B[824]), .B(A[1]), .Z(n5370) );
  NAND U5751 ( .A(n5390), .B(n5391), .Z(n421) );
  NANDN U5752 ( .A(n5392), .B(n5393), .Z(n5391) );
  OR U5753 ( .A(n5394), .B(n5395), .Z(n5393) );
  NAND U5754 ( .A(n5395), .B(n5394), .Z(n5390) );
  XOR U5755 ( .A(n423), .B(n422), .Z(\A1[822] ) );
  XOR U5756 ( .A(n5395), .B(n5396), .Z(n422) );
  XNOR U5757 ( .A(n5394), .B(n5392), .Z(n5396) );
  AND U5758 ( .A(n5397), .B(n5398), .Z(n5392) );
  NANDN U5759 ( .A(n5399), .B(n5400), .Z(n5398) );
  NANDN U5760 ( .A(n5401), .B(n5402), .Z(n5400) );
  AND U5761 ( .A(B[821]), .B(A[3]), .Z(n5394) );
  XNOR U5762 ( .A(n5384), .B(n5403), .Z(n5395) );
  XNOR U5763 ( .A(n5382), .B(n5385), .Z(n5403) );
  NAND U5764 ( .A(A[2]), .B(B[822]), .Z(n5385) );
  NANDN U5765 ( .A(n5404), .B(n5405), .Z(n5382) );
  AND U5766 ( .A(A[0]), .B(B[823]), .Z(n5405) );
  XOR U5767 ( .A(n5387), .B(n5406), .Z(n5384) );
  NAND U5768 ( .A(A[0]), .B(B[824]), .Z(n5406) );
  NAND U5769 ( .A(B[823]), .B(A[1]), .Z(n5387) );
  NAND U5770 ( .A(n5407), .B(n5408), .Z(n423) );
  NANDN U5771 ( .A(n5409), .B(n5410), .Z(n5408) );
  OR U5772 ( .A(n5411), .B(n5412), .Z(n5410) );
  NAND U5773 ( .A(n5412), .B(n5411), .Z(n5407) );
  XOR U5774 ( .A(n425), .B(n424), .Z(\A1[821] ) );
  XOR U5775 ( .A(n5412), .B(n5413), .Z(n424) );
  XNOR U5776 ( .A(n5411), .B(n5409), .Z(n5413) );
  AND U5777 ( .A(n5414), .B(n5415), .Z(n5409) );
  NANDN U5778 ( .A(n5416), .B(n5417), .Z(n5415) );
  NANDN U5779 ( .A(n5418), .B(n5419), .Z(n5417) );
  AND U5780 ( .A(B[820]), .B(A[3]), .Z(n5411) );
  XNOR U5781 ( .A(n5401), .B(n5420), .Z(n5412) );
  XNOR U5782 ( .A(n5399), .B(n5402), .Z(n5420) );
  NAND U5783 ( .A(A[2]), .B(B[821]), .Z(n5402) );
  NANDN U5784 ( .A(n5421), .B(n5422), .Z(n5399) );
  AND U5785 ( .A(A[0]), .B(B[822]), .Z(n5422) );
  XOR U5786 ( .A(n5404), .B(n5423), .Z(n5401) );
  NAND U5787 ( .A(A[0]), .B(B[823]), .Z(n5423) );
  NAND U5788 ( .A(B[822]), .B(A[1]), .Z(n5404) );
  NAND U5789 ( .A(n5424), .B(n5425), .Z(n425) );
  NANDN U5790 ( .A(n5426), .B(n5427), .Z(n5425) );
  OR U5791 ( .A(n5428), .B(n5429), .Z(n5427) );
  NAND U5792 ( .A(n5429), .B(n5428), .Z(n5424) );
  XOR U5793 ( .A(n427), .B(n426), .Z(\A1[820] ) );
  XOR U5794 ( .A(n5429), .B(n5430), .Z(n426) );
  XNOR U5795 ( .A(n5428), .B(n5426), .Z(n5430) );
  AND U5796 ( .A(n5431), .B(n5432), .Z(n5426) );
  NANDN U5797 ( .A(n5433), .B(n5434), .Z(n5432) );
  NANDN U5798 ( .A(n5435), .B(n5436), .Z(n5434) );
  AND U5799 ( .A(B[819]), .B(A[3]), .Z(n5428) );
  XNOR U5800 ( .A(n5418), .B(n5437), .Z(n5429) );
  XNOR U5801 ( .A(n5416), .B(n5419), .Z(n5437) );
  NAND U5802 ( .A(A[2]), .B(B[820]), .Z(n5419) );
  NANDN U5803 ( .A(n5438), .B(n5439), .Z(n5416) );
  AND U5804 ( .A(A[0]), .B(B[821]), .Z(n5439) );
  XOR U5805 ( .A(n5421), .B(n5440), .Z(n5418) );
  NAND U5806 ( .A(A[0]), .B(B[822]), .Z(n5440) );
  NAND U5807 ( .A(B[821]), .B(A[1]), .Z(n5421) );
  NAND U5808 ( .A(n5441), .B(n5442), .Z(n427) );
  NANDN U5809 ( .A(n5443), .B(n5444), .Z(n5442) );
  OR U5810 ( .A(n5445), .B(n5446), .Z(n5444) );
  NAND U5811 ( .A(n5446), .B(n5445), .Z(n5441) );
  XOR U5812 ( .A(n409), .B(n408), .Z(\A1[81] ) );
  XOR U5813 ( .A(n5276), .B(n5447), .Z(n408) );
  XNOR U5814 ( .A(n5275), .B(n5273), .Z(n5447) );
  AND U5815 ( .A(n5448), .B(n5449), .Z(n5273) );
  NANDN U5816 ( .A(n5450), .B(n5451), .Z(n5449) );
  NANDN U5817 ( .A(n5452), .B(n5453), .Z(n5451) );
  AND U5818 ( .A(B[80]), .B(A[3]), .Z(n5275) );
  XNOR U5819 ( .A(n5265), .B(n5454), .Z(n5276) );
  XNOR U5820 ( .A(n5263), .B(n5266), .Z(n5454) );
  NAND U5821 ( .A(A[2]), .B(B[81]), .Z(n5266) );
  NANDN U5822 ( .A(n5455), .B(n5456), .Z(n5263) );
  AND U5823 ( .A(A[0]), .B(B[82]), .Z(n5456) );
  XOR U5824 ( .A(n5268), .B(n5457), .Z(n5265) );
  NAND U5825 ( .A(A[0]), .B(B[83]), .Z(n5457) );
  NAND U5826 ( .A(B[82]), .B(A[1]), .Z(n5268) );
  NAND U5827 ( .A(n5458), .B(n5459), .Z(n409) );
  NANDN U5828 ( .A(n5460), .B(n5461), .Z(n5459) );
  OR U5829 ( .A(n5462), .B(n5463), .Z(n5461) );
  NAND U5830 ( .A(n5463), .B(n5462), .Z(n5458) );
  XOR U5831 ( .A(n429), .B(n428), .Z(\A1[819] ) );
  XOR U5832 ( .A(n5446), .B(n5464), .Z(n428) );
  XNOR U5833 ( .A(n5445), .B(n5443), .Z(n5464) );
  AND U5834 ( .A(n5465), .B(n5466), .Z(n5443) );
  NANDN U5835 ( .A(n5467), .B(n5468), .Z(n5466) );
  NANDN U5836 ( .A(n5469), .B(n5470), .Z(n5468) );
  AND U5837 ( .A(B[818]), .B(A[3]), .Z(n5445) );
  XNOR U5838 ( .A(n5435), .B(n5471), .Z(n5446) );
  XNOR U5839 ( .A(n5433), .B(n5436), .Z(n5471) );
  NAND U5840 ( .A(A[2]), .B(B[819]), .Z(n5436) );
  NANDN U5841 ( .A(n5472), .B(n5473), .Z(n5433) );
  AND U5842 ( .A(A[0]), .B(B[820]), .Z(n5473) );
  XOR U5843 ( .A(n5438), .B(n5474), .Z(n5435) );
  NAND U5844 ( .A(A[0]), .B(B[821]), .Z(n5474) );
  NAND U5845 ( .A(B[820]), .B(A[1]), .Z(n5438) );
  NAND U5846 ( .A(n5475), .B(n5476), .Z(n429) );
  NANDN U5847 ( .A(n5477), .B(n5478), .Z(n5476) );
  OR U5848 ( .A(n5479), .B(n5480), .Z(n5478) );
  NAND U5849 ( .A(n5480), .B(n5479), .Z(n5475) );
  XOR U5850 ( .A(n433), .B(n432), .Z(\A1[818] ) );
  XOR U5851 ( .A(n5480), .B(n5481), .Z(n432) );
  XNOR U5852 ( .A(n5479), .B(n5477), .Z(n5481) );
  AND U5853 ( .A(n5482), .B(n5483), .Z(n5477) );
  NANDN U5854 ( .A(n5484), .B(n5485), .Z(n5483) );
  NANDN U5855 ( .A(n5486), .B(n5487), .Z(n5485) );
  AND U5856 ( .A(B[817]), .B(A[3]), .Z(n5479) );
  XNOR U5857 ( .A(n5469), .B(n5488), .Z(n5480) );
  XNOR U5858 ( .A(n5467), .B(n5470), .Z(n5488) );
  NAND U5859 ( .A(A[2]), .B(B[818]), .Z(n5470) );
  NANDN U5860 ( .A(n5489), .B(n5490), .Z(n5467) );
  AND U5861 ( .A(A[0]), .B(B[819]), .Z(n5490) );
  XOR U5862 ( .A(n5472), .B(n5491), .Z(n5469) );
  NAND U5863 ( .A(A[0]), .B(B[820]), .Z(n5491) );
  NAND U5864 ( .A(B[819]), .B(A[1]), .Z(n5472) );
  NAND U5865 ( .A(n5492), .B(n5493), .Z(n433) );
  NANDN U5866 ( .A(n5494), .B(n5495), .Z(n5493) );
  OR U5867 ( .A(n5496), .B(n5497), .Z(n5495) );
  NAND U5868 ( .A(n5497), .B(n5496), .Z(n5492) );
  XOR U5869 ( .A(n435), .B(n434), .Z(\A1[817] ) );
  XOR U5870 ( .A(n5497), .B(n5498), .Z(n434) );
  XNOR U5871 ( .A(n5496), .B(n5494), .Z(n5498) );
  AND U5872 ( .A(n5499), .B(n5500), .Z(n5494) );
  NANDN U5873 ( .A(n5501), .B(n5502), .Z(n5500) );
  NANDN U5874 ( .A(n5503), .B(n5504), .Z(n5502) );
  AND U5875 ( .A(B[816]), .B(A[3]), .Z(n5496) );
  XNOR U5876 ( .A(n5486), .B(n5505), .Z(n5497) );
  XNOR U5877 ( .A(n5484), .B(n5487), .Z(n5505) );
  NAND U5878 ( .A(A[2]), .B(B[817]), .Z(n5487) );
  NANDN U5879 ( .A(n5506), .B(n5507), .Z(n5484) );
  AND U5880 ( .A(A[0]), .B(B[818]), .Z(n5507) );
  XOR U5881 ( .A(n5489), .B(n5508), .Z(n5486) );
  NAND U5882 ( .A(A[0]), .B(B[819]), .Z(n5508) );
  NAND U5883 ( .A(B[818]), .B(A[1]), .Z(n5489) );
  NAND U5884 ( .A(n5509), .B(n5510), .Z(n435) );
  NANDN U5885 ( .A(n5511), .B(n5512), .Z(n5510) );
  OR U5886 ( .A(n5513), .B(n5514), .Z(n5512) );
  NAND U5887 ( .A(n5514), .B(n5513), .Z(n5509) );
  XOR U5888 ( .A(n437), .B(n436), .Z(\A1[816] ) );
  XOR U5889 ( .A(n5514), .B(n5515), .Z(n436) );
  XNOR U5890 ( .A(n5513), .B(n5511), .Z(n5515) );
  AND U5891 ( .A(n5516), .B(n5517), .Z(n5511) );
  NANDN U5892 ( .A(n5518), .B(n5519), .Z(n5517) );
  NANDN U5893 ( .A(n5520), .B(n5521), .Z(n5519) );
  AND U5894 ( .A(B[815]), .B(A[3]), .Z(n5513) );
  XNOR U5895 ( .A(n5503), .B(n5522), .Z(n5514) );
  XNOR U5896 ( .A(n5501), .B(n5504), .Z(n5522) );
  NAND U5897 ( .A(A[2]), .B(B[816]), .Z(n5504) );
  NANDN U5898 ( .A(n5523), .B(n5524), .Z(n5501) );
  AND U5899 ( .A(A[0]), .B(B[817]), .Z(n5524) );
  XOR U5900 ( .A(n5506), .B(n5525), .Z(n5503) );
  NAND U5901 ( .A(A[0]), .B(B[818]), .Z(n5525) );
  NAND U5902 ( .A(B[817]), .B(A[1]), .Z(n5506) );
  NAND U5903 ( .A(n5526), .B(n5527), .Z(n437) );
  NANDN U5904 ( .A(n5528), .B(n5529), .Z(n5527) );
  OR U5905 ( .A(n5530), .B(n5531), .Z(n5529) );
  NAND U5906 ( .A(n5531), .B(n5530), .Z(n5526) );
  XOR U5907 ( .A(n439), .B(n438), .Z(\A1[815] ) );
  XOR U5908 ( .A(n5531), .B(n5532), .Z(n438) );
  XNOR U5909 ( .A(n5530), .B(n5528), .Z(n5532) );
  AND U5910 ( .A(n5533), .B(n5534), .Z(n5528) );
  NANDN U5911 ( .A(n5535), .B(n5536), .Z(n5534) );
  NANDN U5912 ( .A(n5537), .B(n5538), .Z(n5536) );
  AND U5913 ( .A(B[814]), .B(A[3]), .Z(n5530) );
  XNOR U5914 ( .A(n5520), .B(n5539), .Z(n5531) );
  XNOR U5915 ( .A(n5518), .B(n5521), .Z(n5539) );
  NAND U5916 ( .A(A[2]), .B(B[815]), .Z(n5521) );
  NANDN U5917 ( .A(n5540), .B(n5541), .Z(n5518) );
  AND U5918 ( .A(A[0]), .B(B[816]), .Z(n5541) );
  XOR U5919 ( .A(n5523), .B(n5542), .Z(n5520) );
  NAND U5920 ( .A(A[0]), .B(B[817]), .Z(n5542) );
  NAND U5921 ( .A(B[816]), .B(A[1]), .Z(n5523) );
  NAND U5922 ( .A(n5543), .B(n5544), .Z(n439) );
  NANDN U5923 ( .A(n5545), .B(n5546), .Z(n5544) );
  OR U5924 ( .A(n5547), .B(n5548), .Z(n5546) );
  NAND U5925 ( .A(n5548), .B(n5547), .Z(n5543) );
  XOR U5926 ( .A(n441), .B(n440), .Z(\A1[814] ) );
  XOR U5927 ( .A(n5548), .B(n5549), .Z(n440) );
  XNOR U5928 ( .A(n5547), .B(n5545), .Z(n5549) );
  AND U5929 ( .A(n5550), .B(n5551), .Z(n5545) );
  NANDN U5930 ( .A(n5552), .B(n5553), .Z(n5551) );
  NANDN U5931 ( .A(n5554), .B(n5555), .Z(n5553) );
  AND U5932 ( .A(B[813]), .B(A[3]), .Z(n5547) );
  XNOR U5933 ( .A(n5537), .B(n5556), .Z(n5548) );
  XNOR U5934 ( .A(n5535), .B(n5538), .Z(n5556) );
  NAND U5935 ( .A(A[2]), .B(B[814]), .Z(n5538) );
  NANDN U5936 ( .A(n5557), .B(n5558), .Z(n5535) );
  AND U5937 ( .A(A[0]), .B(B[815]), .Z(n5558) );
  XOR U5938 ( .A(n5540), .B(n5559), .Z(n5537) );
  NAND U5939 ( .A(A[0]), .B(B[816]), .Z(n5559) );
  NAND U5940 ( .A(B[815]), .B(A[1]), .Z(n5540) );
  NAND U5941 ( .A(n5560), .B(n5561), .Z(n441) );
  NANDN U5942 ( .A(n5562), .B(n5563), .Z(n5561) );
  OR U5943 ( .A(n5564), .B(n5565), .Z(n5563) );
  NAND U5944 ( .A(n5565), .B(n5564), .Z(n5560) );
  XOR U5945 ( .A(n443), .B(n442), .Z(\A1[813] ) );
  XOR U5946 ( .A(n5565), .B(n5566), .Z(n442) );
  XNOR U5947 ( .A(n5564), .B(n5562), .Z(n5566) );
  AND U5948 ( .A(n5567), .B(n5568), .Z(n5562) );
  NANDN U5949 ( .A(n5569), .B(n5570), .Z(n5568) );
  NANDN U5950 ( .A(n5571), .B(n5572), .Z(n5570) );
  AND U5951 ( .A(B[812]), .B(A[3]), .Z(n5564) );
  XNOR U5952 ( .A(n5554), .B(n5573), .Z(n5565) );
  XNOR U5953 ( .A(n5552), .B(n5555), .Z(n5573) );
  NAND U5954 ( .A(A[2]), .B(B[813]), .Z(n5555) );
  NANDN U5955 ( .A(n5574), .B(n5575), .Z(n5552) );
  AND U5956 ( .A(A[0]), .B(B[814]), .Z(n5575) );
  XOR U5957 ( .A(n5557), .B(n5576), .Z(n5554) );
  NAND U5958 ( .A(A[0]), .B(B[815]), .Z(n5576) );
  NAND U5959 ( .A(B[814]), .B(A[1]), .Z(n5557) );
  NAND U5960 ( .A(n5577), .B(n5578), .Z(n443) );
  NANDN U5961 ( .A(n5579), .B(n5580), .Z(n5578) );
  OR U5962 ( .A(n5581), .B(n5582), .Z(n5580) );
  NAND U5963 ( .A(n5582), .B(n5581), .Z(n5577) );
  XOR U5964 ( .A(n445), .B(n444), .Z(\A1[812] ) );
  XOR U5965 ( .A(n5582), .B(n5583), .Z(n444) );
  XNOR U5966 ( .A(n5581), .B(n5579), .Z(n5583) );
  AND U5967 ( .A(n5584), .B(n5585), .Z(n5579) );
  NANDN U5968 ( .A(n5586), .B(n5587), .Z(n5585) );
  NANDN U5969 ( .A(n5588), .B(n5589), .Z(n5587) );
  AND U5970 ( .A(B[811]), .B(A[3]), .Z(n5581) );
  XNOR U5971 ( .A(n5571), .B(n5590), .Z(n5582) );
  XNOR U5972 ( .A(n5569), .B(n5572), .Z(n5590) );
  NAND U5973 ( .A(A[2]), .B(B[812]), .Z(n5572) );
  NANDN U5974 ( .A(n5591), .B(n5592), .Z(n5569) );
  AND U5975 ( .A(A[0]), .B(B[813]), .Z(n5592) );
  XOR U5976 ( .A(n5574), .B(n5593), .Z(n5571) );
  NAND U5977 ( .A(A[0]), .B(B[814]), .Z(n5593) );
  NAND U5978 ( .A(B[813]), .B(A[1]), .Z(n5574) );
  NAND U5979 ( .A(n5594), .B(n5595), .Z(n445) );
  NANDN U5980 ( .A(n5596), .B(n5597), .Z(n5595) );
  OR U5981 ( .A(n5598), .B(n5599), .Z(n5597) );
  NAND U5982 ( .A(n5599), .B(n5598), .Z(n5594) );
  XOR U5983 ( .A(n447), .B(n446), .Z(\A1[811] ) );
  XOR U5984 ( .A(n5599), .B(n5600), .Z(n446) );
  XNOR U5985 ( .A(n5598), .B(n5596), .Z(n5600) );
  AND U5986 ( .A(n5601), .B(n5602), .Z(n5596) );
  NANDN U5987 ( .A(n5603), .B(n5604), .Z(n5602) );
  NANDN U5988 ( .A(n5605), .B(n5606), .Z(n5604) );
  AND U5989 ( .A(B[810]), .B(A[3]), .Z(n5598) );
  XNOR U5990 ( .A(n5588), .B(n5607), .Z(n5599) );
  XNOR U5991 ( .A(n5586), .B(n5589), .Z(n5607) );
  NAND U5992 ( .A(A[2]), .B(B[811]), .Z(n5589) );
  NANDN U5993 ( .A(n5608), .B(n5609), .Z(n5586) );
  AND U5994 ( .A(A[0]), .B(B[812]), .Z(n5609) );
  XOR U5995 ( .A(n5591), .B(n5610), .Z(n5588) );
  NAND U5996 ( .A(A[0]), .B(B[813]), .Z(n5610) );
  NAND U5997 ( .A(B[812]), .B(A[1]), .Z(n5591) );
  NAND U5998 ( .A(n5611), .B(n5612), .Z(n447) );
  NANDN U5999 ( .A(n5613), .B(n5614), .Z(n5612) );
  OR U6000 ( .A(n5615), .B(n5616), .Z(n5614) );
  NAND U6001 ( .A(n5616), .B(n5615), .Z(n5611) );
  XOR U6002 ( .A(n449), .B(n448), .Z(\A1[810] ) );
  XOR U6003 ( .A(n5616), .B(n5617), .Z(n448) );
  XNOR U6004 ( .A(n5615), .B(n5613), .Z(n5617) );
  AND U6005 ( .A(n5618), .B(n5619), .Z(n5613) );
  NANDN U6006 ( .A(n5620), .B(n5621), .Z(n5619) );
  NANDN U6007 ( .A(n5622), .B(n5623), .Z(n5621) );
  AND U6008 ( .A(B[809]), .B(A[3]), .Z(n5615) );
  XNOR U6009 ( .A(n5605), .B(n5624), .Z(n5616) );
  XNOR U6010 ( .A(n5603), .B(n5606), .Z(n5624) );
  NAND U6011 ( .A(A[2]), .B(B[810]), .Z(n5606) );
  NANDN U6012 ( .A(n5625), .B(n5626), .Z(n5603) );
  AND U6013 ( .A(A[0]), .B(B[811]), .Z(n5626) );
  XOR U6014 ( .A(n5608), .B(n5627), .Z(n5605) );
  NAND U6015 ( .A(A[0]), .B(B[812]), .Z(n5627) );
  NAND U6016 ( .A(B[811]), .B(A[1]), .Z(n5608) );
  NAND U6017 ( .A(n5628), .B(n5629), .Z(n449) );
  NANDN U6018 ( .A(n5630), .B(n5631), .Z(n5629) );
  OR U6019 ( .A(n5632), .B(n5633), .Z(n5631) );
  NAND U6020 ( .A(n5633), .B(n5632), .Z(n5628) );
  XOR U6021 ( .A(n431), .B(n430), .Z(\A1[80] ) );
  XOR U6022 ( .A(n5463), .B(n5634), .Z(n430) );
  XNOR U6023 ( .A(n5462), .B(n5460), .Z(n5634) );
  AND U6024 ( .A(n5635), .B(n5636), .Z(n5460) );
  NANDN U6025 ( .A(n5637), .B(n5638), .Z(n5636) );
  NANDN U6026 ( .A(n5639), .B(n5640), .Z(n5638) );
  AND U6027 ( .A(B[79]), .B(A[3]), .Z(n5462) );
  XNOR U6028 ( .A(n5452), .B(n5641), .Z(n5463) );
  XNOR U6029 ( .A(n5450), .B(n5453), .Z(n5641) );
  NAND U6030 ( .A(A[2]), .B(B[80]), .Z(n5453) );
  NANDN U6031 ( .A(n5642), .B(n5643), .Z(n5450) );
  AND U6032 ( .A(A[0]), .B(B[81]), .Z(n5643) );
  XOR U6033 ( .A(n5455), .B(n5644), .Z(n5452) );
  NAND U6034 ( .A(A[0]), .B(B[82]), .Z(n5644) );
  NAND U6035 ( .A(B[81]), .B(A[1]), .Z(n5455) );
  NAND U6036 ( .A(n5645), .B(n5646), .Z(n431) );
  NANDN U6037 ( .A(n5647), .B(n5648), .Z(n5646) );
  OR U6038 ( .A(n5649), .B(n5650), .Z(n5648) );
  NAND U6039 ( .A(n5650), .B(n5649), .Z(n5645) );
  XOR U6040 ( .A(n451), .B(n450), .Z(\A1[809] ) );
  XOR U6041 ( .A(n5633), .B(n5651), .Z(n450) );
  XNOR U6042 ( .A(n5632), .B(n5630), .Z(n5651) );
  AND U6043 ( .A(n5652), .B(n5653), .Z(n5630) );
  NANDN U6044 ( .A(n5654), .B(n5655), .Z(n5653) );
  NANDN U6045 ( .A(n5656), .B(n5657), .Z(n5655) );
  AND U6046 ( .A(B[808]), .B(A[3]), .Z(n5632) );
  XNOR U6047 ( .A(n5622), .B(n5658), .Z(n5633) );
  XNOR U6048 ( .A(n5620), .B(n5623), .Z(n5658) );
  NAND U6049 ( .A(A[2]), .B(B[809]), .Z(n5623) );
  NANDN U6050 ( .A(n5659), .B(n5660), .Z(n5620) );
  AND U6051 ( .A(A[0]), .B(B[810]), .Z(n5660) );
  XOR U6052 ( .A(n5625), .B(n5661), .Z(n5622) );
  NAND U6053 ( .A(A[0]), .B(B[811]), .Z(n5661) );
  NAND U6054 ( .A(B[810]), .B(A[1]), .Z(n5625) );
  NAND U6055 ( .A(n5662), .B(n5663), .Z(n451) );
  NANDN U6056 ( .A(n5664), .B(n5665), .Z(n5663) );
  OR U6057 ( .A(n5666), .B(n5667), .Z(n5665) );
  NAND U6058 ( .A(n5667), .B(n5666), .Z(n5662) );
  XOR U6059 ( .A(n455), .B(n454), .Z(\A1[808] ) );
  XOR U6060 ( .A(n5667), .B(n5668), .Z(n454) );
  XNOR U6061 ( .A(n5666), .B(n5664), .Z(n5668) );
  AND U6062 ( .A(n5669), .B(n5670), .Z(n5664) );
  NANDN U6063 ( .A(n5671), .B(n5672), .Z(n5670) );
  NANDN U6064 ( .A(n5673), .B(n5674), .Z(n5672) );
  AND U6065 ( .A(B[807]), .B(A[3]), .Z(n5666) );
  XNOR U6066 ( .A(n5656), .B(n5675), .Z(n5667) );
  XNOR U6067 ( .A(n5654), .B(n5657), .Z(n5675) );
  NAND U6068 ( .A(A[2]), .B(B[808]), .Z(n5657) );
  NANDN U6069 ( .A(n5676), .B(n5677), .Z(n5654) );
  AND U6070 ( .A(A[0]), .B(B[809]), .Z(n5677) );
  XOR U6071 ( .A(n5659), .B(n5678), .Z(n5656) );
  NAND U6072 ( .A(A[0]), .B(B[810]), .Z(n5678) );
  NAND U6073 ( .A(B[809]), .B(A[1]), .Z(n5659) );
  NAND U6074 ( .A(n5679), .B(n5680), .Z(n455) );
  NANDN U6075 ( .A(n5681), .B(n5682), .Z(n5680) );
  OR U6076 ( .A(n5683), .B(n5684), .Z(n5682) );
  NAND U6077 ( .A(n5684), .B(n5683), .Z(n5679) );
  XOR U6078 ( .A(n457), .B(n456), .Z(\A1[807] ) );
  XOR U6079 ( .A(n5684), .B(n5685), .Z(n456) );
  XNOR U6080 ( .A(n5683), .B(n5681), .Z(n5685) );
  AND U6081 ( .A(n5686), .B(n5687), .Z(n5681) );
  NANDN U6082 ( .A(n5688), .B(n5689), .Z(n5687) );
  NANDN U6083 ( .A(n5690), .B(n5691), .Z(n5689) );
  AND U6084 ( .A(B[806]), .B(A[3]), .Z(n5683) );
  XNOR U6085 ( .A(n5673), .B(n5692), .Z(n5684) );
  XNOR U6086 ( .A(n5671), .B(n5674), .Z(n5692) );
  NAND U6087 ( .A(A[2]), .B(B[807]), .Z(n5674) );
  NANDN U6088 ( .A(n5693), .B(n5694), .Z(n5671) );
  AND U6089 ( .A(A[0]), .B(B[808]), .Z(n5694) );
  XOR U6090 ( .A(n5676), .B(n5695), .Z(n5673) );
  NAND U6091 ( .A(A[0]), .B(B[809]), .Z(n5695) );
  NAND U6092 ( .A(B[808]), .B(A[1]), .Z(n5676) );
  NAND U6093 ( .A(n5696), .B(n5697), .Z(n457) );
  NANDN U6094 ( .A(n5698), .B(n5699), .Z(n5697) );
  OR U6095 ( .A(n5700), .B(n5701), .Z(n5699) );
  NAND U6096 ( .A(n5701), .B(n5700), .Z(n5696) );
  XOR U6097 ( .A(n459), .B(n458), .Z(\A1[806] ) );
  XOR U6098 ( .A(n5701), .B(n5702), .Z(n458) );
  XNOR U6099 ( .A(n5700), .B(n5698), .Z(n5702) );
  AND U6100 ( .A(n5703), .B(n5704), .Z(n5698) );
  NANDN U6101 ( .A(n5705), .B(n5706), .Z(n5704) );
  NANDN U6102 ( .A(n5707), .B(n5708), .Z(n5706) );
  AND U6103 ( .A(B[805]), .B(A[3]), .Z(n5700) );
  XNOR U6104 ( .A(n5690), .B(n5709), .Z(n5701) );
  XNOR U6105 ( .A(n5688), .B(n5691), .Z(n5709) );
  NAND U6106 ( .A(A[2]), .B(B[806]), .Z(n5691) );
  NANDN U6107 ( .A(n5710), .B(n5711), .Z(n5688) );
  AND U6108 ( .A(A[0]), .B(B[807]), .Z(n5711) );
  XOR U6109 ( .A(n5693), .B(n5712), .Z(n5690) );
  NAND U6110 ( .A(A[0]), .B(B[808]), .Z(n5712) );
  NAND U6111 ( .A(B[807]), .B(A[1]), .Z(n5693) );
  NAND U6112 ( .A(n5713), .B(n5714), .Z(n459) );
  NANDN U6113 ( .A(n5715), .B(n5716), .Z(n5714) );
  OR U6114 ( .A(n5717), .B(n5718), .Z(n5716) );
  NAND U6115 ( .A(n5718), .B(n5717), .Z(n5713) );
  XOR U6116 ( .A(n461), .B(n460), .Z(\A1[805] ) );
  XOR U6117 ( .A(n5718), .B(n5719), .Z(n460) );
  XNOR U6118 ( .A(n5717), .B(n5715), .Z(n5719) );
  AND U6119 ( .A(n5720), .B(n5721), .Z(n5715) );
  NANDN U6120 ( .A(n5722), .B(n5723), .Z(n5721) );
  NANDN U6121 ( .A(n5724), .B(n5725), .Z(n5723) );
  AND U6122 ( .A(B[804]), .B(A[3]), .Z(n5717) );
  XNOR U6123 ( .A(n5707), .B(n5726), .Z(n5718) );
  XNOR U6124 ( .A(n5705), .B(n5708), .Z(n5726) );
  NAND U6125 ( .A(A[2]), .B(B[805]), .Z(n5708) );
  NANDN U6126 ( .A(n5727), .B(n5728), .Z(n5705) );
  AND U6127 ( .A(A[0]), .B(B[806]), .Z(n5728) );
  XOR U6128 ( .A(n5710), .B(n5729), .Z(n5707) );
  NAND U6129 ( .A(A[0]), .B(B[807]), .Z(n5729) );
  NAND U6130 ( .A(B[806]), .B(A[1]), .Z(n5710) );
  NAND U6131 ( .A(n5730), .B(n5731), .Z(n461) );
  NANDN U6132 ( .A(n5732), .B(n5733), .Z(n5731) );
  OR U6133 ( .A(n5734), .B(n5735), .Z(n5733) );
  NAND U6134 ( .A(n5735), .B(n5734), .Z(n5730) );
  XOR U6135 ( .A(n463), .B(n462), .Z(\A1[804] ) );
  XOR U6136 ( .A(n5735), .B(n5736), .Z(n462) );
  XNOR U6137 ( .A(n5734), .B(n5732), .Z(n5736) );
  AND U6138 ( .A(n5737), .B(n5738), .Z(n5732) );
  NANDN U6139 ( .A(n5739), .B(n5740), .Z(n5738) );
  NANDN U6140 ( .A(n5741), .B(n5742), .Z(n5740) );
  AND U6141 ( .A(B[803]), .B(A[3]), .Z(n5734) );
  XNOR U6142 ( .A(n5724), .B(n5743), .Z(n5735) );
  XNOR U6143 ( .A(n5722), .B(n5725), .Z(n5743) );
  NAND U6144 ( .A(A[2]), .B(B[804]), .Z(n5725) );
  NANDN U6145 ( .A(n5744), .B(n5745), .Z(n5722) );
  AND U6146 ( .A(A[0]), .B(B[805]), .Z(n5745) );
  XOR U6147 ( .A(n5727), .B(n5746), .Z(n5724) );
  NAND U6148 ( .A(A[0]), .B(B[806]), .Z(n5746) );
  NAND U6149 ( .A(B[805]), .B(A[1]), .Z(n5727) );
  NAND U6150 ( .A(n5747), .B(n5748), .Z(n463) );
  NANDN U6151 ( .A(n5749), .B(n5750), .Z(n5748) );
  OR U6152 ( .A(n5751), .B(n5752), .Z(n5750) );
  NAND U6153 ( .A(n5752), .B(n5751), .Z(n5747) );
  XOR U6154 ( .A(n465), .B(n464), .Z(\A1[803] ) );
  XOR U6155 ( .A(n5752), .B(n5753), .Z(n464) );
  XNOR U6156 ( .A(n5751), .B(n5749), .Z(n5753) );
  AND U6157 ( .A(n5754), .B(n5755), .Z(n5749) );
  NANDN U6158 ( .A(n5756), .B(n5757), .Z(n5755) );
  NANDN U6159 ( .A(n5758), .B(n5759), .Z(n5757) );
  AND U6160 ( .A(B[802]), .B(A[3]), .Z(n5751) );
  XNOR U6161 ( .A(n5741), .B(n5760), .Z(n5752) );
  XNOR U6162 ( .A(n5739), .B(n5742), .Z(n5760) );
  NAND U6163 ( .A(A[2]), .B(B[803]), .Z(n5742) );
  NANDN U6164 ( .A(n5761), .B(n5762), .Z(n5739) );
  AND U6165 ( .A(A[0]), .B(B[804]), .Z(n5762) );
  XOR U6166 ( .A(n5744), .B(n5763), .Z(n5741) );
  NAND U6167 ( .A(A[0]), .B(B[805]), .Z(n5763) );
  NAND U6168 ( .A(B[804]), .B(A[1]), .Z(n5744) );
  NAND U6169 ( .A(n5764), .B(n5765), .Z(n465) );
  NANDN U6170 ( .A(n5766), .B(n5767), .Z(n5765) );
  OR U6171 ( .A(n5768), .B(n5769), .Z(n5767) );
  NAND U6172 ( .A(n5769), .B(n5768), .Z(n5764) );
  XOR U6173 ( .A(n467), .B(n466), .Z(\A1[802] ) );
  XOR U6174 ( .A(n5769), .B(n5770), .Z(n466) );
  XNOR U6175 ( .A(n5768), .B(n5766), .Z(n5770) );
  AND U6176 ( .A(n5771), .B(n5772), .Z(n5766) );
  NANDN U6177 ( .A(n5773), .B(n5774), .Z(n5772) );
  NANDN U6178 ( .A(n5775), .B(n5776), .Z(n5774) );
  AND U6179 ( .A(B[801]), .B(A[3]), .Z(n5768) );
  XNOR U6180 ( .A(n5758), .B(n5777), .Z(n5769) );
  XNOR U6181 ( .A(n5756), .B(n5759), .Z(n5777) );
  NAND U6182 ( .A(A[2]), .B(B[802]), .Z(n5759) );
  NANDN U6183 ( .A(n5778), .B(n5779), .Z(n5756) );
  AND U6184 ( .A(A[0]), .B(B[803]), .Z(n5779) );
  XOR U6185 ( .A(n5761), .B(n5780), .Z(n5758) );
  NAND U6186 ( .A(A[0]), .B(B[804]), .Z(n5780) );
  NAND U6187 ( .A(B[803]), .B(A[1]), .Z(n5761) );
  NAND U6188 ( .A(n5781), .B(n5782), .Z(n467) );
  NANDN U6189 ( .A(n5783), .B(n5784), .Z(n5782) );
  OR U6190 ( .A(n5785), .B(n5786), .Z(n5784) );
  NAND U6191 ( .A(n5786), .B(n5785), .Z(n5781) );
  XOR U6192 ( .A(n469), .B(n468), .Z(\A1[801] ) );
  XOR U6193 ( .A(n5786), .B(n5787), .Z(n468) );
  XNOR U6194 ( .A(n5785), .B(n5783), .Z(n5787) );
  AND U6195 ( .A(n5788), .B(n5789), .Z(n5783) );
  NANDN U6196 ( .A(n5790), .B(n5791), .Z(n5789) );
  NANDN U6197 ( .A(n5792), .B(n5793), .Z(n5791) );
  AND U6198 ( .A(B[800]), .B(A[3]), .Z(n5785) );
  XNOR U6199 ( .A(n5775), .B(n5794), .Z(n5786) );
  XNOR U6200 ( .A(n5773), .B(n5776), .Z(n5794) );
  NAND U6201 ( .A(A[2]), .B(B[801]), .Z(n5776) );
  NANDN U6202 ( .A(n5795), .B(n5796), .Z(n5773) );
  AND U6203 ( .A(A[0]), .B(B[802]), .Z(n5796) );
  XOR U6204 ( .A(n5778), .B(n5797), .Z(n5775) );
  NAND U6205 ( .A(A[0]), .B(B[803]), .Z(n5797) );
  NAND U6206 ( .A(B[802]), .B(A[1]), .Z(n5778) );
  NAND U6207 ( .A(n5798), .B(n5799), .Z(n469) );
  NANDN U6208 ( .A(n5800), .B(n5801), .Z(n5799) );
  OR U6209 ( .A(n5802), .B(n5803), .Z(n5801) );
  NAND U6210 ( .A(n5803), .B(n5802), .Z(n5798) );
  XOR U6211 ( .A(n471), .B(n470), .Z(\A1[800] ) );
  XOR U6212 ( .A(n5803), .B(n5804), .Z(n470) );
  XNOR U6213 ( .A(n5802), .B(n5800), .Z(n5804) );
  AND U6214 ( .A(n5805), .B(n5806), .Z(n5800) );
  NANDN U6215 ( .A(n5807), .B(n5808), .Z(n5806) );
  NANDN U6216 ( .A(n5809), .B(n5810), .Z(n5808) );
  AND U6217 ( .A(B[799]), .B(A[3]), .Z(n5802) );
  XNOR U6218 ( .A(n5792), .B(n5811), .Z(n5803) );
  XNOR U6219 ( .A(n5790), .B(n5793), .Z(n5811) );
  NAND U6220 ( .A(A[2]), .B(B[800]), .Z(n5793) );
  NANDN U6221 ( .A(n5812), .B(n5813), .Z(n5790) );
  AND U6222 ( .A(A[0]), .B(B[801]), .Z(n5813) );
  XOR U6223 ( .A(n5795), .B(n5814), .Z(n5792) );
  NAND U6224 ( .A(A[0]), .B(B[802]), .Z(n5814) );
  NAND U6225 ( .A(B[801]), .B(A[1]), .Z(n5795) );
  NAND U6226 ( .A(n5815), .B(n5816), .Z(n471) );
  NANDN U6227 ( .A(n5817), .B(n5818), .Z(n5816) );
  OR U6228 ( .A(n5819), .B(n5820), .Z(n5818) );
  NAND U6229 ( .A(n5820), .B(n5819), .Z(n5815) );
  XOR U6230 ( .A(n253), .B(n252), .Z(\A1[7] ) );
  XNOR U6231 ( .A(n23), .B(n5821), .Z(n252) );
  XNOR U6232 ( .A(n3949), .B(n3947), .Z(n5821) );
  AND U6233 ( .A(n5822), .B(n5823), .Z(n3947) );
  NANDN U6234 ( .A(n5824), .B(n5825), .Z(n5823) );
  NANDN U6235 ( .A(n5826), .B(n5827), .Z(n5825) );
  AND U6236 ( .A(B[6]), .B(A[3]), .Z(n3949) );
  XOR U6237 ( .A(n3939), .B(n5828), .Z(n3950) );
  XOR U6238 ( .A(n3941), .B(n3942), .Z(n5828) );
  NAND U6239 ( .A(B[7]), .B(A[2]), .Z(n3942) );
  ANDN U6240 ( .B(n5829), .A(n5830), .Z(n3941) );
  AND U6241 ( .A(A[0]), .B(B[8]), .Z(n5829) );
  XNOR U6242 ( .A(n5831), .B(n5832), .Z(n3939) );
  NANDN U6243 ( .A(n24), .B(A[0]), .Z(n5832) );
  NAND U6244 ( .A(n5833), .B(n5834), .Z(n253) );
  NANDN U6245 ( .A(n5835), .B(n5836), .Z(n5834) );
  OR U6246 ( .A(n5837), .B(n5838), .Z(n5836) );
  NAND U6247 ( .A(n5838), .B(n5837), .Z(n5833) );
  XOR U6248 ( .A(n453), .B(n452), .Z(\A1[79] ) );
  XOR U6249 ( .A(n5650), .B(n5839), .Z(n452) );
  XNOR U6250 ( .A(n5649), .B(n5647), .Z(n5839) );
  AND U6251 ( .A(n5840), .B(n5841), .Z(n5647) );
  NANDN U6252 ( .A(n5842), .B(n5843), .Z(n5841) );
  NANDN U6253 ( .A(n5844), .B(n5845), .Z(n5843) );
  AND U6254 ( .A(B[78]), .B(A[3]), .Z(n5649) );
  XNOR U6255 ( .A(n5639), .B(n5846), .Z(n5650) );
  XNOR U6256 ( .A(n5637), .B(n5640), .Z(n5846) );
  NAND U6257 ( .A(A[2]), .B(B[79]), .Z(n5640) );
  NANDN U6258 ( .A(n5847), .B(n5848), .Z(n5637) );
  AND U6259 ( .A(A[0]), .B(B[80]), .Z(n5848) );
  XOR U6260 ( .A(n5642), .B(n5849), .Z(n5639) );
  NAND U6261 ( .A(A[0]), .B(B[81]), .Z(n5849) );
  NAND U6262 ( .A(B[80]), .B(A[1]), .Z(n5642) );
  NAND U6263 ( .A(n5850), .B(n5851), .Z(n453) );
  NANDN U6264 ( .A(n5852), .B(n5853), .Z(n5851) );
  OR U6265 ( .A(n5854), .B(n5855), .Z(n5853) );
  NAND U6266 ( .A(n5855), .B(n5854), .Z(n5850) );
  XOR U6267 ( .A(n473), .B(n472), .Z(\A1[799] ) );
  XOR U6268 ( .A(n5820), .B(n5856), .Z(n472) );
  XNOR U6269 ( .A(n5819), .B(n5817), .Z(n5856) );
  AND U6270 ( .A(n5857), .B(n5858), .Z(n5817) );
  NANDN U6271 ( .A(n5859), .B(n5860), .Z(n5858) );
  NANDN U6272 ( .A(n5861), .B(n5862), .Z(n5860) );
  AND U6273 ( .A(B[798]), .B(A[3]), .Z(n5819) );
  XNOR U6274 ( .A(n5809), .B(n5863), .Z(n5820) );
  XNOR U6275 ( .A(n5807), .B(n5810), .Z(n5863) );
  NAND U6276 ( .A(A[2]), .B(B[799]), .Z(n5810) );
  NANDN U6277 ( .A(n5864), .B(n5865), .Z(n5807) );
  AND U6278 ( .A(A[0]), .B(B[800]), .Z(n5865) );
  XOR U6279 ( .A(n5812), .B(n5866), .Z(n5809) );
  NAND U6280 ( .A(A[0]), .B(B[801]), .Z(n5866) );
  NAND U6281 ( .A(B[800]), .B(A[1]), .Z(n5812) );
  NAND U6282 ( .A(n5867), .B(n5868), .Z(n473) );
  NANDN U6283 ( .A(n5869), .B(n5870), .Z(n5868) );
  OR U6284 ( .A(n5871), .B(n5872), .Z(n5870) );
  NAND U6285 ( .A(n5872), .B(n5871), .Z(n5867) );
  XOR U6286 ( .A(n479), .B(n478), .Z(\A1[798] ) );
  XOR U6287 ( .A(n5872), .B(n5873), .Z(n478) );
  XNOR U6288 ( .A(n5871), .B(n5869), .Z(n5873) );
  AND U6289 ( .A(n5874), .B(n5875), .Z(n5869) );
  NANDN U6290 ( .A(n5876), .B(n5877), .Z(n5875) );
  NANDN U6291 ( .A(n5878), .B(n5879), .Z(n5877) );
  AND U6292 ( .A(B[797]), .B(A[3]), .Z(n5871) );
  XNOR U6293 ( .A(n5861), .B(n5880), .Z(n5872) );
  XNOR U6294 ( .A(n5859), .B(n5862), .Z(n5880) );
  NAND U6295 ( .A(A[2]), .B(B[798]), .Z(n5862) );
  NANDN U6296 ( .A(n5881), .B(n5882), .Z(n5859) );
  AND U6297 ( .A(A[0]), .B(B[799]), .Z(n5882) );
  XOR U6298 ( .A(n5864), .B(n5883), .Z(n5861) );
  NAND U6299 ( .A(A[0]), .B(B[800]), .Z(n5883) );
  NAND U6300 ( .A(B[799]), .B(A[1]), .Z(n5864) );
  NAND U6301 ( .A(n5884), .B(n5885), .Z(n479) );
  NANDN U6302 ( .A(n5886), .B(n5887), .Z(n5885) );
  OR U6303 ( .A(n5888), .B(n5889), .Z(n5887) );
  NAND U6304 ( .A(n5889), .B(n5888), .Z(n5884) );
  XOR U6305 ( .A(n481), .B(n480), .Z(\A1[797] ) );
  XOR U6306 ( .A(n5889), .B(n5890), .Z(n480) );
  XNOR U6307 ( .A(n5888), .B(n5886), .Z(n5890) );
  AND U6308 ( .A(n5891), .B(n5892), .Z(n5886) );
  NANDN U6309 ( .A(n5893), .B(n5894), .Z(n5892) );
  NANDN U6310 ( .A(n5895), .B(n5896), .Z(n5894) );
  AND U6311 ( .A(B[796]), .B(A[3]), .Z(n5888) );
  XNOR U6312 ( .A(n5878), .B(n5897), .Z(n5889) );
  XNOR U6313 ( .A(n5876), .B(n5879), .Z(n5897) );
  NAND U6314 ( .A(A[2]), .B(B[797]), .Z(n5879) );
  NANDN U6315 ( .A(n5898), .B(n5899), .Z(n5876) );
  AND U6316 ( .A(A[0]), .B(B[798]), .Z(n5899) );
  XOR U6317 ( .A(n5881), .B(n5900), .Z(n5878) );
  NAND U6318 ( .A(A[0]), .B(B[799]), .Z(n5900) );
  NAND U6319 ( .A(B[798]), .B(A[1]), .Z(n5881) );
  NAND U6320 ( .A(n5901), .B(n5902), .Z(n481) );
  NANDN U6321 ( .A(n5903), .B(n5904), .Z(n5902) );
  OR U6322 ( .A(n5905), .B(n5906), .Z(n5904) );
  NAND U6323 ( .A(n5906), .B(n5905), .Z(n5901) );
  XOR U6324 ( .A(n483), .B(n482), .Z(\A1[796] ) );
  XOR U6325 ( .A(n5906), .B(n5907), .Z(n482) );
  XNOR U6326 ( .A(n5905), .B(n5903), .Z(n5907) );
  AND U6327 ( .A(n5908), .B(n5909), .Z(n5903) );
  NANDN U6328 ( .A(n5910), .B(n5911), .Z(n5909) );
  NANDN U6329 ( .A(n5912), .B(n5913), .Z(n5911) );
  AND U6330 ( .A(B[795]), .B(A[3]), .Z(n5905) );
  XNOR U6331 ( .A(n5895), .B(n5914), .Z(n5906) );
  XNOR U6332 ( .A(n5893), .B(n5896), .Z(n5914) );
  NAND U6333 ( .A(A[2]), .B(B[796]), .Z(n5896) );
  NANDN U6334 ( .A(n5915), .B(n5916), .Z(n5893) );
  AND U6335 ( .A(A[0]), .B(B[797]), .Z(n5916) );
  XOR U6336 ( .A(n5898), .B(n5917), .Z(n5895) );
  NAND U6337 ( .A(A[0]), .B(B[798]), .Z(n5917) );
  NAND U6338 ( .A(B[797]), .B(A[1]), .Z(n5898) );
  NAND U6339 ( .A(n5918), .B(n5919), .Z(n483) );
  NANDN U6340 ( .A(n5920), .B(n5921), .Z(n5919) );
  OR U6341 ( .A(n5922), .B(n5923), .Z(n5921) );
  NAND U6342 ( .A(n5923), .B(n5922), .Z(n5918) );
  XOR U6343 ( .A(n485), .B(n484), .Z(\A1[795] ) );
  XOR U6344 ( .A(n5923), .B(n5924), .Z(n484) );
  XNOR U6345 ( .A(n5922), .B(n5920), .Z(n5924) );
  AND U6346 ( .A(n5925), .B(n5926), .Z(n5920) );
  NANDN U6347 ( .A(n5927), .B(n5928), .Z(n5926) );
  NANDN U6348 ( .A(n5929), .B(n5930), .Z(n5928) );
  AND U6349 ( .A(B[794]), .B(A[3]), .Z(n5922) );
  XNOR U6350 ( .A(n5912), .B(n5931), .Z(n5923) );
  XNOR U6351 ( .A(n5910), .B(n5913), .Z(n5931) );
  NAND U6352 ( .A(A[2]), .B(B[795]), .Z(n5913) );
  NANDN U6353 ( .A(n5932), .B(n5933), .Z(n5910) );
  AND U6354 ( .A(A[0]), .B(B[796]), .Z(n5933) );
  XOR U6355 ( .A(n5915), .B(n5934), .Z(n5912) );
  NAND U6356 ( .A(A[0]), .B(B[797]), .Z(n5934) );
  NAND U6357 ( .A(B[796]), .B(A[1]), .Z(n5915) );
  NAND U6358 ( .A(n5935), .B(n5936), .Z(n485) );
  NANDN U6359 ( .A(n5937), .B(n5938), .Z(n5936) );
  OR U6360 ( .A(n5939), .B(n5940), .Z(n5938) );
  NAND U6361 ( .A(n5940), .B(n5939), .Z(n5935) );
  XOR U6362 ( .A(n487), .B(n486), .Z(\A1[794] ) );
  XOR U6363 ( .A(n5940), .B(n5941), .Z(n486) );
  XNOR U6364 ( .A(n5939), .B(n5937), .Z(n5941) );
  AND U6365 ( .A(n5942), .B(n5943), .Z(n5937) );
  NANDN U6366 ( .A(n5944), .B(n5945), .Z(n5943) );
  NANDN U6367 ( .A(n5946), .B(n5947), .Z(n5945) );
  AND U6368 ( .A(B[793]), .B(A[3]), .Z(n5939) );
  XNOR U6369 ( .A(n5929), .B(n5948), .Z(n5940) );
  XNOR U6370 ( .A(n5927), .B(n5930), .Z(n5948) );
  NAND U6371 ( .A(A[2]), .B(B[794]), .Z(n5930) );
  NANDN U6372 ( .A(n5949), .B(n5950), .Z(n5927) );
  AND U6373 ( .A(A[0]), .B(B[795]), .Z(n5950) );
  XOR U6374 ( .A(n5932), .B(n5951), .Z(n5929) );
  NAND U6375 ( .A(A[0]), .B(B[796]), .Z(n5951) );
  NAND U6376 ( .A(B[795]), .B(A[1]), .Z(n5932) );
  NAND U6377 ( .A(n5952), .B(n5953), .Z(n487) );
  NANDN U6378 ( .A(n5954), .B(n5955), .Z(n5953) );
  OR U6379 ( .A(n5956), .B(n5957), .Z(n5955) );
  NAND U6380 ( .A(n5957), .B(n5956), .Z(n5952) );
  XOR U6381 ( .A(n489), .B(n488), .Z(\A1[793] ) );
  XOR U6382 ( .A(n5957), .B(n5958), .Z(n488) );
  XNOR U6383 ( .A(n5956), .B(n5954), .Z(n5958) );
  AND U6384 ( .A(n5959), .B(n5960), .Z(n5954) );
  NANDN U6385 ( .A(n5961), .B(n5962), .Z(n5960) );
  NANDN U6386 ( .A(n5963), .B(n5964), .Z(n5962) );
  AND U6387 ( .A(B[792]), .B(A[3]), .Z(n5956) );
  XNOR U6388 ( .A(n5946), .B(n5965), .Z(n5957) );
  XNOR U6389 ( .A(n5944), .B(n5947), .Z(n5965) );
  NAND U6390 ( .A(A[2]), .B(B[793]), .Z(n5947) );
  NANDN U6391 ( .A(n5966), .B(n5967), .Z(n5944) );
  AND U6392 ( .A(A[0]), .B(B[794]), .Z(n5967) );
  XOR U6393 ( .A(n5949), .B(n5968), .Z(n5946) );
  NAND U6394 ( .A(A[0]), .B(B[795]), .Z(n5968) );
  NAND U6395 ( .A(B[794]), .B(A[1]), .Z(n5949) );
  NAND U6396 ( .A(n5969), .B(n5970), .Z(n489) );
  NANDN U6397 ( .A(n5971), .B(n5972), .Z(n5970) );
  OR U6398 ( .A(n5973), .B(n5974), .Z(n5972) );
  NAND U6399 ( .A(n5974), .B(n5973), .Z(n5969) );
  XOR U6400 ( .A(n491), .B(n490), .Z(\A1[792] ) );
  XOR U6401 ( .A(n5974), .B(n5975), .Z(n490) );
  XNOR U6402 ( .A(n5973), .B(n5971), .Z(n5975) );
  AND U6403 ( .A(n5976), .B(n5977), .Z(n5971) );
  NANDN U6404 ( .A(n5978), .B(n5979), .Z(n5977) );
  NANDN U6405 ( .A(n5980), .B(n5981), .Z(n5979) );
  AND U6406 ( .A(B[791]), .B(A[3]), .Z(n5973) );
  XNOR U6407 ( .A(n5963), .B(n5982), .Z(n5974) );
  XNOR U6408 ( .A(n5961), .B(n5964), .Z(n5982) );
  NAND U6409 ( .A(A[2]), .B(B[792]), .Z(n5964) );
  NANDN U6410 ( .A(n5983), .B(n5984), .Z(n5961) );
  AND U6411 ( .A(A[0]), .B(B[793]), .Z(n5984) );
  XOR U6412 ( .A(n5966), .B(n5985), .Z(n5963) );
  NAND U6413 ( .A(A[0]), .B(B[794]), .Z(n5985) );
  NAND U6414 ( .A(B[793]), .B(A[1]), .Z(n5966) );
  NAND U6415 ( .A(n5986), .B(n5987), .Z(n491) );
  NANDN U6416 ( .A(n5988), .B(n5989), .Z(n5987) );
  OR U6417 ( .A(n5990), .B(n5991), .Z(n5989) );
  NAND U6418 ( .A(n5991), .B(n5990), .Z(n5986) );
  XOR U6419 ( .A(n493), .B(n492), .Z(\A1[791] ) );
  XOR U6420 ( .A(n5991), .B(n5992), .Z(n492) );
  XNOR U6421 ( .A(n5990), .B(n5988), .Z(n5992) );
  AND U6422 ( .A(n5993), .B(n5994), .Z(n5988) );
  NANDN U6423 ( .A(n5995), .B(n5996), .Z(n5994) );
  NANDN U6424 ( .A(n5997), .B(n5998), .Z(n5996) );
  AND U6425 ( .A(B[790]), .B(A[3]), .Z(n5990) );
  XNOR U6426 ( .A(n5980), .B(n5999), .Z(n5991) );
  XNOR U6427 ( .A(n5978), .B(n5981), .Z(n5999) );
  NAND U6428 ( .A(A[2]), .B(B[791]), .Z(n5981) );
  NANDN U6429 ( .A(n6000), .B(n6001), .Z(n5978) );
  AND U6430 ( .A(A[0]), .B(B[792]), .Z(n6001) );
  XOR U6431 ( .A(n5983), .B(n6002), .Z(n5980) );
  NAND U6432 ( .A(A[0]), .B(B[793]), .Z(n6002) );
  NAND U6433 ( .A(B[792]), .B(A[1]), .Z(n5983) );
  NAND U6434 ( .A(n6003), .B(n6004), .Z(n493) );
  NANDN U6435 ( .A(n6005), .B(n6006), .Z(n6004) );
  OR U6436 ( .A(n6007), .B(n6008), .Z(n6006) );
  NAND U6437 ( .A(n6008), .B(n6007), .Z(n6003) );
  XOR U6438 ( .A(n495), .B(n494), .Z(\A1[790] ) );
  XOR U6439 ( .A(n6008), .B(n6009), .Z(n494) );
  XNOR U6440 ( .A(n6007), .B(n6005), .Z(n6009) );
  AND U6441 ( .A(n6010), .B(n6011), .Z(n6005) );
  NANDN U6442 ( .A(n6012), .B(n6013), .Z(n6011) );
  NANDN U6443 ( .A(n6014), .B(n6015), .Z(n6013) );
  AND U6444 ( .A(B[789]), .B(A[3]), .Z(n6007) );
  XNOR U6445 ( .A(n5997), .B(n6016), .Z(n6008) );
  XNOR U6446 ( .A(n5995), .B(n5998), .Z(n6016) );
  NAND U6447 ( .A(A[2]), .B(B[790]), .Z(n5998) );
  NANDN U6448 ( .A(n6017), .B(n6018), .Z(n5995) );
  AND U6449 ( .A(A[0]), .B(B[791]), .Z(n6018) );
  XOR U6450 ( .A(n6000), .B(n6019), .Z(n5997) );
  NAND U6451 ( .A(A[0]), .B(B[792]), .Z(n6019) );
  NAND U6452 ( .A(B[791]), .B(A[1]), .Z(n6000) );
  NAND U6453 ( .A(n6020), .B(n6021), .Z(n495) );
  NANDN U6454 ( .A(n6022), .B(n6023), .Z(n6021) );
  OR U6455 ( .A(n6024), .B(n6025), .Z(n6023) );
  NAND U6456 ( .A(n6025), .B(n6024), .Z(n6020) );
  XOR U6457 ( .A(n477), .B(n476), .Z(\A1[78] ) );
  XOR U6458 ( .A(n5855), .B(n6026), .Z(n476) );
  XNOR U6459 ( .A(n5854), .B(n5852), .Z(n6026) );
  AND U6460 ( .A(n6027), .B(n6028), .Z(n5852) );
  NANDN U6461 ( .A(n6029), .B(n6030), .Z(n6028) );
  NANDN U6462 ( .A(n6031), .B(n6032), .Z(n6030) );
  AND U6463 ( .A(B[77]), .B(A[3]), .Z(n5854) );
  XNOR U6464 ( .A(n5844), .B(n6033), .Z(n5855) );
  XNOR U6465 ( .A(n5842), .B(n5845), .Z(n6033) );
  NAND U6466 ( .A(A[2]), .B(B[78]), .Z(n5845) );
  NANDN U6467 ( .A(n6034), .B(n6035), .Z(n5842) );
  AND U6468 ( .A(A[0]), .B(B[79]), .Z(n6035) );
  XOR U6469 ( .A(n5847), .B(n6036), .Z(n5844) );
  NAND U6470 ( .A(A[0]), .B(B[80]), .Z(n6036) );
  NAND U6471 ( .A(B[79]), .B(A[1]), .Z(n5847) );
  NAND U6472 ( .A(n6037), .B(n6038), .Z(n477) );
  NANDN U6473 ( .A(n6039), .B(n6040), .Z(n6038) );
  OR U6474 ( .A(n6041), .B(n6042), .Z(n6040) );
  NAND U6475 ( .A(n6042), .B(n6041), .Z(n6037) );
  XOR U6476 ( .A(n497), .B(n496), .Z(\A1[789] ) );
  XOR U6477 ( .A(n6025), .B(n6043), .Z(n496) );
  XNOR U6478 ( .A(n6024), .B(n6022), .Z(n6043) );
  AND U6479 ( .A(n6044), .B(n6045), .Z(n6022) );
  NANDN U6480 ( .A(n6046), .B(n6047), .Z(n6045) );
  NANDN U6481 ( .A(n6048), .B(n6049), .Z(n6047) );
  AND U6482 ( .A(B[788]), .B(A[3]), .Z(n6024) );
  XNOR U6483 ( .A(n6014), .B(n6050), .Z(n6025) );
  XNOR U6484 ( .A(n6012), .B(n6015), .Z(n6050) );
  NAND U6485 ( .A(A[2]), .B(B[789]), .Z(n6015) );
  NANDN U6486 ( .A(n6051), .B(n6052), .Z(n6012) );
  AND U6487 ( .A(A[0]), .B(B[790]), .Z(n6052) );
  XOR U6488 ( .A(n6017), .B(n6053), .Z(n6014) );
  NAND U6489 ( .A(A[0]), .B(B[791]), .Z(n6053) );
  NAND U6490 ( .A(B[790]), .B(A[1]), .Z(n6017) );
  NAND U6491 ( .A(n6054), .B(n6055), .Z(n497) );
  NANDN U6492 ( .A(n6056), .B(n6057), .Z(n6055) );
  OR U6493 ( .A(n6058), .B(n6059), .Z(n6057) );
  NAND U6494 ( .A(n6059), .B(n6058), .Z(n6054) );
  XOR U6495 ( .A(n501), .B(n500), .Z(\A1[788] ) );
  XOR U6496 ( .A(n6059), .B(n6060), .Z(n500) );
  XNOR U6497 ( .A(n6058), .B(n6056), .Z(n6060) );
  AND U6498 ( .A(n6061), .B(n6062), .Z(n6056) );
  NANDN U6499 ( .A(n6063), .B(n6064), .Z(n6062) );
  NANDN U6500 ( .A(n6065), .B(n6066), .Z(n6064) );
  AND U6501 ( .A(B[787]), .B(A[3]), .Z(n6058) );
  XNOR U6502 ( .A(n6048), .B(n6067), .Z(n6059) );
  XNOR U6503 ( .A(n6046), .B(n6049), .Z(n6067) );
  NAND U6504 ( .A(A[2]), .B(B[788]), .Z(n6049) );
  NANDN U6505 ( .A(n6068), .B(n6069), .Z(n6046) );
  AND U6506 ( .A(A[0]), .B(B[789]), .Z(n6069) );
  XOR U6507 ( .A(n6051), .B(n6070), .Z(n6048) );
  NAND U6508 ( .A(A[0]), .B(B[790]), .Z(n6070) );
  NAND U6509 ( .A(B[789]), .B(A[1]), .Z(n6051) );
  NAND U6510 ( .A(n6071), .B(n6072), .Z(n501) );
  NANDN U6511 ( .A(n6073), .B(n6074), .Z(n6072) );
  OR U6512 ( .A(n6075), .B(n6076), .Z(n6074) );
  NAND U6513 ( .A(n6076), .B(n6075), .Z(n6071) );
  XOR U6514 ( .A(n503), .B(n502), .Z(\A1[787] ) );
  XOR U6515 ( .A(n6076), .B(n6077), .Z(n502) );
  XNOR U6516 ( .A(n6075), .B(n6073), .Z(n6077) );
  AND U6517 ( .A(n6078), .B(n6079), .Z(n6073) );
  NANDN U6518 ( .A(n6080), .B(n6081), .Z(n6079) );
  NANDN U6519 ( .A(n6082), .B(n6083), .Z(n6081) );
  AND U6520 ( .A(B[786]), .B(A[3]), .Z(n6075) );
  XNOR U6521 ( .A(n6065), .B(n6084), .Z(n6076) );
  XNOR U6522 ( .A(n6063), .B(n6066), .Z(n6084) );
  NAND U6523 ( .A(A[2]), .B(B[787]), .Z(n6066) );
  NANDN U6524 ( .A(n6085), .B(n6086), .Z(n6063) );
  AND U6525 ( .A(A[0]), .B(B[788]), .Z(n6086) );
  XOR U6526 ( .A(n6068), .B(n6087), .Z(n6065) );
  NAND U6527 ( .A(A[0]), .B(B[789]), .Z(n6087) );
  NAND U6528 ( .A(B[788]), .B(A[1]), .Z(n6068) );
  NAND U6529 ( .A(n6088), .B(n6089), .Z(n503) );
  NANDN U6530 ( .A(n6090), .B(n6091), .Z(n6089) );
  OR U6531 ( .A(n6092), .B(n6093), .Z(n6091) );
  NAND U6532 ( .A(n6093), .B(n6092), .Z(n6088) );
  XOR U6533 ( .A(n505), .B(n504), .Z(\A1[786] ) );
  XOR U6534 ( .A(n6093), .B(n6094), .Z(n504) );
  XNOR U6535 ( .A(n6092), .B(n6090), .Z(n6094) );
  AND U6536 ( .A(n6095), .B(n6096), .Z(n6090) );
  NANDN U6537 ( .A(n6097), .B(n6098), .Z(n6096) );
  NANDN U6538 ( .A(n6099), .B(n6100), .Z(n6098) );
  AND U6539 ( .A(B[785]), .B(A[3]), .Z(n6092) );
  XNOR U6540 ( .A(n6082), .B(n6101), .Z(n6093) );
  XNOR U6541 ( .A(n6080), .B(n6083), .Z(n6101) );
  NAND U6542 ( .A(A[2]), .B(B[786]), .Z(n6083) );
  NANDN U6543 ( .A(n6102), .B(n6103), .Z(n6080) );
  AND U6544 ( .A(A[0]), .B(B[787]), .Z(n6103) );
  XOR U6545 ( .A(n6085), .B(n6104), .Z(n6082) );
  NAND U6546 ( .A(A[0]), .B(B[788]), .Z(n6104) );
  NAND U6547 ( .A(B[787]), .B(A[1]), .Z(n6085) );
  NAND U6548 ( .A(n6105), .B(n6106), .Z(n505) );
  NANDN U6549 ( .A(n6107), .B(n6108), .Z(n6106) );
  OR U6550 ( .A(n6109), .B(n6110), .Z(n6108) );
  NAND U6551 ( .A(n6110), .B(n6109), .Z(n6105) );
  XOR U6552 ( .A(n507), .B(n506), .Z(\A1[785] ) );
  XOR U6553 ( .A(n6110), .B(n6111), .Z(n506) );
  XNOR U6554 ( .A(n6109), .B(n6107), .Z(n6111) );
  AND U6555 ( .A(n6112), .B(n6113), .Z(n6107) );
  NANDN U6556 ( .A(n6114), .B(n6115), .Z(n6113) );
  NANDN U6557 ( .A(n6116), .B(n6117), .Z(n6115) );
  AND U6558 ( .A(B[784]), .B(A[3]), .Z(n6109) );
  XNOR U6559 ( .A(n6099), .B(n6118), .Z(n6110) );
  XNOR U6560 ( .A(n6097), .B(n6100), .Z(n6118) );
  NAND U6561 ( .A(A[2]), .B(B[785]), .Z(n6100) );
  NANDN U6562 ( .A(n6119), .B(n6120), .Z(n6097) );
  AND U6563 ( .A(A[0]), .B(B[786]), .Z(n6120) );
  XOR U6564 ( .A(n6102), .B(n6121), .Z(n6099) );
  NAND U6565 ( .A(A[0]), .B(B[787]), .Z(n6121) );
  NAND U6566 ( .A(B[786]), .B(A[1]), .Z(n6102) );
  NAND U6567 ( .A(n6122), .B(n6123), .Z(n507) );
  NANDN U6568 ( .A(n6124), .B(n6125), .Z(n6123) );
  OR U6569 ( .A(n6126), .B(n6127), .Z(n6125) );
  NAND U6570 ( .A(n6127), .B(n6126), .Z(n6122) );
  XOR U6571 ( .A(n509), .B(n508), .Z(\A1[784] ) );
  XOR U6572 ( .A(n6127), .B(n6128), .Z(n508) );
  XNOR U6573 ( .A(n6126), .B(n6124), .Z(n6128) );
  AND U6574 ( .A(n6129), .B(n6130), .Z(n6124) );
  NANDN U6575 ( .A(n6131), .B(n6132), .Z(n6130) );
  NANDN U6576 ( .A(n6133), .B(n6134), .Z(n6132) );
  AND U6577 ( .A(B[783]), .B(A[3]), .Z(n6126) );
  XNOR U6578 ( .A(n6116), .B(n6135), .Z(n6127) );
  XNOR U6579 ( .A(n6114), .B(n6117), .Z(n6135) );
  NAND U6580 ( .A(A[2]), .B(B[784]), .Z(n6117) );
  NANDN U6581 ( .A(n6136), .B(n6137), .Z(n6114) );
  AND U6582 ( .A(A[0]), .B(B[785]), .Z(n6137) );
  XOR U6583 ( .A(n6119), .B(n6138), .Z(n6116) );
  NAND U6584 ( .A(A[0]), .B(B[786]), .Z(n6138) );
  NAND U6585 ( .A(B[785]), .B(A[1]), .Z(n6119) );
  NAND U6586 ( .A(n6139), .B(n6140), .Z(n509) );
  NANDN U6587 ( .A(n6141), .B(n6142), .Z(n6140) );
  OR U6588 ( .A(n6143), .B(n6144), .Z(n6142) );
  NAND U6589 ( .A(n6144), .B(n6143), .Z(n6139) );
  XOR U6590 ( .A(n511), .B(n510), .Z(\A1[783] ) );
  XOR U6591 ( .A(n6144), .B(n6145), .Z(n510) );
  XNOR U6592 ( .A(n6143), .B(n6141), .Z(n6145) );
  AND U6593 ( .A(n6146), .B(n6147), .Z(n6141) );
  NANDN U6594 ( .A(n6148), .B(n6149), .Z(n6147) );
  NANDN U6595 ( .A(n6150), .B(n6151), .Z(n6149) );
  AND U6596 ( .A(B[782]), .B(A[3]), .Z(n6143) );
  XNOR U6597 ( .A(n6133), .B(n6152), .Z(n6144) );
  XNOR U6598 ( .A(n6131), .B(n6134), .Z(n6152) );
  NAND U6599 ( .A(A[2]), .B(B[783]), .Z(n6134) );
  NANDN U6600 ( .A(n6153), .B(n6154), .Z(n6131) );
  AND U6601 ( .A(A[0]), .B(B[784]), .Z(n6154) );
  XOR U6602 ( .A(n6136), .B(n6155), .Z(n6133) );
  NAND U6603 ( .A(A[0]), .B(B[785]), .Z(n6155) );
  NAND U6604 ( .A(B[784]), .B(A[1]), .Z(n6136) );
  NAND U6605 ( .A(n6156), .B(n6157), .Z(n511) );
  NANDN U6606 ( .A(n6158), .B(n6159), .Z(n6157) );
  OR U6607 ( .A(n6160), .B(n6161), .Z(n6159) );
  NAND U6608 ( .A(n6161), .B(n6160), .Z(n6156) );
  XOR U6609 ( .A(n513), .B(n512), .Z(\A1[782] ) );
  XOR U6610 ( .A(n6161), .B(n6162), .Z(n512) );
  XNOR U6611 ( .A(n6160), .B(n6158), .Z(n6162) );
  AND U6612 ( .A(n6163), .B(n6164), .Z(n6158) );
  NANDN U6613 ( .A(n6165), .B(n6166), .Z(n6164) );
  NANDN U6614 ( .A(n6167), .B(n6168), .Z(n6166) );
  AND U6615 ( .A(B[781]), .B(A[3]), .Z(n6160) );
  XNOR U6616 ( .A(n6150), .B(n6169), .Z(n6161) );
  XNOR U6617 ( .A(n6148), .B(n6151), .Z(n6169) );
  NAND U6618 ( .A(A[2]), .B(B[782]), .Z(n6151) );
  NANDN U6619 ( .A(n6170), .B(n6171), .Z(n6148) );
  AND U6620 ( .A(A[0]), .B(B[783]), .Z(n6171) );
  XOR U6621 ( .A(n6153), .B(n6172), .Z(n6150) );
  NAND U6622 ( .A(A[0]), .B(B[784]), .Z(n6172) );
  NAND U6623 ( .A(B[783]), .B(A[1]), .Z(n6153) );
  NAND U6624 ( .A(n6173), .B(n6174), .Z(n513) );
  NANDN U6625 ( .A(n6175), .B(n6176), .Z(n6174) );
  OR U6626 ( .A(n6177), .B(n6178), .Z(n6176) );
  NAND U6627 ( .A(n6178), .B(n6177), .Z(n6173) );
  XOR U6628 ( .A(n515), .B(n514), .Z(\A1[781] ) );
  XOR U6629 ( .A(n6178), .B(n6179), .Z(n514) );
  XNOR U6630 ( .A(n6177), .B(n6175), .Z(n6179) );
  AND U6631 ( .A(n6180), .B(n6181), .Z(n6175) );
  NANDN U6632 ( .A(n6182), .B(n6183), .Z(n6181) );
  NANDN U6633 ( .A(n6184), .B(n6185), .Z(n6183) );
  AND U6634 ( .A(B[780]), .B(A[3]), .Z(n6177) );
  XNOR U6635 ( .A(n6167), .B(n6186), .Z(n6178) );
  XNOR U6636 ( .A(n6165), .B(n6168), .Z(n6186) );
  NAND U6637 ( .A(A[2]), .B(B[781]), .Z(n6168) );
  NANDN U6638 ( .A(n6187), .B(n6188), .Z(n6165) );
  AND U6639 ( .A(A[0]), .B(B[782]), .Z(n6188) );
  XOR U6640 ( .A(n6170), .B(n6189), .Z(n6167) );
  NAND U6641 ( .A(A[0]), .B(B[783]), .Z(n6189) );
  NAND U6642 ( .A(B[782]), .B(A[1]), .Z(n6170) );
  NAND U6643 ( .A(n6190), .B(n6191), .Z(n515) );
  NANDN U6644 ( .A(n6192), .B(n6193), .Z(n6191) );
  OR U6645 ( .A(n6194), .B(n6195), .Z(n6193) );
  NAND U6646 ( .A(n6195), .B(n6194), .Z(n6190) );
  XOR U6647 ( .A(n517), .B(n516), .Z(\A1[780] ) );
  XOR U6648 ( .A(n6195), .B(n6196), .Z(n516) );
  XNOR U6649 ( .A(n6194), .B(n6192), .Z(n6196) );
  AND U6650 ( .A(n6197), .B(n6198), .Z(n6192) );
  NANDN U6651 ( .A(n6199), .B(n6200), .Z(n6198) );
  NANDN U6652 ( .A(n6201), .B(n6202), .Z(n6200) );
  AND U6653 ( .A(B[779]), .B(A[3]), .Z(n6194) );
  XNOR U6654 ( .A(n6184), .B(n6203), .Z(n6195) );
  XNOR U6655 ( .A(n6182), .B(n6185), .Z(n6203) );
  NAND U6656 ( .A(A[2]), .B(B[780]), .Z(n6185) );
  NANDN U6657 ( .A(n6204), .B(n6205), .Z(n6182) );
  AND U6658 ( .A(A[0]), .B(B[781]), .Z(n6205) );
  XOR U6659 ( .A(n6187), .B(n6206), .Z(n6184) );
  NAND U6660 ( .A(A[0]), .B(B[782]), .Z(n6206) );
  NAND U6661 ( .A(B[781]), .B(A[1]), .Z(n6187) );
  NAND U6662 ( .A(n6207), .B(n6208), .Z(n517) );
  NANDN U6663 ( .A(n6209), .B(n6210), .Z(n6208) );
  OR U6664 ( .A(n6211), .B(n6212), .Z(n6210) );
  NAND U6665 ( .A(n6212), .B(n6211), .Z(n6207) );
  XOR U6666 ( .A(n499), .B(n498), .Z(\A1[77] ) );
  XOR U6667 ( .A(n6042), .B(n6213), .Z(n498) );
  XNOR U6668 ( .A(n6041), .B(n6039), .Z(n6213) );
  AND U6669 ( .A(n6214), .B(n6215), .Z(n6039) );
  NANDN U6670 ( .A(n6216), .B(n6217), .Z(n6215) );
  NANDN U6671 ( .A(n6218), .B(n6219), .Z(n6217) );
  AND U6672 ( .A(B[76]), .B(A[3]), .Z(n6041) );
  XNOR U6673 ( .A(n6031), .B(n6220), .Z(n6042) );
  XNOR U6674 ( .A(n6029), .B(n6032), .Z(n6220) );
  NAND U6675 ( .A(A[2]), .B(B[77]), .Z(n6032) );
  NANDN U6676 ( .A(n6221), .B(n6222), .Z(n6029) );
  AND U6677 ( .A(A[0]), .B(B[78]), .Z(n6222) );
  XOR U6678 ( .A(n6034), .B(n6223), .Z(n6031) );
  NAND U6679 ( .A(A[0]), .B(B[79]), .Z(n6223) );
  NAND U6680 ( .A(B[78]), .B(A[1]), .Z(n6034) );
  NAND U6681 ( .A(n6224), .B(n6225), .Z(n499) );
  NANDN U6682 ( .A(n6226), .B(n6227), .Z(n6225) );
  OR U6683 ( .A(n6228), .B(n6229), .Z(n6227) );
  NAND U6684 ( .A(n6229), .B(n6228), .Z(n6224) );
  XOR U6685 ( .A(n519), .B(n518), .Z(\A1[779] ) );
  XOR U6686 ( .A(n6212), .B(n6230), .Z(n518) );
  XNOR U6687 ( .A(n6211), .B(n6209), .Z(n6230) );
  AND U6688 ( .A(n6231), .B(n6232), .Z(n6209) );
  NANDN U6689 ( .A(n6233), .B(n6234), .Z(n6232) );
  NANDN U6690 ( .A(n6235), .B(n6236), .Z(n6234) );
  AND U6691 ( .A(B[778]), .B(A[3]), .Z(n6211) );
  XNOR U6692 ( .A(n6201), .B(n6237), .Z(n6212) );
  XNOR U6693 ( .A(n6199), .B(n6202), .Z(n6237) );
  NAND U6694 ( .A(A[2]), .B(B[779]), .Z(n6202) );
  NANDN U6695 ( .A(n6238), .B(n6239), .Z(n6199) );
  AND U6696 ( .A(A[0]), .B(B[780]), .Z(n6239) );
  XOR U6697 ( .A(n6204), .B(n6240), .Z(n6201) );
  NAND U6698 ( .A(A[0]), .B(B[781]), .Z(n6240) );
  NAND U6699 ( .A(B[780]), .B(A[1]), .Z(n6204) );
  NAND U6700 ( .A(n6241), .B(n6242), .Z(n519) );
  NANDN U6701 ( .A(n6243), .B(n6244), .Z(n6242) );
  OR U6702 ( .A(n6245), .B(n6246), .Z(n6244) );
  NAND U6703 ( .A(n6246), .B(n6245), .Z(n6241) );
  XOR U6704 ( .A(n523), .B(n522), .Z(\A1[778] ) );
  XOR U6705 ( .A(n6246), .B(n6247), .Z(n522) );
  XNOR U6706 ( .A(n6245), .B(n6243), .Z(n6247) );
  AND U6707 ( .A(n6248), .B(n6249), .Z(n6243) );
  NANDN U6708 ( .A(n6250), .B(n6251), .Z(n6249) );
  NANDN U6709 ( .A(n6252), .B(n6253), .Z(n6251) );
  AND U6710 ( .A(B[777]), .B(A[3]), .Z(n6245) );
  XNOR U6711 ( .A(n6235), .B(n6254), .Z(n6246) );
  XNOR U6712 ( .A(n6233), .B(n6236), .Z(n6254) );
  NAND U6713 ( .A(A[2]), .B(B[778]), .Z(n6236) );
  NANDN U6714 ( .A(n6255), .B(n6256), .Z(n6233) );
  AND U6715 ( .A(A[0]), .B(B[779]), .Z(n6256) );
  XOR U6716 ( .A(n6238), .B(n6257), .Z(n6235) );
  NAND U6717 ( .A(A[0]), .B(B[780]), .Z(n6257) );
  NAND U6718 ( .A(B[779]), .B(A[1]), .Z(n6238) );
  NAND U6719 ( .A(n6258), .B(n6259), .Z(n523) );
  NANDN U6720 ( .A(n6260), .B(n6261), .Z(n6259) );
  OR U6721 ( .A(n6262), .B(n6263), .Z(n6261) );
  NAND U6722 ( .A(n6263), .B(n6262), .Z(n6258) );
  XOR U6723 ( .A(n525), .B(n524), .Z(\A1[777] ) );
  XOR U6724 ( .A(n6263), .B(n6264), .Z(n524) );
  XNOR U6725 ( .A(n6262), .B(n6260), .Z(n6264) );
  AND U6726 ( .A(n6265), .B(n6266), .Z(n6260) );
  NANDN U6727 ( .A(n6267), .B(n6268), .Z(n6266) );
  NANDN U6728 ( .A(n6269), .B(n6270), .Z(n6268) );
  AND U6729 ( .A(B[776]), .B(A[3]), .Z(n6262) );
  XNOR U6730 ( .A(n6252), .B(n6271), .Z(n6263) );
  XNOR U6731 ( .A(n6250), .B(n6253), .Z(n6271) );
  NAND U6732 ( .A(A[2]), .B(B[777]), .Z(n6253) );
  NANDN U6733 ( .A(n6272), .B(n6273), .Z(n6250) );
  AND U6734 ( .A(A[0]), .B(B[778]), .Z(n6273) );
  XOR U6735 ( .A(n6255), .B(n6274), .Z(n6252) );
  NAND U6736 ( .A(A[0]), .B(B[779]), .Z(n6274) );
  NAND U6737 ( .A(B[778]), .B(A[1]), .Z(n6255) );
  NAND U6738 ( .A(n6275), .B(n6276), .Z(n525) );
  NANDN U6739 ( .A(n6277), .B(n6278), .Z(n6276) );
  OR U6740 ( .A(n6279), .B(n6280), .Z(n6278) );
  NAND U6741 ( .A(n6280), .B(n6279), .Z(n6275) );
  XOR U6742 ( .A(n527), .B(n526), .Z(\A1[776] ) );
  XOR U6743 ( .A(n6280), .B(n6281), .Z(n526) );
  XNOR U6744 ( .A(n6279), .B(n6277), .Z(n6281) );
  AND U6745 ( .A(n6282), .B(n6283), .Z(n6277) );
  NANDN U6746 ( .A(n6284), .B(n6285), .Z(n6283) );
  NANDN U6747 ( .A(n6286), .B(n6287), .Z(n6285) );
  AND U6748 ( .A(B[775]), .B(A[3]), .Z(n6279) );
  XNOR U6749 ( .A(n6269), .B(n6288), .Z(n6280) );
  XNOR U6750 ( .A(n6267), .B(n6270), .Z(n6288) );
  NAND U6751 ( .A(A[2]), .B(B[776]), .Z(n6270) );
  NANDN U6752 ( .A(n6289), .B(n6290), .Z(n6267) );
  AND U6753 ( .A(A[0]), .B(B[777]), .Z(n6290) );
  XOR U6754 ( .A(n6272), .B(n6291), .Z(n6269) );
  NAND U6755 ( .A(A[0]), .B(B[778]), .Z(n6291) );
  NAND U6756 ( .A(B[777]), .B(A[1]), .Z(n6272) );
  NAND U6757 ( .A(n6292), .B(n6293), .Z(n527) );
  NANDN U6758 ( .A(n6294), .B(n6295), .Z(n6293) );
  OR U6759 ( .A(n6296), .B(n6297), .Z(n6295) );
  NAND U6760 ( .A(n6297), .B(n6296), .Z(n6292) );
  XOR U6761 ( .A(n529), .B(n528), .Z(\A1[775] ) );
  XOR U6762 ( .A(n6297), .B(n6298), .Z(n528) );
  XNOR U6763 ( .A(n6296), .B(n6294), .Z(n6298) );
  AND U6764 ( .A(n6299), .B(n6300), .Z(n6294) );
  NANDN U6765 ( .A(n6301), .B(n6302), .Z(n6300) );
  NANDN U6766 ( .A(n6303), .B(n6304), .Z(n6302) );
  AND U6767 ( .A(B[774]), .B(A[3]), .Z(n6296) );
  XNOR U6768 ( .A(n6286), .B(n6305), .Z(n6297) );
  XNOR U6769 ( .A(n6284), .B(n6287), .Z(n6305) );
  NAND U6770 ( .A(A[2]), .B(B[775]), .Z(n6287) );
  NANDN U6771 ( .A(n6306), .B(n6307), .Z(n6284) );
  AND U6772 ( .A(A[0]), .B(B[776]), .Z(n6307) );
  XOR U6773 ( .A(n6289), .B(n6308), .Z(n6286) );
  NAND U6774 ( .A(A[0]), .B(B[777]), .Z(n6308) );
  NAND U6775 ( .A(B[776]), .B(A[1]), .Z(n6289) );
  NAND U6776 ( .A(n6309), .B(n6310), .Z(n529) );
  NANDN U6777 ( .A(n6311), .B(n6312), .Z(n6310) );
  OR U6778 ( .A(n6313), .B(n6314), .Z(n6312) );
  NAND U6779 ( .A(n6314), .B(n6313), .Z(n6309) );
  XOR U6780 ( .A(n531), .B(n530), .Z(\A1[774] ) );
  XOR U6781 ( .A(n6314), .B(n6315), .Z(n530) );
  XNOR U6782 ( .A(n6313), .B(n6311), .Z(n6315) );
  AND U6783 ( .A(n6316), .B(n6317), .Z(n6311) );
  NANDN U6784 ( .A(n6318), .B(n6319), .Z(n6317) );
  NANDN U6785 ( .A(n6320), .B(n6321), .Z(n6319) );
  AND U6786 ( .A(B[773]), .B(A[3]), .Z(n6313) );
  XNOR U6787 ( .A(n6303), .B(n6322), .Z(n6314) );
  XNOR U6788 ( .A(n6301), .B(n6304), .Z(n6322) );
  NAND U6789 ( .A(A[2]), .B(B[774]), .Z(n6304) );
  NANDN U6790 ( .A(n6323), .B(n6324), .Z(n6301) );
  AND U6791 ( .A(A[0]), .B(B[775]), .Z(n6324) );
  XOR U6792 ( .A(n6306), .B(n6325), .Z(n6303) );
  NAND U6793 ( .A(A[0]), .B(B[776]), .Z(n6325) );
  NAND U6794 ( .A(B[775]), .B(A[1]), .Z(n6306) );
  NAND U6795 ( .A(n6326), .B(n6327), .Z(n531) );
  NANDN U6796 ( .A(n6328), .B(n6329), .Z(n6327) );
  OR U6797 ( .A(n6330), .B(n6331), .Z(n6329) );
  NAND U6798 ( .A(n6331), .B(n6330), .Z(n6326) );
  XOR U6799 ( .A(n533), .B(n532), .Z(\A1[773] ) );
  XOR U6800 ( .A(n6331), .B(n6332), .Z(n532) );
  XNOR U6801 ( .A(n6330), .B(n6328), .Z(n6332) );
  AND U6802 ( .A(n6333), .B(n6334), .Z(n6328) );
  NANDN U6803 ( .A(n6335), .B(n6336), .Z(n6334) );
  NANDN U6804 ( .A(n6337), .B(n6338), .Z(n6336) );
  AND U6805 ( .A(B[772]), .B(A[3]), .Z(n6330) );
  XNOR U6806 ( .A(n6320), .B(n6339), .Z(n6331) );
  XNOR U6807 ( .A(n6318), .B(n6321), .Z(n6339) );
  NAND U6808 ( .A(A[2]), .B(B[773]), .Z(n6321) );
  NANDN U6809 ( .A(n6340), .B(n6341), .Z(n6318) );
  AND U6810 ( .A(A[0]), .B(B[774]), .Z(n6341) );
  XOR U6811 ( .A(n6323), .B(n6342), .Z(n6320) );
  NAND U6812 ( .A(A[0]), .B(B[775]), .Z(n6342) );
  NAND U6813 ( .A(B[774]), .B(A[1]), .Z(n6323) );
  NAND U6814 ( .A(n6343), .B(n6344), .Z(n533) );
  NANDN U6815 ( .A(n6345), .B(n6346), .Z(n6344) );
  OR U6816 ( .A(n6347), .B(n6348), .Z(n6346) );
  NAND U6817 ( .A(n6348), .B(n6347), .Z(n6343) );
  XOR U6818 ( .A(n535), .B(n534), .Z(\A1[772] ) );
  XOR U6819 ( .A(n6348), .B(n6349), .Z(n534) );
  XNOR U6820 ( .A(n6347), .B(n6345), .Z(n6349) );
  AND U6821 ( .A(n6350), .B(n6351), .Z(n6345) );
  NANDN U6822 ( .A(n6352), .B(n6353), .Z(n6351) );
  NANDN U6823 ( .A(n6354), .B(n6355), .Z(n6353) );
  AND U6824 ( .A(B[771]), .B(A[3]), .Z(n6347) );
  XNOR U6825 ( .A(n6337), .B(n6356), .Z(n6348) );
  XNOR U6826 ( .A(n6335), .B(n6338), .Z(n6356) );
  NAND U6827 ( .A(A[2]), .B(B[772]), .Z(n6338) );
  NANDN U6828 ( .A(n6357), .B(n6358), .Z(n6335) );
  AND U6829 ( .A(A[0]), .B(B[773]), .Z(n6358) );
  XOR U6830 ( .A(n6340), .B(n6359), .Z(n6337) );
  NAND U6831 ( .A(A[0]), .B(B[774]), .Z(n6359) );
  NAND U6832 ( .A(B[773]), .B(A[1]), .Z(n6340) );
  NAND U6833 ( .A(n6360), .B(n6361), .Z(n535) );
  NANDN U6834 ( .A(n6362), .B(n6363), .Z(n6361) );
  OR U6835 ( .A(n6364), .B(n6365), .Z(n6363) );
  NAND U6836 ( .A(n6365), .B(n6364), .Z(n6360) );
  XOR U6837 ( .A(n537), .B(n536), .Z(\A1[771] ) );
  XOR U6838 ( .A(n6365), .B(n6366), .Z(n536) );
  XNOR U6839 ( .A(n6364), .B(n6362), .Z(n6366) );
  AND U6840 ( .A(n6367), .B(n6368), .Z(n6362) );
  NANDN U6841 ( .A(n6369), .B(n6370), .Z(n6368) );
  NANDN U6842 ( .A(n6371), .B(n6372), .Z(n6370) );
  AND U6843 ( .A(B[770]), .B(A[3]), .Z(n6364) );
  XNOR U6844 ( .A(n6354), .B(n6373), .Z(n6365) );
  XNOR U6845 ( .A(n6352), .B(n6355), .Z(n6373) );
  NAND U6846 ( .A(A[2]), .B(B[771]), .Z(n6355) );
  NANDN U6847 ( .A(n6374), .B(n6375), .Z(n6352) );
  AND U6848 ( .A(A[0]), .B(B[772]), .Z(n6375) );
  XOR U6849 ( .A(n6357), .B(n6376), .Z(n6354) );
  NAND U6850 ( .A(A[0]), .B(B[773]), .Z(n6376) );
  NAND U6851 ( .A(B[772]), .B(A[1]), .Z(n6357) );
  NAND U6852 ( .A(n6377), .B(n6378), .Z(n537) );
  NANDN U6853 ( .A(n6379), .B(n6380), .Z(n6378) );
  OR U6854 ( .A(n6381), .B(n6382), .Z(n6380) );
  NAND U6855 ( .A(n6382), .B(n6381), .Z(n6377) );
  XOR U6856 ( .A(n539), .B(n538), .Z(\A1[770] ) );
  XOR U6857 ( .A(n6382), .B(n6383), .Z(n538) );
  XNOR U6858 ( .A(n6381), .B(n6379), .Z(n6383) );
  AND U6859 ( .A(n6384), .B(n6385), .Z(n6379) );
  NANDN U6860 ( .A(n6386), .B(n6387), .Z(n6385) );
  NANDN U6861 ( .A(n6388), .B(n6389), .Z(n6387) );
  AND U6862 ( .A(B[769]), .B(A[3]), .Z(n6381) );
  XNOR U6863 ( .A(n6371), .B(n6390), .Z(n6382) );
  XNOR U6864 ( .A(n6369), .B(n6372), .Z(n6390) );
  NAND U6865 ( .A(A[2]), .B(B[770]), .Z(n6372) );
  NANDN U6866 ( .A(n6391), .B(n6392), .Z(n6369) );
  AND U6867 ( .A(A[0]), .B(B[771]), .Z(n6392) );
  XOR U6868 ( .A(n6374), .B(n6393), .Z(n6371) );
  NAND U6869 ( .A(A[0]), .B(B[772]), .Z(n6393) );
  NAND U6870 ( .A(B[771]), .B(A[1]), .Z(n6374) );
  NAND U6871 ( .A(n6394), .B(n6395), .Z(n539) );
  NANDN U6872 ( .A(n6396), .B(n6397), .Z(n6395) );
  OR U6873 ( .A(n6398), .B(n6399), .Z(n6397) );
  NAND U6874 ( .A(n6399), .B(n6398), .Z(n6394) );
  XOR U6875 ( .A(n521), .B(n520), .Z(\A1[76] ) );
  XOR U6876 ( .A(n6229), .B(n6400), .Z(n520) );
  XNOR U6877 ( .A(n6228), .B(n6226), .Z(n6400) );
  AND U6878 ( .A(n6401), .B(n6402), .Z(n6226) );
  NANDN U6879 ( .A(n6403), .B(n6404), .Z(n6402) );
  NANDN U6880 ( .A(n6405), .B(n6406), .Z(n6404) );
  AND U6881 ( .A(B[75]), .B(A[3]), .Z(n6228) );
  XNOR U6882 ( .A(n6218), .B(n6407), .Z(n6229) );
  XNOR U6883 ( .A(n6216), .B(n6219), .Z(n6407) );
  NAND U6884 ( .A(A[2]), .B(B[76]), .Z(n6219) );
  NANDN U6885 ( .A(n6408), .B(n6409), .Z(n6216) );
  AND U6886 ( .A(A[0]), .B(B[77]), .Z(n6409) );
  XOR U6887 ( .A(n6221), .B(n6410), .Z(n6218) );
  NAND U6888 ( .A(A[0]), .B(B[78]), .Z(n6410) );
  NAND U6889 ( .A(B[77]), .B(A[1]), .Z(n6221) );
  NAND U6890 ( .A(n6411), .B(n6412), .Z(n521) );
  NANDN U6891 ( .A(n6413), .B(n6414), .Z(n6412) );
  OR U6892 ( .A(n6415), .B(n6416), .Z(n6414) );
  NAND U6893 ( .A(n6416), .B(n6415), .Z(n6411) );
  XOR U6894 ( .A(n541), .B(n540), .Z(\A1[769] ) );
  XOR U6895 ( .A(n6399), .B(n6417), .Z(n540) );
  XNOR U6896 ( .A(n6398), .B(n6396), .Z(n6417) );
  AND U6897 ( .A(n6418), .B(n6419), .Z(n6396) );
  NANDN U6898 ( .A(n6420), .B(n6421), .Z(n6419) );
  NANDN U6899 ( .A(n6422), .B(n6423), .Z(n6421) );
  AND U6900 ( .A(B[768]), .B(A[3]), .Z(n6398) );
  XNOR U6901 ( .A(n6388), .B(n6424), .Z(n6399) );
  XNOR U6902 ( .A(n6386), .B(n6389), .Z(n6424) );
  NAND U6903 ( .A(A[2]), .B(B[769]), .Z(n6389) );
  NANDN U6904 ( .A(n6425), .B(n6426), .Z(n6386) );
  AND U6905 ( .A(A[0]), .B(B[770]), .Z(n6426) );
  XOR U6906 ( .A(n6391), .B(n6427), .Z(n6388) );
  NAND U6907 ( .A(A[0]), .B(B[771]), .Z(n6427) );
  NAND U6908 ( .A(B[770]), .B(A[1]), .Z(n6391) );
  NAND U6909 ( .A(n6428), .B(n6429), .Z(n541) );
  NANDN U6910 ( .A(n6430), .B(n6431), .Z(n6429) );
  OR U6911 ( .A(n6432), .B(n6433), .Z(n6431) );
  NAND U6912 ( .A(n6433), .B(n6432), .Z(n6428) );
  XOR U6913 ( .A(n545), .B(n544), .Z(\A1[768] ) );
  XOR U6914 ( .A(n6433), .B(n6434), .Z(n544) );
  XNOR U6915 ( .A(n6432), .B(n6430), .Z(n6434) );
  AND U6916 ( .A(n6435), .B(n6436), .Z(n6430) );
  NANDN U6917 ( .A(n6437), .B(n6438), .Z(n6436) );
  NANDN U6918 ( .A(n6439), .B(n6440), .Z(n6438) );
  AND U6919 ( .A(B[767]), .B(A[3]), .Z(n6432) );
  XNOR U6920 ( .A(n6422), .B(n6441), .Z(n6433) );
  XNOR U6921 ( .A(n6420), .B(n6423), .Z(n6441) );
  NAND U6922 ( .A(A[2]), .B(B[768]), .Z(n6423) );
  NANDN U6923 ( .A(n6442), .B(n6443), .Z(n6420) );
  AND U6924 ( .A(A[0]), .B(B[769]), .Z(n6443) );
  XOR U6925 ( .A(n6425), .B(n6444), .Z(n6422) );
  NAND U6926 ( .A(A[0]), .B(B[770]), .Z(n6444) );
  NAND U6927 ( .A(B[769]), .B(A[1]), .Z(n6425) );
  NAND U6928 ( .A(n6445), .B(n6446), .Z(n545) );
  NANDN U6929 ( .A(n6447), .B(n6448), .Z(n6446) );
  OR U6930 ( .A(n6449), .B(n6450), .Z(n6448) );
  NAND U6931 ( .A(n6450), .B(n6449), .Z(n6445) );
  XOR U6932 ( .A(n547), .B(n546), .Z(\A1[767] ) );
  XOR U6933 ( .A(n6450), .B(n6451), .Z(n546) );
  XNOR U6934 ( .A(n6449), .B(n6447), .Z(n6451) );
  AND U6935 ( .A(n6452), .B(n6453), .Z(n6447) );
  NANDN U6936 ( .A(n6454), .B(n6455), .Z(n6453) );
  NANDN U6937 ( .A(n6456), .B(n6457), .Z(n6455) );
  AND U6938 ( .A(B[766]), .B(A[3]), .Z(n6449) );
  XNOR U6939 ( .A(n6439), .B(n6458), .Z(n6450) );
  XNOR U6940 ( .A(n6437), .B(n6440), .Z(n6458) );
  NAND U6941 ( .A(A[2]), .B(B[767]), .Z(n6440) );
  NANDN U6942 ( .A(n6459), .B(n6460), .Z(n6437) );
  AND U6943 ( .A(A[0]), .B(B[768]), .Z(n6460) );
  XOR U6944 ( .A(n6442), .B(n6461), .Z(n6439) );
  NAND U6945 ( .A(A[0]), .B(B[769]), .Z(n6461) );
  NAND U6946 ( .A(B[768]), .B(A[1]), .Z(n6442) );
  NAND U6947 ( .A(n6462), .B(n6463), .Z(n547) );
  NANDN U6948 ( .A(n6464), .B(n6465), .Z(n6463) );
  OR U6949 ( .A(n6466), .B(n6467), .Z(n6465) );
  NAND U6950 ( .A(n6467), .B(n6466), .Z(n6462) );
  XOR U6951 ( .A(n549), .B(n548), .Z(\A1[766] ) );
  XOR U6952 ( .A(n6467), .B(n6468), .Z(n548) );
  XNOR U6953 ( .A(n6466), .B(n6464), .Z(n6468) );
  AND U6954 ( .A(n6469), .B(n6470), .Z(n6464) );
  NANDN U6955 ( .A(n6471), .B(n6472), .Z(n6470) );
  NANDN U6956 ( .A(n6473), .B(n6474), .Z(n6472) );
  AND U6957 ( .A(B[765]), .B(A[3]), .Z(n6466) );
  XNOR U6958 ( .A(n6456), .B(n6475), .Z(n6467) );
  XNOR U6959 ( .A(n6454), .B(n6457), .Z(n6475) );
  NAND U6960 ( .A(A[2]), .B(B[766]), .Z(n6457) );
  NANDN U6961 ( .A(n6476), .B(n6477), .Z(n6454) );
  AND U6962 ( .A(A[0]), .B(B[767]), .Z(n6477) );
  XOR U6963 ( .A(n6459), .B(n6478), .Z(n6456) );
  NAND U6964 ( .A(A[0]), .B(B[768]), .Z(n6478) );
  NAND U6965 ( .A(B[767]), .B(A[1]), .Z(n6459) );
  NAND U6966 ( .A(n6479), .B(n6480), .Z(n549) );
  NANDN U6967 ( .A(n6481), .B(n6482), .Z(n6480) );
  OR U6968 ( .A(n6483), .B(n6484), .Z(n6482) );
  NAND U6969 ( .A(n6484), .B(n6483), .Z(n6479) );
  XOR U6970 ( .A(n551), .B(n550), .Z(\A1[765] ) );
  XOR U6971 ( .A(n6484), .B(n6485), .Z(n550) );
  XNOR U6972 ( .A(n6483), .B(n6481), .Z(n6485) );
  AND U6973 ( .A(n6486), .B(n6487), .Z(n6481) );
  NANDN U6974 ( .A(n6488), .B(n6489), .Z(n6487) );
  NANDN U6975 ( .A(n6490), .B(n6491), .Z(n6489) );
  AND U6976 ( .A(B[764]), .B(A[3]), .Z(n6483) );
  XNOR U6977 ( .A(n6473), .B(n6492), .Z(n6484) );
  XNOR U6978 ( .A(n6471), .B(n6474), .Z(n6492) );
  NAND U6979 ( .A(A[2]), .B(B[765]), .Z(n6474) );
  NANDN U6980 ( .A(n6493), .B(n6494), .Z(n6471) );
  AND U6981 ( .A(A[0]), .B(B[766]), .Z(n6494) );
  XOR U6982 ( .A(n6476), .B(n6495), .Z(n6473) );
  NAND U6983 ( .A(A[0]), .B(B[767]), .Z(n6495) );
  NAND U6984 ( .A(B[766]), .B(A[1]), .Z(n6476) );
  NAND U6985 ( .A(n6496), .B(n6497), .Z(n551) );
  NANDN U6986 ( .A(n6498), .B(n6499), .Z(n6497) );
  OR U6987 ( .A(n6500), .B(n6501), .Z(n6499) );
  NAND U6988 ( .A(n6501), .B(n6500), .Z(n6496) );
  XOR U6989 ( .A(n553), .B(n552), .Z(\A1[764] ) );
  XOR U6990 ( .A(n6501), .B(n6502), .Z(n552) );
  XNOR U6991 ( .A(n6500), .B(n6498), .Z(n6502) );
  AND U6992 ( .A(n6503), .B(n6504), .Z(n6498) );
  NANDN U6993 ( .A(n6505), .B(n6506), .Z(n6504) );
  NANDN U6994 ( .A(n6507), .B(n6508), .Z(n6506) );
  AND U6995 ( .A(B[763]), .B(A[3]), .Z(n6500) );
  XNOR U6996 ( .A(n6490), .B(n6509), .Z(n6501) );
  XNOR U6997 ( .A(n6488), .B(n6491), .Z(n6509) );
  NAND U6998 ( .A(A[2]), .B(B[764]), .Z(n6491) );
  NANDN U6999 ( .A(n6510), .B(n6511), .Z(n6488) );
  AND U7000 ( .A(A[0]), .B(B[765]), .Z(n6511) );
  XOR U7001 ( .A(n6493), .B(n6512), .Z(n6490) );
  NAND U7002 ( .A(A[0]), .B(B[766]), .Z(n6512) );
  NAND U7003 ( .A(B[765]), .B(A[1]), .Z(n6493) );
  NAND U7004 ( .A(n6513), .B(n6514), .Z(n553) );
  NANDN U7005 ( .A(n6515), .B(n6516), .Z(n6514) );
  OR U7006 ( .A(n6517), .B(n6518), .Z(n6516) );
  NAND U7007 ( .A(n6518), .B(n6517), .Z(n6513) );
  XOR U7008 ( .A(n555), .B(n554), .Z(\A1[763] ) );
  XOR U7009 ( .A(n6518), .B(n6519), .Z(n554) );
  XNOR U7010 ( .A(n6517), .B(n6515), .Z(n6519) );
  AND U7011 ( .A(n6520), .B(n6521), .Z(n6515) );
  NANDN U7012 ( .A(n6522), .B(n6523), .Z(n6521) );
  NANDN U7013 ( .A(n6524), .B(n6525), .Z(n6523) );
  AND U7014 ( .A(B[762]), .B(A[3]), .Z(n6517) );
  XNOR U7015 ( .A(n6507), .B(n6526), .Z(n6518) );
  XNOR U7016 ( .A(n6505), .B(n6508), .Z(n6526) );
  NAND U7017 ( .A(A[2]), .B(B[763]), .Z(n6508) );
  NANDN U7018 ( .A(n6527), .B(n6528), .Z(n6505) );
  AND U7019 ( .A(A[0]), .B(B[764]), .Z(n6528) );
  XOR U7020 ( .A(n6510), .B(n6529), .Z(n6507) );
  NAND U7021 ( .A(A[0]), .B(B[765]), .Z(n6529) );
  NAND U7022 ( .A(B[764]), .B(A[1]), .Z(n6510) );
  NAND U7023 ( .A(n6530), .B(n6531), .Z(n555) );
  NANDN U7024 ( .A(n6532), .B(n6533), .Z(n6531) );
  OR U7025 ( .A(n6534), .B(n6535), .Z(n6533) );
  NAND U7026 ( .A(n6535), .B(n6534), .Z(n6530) );
  XOR U7027 ( .A(n557), .B(n556), .Z(\A1[762] ) );
  XOR U7028 ( .A(n6535), .B(n6536), .Z(n556) );
  XNOR U7029 ( .A(n6534), .B(n6532), .Z(n6536) );
  AND U7030 ( .A(n6537), .B(n6538), .Z(n6532) );
  NANDN U7031 ( .A(n6539), .B(n6540), .Z(n6538) );
  NANDN U7032 ( .A(n6541), .B(n6542), .Z(n6540) );
  AND U7033 ( .A(B[761]), .B(A[3]), .Z(n6534) );
  XNOR U7034 ( .A(n6524), .B(n6543), .Z(n6535) );
  XNOR U7035 ( .A(n6522), .B(n6525), .Z(n6543) );
  NAND U7036 ( .A(A[2]), .B(B[762]), .Z(n6525) );
  NANDN U7037 ( .A(n6544), .B(n6545), .Z(n6522) );
  AND U7038 ( .A(A[0]), .B(B[763]), .Z(n6545) );
  XOR U7039 ( .A(n6527), .B(n6546), .Z(n6524) );
  NAND U7040 ( .A(A[0]), .B(B[764]), .Z(n6546) );
  NAND U7041 ( .A(B[763]), .B(A[1]), .Z(n6527) );
  NAND U7042 ( .A(n6547), .B(n6548), .Z(n557) );
  NANDN U7043 ( .A(n6549), .B(n6550), .Z(n6548) );
  OR U7044 ( .A(n6551), .B(n6552), .Z(n6550) );
  NAND U7045 ( .A(n6552), .B(n6551), .Z(n6547) );
  XOR U7046 ( .A(n559), .B(n558), .Z(\A1[761] ) );
  XOR U7047 ( .A(n6552), .B(n6553), .Z(n558) );
  XNOR U7048 ( .A(n6551), .B(n6549), .Z(n6553) );
  AND U7049 ( .A(n6554), .B(n6555), .Z(n6549) );
  NANDN U7050 ( .A(n6556), .B(n6557), .Z(n6555) );
  NANDN U7051 ( .A(n6558), .B(n6559), .Z(n6557) );
  AND U7052 ( .A(B[760]), .B(A[3]), .Z(n6551) );
  XNOR U7053 ( .A(n6541), .B(n6560), .Z(n6552) );
  XNOR U7054 ( .A(n6539), .B(n6542), .Z(n6560) );
  NAND U7055 ( .A(A[2]), .B(B[761]), .Z(n6542) );
  NANDN U7056 ( .A(n6561), .B(n6562), .Z(n6539) );
  AND U7057 ( .A(A[0]), .B(B[762]), .Z(n6562) );
  XOR U7058 ( .A(n6544), .B(n6563), .Z(n6541) );
  NAND U7059 ( .A(A[0]), .B(B[763]), .Z(n6563) );
  NAND U7060 ( .A(B[762]), .B(A[1]), .Z(n6544) );
  NAND U7061 ( .A(n6564), .B(n6565), .Z(n559) );
  NANDN U7062 ( .A(n6566), .B(n6567), .Z(n6565) );
  OR U7063 ( .A(n6568), .B(n6569), .Z(n6567) );
  NAND U7064 ( .A(n6569), .B(n6568), .Z(n6564) );
  XOR U7065 ( .A(n561), .B(n560), .Z(\A1[760] ) );
  XOR U7066 ( .A(n6569), .B(n6570), .Z(n560) );
  XNOR U7067 ( .A(n6568), .B(n6566), .Z(n6570) );
  AND U7068 ( .A(n6571), .B(n6572), .Z(n6566) );
  NANDN U7069 ( .A(n6573), .B(n6574), .Z(n6572) );
  NANDN U7070 ( .A(n6575), .B(n6576), .Z(n6574) );
  AND U7071 ( .A(B[759]), .B(A[3]), .Z(n6568) );
  XNOR U7072 ( .A(n6558), .B(n6577), .Z(n6569) );
  XNOR U7073 ( .A(n6556), .B(n6559), .Z(n6577) );
  NAND U7074 ( .A(A[2]), .B(B[760]), .Z(n6559) );
  NANDN U7075 ( .A(n6578), .B(n6579), .Z(n6556) );
  AND U7076 ( .A(A[0]), .B(B[761]), .Z(n6579) );
  XOR U7077 ( .A(n6561), .B(n6580), .Z(n6558) );
  NAND U7078 ( .A(A[0]), .B(B[762]), .Z(n6580) );
  NAND U7079 ( .A(B[761]), .B(A[1]), .Z(n6561) );
  NAND U7080 ( .A(n6581), .B(n6582), .Z(n561) );
  NANDN U7081 ( .A(n6583), .B(n6584), .Z(n6582) );
  OR U7082 ( .A(n6585), .B(n6586), .Z(n6584) );
  NAND U7083 ( .A(n6586), .B(n6585), .Z(n6581) );
  XOR U7084 ( .A(n543), .B(n542), .Z(\A1[75] ) );
  XOR U7085 ( .A(n6416), .B(n6587), .Z(n542) );
  XNOR U7086 ( .A(n6415), .B(n6413), .Z(n6587) );
  AND U7087 ( .A(n6588), .B(n6589), .Z(n6413) );
  NANDN U7088 ( .A(n6590), .B(n6591), .Z(n6589) );
  NANDN U7089 ( .A(n6592), .B(n6593), .Z(n6591) );
  AND U7090 ( .A(B[74]), .B(A[3]), .Z(n6415) );
  XNOR U7091 ( .A(n6405), .B(n6594), .Z(n6416) );
  XNOR U7092 ( .A(n6403), .B(n6406), .Z(n6594) );
  NAND U7093 ( .A(A[2]), .B(B[75]), .Z(n6406) );
  NANDN U7094 ( .A(n6595), .B(n6596), .Z(n6403) );
  AND U7095 ( .A(A[0]), .B(B[76]), .Z(n6596) );
  XOR U7096 ( .A(n6408), .B(n6597), .Z(n6405) );
  NAND U7097 ( .A(A[0]), .B(B[77]), .Z(n6597) );
  NAND U7098 ( .A(B[76]), .B(A[1]), .Z(n6408) );
  NAND U7099 ( .A(n6598), .B(n6599), .Z(n543) );
  NANDN U7100 ( .A(n6600), .B(n6601), .Z(n6599) );
  OR U7101 ( .A(n6602), .B(n6603), .Z(n6601) );
  NAND U7102 ( .A(n6603), .B(n6602), .Z(n6598) );
  XOR U7103 ( .A(n563), .B(n562), .Z(\A1[759] ) );
  XOR U7104 ( .A(n6586), .B(n6604), .Z(n562) );
  XNOR U7105 ( .A(n6585), .B(n6583), .Z(n6604) );
  AND U7106 ( .A(n6605), .B(n6606), .Z(n6583) );
  NANDN U7107 ( .A(n6607), .B(n6608), .Z(n6606) );
  NANDN U7108 ( .A(n6609), .B(n6610), .Z(n6608) );
  AND U7109 ( .A(B[758]), .B(A[3]), .Z(n6585) );
  XNOR U7110 ( .A(n6575), .B(n6611), .Z(n6586) );
  XNOR U7111 ( .A(n6573), .B(n6576), .Z(n6611) );
  NAND U7112 ( .A(A[2]), .B(B[759]), .Z(n6576) );
  NANDN U7113 ( .A(n6612), .B(n6613), .Z(n6573) );
  AND U7114 ( .A(A[0]), .B(B[760]), .Z(n6613) );
  XOR U7115 ( .A(n6578), .B(n6614), .Z(n6575) );
  NAND U7116 ( .A(A[0]), .B(B[761]), .Z(n6614) );
  NAND U7117 ( .A(B[760]), .B(A[1]), .Z(n6578) );
  NAND U7118 ( .A(n6615), .B(n6616), .Z(n563) );
  NANDN U7119 ( .A(n6617), .B(n6618), .Z(n6616) );
  OR U7120 ( .A(n6619), .B(n6620), .Z(n6618) );
  NAND U7121 ( .A(n6620), .B(n6619), .Z(n6615) );
  XOR U7122 ( .A(n567), .B(n566), .Z(\A1[758] ) );
  XOR U7123 ( .A(n6620), .B(n6621), .Z(n566) );
  XNOR U7124 ( .A(n6619), .B(n6617), .Z(n6621) );
  AND U7125 ( .A(n6622), .B(n6623), .Z(n6617) );
  NANDN U7126 ( .A(n6624), .B(n6625), .Z(n6623) );
  NANDN U7127 ( .A(n6626), .B(n6627), .Z(n6625) );
  AND U7128 ( .A(B[757]), .B(A[3]), .Z(n6619) );
  XNOR U7129 ( .A(n6609), .B(n6628), .Z(n6620) );
  XNOR U7130 ( .A(n6607), .B(n6610), .Z(n6628) );
  NAND U7131 ( .A(A[2]), .B(B[758]), .Z(n6610) );
  NANDN U7132 ( .A(n6629), .B(n6630), .Z(n6607) );
  AND U7133 ( .A(A[0]), .B(B[759]), .Z(n6630) );
  XOR U7134 ( .A(n6612), .B(n6631), .Z(n6609) );
  NAND U7135 ( .A(A[0]), .B(B[760]), .Z(n6631) );
  NAND U7136 ( .A(B[759]), .B(A[1]), .Z(n6612) );
  NAND U7137 ( .A(n6632), .B(n6633), .Z(n567) );
  NANDN U7138 ( .A(n6634), .B(n6635), .Z(n6633) );
  OR U7139 ( .A(n6636), .B(n6637), .Z(n6635) );
  NAND U7140 ( .A(n6637), .B(n6636), .Z(n6632) );
  XOR U7141 ( .A(n569), .B(n568), .Z(\A1[757] ) );
  XOR U7142 ( .A(n6637), .B(n6638), .Z(n568) );
  XNOR U7143 ( .A(n6636), .B(n6634), .Z(n6638) );
  AND U7144 ( .A(n6639), .B(n6640), .Z(n6634) );
  NANDN U7145 ( .A(n6641), .B(n6642), .Z(n6640) );
  NANDN U7146 ( .A(n6643), .B(n6644), .Z(n6642) );
  AND U7147 ( .A(B[756]), .B(A[3]), .Z(n6636) );
  XNOR U7148 ( .A(n6626), .B(n6645), .Z(n6637) );
  XNOR U7149 ( .A(n6624), .B(n6627), .Z(n6645) );
  NAND U7150 ( .A(A[2]), .B(B[757]), .Z(n6627) );
  NANDN U7151 ( .A(n6646), .B(n6647), .Z(n6624) );
  AND U7152 ( .A(A[0]), .B(B[758]), .Z(n6647) );
  XOR U7153 ( .A(n6629), .B(n6648), .Z(n6626) );
  NAND U7154 ( .A(A[0]), .B(B[759]), .Z(n6648) );
  NAND U7155 ( .A(B[758]), .B(A[1]), .Z(n6629) );
  NAND U7156 ( .A(n6649), .B(n6650), .Z(n569) );
  NANDN U7157 ( .A(n6651), .B(n6652), .Z(n6650) );
  OR U7158 ( .A(n6653), .B(n6654), .Z(n6652) );
  NAND U7159 ( .A(n6654), .B(n6653), .Z(n6649) );
  XOR U7160 ( .A(n571), .B(n570), .Z(\A1[756] ) );
  XOR U7161 ( .A(n6654), .B(n6655), .Z(n570) );
  XNOR U7162 ( .A(n6653), .B(n6651), .Z(n6655) );
  AND U7163 ( .A(n6656), .B(n6657), .Z(n6651) );
  NANDN U7164 ( .A(n6658), .B(n6659), .Z(n6657) );
  NANDN U7165 ( .A(n6660), .B(n6661), .Z(n6659) );
  AND U7166 ( .A(B[755]), .B(A[3]), .Z(n6653) );
  XNOR U7167 ( .A(n6643), .B(n6662), .Z(n6654) );
  XNOR U7168 ( .A(n6641), .B(n6644), .Z(n6662) );
  NAND U7169 ( .A(A[2]), .B(B[756]), .Z(n6644) );
  NANDN U7170 ( .A(n6663), .B(n6664), .Z(n6641) );
  AND U7171 ( .A(A[0]), .B(B[757]), .Z(n6664) );
  XOR U7172 ( .A(n6646), .B(n6665), .Z(n6643) );
  NAND U7173 ( .A(A[0]), .B(B[758]), .Z(n6665) );
  NAND U7174 ( .A(B[757]), .B(A[1]), .Z(n6646) );
  NAND U7175 ( .A(n6666), .B(n6667), .Z(n571) );
  NANDN U7176 ( .A(n6668), .B(n6669), .Z(n6667) );
  OR U7177 ( .A(n6670), .B(n6671), .Z(n6669) );
  NAND U7178 ( .A(n6671), .B(n6670), .Z(n6666) );
  XOR U7179 ( .A(n573), .B(n572), .Z(\A1[755] ) );
  XOR U7180 ( .A(n6671), .B(n6672), .Z(n572) );
  XNOR U7181 ( .A(n6670), .B(n6668), .Z(n6672) );
  AND U7182 ( .A(n6673), .B(n6674), .Z(n6668) );
  NANDN U7183 ( .A(n6675), .B(n6676), .Z(n6674) );
  NANDN U7184 ( .A(n6677), .B(n6678), .Z(n6676) );
  AND U7185 ( .A(B[754]), .B(A[3]), .Z(n6670) );
  XNOR U7186 ( .A(n6660), .B(n6679), .Z(n6671) );
  XNOR U7187 ( .A(n6658), .B(n6661), .Z(n6679) );
  NAND U7188 ( .A(A[2]), .B(B[755]), .Z(n6661) );
  NANDN U7189 ( .A(n6680), .B(n6681), .Z(n6658) );
  AND U7190 ( .A(A[0]), .B(B[756]), .Z(n6681) );
  XOR U7191 ( .A(n6663), .B(n6682), .Z(n6660) );
  NAND U7192 ( .A(A[0]), .B(B[757]), .Z(n6682) );
  NAND U7193 ( .A(B[756]), .B(A[1]), .Z(n6663) );
  NAND U7194 ( .A(n6683), .B(n6684), .Z(n573) );
  NANDN U7195 ( .A(n6685), .B(n6686), .Z(n6684) );
  OR U7196 ( .A(n6687), .B(n6688), .Z(n6686) );
  NAND U7197 ( .A(n6688), .B(n6687), .Z(n6683) );
  XOR U7198 ( .A(n575), .B(n574), .Z(\A1[754] ) );
  XOR U7199 ( .A(n6688), .B(n6689), .Z(n574) );
  XNOR U7200 ( .A(n6687), .B(n6685), .Z(n6689) );
  AND U7201 ( .A(n6690), .B(n6691), .Z(n6685) );
  NANDN U7202 ( .A(n6692), .B(n6693), .Z(n6691) );
  NANDN U7203 ( .A(n6694), .B(n6695), .Z(n6693) );
  AND U7204 ( .A(B[753]), .B(A[3]), .Z(n6687) );
  XNOR U7205 ( .A(n6677), .B(n6696), .Z(n6688) );
  XNOR U7206 ( .A(n6675), .B(n6678), .Z(n6696) );
  NAND U7207 ( .A(A[2]), .B(B[754]), .Z(n6678) );
  NANDN U7208 ( .A(n6697), .B(n6698), .Z(n6675) );
  AND U7209 ( .A(A[0]), .B(B[755]), .Z(n6698) );
  XOR U7210 ( .A(n6680), .B(n6699), .Z(n6677) );
  NAND U7211 ( .A(A[0]), .B(B[756]), .Z(n6699) );
  NAND U7212 ( .A(B[755]), .B(A[1]), .Z(n6680) );
  NAND U7213 ( .A(n6700), .B(n6701), .Z(n575) );
  NANDN U7214 ( .A(n6702), .B(n6703), .Z(n6701) );
  OR U7215 ( .A(n6704), .B(n6705), .Z(n6703) );
  NAND U7216 ( .A(n6705), .B(n6704), .Z(n6700) );
  XOR U7217 ( .A(n577), .B(n576), .Z(\A1[753] ) );
  XOR U7218 ( .A(n6705), .B(n6706), .Z(n576) );
  XNOR U7219 ( .A(n6704), .B(n6702), .Z(n6706) );
  AND U7220 ( .A(n6707), .B(n6708), .Z(n6702) );
  NANDN U7221 ( .A(n6709), .B(n6710), .Z(n6708) );
  NANDN U7222 ( .A(n6711), .B(n6712), .Z(n6710) );
  AND U7223 ( .A(B[752]), .B(A[3]), .Z(n6704) );
  XNOR U7224 ( .A(n6694), .B(n6713), .Z(n6705) );
  XNOR U7225 ( .A(n6692), .B(n6695), .Z(n6713) );
  NAND U7226 ( .A(A[2]), .B(B[753]), .Z(n6695) );
  NANDN U7227 ( .A(n6714), .B(n6715), .Z(n6692) );
  AND U7228 ( .A(A[0]), .B(B[754]), .Z(n6715) );
  XOR U7229 ( .A(n6697), .B(n6716), .Z(n6694) );
  NAND U7230 ( .A(A[0]), .B(B[755]), .Z(n6716) );
  NAND U7231 ( .A(B[754]), .B(A[1]), .Z(n6697) );
  NAND U7232 ( .A(n6717), .B(n6718), .Z(n577) );
  NANDN U7233 ( .A(n6719), .B(n6720), .Z(n6718) );
  OR U7234 ( .A(n6721), .B(n6722), .Z(n6720) );
  NAND U7235 ( .A(n6722), .B(n6721), .Z(n6717) );
  XOR U7236 ( .A(n579), .B(n578), .Z(\A1[752] ) );
  XOR U7237 ( .A(n6722), .B(n6723), .Z(n578) );
  XNOR U7238 ( .A(n6721), .B(n6719), .Z(n6723) );
  AND U7239 ( .A(n6724), .B(n6725), .Z(n6719) );
  NANDN U7240 ( .A(n6726), .B(n6727), .Z(n6725) );
  NANDN U7241 ( .A(n6728), .B(n6729), .Z(n6727) );
  AND U7242 ( .A(B[751]), .B(A[3]), .Z(n6721) );
  XNOR U7243 ( .A(n6711), .B(n6730), .Z(n6722) );
  XNOR U7244 ( .A(n6709), .B(n6712), .Z(n6730) );
  NAND U7245 ( .A(A[2]), .B(B[752]), .Z(n6712) );
  NANDN U7246 ( .A(n6731), .B(n6732), .Z(n6709) );
  AND U7247 ( .A(A[0]), .B(B[753]), .Z(n6732) );
  XOR U7248 ( .A(n6714), .B(n6733), .Z(n6711) );
  NAND U7249 ( .A(A[0]), .B(B[754]), .Z(n6733) );
  NAND U7250 ( .A(B[753]), .B(A[1]), .Z(n6714) );
  NAND U7251 ( .A(n6734), .B(n6735), .Z(n579) );
  NANDN U7252 ( .A(n6736), .B(n6737), .Z(n6735) );
  OR U7253 ( .A(n6738), .B(n6739), .Z(n6737) );
  NAND U7254 ( .A(n6739), .B(n6738), .Z(n6734) );
  XOR U7255 ( .A(n581), .B(n580), .Z(\A1[751] ) );
  XOR U7256 ( .A(n6739), .B(n6740), .Z(n580) );
  XNOR U7257 ( .A(n6738), .B(n6736), .Z(n6740) );
  AND U7258 ( .A(n6741), .B(n6742), .Z(n6736) );
  NANDN U7259 ( .A(n6743), .B(n6744), .Z(n6742) );
  NANDN U7260 ( .A(n6745), .B(n6746), .Z(n6744) );
  AND U7261 ( .A(B[750]), .B(A[3]), .Z(n6738) );
  XNOR U7262 ( .A(n6728), .B(n6747), .Z(n6739) );
  XNOR U7263 ( .A(n6726), .B(n6729), .Z(n6747) );
  NAND U7264 ( .A(A[2]), .B(B[751]), .Z(n6729) );
  NANDN U7265 ( .A(n6748), .B(n6749), .Z(n6726) );
  AND U7266 ( .A(A[0]), .B(B[752]), .Z(n6749) );
  XOR U7267 ( .A(n6731), .B(n6750), .Z(n6728) );
  NAND U7268 ( .A(A[0]), .B(B[753]), .Z(n6750) );
  NAND U7269 ( .A(B[752]), .B(A[1]), .Z(n6731) );
  NAND U7270 ( .A(n6751), .B(n6752), .Z(n581) );
  NANDN U7271 ( .A(n6753), .B(n6754), .Z(n6752) );
  OR U7272 ( .A(n6755), .B(n6756), .Z(n6754) );
  NAND U7273 ( .A(n6756), .B(n6755), .Z(n6751) );
  XOR U7274 ( .A(n583), .B(n582), .Z(\A1[750] ) );
  XOR U7275 ( .A(n6756), .B(n6757), .Z(n582) );
  XNOR U7276 ( .A(n6755), .B(n6753), .Z(n6757) );
  AND U7277 ( .A(n6758), .B(n6759), .Z(n6753) );
  NANDN U7278 ( .A(n6760), .B(n6761), .Z(n6759) );
  NANDN U7279 ( .A(n6762), .B(n6763), .Z(n6761) );
  AND U7280 ( .A(B[749]), .B(A[3]), .Z(n6755) );
  XNOR U7281 ( .A(n6745), .B(n6764), .Z(n6756) );
  XNOR U7282 ( .A(n6743), .B(n6746), .Z(n6764) );
  NAND U7283 ( .A(A[2]), .B(B[750]), .Z(n6746) );
  NANDN U7284 ( .A(n6765), .B(n6766), .Z(n6743) );
  AND U7285 ( .A(A[0]), .B(B[751]), .Z(n6766) );
  XOR U7286 ( .A(n6748), .B(n6767), .Z(n6745) );
  NAND U7287 ( .A(A[0]), .B(B[752]), .Z(n6767) );
  NAND U7288 ( .A(B[751]), .B(A[1]), .Z(n6748) );
  NAND U7289 ( .A(n6768), .B(n6769), .Z(n583) );
  NANDN U7290 ( .A(n6770), .B(n6771), .Z(n6769) );
  OR U7291 ( .A(n6772), .B(n6773), .Z(n6771) );
  NAND U7292 ( .A(n6773), .B(n6772), .Z(n6768) );
  XOR U7293 ( .A(n565), .B(n564), .Z(\A1[74] ) );
  XOR U7294 ( .A(n6603), .B(n6774), .Z(n564) );
  XNOR U7295 ( .A(n6602), .B(n6600), .Z(n6774) );
  AND U7296 ( .A(n6775), .B(n6776), .Z(n6600) );
  NANDN U7297 ( .A(n6777), .B(n6778), .Z(n6776) );
  NANDN U7298 ( .A(n6779), .B(n6780), .Z(n6778) );
  AND U7299 ( .A(B[73]), .B(A[3]), .Z(n6602) );
  XNOR U7300 ( .A(n6592), .B(n6781), .Z(n6603) );
  XNOR U7301 ( .A(n6590), .B(n6593), .Z(n6781) );
  NAND U7302 ( .A(A[2]), .B(B[74]), .Z(n6593) );
  NANDN U7303 ( .A(n6782), .B(n6783), .Z(n6590) );
  AND U7304 ( .A(A[0]), .B(B[75]), .Z(n6783) );
  XOR U7305 ( .A(n6595), .B(n6784), .Z(n6592) );
  NAND U7306 ( .A(A[0]), .B(B[76]), .Z(n6784) );
  NAND U7307 ( .A(B[75]), .B(A[1]), .Z(n6595) );
  NAND U7308 ( .A(n6785), .B(n6786), .Z(n565) );
  NANDN U7309 ( .A(n6787), .B(n6788), .Z(n6786) );
  OR U7310 ( .A(n6789), .B(n6790), .Z(n6788) );
  NAND U7311 ( .A(n6790), .B(n6789), .Z(n6785) );
  XOR U7312 ( .A(n585), .B(n584), .Z(\A1[749] ) );
  XOR U7313 ( .A(n6773), .B(n6791), .Z(n584) );
  XNOR U7314 ( .A(n6772), .B(n6770), .Z(n6791) );
  AND U7315 ( .A(n6792), .B(n6793), .Z(n6770) );
  NANDN U7316 ( .A(n6794), .B(n6795), .Z(n6793) );
  NANDN U7317 ( .A(n6796), .B(n6797), .Z(n6795) );
  AND U7318 ( .A(B[748]), .B(A[3]), .Z(n6772) );
  XNOR U7319 ( .A(n6762), .B(n6798), .Z(n6773) );
  XNOR U7320 ( .A(n6760), .B(n6763), .Z(n6798) );
  NAND U7321 ( .A(A[2]), .B(B[749]), .Z(n6763) );
  NANDN U7322 ( .A(n6799), .B(n6800), .Z(n6760) );
  AND U7323 ( .A(A[0]), .B(B[750]), .Z(n6800) );
  XOR U7324 ( .A(n6765), .B(n6801), .Z(n6762) );
  NAND U7325 ( .A(A[0]), .B(B[751]), .Z(n6801) );
  NAND U7326 ( .A(B[750]), .B(A[1]), .Z(n6765) );
  NAND U7327 ( .A(n6802), .B(n6803), .Z(n585) );
  NANDN U7328 ( .A(n6804), .B(n6805), .Z(n6803) );
  OR U7329 ( .A(n6806), .B(n6807), .Z(n6805) );
  NAND U7330 ( .A(n6807), .B(n6806), .Z(n6802) );
  XOR U7331 ( .A(n589), .B(n588), .Z(\A1[748] ) );
  XOR U7332 ( .A(n6807), .B(n6808), .Z(n588) );
  XNOR U7333 ( .A(n6806), .B(n6804), .Z(n6808) );
  AND U7334 ( .A(n6809), .B(n6810), .Z(n6804) );
  NANDN U7335 ( .A(n6811), .B(n6812), .Z(n6810) );
  NANDN U7336 ( .A(n6813), .B(n6814), .Z(n6812) );
  AND U7337 ( .A(B[747]), .B(A[3]), .Z(n6806) );
  XNOR U7338 ( .A(n6796), .B(n6815), .Z(n6807) );
  XNOR U7339 ( .A(n6794), .B(n6797), .Z(n6815) );
  NAND U7340 ( .A(A[2]), .B(B[748]), .Z(n6797) );
  NANDN U7341 ( .A(n6816), .B(n6817), .Z(n6794) );
  AND U7342 ( .A(A[0]), .B(B[749]), .Z(n6817) );
  XOR U7343 ( .A(n6799), .B(n6818), .Z(n6796) );
  NAND U7344 ( .A(A[0]), .B(B[750]), .Z(n6818) );
  NAND U7345 ( .A(B[749]), .B(A[1]), .Z(n6799) );
  NAND U7346 ( .A(n6819), .B(n6820), .Z(n589) );
  NANDN U7347 ( .A(n6821), .B(n6822), .Z(n6820) );
  OR U7348 ( .A(n6823), .B(n6824), .Z(n6822) );
  NAND U7349 ( .A(n6824), .B(n6823), .Z(n6819) );
  XOR U7350 ( .A(n591), .B(n590), .Z(\A1[747] ) );
  XOR U7351 ( .A(n6824), .B(n6825), .Z(n590) );
  XNOR U7352 ( .A(n6823), .B(n6821), .Z(n6825) );
  AND U7353 ( .A(n6826), .B(n6827), .Z(n6821) );
  NANDN U7354 ( .A(n6828), .B(n6829), .Z(n6827) );
  NANDN U7355 ( .A(n6830), .B(n6831), .Z(n6829) );
  AND U7356 ( .A(B[746]), .B(A[3]), .Z(n6823) );
  XNOR U7357 ( .A(n6813), .B(n6832), .Z(n6824) );
  XNOR U7358 ( .A(n6811), .B(n6814), .Z(n6832) );
  NAND U7359 ( .A(A[2]), .B(B[747]), .Z(n6814) );
  NANDN U7360 ( .A(n6833), .B(n6834), .Z(n6811) );
  AND U7361 ( .A(A[0]), .B(B[748]), .Z(n6834) );
  XOR U7362 ( .A(n6816), .B(n6835), .Z(n6813) );
  NAND U7363 ( .A(A[0]), .B(B[749]), .Z(n6835) );
  NAND U7364 ( .A(B[748]), .B(A[1]), .Z(n6816) );
  NAND U7365 ( .A(n6836), .B(n6837), .Z(n591) );
  NANDN U7366 ( .A(n6838), .B(n6839), .Z(n6837) );
  OR U7367 ( .A(n6840), .B(n6841), .Z(n6839) );
  NAND U7368 ( .A(n6841), .B(n6840), .Z(n6836) );
  XOR U7369 ( .A(n593), .B(n592), .Z(\A1[746] ) );
  XOR U7370 ( .A(n6841), .B(n6842), .Z(n592) );
  XNOR U7371 ( .A(n6840), .B(n6838), .Z(n6842) );
  AND U7372 ( .A(n6843), .B(n6844), .Z(n6838) );
  NANDN U7373 ( .A(n6845), .B(n6846), .Z(n6844) );
  NANDN U7374 ( .A(n6847), .B(n6848), .Z(n6846) );
  AND U7375 ( .A(B[745]), .B(A[3]), .Z(n6840) );
  XNOR U7376 ( .A(n6830), .B(n6849), .Z(n6841) );
  XNOR U7377 ( .A(n6828), .B(n6831), .Z(n6849) );
  NAND U7378 ( .A(A[2]), .B(B[746]), .Z(n6831) );
  NANDN U7379 ( .A(n6850), .B(n6851), .Z(n6828) );
  AND U7380 ( .A(A[0]), .B(B[747]), .Z(n6851) );
  XOR U7381 ( .A(n6833), .B(n6852), .Z(n6830) );
  NAND U7382 ( .A(A[0]), .B(B[748]), .Z(n6852) );
  NAND U7383 ( .A(B[747]), .B(A[1]), .Z(n6833) );
  NAND U7384 ( .A(n6853), .B(n6854), .Z(n593) );
  NANDN U7385 ( .A(n6855), .B(n6856), .Z(n6854) );
  OR U7386 ( .A(n6857), .B(n6858), .Z(n6856) );
  NAND U7387 ( .A(n6858), .B(n6857), .Z(n6853) );
  XOR U7388 ( .A(n595), .B(n594), .Z(\A1[745] ) );
  XOR U7389 ( .A(n6858), .B(n6859), .Z(n594) );
  XNOR U7390 ( .A(n6857), .B(n6855), .Z(n6859) );
  AND U7391 ( .A(n6860), .B(n6861), .Z(n6855) );
  NANDN U7392 ( .A(n6862), .B(n6863), .Z(n6861) );
  NANDN U7393 ( .A(n6864), .B(n6865), .Z(n6863) );
  AND U7394 ( .A(B[744]), .B(A[3]), .Z(n6857) );
  XNOR U7395 ( .A(n6847), .B(n6866), .Z(n6858) );
  XNOR U7396 ( .A(n6845), .B(n6848), .Z(n6866) );
  NAND U7397 ( .A(A[2]), .B(B[745]), .Z(n6848) );
  NANDN U7398 ( .A(n6867), .B(n6868), .Z(n6845) );
  AND U7399 ( .A(A[0]), .B(B[746]), .Z(n6868) );
  XOR U7400 ( .A(n6850), .B(n6869), .Z(n6847) );
  NAND U7401 ( .A(A[0]), .B(B[747]), .Z(n6869) );
  NAND U7402 ( .A(B[746]), .B(A[1]), .Z(n6850) );
  NAND U7403 ( .A(n6870), .B(n6871), .Z(n595) );
  NANDN U7404 ( .A(n6872), .B(n6873), .Z(n6871) );
  OR U7405 ( .A(n6874), .B(n6875), .Z(n6873) );
  NAND U7406 ( .A(n6875), .B(n6874), .Z(n6870) );
  XOR U7407 ( .A(n597), .B(n596), .Z(\A1[744] ) );
  XOR U7408 ( .A(n6875), .B(n6876), .Z(n596) );
  XNOR U7409 ( .A(n6874), .B(n6872), .Z(n6876) );
  AND U7410 ( .A(n6877), .B(n6878), .Z(n6872) );
  NANDN U7411 ( .A(n6879), .B(n6880), .Z(n6878) );
  NANDN U7412 ( .A(n6881), .B(n6882), .Z(n6880) );
  AND U7413 ( .A(B[743]), .B(A[3]), .Z(n6874) );
  XNOR U7414 ( .A(n6864), .B(n6883), .Z(n6875) );
  XNOR U7415 ( .A(n6862), .B(n6865), .Z(n6883) );
  NAND U7416 ( .A(A[2]), .B(B[744]), .Z(n6865) );
  NANDN U7417 ( .A(n6884), .B(n6885), .Z(n6862) );
  AND U7418 ( .A(A[0]), .B(B[745]), .Z(n6885) );
  XOR U7419 ( .A(n6867), .B(n6886), .Z(n6864) );
  NAND U7420 ( .A(A[0]), .B(B[746]), .Z(n6886) );
  NAND U7421 ( .A(B[745]), .B(A[1]), .Z(n6867) );
  NAND U7422 ( .A(n6887), .B(n6888), .Z(n597) );
  NANDN U7423 ( .A(n6889), .B(n6890), .Z(n6888) );
  OR U7424 ( .A(n6891), .B(n6892), .Z(n6890) );
  NAND U7425 ( .A(n6892), .B(n6891), .Z(n6887) );
  XOR U7426 ( .A(n599), .B(n598), .Z(\A1[743] ) );
  XOR U7427 ( .A(n6892), .B(n6893), .Z(n598) );
  XNOR U7428 ( .A(n6891), .B(n6889), .Z(n6893) );
  AND U7429 ( .A(n6894), .B(n6895), .Z(n6889) );
  NANDN U7430 ( .A(n6896), .B(n6897), .Z(n6895) );
  NANDN U7431 ( .A(n6898), .B(n6899), .Z(n6897) );
  AND U7432 ( .A(B[742]), .B(A[3]), .Z(n6891) );
  XNOR U7433 ( .A(n6881), .B(n6900), .Z(n6892) );
  XNOR U7434 ( .A(n6879), .B(n6882), .Z(n6900) );
  NAND U7435 ( .A(A[2]), .B(B[743]), .Z(n6882) );
  NANDN U7436 ( .A(n6901), .B(n6902), .Z(n6879) );
  AND U7437 ( .A(A[0]), .B(B[744]), .Z(n6902) );
  XOR U7438 ( .A(n6884), .B(n6903), .Z(n6881) );
  NAND U7439 ( .A(A[0]), .B(B[745]), .Z(n6903) );
  NAND U7440 ( .A(B[744]), .B(A[1]), .Z(n6884) );
  NAND U7441 ( .A(n6904), .B(n6905), .Z(n599) );
  NANDN U7442 ( .A(n6906), .B(n6907), .Z(n6905) );
  OR U7443 ( .A(n6908), .B(n6909), .Z(n6907) );
  NAND U7444 ( .A(n6909), .B(n6908), .Z(n6904) );
  XOR U7445 ( .A(n601), .B(n600), .Z(\A1[742] ) );
  XOR U7446 ( .A(n6909), .B(n6910), .Z(n600) );
  XNOR U7447 ( .A(n6908), .B(n6906), .Z(n6910) );
  AND U7448 ( .A(n6911), .B(n6912), .Z(n6906) );
  NANDN U7449 ( .A(n6913), .B(n6914), .Z(n6912) );
  NANDN U7450 ( .A(n6915), .B(n6916), .Z(n6914) );
  AND U7451 ( .A(B[741]), .B(A[3]), .Z(n6908) );
  XNOR U7452 ( .A(n6898), .B(n6917), .Z(n6909) );
  XNOR U7453 ( .A(n6896), .B(n6899), .Z(n6917) );
  NAND U7454 ( .A(A[2]), .B(B[742]), .Z(n6899) );
  NANDN U7455 ( .A(n6918), .B(n6919), .Z(n6896) );
  AND U7456 ( .A(A[0]), .B(B[743]), .Z(n6919) );
  XOR U7457 ( .A(n6901), .B(n6920), .Z(n6898) );
  NAND U7458 ( .A(A[0]), .B(B[744]), .Z(n6920) );
  NAND U7459 ( .A(B[743]), .B(A[1]), .Z(n6901) );
  NAND U7460 ( .A(n6921), .B(n6922), .Z(n601) );
  NANDN U7461 ( .A(n6923), .B(n6924), .Z(n6922) );
  OR U7462 ( .A(n6925), .B(n6926), .Z(n6924) );
  NAND U7463 ( .A(n6926), .B(n6925), .Z(n6921) );
  XOR U7464 ( .A(n603), .B(n602), .Z(\A1[741] ) );
  XOR U7465 ( .A(n6926), .B(n6927), .Z(n602) );
  XNOR U7466 ( .A(n6925), .B(n6923), .Z(n6927) );
  AND U7467 ( .A(n6928), .B(n6929), .Z(n6923) );
  NANDN U7468 ( .A(n6930), .B(n6931), .Z(n6929) );
  NANDN U7469 ( .A(n6932), .B(n6933), .Z(n6931) );
  AND U7470 ( .A(B[740]), .B(A[3]), .Z(n6925) );
  XNOR U7471 ( .A(n6915), .B(n6934), .Z(n6926) );
  XNOR U7472 ( .A(n6913), .B(n6916), .Z(n6934) );
  NAND U7473 ( .A(A[2]), .B(B[741]), .Z(n6916) );
  NANDN U7474 ( .A(n6935), .B(n6936), .Z(n6913) );
  AND U7475 ( .A(A[0]), .B(B[742]), .Z(n6936) );
  XOR U7476 ( .A(n6918), .B(n6937), .Z(n6915) );
  NAND U7477 ( .A(A[0]), .B(B[743]), .Z(n6937) );
  NAND U7478 ( .A(B[742]), .B(A[1]), .Z(n6918) );
  NAND U7479 ( .A(n6938), .B(n6939), .Z(n603) );
  NANDN U7480 ( .A(n6940), .B(n6941), .Z(n6939) );
  OR U7481 ( .A(n6942), .B(n6943), .Z(n6941) );
  NAND U7482 ( .A(n6943), .B(n6942), .Z(n6938) );
  XOR U7483 ( .A(n605), .B(n604), .Z(\A1[740] ) );
  XOR U7484 ( .A(n6943), .B(n6944), .Z(n604) );
  XNOR U7485 ( .A(n6942), .B(n6940), .Z(n6944) );
  AND U7486 ( .A(n6945), .B(n6946), .Z(n6940) );
  NANDN U7487 ( .A(n6947), .B(n6948), .Z(n6946) );
  NANDN U7488 ( .A(n6949), .B(n6950), .Z(n6948) );
  AND U7489 ( .A(B[739]), .B(A[3]), .Z(n6942) );
  XNOR U7490 ( .A(n6932), .B(n6951), .Z(n6943) );
  XNOR U7491 ( .A(n6930), .B(n6933), .Z(n6951) );
  NAND U7492 ( .A(A[2]), .B(B[740]), .Z(n6933) );
  NANDN U7493 ( .A(n6952), .B(n6953), .Z(n6930) );
  AND U7494 ( .A(A[0]), .B(B[741]), .Z(n6953) );
  XOR U7495 ( .A(n6935), .B(n6954), .Z(n6932) );
  NAND U7496 ( .A(A[0]), .B(B[742]), .Z(n6954) );
  NAND U7497 ( .A(B[741]), .B(A[1]), .Z(n6935) );
  NAND U7498 ( .A(n6955), .B(n6956), .Z(n605) );
  NANDN U7499 ( .A(n6957), .B(n6958), .Z(n6956) );
  OR U7500 ( .A(n6959), .B(n6960), .Z(n6958) );
  NAND U7501 ( .A(n6960), .B(n6959), .Z(n6955) );
  XOR U7502 ( .A(n587), .B(n586), .Z(\A1[73] ) );
  XOR U7503 ( .A(n6790), .B(n6961), .Z(n586) );
  XNOR U7504 ( .A(n6789), .B(n6787), .Z(n6961) );
  AND U7505 ( .A(n6962), .B(n6963), .Z(n6787) );
  NANDN U7506 ( .A(n6964), .B(n6965), .Z(n6963) );
  NANDN U7507 ( .A(n6966), .B(n6967), .Z(n6965) );
  AND U7508 ( .A(B[72]), .B(A[3]), .Z(n6789) );
  XNOR U7509 ( .A(n6779), .B(n6968), .Z(n6790) );
  XNOR U7510 ( .A(n6777), .B(n6780), .Z(n6968) );
  NAND U7511 ( .A(A[2]), .B(B[73]), .Z(n6780) );
  NANDN U7512 ( .A(n6969), .B(n6970), .Z(n6777) );
  AND U7513 ( .A(A[0]), .B(B[74]), .Z(n6970) );
  XOR U7514 ( .A(n6782), .B(n6971), .Z(n6779) );
  NAND U7515 ( .A(A[0]), .B(B[75]), .Z(n6971) );
  NAND U7516 ( .A(B[74]), .B(A[1]), .Z(n6782) );
  NAND U7517 ( .A(n6972), .B(n6973), .Z(n587) );
  NANDN U7518 ( .A(n6974), .B(n6975), .Z(n6973) );
  OR U7519 ( .A(n6976), .B(n6977), .Z(n6975) );
  NAND U7520 ( .A(n6977), .B(n6976), .Z(n6972) );
  XOR U7521 ( .A(n607), .B(n606), .Z(\A1[739] ) );
  XOR U7522 ( .A(n6960), .B(n6978), .Z(n606) );
  XNOR U7523 ( .A(n6959), .B(n6957), .Z(n6978) );
  AND U7524 ( .A(n6979), .B(n6980), .Z(n6957) );
  NANDN U7525 ( .A(n6981), .B(n6982), .Z(n6980) );
  NANDN U7526 ( .A(n6983), .B(n6984), .Z(n6982) );
  AND U7527 ( .A(B[738]), .B(A[3]), .Z(n6959) );
  XNOR U7528 ( .A(n6949), .B(n6985), .Z(n6960) );
  XNOR U7529 ( .A(n6947), .B(n6950), .Z(n6985) );
  NAND U7530 ( .A(A[2]), .B(B[739]), .Z(n6950) );
  NANDN U7531 ( .A(n6986), .B(n6987), .Z(n6947) );
  AND U7532 ( .A(A[0]), .B(B[740]), .Z(n6987) );
  XOR U7533 ( .A(n6952), .B(n6988), .Z(n6949) );
  NAND U7534 ( .A(A[0]), .B(B[741]), .Z(n6988) );
  NAND U7535 ( .A(B[740]), .B(A[1]), .Z(n6952) );
  NAND U7536 ( .A(n6989), .B(n6990), .Z(n607) );
  NANDN U7537 ( .A(n6991), .B(n6992), .Z(n6990) );
  OR U7538 ( .A(n6993), .B(n6994), .Z(n6992) );
  NAND U7539 ( .A(n6994), .B(n6993), .Z(n6989) );
  XOR U7540 ( .A(n611), .B(n610), .Z(\A1[738] ) );
  XOR U7541 ( .A(n6994), .B(n6995), .Z(n610) );
  XNOR U7542 ( .A(n6993), .B(n6991), .Z(n6995) );
  AND U7543 ( .A(n6996), .B(n6997), .Z(n6991) );
  NANDN U7544 ( .A(n6998), .B(n6999), .Z(n6997) );
  NANDN U7545 ( .A(n7000), .B(n7001), .Z(n6999) );
  AND U7546 ( .A(B[737]), .B(A[3]), .Z(n6993) );
  XNOR U7547 ( .A(n6983), .B(n7002), .Z(n6994) );
  XNOR U7548 ( .A(n6981), .B(n6984), .Z(n7002) );
  NAND U7549 ( .A(A[2]), .B(B[738]), .Z(n6984) );
  NANDN U7550 ( .A(n7003), .B(n7004), .Z(n6981) );
  AND U7551 ( .A(A[0]), .B(B[739]), .Z(n7004) );
  XOR U7552 ( .A(n6986), .B(n7005), .Z(n6983) );
  NAND U7553 ( .A(A[0]), .B(B[740]), .Z(n7005) );
  NAND U7554 ( .A(B[739]), .B(A[1]), .Z(n6986) );
  NAND U7555 ( .A(n7006), .B(n7007), .Z(n611) );
  NANDN U7556 ( .A(n7008), .B(n7009), .Z(n7007) );
  OR U7557 ( .A(n7010), .B(n7011), .Z(n7009) );
  NAND U7558 ( .A(n7011), .B(n7010), .Z(n7006) );
  XOR U7559 ( .A(n613), .B(n612), .Z(\A1[737] ) );
  XOR U7560 ( .A(n7011), .B(n7012), .Z(n612) );
  XNOR U7561 ( .A(n7010), .B(n7008), .Z(n7012) );
  AND U7562 ( .A(n7013), .B(n7014), .Z(n7008) );
  NANDN U7563 ( .A(n7015), .B(n7016), .Z(n7014) );
  NANDN U7564 ( .A(n7017), .B(n7018), .Z(n7016) );
  AND U7565 ( .A(B[736]), .B(A[3]), .Z(n7010) );
  XNOR U7566 ( .A(n7000), .B(n7019), .Z(n7011) );
  XNOR U7567 ( .A(n6998), .B(n7001), .Z(n7019) );
  NAND U7568 ( .A(A[2]), .B(B[737]), .Z(n7001) );
  NANDN U7569 ( .A(n7020), .B(n7021), .Z(n6998) );
  AND U7570 ( .A(A[0]), .B(B[738]), .Z(n7021) );
  XOR U7571 ( .A(n7003), .B(n7022), .Z(n7000) );
  NAND U7572 ( .A(A[0]), .B(B[739]), .Z(n7022) );
  NAND U7573 ( .A(B[738]), .B(A[1]), .Z(n7003) );
  NAND U7574 ( .A(n7023), .B(n7024), .Z(n613) );
  NANDN U7575 ( .A(n7025), .B(n7026), .Z(n7024) );
  OR U7576 ( .A(n7027), .B(n7028), .Z(n7026) );
  NAND U7577 ( .A(n7028), .B(n7027), .Z(n7023) );
  XOR U7578 ( .A(n615), .B(n614), .Z(\A1[736] ) );
  XOR U7579 ( .A(n7028), .B(n7029), .Z(n614) );
  XNOR U7580 ( .A(n7027), .B(n7025), .Z(n7029) );
  AND U7581 ( .A(n7030), .B(n7031), .Z(n7025) );
  NANDN U7582 ( .A(n7032), .B(n7033), .Z(n7031) );
  NANDN U7583 ( .A(n7034), .B(n7035), .Z(n7033) );
  AND U7584 ( .A(B[735]), .B(A[3]), .Z(n7027) );
  XNOR U7585 ( .A(n7017), .B(n7036), .Z(n7028) );
  XNOR U7586 ( .A(n7015), .B(n7018), .Z(n7036) );
  NAND U7587 ( .A(A[2]), .B(B[736]), .Z(n7018) );
  NANDN U7588 ( .A(n7037), .B(n7038), .Z(n7015) );
  AND U7589 ( .A(A[0]), .B(B[737]), .Z(n7038) );
  XOR U7590 ( .A(n7020), .B(n7039), .Z(n7017) );
  NAND U7591 ( .A(A[0]), .B(B[738]), .Z(n7039) );
  NAND U7592 ( .A(B[737]), .B(A[1]), .Z(n7020) );
  NAND U7593 ( .A(n7040), .B(n7041), .Z(n615) );
  NANDN U7594 ( .A(n7042), .B(n7043), .Z(n7041) );
  OR U7595 ( .A(n7044), .B(n7045), .Z(n7043) );
  NAND U7596 ( .A(n7045), .B(n7044), .Z(n7040) );
  XOR U7597 ( .A(n617), .B(n616), .Z(\A1[735] ) );
  XOR U7598 ( .A(n7045), .B(n7046), .Z(n616) );
  XNOR U7599 ( .A(n7044), .B(n7042), .Z(n7046) );
  AND U7600 ( .A(n7047), .B(n7048), .Z(n7042) );
  NANDN U7601 ( .A(n7049), .B(n7050), .Z(n7048) );
  NANDN U7602 ( .A(n7051), .B(n7052), .Z(n7050) );
  AND U7603 ( .A(B[734]), .B(A[3]), .Z(n7044) );
  XNOR U7604 ( .A(n7034), .B(n7053), .Z(n7045) );
  XNOR U7605 ( .A(n7032), .B(n7035), .Z(n7053) );
  NAND U7606 ( .A(A[2]), .B(B[735]), .Z(n7035) );
  NANDN U7607 ( .A(n7054), .B(n7055), .Z(n7032) );
  AND U7608 ( .A(A[0]), .B(B[736]), .Z(n7055) );
  XOR U7609 ( .A(n7037), .B(n7056), .Z(n7034) );
  NAND U7610 ( .A(A[0]), .B(B[737]), .Z(n7056) );
  NAND U7611 ( .A(B[736]), .B(A[1]), .Z(n7037) );
  NAND U7612 ( .A(n7057), .B(n7058), .Z(n617) );
  NANDN U7613 ( .A(n7059), .B(n7060), .Z(n7058) );
  OR U7614 ( .A(n7061), .B(n7062), .Z(n7060) );
  NAND U7615 ( .A(n7062), .B(n7061), .Z(n7057) );
  XOR U7616 ( .A(n619), .B(n618), .Z(\A1[734] ) );
  XOR U7617 ( .A(n7062), .B(n7063), .Z(n618) );
  XNOR U7618 ( .A(n7061), .B(n7059), .Z(n7063) );
  AND U7619 ( .A(n7064), .B(n7065), .Z(n7059) );
  NANDN U7620 ( .A(n7066), .B(n7067), .Z(n7065) );
  NANDN U7621 ( .A(n7068), .B(n7069), .Z(n7067) );
  AND U7622 ( .A(B[733]), .B(A[3]), .Z(n7061) );
  XNOR U7623 ( .A(n7051), .B(n7070), .Z(n7062) );
  XNOR U7624 ( .A(n7049), .B(n7052), .Z(n7070) );
  NAND U7625 ( .A(A[2]), .B(B[734]), .Z(n7052) );
  NANDN U7626 ( .A(n7071), .B(n7072), .Z(n7049) );
  AND U7627 ( .A(A[0]), .B(B[735]), .Z(n7072) );
  XOR U7628 ( .A(n7054), .B(n7073), .Z(n7051) );
  NAND U7629 ( .A(A[0]), .B(B[736]), .Z(n7073) );
  NAND U7630 ( .A(B[735]), .B(A[1]), .Z(n7054) );
  NAND U7631 ( .A(n7074), .B(n7075), .Z(n619) );
  NANDN U7632 ( .A(n7076), .B(n7077), .Z(n7075) );
  OR U7633 ( .A(n7078), .B(n7079), .Z(n7077) );
  NAND U7634 ( .A(n7079), .B(n7078), .Z(n7074) );
  XOR U7635 ( .A(n621), .B(n620), .Z(\A1[733] ) );
  XOR U7636 ( .A(n7079), .B(n7080), .Z(n620) );
  XNOR U7637 ( .A(n7078), .B(n7076), .Z(n7080) );
  AND U7638 ( .A(n7081), .B(n7082), .Z(n7076) );
  NANDN U7639 ( .A(n7083), .B(n7084), .Z(n7082) );
  NANDN U7640 ( .A(n7085), .B(n7086), .Z(n7084) );
  AND U7641 ( .A(B[732]), .B(A[3]), .Z(n7078) );
  XNOR U7642 ( .A(n7068), .B(n7087), .Z(n7079) );
  XNOR U7643 ( .A(n7066), .B(n7069), .Z(n7087) );
  NAND U7644 ( .A(A[2]), .B(B[733]), .Z(n7069) );
  NANDN U7645 ( .A(n7088), .B(n7089), .Z(n7066) );
  AND U7646 ( .A(A[0]), .B(B[734]), .Z(n7089) );
  XOR U7647 ( .A(n7071), .B(n7090), .Z(n7068) );
  NAND U7648 ( .A(A[0]), .B(B[735]), .Z(n7090) );
  NAND U7649 ( .A(B[734]), .B(A[1]), .Z(n7071) );
  NAND U7650 ( .A(n7091), .B(n7092), .Z(n621) );
  NANDN U7651 ( .A(n7093), .B(n7094), .Z(n7092) );
  OR U7652 ( .A(n7095), .B(n7096), .Z(n7094) );
  NAND U7653 ( .A(n7096), .B(n7095), .Z(n7091) );
  XOR U7654 ( .A(n623), .B(n622), .Z(\A1[732] ) );
  XOR U7655 ( .A(n7096), .B(n7097), .Z(n622) );
  XNOR U7656 ( .A(n7095), .B(n7093), .Z(n7097) );
  AND U7657 ( .A(n7098), .B(n7099), .Z(n7093) );
  NANDN U7658 ( .A(n7100), .B(n7101), .Z(n7099) );
  NANDN U7659 ( .A(n7102), .B(n7103), .Z(n7101) );
  AND U7660 ( .A(B[731]), .B(A[3]), .Z(n7095) );
  XNOR U7661 ( .A(n7085), .B(n7104), .Z(n7096) );
  XNOR U7662 ( .A(n7083), .B(n7086), .Z(n7104) );
  NAND U7663 ( .A(A[2]), .B(B[732]), .Z(n7086) );
  NANDN U7664 ( .A(n7105), .B(n7106), .Z(n7083) );
  AND U7665 ( .A(A[0]), .B(B[733]), .Z(n7106) );
  XOR U7666 ( .A(n7088), .B(n7107), .Z(n7085) );
  NAND U7667 ( .A(A[0]), .B(B[734]), .Z(n7107) );
  NAND U7668 ( .A(B[733]), .B(A[1]), .Z(n7088) );
  NAND U7669 ( .A(n7108), .B(n7109), .Z(n623) );
  NANDN U7670 ( .A(n7110), .B(n7111), .Z(n7109) );
  OR U7671 ( .A(n7112), .B(n7113), .Z(n7111) );
  NAND U7672 ( .A(n7113), .B(n7112), .Z(n7108) );
  XOR U7673 ( .A(n625), .B(n624), .Z(\A1[731] ) );
  XOR U7674 ( .A(n7113), .B(n7114), .Z(n624) );
  XNOR U7675 ( .A(n7112), .B(n7110), .Z(n7114) );
  AND U7676 ( .A(n7115), .B(n7116), .Z(n7110) );
  NANDN U7677 ( .A(n7117), .B(n7118), .Z(n7116) );
  NANDN U7678 ( .A(n7119), .B(n7120), .Z(n7118) );
  AND U7679 ( .A(B[730]), .B(A[3]), .Z(n7112) );
  XNOR U7680 ( .A(n7102), .B(n7121), .Z(n7113) );
  XNOR U7681 ( .A(n7100), .B(n7103), .Z(n7121) );
  NAND U7682 ( .A(A[2]), .B(B[731]), .Z(n7103) );
  NANDN U7683 ( .A(n7122), .B(n7123), .Z(n7100) );
  AND U7684 ( .A(A[0]), .B(B[732]), .Z(n7123) );
  XOR U7685 ( .A(n7105), .B(n7124), .Z(n7102) );
  NAND U7686 ( .A(A[0]), .B(B[733]), .Z(n7124) );
  NAND U7687 ( .A(B[732]), .B(A[1]), .Z(n7105) );
  NAND U7688 ( .A(n7125), .B(n7126), .Z(n625) );
  NANDN U7689 ( .A(n7127), .B(n7128), .Z(n7126) );
  OR U7690 ( .A(n7129), .B(n7130), .Z(n7128) );
  NAND U7691 ( .A(n7130), .B(n7129), .Z(n7125) );
  XOR U7692 ( .A(n627), .B(n626), .Z(\A1[730] ) );
  XOR U7693 ( .A(n7130), .B(n7131), .Z(n626) );
  XNOR U7694 ( .A(n7129), .B(n7127), .Z(n7131) );
  AND U7695 ( .A(n7132), .B(n7133), .Z(n7127) );
  NANDN U7696 ( .A(n7134), .B(n7135), .Z(n7133) );
  NANDN U7697 ( .A(n7136), .B(n7137), .Z(n7135) );
  AND U7698 ( .A(B[729]), .B(A[3]), .Z(n7129) );
  XNOR U7699 ( .A(n7119), .B(n7138), .Z(n7130) );
  XNOR U7700 ( .A(n7117), .B(n7120), .Z(n7138) );
  NAND U7701 ( .A(A[2]), .B(B[730]), .Z(n7120) );
  NANDN U7702 ( .A(n7139), .B(n7140), .Z(n7117) );
  AND U7703 ( .A(A[0]), .B(B[731]), .Z(n7140) );
  XOR U7704 ( .A(n7122), .B(n7141), .Z(n7119) );
  NAND U7705 ( .A(A[0]), .B(B[732]), .Z(n7141) );
  NAND U7706 ( .A(B[731]), .B(A[1]), .Z(n7122) );
  NAND U7707 ( .A(n7142), .B(n7143), .Z(n627) );
  NANDN U7708 ( .A(n7144), .B(n7145), .Z(n7143) );
  OR U7709 ( .A(n7146), .B(n7147), .Z(n7145) );
  NAND U7710 ( .A(n7147), .B(n7146), .Z(n7142) );
  XOR U7711 ( .A(n609), .B(n608), .Z(\A1[72] ) );
  XOR U7712 ( .A(n6977), .B(n7148), .Z(n608) );
  XNOR U7713 ( .A(n6976), .B(n6974), .Z(n7148) );
  AND U7714 ( .A(n7149), .B(n7150), .Z(n6974) );
  NANDN U7715 ( .A(n7151), .B(n7152), .Z(n7150) );
  NANDN U7716 ( .A(n7153), .B(n7154), .Z(n7152) );
  AND U7717 ( .A(B[71]), .B(A[3]), .Z(n6976) );
  XNOR U7718 ( .A(n6966), .B(n7155), .Z(n6977) );
  XNOR U7719 ( .A(n6964), .B(n6967), .Z(n7155) );
  NAND U7720 ( .A(A[2]), .B(B[72]), .Z(n6967) );
  NANDN U7721 ( .A(n7156), .B(n7157), .Z(n6964) );
  AND U7722 ( .A(A[0]), .B(B[73]), .Z(n7157) );
  XOR U7723 ( .A(n6969), .B(n7158), .Z(n6966) );
  NAND U7724 ( .A(A[0]), .B(B[74]), .Z(n7158) );
  NAND U7725 ( .A(B[73]), .B(A[1]), .Z(n6969) );
  NAND U7726 ( .A(n7159), .B(n7160), .Z(n609) );
  NANDN U7727 ( .A(n7161), .B(n7162), .Z(n7160) );
  OR U7728 ( .A(n7163), .B(n7164), .Z(n7162) );
  NAND U7729 ( .A(n7164), .B(n7163), .Z(n7159) );
  XOR U7730 ( .A(n629), .B(n628), .Z(\A1[729] ) );
  XOR U7731 ( .A(n7147), .B(n7165), .Z(n628) );
  XNOR U7732 ( .A(n7146), .B(n7144), .Z(n7165) );
  AND U7733 ( .A(n7166), .B(n7167), .Z(n7144) );
  NANDN U7734 ( .A(n7168), .B(n7169), .Z(n7167) );
  NANDN U7735 ( .A(n7170), .B(n7171), .Z(n7169) );
  AND U7736 ( .A(B[728]), .B(A[3]), .Z(n7146) );
  XNOR U7737 ( .A(n7136), .B(n7172), .Z(n7147) );
  XNOR U7738 ( .A(n7134), .B(n7137), .Z(n7172) );
  NAND U7739 ( .A(A[2]), .B(B[729]), .Z(n7137) );
  NANDN U7740 ( .A(n7173), .B(n7174), .Z(n7134) );
  AND U7741 ( .A(A[0]), .B(B[730]), .Z(n7174) );
  XOR U7742 ( .A(n7139), .B(n7175), .Z(n7136) );
  NAND U7743 ( .A(A[0]), .B(B[731]), .Z(n7175) );
  NAND U7744 ( .A(B[730]), .B(A[1]), .Z(n7139) );
  NAND U7745 ( .A(n7176), .B(n7177), .Z(n629) );
  NANDN U7746 ( .A(n7178), .B(n7179), .Z(n7177) );
  OR U7747 ( .A(n7180), .B(n7181), .Z(n7179) );
  NAND U7748 ( .A(n7181), .B(n7180), .Z(n7176) );
  XOR U7749 ( .A(n633), .B(n632), .Z(\A1[728] ) );
  XOR U7750 ( .A(n7181), .B(n7182), .Z(n632) );
  XNOR U7751 ( .A(n7180), .B(n7178), .Z(n7182) );
  AND U7752 ( .A(n7183), .B(n7184), .Z(n7178) );
  NANDN U7753 ( .A(n7185), .B(n7186), .Z(n7184) );
  NANDN U7754 ( .A(n7187), .B(n7188), .Z(n7186) );
  AND U7755 ( .A(B[727]), .B(A[3]), .Z(n7180) );
  XNOR U7756 ( .A(n7170), .B(n7189), .Z(n7181) );
  XNOR U7757 ( .A(n7168), .B(n7171), .Z(n7189) );
  NAND U7758 ( .A(A[2]), .B(B[728]), .Z(n7171) );
  NANDN U7759 ( .A(n7190), .B(n7191), .Z(n7168) );
  AND U7760 ( .A(A[0]), .B(B[729]), .Z(n7191) );
  XOR U7761 ( .A(n7173), .B(n7192), .Z(n7170) );
  NAND U7762 ( .A(A[0]), .B(B[730]), .Z(n7192) );
  NAND U7763 ( .A(B[729]), .B(A[1]), .Z(n7173) );
  NAND U7764 ( .A(n7193), .B(n7194), .Z(n633) );
  NANDN U7765 ( .A(n7195), .B(n7196), .Z(n7194) );
  OR U7766 ( .A(n7197), .B(n7198), .Z(n7196) );
  NAND U7767 ( .A(n7198), .B(n7197), .Z(n7193) );
  XOR U7768 ( .A(n635), .B(n634), .Z(\A1[727] ) );
  XOR U7769 ( .A(n7198), .B(n7199), .Z(n634) );
  XNOR U7770 ( .A(n7197), .B(n7195), .Z(n7199) );
  AND U7771 ( .A(n7200), .B(n7201), .Z(n7195) );
  NANDN U7772 ( .A(n7202), .B(n7203), .Z(n7201) );
  NANDN U7773 ( .A(n7204), .B(n7205), .Z(n7203) );
  AND U7774 ( .A(B[726]), .B(A[3]), .Z(n7197) );
  XNOR U7775 ( .A(n7187), .B(n7206), .Z(n7198) );
  XNOR U7776 ( .A(n7185), .B(n7188), .Z(n7206) );
  NAND U7777 ( .A(A[2]), .B(B[727]), .Z(n7188) );
  NANDN U7778 ( .A(n7207), .B(n7208), .Z(n7185) );
  AND U7779 ( .A(A[0]), .B(B[728]), .Z(n7208) );
  XOR U7780 ( .A(n7190), .B(n7209), .Z(n7187) );
  NAND U7781 ( .A(A[0]), .B(B[729]), .Z(n7209) );
  NAND U7782 ( .A(B[728]), .B(A[1]), .Z(n7190) );
  NAND U7783 ( .A(n7210), .B(n7211), .Z(n635) );
  NANDN U7784 ( .A(n7212), .B(n7213), .Z(n7211) );
  OR U7785 ( .A(n7214), .B(n7215), .Z(n7213) );
  NAND U7786 ( .A(n7215), .B(n7214), .Z(n7210) );
  XOR U7787 ( .A(n637), .B(n636), .Z(\A1[726] ) );
  XOR U7788 ( .A(n7215), .B(n7216), .Z(n636) );
  XNOR U7789 ( .A(n7214), .B(n7212), .Z(n7216) );
  AND U7790 ( .A(n7217), .B(n7218), .Z(n7212) );
  NANDN U7791 ( .A(n7219), .B(n7220), .Z(n7218) );
  NANDN U7792 ( .A(n7221), .B(n7222), .Z(n7220) );
  AND U7793 ( .A(B[725]), .B(A[3]), .Z(n7214) );
  XNOR U7794 ( .A(n7204), .B(n7223), .Z(n7215) );
  XNOR U7795 ( .A(n7202), .B(n7205), .Z(n7223) );
  NAND U7796 ( .A(A[2]), .B(B[726]), .Z(n7205) );
  NANDN U7797 ( .A(n7224), .B(n7225), .Z(n7202) );
  AND U7798 ( .A(A[0]), .B(B[727]), .Z(n7225) );
  XOR U7799 ( .A(n7207), .B(n7226), .Z(n7204) );
  NAND U7800 ( .A(A[0]), .B(B[728]), .Z(n7226) );
  NAND U7801 ( .A(B[727]), .B(A[1]), .Z(n7207) );
  NAND U7802 ( .A(n7227), .B(n7228), .Z(n637) );
  NANDN U7803 ( .A(n7229), .B(n7230), .Z(n7228) );
  OR U7804 ( .A(n7231), .B(n7232), .Z(n7230) );
  NAND U7805 ( .A(n7232), .B(n7231), .Z(n7227) );
  XOR U7806 ( .A(n639), .B(n638), .Z(\A1[725] ) );
  XOR U7807 ( .A(n7232), .B(n7233), .Z(n638) );
  XNOR U7808 ( .A(n7231), .B(n7229), .Z(n7233) );
  AND U7809 ( .A(n7234), .B(n7235), .Z(n7229) );
  NANDN U7810 ( .A(n7236), .B(n7237), .Z(n7235) );
  NANDN U7811 ( .A(n7238), .B(n7239), .Z(n7237) );
  AND U7812 ( .A(B[724]), .B(A[3]), .Z(n7231) );
  XNOR U7813 ( .A(n7221), .B(n7240), .Z(n7232) );
  XNOR U7814 ( .A(n7219), .B(n7222), .Z(n7240) );
  NAND U7815 ( .A(A[2]), .B(B[725]), .Z(n7222) );
  NANDN U7816 ( .A(n7241), .B(n7242), .Z(n7219) );
  AND U7817 ( .A(A[0]), .B(B[726]), .Z(n7242) );
  XOR U7818 ( .A(n7224), .B(n7243), .Z(n7221) );
  NAND U7819 ( .A(A[0]), .B(B[727]), .Z(n7243) );
  NAND U7820 ( .A(B[726]), .B(A[1]), .Z(n7224) );
  NAND U7821 ( .A(n7244), .B(n7245), .Z(n639) );
  NANDN U7822 ( .A(n7246), .B(n7247), .Z(n7245) );
  OR U7823 ( .A(n7248), .B(n7249), .Z(n7247) );
  NAND U7824 ( .A(n7249), .B(n7248), .Z(n7244) );
  XOR U7825 ( .A(n641), .B(n640), .Z(\A1[724] ) );
  XOR U7826 ( .A(n7249), .B(n7250), .Z(n640) );
  XNOR U7827 ( .A(n7248), .B(n7246), .Z(n7250) );
  AND U7828 ( .A(n7251), .B(n7252), .Z(n7246) );
  NANDN U7829 ( .A(n7253), .B(n7254), .Z(n7252) );
  NANDN U7830 ( .A(n7255), .B(n7256), .Z(n7254) );
  AND U7831 ( .A(B[723]), .B(A[3]), .Z(n7248) );
  XNOR U7832 ( .A(n7238), .B(n7257), .Z(n7249) );
  XNOR U7833 ( .A(n7236), .B(n7239), .Z(n7257) );
  NAND U7834 ( .A(A[2]), .B(B[724]), .Z(n7239) );
  NANDN U7835 ( .A(n7258), .B(n7259), .Z(n7236) );
  AND U7836 ( .A(A[0]), .B(B[725]), .Z(n7259) );
  XOR U7837 ( .A(n7241), .B(n7260), .Z(n7238) );
  NAND U7838 ( .A(A[0]), .B(B[726]), .Z(n7260) );
  NAND U7839 ( .A(B[725]), .B(A[1]), .Z(n7241) );
  NAND U7840 ( .A(n7261), .B(n7262), .Z(n641) );
  NANDN U7841 ( .A(n7263), .B(n7264), .Z(n7262) );
  OR U7842 ( .A(n7265), .B(n7266), .Z(n7264) );
  NAND U7843 ( .A(n7266), .B(n7265), .Z(n7261) );
  XOR U7844 ( .A(n643), .B(n642), .Z(\A1[723] ) );
  XOR U7845 ( .A(n7266), .B(n7267), .Z(n642) );
  XNOR U7846 ( .A(n7265), .B(n7263), .Z(n7267) );
  AND U7847 ( .A(n7268), .B(n7269), .Z(n7263) );
  NANDN U7848 ( .A(n7270), .B(n7271), .Z(n7269) );
  NANDN U7849 ( .A(n7272), .B(n7273), .Z(n7271) );
  AND U7850 ( .A(B[722]), .B(A[3]), .Z(n7265) );
  XNOR U7851 ( .A(n7255), .B(n7274), .Z(n7266) );
  XNOR U7852 ( .A(n7253), .B(n7256), .Z(n7274) );
  NAND U7853 ( .A(A[2]), .B(B[723]), .Z(n7256) );
  NANDN U7854 ( .A(n7275), .B(n7276), .Z(n7253) );
  AND U7855 ( .A(A[0]), .B(B[724]), .Z(n7276) );
  XOR U7856 ( .A(n7258), .B(n7277), .Z(n7255) );
  NAND U7857 ( .A(A[0]), .B(B[725]), .Z(n7277) );
  NAND U7858 ( .A(B[724]), .B(A[1]), .Z(n7258) );
  NAND U7859 ( .A(n7278), .B(n7279), .Z(n643) );
  NANDN U7860 ( .A(n7280), .B(n7281), .Z(n7279) );
  OR U7861 ( .A(n7282), .B(n7283), .Z(n7281) );
  NAND U7862 ( .A(n7283), .B(n7282), .Z(n7278) );
  XOR U7863 ( .A(n645), .B(n644), .Z(\A1[722] ) );
  XOR U7864 ( .A(n7283), .B(n7284), .Z(n644) );
  XNOR U7865 ( .A(n7282), .B(n7280), .Z(n7284) );
  AND U7866 ( .A(n7285), .B(n7286), .Z(n7280) );
  NANDN U7867 ( .A(n7287), .B(n7288), .Z(n7286) );
  NANDN U7868 ( .A(n7289), .B(n7290), .Z(n7288) );
  AND U7869 ( .A(B[721]), .B(A[3]), .Z(n7282) );
  XNOR U7870 ( .A(n7272), .B(n7291), .Z(n7283) );
  XNOR U7871 ( .A(n7270), .B(n7273), .Z(n7291) );
  NAND U7872 ( .A(A[2]), .B(B[722]), .Z(n7273) );
  NANDN U7873 ( .A(n7292), .B(n7293), .Z(n7270) );
  AND U7874 ( .A(A[0]), .B(B[723]), .Z(n7293) );
  XOR U7875 ( .A(n7275), .B(n7294), .Z(n7272) );
  NAND U7876 ( .A(A[0]), .B(B[724]), .Z(n7294) );
  NAND U7877 ( .A(B[723]), .B(A[1]), .Z(n7275) );
  NAND U7878 ( .A(n7295), .B(n7296), .Z(n645) );
  NANDN U7879 ( .A(n7297), .B(n7298), .Z(n7296) );
  OR U7880 ( .A(n7299), .B(n7300), .Z(n7298) );
  NAND U7881 ( .A(n7300), .B(n7299), .Z(n7295) );
  XOR U7882 ( .A(n647), .B(n646), .Z(\A1[721] ) );
  XOR U7883 ( .A(n7300), .B(n7301), .Z(n646) );
  XNOR U7884 ( .A(n7299), .B(n7297), .Z(n7301) );
  AND U7885 ( .A(n7302), .B(n7303), .Z(n7297) );
  NANDN U7886 ( .A(n7304), .B(n7305), .Z(n7303) );
  NANDN U7887 ( .A(n7306), .B(n7307), .Z(n7305) );
  AND U7888 ( .A(B[720]), .B(A[3]), .Z(n7299) );
  XNOR U7889 ( .A(n7289), .B(n7308), .Z(n7300) );
  XNOR U7890 ( .A(n7287), .B(n7290), .Z(n7308) );
  NAND U7891 ( .A(A[2]), .B(B[721]), .Z(n7290) );
  NANDN U7892 ( .A(n7309), .B(n7310), .Z(n7287) );
  AND U7893 ( .A(A[0]), .B(B[722]), .Z(n7310) );
  XOR U7894 ( .A(n7292), .B(n7311), .Z(n7289) );
  NAND U7895 ( .A(A[0]), .B(B[723]), .Z(n7311) );
  NAND U7896 ( .A(B[722]), .B(A[1]), .Z(n7292) );
  NAND U7897 ( .A(n7312), .B(n7313), .Z(n647) );
  NANDN U7898 ( .A(n7314), .B(n7315), .Z(n7313) );
  OR U7899 ( .A(n7316), .B(n7317), .Z(n7315) );
  NAND U7900 ( .A(n7317), .B(n7316), .Z(n7312) );
  XOR U7901 ( .A(n649), .B(n648), .Z(\A1[720] ) );
  XOR U7902 ( .A(n7317), .B(n7318), .Z(n648) );
  XNOR U7903 ( .A(n7316), .B(n7314), .Z(n7318) );
  AND U7904 ( .A(n7319), .B(n7320), .Z(n7314) );
  NANDN U7905 ( .A(n7321), .B(n7322), .Z(n7320) );
  NANDN U7906 ( .A(n7323), .B(n7324), .Z(n7322) );
  AND U7907 ( .A(B[719]), .B(A[3]), .Z(n7316) );
  XNOR U7908 ( .A(n7306), .B(n7325), .Z(n7317) );
  XNOR U7909 ( .A(n7304), .B(n7307), .Z(n7325) );
  NAND U7910 ( .A(A[2]), .B(B[720]), .Z(n7307) );
  NANDN U7911 ( .A(n7326), .B(n7327), .Z(n7304) );
  AND U7912 ( .A(A[0]), .B(B[721]), .Z(n7327) );
  XOR U7913 ( .A(n7309), .B(n7328), .Z(n7306) );
  NAND U7914 ( .A(A[0]), .B(B[722]), .Z(n7328) );
  NAND U7915 ( .A(B[721]), .B(A[1]), .Z(n7309) );
  NAND U7916 ( .A(n7329), .B(n7330), .Z(n649) );
  NANDN U7917 ( .A(n7331), .B(n7332), .Z(n7330) );
  OR U7918 ( .A(n7333), .B(n7334), .Z(n7332) );
  NAND U7919 ( .A(n7334), .B(n7333), .Z(n7329) );
  XOR U7920 ( .A(n631), .B(n630), .Z(\A1[71] ) );
  XOR U7921 ( .A(n7164), .B(n7335), .Z(n630) );
  XNOR U7922 ( .A(n7163), .B(n7161), .Z(n7335) );
  AND U7923 ( .A(n7336), .B(n7337), .Z(n7161) );
  NANDN U7924 ( .A(n7338), .B(n7339), .Z(n7337) );
  NANDN U7925 ( .A(n7340), .B(n7341), .Z(n7339) );
  AND U7926 ( .A(B[70]), .B(A[3]), .Z(n7163) );
  XNOR U7927 ( .A(n7153), .B(n7342), .Z(n7164) );
  XNOR U7928 ( .A(n7151), .B(n7154), .Z(n7342) );
  NAND U7929 ( .A(A[2]), .B(B[71]), .Z(n7154) );
  NANDN U7930 ( .A(n7343), .B(n7344), .Z(n7151) );
  AND U7931 ( .A(A[0]), .B(B[72]), .Z(n7344) );
  XOR U7932 ( .A(n7156), .B(n7345), .Z(n7153) );
  NAND U7933 ( .A(A[0]), .B(B[73]), .Z(n7345) );
  NAND U7934 ( .A(B[72]), .B(A[1]), .Z(n7156) );
  NAND U7935 ( .A(n7346), .B(n7347), .Z(n631) );
  NANDN U7936 ( .A(n7348), .B(n7349), .Z(n7347) );
  OR U7937 ( .A(n7350), .B(n7351), .Z(n7349) );
  NAND U7938 ( .A(n7351), .B(n7350), .Z(n7346) );
  XOR U7939 ( .A(n651), .B(n650), .Z(\A1[719] ) );
  XOR U7940 ( .A(n7334), .B(n7352), .Z(n650) );
  XNOR U7941 ( .A(n7333), .B(n7331), .Z(n7352) );
  AND U7942 ( .A(n7353), .B(n7354), .Z(n7331) );
  NANDN U7943 ( .A(n7355), .B(n7356), .Z(n7354) );
  NANDN U7944 ( .A(n7357), .B(n7358), .Z(n7356) );
  AND U7945 ( .A(B[718]), .B(A[3]), .Z(n7333) );
  XNOR U7946 ( .A(n7323), .B(n7359), .Z(n7334) );
  XNOR U7947 ( .A(n7321), .B(n7324), .Z(n7359) );
  NAND U7948 ( .A(A[2]), .B(B[719]), .Z(n7324) );
  NANDN U7949 ( .A(n7360), .B(n7361), .Z(n7321) );
  AND U7950 ( .A(A[0]), .B(B[720]), .Z(n7361) );
  XOR U7951 ( .A(n7326), .B(n7362), .Z(n7323) );
  NAND U7952 ( .A(A[0]), .B(B[721]), .Z(n7362) );
  NAND U7953 ( .A(B[720]), .B(A[1]), .Z(n7326) );
  NAND U7954 ( .A(n7363), .B(n7364), .Z(n651) );
  NANDN U7955 ( .A(n7365), .B(n7366), .Z(n7364) );
  OR U7956 ( .A(n7367), .B(n7368), .Z(n7366) );
  NAND U7957 ( .A(n7368), .B(n7367), .Z(n7363) );
  XOR U7958 ( .A(n655), .B(n654), .Z(\A1[718] ) );
  XOR U7959 ( .A(n7368), .B(n7369), .Z(n654) );
  XNOR U7960 ( .A(n7367), .B(n7365), .Z(n7369) );
  AND U7961 ( .A(n7370), .B(n7371), .Z(n7365) );
  NANDN U7962 ( .A(n7372), .B(n7373), .Z(n7371) );
  NANDN U7963 ( .A(n7374), .B(n7375), .Z(n7373) );
  AND U7964 ( .A(B[717]), .B(A[3]), .Z(n7367) );
  XNOR U7965 ( .A(n7357), .B(n7376), .Z(n7368) );
  XNOR U7966 ( .A(n7355), .B(n7358), .Z(n7376) );
  NAND U7967 ( .A(A[2]), .B(B[718]), .Z(n7358) );
  NANDN U7968 ( .A(n7377), .B(n7378), .Z(n7355) );
  AND U7969 ( .A(A[0]), .B(B[719]), .Z(n7378) );
  XOR U7970 ( .A(n7360), .B(n7379), .Z(n7357) );
  NAND U7971 ( .A(A[0]), .B(B[720]), .Z(n7379) );
  NAND U7972 ( .A(B[719]), .B(A[1]), .Z(n7360) );
  NAND U7973 ( .A(n7380), .B(n7381), .Z(n655) );
  NANDN U7974 ( .A(n7382), .B(n7383), .Z(n7381) );
  OR U7975 ( .A(n7384), .B(n7385), .Z(n7383) );
  NAND U7976 ( .A(n7385), .B(n7384), .Z(n7380) );
  XOR U7977 ( .A(n657), .B(n656), .Z(\A1[717] ) );
  XOR U7978 ( .A(n7385), .B(n7386), .Z(n656) );
  XNOR U7979 ( .A(n7384), .B(n7382), .Z(n7386) );
  AND U7980 ( .A(n7387), .B(n7388), .Z(n7382) );
  NANDN U7981 ( .A(n7389), .B(n7390), .Z(n7388) );
  NANDN U7982 ( .A(n7391), .B(n7392), .Z(n7390) );
  AND U7983 ( .A(B[716]), .B(A[3]), .Z(n7384) );
  XNOR U7984 ( .A(n7374), .B(n7393), .Z(n7385) );
  XNOR U7985 ( .A(n7372), .B(n7375), .Z(n7393) );
  NAND U7986 ( .A(A[2]), .B(B[717]), .Z(n7375) );
  NANDN U7987 ( .A(n7394), .B(n7395), .Z(n7372) );
  AND U7988 ( .A(A[0]), .B(B[718]), .Z(n7395) );
  XOR U7989 ( .A(n7377), .B(n7396), .Z(n7374) );
  NAND U7990 ( .A(A[0]), .B(B[719]), .Z(n7396) );
  NAND U7991 ( .A(B[718]), .B(A[1]), .Z(n7377) );
  NAND U7992 ( .A(n7397), .B(n7398), .Z(n657) );
  NANDN U7993 ( .A(n7399), .B(n7400), .Z(n7398) );
  OR U7994 ( .A(n7401), .B(n7402), .Z(n7400) );
  NAND U7995 ( .A(n7402), .B(n7401), .Z(n7397) );
  XOR U7996 ( .A(n659), .B(n658), .Z(\A1[716] ) );
  XOR U7997 ( .A(n7402), .B(n7403), .Z(n658) );
  XNOR U7998 ( .A(n7401), .B(n7399), .Z(n7403) );
  AND U7999 ( .A(n7404), .B(n7405), .Z(n7399) );
  NANDN U8000 ( .A(n7406), .B(n7407), .Z(n7405) );
  NANDN U8001 ( .A(n7408), .B(n7409), .Z(n7407) );
  AND U8002 ( .A(B[715]), .B(A[3]), .Z(n7401) );
  XNOR U8003 ( .A(n7391), .B(n7410), .Z(n7402) );
  XNOR U8004 ( .A(n7389), .B(n7392), .Z(n7410) );
  NAND U8005 ( .A(A[2]), .B(B[716]), .Z(n7392) );
  NANDN U8006 ( .A(n7411), .B(n7412), .Z(n7389) );
  AND U8007 ( .A(A[0]), .B(B[717]), .Z(n7412) );
  XOR U8008 ( .A(n7394), .B(n7413), .Z(n7391) );
  NAND U8009 ( .A(A[0]), .B(B[718]), .Z(n7413) );
  NAND U8010 ( .A(B[717]), .B(A[1]), .Z(n7394) );
  NAND U8011 ( .A(n7414), .B(n7415), .Z(n659) );
  NANDN U8012 ( .A(n7416), .B(n7417), .Z(n7415) );
  OR U8013 ( .A(n7418), .B(n7419), .Z(n7417) );
  NAND U8014 ( .A(n7419), .B(n7418), .Z(n7414) );
  XOR U8015 ( .A(n661), .B(n660), .Z(\A1[715] ) );
  XOR U8016 ( .A(n7419), .B(n7420), .Z(n660) );
  XNOR U8017 ( .A(n7418), .B(n7416), .Z(n7420) );
  AND U8018 ( .A(n7421), .B(n7422), .Z(n7416) );
  NANDN U8019 ( .A(n7423), .B(n7424), .Z(n7422) );
  NANDN U8020 ( .A(n7425), .B(n7426), .Z(n7424) );
  AND U8021 ( .A(B[714]), .B(A[3]), .Z(n7418) );
  XNOR U8022 ( .A(n7408), .B(n7427), .Z(n7419) );
  XNOR U8023 ( .A(n7406), .B(n7409), .Z(n7427) );
  NAND U8024 ( .A(A[2]), .B(B[715]), .Z(n7409) );
  NANDN U8025 ( .A(n7428), .B(n7429), .Z(n7406) );
  AND U8026 ( .A(A[0]), .B(B[716]), .Z(n7429) );
  XOR U8027 ( .A(n7411), .B(n7430), .Z(n7408) );
  NAND U8028 ( .A(A[0]), .B(B[717]), .Z(n7430) );
  NAND U8029 ( .A(B[716]), .B(A[1]), .Z(n7411) );
  NAND U8030 ( .A(n7431), .B(n7432), .Z(n661) );
  NANDN U8031 ( .A(n7433), .B(n7434), .Z(n7432) );
  OR U8032 ( .A(n7435), .B(n7436), .Z(n7434) );
  NAND U8033 ( .A(n7436), .B(n7435), .Z(n7431) );
  XOR U8034 ( .A(n663), .B(n662), .Z(\A1[714] ) );
  XOR U8035 ( .A(n7436), .B(n7437), .Z(n662) );
  XNOR U8036 ( .A(n7435), .B(n7433), .Z(n7437) );
  AND U8037 ( .A(n7438), .B(n7439), .Z(n7433) );
  NANDN U8038 ( .A(n7440), .B(n7441), .Z(n7439) );
  NANDN U8039 ( .A(n7442), .B(n7443), .Z(n7441) );
  AND U8040 ( .A(B[713]), .B(A[3]), .Z(n7435) );
  XNOR U8041 ( .A(n7425), .B(n7444), .Z(n7436) );
  XNOR U8042 ( .A(n7423), .B(n7426), .Z(n7444) );
  NAND U8043 ( .A(A[2]), .B(B[714]), .Z(n7426) );
  NANDN U8044 ( .A(n7445), .B(n7446), .Z(n7423) );
  AND U8045 ( .A(A[0]), .B(B[715]), .Z(n7446) );
  XOR U8046 ( .A(n7428), .B(n7447), .Z(n7425) );
  NAND U8047 ( .A(A[0]), .B(B[716]), .Z(n7447) );
  NAND U8048 ( .A(B[715]), .B(A[1]), .Z(n7428) );
  NAND U8049 ( .A(n7448), .B(n7449), .Z(n663) );
  NANDN U8050 ( .A(n7450), .B(n7451), .Z(n7449) );
  OR U8051 ( .A(n7452), .B(n7453), .Z(n7451) );
  NAND U8052 ( .A(n7453), .B(n7452), .Z(n7448) );
  XOR U8053 ( .A(n665), .B(n664), .Z(\A1[713] ) );
  XOR U8054 ( .A(n7453), .B(n7454), .Z(n664) );
  XNOR U8055 ( .A(n7452), .B(n7450), .Z(n7454) );
  AND U8056 ( .A(n7455), .B(n7456), .Z(n7450) );
  NANDN U8057 ( .A(n7457), .B(n7458), .Z(n7456) );
  NANDN U8058 ( .A(n7459), .B(n7460), .Z(n7458) );
  AND U8059 ( .A(B[712]), .B(A[3]), .Z(n7452) );
  XNOR U8060 ( .A(n7442), .B(n7461), .Z(n7453) );
  XNOR U8061 ( .A(n7440), .B(n7443), .Z(n7461) );
  NAND U8062 ( .A(A[2]), .B(B[713]), .Z(n7443) );
  NANDN U8063 ( .A(n7462), .B(n7463), .Z(n7440) );
  AND U8064 ( .A(A[0]), .B(B[714]), .Z(n7463) );
  XOR U8065 ( .A(n7445), .B(n7464), .Z(n7442) );
  NAND U8066 ( .A(A[0]), .B(B[715]), .Z(n7464) );
  NAND U8067 ( .A(B[714]), .B(A[1]), .Z(n7445) );
  NAND U8068 ( .A(n7465), .B(n7466), .Z(n665) );
  NANDN U8069 ( .A(n7467), .B(n7468), .Z(n7466) );
  OR U8070 ( .A(n7469), .B(n7470), .Z(n7468) );
  NAND U8071 ( .A(n7470), .B(n7469), .Z(n7465) );
  XOR U8072 ( .A(n667), .B(n666), .Z(\A1[712] ) );
  XOR U8073 ( .A(n7470), .B(n7471), .Z(n666) );
  XNOR U8074 ( .A(n7469), .B(n7467), .Z(n7471) );
  AND U8075 ( .A(n7472), .B(n7473), .Z(n7467) );
  NANDN U8076 ( .A(n7474), .B(n7475), .Z(n7473) );
  NANDN U8077 ( .A(n7476), .B(n7477), .Z(n7475) );
  AND U8078 ( .A(B[711]), .B(A[3]), .Z(n7469) );
  XNOR U8079 ( .A(n7459), .B(n7478), .Z(n7470) );
  XNOR U8080 ( .A(n7457), .B(n7460), .Z(n7478) );
  NAND U8081 ( .A(A[2]), .B(B[712]), .Z(n7460) );
  NANDN U8082 ( .A(n7479), .B(n7480), .Z(n7457) );
  AND U8083 ( .A(A[0]), .B(B[713]), .Z(n7480) );
  XOR U8084 ( .A(n7462), .B(n7481), .Z(n7459) );
  NAND U8085 ( .A(A[0]), .B(B[714]), .Z(n7481) );
  NAND U8086 ( .A(B[713]), .B(A[1]), .Z(n7462) );
  NAND U8087 ( .A(n7482), .B(n7483), .Z(n667) );
  NANDN U8088 ( .A(n7484), .B(n7485), .Z(n7483) );
  OR U8089 ( .A(n7486), .B(n7487), .Z(n7485) );
  NAND U8090 ( .A(n7487), .B(n7486), .Z(n7482) );
  XOR U8091 ( .A(n669), .B(n668), .Z(\A1[711] ) );
  XOR U8092 ( .A(n7487), .B(n7488), .Z(n668) );
  XNOR U8093 ( .A(n7486), .B(n7484), .Z(n7488) );
  AND U8094 ( .A(n7489), .B(n7490), .Z(n7484) );
  NANDN U8095 ( .A(n7491), .B(n7492), .Z(n7490) );
  NANDN U8096 ( .A(n7493), .B(n7494), .Z(n7492) );
  AND U8097 ( .A(B[710]), .B(A[3]), .Z(n7486) );
  XNOR U8098 ( .A(n7476), .B(n7495), .Z(n7487) );
  XNOR U8099 ( .A(n7474), .B(n7477), .Z(n7495) );
  NAND U8100 ( .A(A[2]), .B(B[711]), .Z(n7477) );
  NANDN U8101 ( .A(n7496), .B(n7497), .Z(n7474) );
  AND U8102 ( .A(A[0]), .B(B[712]), .Z(n7497) );
  XOR U8103 ( .A(n7479), .B(n7498), .Z(n7476) );
  NAND U8104 ( .A(A[0]), .B(B[713]), .Z(n7498) );
  NAND U8105 ( .A(B[712]), .B(A[1]), .Z(n7479) );
  NAND U8106 ( .A(n7499), .B(n7500), .Z(n669) );
  NANDN U8107 ( .A(n7501), .B(n7502), .Z(n7500) );
  OR U8108 ( .A(n7503), .B(n7504), .Z(n7502) );
  NAND U8109 ( .A(n7504), .B(n7503), .Z(n7499) );
  XOR U8110 ( .A(n671), .B(n670), .Z(\A1[710] ) );
  XOR U8111 ( .A(n7504), .B(n7505), .Z(n670) );
  XNOR U8112 ( .A(n7503), .B(n7501), .Z(n7505) );
  AND U8113 ( .A(n7506), .B(n7507), .Z(n7501) );
  NANDN U8114 ( .A(n7508), .B(n7509), .Z(n7507) );
  NANDN U8115 ( .A(n7510), .B(n7511), .Z(n7509) );
  AND U8116 ( .A(B[709]), .B(A[3]), .Z(n7503) );
  XNOR U8117 ( .A(n7493), .B(n7512), .Z(n7504) );
  XNOR U8118 ( .A(n7491), .B(n7494), .Z(n7512) );
  NAND U8119 ( .A(A[2]), .B(B[710]), .Z(n7494) );
  NANDN U8120 ( .A(n7513), .B(n7514), .Z(n7491) );
  AND U8121 ( .A(A[0]), .B(B[711]), .Z(n7514) );
  XOR U8122 ( .A(n7496), .B(n7515), .Z(n7493) );
  NAND U8123 ( .A(A[0]), .B(B[712]), .Z(n7515) );
  NAND U8124 ( .A(B[711]), .B(A[1]), .Z(n7496) );
  NAND U8125 ( .A(n7516), .B(n7517), .Z(n671) );
  NANDN U8126 ( .A(n7518), .B(n7519), .Z(n7517) );
  OR U8127 ( .A(n7520), .B(n7521), .Z(n7519) );
  NAND U8128 ( .A(n7521), .B(n7520), .Z(n7516) );
  XOR U8129 ( .A(n653), .B(n652), .Z(\A1[70] ) );
  XOR U8130 ( .A(n7351), .B(n7522), .Z(n652) );
  XNOR U8131 ( .A(n7350), .B(n7348), .Z(n7522) );
  AND U8132 ( .A(n7523), .B(n7524), .Z(n7348) );
  NANDN U8133 ( .A(n7525), .B(n7526), .Z(n7524) );
  NANDN U8134 ( .A(n7527), .B(n7528), .Z(n7526) );
  AND U8135 ( .A(B[69]), .B(A[3]), .Z(n7350) );
  XNOR U8136 ( .A(n7340), .B(n7529), .Z(n7351) );
  XNOR U8137 ( .A(n7338), .B(n7341), .Z(n7529) );
  NAND U8138 ( .A(A[2]), .B(B[70]), .Z(n7341) );
  NANDN U8139 ( .A(n7530), .B(n7531), .Z(n7338) );
  AND U8140 ( .A(A[0]), .B(B[71]), .Z(n7531) );
  XOR U8141 ( .A(n7343), .B(n7532), .Z(n7340) );
  NAND U8142 ( .A(A[0]), .B(B[72]), .Z(n7532) );
  NAND U8143 ( .A(B[71]), .B(A[1]), .Z(n7343) );
  NAND U8144 ( .A(n7533), .B(n7534), .Z(n653) );
  NANDN U8145 ( .A(n7535), .B(n7536), .Z(n7534) );
  OR U8146 ( .A(n7537), .B(n7538), .Z(n7536) );
  NAND U8147 ( .A(n7538), .B(n7537), .Z(n7533) );
  XOR U8148 ( .A(n673), .B(n672), .Z(\A1[709] ) );
  XOR U8149 ( .A(n7521), .B(n7539), .Z(n672) );
  XNOR U8150 ( .A(n7520), .B(n7518), .Z(n7539) );
  AND U8151 ( .A(n7540), .B(n7541), .Z(n7518) );
  NANDN U8152 ( .A(n7542), .B(n7543), .Z(n7541) );
  NANDN U8153 ( .A(n7544), .B(n7545), .Z(n7543) );
  AND U8154 ( .A(B[708]), .B(A[3]), .Z(n7520) );
  XNOR U8155 ( .A(n7510), .B(n7546), .Z(n7521) );
  XNOR U8156 ( .A(n7508), .B(n7511), .Z(n7546) );
  NAND U8157 ( .A(A[2]), .B(B[709]), .Z(n7511) );
  NANDN U8158 ( .A(n7547), .B(n7548), .Z(n7508) );
  AND U8159 ( .A(A[0]), .B(B[710]), .Z(n7548) );
  XOR U8160 ( .A(n7513), .B(n7549), .Z(n7510) );
  NAND U8161 ( .A(A[0]), .B(B[711]), .Z(n7549) );
  NAND U8162 ( .A(B[710]), .B(A[1]), .Z(n7513) );
  NAND U8163 ( .A(n7550), .B(n7551), .Z(n673) );
  NANDN U8164 ( .A(n7552), .B(n7553), .Z(n7551) );
  OR U8165 ( .A(n7554), .B(n7555), .Z(n7553) );
  NAND U8166 ( .A(n7555), .B(n7554), .Z(n7550) );
  XOR U8167 ( .A(n677), .B(n676), .Z(\A1[708] ) );
  XOR U8168 ( .A(n7555), .B(n7556), .Z(n676) );
  XNOR U8169 ( .A(n7554), .B(n7552), .Z(n7556) );
  AND U8170 ( .A(n7557), .B(n7558), .Z(n7552) );
  NANDN U8171 ( .A(n7559), .B(n7560), .Z(n7558) );
  NANDN U8172 ( .A(n7561), .B(n7562), .Z(n7560) );
  AND U8173 ( .A(B[707]), .B(A[3]), .Z(n7554) );
  XNOR U8174 ( .A(n7544), .B(n7563), .Z(n7555) );
  XNOR U8175 ( .A(n7542), .B(n7545), .Z(n7563) );
  NAND U8176 ( .A(A[2]), .B(B[708]), .Z(n7545) );
  NANDN U8177 ( .A(n7564), .B(n7565), .Z(n7542) );
  AND U8178 ( .A(A[0]), .B(B[709]), .Z(n7565) );
  XOR U8179 ( .A(n7547), .B(n7566), .Z(n7544) );
  NAND U8180 ( .A(A[0]), .B(B[710]), .Z(n7566) );
  NAND U8181 ( .A(B[709]), .B(A[1]), .Z(n7547) );
  NAND U8182 ( .A(n7567), .B(n7568), .Z(n677) );
  NANDN U8183 ( .A(n7569), .B(n7570), .Z(n7568) );
  OR U8184 ( .A(n7571), .B(n7572), .Z(n7570) );
  NAND U8185 ( .A(n7572), .B(n7571), .Z(n7567) );
  XOR U8186 ( .A(n679), .B(n678), .Z(\A1[707] ) );
  XOR U8187 ( .A(n7572), .B(n7573), .Z(n678) );
  XNOR U8188 ( .A(n7571), .B(n7569), .Z(n7573) );
  AND U8189 ( .A(n7574), .B(n7575), .Z(n7569) );
  NANDN U8190 ( .A(n7576), .B(n7577), .Z(n7575) );
  NANDN U8191 ( .A(n7578), .B(n7579), .Z(n7577) );
  AND U8192 ( .A(B[706]), .B(A[3]), .Z(n7571) );
  XNOR U8193 ( .A(n7561), .B(n7580), .Z(n7572) );
  XNOR U8194 ( .A(n7559), .B(n7562), .Z(n7580) );
  NAND U8195 ( .A(A[2]), .B(B[707]), .Z(n7562) );
  NANDN U8196 ( .A(n7581), .B(n7582), .Z(n7559) );
  AND U8197 ( .A(A[0]), .B(B[708]), .Z(n7582) );
  XOR U8198 ( .A(n7564), .B(n7583), .Z(n7561) );
  NAND U8199 ( .A(A[0]), .B(B[709]), .Z(n7583) );
  NAND U8200 ( .A(B[708]), .B(A[1]), .Z(n7564) );
  NAND U8201 ( .A(n7584), .B(n7585), .Z(n679) );
  NANDN U8202 ( .A(n7586), .B(n7587), .Z(n7585) );
  OR U8203 ( .A(n7588), .B(n7589), .Z(n7587) );
  NAND U8204 ( .A(n7589), .B(n7588), .Z(n7584) );
  XOR U8205 ( .A(n681), .B(n680), .Z(\A1[706] ) );
  XOR U8206 ( .A(n7589), .B(n7590), .Z(n680) );
  XNOR U8207 ( .A(n7588), .B(n7586), .Z(n7590) );
  AND U8208 ( .A(n7591), .B(n7592), .Z(n7586) );
  NANDN U8209 ( .A(n7593), .B(n7594), .Z(n7592) );
  NANDN U8210 ( .A(n7595), .B(n7596), .Z(n7594) );
  AND U8211 ( .A(B[705]), .B(A[3]), .Z(n7588) );
  XNOR U8212 ( .A(n7578), .B(n7597), .Z(n7589) );
  XNOR U8213 ( .A(n7576), .B(n7579), .Z(n7597) );
  NAND U8214 ( .A(A[2]), .B(B[706]), .Z(n7579) );
  NANDN U8215 ( .A(n7598), .B(n7599), .Z(n7576) );
  AND U8216 ( .A(A[0]), .B(B[707]), .Z(n7599) );
  XOR U8217 ( .A(n7581), .B(n7600), .Z(n7578) );
  NAND U8218 ( .A(A[0]), .B(B[708]), .Z(n7600) );
  NAND U8219 ( .A(B[707]), .B(A[1]), .Z(n7581) );
  NAND U8220 ( .A(n7601), .B(n7602), .Z(n681) );
  NANDN U8221 ( .A(n7603), .B(n7604), .Z(n7602) );
  OR U8222 ( .A(n7605), .B(n7606), .Z(n7604) );
  NAND U8223 ( .A(n7606), .B(n7605), .Z(n7601) );
  XOR U8224 ( .A(n683), .B(n682), .Z(\A1[705] ) );
  XOR U8225 ( .A(n7606), .B(n7607), .Z(n682) );
  XNOR U8226 ( .A(n7605), .B(n7603), .Z(n7607) );
  AND U8227 ( .A(n7608), .B(n7609), .Z(n7603) );
  NANDN U8228 ( .A(n7610), .B(n7611), .Z(n7609) );
  NANDN U8229 ( .A(n7612), .B(n7613), .Z(n7611) );
  AND U8230 ( .A(B[704]), .B(A[3]), .Z(n7605) );
  XNOR U8231 ( .A(n7595), .B(n7614), .Z(n7606) );
  XNOR U8232 ( .A(n7593), .B(n7596), .Z(n7614) );
  NAND U8233 ( .A(A[2]), .B(B[705]), .Z(n7596) );
  NANDN U8234 ( .A(n7615), .B(n7616), .Z(n7593) );
  AND U8235 ( .A(A[0]), .B(B[706]), .Z(n7616) );
  XOR U8236 ( .A(n7598), .B(n7617), .Z(n7595) );
  NAND U8237 ( .A(A[0]), .B(B[707]), .Z(n7617) );
  NAND U8238 ( .A(B[706]), .B(A[1]), .Z(n7598) );
  NAND U8239 ( .A(n7618), .B(n7619), .Z(n683) );
  NANDN U8240 ( .A(n7620), .B(n7621), .Z(n7619) );
  OR U8241 ( .A(n7622), .B(n7623), .Z(n7621) );
  NAND U8242 ( .A(n7623), .B(n7622), .Z(n7618) );
  XOR U8243 ( .A(n685), .B(n684), .Z(\A1[704] ) );
  XOR U8244 ( .A(n7623), .B(n7624), .Z(n684) );
  XNOR U8245 ( .A(n7622), .B(n7620), .Z(n7624) );
  AND U8246 ( .A(n7625), .B(n7626), .Z(n7620) );
  NANDN U8247 ( .A(n7627), .B(n7628), .Z(n7626) );
  NANDN U8248 ( .A(n7629), .B(n7630), .Z(n7628) );
  AND U8249 ( .A(B[703]), .B(A[3]), .Z(n7622) );
  XNOR U8250 ( .A(n7612), .B(n7631), .Z(n7623) );
  XNOR U8251 ( .A(n7610), .B(n7613), .Z(n7631) );
  NAND U8252 ( .A(A[2]), .B(B[704]), .Z(n7613) );
  NANDN U8253 ( .A(n7632), .B(n7633), .Z(n7610) );
  AND U8254 ( .A(A[0]), .B(B[705]), .Z(n7633) );
  XOR U8255 ( .A(n7615), .B(n7634), .Z(n7612) );
  NAND U8256 ( .A(A[0]), .B(B[706]), .Z(n7634) );
  NAND U8257 ( .A(B[705]), .B(A[1]), .Z(n7615) );
  NAND U8258 ( .A(n7635), .B(n7636), .Z(n685) );
  NANDN U8259 ( .A(n7637), .B(n7638), .Z(n7636) );
  OR U8260 ( .A(n7639), .B(n7640), .Z(n7638) );
  NAND U8261 ( .A(n7640), .B(n7639), .Z(n7635) );
  XOR U8262 ( .A(n687), .B(n686), .Z(\A1[703] ) );
  XOR U8263 ( .A(n7640), .B(n7641), .Z(n686) );
  XNOR U8264 ( .A(n7639), .B(n7637), .Z(n7641) );
  AND U8265 ( .A(n7642), .B(n7643), .Z(n7637) );
  NANDN U8266 ( .A(n7644), .B(n7645), .Z(n7643) );
  NANDN U8267 ( .A(n7646), .B(n7647), .Z(n7645) );
  AND U8268 ( .A(B[702]), .B(A[3]), .Z(n7639) );
  XNOR U8269 ( .A(n7629), .B(n7648), .Z(n7640) );
  XNOR U8270 ( .A(n7627), .B(n7630), .Z(n7648) );
  NAND U8271 ( .A(A[2]), .B(B[703]), .Z(n7630) );
  NANDN U8272 ( .A(n7649), .B(n7650), .Z(n7627) );
  AND U8273 ( .A(A[0]), .B(B[704]), .Z(n7650) );
  XOR U8274 ( .A(n7632), .B(n7651), .Z(n7629) );
  NAND U8275 ( .A(A[0]), .B(B[705]), .Z(n7651) );
  NAND U8276 ( .A(B[704]), .B(A[1]), .Z(n7632) );
  NAND U8277 ( .A(n7652), .B(n7653), .Z(n687) );
  NANDN U8278 ( .A(n7654), .B(n7655), .Z(n7653) );
  OR U8279 ( .A(n7656), .B(n7657), .Z(n7655) );
  NAND U8280 ( .A(n7657), .B(n7656), .Z(n7652) );
  XOR U8281 ( .A(n689), .B(n688), .Z(\A1[702] ) );
  XOR U8282 ( .A(n7657), .B(n7658), .Z(n688) );
  XNOR U8283 ( .A(n7656), .B(n7654), .Z(n7658) );
  AND U8284 ( .A(n7659), .B(n7660), .Z(n7654) );
  NANDN U8285 ( .A(n7661), .B(n7662), .Z(n7660) );
  NANDN U8286 ( .A(n7663), .B(n7664), .Z(n7662) );
  AND U8287 ( .A(B[701]), .B(A[3]), .Z(n7656) );
  XNOR U8288 ( .A(n7646), .B(n7665), .Z(n7657) );
  XNOR U8289 ( .A(n7644), .B(n7647), .Z(n7665) );
  NAND U8290 ( .A(A[2]), .B(B[702]), .Z(n7647) );
  NANDN U8291 ( .A(n7666), .B(n7667), .Z(n7644) );
  AND U8292 ( .A(A[0]), .B(B[703]), .Z(n7667) );
  XOR U8293 ( .A(n7649), .B(n7668), .Z(n7646) );
  NAND U8294 ( .A(A[0]), .B(B[704]), .Z(n7668) );
  NAND U8295 ( .A(B[703]), .B(A[1]), .Z(n7649) );
  NAND U8296 ( .A(n7669), .B(n7670), .Z(n689) );
  NANDN U8297 ( .A(n7671), .B(n7672), .Z(n7670) );
  OR U8298 ( .A(n7673), .B(n7674), .Z(n7672) );
  NAND U8299 ( .A(n7674), .B(n7673), .Z(n7669) );
  XOR U8300 ( .A(n691), .B(n690), .Z(\A1[701] ) );
  XOR U8301 ( .A(n7674), .B(n7675), .Z(n690) );
  XNOR U8302 ( .A(n7673), .B(n7671), .Z(n7675) );
  AND U8303 ( .A(n7676), .B(n7677), .Z(n7671) );
  NANDN U8304 ( .A(n7678), .B(n7679), .Z(n7677) );
  NANDN U8305 ( .A(n7680), .B(n7681), .Z(n7679) );
  AND U8306 ( .A(B[700]), .B(A[3]), .Z(n7673) );
  XNOR U8307 ( .A(n7663), .B(n7682), .Z(n7674) );
  XNOR U8308 ( .A(n7661), .B(n7664), .Z(n7682) );
  NAND U8309 ( .A(A[2]), .B(B[701]), .Z(n7664) );
  NANDN U8310 ( .A(n7683), .B(n7684), .Z(n7661) );
  AND U8311 ( .A(A[0]), .B(B[702]), .Z(n7684) );
  XOR U8312 ( .A(n7666), .B(n7685), .Z(n7663) );
  NAND U8313 ( .A(A[0]), .B(B[703]), .Z(n7685) );
  NAND U8314 ( .A(B[702]), .B(A[1]), .Z(n7666) );
  NAND U8315 ( .A(n7686), .B(n7687), .Z(n691) );
  NANDN U8316 ( .A(n7688), .B(n7689), .Z(n7687) );
  OR U8317 ( .A(n7690), .B(n7691), .Z(n7689) );
  NAND U8318 ( .A(n7691), .B(n7690), .Z(n7686) );
  XOR U8319 ( .A(n693), .B(n692), .Z(\A1[700] ) );
  XOR U8320 ( .A(n7691), .B(n7692), .Z(n692) );
  XNOR U8321 ( .A(n7690), .B(n7688), .Z(n7692) );
  AND U8322 ( .A(n7693), .B(n7694), .Z(n7688) );
  NANDN U8323 ( .A(n7695), .B(n7696), .Z(n7694) );
  NANDN U8324 ( .A(n7697), .B(n7698), .Z(n7696) );
  AND U8325 ( .A(B[699]), .B(A[3]), .Z(n7690) );
  XNOR U8326 ( .A(n7680), .B(n7699), .Z(n7691) );
  XNOR U8327 ( .A(n7678), .B(n7681), .Z(n7699) );
  NAND U8328 ( .A(A[2]), .B(B[700]), .Z(n7681) );
  NANDN U8329 ( .A(n7700), .B(n7701), .Z(n7678) );
  AND U8330 ( .A(A[0]), .B(B[701]), .Z(n7701) );
  XOR U8331 ( .A(n7683), .B(n7702), .Z(n7680) );
  NAND U8332 ( .A(A[0]), .B(B[702]), .Z(n7702) );
  NAND U8333 ( .A(B[701]), .B(A[1]), .Z(n7683) );
  NAND U8334 ( .A(n7703), .B(n7704), .Z(n693) );
  NANDN U8335 ( .A(n7705), .B(n7706), .Z(n7704) );
  OR U8336 ( .A(n7707), .B(n7708), .Z(n7706) );
  NAND U8337 ( .A(n7708), .B(n7707), .Z(n7703) );
  XOR U8338 ( .A(n475), .B(n474), .Z(\A1[6] ) );
  XOR U8339 ( .A(n5838), .B(n7709), .Z(n474) );
  XNOR U8340 ( .A(n5837), .B(n5835), .Z(n7709) );
  AND U8341 ( .A(n7710), .B(n7711), .Z(n5835) );
  NANDN U8342 ( .A(n7712), .B(n7713), .Z(n7711) );
  NANDN U8343 ( .A(n7714), .B(n7715), .Z(n7713) );
  AND U8344 ( .A(B[5]), .B(A[3]), .Z(n5837) );
  XNOR U8345 ( .A(n5826), .B(n7716), .Z(n5838) );
  XNOR U8346 ( .A(n5824), .B(n5827), .Z(n7716) );
  NAND U8347 ( .A(B[6]), .B(A[2]), .Z(n5827) );
  NAND U8348 ( .A(n7717), .B(B[7]), .Z(n5824) );
  ANDN U8349 ( .B(A[0]), .A(n7718), .Z(n7717) );
  XOR U8350 ( .A(n5830), .B(n7719), .Z(n5826) );
  NAND U8351 ( .A(A[0]), .B(B[8]), .Z(n7719) );
  NAND U8352 ( .A(B[7]), .B(A[1]), .Z(n5830) );
  NAND U8353 ( .A(n7720), .B(n7721), .Z(n475) );
  NANDN U8354 ( .A(n7722), .B(n7723), .Z(n7721) );
  OR U8355 ( .A(n7724), .B(n7725), .Z(n7723) );
  NAND U8356 ( .A(n7725), .B(n7724), .Z(n7720) );
  XOR U8357 ( .A(n675), .B(n674), .Z(\A1[69] ) );
  XOR U8358 ( .A(n7538), .B(n7726), .Z(n674) );
  XNOR U8359 ( .A(n7537), .B(n7535), .Z(n7726) );
  AND U8360 ( .A(n7727), .B(n7728), .Z(n7535) );
  NANDN U8361 ( .A(n7729), .B(n7730), .Z(n7728) );
  NANDN U8362 ( .A(n7731), .B(n7732), .Z(n7730) );
  AND U8363 ( .A(B[68]), .B(A[3]), .Z(n7537) );
  XNOR U8364 ( .A(n7527), .B(n7733), .Z(n7538) );
  XNOR U8365 ( .A(n7525), .B(n7528), .Z(n7733) );
  NAND U8366 ( .A(A[2]), .B(B[69]), .Z(n7528) );
  NANDN U8367 ( .A(n7734), .B(n7735), .Z(n7525) );
  AND U8368 ( .A(A[0]), .B(B[70]), .Z(n7735) );
  XOR U8369 ( .A(n7530), .B(n7736), .Z(n7527) );
  NAND U8370 ( .A(A[0]), .B(B[71]), .Z(n7736) );
  NAND U8371 ( .A(B[70]), .B(A[1]), .Z(n7530) );
  NAND U8372 ( .A(n7737), .B(n7738), .Z(n675) );
  NANDN U8373 ( .A(n7739), .B(n7740), .Z(n7738) );
  OR U8374 ( .A(n7741), .B(n7742), .Z(n7740) );
  NAND U8375 ( .A(n7742), .B(n7741), .Z(n7737) );
  XOR U8376 ( .A(n695), .B(n694), .Z(\A1[699] ) );
  XOR U8377 ( .A(n7708), .B(n7743), .Z(n694) );
  XNOR U8378 ( .A(n7707), .B(n7705), .Z(n7743) );
  AND U8379 ( .A(n7744), .B(n7745), .Z(n7705) );
  NANDN U8380 ( .A(n7746), .B(n7747), .Z(n7745) );
  NANDN U8381 ( .A(n7748), .B(n7749), .Z(n7747) );
  AND U8382 ( .A(B[698]), .B(A[3]), .Z(n7707) );
  XNOR U8383 ( .A(n7697), .B(n7750), .Z(n7708) );
  XNOR U8384 ( .A(n7695), .B(n7698), .Z(n7750) );
  NAND U8385 ( .A(A[2]), .B(B[699]), .Z(n7698) );
  NANDN U8386 ( .A(n7751), .B(n7752), .Z(n7695) );
  AND U8387 ( .A(A[0]), .B(B[700]), .Z(n7752) );
  XOR U8388 ( .A(n7700), .B(n7753), .Z(n7697) );
  NAND U8389 ( .A(A[0]), .B(B[701]), .Z(n7753) );
  NAND U8390 ( .A(B[700]), .B(A[1]), .Z(n7700) );
  NAND U8391 ( .A(n7754), .B(n7755), .Z(n695) );
  NANDN U8392 ( .A(n7756), .B(n7757), .Z(n7755) );
  OR U8393 ( .A(n7758), .B(n7759), .Z(n7757) );
  NAND U8394 ( .A(n7759), .B(n7758), .Z(n7754) );
  XOR U8395 ( .A(n701), .B(n700), .Z(\A1[698] ) );
  XOR U8396 ( .A(n7759), .B(n7760), .Z(n700) );
  XNOR U8397 ( .A(n7758), .B(n7756), .Z(n7760) );
  AND U8398 ( .A(n7761), .B(n7762), .Z(n7756) );
  NANDN U8399 ( .A(n7763), .B(n7764), .Z(n7762) );
  NANDN U8400 ( .A(n7765), .B(n7766), .Z(n7764) );
  AND U8401 ( .A(B[697]), .B(A[3]), .Z(n7758) );
  XNOR U8402 ( .A(n7748), .B(n7767), .Z(n7759) );
  XNOR U8403 ( .A(n7746), .B(n7749), .Z(n7767) );
  NAND U8404 ( .A(A[2]), .B(B[698]), .Z(n7749) );
  NANDN U8405 ( .A(n7768), .B(n7769), .Z(n7746) );
  AND U8406 ( .A(A[0]), .B(B[699]), .Z(n7769) );
  XOR U8407 ( .A(n7751), .B(n7770), .Z(n7748) );
  NAND U8408 ( .A(A[0]), .B(B[700]), .Z(n7770) );
  NAND U8409 ( .A(B[699]), .B(A[1]), .Z(n7751) );
  NAND U8410 ( .A(n7771), .B(n7772), .Z(n701) );
  NANDN U8411 ( .A(n7773), .B(n7774), .Z(n7772) );
  OR U8412 ( .A(n7775), .B(n7776), .Z(n7774) );
  NAND U8413 ( .A(n7776), .B(n7775), .Z(n7771) );
  XOR U8414 ( .A(n703), .B(n702), .Z(\A1[697] ) );
  XOR U8415 ( .A(n7776), .B(n7777), .Z(n702) );
  XNOR U8416 ( .A(n7775), .B(n7773), .Z(n7777) );
  AND U8417 ( .A(n7778), .B(n7779), .Z(n7773) );
  NANDN U8418 ( .A(n7780), .B(n7781), .Z(n7779) );
  NANDN U8419 ( .A(n7782), .B(n7783), .Z(n7781) );
  AND U8420 ( .A(B[696]), .B(A[3]), .Z(n7775) );
  XNOR U8421 ( .A(n7765), .B(n7784), .Z(n7776) );
  XNOR U8422 ( .A(n7763), .B(n7766), .Z(n7784) );
  NAND U8423 ( .A(A[2]), .B(B[697]), .Z(n7766) );
  NANDN U8424 ( .A(n7785), .B(n7786), .Z(n7763) );
  AND U8425 ( .A(A[0]), .B(B[698]), .Z(n7786) );
  XOR U8426 ( .A(n7768), .B(n7787), .Z(n7765) );
  NAND U8427 ( .A(A[0]), .B(B[699]), .Z(n7787) );
  NAND U8428 ( .A(B[698]), .B(A[1]), .Z(n7768) );
  NAND U8429 ( .A(n7788), .B(n7789), .Z(n703) );
  NANDN U8430 ( .A(n7790), .B(n7791), .Z(n7789) );
  OR U8431 ( .A(n7792), .B(n7793), .Z(n7791) );
  NAND U8432 ( .A(n7793), .B(n7792), .Z(n7788) );
  XOR U8433 ( .A(n705), .B(n704), .Z(\A1[696] ) );
  XOR U8434 ( .A(n7793), .B(n7794), .Z(n704) );
  XNOR U8435 ( .A(n7792), .B(n7790), .Z(n7794) );
  AND U8436 ( .A(n7795), .B(n7796), .Z(n7790) );
  NANDN U8437 ( .A(n7797), .B(n7798), .Z(n7796) );
  NANDN U8438 ( .A(n7799), .B(n7800), .Z(n7798) );
  AND U8439 ( .A(B[695]), .B(A[3]), .Z(n7792) );
  XNOR U8440 ( .A(n7782), .B(n7801), .Z(n7793) );
  XNOR U8441 ( .A(n7780), .B(n7783), .Z(n7801) );
  NAND U8442 ( .A(A[2]), .B(B[696]), .Z(n7783) );
  NANDN U8443 ( .A(n7802), .B(n7803), .Z(n7780) );
  AND U8444 ( .A(A[0]), .B(B[697]), .Z(n7803) );
  XOR U8445 ( .A(n7785), .B(n7804), .Z(n7782) );
  NAND U8446 ( .A(A[0]), .B(B[698]), .Z(n7804) );
  NAND U8447 ( .A(B[697]), .B(A[1]), .Z(n7785) );
  NAND U8448 ( .A(n7805), .B(n7806), .Z(n705) );
  NANDN U8449 ( .A(n7807), .B(n7808), .Z(n7806) );
  OR U8450 ( .A(n7809), .B(n7810), .Z(n7808) );
  NAND U8451 ( .A(n7810), .B(n7809), .Z(n7805) );
  XOR U8452 ( .A(n707), .B(n706), .Z(\A1[695] ) );
  XOR U8453 ( .A(n7810), .B(n7811), .Z(n706) );
  XNOR U8454 ( .A(n7809), .B(n7807), .Z(n7811) );
  AND U8455 ( .A(n7812), .B(n7813), .Z(n7807) );
  NANDN U8456 ( .A(n7814), .B(n7815), .Z(n7813) );
  NANDN U8457 ( .A(n7816), .B(n7817), .Z(n7815) );
  AND U8458 ( .A(B[694]), .B(A[3]), .Z(n7809) );
  XNOR U8459 ( .A(n7799), .B(n7818), .Z(n7810) );
  XNOR U8460 ( .A(n7797), .B(n7800), .Z(n7818) );
  NAND U8461 ( .A(A[2]), .B(B[695]), .Z(n7800) );
  NANDN U8462 ( .A(n7819), .B(n7820), .Z(n7797) );
  AND U8463 ( .A(A[0]), .B(B[696]), .Z(n7820) );
  XOR U8464 ( .A(n7802), .B(n7821), .Z(n7799) );
  NAND U8465 ( .A(A[0]), .B(B[697]), .Z(n7821) );
  NAND U8466 ( .A(B[696]), .B(A[1]), .Z(n7802) );
  NAND U8467 ( .A(n7822), .B(n7823), .Z(n707) );
  NANDN U8468 ( .A(n7824), .B(n7825), .Z(n7823) );
  OR U8469 ( .A(n7826), .B(n7827), .Z(n7825) );
  NAND U8470 ( .A(n7827), .B(n7826), .Z(n7822) );
  XOR U8471 ( .A(n709), .B(n708), .Z(\A1[694] ) );
  XOR U8472 ( .A(n7827), .B(n7828), .Z(n708) );
  XNOR U8473 ( .A(n7826), .B(n7824), .Z(n7828) );
  AND U8474 ( .A(n7829), .B(n7830), .Z(n7824) );
  NANDN U8475 ( .A(n7831), .B(n7832), .Z(n7830) );
  NANDN U8476 ( .A(n7833), .B(n7834), .Z(n7832) );
  AND U8477 ( .A(B[693]), .B(A[3]), .Z(n7826) );
  XNOR U8478 ( .A(n7816), .B(n7835), .Z(n7827) );
  XNOR U8479 ( .A(n7814), .B(n7817), .Z(n7835) );
  NAND U8480 ( .A(A[2]), .B(B[694]), .Z(n7817) );
  NANDN U8481 ( .A(n7836), .B(n7837), .Z(n7814) );
  AND U8482 ( .A(A[0]), .B(B[695]), .Z(n7837) );
  XOR U8483 ( .A(n7819), .B(n7838), .Z(n7816) );
  NAND U8484 ( .A(A[0]), .B(B[696]), .Z(n7838) );
  NAND U8485 ( .A(B[695]), .B(A[1]), .Z(n7819) );
  NAND U8486 ( .A(n7839), .B(n7840), .Z(n709) );
  NANDN U8487 ( .A(n7841), .B(n7842), .Z(n7840) );
  OR U8488 ( .A(n7843), .B(n7844), .Z(n7842) );
  NAND U8489 ( .A(n7844), .B(n7843), .Z(n7839) );
  XOR U8490 ( .A(n711), .B(n710), .Z(\A1[693] ) );
  XOR U8491 ( .A(n7844), .B(n7845), .Z(n710) );
  XNOR U8492 ( .A(n7843), .B(n7841), .Z(n7845) );
  AND U8493 ( .A(n7846), .B(n7847), .Z(n7841) );
  NANDN U8494 ( .A(n7848), .B(n7849), .Z(n7847) );
  NANDN U8495 ( .A(n7850), .B(n7851), .Z(n7849) );
  AND U8496 ( .A(B[692]), .B(A[3]), .Z(n7843) );
  XNOR U8497 ( .A(n7833), .B(n7852), .Z(n7844) );
  XNOR U8498 ( .A(n7831), .B(n7834), .Z(n7852) );
  NAND U8499 ( .A(A[2]), .B(B[693]), .Z(n7834) );
  NANDN U8500 ( .A(n7853), .B(n7854), .Z(n7831) );
  AND U8501 ( .A(A[0]), .B(B[694]), .Z(n7854) );
  XOR U8502 ( .A(n7836), .B(n7855), .Z(n7833) );
  NAND U8503 ( .A(A[0]), .B(B[695]), .Z(n7855) );
  NAND U8504 ( .A(B[694]), .B(A[1]), .Z(n7836) );
  NAND U8505 ( .A(n7856), .B(n7857), .Z(n711) );
  NANDN U8506 ( .A(n7858), .B(n7859), .Z(n7857) );
  OR U8507 ( .A(n7860), .B(n7861), .Z(n7859) );
  NAND U8508 ( .A(n7861), .B(n7860), .Z(n7856) );
  XOR U8509 ( .A(n713), .B(n712), .Z(\A1[692] ) );
  XOR U8510 ( .A(n7861), .B(n7862), .Z(n712) );
  XNOR U8511 ( .A(n7860), .B(n7858), .Z(n7862) );
  AND U8512 ( .A(n7863), .B(n7864), .Z(n7858) );
  NANDN U8513 ( .A(n7865), .B(n7866), .Z(n7864) );
  NANDN U8514 ( .A(n7867), .B(n7868), .Z(n7866) );
  AND U8515 ( .A(B[691]), .B(A[3]), .Z(n7860) );
  XNOR U8516 ( .A(n7850), .B(n7869), .Z(n7861) );
  XNOR U8517 ( .A(n7848), .B(n7851), .Z(n7869) );
  NAND U8518 ( .A(A[2]), .B(B[692]), .Z(n7851) );
  NANDN U8519 ( .A(n7870), .B(n7871), .Z(n7848) );
  AND U8520 ( .A(A[0]), .B(B[693]), .Z(n7871) );
  XOR U8521 ( .A(n7853), .B(n7872), .Z(n7850) );
  NAND U8522 ( .A(A[0]), .B(B[694]), .Z(n7872) );
  NAND U8523 ( .A(B[693]), .B(A[1]), .Z(n7853) );
  NAND U8524 ( .A(n7873), .B(n7874), .Z(n713) );
  NANDN U8525 ( .A(n7875), .B(n7876), .Z(n7874) );
  OR U8526 ( .A(n7877), .B(n7878), .Z(n7876) );
  NAND U8527 ( .A(n7878), .B(n7877), .Z(n7873) );
  XOR U8528 ( .A(n715), .B(n714), .Z(\A1[691] ) );
  XOR U8529 ( .A(n7878), .B(n7879), .Z(n714) );
  XNOR U8530 ( .A(n7877), .B(n7875), .Z(n7879) );
  AND U8531 ( .A(n7880), .B(n7881), .Z(n7875) );
  NANDN U8532 ( .A(n7882), .B(n7883), .Z(n7881) );
  NANDN U8533 ( .A(n7884), .B(n7885), .Z(n7883) );
  AND U8534 ( .A(B[690]), .B(A[3]), .Z(n7877) );
  XNOR U8535 ( .A(n7867), .B(n7886), .Z(n7878) );
  XNOR U8536 ( .A(n7865), .B(n7868), .Z(n7886) );
  NAND U8537 ( .A(A[2]), .B(B[691]), .Z(n7868) );
  NANDN U8538 ( .A(n7887), .B(n7888), .Z(n7865) );
  AND U8539 ( .A(A[0]), .B(B[692]), .Z(n7888) );
  XOR U8540 ( .A(n7870), .B(n7889), .Z(n7867) );
  NAND U8541 ( .A(A[0]), .B(B[693]), .Z(n7889) );
  NAND U8542 ( .A(B[692]), .B(A[1]), .Z(n7870) );
  NAND U8543 ( .A(n7890), .B(n7891), .Z(n715) );
  NANDN U8544 ( .A(n7892), .B(n7893), .Z(n7891) );
  OR U8545 ( .A(n7894), .B(n7895), .Z(n7893) );
  NAND U8546 ( .A(n7895), .B(n7894), .Z(n7890) );
  XOR U8547 ( .A(n717), .B(n716), .Z(\A1[690] ) );
  XOR U8548 ( .A(n7895), .B(n7896), .Z(n716) );
  XNOR U8549 ( .A(n7894), .B(n7892), .Z(n7896) );
  AND U8550 ( .A(n7897), .B(n7898), .Z(n7892) );
  NANDN U8551 ( .A(n7899), .B(n7900), .Z(n7898) );
  NANDN U8552 ( .A(n7901), .B(n7902), .Z(n7900) );
  AND U8553 ( .A(B[689]), .B(A[3]), .Z(n7894) );
  XNOR U8554 ( .A(n7884), .B(n7903), .Z(n7895) );
  XNOR U8555 ( .A(n7882), .B(n7885), .Z(n7903) );
  NAND U8556 ( .A(A[2]), .B(B[690]), .Z(n7885) );
  NANDN U8557 ( .A(n7904), .B(n7905), .Z(n7882) );
  AND U8558 ( .A(A[0]), .B(B[691]), .Z(n7905) );
  XOR U8559 ( .A(n7887), .B(n7906), .Z(n7884) );
  NAND U8560 ( .A(A[0]), .B(B[692]), .Z(n7906) );
  NAND U8561 ( .A(B[691]), .B(A[1]), .Z(n7887) );
  NAND U8562 ( .A(n7907), .B(n7908), .Z(n717) );
  NANDN U8563 ( .A(n7909), .B(n7910), .Z(n7908) );
  OR U8564 ( .A(n7911), .B(n7912), .Z(n7910) );
  NAND U8565 ( .A(n7912), .B(n7911), .Z(n7907) );
  XOR U8566 ( .A(n699), .B(n698), .Z(\A1[68] ) );
  XOR U8567 ( .A(n7742), .B(n7913), .Z(n698) );
  XNOR U8568 ( .A(n7741), .B(n7739), .Z(n7913) );
  AND U8569 ( .A(n7914), .B(n7915), .Z(n7739) );
  NANDN U8570 ( .A(n7916), .B(n7917), .Z(n7915) );
  NANDN U8571 ( .A(n7918), .B(n7919), .Z(n7917) );
  AND U8572 ( .A(B[67]), .B(A[3]), .Z(n7741) );
  XNOR U8573 ( .A(n7731), .B(n7920), .Z(n7742) );
  XNOR U8574 ( .A(n7729), .B(n7732), .Z(n7920) );
  NAND U8575 ( .A(A[2]), .B(B[68]), .Z(n7732) );
  NANDN U8576 ( .A(n7921), .B(n7922), .Z(n7729) );
  AND U8577 ( .A(A[0]), .B(B[69]), .Z(n7922) );
  XOR U8578 ( .A(n7734), .B(n7923), .Z(n7731) );
  NAND U8579 ( .A(A[0]), .B(B[70]), .Z(n7923) );
  NAND U8580 ( .A(B[69]), .B(A[1]), .Z(n7734) );
  NAND U8581 ( .A(n7924), .B(n7925), .Z(n699) );
  NANDN U8582 ( .A(n7926), .B(n7927), .Z(n7925) );
  OR U8583 ( .A(n7928), .B(n7929), .Z(n7927) );
  NAND U8584 ( .A(n7929), .B(n7928), .Z(n7924) );
  XOR U8585 ( .A(n719), .B(n718), .Z(\A1[689] ) );
  XOR U8586 ( .A(n7912), .B(n7930), .Z(n718) );
  XNOR U8587 ( .A(n7911), .B(n7909), .Z(n7930) );
  AND U8588 ( .A(n7931), .B(n7932), .Z(n7909) );
  NANDN U8589 ( .A(n7933), .B(n7934), .Z(n7932) );
  NANDN U8590 ( .A(n7935), .B(n7936), .Z(n7934) );
  AND U8591 ( .A(B[688]), .B(A[3]), .Z(n7911) );
  XNOR U8592 ( .A(n7901), .B(n7937), .Z(n7912) );
  XNOR U8593 ( .A(n7899), .B(n7902), .Z(n7937) );
  NAND U8594 ( .A(A[2]), .B(B[689]), .Z(n7902) );
  NANDN U8595 ( .A(n7938), .B(n7939), .Z(n7899) );
  AND U8596 ( .A(A[0]), .B(B[690]), .Z(n7939) );
  XOR U8597 ( .A(n7904), .B(n7940), .Z(n7901) );
  NAND U8598 ( .A(A[0]), .B(B[691]), .Z(n7940) );
  NAND U8599 ( .A(B[690]), .B(A[1]), .Z(n7904) );
  NAND U8600 ( .A(n7941), .B(n7942), .Z(n719) );
  NANDN U8601 ( .A(n7943), .B(n7944), .Z(n7942) );
  OR U8602 ( .A(n7945), .B(n7946), .Z(n7944) );
  NAND U8603 ( .A(n7946), .B(n7945), .Z(n7941) );
  XOR U8604 ( .A(n723), .B(n722), .Z(\A1[688] ) );
  XOR U8605 ( .A(n7946), .B(n7947), .Z(n722) );
  XNOR U8606 ( .A(n7945), .B(n7943), .Z(n7947) );
  AND U8607 ( .A(n7948), .B(n7949), .Z(n7943) );
  NANDN U8608 ( .A(n7950), .B(n7951), .Z(n7949) );
  NANDN U8609 ( .A(n7952), .B(n7953), .Z(n7951) );
  AND U8610 ( .A(B[687]), .B(A[3]), .Z(n7945) );
  XNOR U8611 ( .A(n7935), .B(n7954), .Z(n7946) );
  XNOR U8612 ( .A(n7933), .B(n7936), .Z(n7954) );
  NAND U8613 ( .A(A[2]), .B(B[688]), .Z(n7936) );
  NANDN U8614 ( .A(n7955), .B(n7956), .Z(n7933) );
  AND U8615 ( .A(A[0]), .B(B[689]), .Z(n7956) );
  XOR U8616 ( .A(n7938), .B(n7957), .Z(n7935) );
  NAND U8617 ( .A(A[0]), .B(B[690]), .Z(n7957) );
  NAND U8618 ( .A(B[689]), .B(A[1]), .Z(n7938) );
  NAND U8619 ( .A(n7958), .B(n7959), .Z(n723) );
  NANDN U8620 ( .A(n7960), .B(n7961), .Z(n7959) );
  OR U8621 ( .A(n7962), .B(n7963), .Z(n7961) );
  NAND U8622 ( .A(n7963), .B(n7962), .Z(n7958) );
  XOR U8623 ( .A(n725), .B(n724), .Z(\A1[687] ) );
  XOR U8624 ( .A(n7963), .B(n7964), .Z(n724) );
  XNOR U8625 ( .A(n7962), .B(n7960), .Z(n7964) );
  AND U8626 ( .A(n7965), .B(n7966), .Z(n7960) );
  NANDN U8627 ( .A(n7967), .B(n7968), .Z(n7966) );
  NANDN U8628 ( .A(n7969), .B(n7970), .Z(n7968) );
  AND U8629 ( .A(B[686]), .B(A[3]), .Z(n7962) );
  XNOR U8630 ( .A(n7952), .B(n7971), .Z(n7963) );
  XNOR U8631 ( .A(n7950), .B(n7953), .Z(n7971) );
  NAND U8632 ( .A(A[2]), .B(B[687]), .Z(n7953) );
  NANDN U8633 ( .A(n7972), .B(n7973), .Z(n7950) );
  AND U8634 ( .A(A[0]), .B(B[688]), .Z(n7973) );
  XOR U8635 ( .A(n7955), .B(n7974), .Z(n7952) );
  NAND U8636 ( .A(A[0]), .B(B[689]), .Z(n7974) );
  NAND U8637 ( .A(B[688]), .B(A[1]), .Z(n7955) );
  NAND U8638 ( .A(n7975), .B(n7976), .Z(n725) );
  NANDN U8639 ( .A(n7977), .B(n7978), .Z(n7976) );
  OR U8640 ( .A(n7979), .B(n7980), .Z(n7978) );
  NAND U8641 ( .A(n7980), .B(n7979), .Z(n7975) );
  XOR U8642 ( .A(n727), .B(n726), .Z(\A1[686] ) );
  XOR U8643 ( .A(n7980), .B(n7981), .Z(n726) );
  XNOR U8644 ( .A(n7979), .B(n7977), .Z(n7981) );
  AND U8645 ( .A(n7982), .B(n7983), .Z(n7977) );
  NANDN U8646 ( .A(n7984), .B(n7985), .Z(n7983) );
  NANDN U8647 ( .A(n7986), .B(n7987), .Z(n7985) );
  AND U8648 ( .A(B[685]), .B(A[3]), .Z(n7979) );
  XNOR U8649 ( .A(n7969), .B(n7988), .Z(n7980) );
  XNOR U8650 ( .A(n7967), .B(n7970), .Z(n7988) );
  NAND U8651 ( .A(A[2]), .B(B[686]), .Z(n7970) );
  NANDN U8652 ( .A(n7989), .B(n7990), .Z(n7967) );
  AND U8653 ( .A(A[0]), .B(B[687]), .Z(n7990) );
  XOR U8654 ( .A(n7972), .B(n7991), .Z(n7969) );
  NAND U8655 ( .A(A[0]), .B(B[688]), .Z(n7991) );
  NAND U8656 ( .A(B[687]), .B(A[1]), .Z(n7972) );
  NAND U8657 ( .A(n7992), .B(n7993), .Z(n727) );
  NANDN U8658 ( .A(n7994), .B(n7995), .Z(n7993) );
  OR U8659 ( .A(n7996), .B(n7997), .Z(n7995) );
  NAND U8660 ( .A(n7997), .B(n7996), .Z(n7992) );
  XOR U8661 ( .A(n729), .B(n728), .Z(\A1[685] ) );
  XOR U8662 ( .A(n7997), .B(n7998), .Z(n728) );
  XNOR U8663 ( .A(n7996), .B(n7994), .Z(n7998) );
  AND U8664 ( .A(n7999), .B(n8000), .Z(n7994) );
  NANDN U8665 ( .A(n8001), .B(n8002), .Z(n8000) );
  NANDN U8666 ( .A(n8003), .B(n8004), .Z(n8002) );
  AND U8667 ( .A(B[684]), .B(A[3]), .Z(n7996) );
  XNOR U8668 ( .A(n7986), .B(n8005), .Z(n7997) );
  XNOR U8669 ( .A(n7984), .B(n7987), .Z(n8005) );
  NAND U8670 ( .A(A[2]), .B(B[685]), .Z(n7987) );
  NANDN U8671 ( .A(n8006), .B(n8007), .Z(n7984) );
  AND U8672 ( .A(A[0]), .B(B[686]), .Z(n8007) );
  XOR U8673 ( .A(n7989), .B(n8008), .Z(n7986) );
  NAND U8674 ( .A(A[0]), .B(B[687]), .Z(n8008) );
  NAND U8675 ( .A(B[686]), .B(A[1]), .Z(n7989) );
  NAND U8676 ( .A(n8009), .B(n8010), .Z(n729) );
  NANDN U8677 ( .A(n8011), .B(n8012), .Z(n8010) );
  OR U8678 ( .A(n8013), .B(n8014), .Z(n8012) );
  NAND U8679 ( .A(n8014), .B(n8013), .Z(n8009) );
  XOR U8680 ( .A(n731), .B(n730), .Z(\A1[684] ) );
  XOR U8681 ( .A(n8014), .B(n8015), .Z(n730) );
  XNOR U8682 ( .A(n8013), .B(n8011), .Z(n8015) );
  AND U8683 ( .A(n8016), .B(n8017), .Z(n8011) );
  NANDN U8684 ( .A(n8018), .B(n8019), .Z(n8017) );
  NANDN U8685 ( .A(n8020), .B(n8021), .Z(n8019) );
  AND U8686 ( .A(B[683]), .B(A[3]), .Z(n8013) );
  XNOR U8687 ( .A(n8003), .B(n8022), .Z(n8014) );
  XNOR U8688 ( .A(n8001), .B(n8004), .Z(n8022) );
  NAND U8689 ( .A(A[2]), .B(B[684]), .Z(n8004) );
  NANDN U8690 ( .A(n8023), .B(n8024), .Z(n8001) );
  AND U8691 ( .A(A[0]), .B(B[685]), .Z(n8024) );
  XOR U8692 ( .A(n8006), .B(n8025), .Z(n8003) );
  NAND U8693 ( .A(A[0]), .B(B[686]), .Z(n8025) );
  NAND U8694 ( .A(B[685]), .B(A[1]), .Z(n8006) );
  NAND U8695 ( .A(n8026), .B(n8027), .Z(n731) );
  NANDN U8696 ( .A(n8028), .B(n8029), .Z(n8027) );
  OR U8697 ( .A(n8030), .B(n8031), .Z(n8029) );
  NAND U8698 ( .A(n8031), .B(n8030), .Z(n8026) );
  XOR U8699 ( .A(n733), .B(n732), .Z(\A1[683] ) );
  XOR U8700 ( .A(n8031), .B(n8032), .Z(n732) );
  XNOR U8701 ( .A(n8030), .B(n8028), .Z(n8032) );
  AND U8702 ( .A(n8033), .B(n8034), .Z(n8028) );
  NANDN U8703 ( .A(n8035), .B(n8036), .Z(n8034) );
  NANDN U8704 ( .A(n8037), .B(n8038), .Z(n8036) );
  AND U8705 ( .A(B[682]), .B(A[3]), .Z(n8030) );
  XNOR U8706 ( .A(n8020), .B(n8039), .Z(n8031) );
  XNOR U8707 ( .A(n8018), .B(n8021), .Z(n8039) );
  NAND U8708 ( .A(A[2]), .B(B[683]), .Z(n8021) );
  NANDN U8709 ( .A(n8040), .B(n8041), .Z(n8018) );
  AND U8710 ( .A(A[0]), .B(B[684]), .Z(n8041) );
  XOR U8711 ( .A(n8023), .B(n8042), .Z(n8020) );
  NAND U8712 ( .A(A[0]), .B(B[685]), .Z(n8042) );
  NAND U8713 ( .A(B[684]), .B(A[1]), .Z(n8023) );
  NAND U8714 ( .A(n8043), .B(n8044), .Z(n733) );
  NANDN U8715 ( .A(n8045), .B(n8046), .Z(n8044) );
  OR U8716 ( .A(n8047), .B(n8048), .Z(n8046) );
  NAND U8717 ( .A(n8048), .B(n8047), .Z(n8043) );
  XOR U8718 ( .A(n735), .B(n734), .Z(\A1[682] ) );
  XOR U8719 ( .A(n8048), .B(n8049), .Z(n734) );
  XNOR U8720 ( .A(n8047), .B(n8045), .Z(n8049) );
  AND U8721 ( .A(n8050), .B(n8051), .Z(n8045) );
  NANDN U8722 ( .A(n8052), .B(n8053), .Z(n8051) );
  NANDN U8723 ( .A(n8054), .B(n8055), .Z(n8053) );
  AND U8724 ( .A(B[681]), .B(A[3]), .Z(n8047) );
  XNOR U8725 ( .A(n8037), .B(n8056), .Z(n8048) );
  XNOR U8726 ( .A(n8035), .B(n8038), .Z(n8056) );
  NAND U8727 ( .A(A[2]), .B(B[682]), .Z(n8038) );
  NANDN U8728 ( .A(n8057), .B(n8058), .Z(n8035) );
  AND U8729 ( .A(A[0]), .B(B[683]), .Z(n8058) );
  XOR U8730 ( .A(n8040), .B(n8059), .Z(n8037) );
  NAND U8731 ( .A(A[0]), .B(B[684]), .Z(n8059) );
  NAND U8732 ( .A(B[683]), .B(A[1]), .Z(n8040) );
  NAND U8733 ( .A(n8060), .B(n8061), .Z(n735) );
  NANDN U8734 ( .A(n8062), .B(n8063), .Z(n8061) );
  OR U8735 ( .A(n8064), .B(n8065), .Z(n8063) );
  NAND U8736 ( .A(n8065), .B(n8064), .Z(n8060) );
  XOR U8737 ( .A(n737), .B(n736), .Z(\A1[681] ) );
  XOR U8738 ( .A(n8065), .B(n8066), .Z(n736) );
  XNOR U8739 ( .A(n8064), .B(n8062), .Z(n8066) );
  AND U8740 ( .A(n8067), .B(n8068), .Z(n8062) );
  NANDN U8741 ( .A(n8069), .B(n8070), .Z(n8068) );
  NANDN U8742 ( .A(n8071), .B(n8072), .Z(n8070) );
  AND U8743 ( .A(B[680]), .B(A[3]), .Z(n8064) );
  XNOR U8744 ( .A(n8054), .B(n8073), .Z(n8065) );
  XNOR U8745 ( .A(n8052), .B(n8055), .Z(n8073) );
  NAND U8746 ( .A(A[2]), .B(B[681]), .Z(n8055) );
  NANDN U8747 ( .A(n8074), .B(n8075), .Z(n8052) );
  AND U8748 ( .A(A[0]), .B(B[682]), .Z(n8075) );
  XOR U8749 ( .A(n8057), .B(n8076), .Z(n8054) );
  NAND U8750 ( .A(A[0]), .B(B[683]), .Z(n8076) );
  NAND U8751 ( .A(B[682]), .B(A[1]), .Z(n8057) );
  NAND U8752 ( .A(n8077), .B(n8078), .Z(n737) );
  NANDN U8753 ( .A(n8079), .B(n8080), .Z(n8078) );
  OR U8754 ( .A(n8081), .B(n8082), .Z(n8080) );
  NAND U8755 ( .A(n8082), .B(n8081), .Z(n8077) );
  XOR U8756 ( .A(n739), .B(n738), .Z(\A1[680] ) );
  XOR U8757 ( .A(n8082), .B(n8083), .Z(n738) );
  XNOR U8758 ( .A(n8081), .B(n8079), .Z(n8083) );
  AND U8759 ( .A(n8084), .B(n8085), .Z(n8079) );
  NANDN U8760 ( .A(n8086), .B(n8087), .Z(n8085) );
  NANDN U8761 ( .A(n8088), .B(n8089), .Z(n8087) );
  AND U8762 ( .A(B[679]), .B(A[3]), .Z(n8081) );
  XNOR U8763 ( .A(n8071), .B(n8090), .Z(n8082) );
  XNOR U8764 ( .A(n8069), .B(n8072), .Z(n8090) );
  NAND U8765 ( .A(A[2]), .B(B[680]), .Z(n8072) );
  NANDN U8766 ( .A(n8091), .B(n8092), .Z(n8069) );
  AND U8767 ( .A(A[0]), .B(B[681]), .Z(n8092) );
  XOR U8768 ( .A(n8074), .B(n8093), .Z(n8071) );
  NAND U8769 ( .A(A[0]), .B(B[682]), .Z(n8093) );
  NAND U8770 ( .A(B[681]), .B(A[1]), .Z(n8074) );
  NAND U8771 ( .A(n8094), .B(n8095), .Z(n739) );
  NANDN U8772 ( .A(n8096), .B(n8097), .Z(n8095) );
  OR U8773 ( .A(n8098), .B(n8099), .Z(n8097) );
  NAND U8774 ( .A(n8099), .B(n8098), .Z(n8094) );
  XOR U8775 ( .A(n721), .B(n720), .Z(\A1[67] ) );
  XOR U8776 ( .A(n7929), .B(n8100), .Z(n720) );
  XNOR U8777 ( .A(n7928), .B(n7926), .Z(n8100) );
  AND U8778 ( .A(n8101), .B(n8102), .Z(n7926) );
  NANDN U8779 ( .A(n8103), .B(n8104), .Z(n8102) );
  NANDN U8780 ( .A(n8105), .B(n8106), .Z(n8104) );
  AND U8781 ( .A(B[66]), .B(A[3]), .Z(n7928) );
  XNOR U8782 ( .A(n7918), .B(n8107), .Z(n7929) );
  XNOR U8783 ( .A(n7916), .B(n7919), .Z(n8107) );
  NAND U8784 ( .A(A[2]), .B(B[67]), .Z(n7919) );
  NANDN U8785 ( .A(n8108), .B(n8109), .Z(n7916) );
  AND U8786 ( .A(A[0]), .B(B[68]), .Z(n8109) );
  XOR U8787 ( .A(n7921), .B(n8110), .Z(n7918) );
  NAND U8788 ( .A(A[0]), .B(B[69]), .Z(n8110) );
  NAND U8789 ( .A(B[68]), .B(A[1]), .Z(n7921) );
  NAND U8790 ( .A(n8111), .B(n8112), .Z(n721) );
  NANDN U8791 ( .A(n8113), .B(n8114), .Z(n8112) );
  OR U8792 ( .A(n8115), .B(n8116), .Z(n8114) );
  NAND U8793 ( .A(n8116), .B(n8115), .Z(n8111) );
  XOR U8794 ( .A(n741), .B(n740), .Z(\A1[679] ) );
  XOR U8795 ( .A(n8099), .B(n8117), .Z(n740) );
  XNOR U8796 ( .A(n8098), .B(n8096), .Z(n8117) );
  AND U8797 ( .A(n8118), .B(n8119), .Z(n8096) );
  NANDN U8798 ( .A(n8120), .B(n8121), .Z(n8119) );
  NANDN U8799 ( .A(n8122), .B(n8123), .Z(n8121) );
  AND U8800 ( .A(B[678]), .B(A[3]), .Z(n8098) );
  XNOR U8801 ( .A(n8088), .B(n8124), .Z(n8099) );
  XNOR U8802 ( .A(n8086), .B(n8089), .Z(n8124) );
  NAND U8803 ( .A(A[2]), .B(B[679]), .Z(n8089) );
  NANDN U8804 ( .A(n8125), .B(n8126), .Z(n8086) );
  AND U8805 ( .A(A[0]), .B(B[680]), .Z(n8126) );
  XOR U8806 ( .A(n8091), .B(n8127), .Z(n8088) );
  NAND U8807 ( .A(A[0]), .B(B[681]), .Z(n8127) );
  NAND U8808 ( .A(B[680]), .B(A[1]), .Z(n8091) );
  NAND U8809 ( .A(n8128), .B(n8129), .Z(n741) );
  NANDN U8810 ( .A(n8130), .B(n8131), .Z(n8129) );
  OR U8811 ( .A(n8132), .B(n8133), .Z(n8131) );
  NAND U8812 ( .A(n8133), .B(n8132), .Z(n8128) );
  XOR U8813 ( .A(n745), .B(n744), .Z(\A1[678] ) );
  XOR U8814 ( .A(n8133), .B(n8134), .Z(n744) );
  XNOR U8815 ( .A(n8132), .B(n8130), .Z(n8134) );
  AND U8816 ( .A(n8135), .B(n8136), .Z(n8130) );
  NANDN U8817 ( .A(n8137), .B(n8138), .Z(n8136) );
  NANDN U8818 ( .A(n8139), .B(n8140), .Z(n8138) );
  AND U8819 ( .A(B[677]), .B(A[3]), .Z(n8132) );
  XNOR U8820 ( .A(n8122), .B(n8141), .Z(n8133) );
  XNOR U8821 ( .A(n8120), .B(n8123), .Z(n8141) );
  NAND U8822 ( .A(A[2]), .B(B[678]), .Z(n8123) );
  NANDN U8823 ( .A(n8142), .B(n8143), .Z(n8120) );
  AND U8824 ( .A(A[0]), .B(B[679]), .Z(n8143) );
  XOR U8825 ( .A(n8125), .B(n8144), .Z(n8122) );
  NAND U8826 ( .A(A[0]), .B(B[680]), .Z(n8144) );
  NAND U8827 ( .A(B[679]), .B(A[1]), .Z(n8125) );
  NAND U8828 ( .A(n8145), .B(n8146), .Z(n745) );
  NANDN U8829 ( .A(n8147), .B(n8148), .Z(n8146) );
  OR U8830 ( .A(n8149), .B(n8150), .Z(n8148) );
  NAND U8831 ( .A(n8150), .B(n8149), .Z(n8145) );
  XOR U8832 ( .A(n747), .B(n746), .Z(\A1[677] ) );
  XOR U8833 ( .A(n8150), .B(n8151), .Z(n746) );
  XNOR U8834 ( .A(n8149), .B(n8147), .Z(n8151) );
  AND U8835 ( .A(n8152), .B(n8153), .Z(n8147) );
  NANDN U8836 ( .A(n8154), .B(n8155), .Z(n8153) );
  NANDN U8837 ( .A(n8156), .B(n8157), .Z(n8155) );
  AND U8838 ( .A(B[676]), .B(A[3]), .Z(n8149) );
  XNOR U8839 ( .A(n8139), .B(n8158), .Z(n8150) );
  XNOR U8840 ( .A(n8137), .B(n8140), .Z(n8158) );
  NAND U8841 ( .A(A[2]), .B(B[677]), .Z(n8140) );
  NANDN U8842 ( .A(n8159), .B(n8160), .Z(n8137) );
  AND U8843 ( .A(A[0]), .B(B[678]), .Z(n8160) );
  XOR U8844 ( .A(n8142), .B(n8161), .Z(n8139) );
  NAND U8845 ( .A(A[0]), .B(B[679]), .Z(n8161) );
  NAND U8846 ( .A(B[678]), .B(A[1]), .Z(n8142) );
  NAND U8847 ( .A(n8162), .B(n8163), .Z(n747) );
  NANDN U8848 ( .A(n8164), .B(n8165), .Z(n8163) );
  OR U8849 ( .A(n8166), .B(n8167), .Z(n8165) );
  NAND U8850 ( .A(n8167), .B(n8166), .Z(n8162) );
  XOR U8851 ( .A(n749), .B(n748), .Z(\A1[676] ) );
  XOR U8852 ( .A(n8167), .B(n8168), .Z(n748) );
  XNOR U8853 ( .A(n8166), .B(n8164), .Z(n8168) );
  AND U8854 ( .A(n8169), .B(n8170), .Z(n8164) );
  NANDN U8855 ( .A(n8171), .B(n8172), .Z(n8170) );
  NANDN U8856 ( .A(n8173), .B(n8174), .Z(n8172) );
  AND U8857 ( .A(B[675]), .B(A[3]), .Z(n8166) );
  XNOR U8858 ( .A(n8156), .B(n8175), .Z(n8167) );
  XNOR U8859 ( .A(n8154), .B(n8157), .Z(n8175) );
  NAND U8860 ( .A(A[2]), .B(B[676]), .Z(n8157) );
  NANDN U8861 ( .A(n8176), .B(n8177), .Z(n8154) );
  AND U8862 ( .A(A[0]), .B(B[677]), .Z(n8177) );
  XOR U8863 ( .A(n8159), .B(n8178), .Z(n8156) );
  NAND U8864 ( .A(A[0]), .B(B[678]), .Z(n8178) );
  NAND U8865 ( .A(B[677]), .B(A[1]), .Z(n8159) );
  NAND U8866 ( .A(n8179), .B(n8180), .Z(n749) );
  NANDN U8867 ( .A(n8181), .B(n8182), .Z(n8180) );
  OR U8868 ( .A(n8183), .B(n8184), .Z(n8182) );
  NAND U8869 ( .A(n8184), .B(n8183), .Z(n8179) );
  XOR U8870 ( .A(n751), .B(n750), .Z(\A1[675] ) );
  XOR U8871 ( .A(n8184), .B(n8185), .Z(n750) );
  XNOR U8872 ( .A(n8183), .B(n8181), .Z(n8185) );
  AND U8873 ( .A(n8186), .B(n8187), .Z(n8181) );
  NANDN U8874 ( .A(n8188), .B(n8189), .Z(n8187) );
  NANDN U8875 ( .A(n8190), .B(n8191), .Z(n8189) );
  AND U8876 ( .A(B[674]), .B(A[3]), .Z(n8183) );
  XNOR U8877 ( .A(n8173), .B(n8192), .Z(n8184) );
  XNOR U8878 ( .A(n8171), .B(n8174), .Z(n8192) );
  NAND U8879 ( .A(A[2]), .B(B[675]), .Z(n8174) );
  NANDN U8880 ( .A(n8193), .B(n8194), .Z(n8171) );
  AND U8881 ( .A(A[0]), .B(B[676]), .Z(n8194) );
  XOR U8882 ( .A(n8176), .B(n8195), .Z(n8173) );
  NAND U8883 ( .A(A[0]), .B(B[677]), .Z(n8195) );
  NAND U8884 ( .A(B[676]), .B(A[1]), .Z(n8176) );
  NAND U8885 ( .A(n8196), .B(n8197), .Z(n751) );
  NANDN U8886 ( .A(n8198), .B(n8199), .Z(n8197) );
  OR U8887 ( .A(n8200), .B(n8201), .Z(n8199) );
  NAND U8888 ( .A(n8201), .B(n8200), .Z(n8196) );
  XOR U8889 ( .A(n753), .B(n752), .Z(\A1[674] ) );
  XOR U8890 ( .A(n8201), .B(n8202), .Z(n752) );
  XNOR U8891 ( .A(n8200), .B(n8198), .Z(n8202) );
  AND U8892 ( .A(n8203), .B(n8204), .Z(n8198) );
  NANDN U8893 ( .A(n8205), .B(n8206), .Z(n8204) );
  NANDN U8894 ( .A(n8207), .B(n8208), .Z(n8206) );
  AND U8895 ( .A(B[673]), .B(A[3]), .Z(n8200) );
  XNOR U8896 ( .A(n8190), .B(n8209), .Z(n8201) );
  XNOR U8897 ( .A(n8188), .B(n8191), .Z(n8209) );
  NAND U8898 ( .A(A[2]), .B(B[674]), .Z(n8191) );
  NANDN U8899 ( .A(n8210), .B(n8211), .Z(n8188) );
  AND U8900 ( .A(A[0]), .B(B[675]), .Z(n8211) );
  XOR U8901 ( .A(n8193), .B(n8212), .Z(n8190) );
  NAND U8902 ( .A(A[0]), .B(B[676]), .Z(n8212) );
  NAND U8903 ( .A(B[675]), .B(A[1]), .Z(n8193) );
  NAND U8904 ( .A(n8213), .B(n8214), .Z(n753) );
  NANDN U8905 ( .A(n8215), .B(n8216), .Z(n8214) );
  OR U8906 ( .A(n8217), .B(n8218), .Z(n8216) );
  NAND U8907 ( .A(n8218), .B(n8217), .Z(n8213) );
  XOR U8908 ( .A(n755), .B(n754), .Z(\A1[673] ) );
  XOR U8909 ( .A(n8218), .B(n8219), .Z(n754) );
  XNOR U8910 ( .A(n8217), .B(n8215), .Z(n8219) );
  AND U8911 ( .A(n8220), .B(n8221), .Z(n8215) );
  NANDN U8912 ( .A(n8222), .B(n8223), .Z(n8221) );
  NANDN U8913 ( .A(n8224), .B(n8225), .Z(n8223) );
  AND U8914 ( .A(B[672]), .B(A[3]), .Z(n8217) );
  XNOR U8915 ( .A(n8207), .B(n8226), .Z(n8218) );
  XNOR U8916 ( .A(n8205), .B(n8208), .Z(n8226) );
  NAND U8917 ( .A(A[2]), .B(B[673]), .Z(n8208) );
  NANDN U8918 ( .A(n8227), .B(n8228), .Z(n8205) );
  AND U8919 ( .A(A[0]), .B(B[674]), .Z(n8228) );
  XOR U8920 ( .A(n8210), .B(n8229), .Z(n8207) );
  NAND U8921 ( .A(A[0]), .B(B[675]), .Z(n8229) );
  NAND U8922 ( .A(B[674]), .B(A[1]), .Z(n8210) );
  NAND U8923 ( .A(n8230), .B(n8231), .Z(n755) );
  NANDN U8924 ( .A(n8232), .B(n8233), .Z(n8231) );
  OR U8925 ( .A(n8234), .B(n8235), .Z(n8233) );
  NAND U8926 ( .A(n8235), .B(n8234), .Z(n8230) );
  XOR U8927 ( .A(n757), .B(n756), .Z(\A1[672] ) );
  XOR U8928 ( .A(n8235), .B(n8236), .Z(n756) );
  XNOR U8929 ( .A(n8234), .B(n8232), .Z(n8236) );
  AND U8930 ( .A(n8237), .B(n8238), .Z(n8232) );
  NANDN U8931 ( .A(n8239), .B(n8240), .Z(n8238) );
  NANDN U8932 ( .A(n8241), .B(n8242), .Z(n8240) );
  AND U8933 ( .A(B[671]), .B(A[3]), .Z(n8234) );
  XNOR U8934 ( .A(n8224), .B(n8243), .Z(n8235) );
  XNOR U8935 ( .A(n8222), .B(n8225), .Z(n8243) );
  NAND U8936 ( .A(A[2]), .B(B[672]), .Z(n8225) );
  NANDN U8937 ( .A(n8244), .B(n8245), .Z(n8222) );
  AND U8938 ( .A(A[0]), .B(B[673]), .Z(n8245) );
  XOR U8939 ( .A(n8227), .B(n8246), .Z(n8224) );
  NAND U8940 ( .A(A[0]), .B(B[674]), .Z(n8246) );
  NAND U8941 ( .A(B[673]), .B(A[1]), .Z(n8227) );
  NAND U8942 ( .A(n8247), .B(n8248), .Z(n757) );
  NANDN U8943 ( .A(n8249), .B(n8250), .Z(n8248) );
  OR U8944 ( .A(n8251), .B(n8252), .Z(n8250) );
  NAND U8945 ( .A(n8252), .B(n8251), .Z(n8247) );
  XOR U8946 ( .A(n759), .B(n758), .Z(\A1[671] ) );
  XOR U8947 ( .A(n8252), .B(n8253), .Z(n758) );
  XNOR U8948 ( .A(n8251), .B(n8249), .Z(n8253) );
  AND U8949 ( .A(n8254), .B(n8255), .Z(n8249) );
  NANDN U8950 ( .A(n8256), .B(n8257), .Z(n8255) );
  NANDN U8951 ( .A(n8258), .B(n8259), .Z(n8257) );
  AND U8952 ( .A(B[670]), .B(A[3]), .Z(n8251) );
  XNOR U8953 ( .A(n8241), .B(n8260), .Z(n8252) );
  XNOR U8954 ( .A(n8239), .B(n8242), .Z(n8260) );
  NAND U8955 ( .A(A[2]), .B(B[671]), .Z(n8242) );
  NANDN U8956 ( .A(n8261), .B(n8262), .Z(n8239) );
  AND U8957 ( .A(A[0]), .B(B[672]), .Z(n8262) );
  XOR U8958 ( .A(n8244), .B(n8263), .Z(n8241) );
  NAND U8959 ( .A(A[0]), .B(B[673]), .Z(n8263) );
  NAND U8960 ( .A(B[672]), .B(A[1]), .Z(n8244) );
  NAND U8961 ( .A(n8264), .B(n8265), .Z(n759) );
  NANDN U8962 ( .A(n8266), .B(n8267), .Z(n8265) );
  OR U8963 ( .A(n8268), .B(n8269), .Z(n8267) );
  NAND U8964 ( .A(n8269), .B(n8268), .Z(n8264) );
  XOR U8965 ( .A(n761), .B(n760), .Z(\A1[670] ) );
  XOR U8966 ( .A(n8269), .B(n8270), .Z(n760) );
  XNOR U8967 ( .A(n8268), .B(n8266), .Z(n8270) );
  AND U8968 ( .A(n8271), .B(n8272), .Z(n8266) );
  NANDN U8969 ( .A(n8273), .B(n8274), .Z(n8272) );
  NANDN U8970 ( .A(n8275), .B(n8276), .Z(n8274) );
  AND U8971 ( .A(B[669]), .B(A[3]), .Z(n8268) );
  XNOR U8972 ( .A(n8258), .B(n8277), .Z(n8269) );
  XNOR U8973 ( .A(n8256), .B(n8259), .Z(n8277) );
  NAND U8974 ( .A(A[2]), .B(B[670]), .Z(n8259) );
  NANDN U8975 ( .A(n8278), .B(n8279), .Z(n8256) );
  AND U8976 ( .A(A[0]), .B(B[671]), .Z(n8279) );
  XOR U8977 ( .A(n8261), .B(n8280), .Z(n8258) );
  NAND U8978 ( .A(A[0]), .B(B[672]), .Z(n8280) );
  NAND U8979 ( .A(B[671]), .B(A[1]), .Z(n8261) );
  NAND U8980 ( .A(n8281), .B(n8282), .Z(n761) );
  NANDN U8981 ( .A(n8283), .B(n8284), .Z(n8282) );
  OR U8982 ( .A(n8285), .B(n8286), .Z(n8284) );
  NAND U8983 ( .A(n8286), .B(n8285), .Z(n8281) );
  XOR U8984 ( .A(n743), .B(n742), .Z(\A1[66] ) );
  XOR U8985 ( .A(n8116), .B(n8287), .Z(n742) );
  XNOR U8986 ( .A(n8115), .B(n8113), .Z(n8287) );
  AND U8987 ( .A(n8288), .B(n8289), .Z(n8113) );
  NANDN U8988 ( .A(n8290), .B(n8291), .Z(n8289) );
  NANDN U8989 ( .A(n8292), .B(n8293), .Z(n8291) );
  AND U8990 ( .A(B[65]), .B(A[3]), .Z(n8115) );
  XNOR U8991 ( .A(n8105), .B(n8294), .Z(n8116) );
  XNOR U8992 ( .A(n8103), .B(n8106), .Z(n8294) );
  NAND U8993 ( .A(A[2]), .B(B[66]), .Z(n8106) );
  NANDN U8994 ( .A(n8295), .B(n8296), .Z(n8103) );
  AND U8995 ( .A(A[0]), .B(B[67]), .Z(n8296) );
  XOR U8996 ( .A(n8108), .B(n8297), .Z(n8105) );
  NAND U8997 ( .A(A[0]), .B(B[68]), .Z(n8297) );
  NAND U8998 ( .A(B[67]), .B(A[1]), .Z(n8108) );
  NAND U8999 ( .A(n8298), .B(n8299), .Z(n743) );
  NANDN U9000 ( .A(n8300), .B(n8301), .Z(n8299) );
  OR U9001 ( .A(n8302), .B(n8303), .Z(n8301) );
  NAND U9002 ( .A(n8303), .B(n8302), .Z(n8298) );
  XOR U9003 ( .A(n763), .B(n762), .Z(\A1[669] ) );
  XOR U9004 ( .A(n8286), .B(n8304), .Z(n762) );
  XNOR U9005 ( .A(n8285), .B(n8283), .Z(n8304) );
  AND U9006 ( .A(n8305), .B(n8306), .Z(n8283) );
  NANDN U9007 ( .A(n8307), .B(n8308), .Z(n8306) );
  NANDN U9008 ( .A(n8309), .B(n8310), .Z(n8308) );
  AND U9009 ( .A(B[668]), .B(A[3]), .Z(n8285) );
  XNOR U9010 ( .A(n8275), .B(n8311), .Z(n8286) );
  XNOR U9011 ( .A(n8273), .B(n8276), .Z(n8311) );
  NAND U9012 ( .A(A[2]), .B(B[669]), .Z(n8276) );
  NANDN U9013 ( .A(n8312), .B(n8313), .Z(n8273) );
  AND U9014 ( .A(A[0]), .B(B[670]), .Z(n8313) );
  XOR U9015 ( .A(n8278), .B(n8314), .Z(n8275) );
  NAND U9016 ( .A(A[0]), .B(B[671]), .Z(n8314) );
  NAND U9017 ( .A(B[670]), .B(A[1]), .Z(n8278) );
  NAND U9018 ( .A(n8315), .B(n8316), .Z(n763) );
  NANDN U9019 ( .A(n8317), .B(n8318), .Z(n8316) );
  OR U9020 ( .A(n8319), .B(n8320), .Z(n8318) );
  NAND U9021 ( .A(n8320), .B(n8319), .Z(n8315) );
  XOR U9022 ( .A(n767), .B(n766), .Z(\A1[668] ) );
  XOR U9023 ( .A(n8320), .B(n8321), .Z(n766) );
  XNOR U9024 ( .A(n8319), .B(n8317), .Z(n8321) );
  AND U9025 ( .A(n8322), .B(n8323), .Z(n8317) );
  NANDN U9026 ( .A(n8324), .B(n8325), .Z(n8323) );
  NANDN U9027 ( .A(n8326), .B(n8327), .Z(n8325) );
  AND U9028 ( .A(B[667]), .B(A[3]), .Z(n8319) );
  XNOR U9029 ( .A(n8309), .B(n8328), .Z(n8320) );
  XNOR U9030 ( .A(n8307), .B(n8310), .Z(n8328) );
  NAND U9031 ( .A(A[2]), .B(B[668]), .Z(n8310) );
  NANDN U9032 ( .A(n8329), .B(n8330), .Z(n8307) );
  AND U9033 ( .A(A[0]), .B(B[669]), .Z(n8330) );
  XOR U9034 ( .A(n8312), .B(n8331), .Z(n8309) );
  NAND U9035 ( .A(A[0]), .B(B[670]), .Z(n8331) );
  NAND U9036 ( .A(B[669]), .B(A[1]), .Z(n8312) );
  NAND U9037 ( .A(n8332), .B(n8333), .Z(n767) );
  NANDN U9038 ( .A(n8334), .B(n8335), .Z(n8333) );
  OR U9039 ( .A(n8336), .B(n8337), .Z(n8335) );
  NAND U9040 ( .A(n8337), .B(n8336), .Z(n8332) );
  XOR U9041 ( .A(n769), .B(n768), .Z(\A1[667] ) );
  XOR U9042 ( .A(n8337), .B(n8338), .Z(n768) );
  XNOR U9043 ( .A(n8336), .B(n8334), .Z(n8338) );
  AND U9044 ( .A(n8339), .B(n8340), .Z(n8334) );
  NANDN U9045 ( .A(n8341), .B(n8342), .Z(n8340) );
  NANDN U9046 ( .A(n8343), .B(n8344), .Z(n8342) );
  AND U9047 ( .A(B[666]), .B(A[3]), .Z(n8336) );
  XNOR U9048 ( .A(n8326), .B(n8345), .Z(n8337) );
  XNOR U9049 ( .A(n8324), .B(n8327), .Z(n8345) );
  NAND U9050 ( .A(A[2]), .B(B[667]), .Z(n8327) );
  NANDN U9051 ( .A(n8346), .B(n8347), .Z(n8324) );
  AND U9052 ( .A(A[0]), .B(B[668]), .Z(n8347) );
  XOR U9053 ( .A(n8329), .B(n8348), .Z(n8326) );
  NAND U9054 ( .A(A[0]), .B(B[669]), .Z(n8348) );
  NAND U9055 ( .A(B[668]), .B(A[1]), .Z(n8329) );
  NAND U9056 ( .A(n8349), .B(n8350), .Z(n769) );
  NANDN U9057 ( .A(n8351), .B(n8352), .Z(n8350) );
  OR U9058 ( .A(n8353), .B(n8354), .Z(n8352) );
  NAND U9059 ( .A(n8354), .B(n8353), .Z(n8349) );
  XOR U9060 ( .A(n771), .B(n770), .Z(\A1[666] ) );
  XOR U9061 ( .A(n8354), .B(n8355), .Z(n770) );
  XNOR U9062 ( .A(n8353), .B(n8351), .Z(n8355) );
  AND U9063 ( .A(n8356), .B(n8357), .Z(n8351) );
  NANDN U9064 ( .A(n8358), .B(n8359), .Z(n8357) );
  NANDN U9065 ( .A(n8360), .B(n8361), .Z(n8359) );
  AND U9066 ( .A(B[665]), .B(A[3]), .Z(n8353) );
  XNOR U9067 ( .A(n8343), .B(n8362), .Z(n8354) );
  XNOR U9068 ( .A(n8341), .B(n8344), .Z(n8362) );
  NAND U9069 ( .A(A[2]), .B(B[666]), .Z(n8344) );
  NANDN U9070 ( .A(n8363), .B(n8364), .Z(n8341) );
  AND U9071 ( .A(A[0]), .B(B[667]), .Z(n8364) );
  XOR U9072 ( .A(n8346), .B(n8365), .Z(n8343) );
  NAND U9073 ( .A(A[0]), .B(B[668]), .Z(n8365) );
  NAND U9074 ( .A(B[667]), .B(A[1]), .Z(n8346) );
  NAND U9075 ( .A(n8366), .B(n8367), .Z(n771) );
  NANDN U9076 ( .A(n8368), .B(n8369), .Z(n8367) );
  OR U9077 ( .A(n8370), .B(n8371), .Z(n8369) );
  NAND U9078 ( .A(n8371), .B(n8370), .Z(n8366) );
  XOR U9079 ( .A(n773), .B(n772), .Z(\A1[665] ) );
  XOR U9080 ( .A(n8371), .B(n8372), .Z(n772) );
  XNOR U9081 ( .A(n8370), .B(n8368), .Z(n8372) );
  AND U9082 ( .A(n8373), .B(n8374), .Z(n8368) );
  NANDN U9083 ( .A(n8375), .B(n8376), .Z(n8374) );
  NANDN U9084 ( .A(n8377), .B(n8378), .Z(n8376) );
  AND U9085 ( .A(B[664]), .B(A[3]), .Z(n8370) );
  XNOR U9086 ( .A(n8360), .B(n8379), .Z(n8371) );
  XNOR U9087 ( .A(n8358), .B(n8361), .Z(n8379) );
  NAND U9088 ( .A(A[2]), .B(B[665]), .Z(n8361) );
  NANDN U9089 ( .A(n8380), .B(n8381), .Z(n8358) );
  AND U9090 ( .A(A[0]), .B(B[666]), .Z(n8381) );
  XOR U9091 ( .A(n8363), .B(n8382), .Z(n8360) );
  NAND U9092 ( .A(A[0]), .B(B[667]), .Z(n8382) );
  NAND U9093 ( .A(B[666]), .B(A[1]), .Z(n8363) );
  NAND U9094 ( .A(n8383), .B(n8384), .Z(n773) );
  NANDN U9095 ( .A(n8385), .B(n8386), .Z(n8384) );
  OR U9096 ( .A(n8387), .B(n8388), .Z(n8386) );
  NAND U9097 ( .A(n8388), .B(n8387), .Z(n8383) );
  XOR U9098 ( .A(n775), .B(n774), .Z(\A1[664] ) );
  XOR U9099 ( .A(n8388), .B(n8389), .Z(n774) );
  XNOR U9100 ( .A(n8387), .B(n8385), .Z(n8389) );
  AND U9101 ( .A(n8390), .B(n8391), .Z(n8385) );
  NANDN U9102 ( .A(n8392), .B(n8393), .Z(n8391) );
  NANDN U9103 ( .A(n8394), .B(n8395), .Z(n8393) );
  AND U9104 ( .A(B[663]), .B(A[3]), .Z(n8387) );
  XNOR U9105 ( .A(n8377), .B(n8396), .Z(n8388) );
  XNOR U9106 ( .A(n8375), .B(n8378), .Z(n8396) );
  NAND U9107 ( .A(A[2]), .B(B[664]), .Z(n8378) );
  NANDN U9108 ( .A(n8397), .B(n8398), .Z(n8375) );
  AND U9109 ( .A(A[0]), .B(B[665]), .Z(n8398) );
  XOR U9110 ( .A(n8380), .B(n8399), .Z(n8377) );
  NAND U9111 ( .A(A[0]), .B(B[666]), .Z(n8399) );
  NAND U9112 ( .A(B[665]), .B(A[1]), .Z(n8380) );
  NAND U9113 ( .A(n8400), .B(n8401), .Z(n775) );
  NANDN U9114 ( .A(n8402), .B(n8403), .Z(n8401) );
  OR U9115 ( .A(n8404), .B(n8405), .Z(n8403) );
  NAND U9116 ( .A(n8405), .B(n8404), .Z(n8400) );
  XOR U9117 ( .A(n777), .B(n776), .Z(\A1[663] ) );
  XOR U9118 ( .A(n8405), .B(n8406), .Z(n776) );
  XNOR U9119 ( .A(n8404), .B(n8402), .Z(n8406) );
  AND U9120 ( .A(n8407), .B(n8408), .Z(n8402) );
  NANDN U9121 ( .A(n8409), .B(n8410), .Z(n8408) );
  NANDN U9122 ( .A(n8411), .B(n8412), .Z(n8410) );
  AND U9123 ( .A(B[662]), .B(A[3]), .Z(n8404) );
  XNOR U9124 ( .A(n8394), .B(n8413), .Z(n8405) );
  XNOR U9125 ( .A(n8392), .B(n8395), .Z(n8413) );
  NAND U9126 ( .A(A[2]), .B(B[663]), .Z(n8395) );
  NANDN U9127 ( .A(n8414), .B(n8415), .Z(n8392) );
  AND U9128 ( .A(A[0]), .B(B[664]), .Z(n8415) );
  XOR U9129 ( .A(n8397), .B(n8416), .Z(n8394) );
  NAND U9130 ( .A(A[0]), .B(B[665]), .Z(n8416) );
  NAND U9131 ( .A(B[664]), .B(A[1]), .Z(n8397) );
  NAND U9132 ( .A(n8417), .B(n8418), .Z(n777) );
  NANDN U9133 ( .A(n8419), .B(n8420), .Z(n8418) );
  OR U9134 ( .A(n8421), .B(n8422), .Z(n8420) );
  NAND U9135 ( .A(n8422), .B(n8421), .Z(n8417) );
  XOR U9136 ( .A(n779), .B(n778), .Z(\A1[662] ) );
  XOR U9137 ( .A(n8422), .B(n8423), .Z(n778) );
  XNOR U9138 ( .A(n8421), .B(n8419), .Z(n8423) );
  AND U9139 ( .A(n8424), .B(n8425), .Z(n8419) );
  NANDN U9140 ( .A(n8426), .B(n8427), .Z(n8425) );
  NANDN U9141 ( .A(n8428), .B(n8429), .Z(n8427) );
  AND U9142 ( .A(B[661]), .B(A[3]), .Z(n8421) );
  XNOR U9143 ( .A(n8411), .B(n8430), .Z(n8422) );
  XNOR U9144 ( .A(n8409), .B(n8412), .Z(n8430) );
  NAND U9145 ( .A(A[2]), .B(B[662]), .Z(n8412) );
  NANDN U9146 ( .A(n8431), .B(n8432), .Z(n8409) );
  AND U9147 ( .A(A[0]), .B(B[663]), .Z(n8432) );
  XOR U9148 ( .A(n8414), .B(n8433), .Z(n8411) );
  NAND U9149 ( .A(A[0]), .B(B[664]), .Z(n8433) );
  NAND U9150 ( .A(B[663]), .B(A[1]), .Z(n8414) );
  NAND U9151 ( .A(n8434), .B(n8435), .Z(n779) );
  NANDN U9152 ( .A(n8436), .B(n8437), .Z(n8435) );
  OR U9153 ( .A(n8438), .B(n8439), .Z(n8437) );
  NAND U9154 ( .A(n8439), .B(n8438), .Z(n8434) );
  XOR U9155 ( .A(n781), .B(n780), .Z(\A1[661] ) );
  XOR U9156 ( .A(n8439), .B(n8440), .Z(n780) );
  XNOR U9157 ( .A(n8438), .B(n8436), .Z(n8440) );
  AND U9158 ( .A(n8441), .B(n8442), .Z(n8436) );
  NANDN U9159 ( .A(n8443), .B(n8444), .Z(n8442) );
  NANDN U9160 ( .A(n8445), .B(n8446), .Z(n8444) );
  AND U9161 ( .A(B[660]), .B(A[3]), .Z(n8438) );
  XNOR U9162 ( .A(n8428), .B(n8447), .Z(n8439) );
  XNOR U9163 ( .A(n8426), .B(n8429), .Z(n8447) );
  NAND U9164 ( .A(A[2]), .B(B[661]), .Z(n8429) );
  NANDN U9165 ( .A(n8448), .B(n8449), .Z(n8426) );
  AND U9166 ( .A(A[0]), .B(B[662]), .Z(n8449) );
  XOR U9167 ( .A(n8431), .B(n8450), .Z(n8428) );
  NAND U9168 ( .A(A[0]), .B(B[663]), .Z(n8450) );
  NAND U9169 ( .A(B[662]), .B(A[1]), .Z(n8431) );
  NAND U9170 ( .A(n8451), .B(n8452), .Z(n781) );
  NANDN U9171 ( .A(n8453), .B(n8454), .Z(n8452) );
  OR U9172 ( .A(n8455), .B(n8456), .Z(n8454) );
  NAND U9173 ( .A(n8456), .B(n8455), .Z(n8451) );
  XOR U9174 ( .A(n783), .B(n782), .Z(\A1[660] ) );
  XOR U9175 ( .A(n8456), .B(n8457), .Z(n782) );
  XNOR U9176 ( .A(n8455), .B(n8453), .Z(n8457) );
  AND U9177 ( .A(n8458), .B(n8459), .Z(n8453) );
  NANDN U9178 ( .A(n8460), .B(n8461), .Z(n8459) );
  NANDN U9179 ( .A(n8462), .B(n8463), .Z(n8461) );
  AND U9180 ( .A(B[659]), .B(A[3]), .Z(n8455) );
  XNOR U9181 ( .A(n8445), .B(n8464), .Z(n8456) );
  XNOR U9182 ( .A(n8443), .B(n8446), .Z(n8464) );
  NAND U9183 ( .A(A[2]), .B(B[660]), .Z(n8446) );
  NANDN U9184 ( .A(n8465), .B(n8466), .Z(n8443) );
  AND U9185 ( .A(A[0]), .B(B[661]), .Z(n8466) );
  XOR U9186 ( .A(n8448), .B(n8467), .Z(n8445) );
  NAND U9187 ( .A(A[0]), .B(B[662]), .Z(n8467) );
  NAND U9188 ( .A(B[661]), .B(A[1]), .Z(n8448) );
  NAND U9189 ( .A(n8468), .B(n8469), .Z(n783) );
  NANDN U9190 ( .A(n8470), .B(n8471), .Z(n8469) );
  OR U9191 ( .A(n8472), .B(n8473), .Z(n8471) );
  NAND U9192 ( .A(n8473), .B(n8472), .Z(n8468) );
  XOR U9193 ( .A(n765), .B(n764), .Z(\A1[65] ) );
  XOR U9194 ( .A(n8303), .B(n8474), .Z(n764) );
  XNOR U9195 ( .A(n8302), .B(n8300), .Z(n8474) );
  AND U9196 ( .A(n8475), .B(n8476), .Z(n8300) );
  NANDN U9197 ( .A(n8477), .B(n8478), .Z(n8476) );
  NANDN U9198 ( .A(n8479), .B(n8480), .Z(n8478) );
  AND U9199 ( .A(B[64]), .B(A[3]), .Z(n8302) );
  XNOR U9200 ( .A(n8292), .B(n8481), .Z(n8303) );
  XNOR U9201 ( .A(n8290), .B(n8293), .Z(n8481) );
  NAND U9202 ( .A(A[2]), .B(B[65]), .Z(n8293) );
  NANDN U9203 ( .A(n8482), .B(n8483), .Z(n8290) );
  AND U9204 ( .A(A[0]), .B(B[66]), .Z(n8483) );
  XOR U9205 ( .A(n8295), .B(n8484), .Z(n8292) );
  NAND U9206 ( .A(A[0]), .B(B[67]), .Z(n8484) );
  NAND U9207 ( .A(B[66]), .B(A[1]), .Z(n8295) );
  NAND U9208 ( .A(n8485), .B(n8486), .Z(n765) );
  NANDN U9209 ( .A(n8487), .B(n8488), .Z(n8486) );
  OR U9210 ( .A(n8489), .B(n8490), .Z(n8488) );
  NAND U9211 ( .A(n8490), .B(n8489), .Z(n8485) );
  XOR U9212 ( .A(n785), .B(n784), .Z(\A1[659] ) );
  XOR U9213 ( .A(n8473), .B(n8491), .Z(n784) );
  XNOR U9214 ( .A(n8472), .B(n8470), .Z(n8491) );
  AND U9215 ( .A(n8492), .B(n8493), .Z(n8470) );
  NANDN U9216 ( .A(n8494), .B(n8495), .Z(n8493) );
  NANDN U9217 ( .A(n8496), .B(n8497), .Z(n8495) );
  AND U9218 ( .A(B[658]), .B(A[3]), .Z(n8472) );
  XNOR U9219 ( .A(n8462), .B(n8498), .Z(n8473) );
  XNOR U9220 ( .A(n8460), .B(n8463), .Z(n8498) );
  NAND U9221 ( .A(A[2]), .B(B[659]), .Z(n8463) );
  NANDN U9222 ( .A(n8499), .B(n8500), .Z(n8460) );
  AND U9223 ( .A(A[0]), .B(B[660]), .Z(n8500) );
  XOR U9224 ( .A(n8465), .B(n8501), .Z(n8462) );
  NAND U9225 ( .A(A[0]), .B(B[661]), .Z(n8501) );
  NAND U9226 ( .A(B[660]), .B(A[1]), .Z(n8465) );
  NAND U9227 ( .A(n8502), .B(n8503), .Z(n785) );
  NANDN U9228 ( .A(n8504), .B(n8505), .Z(n8503) );
  OR U9229 ( .A(n8506), .B(n8507), .Z(n8505) );
  NAND U9230 ( .A(n8507), .B(n8506), .Z(n8502) );
  XOR U9231 ( .A(n789), .B(n788), .Z(\A1[658] ) );
  XOR U9232 ( .A(n8507), .B(n8508), .Z(n788) );
  XNOR U9233 ( .A(n8506), .B(n8504), .Z(n8508) );
  AND U9234 ( .A(n8509), .B(n8510), .Z(n8504) );
  NANDN U9235 ( .A(n8511), .B(n8512), .Z(n8510) );
  NANDN U9236 ( .A(n8513), .B(n8514), .Z(n8512) );
  AND U9237 ( .A(B[657]), .B(A[3]), .Z(n8506) );
  XNOR U9238 ( .A(n8496), .B(n8515), .Z(n8507) );
  XNOR U9239 ( .A(n8494), .B(n8497), .Z(n8515) );
  NAND U9240 ( .A(A[2]), .B(B[658]), .Z(n8497) );
  NANDN U9241 ( .A(n8516), .B(n8517), .Z(n8494) );
  AND U9242 ( .A(A[0]), .B(B[659]), .Z(n8517) );
  XOR U9243 ( .A(n8499), .B(n8518), .Z(n8496) );
  NAND U9244 ( .A(A[0]), .B(B[660]), .Z(n8518) );
  NAND U9245 ( .A(B[659]), .B(A[1]), .Z(n8499) );
  NAND U9246 ( .A(n8519), .B(n8520), .Z(n789) );
  NANDN U9247 ( .A(n8521), .B(n8522), .Z(n8520) );
  OR U9248 ( .A(n8523), .B(n8524), .Z(n8522) );
  NAND U9249 ( .A(n8524), .B(n8523), .Z(n8519) );
  XOR U9250 ( .A(n791), .B(n790), .Z(\A1[657] ) );
  XOR U9251 ( .A(n8524), .B(n8525), .Z(n790) );
  XNOR U9252 ( .A(n8523), .B(n8521), .Z(n8525) );
  AND U9253 ( .A(n8526), .B(n8527), .Z(n8521) );
  NANDN U9254 ( .A(n8528), .B(n8529), .Z(n8527) );
  NANDN U9255 ( .A(n8530), .B(n8531), .Z(n8529) );
  AND U9256 ( .A(B[656]), .B(A[3]), .Z(n8523) );
  XNOR U9257 ( .A(n8513), .B(n8532), .Z(n8524) );
  XNOR U9258 ( .A(n8511), .B(n8514), .Z(n8532) );
  NAND U9259 ( .A(A[2]), .B(B[657]), .Z(n8514) );
  NANDN U9260 ( .A(n8533), .B(n8534), .Z(n8511) );
  AND U9261 ( .A(A[0]), .B(B[658]), .Z(n8534) );
  XOR U9262 ( .A(n8516), .B(n8535), .Z(n8513) );
  NAND U9263 ( .A(A[0]), .B(B[659]), .Z(n8535) );
  NAND U9264 ( .A(B[658]), .B(A[1]), .Z(n8516) );
  NAND U9265 ( .A(n8536), .B(n8537), .Z(n791) );
  NANDN U9266 ( .A(n8538), .B(n8539), .Z(n8537) );
  OR U9267 ( .A(n8540), .B(n8541), .Z(n8539) );
  NAND U9268 ( .A(n8541), .B(n8540), .Z(n8536) );
  XOR U9269 ( .A(n793), .B(n792), .Z(\A1[656] ) );
  XOR U9270 ( .A(n8541), .B(n8542), .Z(n792) );
  XNOR U9271 ( .A(n8540), .B(n8538), .Z(n8542) );
  AND U9272 ( .A(n8543), .B(n8544), .Z(n8538) );
  NANDN U9273 ( .A(n8545), .B(n8546), .Z(n8544) );
  NANDN U9274 ( .A(n8547), .B(n8548), .Z(n8546) );
  AND U9275 ( .A(B[655]), .B(A[3]), .Z(n8540) );
  XNOR U9276 ( .A(n8530), .B(n8549), .Z(n8541) );
  XNOR U9277 ( .A(n8528), .B(n8531), .Z(n8549) );
  NAND U9278 ( .A(A[2]), .B(B[656]), .Z(n8531) );
  NANDN U9279 ( .A(n8550), .B(n8551), .Z(n8528) );
  AND U9280 ( .A(A[0]), .B(B[657]), .Z(n8551) );
  XOR U9281 ( .A(n8533), .B(n8552), .Z(n8530) );
  NAND U9282 ( .A(A[0]), .B(B[658]), .Z(n8552) );
  NAND U9283 ( .A(B[657]), .B(A[1]), .Z(n8533) );
  NAND U9284 ( .A(n8553), .B(n8554), .Z(n793) );
  NANDN U9285 ( .A(n8555), .B(n8556), .Z(n8554) );
  OR U9286 ( .A(n8557), .B(n8558), .Z(n8556) );
  NAND U9287 ( .A(n8558), .B(n8557), .Z(n8553) );
  XOR U9288 ( .A(n795), .B(n794), .Z(\A1[655] ) );
  XOR U9289 ( .A(n8558), .B(n8559), .Z(n794) );
  XNOR U9290 ( .A(n8557), .B(n8555), .Z(n8559) );
  AND U9291 ( .A(n8560), .B(n8561), .Z(n8555) );
  NANDN U9292 ( .A(n8562), .B(n8563), .Z(n8561) );
  NANDN U9293 ( .A(n8564), .B(n8565), .Z(n8563) );
  AND U9294 ( .A(B[654]), .B(A[3]), .Z(n8557) );
  XNOR U9295 ( .A(n8547), .B(n8566), .Z(n8558) );
  XNOR U9296 ( .A(n8545), .B(n8548), .Z(n8566) );
  NAND U9297 ( .A(A[2]), .B(B[655]), .Z(n8548) );
  NANDN U9298 ( .A(n8567), .B(n8568), .Z(n8545) );
  AND U9299 ( .A(A[0]), .B(B[656]), .Z(n8568) );
  XOR U9300 ( .A(n8550), .B(n8569), .Z(n8547) );
  NAND U9301 ( .A(A[0]), .B(B[657]), .Z(n8569) );
  NAND U9302 ( .A(B[656]), .B(A[1]), .Z(n8550) );
  NAND U9303 ( .A(n8570), .B(n8571), .Z(n795) );
  NANDN U9304 ( .A(n8572), .B(n8573), .Z(n8571) );
  OR U9305 ( .A(n8574), .B(n8575), .Z(n8573) );
  NAND U9306 ( .A(n8575), .B(n8574), .Z(n8570) );
  XOR U9307 ( .A(n797), .B(n796), .Z(\A1[654] ) );
  XOR U9308 ( .A(n8575), .B(n8576), .Z(n796) );
  XNOR U9309 ( .A(n8574), .B(n8572), .Z(n8576) );
  AND U9310 ( .A(n8577), .B(n8578), .Z(n8572) );
  NANDN U9311 ( .A(n8579), .B(n8580), .Z(n8578) );
  NANDN U9312 ( .A(n8581), .B(n8582), .Z(n8580) );
  AND U9313 ( .A(B[653]), .B(A[3]), .Z(n8574) );
  XNOR U9314 ( .A(n8564), .B(n8583), .Z(n8575) );
  XNOR U9315 ( .A(n8562), .B(n8565), .Z(n8583) );
  NAND U9316 ( .A(A[2]), .B(B[654]), .Z(n8565) );
  NANDN U9317 ( .A(n8584), .B(n8585), .Z(n8562) );
  AND U9318 ( .A(A[0]), .B(B[655]), .Z(n8585) );
  XOR U9319 ( .A(n8567), .B(n8586), .Z(n8564) );
  NAND U9320 ( .A(A[0]), .B(B[656]), .Z(n8586) );
  NAND U9321 ( .A(B[655]), .B(A[1]), .Z(n8567) );
  NAND U9322 ( .A(n8587), .B(n8588), .Z(n797) );
  NANDN U9323 ( .A(n8589), .B(n8590), .Z(n8588) );
  OR U9324 ( .A(n8591), .B(n8592), .Z(n8590) );
  NAND U9325 ( .A(n8592), .B(n8591), .Z(n8587) );
  XOR U9326 ( .A(n799), .B(n798), .Z(\A1[653] ) );
  XOR U9327 ( .A(n8592), .B(n8593), .Z(n798) );
  XNOR U9328 ( .A(n8591), .B(n8589), .Z(n8593) );
  AND U9329 ( .A(n8594), .B(n8595), .Z(n8589) );
  NANDN U9330 ( .A(n8596), .B(n8597), .Z(n8595) );
  NANDN U9331 ( .A(n8598), .B(n8599), .Z(n8597) );
  AND U9332 ( .A(B[652]), .B(A[3]), .Z(n8591) );
  XNOR U9333 ( .A(n8581), .B(n8600), .Z(n8592) );
  XNOR U9334 ( .A(n8579), .B(n8582), .Z(n8600) );
  NAND U9335 ( .A(A[2]), .B(B[653]), .Z(n8582) );
  NANDN U9336 ( .A(n8601), .B(n8602), .Z(n8579) );
  AND U9337 ( .A(A[0]), .B(B[654]), .Z(n8602) );
  XOR U9338 ( .A(n8584), .B(n8603), .Z(n8581) );
  NAND U9339 ( .A(A[0]), .B(B[655]), .Z(n8603) );
  NAND U9340 ( .A(B[654]), .B(A[1]), .Z(n8584) );
  NAND U9341 ( .A(n8604), .B(n8605), .Z(n799) );
  NANDN U9342 ( .A(n8606), .B(n8607), .Z(n8605) );
  OR U9343 ( .A(n8608), .B(n8609), .Z(n8607) );
  NAND U9344 ( .A(n8609), .B(n8608), .Z(n8604) );
  XOR U9345 ( .A(n801), .B(n800), .Z(\A1[652] ) );
  XOR U9346 ( .A(n8609), .B(n8610), .Z(n800) );
  XNOR U9347 ( .A(n8608), .B(n8606), .Z(n8610) );
  AND U9348 ( .A(n8611), .B(n8612), .Z(n8606) );
  NANDN U9349 ( .A(n8613), .B(n8614), .Z(n8612) );
  NANDN U9350 ( .A(n8615), .B(n8616), .Z(n8614) );
  AND U9351 ( .A(B[651]), .B(A[3]), .Z(n8608) );
  XNOR U9352 ( .A(n8598), .B(n8617), .Z(n8609) );
  XNOR U9353 ( .A(n8596), .B(n8599), .Z(n8617) );
  NAND U9354 ( .A(A[2]), .B(B[652]), .Z(n8599) );
  NANDN U9355 ( .A(n8618), .B(n8619), .Z(n8596) );
  AND U9356 ( .A(A[0]), .B(B[653]), .Z(n8619) );
  XOR U9357 ( .A(n8601), .B(n8620), .Z(n8598) );
  NAND U9358 ( .A(A[0]), .B(B[654]), .Z(n8620) );
  NAND U9359 ( .A(B[653]), .B(A[1]), .Z(n8601) );
  NAND U9360 ( .A(n8621), .B(n8622), .Z(n801) );
  NANDN U9361 ( .A(n8623), .B(n8624), .Z(n8622) );
  OR U9362 ( .A(n8625), .B(n8626), .Z(n8624) );
  NAND U9363 ( .A(n8626), .B(n8625), .Z(n8621) );
  XOR U9364 ( .A(n803), .B(n802), .Z(\A1[651] ) );
  XOR U9365 ( .A(n8626), .B(n8627), .Z(n802) );
  XNOR U9366 ( .A(n8625), .B(n8623), .Z(n8627) );
  AND U9367 ( .A(n8628), .B(n8629), .Z(n8623) );
  NANDN U9368 ( .A(n8630), .B(n8631), .Z(n8629) );
  NANDN U9369 ( .A(n8632), .B(n8633), .Z(n8631) );
  AND U9370 ( .A(B[650]), .B(A[3]), .Z(n8625) );
  XNOR U9371 ( .A(n8615), .B(n8634), .Z(n8626) );
  XNOR U9372 ( .A(n8613), .B(n8616), .Z(n8634) );
  NAND U9373 ( .A(A[2]), .B(B[651]), .Z(n8616) );
  NANDN U9374 ( .A(n8635), .B(n8636), .Z(n8613) );
  AND U9375 ( .A(A[0]), .B(B[652]), .Z(n8636) );
  XOR U9376 ( .A(n8618), .B(n8637), .Z(n8615) );
  NAND U9377 ( .A(A[0]), .B(B[653]), .Z(n8637) );
  NAND U9378 ( .A(B[652]), .B(A[1]), .Z(n8618) );
  NAND U9379 ( .A(n8638), .B(n8639), .Z(n803) );
  NANDN U9380 ( .A(n8640), .B(n8641), .Z(n8639) );
  OR U9381 ( .A(n8642), .B(n8643), .Z(n8641) );
  NAND U9382 ( .A(n8643), .B(n8642), .Z(n8638) );
  XOR U9383 ( .A(n805), .B(n804), .Z(\A1[650] ) );
  XOR U9384 ( .A(n8643), .B(n8644), .Z(n804) );
  XNOR U9385 ( .A(n8642), .B(n8640), .Z(n8644) );
  AND U9386 ( .A(n8645), .B(n8646), .Z(n8640) );
  NANDN U9387 ( .A(n8647), .B(n8648), .Z(n8646) );
  NANDN U9388 ( .A(n8649), .B(n8650), .Z(n8648) );
  AND U9389 ( .A(B[649]), .B(A[3]), .Z(n8642) );
  XNOR U9390 ( .A(n8632), .B(n8651), .Z(n8643) );
  XNOR U9391 ( .A(n8630), .B(n8633), .Z(n8651) );
  NAND U9392 ( .A(A[2]), .B(B[650]), .Z(n8633) );
  NANDN U9393 ( .A(n8652), .B(n8653), .Z(n8630) );
  AND U9394 ( .A(A[0]), .B(B[651]), .Z(n8653) );
  XOR U9395 ( .A(n8635), .B(n8654), .Z(n8632) );
  NAND U9396 ( .A(A[0]), .B(B[652]), .Z(n8654) );
  NAND U9397 ( .A(B[651]), .B(A[1]), .Z(n8635) );
  NAND U9398 ( .A(n8655), .B(n8656), .Z(n805) );
  NANDN U9399 ( .A(n8657), .B(n8658), .Z(n8656) );
  OR U9400 ( .A(n8659), .B(n8660), .Z(n8658) );
  NAND U9401 ( .A(n8660), .B(n8659), .Z(n8655) );
  XOR U9402 ( .A(n787), .B(n786), .Z(\A1[64] ) );
  XOR U9403 ( .A(n8490), .B(n8661), .Z(n786) );
  XNOR U9404 ( .A(n8489), .B(n8487), .Z(n8661) );
  AND U9405 ( .A(n8662), .B(n8663), .Z(n8487) );
  NANDN U9406 ( .A(n8664), .B(n8665), .Z(n8663) );
  NANDN U9407 ( .A(n8666), .B(n8667), .Z(n8665) );
  AND U9408 ( .A(B[63]), .B(A[3]), .Z(n8489) );
  XNOR U9409 ( .A(n8479), .B(n8668), .Z(n8490) );
  XNOR U9410 ( .A(n8477), .B(n8480), .Z(n8668) );
  NAND U9411 ( .A(A[2]), .B(B[64]), .Z(n8480) );
  NANDN U9412 ( .A(n8669), .B(n8670), .Z(n8477) );
  AND U9413 ( .A(A[0]), .B(B[65]), .Z(n8670) );
  XOR U9414 ( .A(n8482), .B(n8671), .Z(n8479) );
  NAND U9415 ( .A(A[0]), .B(B[66]), .Z(n8671) );
  NAND U9416 ( .A(B[65]), .B(A[1]), .Z(n8482) );
  NAND U9417 ( .A(n8672), .B(n8673), .Z(n787) );
  NANDN U9418 ( .A(n8674), .B(n8675), .Z(n8673) );
  OR U9419 ( .A(n8676), .B(n8677), .Z(n8675) );
  NAND U9420 ( .A(n8677), .B(n8676), .Z(n8672) );
  XOR U9421 ( .A(n807), .B(n806), .Z(\A1[649] ) );
  XOR U9422 ( .A(n8660), .B(n8678), .Z(n806) );
  XNOR U9423 ( .A(n8659), .B(n8657), .Z(n8678) );
  AND U9424 ( .A(n8679), .B(n8680), .Z(n8657) );
  NANDN U9425 ( .A(n8681), .B(n8682), .Z(n8680) );
  NANDN U9426 ( .A(n8683), .B(n8684), .Z(n8682) );
  AND U9427 ( .A(B[648]), .B(A[3]), .Z(n8659) );
  XNOR U9428 ( .A(n8649), .B(n8685), .Z(n8660) );
  XNOR U9429 ( .A(n8647), .B(n8650), .Z(n8685) );
  NAND U9430 ( .A(A[2]), .B(B[649]), .Z(n8650) );
  NANDN U9431 ( .A(n8686), .B(n8687), .Z(n8647) );
  AND U9432 ( .A(A[0]), .B(B[650]), .Z(n8687) );
  XOR U9433 ( .A(n8652), .B(n8688), .Z(n8649) );
  NAND U9434 ( .A(A[0]), .B(B[651]), .Z(n8688) );
  NAND U9435 ( .A(B[650]), .B(A[1]), .Z(n8652) );
  NAND U9436 ( .A(n8689), .B(n8690), .Z(n807) );
  NANDN U9437 ( .A(n8691), .B(n8692), .Z(n8690) );
  OR U9438 ( .A(n8693), .B(n8694), .Z(n8692) );
  NAND U9439 ( .A(n8694), .B(n8693), .Z(n8689) );
  XOR U9440 ( .A(n811), .B(n810), .Z(\A1[648] ) );
  XOR U9441 ( .A(n8694), .B(n8695), .Z(n810) );
  XNOR U9442 ( .A(n8693), .B(n8691), .Z(n8695) );
  AND U9443 ( .A(n8696), .B(n8697), .Z(n8691) );
  NANDN U9444 ( .A(n8698), .B(n8699), .Z(n8697) );
  NANDN U9445 ( .A(n8700), .B(n8701), .Z(n8699) );
  AND U9446 ( .A(B[647]), .B(A[3]), .Z(n8693) );
  XNOR U9447 ( .A(n8683), .B(n8702), .Z(n8694) );
  XNOR U9448 ( .A(n8681), .B(n8684), .Z(n8702) );
  NAND U9449 ( .A(A[2]), .B(B[648]), .Z(n8684) );
  NANDN U9450 ( .A(n8703), .B(n8704), .Z(n8681) );
  AND U9451 ( .A(A[0]), .B(B[649]), .Z(n8704) );
  XOR U9452 ( .A(n8686), .B(n8705), .Z(n8683) );
  NAND U9453 ( .A(A[0]), .B(B[650]), .Z(n8705) );
  NAND U9454 ( .A(B[649]), .B(A[1]), .Z(n8686) );
  NAND U9455 ( .A(n8706), .B(n8707), .Z(n811) );
  NANDN U9456 ( .A(n8708), .B(n8709), .Z(n8707) );
  OR U9457 ( .A(n8710), .B(n8711), .Z(n8709) );
  NAND U9458 ( .A(n8711), .B(n8710), .Z(n8706) );
  XOR U9459 ( .A(n813), .B(n812), .Z(\A1[647] ) );
  XOR U9460 ( .A(n8711), .B(n8712), .Z(n812) );
  XNOR U9461 ( .A(n8710), .B(n8708), .Z(n8712) );
  AND U9462 ( .A(n8713), .B(n8714), .Z(n8708) );
  NANDN U9463 ( .A(n8715), .B(n8716), .Z(n8714) );
  NANDN U9464 ( .A(n8717), .B(n8718), .Z(n8716) );
  AND U9465 ( .A(B[646]), .B(A[3]), .Z(n8710) );
  XNOR U9466 ( .A(n8700), .B(n8719), .Z(n8711) );
  XNOR U9467 ( .A(n8698), .B(n8701), .Z(n8719) );
  NAND U9468 ( .A(A[2]), .B(B[647]), .Z(n8701) );
  NANDN U9469 ( .A(n8720), .B(n8721), .Z(n8698) );
  AND U9470 ( .A(A[0]), .B(B[648]), .Z(n8721) );
  XOR U9471 ( .A(n8703), .B(n8722), .Z(n8700) );
  NAND U9472 ( .A(A[0]), .B(B[649]), .Z(n8722) );
  NAND U9473 ( .A(B[648]), .B(A[1]), .Z(n8703) );
  NAND U9474 ( .A(n8723), .B(n8724), .Z(n813) );
  NANDN U9475 ( .A(n8725), .B(n8726), .Z(n8724) );
  OR U9476 ( .A(n8727), .B(n8728), .Z(n8726) );
  NAND U9477 ( .A(n8728), .B(n8727), .Z(n8723) );
  XOR U9478 ( .A(n815), .B(n814), .Z(\A1[646] ) );
  XOR U9479 ( .A(n8728), .B(n8729), .Z(n814) );
  XNOR U9480 ( .A(n8727), .B(n8725), .Z(n8729) );
  AND U9481 ( .A(n8730), .B(n8731), .Z(n8725) );
  NANDN U9482 ( .A(n8732), .B(n8733), .Z(n8731) );
  NANDN U9483 ( .A(n8734), .B(n8735), .Z(n8733) );
  AND U9484 ( .A(B[645]), .B(A[3]), .Z(n8727) );
  XNOR U9485 ( .A(n8717), .B(n8736), .Z(n8728) );
  XNOR U9486 ( .A(n8715), .B(n8718), .Z(n8736) );
  NAND U9487 ( .A(A[2]), .B(B[646]), .Z(n8718) );
  NANDN U9488 ( .A(n8737), .B(n8738), .Z(n8715) );
  AND U9489 ( .A(A[0]), .B(B[647]), .Z(n8738) );
  XOR U9490 ( .A(n8720), .B(n8739), .Z(n8717) );
  NAND U9491 ( .A(A[0]), .B(B[648]), .Z(n8739) );
  NAND U9492 ( .A(B[647]), .B(A[1]), .Z(n8720) );
  NAND U9493 ( .A(n8740), .B(n8741), .Z(n815) );
  NANDN U9494 ( .A(n8742), .B(n8743), .Z(n8741) );
  OR U9495 ( .A(n8744), .B(n8745), .Z(n8743) );
  NAND U9496 ( .A(n8745), .B(n8744), .Z(n8740) );
  XOR U9497 ( .A(n817), .B(n816), .Z(\A1[645] ) );
  XOR U9498 ( .A(n8745), .B(n8746), .Z(n816) );
  XNOR U9499 ( .A(n8744), .B(n8742), .Z(n8746) );
  AND U9500 ( .A(n8747), .B(n8748), .Z(n8742) );
  NANDN U9501 ( .A(n8749), .B(n8750), .Z(n8748) );
  NANDN U9502 ( .A(n8751), .B(n8752), .Z(n8750) );
  AND U9503 ( .A(B[644]), .B(A[3]), .Z(n8744) );
  XNOR U9504 ( .A(n8734), .B(n8753), .Z(n8745) );
  XNOR U9505 ( .A(n8732), .B(n8735), .Z(n8753) );
  NAND U9506 ( .A(A[2]), .B(B[645]), .Z(n8735) );
  NANDN U9507 ( .A(n8754), .B(n8755), .Z(n8732) );
  AND U9508 ( .A(A[0]), .B(B[646]), .Z(n8755) );
  XOR U9509 ( .A(n8737), .B(n8756), .Z(n8734) );
  NAND U9510 ( .A(A[0]), .B(B[647]), .Z(n8756) );
  NAND U9511 ( .A(B[646]), .B(A[1]), .Z(n8737) );
  NAND U9512 ( .A(n8757), .B(n8758), .Z(n817) );
  NANDN U9513 ( .A(n8759), .B(n8760), .Z(n8758) );
  OR U9514 ( .A(n8761), .B(n8762), .Z(n8760) );
  NAND U9515 ( .A(n8762), .B(n8761), .Z(n8757) );
  XOR U9516 ( .A(n819), .B(n818), .Z(\A1[644] ) );
  XOR U9517 ( .A(n8762), .B(n8763), .Z(n818) );
  XNOR U9518 ( .A(n8761), .B(n8759), .Z(n8763) );
  AND U9519 ( .A(n8764), .B(n8765), .Z(n8759) );
  NANDN U9520 ( .A(n8766), .B(n8767), .Z(n8765) );
  NANDN U9521 ( .A(n8768), .B(n8769), .Z(n8767) );
  AND U9522 ( .A(B[643]), .B(A[3]), .Z(n8761) );
  XNOR U9523 ( .A(n8751), .B(n8770), .Z(n8762) );
  XNOR U9524 ( .A(n8749), .B(n8752), .Z(n8770) );
  NAND U9525 ( .A(A[2]), .B(B[644]), .Z(n8752) );
  NANDN U9526 ( .A(n8771), .B(n8772), .Z(n8749) );
  AND U9527 ( .A(A[0]), .B(B[645]), .Z(n8772) );
  XOR U9528 ( .A(n8754), .B(n8773), .Z(n8751) );
  NAND U9529 ( .A(A[0]), .B(B[646]), .Z(n8773) );
  NAND U9530 ( .A(B[645]), .B(A[1]), .Z(n8754) );
  NAND U9531 ( .A(n8774), .B(n8775), .Z(n819) );
  NANDN U9532 ( .A(n8776), .B(n8777), .Z(n8775) );
  OR U9533 ( .A(n8778), .B(n8779), .Z(n8777) );
  NAND U9534 ( .A(n8779), .B(n8778), .Z(n8774) );
  XOR U9535 ( .A(n821), .B(n820), .Z(\A1[643] ) );
  XOR U9536 ( .A(n8779), .B(n8780), .Z(n820) );
  XNOR U9537 ( .A(n8778), .B(n8776), .Z(n8780) );
  AND U9538 ( .A(n8781), .B(n8782), .Z(n8776) );
  NANDN U9539 ( .A(n8783), .B(n8784), .Z(n8782) );
  NANDN U9540 ( .A(n8785), .B(n8786), .Z(n8784) );
  AND U9541 ( .A(B[642]), .B(A[3]), .Z(n8778) );
  XNOR U9542 ( .A(n8768), .B(n8787), .Z(n8779) );
  XNOR U9543 ( .A(n8766), .B(n8769), .Z(n8787) );
  NAND U9544 ( .A(A[2]), .B(B[643]), .Z(n8769) );
  NANDN U9545 ( .A(n8788), .B(n8789), .Z(n8766) );
  AND U9546 ( .A(A[0]), .B(B[644]), .Z(n8789) );
  XOR U9547 ( .A(n8771), .B(n8790), .Z(n8768) );
  NAND U9548 ( .A(A[0]), .B(B[645]), .Z(n8790) );
  NAND U9549 ( .A(B[644]), .B(A[1]), .Z(n8771) );
  NAND U9550 ( .A(n8791), .B(n8792), .Z(n821) );
  NANDN U9551 ( .A(n8793), .B(n8794), .Z(n8792) );
  OR U9552 ( .A(n8795), .B(n8796), .Z(n8794) );
  NAND U9553 ( .A(n8796), .B(n8795), .Z(n8791) );
  XOR U9554 ( .A(n823), .B(n822), .Z(\A1[642] ) );
  XOR U9555 ( .A(n8796), .B(n8797), .Z(n822) );
  XNOR U9556 ( .A(n8795), .B(n8793), .Z(n8797) );
  AND U9557 ( .A(n8798), .B(n8799), .Z(n8793) );
  NANDN U9558 ( .A(n8800), .B(n8801), .Z(n8799) );
  NANDN U9559 ( .A(n8802), .B(n8803), .Z(n8801) );
  AND U9560 ( .A(B[641]), .B(A[3]), .Z(n8795) );
  XNOR U9561 ( .A(n8785), .B(n8804), .Z(n8796) );
  XNOR U9562 ( .A(n8783), .B(n8786), .Z(n8804) );
  NAND U9563 ( .A(A[2]), .B(B[642]), .Z(n8786) );
  NANDN U9564 ( .A(n8805), .B(n8806), .Z(n8783) );
  AND U9565 ( .A(A[0]), .B(B[643]), .Z(n8806) );
  XOR U9566 ( .A(n8788), .B(n8807), .Z(n8785) );
  NAND U9567 ( .A(A[0]), .B(B[644]), .Z(n8807) );
  NAND U9568 ( .A(B[643]), .B(A[1]), .Z(n8788) );
  NAND U9569 ( .A(n8808), .B(n8809), .Z(n823) );
  NANDN U9570 ( .A(n8810), .B(n8811), .Z(n8809) );
  OR U9571 ( .A(n8812), .B(n8813), .Z(n8811) );
  NAND U9572 ( .A(n8813), .B(n8812), .Z(n8808) );
  XOR U9573 ( .A(n825), .B(n824), .Z(\A1[641] ) );
  XOR U9574 ( .A(n8813), .B(n8814), .Z(n824) );
  XNOR U9575 ( .A(n8812), .B(n8810), .Z(n8814) );
  AND U9576 ( .A(n8815), .B(n8816), .Z(n8810) );
  NANDN U9577 ( .A(n8817), .B(n8818), .Z(n8816) );
  NANDN U9578 ( .A(n8819), .B(n8820), .Z(n8818) );
  AND U9579 ( .A(B[640]), .B(A[3]), .Z(n8812) );
  XNOR U9580 ( .A(n8802), .B(n8821), .Z(n8813) );
  XNOR U9581 ( .A(n8800), .B(n8803), .Z(n8821) );
  NAND U9582 ( .A(A[2]), .B(B[641]), .Z(n8803) );
  NANDN U9583 ( .A(n8822), .B(n8823), .Z(n8800) );
  AND U9584 ( .A(A[0]), .B(B[642]), .Z(n8823) );
  XOR U9585 ( .A(n8805), .B(n8824), .Z(n8802) );
  NAND U9586 ( .A(A[0]), .B(B[643]), .Z(n8824) );
  NAND U9587 ( .A(B[642]), .B(A[1]), .Z(n8805) );
  NAND U9588 ( .A(n8825), .B(n8826), .Z(n825) );
  NANDN U9589 ( .A(n8827), .B(n8828), .Z(n8826) );
  OR U9590 ( .A(n8829), .B(n8830), .Z(n8828) );
  NAND U9591 ( .A(n8830), .B(n8829), .Z(n8825) );
  XOR U9592 ( .A(n827), .B(n826), .Z(\A1[640] ) );
  XOR U9593 ( .A(n8830), .B(n8831), .Z(n826) );
  XNOR U9594 ( .A(n8829), .B(n8827), .Z(n8831) );
  AND U9595 ( .A(n8832), .B(n8833), .Z(n8827) );
  NANDN U9596 ( .A(n8834), .B(n8835), .Z(n8833) );
  NANDN U9597 ( .A(n8836), .B(n8837), .Z(n8835) );
  AND U9598 ( .A(B[639]), .B(A[3]), .Z(n8829) );
  XNOR U9599 ( .A(n8819), .B(n8838), .Z(n8830) );
  XNOR U9600 ( .A(n8817), .B(n8820), .Z(n8838) );
  NAND U9601 ( .A(A[2]), .B(B[640]), .Z(n8820) );
  NANDN U9602 ( .A(n8839), .B(n8840), .Z(n8817) );
  AND U9603 ( .A(A[0]), .B(B[641]), .Z(n8840) );
  XOR U9604 ( .A(n8822), .B(n8841), .Z(n8819) );
  NAND U9605 ( .A(A[0]), .B(B[642]), .Z(n8841) );
  NAND U9606 ( .A(B[641]), .B(A[1]), .Z(n8822) );
  NAND U9607 ( .A(n8842), .B(n8843), .Z(n827) );
  NANDN U9608 ( .A(n8844), .B(n8845), .Z(n8843) );
  OR U9609 ( .A(n8846), .B(n8847), .Z(n8845) );
  NAND U9610 ( .A(n8847), .B(n8846), .Z(n8842) );
  XOR U9611 ( .A(n809), .B(n808), .Z(\A1[63] ) );
  XOR U9612 ( .A(n8677), .B(n8848), .Z(n808) );
  XNOR U9613 ( .A(n8676), .B(n8674), .Z(n8848) );
  AND U9614 ( .A(n8849), .B(n8850), .Z(n8674) );
  NANDN U9615 ( .A(n8851), .B(n8852), .Z(n8850) );
  NANDN U9616 ( .A(n8853), .B(n8854), .Z(n8852) );
  AND U9617 ( .A(B[62]), .B(A[3]), .Z(n8676) );
  XNOR U9618 ( .A(n8666), .B(n8855), .Z(n8677) );
  XNOR U9619 ( .A(n8664), .B(n8667), .Z(n8855) );
  NAND U9620 ( .A(A[2]), .B(B[63]), .Z(n8667) );
  NANDN U9621 ( .A(n8856), .B(n8857), .Z(n8664) );
  AND U9622 ( .A(A[0]), .B(B[64]), .Z(n8857) );
  XOR U9623 ( .A(n8669), .B(n8858), .Z(n8666) );
  NAND U9624 ( .A(A[0]), .B(B[65]), .Z(n8858) );
  NAND U9625 ( .A(B[64]), .B(A[1]), .Z(n8669) );
  NAND U9626 ( .A(n8859), .B(n8860), .Z(n809) );
  NANDN U9627 ( .A(n8861), .B(n8862), .Z(n8860) );
  OR U9628 ( .A(n8863), .B(n8864), .Z(n8862) );
  NAND U9629 ( .A(n8864), .B(n8863), .Z(n8859) );
  XOR U9630 ( .A(n829), .B(n828), .Z(\A1[639] ) );
  XOR U9631 ( .A(n8847), .B(n8865), .Z(n828) );
  XNOR U9632 ( .A(n8846), .B(n8844), .Z(n8865) );
  AND U9633 ( .A(n8866), .B(n8867), .Z(n8844) );
  NANDN U9634 ( .A(n8868), .B(n8869), .Z(n8867) );
  NANDN U9635 ( .A(n8870), .B(n8871), .Z(n8869) );
  AND U9636 ( .A(B[638]), .B(A[3]), .Z(n8846) );
  XNOR U9637 ( .A(n8836), .B(n8872), .Z(n8847) );
  XNOR U9638 ( .A(n8834), .B(n8837), .Z(n8872) );
  NAND U9639 ( .A(A[2]), .B(B[639]), .Z(n8837) );
  NANDN U9640 ( .A(n8873), .B(n8874), .Z(n8834) );
  AND U9641 ( .A(A[0]), .B(B[640]), .Z(n8874) );
  XOR U9642 ( .A(n8839), .B(n8875), .Z(n8836) );
  NAND U9643 ( .A(A[0]), .B(B[641]), .Z(n8875) );
  NAND U9644 ( .A(B[640]), .B(A[1]), .Z(n8839) );
  NAND U9645 ( .A(n8876), .B(n8877), .Z(n829) );
  NANDN U9646 ( .A(n8878), .B(n8879), .Z(n8877) );
  OR U9647 ( .A(n8880), .B(n8881), .Z(n8879) );
  NAND U9648 ( .A(n8881), .B(n8880), .Z(n8876) );
  XOR U9649 ( .A(n833), .B(n832), .Z(\A1[638] ) );
  XOR U9650 ( .A(n8881), .B(n8882), .Z(n832) );
  XNOR U9651 ( .A(n8880), .B(n8878), .Z(n8882) );
  AND U9652 ( .A(n8883), .B(n8884), .Z(n8878) );
  NANDN U9653 ( .A(n8885), .B(n8886), .Z(n8884) );
  NANDN U9654 ( .A(n8887), .B(n8888), .Z(n8886) );
  AND U9655 ( .A(B[637]), .B(A[3]), .Z(n8880) );
  XNOR U9656 ( .A(n8870), .B(n8889), .Z(n8881) );
  XNOR U9657 ( .A(n8868), .B(n8871), .Z(n8889) );
  NAND U9658 ( .A(A[2]), .B(B[638]), .Z(n8871) );
  NANDN U9659 ( .A(n8890), .B(n8891), .Z(n8868) );
  AND U9660 ( .A(A[0]), .B(B[639]), .Z(n8891) );
  XOR U9661 ( .A(n8873), .B(n8892), .Z(n8870) );
  NAND U9662 ( .A(A[0]), .B(B[640]), .Z(n8892) );
  NAND U9663 ( .A(B[639]), .B(A[1]), .Z(n8873) );
  NAND U9664 ( .A(n8893), .B(n8894), .Z(n833) );
  NANDN U9665 ( .A(n8895), .B(n8896), .Z(n8894) );
  OR U9666 ( .A(n8897), .B(n8898), .Z(n8896) );
  NAND U9667 ( .A(n8898), .B(n8897), .Z(n8893) );
  XOR U9668 ( .A(n835), .B(n834), .Z(\A1[637] ) );
  XOR U9669 ( .A(n8898), .B(n8899), .Z(n834) );
  XNOR U9670 ( .A(n8897), .B(n8895), .Z(n8899) );
  AND U9671 ( .A(n8900), .B(n8901), .Z(n8895) );
  NANDN U9672 ( .A(n8902), .B(n8903), .Z(n8901) );
  NANDN U9673 ( .A(n8904), .B(n8905), .Z(n8903) );
  AND U9674 ( .A(B[636]), .B(A[3]), .Z(n8897) );
  XNOR U9675 ( .A(n8887), .B(n8906), .Z(n8898) );
  XNOR U9676 ( .A(n8885), .B(n8888), .Z(n8906) );
  NAND U9677 ( .A(A[2]), .B(B[637]), .Z(n8888) );
  NANDN U9678 ( .A(n8907), .B(n8908), .Z(n8885) );
  AND U9679 ( .A(A[0]), .B(B[638]), .Z(n8908) );
  XOR U9680 ( .A(n8890), .B(n8909), .Z(n8887) );
  NAND U9681 ( .A(A[0]), .B(B[639]), .Z(n8909) );
  NAND U9682 ( .A(B[638]), .B(A[1]), .Z(n8890) );
  NAND U9683 ( .A(n8910), .B(n8911), .Z(n835) );
  NANDN U9684 ( .A(n8912), .B(n8913), .Z(n8911) );
  OR U9685 ( .A(n8914), .B(n8915), .Z(n8913) );
  NAND U9686 ( .A(n8915), .B(n8914), .Z(n8910) );
  XOR U9687 ( .A(n837), .B(n836), .Z(\A1[636] ) );
  XOR U9688 ( .A(n8915), .B(n8916), .Z(n836) );
  XNOR U9689 ( .A(n8914), .B(n8912), .Z(n8916) );
  AND U9690 ( .A(n8917), .B(n8918), .Z(n8912) );
  NANDN U9691 ( .A(n8919), .B(n8920), .Z(n8918) );
  NANDN U9692 ( .A(n8921), .B(n8922), .Z(n8920) );
  AND U9693 ( .A(B[635]), .B(A[3]), .Z(n8914) );
  XNOR U9694 ( .A(n8904), .B(n8923), .Z(n8915) );
  XNOR U9695 ( .A(n8902), .B(n8905), .Z(n8923) );
  NAND U9696 ( .A(A[2]), .B(B[636]), .Z(n8905) );
  NANDN U9697 ( .A(n8924), .B(n8925), .Z(n8902) );
  AND U9698 ( .A(A[0]), .B(B[637]), .Z(n8925) );
  XOR U9699 ( .A(n8907), .B(n8926), .Z(n8904) );
  NAND U9700 ( .A(A[0]), .B(B[638]), .Z(n8926) );
  NAND U9701 ( .A(B[637]), .B(A[1]), .Z(n8907) );
  NAND U9702 ( .A(n8927), .B(n8928), .Z(n837) );
  NANDN U9703 ( .A(n8929), .B(n8930), .Z(n8928) );
  OR U9704 ( .A(n8931), .B(n8932), .Z(n8930) );
  NAND U9705 ( .A(n8932), .B(n8931), .Z(n8927) );
  XOR U9706 ( .A(n839), .B(n838), .Z(\A1[635] ) );
  XOR U9707 ( .A(n8932), .B(n8933), .Z(n838) );
  XNOR U9708 ( .A(n8931), .B(n8929), .Z(n8933) );
  AND U9709 ( .A(n8934), .B(n8935), .Z(n8929) );
  NANDN U9710 ( .A(n8936), .B(n8937), .Z(n8935) );
  NANDN U9711 ( .A(n8938), .B(n8939), .Z(n8937) );
  AND U9712 ( .A(B[634]), .B(A[3]), .Z(n8931) );
  XNOR U9713 ( .A(n8921), .B(n8940), .Z(n8932) );
  XNOR U9714 ( .A(n8919), .B(n8922), .Z(n8940) );
  NAND U9715 ( .A(A[2]), .B(B[635]), .Z(n8922) );
  NANDN U9716 ( .A(n8941), .B(n8942), .Z(n8919) );
  AND U9717 ( .A(A[0]), .B(B[636]), .Z(n8942) );
  XOR U9718 ( .A(n8924), .B(n8943), .Z(n8921) );
  NAND U9719 ( .A(A[0]), .B(B[637]), .Z(n8943) );
  NAND U9720 ( .A(B[636]), .B(A[1]), .Z(n8924) );
  NAND U9721 ( .A(n8944), .B(n8945), .Z(n839) );
  NANDN U9722 ( .A(n8946), .B(n8947), .Z(n8945) );
  OR U9723 ( .A(n8948), .B(n8949), .Z(n8947) );
  NAND U9724 ( .A(n8949), .B(n8948), .Z(n8944) );
  XOR U9725 ( .A(n841), .B(n840), .Z(\A1[634] ) );
  XOR U9726 ( .A(n8949), .B(n8950), .Z(n840) );
  XNOR U9727 ( .A(n8948), .B(n8946), .Z(n8950) );
  AND U9728 ( .A(n8951), .B(n8952), .Z(n8946) );
  NANDN U9729 ( .A(n8953), .B(n8954), .Z(n8952) );
  NANDN U9730 ( .A(n8955), .B(n8956), .Z(n8954) );
  AND U9731 ( .A(B[633]), .B(A[3]), .Z(n8948) );
  XNOR U9732 ( .A(n8938), .B(n8957), .Z(n8949) );
  XNOR U9733 ( .A(n8936), .B(n8939), .Z(n8957) );
  NAND U9734 ( .A(A[2]), .B(B[634]), .Z(n8939) );
  NANDN U9735 ( .A(n8958), .B(n8959), .Z(n8936) );
  AND U9736 ( .A(A[0]), .B(B[635]), .Z(n8959) );
  XOR U9737 ( .A(n8941), .B(n8960), .Z(n8938) );
  NAND U9738 ( .A(A[0]), .B(B[636]), .Z(n8960) );
  NAND U9739 ( .A(B[635]), .B(A[1]), .Z(n8941) );
  NAND U9740 ( .A(n8961), .B(n8962), .Z(n841) );
  NANDN U9741 ( .A(n8963), .B(n8964), .Z(n8962) );
  OR U9742 ( .A(n8965), .B(n8966), .Z(n8964) );
  NAND U9743 ( .A(n8966), .B(n8965), .Z(n8961) );
  XOR U9744 ( .A(n843), .B(n842), .Z(\A1[633] ) );
  XOR U9745 ( .A(n8966), .B(n8967), .Z(n842) );
  XNOR U9746 ( .A(n8965), .B(n8963), .Z(n8967) );
  AND U9747 ( .A(n8968), .B(n8969), .Z(n8963) );
  NANDN U9748 ( .A(n8970), .B(n8971), .Z(n8969) );
  NANDN U9749 ( .A(n8972), .B(n8973), .Z(n8971) );
  AND U9750 ( .A(B[632]), .B(A[3]), .Z(n8965) );
  XNOR U9751 ( .A(n8955), .B(n8974), .Z(n8966) );
  XNOR U9752 ( .A(n8953), .B(n8956), .Z(n8974) );
  NAND U9753 ( .A(A[2]), .B(B[633]), .Z(n8956) );
  NANDN U9754 ( .A(n8975), .B(n8976), .Z(n8953) );
  AND U9755 ( .A(A[0]), .B(B[634]), .Z(n8976) );
  XOR U9756 ( .A(n8958), .B(n8977), .Z(n8955) );
  NAND U9757 ( .A(A[0]), .B(B[635]), .Z(n8977) );
  NAND U9758 ( .A(B[634]), .B(A[1]), .Z(n8958) );
  NAND U9759 ( .A(n8978), .B(n8979), .Z(n843) );
  NANDN U9760 ( .A(n8980), .B(n8981), .Z(n8979) );
  OR U9761 ( .A(n8982), .B(n8983), .Z(n8981) );
  NAND U9762 ( .A(n8983), .B(n8982), .Z(n8978) );
  XOR U9763 ( .A(n845), .B(n844), .Z(\A1[632] ) );
  XOR U9764 ( .A(n8983), .B(n8984), .Z(n844) );
  XNOR U9765 ( .A(n8982), .B(n8980), .Z(n8984) );
  AND U9766 ( .A(n8985), .B(n8986), .Z(n8980) );
  NANDN U9767 ( .A(n8987), .B(n8988), .Z(n8986) );
  NANDN U9768 ( .A(n8989), .B(n8990), .Z(n8988) );
  AND U9769 ( .A(B[631]), .B(A[3]), .Z(n8982) );
  XNOR U9770 ( .A(n8972), .B(n8991), .Z(n8983) );
  XNOR U9771 ( .A(n8970), .B(n8973), .Z(n8991) );
  NAND U9772 ( .A(A[2]), .B(B[632]), .Z(n8973) );
  NANDN U9773 ( .A(n8992), .B(n8993), .Z(n8970) );
  AND U9774 ( .A(A[0]), .B(B[633]), .Z(n8993) );
  XOR U9775 ( .A(n8975), .B(n8994), .Z(n8972) );
  NAND U9776 ( .A(A[0]), .B(B[634]), .Z(n8994) );
  NAND U9777 ( .A(B[633]), .B(A[1]), .Z(n8975) );
  NAND U9778 ( .A(n8995), .B(n8996), .Z(n845) );
  NANDN U9779 ( .A(n8997), .B(n8998), .Z(n8996) );
  OR U9780 ( .A(n8999), .B(n9000), .Z(n8998) );
  NAND U9781 ( .A(n9000), .B(n8999), .Z(n8995) );
  XOR U9782 ( .A(n847), .B(n846), .Z(\A1[631] ) );
  XOR U9783 ( .A(n9000), .B(n9001), .Z(n846) );
  XNOR U9784 ( .A(n8999), .B(n8997), .Z(n9001) );
  AND U9785 ( .A(n9002), .B(n9003), .Z(n8997) );
  NANDN U9786 ( .A(n9004), .B(n9005), .Z(n9003) );
  NANDN U9787 ( .A(n9006), .B(n9007), .Z(n9005) );
  AND U9788 ( .A(B[630]), .B(A[3]), .Z(n8999) );
  XNOR U9789 ( .A(n8989), .B(n9008), .Z(n9000) );
  XNOR U9790 ( .A(n8987), .B(n8990), .Z(n9008) );
  NAND U9791 ( .A(A[2]), .B(B[631]), .Z(n8990) );
  NANDN U9792 ( .A(n9009), .B(n9010), .Z(n8987) );
  AND U9793 ( .A(A[0]), .B(B[632]), .Z(n9010) );
  XOR U9794 ( .A(n8992), .B(n9011), .Z(n8989) );
  NAND U9795 ( .A(A[0]), .B(B[633]), .Z(n9011) );
  NAND U9796 ( .A(B[632]), .B(A[1]), .Z(n8992) );
  NAND U9797 ( .A(n9012), .B(n9013), .Z(n847) );
  NANDN U9798 ( .A(n9014), .B(n9015), .Z(n9013) );
  OR U9799 ( .A(n9016), .B(n9017), .Z(n9015) );
  NAND U9800 ( .A(n9017), .B(n9016), .Z(n9012) );
  XOR U9801 ( .A(n849), .B(n848), .Z(\A1[630] ) );
  XOR U9802 ( .A(n9017), .B(n9018), .Z(n848) );
  XNOR U9803 ( .A(n9016), .B(n9014), .Z(n9018) );
  AND U9804 ( .A(n9019), .B(n9020), .Z(n9014) );
  NANDN U9805 ( .A(n9021), .B(n9022), .Z(n9020) );
  NANDN U9806 ( .A(n9023), .B(n9024), .Z(n9022) );
  AND U9807 ( .A(B[629]), .B(A[3]), .Z(n9016) );
  XNOR U9808 ( .A(n9006), .B(n9025), .Z(n9017) );
  XNOR U9809 ( .A(n9004), .B(n9007), .Z(n9025) );
  NAND U9810 ( .A(A[2]), .B(B[630]), .Z(n9007) );
  NANDN U9811 ( .A(n9026), .B(n9027), .Z(n9004) );
  AND U9812 ( .A(A[0]), .B(B[631]), .Z(n9027) );
  XOR U9813 ( .A(n9009), .B(n9028), .Z(n9006) );
  NAND U9814 ( .A(A[0]), .B(B[632]), .Z(n9028) );
  NAND U9815 ( .A(B[631]), .B(A[1]), .Z(n9009) );
  NAND U9816 ( .A(n9029), .B(n9030), .Z(n849) );
  NANDN U9817 ( .A(n9031), .B(n9032), .Z(n9030) );
  OR U9818 ( .A(n9033), .B(n9034), .Z(n9032) );
  NAND U9819 ( .A(n9034), .B(n9033), .Z(n9029) );
  XOR U9820 ( .A(n831), .B(n830), .Z(\A1[62] ) );
  XOR U9821 ( .A(n8864), .B(n9035), .Z(n830) );
  XNOR U9822 ( .A(n8863), .B(n8861), .Z(n9035) );
  AND U9823 ( .A(n9036), .B(n9037), .Z(n8861) );
  NANDN U9824 ( .A(n9038), .B(n9039), .Z(n9037) );
  NANDN U9825 ( .A(n9040), .B(n9041), .Z(n9039) );
  AND U9826 ( .A(B[61]), .B(A[3]), .Z(n8863) );
  XNOR U9827 ( .A(n8853), .B(n9042), .Z(n8864) );
  XNOR U9828 ( .A(n8851), .B(n8854), .Z(n9042) );
  NAND U9829 ( .A(A[2]), .B(B[62]), .Z(n8854) );
  NANDN U9830 ( .A(n9043), .B(n9044), .Z(n8851) );
  AND U9831 ( .A(A[0]), .B(B[63]), .Z(n9044) );
  XOR U9832 ( .A(n8856), .B(n9045), .Z(n8853) );
  NAND U9833 ( .A(A[0]), .B(B[64]), .Z(n9045) );
  NAND U9834 ( .A(B[63]), .B(A[1]), .Z(n8856) );
  NAND U9835 ( .A(n9046), .B(n9047), .Z(n831) );
  NANDN U9836 ( .A(n9048), .B(n9049), .Z(n9047) );
  OR U9837 ( .A(n9050), .B(n9051), .Z(n9049) );
  NAND U9838 ( .A(n9051), .B(n9050), .Z(n9046) );
  XOR U9839 ( .A(n851), .B(n850), .Z(\A1[629] ) );
  XOR U9840 ( .A(n9034), .B(n9052), .Z(n850) );
  XNOR U9841 ( .A(n9033), .B(n9031), .Z(n9052) );
  AND U9842 ( .A(n9053), .B(n9054), .Z(n9031) );
  NANDN U9843 ( .A(n9055), .B(n9056), .Z(n9054) );
  NANDN U9844 ( .A(n9057), .B(n9058), .Z(n9056) );
  AND U9845 ( .A(B[628]), .B(A[3]), .Z(n9033) );
  XNOR U9846 ( .A(n9023), .B(n9059), .Z(n9034) );
  XNOR U9847 ( .A(n9021), .B(n9024), .Z(n9059) );
  NAND U9848 ( .A(A[2]), .B(B[629]), .Z(n9024) );
  NANDN U9849 ( .A(n9060), .B(n9061), .Z(n9021) );
  AND U9850 ( .A(A[0]), .B(B[630]), .Z(n9061) );
  XOR U9851 ( .A(n9026), .B(n9062), .Z(n9023) );
  NAND U9852 ( .A(A[0]), .B(B[631]), .Z(n9062) );
  NAND U9853 ( .A(B[630]), .B(A[1]), .Z(n9026) );
  NAND U9854 ( .A(n9063), .B(n9064), .Z(n851) );
  NANDN U9855 ( .A(n9065), .B(n9066), .Z(n9064) );
  OR U9856 ( .A(n9067), .B(n9068), .Z(n9066) );
  NAND U9857 ( .A(n9068), .B(n9067), .Z(n9063) );
  XOR U9858 ( .A(n855), .B(n854), .Z(\A1[628] ) );
  XOR U9859 ( .A(n9068), .B(n9069), .Z(n854) );
  XNOR U9860 ( .A(n9067), .B(n9065), .Z(n9069) );
  AND U9861 ( .A(n9070), .B(n9071), .Z(n9065) );
  NANDN U9862 ( .A(n9072), .B(n9073), .Z(n9071) );
  NANDN U9863 ( .A(n9074), .B(n9075), .Z(n9073) );
  AND U9864 ( .A(B[627]), .B(A[3]), .Z(n9067) );
  XNOR U9865 ( .A(n9057), .B(n9076), .Z(n9068) );
  XNOR U9866 ( .A(n9055), .B(n9058), .Z(n9076) );
  NAND U9867 ( .A(A[2]), .B(B[628]), .Z(n9058) );
  NANDN U9868 ( .A(n9077), .B(n9078), .Z(n9055) );
  AND U9869 ( .A(A[0]), .B(B[629]), .Z(n9078) );
  XOR U9870 ( .A(n9060), .B(n9079), .Z(n9057) );
  NAND U9871 ( .A(A[0]), .B(B[630]), .Z(n9079) );
  NAND U9872 ( .A(B[629]), .B(A[1]), .Z(n9060) );
  NAND U9873 ( .A(n9080), .B(n9081), .Z(n855) );
  NANDN U9874 ( .A(n9082), .B(n9083), .Z(n9081) );
  OR U9875 ( .A(n9084), .B(n9085), .Z(n9083) );
  NAND U9876 ( .A(n9085), .B(n9084), .Z(n9080) );
  XOR U9877 ( .A(n857), .B(n856), .Z(\A1[627] ) );
  XOR U9878 ( .A(n9085), .B(n9086), .Z(n856) );
  XNOR U9879 ( .A(n9084), .B(n9082), .Z(n9086) );
  AND U9880 ( .A(n9087), .B(n9088), .Z(n9082) );
  NANDN U9881 ( .A(n9089), .B(n9090), .Z(n9088) );
  NANDN U9882 ( .A(n9091), .B(n9092), .Z(n9090) );
  AND U9883 ( .A(B[626]), .B(A[3]), .Z(n9084) );
  XNOR U9884 ( .A(n9074), .B(n9093), .Z(n9085) );
  XNOR U9885 ( .A(n9072), .B(n9075), .Z(n9093) );
  NAND U9886 ( .A(A[2]), .B(B[627]), .Z(n9075) );
  NANDN U9887 ( .A(n9094), .B(n9095), .Z(n9072) );
  AND U9888 ( .A(A[0]), .B(B[628]), .Z(n9095) );
  XOR U9889 ( .A(n9077), .B(n9096), .Z(n9074) );
  NAND U9890 ( .A(A[0]), .B(B[629]), .Z(n9096) );
  NAND U9891 ( .A(B[628]), .B(A[1]), .Z(n9077) );
  NAND U9892 ( .A(n9097), .B(n9098), .Z(n857) );
  NANDN U9893 ( .A(n9099), .B(n9100), .Z(n9098) );
  OR U9894 ( .A(n9101), .B(n9102), .Z(n9100) );
  NAND U9895 ( .A(n9102), .B(n9101), .Z(n9097) );
  XOR U9896 ( .A(n859), .B(n858), .Z(\A1[626] ) );
  XOR U9897 ( .A(n9102), .B(n9103), .Z(n858) );
  XNOR U9898 ( .A(n9101), .B(n9099), .Z(n9103) );
  AND U9899 ( .A(n9104), .B(n9105), .Z(n9099) );
  NANDN U9900 ( .A(n9106), .B(n9107), .Z(n9105) );
  NANDN U9901 ( .A(n9108), .B(n9109), .Z(n9107) );
  AND U9902 ( .A(B[625]), .B(A[3]), .Z(n9101) );
  XNOR U9903 ( .A(n9091), .B(n9110), .Z(n9102) );
  XNOR U9904 ( .A(n9089), .B(n9092), .Z(n9110) );
  NAND U9905 ( .A(A[2]), .B(B[626]), .Z(n9092) );
  NANDN U9906 ( .A(n9111), .B(n9112), .Z(n9089) );
  AND U9907 ( .A(A[0]), .B(B[627]), .Z(n9112) );
  XOR U9908 ( .A(n9094), .B(n9113), .Z(n9091) );
  NAND U9909 ( .A(A[0]), .B(B[628]), .Z(n9113) );
  NAND U9910 ( .A(B[627]), .B(A[1]), .Z(n9094) );
  NAND U9911 ( .A(n9114), .B(n9115), .Z(n859) );
  NANDN U9912 ( .A(n9116), .B(n9117), .Z(n9115) );
  OR U9913 ( .A(n9118), .B(n9119), .Z(n9117) );
  NAND U9914 ( .A(n9119), .B(n9118), .Z(n9114) );
  XOR U9915 ( .A(n861), .B(n860), .Z(\A1[625] ) );
  XOR U9916 ( .A(n9119), .B(n9120), .Z(n860) );
  XNOR U9917 ( .A(n9118), .B(n9116), .Z(n9120) );
  AND U9918 ( .A(n9121), .B(n9122), .Z(n9116) );
  NANDN U9919 ( .A(n9123), .B(n9124), .Z(n9122) );
  NANDN U9920 ( .A(n9125), .B(n9126), .Z(n9124) );
  AND U9921 ( .A(B[624]), .B(A[3]), .Z(n9118) );
  XNOR U9922 ( .A(n9108), .B(n9127), .Z(n9119) );
  XNOR U9923 ( .A(n9106), .B(n9109), .Z(n9127) );
  NAND U9924 ( .A(A[2]), .B(B[625]), .Z(n9109) );
  NANDN U9925 ( .A(n9128), .B(n9129), .Z(n9106) );
  AND U9926 ( .A(A[0]), .B(B[626]), .Z(n9129) );
  XOR U9927 ( .A(n9111), .B(n9130), .Z(n9108) );
  NAND U9928 ( .A(A[0]), .B(B[627]), .Z(n9130) );
  NAND U9929 ( .A(B[626]), .B(A[1]), .Z(n9111) );
  NAND U9930 ( .A(n9131), .B(n9132), .Z(n861) );
  NANDN U9931 ( .A(n9133), .B(n9134), .Z(n9132) );
  OR U9932 ( .A(n9135), .B(n9136), .Z(n9134) );
  NAND U9933 ( .A(n9136), .B(n9135), .Z(n9131) );
  XOR U9934 ( .A(n863), .B(n862), .Z(\A1[624] ) );
  XOR U9935 ( .A(n9136), .B(n9137), .Z(n862) );
  XNOR U9936 ( .A(n9135), .B(n9133), .Z(n9137) );
  AND U9937 ( .A(n9138), .B(n9139), .Z(n9133) );
  NANDN U9938 ( .A(n9140), .B(n9141), .Z(n9139) );
  NANDN U9939 ( .A(n9142), .B(n9143), .Z(n9141) );
  AND U9940 ( .A(B[623]), .B(A[3]), .Z(n9135) );
  XNOR U9941 ( .A(n9125), .B(n9144), .Z(n9136) );
  XNOR U9942 ( .A(n9123), .B(n9126), .Z(n9144) );
  NAND U9943 ( .A(A[2]), .B(B[624]), .Z(n9126) );
  NANDN U9944 ( .A(n9145), .B(n9146), .Z(n9123) );
  AND U9945 ( .A(A[0]), .B(B[625]), .Z(n9146) );
  XOR U9946 ( .A(n9128), .B(n9147), .Z(n9125) );
  NAND U9947 ( .A(A[0]), .B(B[626]), .Z(n9147) );
  NAND U9948 ( .A(B[625]), .B(A[1]), .Z(n9128) );
  NAND U9949 ( .A(n9148), .B(n9149), .Z(n863) );
  NANDN U9950 ( .A(n9150), .B(n9151), .Z(n9149) );
  OR U9951 ( .A(n9152), .B(n9153), .Z(n9151) );
  NAND U9952 ( .A(n9153), .B(n9152), .Z(n9148) );
  XOR U9953 ( .A(n865), .B(n864), .Z(\A1[623] ) );
  XOR U9954 ( .A(n9153), .B(n9154), .Z(n864) );
  XNOR U9955 ( .A(n9152), .B(n9150), .Z(n9154) );
  AND U9956 ( .A(n9155), .B(n9156), .Z(n9150) );
  NANDN U9957 ( .A(n9157), .B(n9158), .Z(n9156) );
  NANDN U9958 ( .A(n9159), .B(n9160), .Z(n9158) );
  AND U9959 ( .A(B[622]), .B(A[3]), .Z(n9152) );
  XNOR U9960 ( .A(n9142), .B(n9161), .Z(n9153) );
  XNOR U9961 ( .A(n9140), .B(n9143), .Z(n9161) );
  NAND U9962 ( .A(A[2]), .B(B[623]), .Z(n9143) );
  NANDN U9963 ( .A(n9162), .B(n9163), .Z(n9140) );
  AND U9964 ( .A(A[0]), .B(B[624]), .Z(n9163) );
  XOR U9965 ( .A(n9145), .B(n9164), .Z(n9142) );
  NAND U9966 ( .A(A[0]), .B(B[625]), .Z(n9164) );
  NAND U9967 ( .A(B[624]), .B(A[1]), .Z(n9145) );
  NAND U9968 ( .A(n9165), .B(n9166), .Z(n865) );
  NANDN U9969 ( .A(n9167), .B(n9168), .Z(n9166) );
  OR U9970 ( .A(n9169), .B(n9170), .Z(n9168) );
  NAND U9971 ( .A(n9170), .B(n9169), .Z(n9165) );
  XOR U9972 ( .A(n867), .B(n866), .Z(\A1[622] ) );
  XOR U9973 ( .A(n9170), .B(n9171), .Z(n866) );
  XNOR U9974 ( .A(n9169), .B(n9167), .Z(n9171) );
  AND U9975 ( .A(n9172), .B(n9173), .Z(n9167) );
  NANDN U9976 ( .A(n9174), .B(n9175), .Z(n9173) );
  NANDN U9977 ( .A(n9176), .B(n9177), .Z(n9175) );
  AND U9978 ( .A(B[621]), .B(A[3]), .Z(n9169) );
  XNOR U9979 ( .A(n9159), .B(n9178), .Z(n9170) );
  XNOR U9980 ( .A(n9157), .B(n9160), .Z(n9178) );
  NAND U9981 ( .A(A[2]), .B(B[622]), .Z(n9160) );
  NANDN U9982 ( .A(n9179), .B(n9180), .Z(n9157) );
  AND U9983 ( .A(A[0]), .B(B[623]), .Z(n9180) );
  XOR U9984 ( .A(n9162), .B(n9181), .Z(n9159) );
  NAND U9985 ( .A(A[0]), .B(B[624]), .Z(n9181) );
  NAND U9986 ( .A(B[623]), .B(A[1]), .Z(n9162) );
  NAND U9987 ( .A(n9182), .B(n9183), .Z(n867) );
  NANDN U9988 ( .A(n9184), .B(n9185), .Z(n9183) );
  OR U9989 ( .A(n9186), .B(n9187), .Z(n9185) );
  NAND U9990 ( .A(n9187), .B(n9186), .Z(n9182) );
  XOR U9991 ( .A(n869), .B(n868), .Z(\A1[621] ) );
  XOR U9992 ( .A(n9187), .B(n9188), .Z(n868) );
  XNOR U9993 ( .A(n9186), .B(n9184), .Z(n9188) );
  AND U9994 ( .A(n9189), .B(n9190), .Z(n9184) );
  NANDN U9995 ( .A(n9191), .B(n9192), .Z(n9190) );
  NANDN U9996 ( .A(n9193), .B(n9194), .Z(n9192) );
  AND U9997 ( .A(B[620]), .B(A[3]), .Z(n9186) );
  XNOR U9998 ( .A(n9176), .B(n9195), .Z(n9187) );
  XNOR U9999 ( .A(n9174), .B(n9177), .Z(n9195) );
  NAND U10000 ( .A(A[2]), .B(B[621]), .Z(n9177) );
  NANDN U10001 ( .A(n9196), .B(n9197), .Z(n9174) );
  AND U10002 ( .A(A[0]), .B(B[622]), .Z(n9197) );
  XOR U10003 ( .A(n9179), .B(n9198), .Z(n9176) );
  NAND U10004 ( .A(A[0]), .B(B[623]), .Z(n9198) );
  NAND U10005 ( .A(B[622]), .B(A[1]), .Z(n9179) );
  NAND U10006 ( .A(n9199), .B(n9200), .Z(n869) );
  NANDN U10007 ( .A(n9201), .B(n9202), .Z(n9200) );
  OR U10008 ( .A(n9203), .B(n9204), .Z(n9202) );
  NAND U10009 ( .A(n9204), .B(n9203), .Z(n9199) );
  XOR U10010 ( .A(n871), .B(n870), .Z(\A1[620] ) );
  XOR U10011 ( .A(n9204), .B(n9205), .Z(n870) );
  XNOR U10012 ( .A(n9203), .B(n9201), .Z(n9205) );
  AND U10013 ( .A(n9206), .B(n9207), .Z(n9201) );
  NANDN U10014 ( .A(n9208), .B(n9209), .Z(n9207) );
  NANDN U10015 ( .A(n9210), .B(n9211), .Z(n9209) );
  AND U10016 ( .A(B[619]), .B(A[3]), .Z(n9203) );
  XNOR U10017 ( .A(n9193), .B(n9212), .Z(n9204) );
  XNOR U10018 ( .A(n9191), .B(n9194), .Z(n9212) );
  NAND U10019 ( .A(A[2]), .B(B[620]), .Z(n9194) );
  NANDN U10020 ( .A(n9213), .B(n9214), .Z(n9191) );
  AND U10021 ( .A(A[0]), .B(B[621]), .Z(n9214) );
  XOR U10022 ( .A(n9196), .B(n9215), .Z(n9193) );
  NAND U10023 ( .A(A[0]), .B(B[622]), .Z(n9215) );
  NAND U10024 ( .A(B[621]), .B(A[1]), .Z(n9196) );
  NAND U10025 ( .A(n9216), .B(n9217), .Z(n871) );
  NANDN U10026 ( .A(n9218), .B(n9219), .Z(n9217) );
  OR U10027 ( .A(n9220), .B(n9221), .Z(n9219) );
  NAND U10028 ( .A(n9221), .B(n9220), .Z(n9216) );
  XOR U10029 ( .A(n853), .B(n852), .Z(\A1[61] ) );
  XOR U10030 ( .A(n9051), .B(n9222), .Z(n852) );
  XNOR U10031 ( .A(n9050), .B(n9048), .Z(n9222) );
  AND U10032 ( .A(n9223), .B(n9224), .Z(n9048) );
  NANDN U10033 ( .A(n9225), .B(n9226), .Z(n9224) );
  NANDN U10034 ( .A(n9227), .B(n9228), .Z(n9226) );
  AND U10035 ( .A(B[60]), .B(A[3]), .Z(n9050) );
  XNOR U10036 ( .A(n9040), .B(n9229), .Z(n9051) );
  XNOR U10037 ( .A(n9038), .B(n9041), .Z(n9229) );
  NAND U10038 ( .A(A[2]), .B(B[61]), .Z(n9041) );
  NANDN U10039 ( .A(n9230), .B(n9231), .Z(n9038) );
  AND U10040 ( .A(A[0]), .B(B[62]), .Z(n9231) );
  XOR U10041 ( .A(n9043), .B(n9232), .Z(n9040) );
  NAND U10042 ( .A(A[0]), .B(B[63]), .Z(n9232) );
  NAND U10043 ( .A(B[62]), .B(A[1]), .Z(n9043) );
  NAND U10044 ( .A(n9233), .B(n9234), .Z(n853) );
  NANDN U10045 ( .A(n9235), .B(n9236), .Z(n9234) );
  OR U10046 ( .A(n9237), .B(n9238), .Z(n9236) );
  NAND U10047 ( .A(n9238), .B(n9237), .Z(n9233) );
  XOR U10048 ( .A(n873), .B(n872), .Z(\A1[619] ) );
  XOR U10049 ( .A(n9221), .B(n9239), .Z(n872) );
  XNOR U10050 ( .A(n9220), .B(n9218), .Z(n9239) );
  AND U10051 ( .A(n9240), .B(n9241), .Z(n9218) );
  NANDN U10052 ( .A(n9242), .B(n9243), .Z(n9241) );
  NANDN U10053 ( .A(n9244), .B(n9245), .Z(n9243) );
  AND U10054 ( .A(B[618]), .B(A[3]), .Z(n9220) );
  XNOR U10055 ( .A(n9210), .B(n9246), .Z(n9221) );
  XNOR U10056 ( .A(n9208), .B(n9211), .Z(n9246) );
  NAND U10057 ( .A(A[2]), .B(B[619]), .Z(n9211) );
  NANDN U10058 ( .A(n9247), .B(n9248), .Z(n9208) );
  AND U10059 ( .A(A[0]), .B(B[620]), .Z(n9248) );
  XOR U10060 ( .A(n9213), .B(n9249), .Z(n9210) );
  NAND U10061 ( .A(A[0]), .B(B[621]), .Z(n9249) );
  NAND U10062 ( .A(B[620]), .B(A[1]), .Z(n9213) );
  NAND U10063 ( .A(n9250), .B(n9251), .Z(n873) );
  NANDN U10064 ( .A(n9252), .B(n9253), .Z(n9251) );
  OR U10065 ( .A(n9254), .B(n9255), .Z(n9253) );
  NAND U10066 ( .A(n9255), .B(n9254), .Z(n9250) );
  XOR U10067 ( .A(n877), .B(n876), .Z(\A1[618] ) );
  XOR U10068 ( .A(n9255), .B(n9256), .Z(n876) );
  XNOR U10069 ( .A(n9254), .B(n9252), .Z(n9256) );
  AND U10070 ( .A(n9257), .B(n9258), .Z(n9252) );
  NANDN U10071 ( .A(n9259), .B(n9260), .Z(n9258) );
  NANDN U10072 ( .A(n9261), .B(n9262), .Z(n9260) );
  AND U10073 ( .A(B[617]), .B(A[3]), .Z(n9254) );
  XNOR U10074 ( .A(n9244), .B(n9263), .Z(n9255) );
  XNOR U10075 ( .A(n9242), .B(n9245), .Z(n9263) );
  NAND U10076 ( .A(A[2]), .B(B[618]), .Z(n9245) );
  NANDN U10077 ( .A(n9264), .B(n9265), .Z(n9242) );
  AND U10078 ( .A(A[0]), .B(B[619]), .Z(n9265) );
  XOR U10079 ( .A(n9247), .B(n9266), .Z(n9244) );
  NAND U10080 ( .A(A[0]), .B(B[620]), .Z(n9266) );
  NAND U10081 ( .A(B[619]), .B(A[1]), .Z(n9247) );
  NAND U10082 ( .A(n9267), .B(n9268), .Z(n877) );
  NANDN U10083 ( .A(n9269), .B(n9270), .Z(n9268) );
  OR U10084 ( .A(n9271), .B(n9272), .Z(n9270) );
  NAND U10085 ( .A(n9272), .B(n9271), .Z(n9267) );
  XOR U10086 ( .A(n879), .B(n878), .Z(\A1[617] ) );
  XOR U10087 ( .A(n9272), .B(n9273), .Z(n878) );
  XNOR U10088 ( .A(n9271), .B(n9269), .Z(n9273) );
  AND U10089 ( .A(n9274), .B(n9275), .Z(n9269) );
  NANDN U10090 ( .A(n9276), .B(n9277), .Z(n9275) );
  NANDN U10091 ( .A(n9278), .B(n9279), .Z(n9277) );
  AND U10092 ( .A(B[616]), .B(A[3]), .Z(n9271) );
  XNOR U10093 ( .A(n9261), .B(n9280), .Z(n9272) );
  XNOR U10094 ( .A(n9259), .B(n9262), .Z(n9280) );
  NAND U10095 ( .A(A[2]), .B(B[617]), .Z(n9262) );
  NANDN U10096 ( .A(n9281), .B(n9282), .Z(n9259) );
  AND U10097 ( .A(A[0]), .B(B[618]), .Z(n9282) );
  XOR U10098 ( .A(n9264), .B(n9283), .Z(n9261) );
  NAND U10099 ( .A(A[0]), .B(B[619]), .Z(n9283) );
  NAND U10100 ( .A(B[618]), .B(A[1]), .Z(n9264) );
  NAND U10101 ( .A(n9284), .B(n9285), .Z(n879) );
  NANDN U10102 ( .A(n9286), .B(n9287), .Z(n9285) );
  OR U10103 ( .A(n9288), .B(n9289), .Z(n9287) );
  NAND U10104 ( .A(n9289), .B(n9288), .Z(n9284) );
  XOR U10105 ( .A(n881), .B(n880), .Z(\A1[616] ) );
  XOR U10106 ( .A(n9289), .B(n9290), .Z(n880) );
  XNOR U10107 ( .A(n9288), .B(n9286), .Z(n9290) );
  AND U10108 ( .A(n9291), .B(n9292), .Z(n9286) );
  NANDN U10109 ( .A(n9293), .B(n9294), .Z(n9292) );
  NANDN U10110 ( .A(n9295), .B(n9296), .Z(n9294) );
  AND U10111 ( .A(B[615]), .B(A[3]), .Z(n9288) );
  XNOR U10112 ( .A(n9278), .B(n9297), .Z(n9289) );
  XNOR U10113 ( .A(n9276), .B(n9279), .Z(n9297) );
  NAND U10114 ( .A(A[2]), .B(B[616]), .Z(n9279) );
  NANDN U10115 ( .A(n9298), .B(n9299), .Z(n9276) );
  AND U10116 ( .A(A[0]), .B(B[617]), .Z(n9299) );
  XOR U10117 ( .A(n9281), .B(n9300), .Z(n9278) );
  NAND U10118 ( .A(A[0]), .B(B[618]), .Z(n9300) );
  NAND U10119 ( .A(B[617]), .B(A[1]), .Z(n9281) );
  NAND U10120 ( .A(n9301), .B(n9302), .Z(n881) );
  NANDN U10121 ( .A(n9303), .B(n9304), .Z(n9302) );
  OR U10122 ( .A(n9305), .B(n9306), .Z(n9304) );
  NAND U10123 ( .A(n9306), .B(n9305), .Z(n9301) );
  XOR U10124 ( .A(n883), .B(n882), .Z(\A1[615] ) );
  XOR U10125 ( .A(n9306), .B(n9307), .Z(n882) );
  XNOR U10126 ( .A(n9305), .B(n9303), .Z(n9307) );
  AND U10127 ( .A(n9308), .B(n9309), .Z(n9303) );
  NANDN U10128 ( .A(n9310), .B(n9311), .Z(n9309) );
  NANDN U10129 ( .A(n9312), .B(n9313), .Z(n9311) );
  AND U10130 ( .A(B[614]), .B(A[3]), .Z(n9305) );
  XNOR U10131 ( .A(n9295), .B(n9314), .Z(n9306) );
  XNOR U10132 ( .A(n9293), .B(n9296), .Z(n9314) );
  NAND U10133 ( .A(A[2]), .B(B[615]), .Z(n9296) );
  NANDN U10134 ( .A(n9315), .B(n9316), .Z(n9293) );
  AND U10135 ( .A(A[0]), .B(B[616]), .Z(n9316) );
  XOR U10136 ( .A(n9298), .B(n9317), .Z(n9295) );
  NAND U10137 ( .A(A[0]), .B(B[617]), .Z(n9317) );
  NAND U10138 ( .A(B[616]), .B(A[1]), .Z(n9298) );
  NAND U10139 ( .A(n9318), .B(n9319), .Z(n883) );
  NANDN U10140 ( .A(n9320), .B(n9321), .Z(n9319) );
  OR U10141 ( .A(n9322), .B(n9323), .Z(n9321) );
  NAND U10142 ( .A(n9323), .B(n9322), .Z(n9318) );
  XOR U10143 ( .A(n885), .B(n884), .Z(\A1[614] ) );
  XOR U10144 ( .A(n9323), .B(n9324), .Z(n884) );
  XNOR U10145 ( .A(n9322), .B(n9320), .Z(n9324) );
  AND U10146 ( .A(n9325), .B(n9326), .Z(n9320) );
  NANDN U10147 ( .A(n9327), .B(n9328), .Z(n9326) );
  NANDN U10148 ( .A(n9329), .B(n9330), .Z(n9328) );
  AND U10149 ( .A(B[613]), .B(A[3]), .Z(n9322) );
  XNOR U10150 ( .A(n9312), .B(n9331), .Z(n9323) );
  XNOR U10151 ( .A(n9310), .B(n9313), .Z(n9331) );
  NAND U10152 ( .A(A[2]), .B(B[614]), .Z(n9313) );
  NANDN U10153 ( .A(n9332), .B(n9333), .Z(n9310) );
  AND U10154 ( .A(A[0]), .B(B[615]), .Z(n9333) );
  XOR U10155 ( .A(n9315), .B(n9334), .Z(n9312) );
  NAND U10156 ( .A(A[0]), .B(B[616]), .Z(n9334) );
  NAND U10157 ( .A(B[615]), .B(A[1]), .Z(n9315) );
  NAND U10158 ( .A(n9335), .B(n9336), .Z(n885) );
  NANDN U10159 ( .A(n9337), .B(n9338), .Z(n9336) );
  OR U10160 ( .A(n9339), .B(n9340), .Z(n9338) );
  NAND U10161 ( .A(n9340), .B(n9339), .Z(n9335) );
  XOR U10162 ( .A(n887), .B(n886), .Z(\A1[613] ) );
  XOR U10163 ( .A(n9340), .B(n9341), .Z(n886) );
  XNOR U10164 ( .A(n9339), .B(n9337), .Z(n9341) );
  AND U10165 ( .A(n9342), .B(n9343), .Z(n9337) );
  NANDN U10166 ( .A(n9344), .B(n9345), .Z(n9343) );
  NANDN U10167 ( .A(n9346), .B(n9347), .Z(n9345) );
  AND U10168 ( .A(B[612]), .B(A[3]), .Z(n9339) );
  XNOR U10169 ( .A(n9329), .B(n9348), .Z(n9340) );
  XNOR U10170 ( .A(n9327), .B(n9330), .Z(n9348) );
  NAND U10171 ( .A(A[2]), .B(B[613]), .Z(n9330) );
  NANDN U10172 ( .A(n9349), .B(n9350), .Z(n9327) );
  AND U10173 ( .A(A[0]), .B(B[614]), .Z(n9350) );
  XOR U10174 ( .A(n9332), .B(n9351), .Z(n9329) );
  NAND U10175 ( .A(A[0]), .B(B[615]), .Z(n9351) );
  NAND U10176 ( .A(B[614]), .B(A[1]), .Z(n9332) );
  NAND U10177 ( .A(n9352), .B(n9353), .Z(n887) );
  NANDN U10178 ( .A(n9354), .B(n9355), .Z(n9353) );
  OR U10179 ( .A(n9356), .B(n9357), .Z(n9355) );
  NAND U10180 ( .A(n9357), .B(n9356), .Z(n9352) );
  XOR U10181 ( .A(n889), .B(n888), .Z(\A1[612] ) );
  XOR U10182 ( .A(n9357), .B(n9358), .Z(n888) );
  XNOR U10183 ( .A(n9356), .B(n9354), .Z(n9358) );
  AND U10184 ( .A(n9359), .B(n9360), .Z(n9354) );
  NANDN U10185 ( .A(n9361), .B(n9362), .Z(n9360) );
  NANDN U10186 ( .A(n9363), .B(n9364), .Z(n9362) );
  AND U10187 ( .A(B[611]), .B(A[3]), .Z(n9356) );
  XNOR U10188 ( .A(n9346), .B(n9365), .Z(n9357) );
  XNOR U10189 ( .A(n9344), .B(n9347), .Z(n9365) );
  NAND U10190 ( .A(A[2]), .B(B[612]), .Z(n9347) );
  NANDN U10191 ( .A(n9366), .B(n9367), .Z(n9344) );
  AND U10192 ( .A(A[0]), .B(B[613]), .Z(n9367) );
  XOR U10193 ( .A(n9349), .B(n9368), .Z(n9346) );
  NAND U10194 ( .A(A[0]), .B(B[614]), .Z(n9368) );
  NAND U10195 ( .A(B[613]), .B(A[1]), .Z(n9349) );
  NAND U10196 ( .A(n9369), .B(n9370), .Z(n889) );
  NANDN U10197 ( .A(n9371), .B(n9372), .Z(n9370) );
  OR U10198 ( .A(n9373), .B(n9374), .Z(n9372) );
  NAND U10199 ( .A(n9374), .B(n9373), .Z(n9369) );
  XOR U10200 ( .A(n891), .B(n890), .Z(\A1[611] ) );
  XOR U10201 ( .A(n9374), .B(n9375), .Z(n890) );
  XNOR U10202 ( .A(n9373), .B(n9371), .Z(n9375) );
  AND U10203 ( .A(n9376), .B(n9377), .Z(n9371) );
  NANDN U10204 ( .A(n9378), .B(n9379), .Z(n9377) );
  NANDN U10205 ( .A(n9380), .B(n9381), .Z(n9379) );
  AND U10206 ( .A(B[610]), .B(A[3]), .Z(n9373) );
  XNOR U10207 ( .A(n9363), .B(n9382), .Z(n9374) );
  XNOR U10208 ( .A(n9361), .B(n9364), .Z(n9382) );
  NAND U10209 ( .A(A[2]), .B(B[611]), .Z(n9364) );
  NANDN U10210 ( .A(n9383), .B(n9384), .Z(n9361) );
  AND U10211 ( .A(A[0]), .B(B[612]), .Z(n9384) );
  XOR U10212 ( .A(n9366), .B(n9385), .Z(n9363) );
  NAND U10213 ( .A(A[0]), .B(B[613]), .Z(n9385) );
  NAND U10214 ( .A(B[612]), .B(A[1]), .Z(n9366) );
  NAND U10215 ( .A(n9386), .B(n9387), .Z(n891) );
  NANDN U10216 ( .A(n9388), .B(n9389), .Z(n9387) );
  OR U10217 ( .A(n9390), .B(n9391), .Z(n9389) );
  NAND U10218 ( .A(n9391), .B(n9390), .Z(n9386) );
  XOR U10219 ( .A(n893), .B(n892), .Z(\A1[610] ) );
  XOR U10220 ( .A(n9391), .B(n9392), .Z(n892) );
  XNOR U10221 ( .A(n9390), .B(n9388), .Z(n9392) );
  AND U10222 ( .A(n9393), .B(n9394), .Z(n9388) );
  NANDN U10223 ( .A(n9395), .B(n9396), .Z(n9394) );
  NANDN U10224 ( .A(n9397), .B(n9398), .Z(n9396) );
  AND U10225 ( .A(B[609]), .B(A[3]), .Z(n9390) );
  XNOR U10226 ( .A(n9380), .B(n9399), .Z(n9391) );
  XNOR U10227 ( .A(n9378), .B(n9381), .Z(n9399) );
  NAND U10228 ( .A(A[2]), .B(B[610]), .Z(n9381) );
  NANDN U10229 ( .A(n9400), .B(n9401), .Z(n9378) );
  AND U10230 ( .A(A[0]), .B(B[611]), .Z(n9401) );
  XOR U10231 ( .A(n9383), .B(n9402), .Z(n9380) );
  NAND U10232 ( .A(A[0]), .B(B[612]), .Z(n9402) );
  NAND U10233 ( .A(B[611]), .B(A[1]), .Z(n9383) );
  NAND U10234 ( .A(n9403), .B(n9404), .Z(n893) );
  NANDN U10235 ( .A(n9405), .B(n9406), .Z(n9404) );
  OR U10236 ( .A(n9407), .B(n9408), .Z(n9406) );
  NAND U10237 ( .A(n9408), .B(n9407), .Z(n9403) );
  XOR U10238 ( .A(n875), .B(n874), .Z(\A1[60] ) );
  XOR U10239 ( .A(n9238), .B(n9409), .Z(n874) );
  XNOR U10240 ( .A(n9237), .B(n9235), .Z(n9409) );
  AND U10241 ( .A(n9410), .B(n9411), .Z(n9235) );
  NANDN U10242 ( .A(n9412), .B(n9413), .Z(n9411) );
  NANDN U10243 ( .A(n9414), .B(n9415), .Z(n9413) );
  AND U10244 ( .A(B[59]), .B(A[3]), .Z(n9237) );
  XNOR U10245 ( .A(n9227), .B(n9416), .Z(n9238) );
  XNOR U10246 ( .A(n9225), .B(n9228), .Z(n9416) );
  NAND U10247 ( .A(A[2]), .B(B[60]), .Z(n9228) );
  NANDN U10248 ( .A(n9417), .B(n9418), .Z(n9225) );
  AND U10249 ( .A(A[0]), .B(B[61]), .Z(n9418) );
  XOR U10250 ( .A(n9230), .B(n9419), .Z(n9227) );
  NAND U10251 ( .A(A[0]), .B(B[62]), .Z(n9419) );
  NAND U10252 ( .A(B[61]), .B(A[1]), .Z(n9230) );
  NAND U10253 ( .A(n9420), .B(n9421), .Z(n875) );
  NANDN U10254 ( .A(n9422), .B(n9423), .Z(n9421) );
  OR U10255 ( .A(n9424), .B(n9425), .Z(n9423) );
  NAND U10256 ( .A(n9425), .B(n9424), .Z(n9420) );
  XOR U10257 ( .A(n895), .B(n894), .Z(\A1[609] ) );
  XOR U10258 ( .A(n9408), .B(n9426), .Z(n894) );
  XNOR U10259 ( .A(n9407), .B(n9405), .Z(n9426) );
  AND U10260 ( .A(n9427), .B(n9428), .Z(n9405) );
  NANDN U10261 ( .A(n9429), .B(n9430), .Z(n9428) );
  NANDN U10262 ( .A(n9431), .B(n9432), .Z(n9430) );
  AND U10263 ( .A(B[608]), .B(A[3]), .Z(n9407) );
  XNOR U10264 ( .A(n9397), .B(n9433), .Z(n9408) );
  XNOR U10265 ( .A(n9395), .B(n9398), .Z(n9433) );
  NAND U10266 ( .A(A[2]), .B(B[609]), .Z(n9398) );
  NANDN U10267 ( .A(n9434), .B(n9435), .Z(n9395) );
  AND U10268 ( .A(A[0]), .B(B[610]), .Z(n9435) );
  XOR U10269 ( .A(n9400), .B(n9436), .Z(n9397) );
  NAND U10270 ( .A(A[0]), .B(B[611]), .Z(n9436) );
  NAND U10271 ( .A(B[610]), .B(A[1]), .Z(n9400) );
  NAND U10272 ( .A(n9437), .B(n9438), .Z(n895) );
  NANDN U10273 ( .A(n9439), .B(n9440), .Z(n9438) );
  OR U10274 ( .A(n9441), .B(n9442), .Z(n9440) );
  NAND U10275 ( .A(n9442), .B(n9441), .Z(n9437) );
  XOR U10276 ( .A(n899), .B(n898), .Z(\A1[608] ) );
  XOR U10277 ( .A(n9442), .B(n9443), .Z(n898) );
  XNOR U10278 ( .A(n9441), .B(n9439), .Z(n9443) );
  AND U10279 ( .A(n9444), .B(n9445), .Z(n9439) );
  NANDN U10280 ( .A(n9446), .B(n9447), .Z(n9445) );
  NANDN U10281 ( .A(n9448), .B(n9449), .Z(n9447) );
  AND U10282 ( .A(B[607]), .B(A[3]), .Z(n9441) );
  XNOR U10283 ( .A(n9431), .B(n9450), .Z(n9442) );
  XNOR U10284 ( .A(n9429), .B(n9432), .Z(n9450) );
  NAND U10285 ( .A(A[2]), .B(B[608]), .Z(n9432) );
  NANDN U10286 ( .A(n9451), .B(n9452), .Z(n9429) );
  AND U10287 ( .A(A[0]), .B(B[609]), .Z(n9452) );
  XOR U10288 ( .A(n9434), .B(n9453), .Z(n9431) );
  NAND U10289 ( .A(A[0]), .B(B[610]), .Z(n9453) );
  NAND U10290 ( .A(B[609]), .B(A[1]), .Z(n9434) );
  NAND U10291 ( .A(n9454), .B(n9455), .Z(n899) );
  NANDN U10292 ( .A(n9456), .B(n9457), .Z(n9455) );
  OR U10293 ( .A(n9458), .B(n9459), .Z(n9457) );
  NAND U10294 ( .A(n9459), .B(n9458), .Z(n9454) );
  XOR U10295 ( .A(n901), .B(n900), .Z(\A1[607] ) );
  XOR U10296 ( .A(n9459), .B(n9460), .Z(n900) );
  XNOR U10297 ( .A(n9458), .B(n9456), .Z(n9460) );
  AND U10298 ( .A(n9461), .B(n9462), .Z(n9456) );
  NANDN U10299 ( .A(n9463), .B(n9464), .Z(n9462) );
  NANDN U10300 ( .A(n9465), .B(n9466), .Z(n9464) );
  AND U10301 ( .A(B[606]), .B(A[3]), .Z(n9458) );
  XNOR U10302 ( .A(n9448), .B(n9467), .Z(n9459) );
  XNOR U10303 ( .A(n9446), .B(n9449), .Z(n9467) );
  NAND U10304 ( .A(A[2]), .B(B[607]), .Z(n9449) );
  NANDN U10305 ( .A(n9468), .B(n9469), .Z(n9446) );
  AND U10306 ( .A(A[0]), .B(B[608]), .Z(n9469) );
  XOR U10307 ( .A(n9451), .B(n9470), .Z(n9448) );
  NAND U10308 ( .A(A[0]), .B(B[609]), .Z(n9470) );
  NAND U10309 ( .A(B[608]), .B(A[1]), .Z(n9451) );
  NAND U10310 ( .A(n9471), .B(n9472), .Z(n901) );
  NANDN U10311 ( .A(n9473), .B(n9474), .Z(n9472) );
  OR U10312 ( .A(n9475), .B(n9476), .Z(n9474) );
  NAND U10313 ( .A(n9476), .B(n9475), .Z(n9471) );
  XOR U10314 ( .A(n903), .B(n902), .Z(\A1[606] ) );
  XOR U10315 ( .A(n9476), .B(n9477), .Z(n902) );
  XNOR U10316 ( .A(n9475), .B(n9473), .Z(n9477) );
  AND U10317 ( .A(n9478), .B(n9479), .Z(n9473) );
  NANDN U10318 ( .A(n9480), .B(n9481), .Z(n9479) );
  NANDN U10319 ( .A(n9482), .B(n9483), .Z(n9481) );
  AND U10320 ( .A(B[605]), .B(A[3]), .Z(n9475) );
  XNOR U10321 ( .A(n9465), .B(n9484), .Z(n9476) );
  XNOR U10322 ( .A(n9463), .B(n9466), .Z(n9484) );
  NAND U10323 ( .A(A[2]), .B(B[606]), .Z(n9466) );
  NANDN U10324 ( .A(n9485), .B(n9486), .Z(n9463) );
  AND U10325 ( .A(A[0]), .B(B[607]), .Z(n9486) );
  XOR U10326 ( .A(n9468), .B(n9487), .Z(n9465) );
  NAND U10327 ( .A(A[0]), .B(B[608]), .Z(n9487) );
  NAND U10328 ( .A(B[607]), .B(A[1]), .Z(n9468) );
  NAND U10329 ( .A(n9488), .B(n9489), .Z(n903) );
  NANDN U10330 ( .A(n9490), .B(n9491), .Z(n9489) );
  OR U10331 ( .A(n9492), .B(n9493), .Z(n9491) );
  NAND U10332 ( .A(n9493), .B(n9492), .Z(n9488) );
  XOR U10333 ( .A(n905), .B(n904), .Z(\A1[605] ) );
  XOR U10334 ( .A(n9493), .B(n9494), .Z(n904) );
  XNOR U10335 ( .A(n9492), .B(n9490), .Z(n9494) );
  AND U10336 ( .A(n9495), .B(n9496), .Z(n9490) );
  NANDN U10337 ( .A(n9497), .B(n9498), .Z(n9496) );
  NANDN U10338 ( .A(n9499), .B(n9500), .Z(n9498) );
  AND U10339 ( .A(B[604]), .B(A[3]), .Z(n9492) );
  XNOR U10340 ( .A(n9482), .B(n9501), .Z(n9493) );
  XNOR U10341 ( .A(n9480), .B(n9483), .Z(n9501) );
  NAND U10342 ( .A(A[2]), .B(B[605]), .Z(n9483) );
  NANDN U10343 ( .A(n9502), .B(n9503), .Z(n9480) );
  AND U10344 ( .A(A[0]), .B(B[606]), .Z(n9503) );
  XOR U10345 ( .A(n9485), .B(n9504), .Z(n9482) );
  NAND U10346 ( .A(A[0]), .B(B[607]), .Z(n9504) );
  NAND U10347 ( .A(B[606]), .B(A[1]), .Z(n9485) );
  NAND U10348 ( .A(n9505), .B(n9506), .Z(n905) );
  NANDN U10349 ( .A(n9507), .B(n9508), .Z(n9506) );
  OR U10350 ( .A(n9509), .B(n9510), .Z(n9508) );
  NAND U10351 ( .A(n9510), .B(n9509), .Z(n9505) );
  XOR U10352 ( .A(n907), .B(n906), .Z(\A1[604] ) );
  XOR U10353 ( .A(n9510), .B(n9511), .Z(n906) );
  XNOR U10354 ( .A(n9509), .B(n9507), .Z(n9511) );
  AND U10355 ( .A(n9512), .B(n9513), .Z(n9507) );
  NANDN U10356 ( .A(n9514), .B(n9515), .Z(n9513) );
  NANDN U10357 ( .A(n9516), .B(n9517), .Z(n9515) );
  AND U10358 ( .A(B[603]), .B(A[3]), .Z(n9509) );
  XNOR U10359 ( .A(n9499), .B(n9518), .Z(n9510) );
  XNOR U10360 ( .A(n9497), .B(n9500), .Z(n9518) );
  NAND U10361 ( .A(A[2]), .B(B[604]), .Z(n9500) );
  NANDN U10362 ( .A(n9519), .B(n9520), .Z(n9497) );
  AND U10363 ( .A(A[0]), .B(B[605]), .Z(n9520) );
  XOR U10364 ( .A(n9502), .B(n9521), .Z(n9499) );
  NAND U10365 ( .A(A[0]), .B(B[606]), .Z(n9521) );
  NAND U10366 ( .A(B[605]), .B(A[1]), .Z(n9502) );
  NAND U10367 ( .A(n9522), .B(n9523), .Z(n907) );
  NANDN U10368 ( .A(n9524), .B(n9525), .Z(n9523) );
  OR U10369 ( .A(n9526), .B(n9527), .Z(n9525) );
  NAND U10370 ( .A(n9527), .B(n9526), .Z(n9522) );
  XOR U10371 ( .A(n909), .B(n908), .Z(\A1[603] ) );
  XOR U10372 ( .A(n9527), .B(n9528), .Z(n908) );
  XNOR U10373 ( .A(n9526), .B(n9524), .Z(n9528) );
  AND U10374 ( .A(n9529), .B(n9530), .Z(n9524) );
  NANDN U10375 ( .A(n9531), .B(n9532), .Z(n9530) );
  NANDN U10376 ( .A(n9533), .B(n9534), .Z(n9532) );
  AND U10377 ( .A(B[602]), .B(A[3]), .Z(n9526) );
  XNOR U10378 ( .A(n9516), .B(n9535), .Z(n9527) );
  XNOR U10379 ( .A(n9514), .B(n9517), .Z(n9535) );
  NAND U10380 ( .A(A[2]), .B(B[603]), .Z(n9517) );
  NANDN U10381 ( .A(n9536), .B(n9537), .Z(n9514) );
  AND U10382 ( .A(A[0]), .B(B[604]), .Z(n9537) );
  XOR U10383 ( .A(n9519), .B(n9538), .Z(n9516) );
  NAND U10384 ( .A(A[0]), .B(B[605]), .Z(n9538) );
  NAND U10385 ( .A(B[604]), .B(A[1]), .Z(n9519) );
  NAND U10386 ( .A(n9539), .B(n9540), .Z(n909) );
  NANDN U10387 ( .A(n9541), .B(n9542), .Z(n9540) );
  OR U10388 ( .A(n9543), .B(n9544), .Z(n9542) );
  NAND U10389 ( .A(n9544), .B(n9543), .Z(n9539) );
  XOR U10390 ( .A(n911), .B(n910), .Z(\A1[602] ) );
  XOR U10391 ( .A(n9544), .B(n9545), .Z(n910) );
  XNOR U10392 ( .A(n9543), .B(n9541), .Z(n9545) );
  AND U10393 ( .A(n9546), .B(n9547), .Z(n9541) );
  NANDN U10394 ( .A(n9548), .B(n9549), .Z(n9547) );
  NANDN U10395 ( .A(n9550), .B(n9551), .Z(n9549) );
  AND U10396 ( .A(B[601]), .B(A[3]), .Z(n9543) );
  XNOR U10397 ( .A(n9533), .B(n9552), .Z(n9544) );
  XNOR U10398 ( .A(n9531), .B(n9534), .Z(n9552) );
  NAND U10399 ( .A(A[2]), .B(B[602]), .Z(n9534) );
  NANDN U10400 ( .A(n9553), .B(n9554), .Z(n9531) );
  AND U10401 ( .A(A[0]), .B(B[603]), .Z(n9554) );
  XOR U10402 ( .A(n9536), .B(n9555), .Z(n9533) );
  NAND U10403 ( .A(A[0]), .B(B[604]), .Z(n9555) );
  NAND U10404 ( .A(B[603]), .B(A[1]), .Z(n9536) );
  NAND U10405 ( .A(n9556), .B(n9557), .Z(n911) );
  NANDN U10406 ( .A(n9558), .B(n9559), .Z(n9557) );
  OR U10407 ( .A(n9560), .B(n9561), .Z(n9559) );
  NAND U10408 ( .A(n9561), .B(n9560), .Z(n9556) );
  XOR U10409 ( .A(n913), .B(n912), .Z(\A1[601] ) );
  XOR U10410 ( .A(n9561), .B(n9562), .Z(n912) );
  XNOR U10411 ( .A(n9560), .B(n9558), .Z(n9562) );
  AND U10412 ( .A(n9563), .B(n9564), .Z(n9558) );
  NANDN U10413 ( .A(n9565), .B(n9566), .Z(n9564) );
  NANDN U10414 ( .A(n9567), .B(n9568), .Z(n9566) );
  AND U10415 ( .A(B[600]), .B(A[3]), .Z(n9560) );
  XNOR U10416 ( .A(n9550), .B(n9569), .Z(n9561) );
  XNOR U10417 ( .A(n9548), .B(n9551), .Z(n9569) );
  NAND U10418 ( .A(A[2]), .B(B[601]), .Z(n9551) );
  NANDN U10419 ( .A(n9570), .B(n9571), .Z(n9548) );
  AND U10420 ( .A(A[0]), .B(B[602]), .Z(n9571) );
  XOR U10421 ( .A(n9553), .B(n9572), .Z(n9550) );
  NAND U10422 ( .A(A[0]), .B(B[603]), .Z(n9572) );
  NAND U10423 ( .A(B[602]), .B(A[1]), .Z(n9553) );
  NAND U10424 ( .A(n9573), .B(n9574), .Z(n913) );
  NANDN U10425 ( .A(n9575), .B(n9576), .Z(n9574) );
  OR U10426 ( .A(n9577), .B(n9578), .Z(n9576) );
  NAND U10427 ( .A(n9578), .B(n9577), .Z(n9573) );
  XOR U10428 ( .A(n915), .B(n914), .Z(\A1[600] ) );
  XOR U10429 ( .A(n9578), .B(n9579), .Z(n914) );
  XNOR U10430 ( .A(n9577), .B(n9575), .Z(n9579) );
  AND U10431 ( .A(n9580), .B(n9581), .Z(n9575) );
  NANDN U10432 ( .A(n9582), .B(n9583), .Z(n9581) );
  NANDN U10433 ( .A(n9584), .B(n9585), .Z(n9583) );
  AND U10434 ( .A(B[599]), .B(A[3]), .Z(n9577) );
  XNOR U10435 ( .A(n9567), .B(n9586), .Z(n9578) );
  XNOR U10436 ( .A(n9565), .B(n9568), .Z(n9586) );
  NAND U10437 ( .A(A[2]), .B(B[600]), .Z(n9568) );
  NANDN U10438 ( .A(n9587), .B(n9588), .Z(n9565) );
  AND U10439 ( .A(A[0]), .B(B[601]), .Z(n9588) );
  XOR U10440 ( .A(n9570), .B(n9589), .Z(n9567) );
  NAND U10441 ( .A(A[0]), .B(B[602]), .Z(n9589) );
  NAND U10442 ( .A(B[601]), .B(A[1]), .Z(n9570) );
  NAND U10443 ( .A(n9590), .B(n9591), .Z(n915) );
  NANDN U10444 ( .A(n9592), .B(n9593), .Z(n9591) );
  OR U10445 ( .A(n9594), .B(n9595), .Z(n9593) );
  NAND U10446 ( .A(n9595), .B(n9594), .Z(n9590) );
  XOR U10447 ( .A(n697), .B(n696), .Z(\A1[5] ) );
  XOR U10448 ( .A(n7725), .B(n9596), .Z(n696) );
  XNOR U10449 ( .A(n7724), .B(n7722), .Z(n9596) );
  AND U10450 ( .A(n9597), .B(n9598), .Z(n7722) );
  NANDN U10451 ( .A(n9599), .B(n9600), .Z(n9598) );
  NANDN U10452 ( .A(n9601), .B(n9602), .Z(n9600) );
  AND U10453 ( .A(B[4]), .B(A[3]), .Z(n7724) );
  XNOR U10454 ( .A(n7714), .B(n9603), .Z(n7725) );
  XNOR U10455 ( .A(n7712), .B(n7715), .Z(n9603) );
  NAND U10456 ( .A(A[2]), .B(B[5]), .Z(n7715) );
  NANDN U10457 ( .A(n9604), .B(n9605), .Z(n7712) );
  AND U10458 ( .A(A[0]), .B(B[6]), .Z(n9605) );
  XOR U10459 ( .A(n7718), .B(n9606), .Z(n7714) );
  NAND U10460 ( .A(A[0]), .B(B[7]), .Z(n9606) );
  NAND U10461 ( .A(B[6]), .B(A[1]), .Z(n7718) );
  NAND U10462 ( .A(n9607), .B(n9608), .Z(n697) );
  NANDN U10463 ( .A(n9609), .B(n9610), .Z(n9608) );
  OR U10464 ( .A(n9611), .B(n9612), .Z(n9610) );
  NAND U10465 ( .A(n9612), .B(n9611), .Z(n9607) );
  XOR U10466 ( .A(n897), .B(n896), .Z(\A1[59] ) );
  XOR U10467 ( .A(n9425), .B(n9613), .Z(n896) );
  XNOR U10468 ( .A(n9424), .B(n9422), .Z(n9613) );
  AND U10469 ( .A(n9614), .B(n9615), .Z(n9422) );
  NANDN U10470 ( .A(n9616), .B(n9617), .Z(n9615) );
  NANDN U10471 ( .A(n9618), .B(n9619), .Z(n9617) );
  AND U10472 ( .A(B[58]), .B(A[3]), .Z(n9424) );
  XNOR U10473 ( .A(n9414), .B(n9620), .Z(n9425) );
  XNOR U10474 ( .A(n9412), .B(n9415), .Z(n9620) );
  NAND U10475 ( .A(A[2]), .B(B[59]), .Z(n9415) );
  NANDN U10476 ( .A(n9621), .B(n9622), .Z(n9412) );
  AND U10477 ( .A(A[0]), .B(B[60]), .Z(n9622) );
  XOR U10478 ( .A(n9417), .B(n9623), .Z(n9414) );
  NAND U10479 ( .A(A[0]), .B(B[61]), .Z(n9623) );
  NAND U10480 ( .A(B[60]), .B(A[1]), .Z(n9417) );
  NAND U10481 ( .A(n9624), .B(n9625), .Z(n897) );
  NANDN U10482 ( .A(n9626), .B(n9627), .Z(n9625) );
  OR U10483 ( .A(n9628), .B(n9629), .Z(n9627) );
  NAND U10484 ( .A(n9629), .B(n9628), .Z(n9624) );
  XOR U10485 ( .A(n917), .B(n916), .Z(\A1[599] ) );
  XOR U10486 ( .A(n9595), .B(n9630), .Z(n916) );
  XNOR U10487 ( .A(n9594), .B(n9592), .Z(n9630) );
  AND U10488 ( .A(n9631), .B(n9632), .Z(n9592) );
  NANDN U10489 ( .A(n9633), .B(n9634), .Z(n9632) );
  NANDN U10490 ( .A(n9635), .B(n9636), .Z(n9634) );
  AND U10491 ( .A(B[598]), .B(A[3]), .Z(n9594) );
  XNOR U10492 ( .A(n9584), .B(n9637), .Z(n9595) );
  XNOR U10493 ( .A(n9582), .B(n9585), .Z(n9637) );
  NAND U10494 ( .A(A[2]), .B(B[599]), .Z(n9585) );
  NANDN U10495 ( .A(n9638), .B(n9639), .Z(n9582) );
  AND U10496 ( .A(A[0]), .B(B[600]), .Z(n9639) );
  XOR U10497 ( .A(n9587), .B(n9640), .Z(n9584) );
  NAND U10498 ( .A(A[0]), .B(B[601]), .Z(n9640) );
  NAND U10499 ( .A(B[600]), .B(A[1]), .Z(n9587) );
  NAND U10500 ( .A(n9641), .B(n9642), .Z(n917) );
  NANDN U10501 ( .A(n9643), .B(n9644), .Z(n9642) );
  OR U10502 ( .A(n9645), .B(n9646), .Z(n9644) );
  NAND U10503 ( .A(n9646), .B(n9645), .Z(n9641) );
  XOR U10504 ( .A(n923), .B(n922), .Z(\A1[598] ) );
  XOR U10505 ( .A(n9646), .B(n9647), .Z(n922) );
  XNOR U10506 ( .A(n9645), .B(n9643), .Z(n9647) );
  AND U10507 ( .A(n9648), .B(n9649), .Z(n9643) );
  NANDN U10508 ( .A(n9650), .B(n9651), .Z(n9649) );
  NANDN U10509 ( .A(n9652), .B(n9653), .Z(n9651) );
  AND U10510 ( .A(B[597]), .B(A[3]), .Z(n9645) );
  XNOR U10511 ( .A(n9635), .B(n9654), .Z(n9646) );
  XNOR U10512 ( .A(n9633), .B(n9636), .Z(n9654) );
  NAND U10513 ( .A(A[2]), .B(B[598]), .Z(n9636) );
  NANDN U10514 ( .A(n9655), .B(n9656), .Z(n9633) );
  AND U10515 ( .A(A[0]), .B(B[599]), .Z(n9656) );
  XOR U10516 ( .A(n9638), .B(n9657), .Z(n9635) );
  NAND U10517 ( .A(A[0]), .B(B[600]), .Z(n9657) );
  NAND U10518 ( .A(B[599]), .B(A[1]), .Z(n9638) );
  NAND U10519 ( .A(n9658), .B(n9659), .Z(n923) );
  NANDN U10520 ( .A(n9660), .B(n9661), .Z(n9659) );
  OR U10521 ( .A(n9662), .B(n9663), .Z(n9661) );
  NAND U10522 ( .A(n9663), .B(n9662), .Z(n9658) );
  XOR U10523 ( .A(n925), .B(n924), .Z(\A1[597] ) );
  XOR U10524 ( .A(n9663), .B(n9664), .Z(n924) );
  XNOR U10525 ( .A(n9662), .B(n9660), .Z(n9664) );
  AND U10526 ( .A(n9665), .B(n9666), .Z(n9660) );
  NANDN U10527 ( .A(n9667), .B(n9668), .Z(n9666) );
  NANDN U10528 ( .A(n9669), .B(n9670), .Z(n9668) );
  AND U10529 ( .A(B[596]), .B(A[3]), .Z(n9662) );
  XNOR U10530 ( .A(n9652), .B(n9671), .Z(n9663) );
  XNOR U10531 ( .A(n9650), .B(n9653), .Z(n9671) );
  NAND U10532 ( .A(A[2]), .B(B[597]), .Z(n9653) );
  NANDN U10533 ( .A(n9672), .B(n9673), .Z(n9650) );
  AND U10534 ( .A(A[0]), .B(B[598]), .Z(n9673) );
  XOR U10535 ( .A(n9655), .B(n9674), .Z(n9652) );
  NAND U10536 ( .A(A[0]), .B(B[599]), .Z(n9674) );
  NAND U10537 ( .A(B[598]), .B(A[1]), .Z(n9655) );
  NAND U10538 ( .A(n9675), .B(n9676), .Z(n925) );
  NANDN U10539 ( .A(n9677), .B(n9678), .Z(n9676) );
  OR U10540 ( .A(n9679), .B(n9680), .Z(n9678) );
  NAND U10541 ( .A(n9680), .B(n9679), .Z(n9675) );
  XOR U10542 ( .A(n927), .B(n926), .Z(\A1[596] ) );
  XOR U10543 ( .A(n9680), .B(n9681), .Z(n926) );
  XNOR U10544 ( .A(n9679), .B(n9677), .Z(n9681) );
  AND U10545 ( .A(n9682), .B(n9683), .Z(n9677) );
  NANDN U10546 ( .A(n9684), .B(n9685), .Z(n9683) );
  NANDN U10547 ( .A(n9686), .B(n9687), .Z(n9685) );
  AND U10548 ( .A(B[595]), .B(A[3]), .Z(n9679) );
  XNOR U10549 ( .A(n9669), .B(n9688), .Z(n9680) );
  XNOR U10550 ( .A(n9667), .B(n9670), .Z(n9688) );
  NAND U10551 ( .A(A[2]), .B(B[596]), .Z(n9670) );
  NANDN U10552 ( .A(n9689), .B(n9690), .Z(n9667) );
  AND U10553 ( .A(A[0]), .B(B[597]), .Z(n9690) );
  XOR U10554 ( .A(n9672), .B(n9691), .Z(n9669) );
  NAND U10555 ( .A(A[0]), .B(B[598]), .Z(n9691) );
  NAND U10556 ( .A(B[597]), .B(A[1]), .Z(n9672) );
  NAND U10557 ( .A(n9692), .B(n9693), .Z(n927) );
  NANDN U10558 ( .A(n9694), .B(n9695), .Z(n9693) );
  OR U10559 ( .A(n9696), .B(n9697), .Z(n9695) );
  NAND U10560 ( .A(n9697), .B(n9696), .Z(n9692) );
  XOR U10561 ( .A(n929), .B(n928), .Z(\A1[595] ) );
  XOR U10562 ( .A(n9697), .B(n9698), .Z(n928) );
  XNOR U10563 ( .A(n9696), .B(n9694), .Z(n9698) );
  AND U10564 ( .A(n9699), .B(n9700), .Z(n9694) );
  NANDN U10565 ( .A(n9701), .B(n9702), .Z(n9700) );
  NANDN U10566 ( .A(n9703), .B(n9704), .Z(n9702) );
  AND U10567 ( .A(B[594]), .B(A[3]), .Z(n9696) );
  XNOR U10568 ( .A(n9686), .B(n9705), .Z(n9697) );
  XNOR U10569 ( .A(n9684), .B(n9687), .Z(n9705) );
  NAND U10570 ( .A(A[2]), .B(B[595]), .Z(n9687) );
  NANDN U10571 ( .A(n9706), .B(n9707), .Z(n9684) );
  AND U10572 ( .A(A[0]), .B(B[596]), .Z(n9707) );
  XOR U10573 ( .A(n9689), .B(n9708), .Z(n9686) );
  NAND U10574 ( .A(A[0]), .B(B[597]), .Z(n9708) );
  NAND U10575 ( .A(B[596]), .B(A[1]), .Z(n9689) );
  NAND U10576 ( .A(n9709), .B(n9710), .Z(n929) );
  NANDN U10577 ( .A(n9711), .B(n9712), .Z(n9710) );
  OR U10578 ( .A(n9713), .B(n9714), .Z(n9712) );
  NAND U10579 ( .A(n9714), .B(n9713), .Z(n9709) );
  XOR U10580 ( .A(n931), .B(n930), .Z(\A1[594] ) );
  XOR U10581 ( .A(n9714), .B(n9715), .Z(n930) );
  XNOR U10582 ( .A(n9713), .B(n9711), .Z(n9715) );
  AND U10583 ( .A(n9716), .B(n9717), .Z(n9711) );
  NANDN U10584 ( .A(n9718), .B(n9719), .Z(n9717) );
  NANDN U10585 ( .A(n9720), .B(n9721), .Z(n9719) );
  AND U10586 ( .A(B[593]), .B(A[3]), .Z(n9713) );
  XNOR U10587 ( .A(n9703), .B(n9722), .Z(n9714) );
  XNOR U10588 ( .A(n9701), .B(n9704), .Z(n9722) );
  NAND U10589 ( .A(A[2]), .B(B[594]), .Z(n9704) );
  NANDN U10590 ( .A(n9723), .B(n9724), .Z(n9701) );
  AND U10591 ( .A(A[0]), .B(B[595]), .Z(n9724) );
  XOR U10592 ( .A(n9706), .B(n9725), .Z(n9703) );
  NAND U10593 ( .A(A[0]), .B(B[596]), .Z(n9725) );
  NAND U10594 ( .A(B[595]), .B(A[1]), .Z(n9706) );
  NAND U10595 ( .A(n9726), .B(n9727), .Z(n931) );
  NANDN U10596 ( .A(n9728), .B(n9729), .Z(n9727) );
  OR U10597 ( .A(n9730), .B(n9731), .Z(n9729) );
  NAND U10598 ( .A(n9731), .B(n9730), .Z(n9726) );
  XOR U10599 ( .A(n933), .B(n932), .Z(\A1[593] ) );
  XOR U10600 ( .A(n9731), .B(n9732), .Z(n932) );
  XNOR U10601 ( .A(n9730), .B(n9728), .Z(n9732) );
  AND U10602 ( .A(n9733), .B(n9734), .Z(n9728) );
  NANDN U10603 ( .A(n9735), .B(n9736), .Z(n9734) );
  NANDN U10604 ( .A(n9737), .B(n9738), .Z(n9736) );
  AND U10605 ( .A(B[592]), .B(A[3]), .Z(n9730) );
  XNOR U10606 ( .A(n9720), .B(n9739), .Z(n9731) );
  XNOR U10607 ( .A(n9718), .B(n9721), .Z(n9739) );
  NAND U10608 ( .A(A[2]), .B(B[593]), .Z(n9721) );
  NANDN U10609 ( .A(n9740), .B(n9741), .Z(n9718) );
  AND U10610 ( .A(A[0]), .B(B[594]), .Z(n9741) );
  XOR U10611 ( .A(n9723), .B(n9742), .Z(n9720) );
  NAND U10612 ( .A(A[0]), .B(B[595]), .Z(n9742) );
  NAND U10613 ( .A(B[594]), .B(A[1]), .Z(n9723) );
  NAND U10614 ( .A(n9743), .B(n9744), .Z(n933) );
  NANDN U10615 ( .A(n9745), .B(n9746), .Z(n9744) );
  OR U10616 ( .A(n9747), .B(n9748), .Z(n9746) );
  NAND U10617 ( .A(n9748), .B(n9747), .Z(n9743) );
  XOR U10618 ( .A(n935), .B(n934), .Z(\A1[592] ) );
  XOR U10619 ( .A(n9748), .B(n9749), .Z(n934) );
  XNOR U10620 ( .A(n9747), .B(n9745), .Z(n9749) );
  AND U10621 ( .A(n9750), .B(n9751), .Z(n9745) );
  NANDN U10622 ( .A(n9752), .B(n9753), .Z(n9751) );
  NANDN U10623 ( .A(n9754), .B(n9755), .Z(n9753) );
  AND U10624 ( .A(B[591]), .B(A[3]), .Z(n9747) );
  XNOR U10625 ( .A(n9737), .B(n9756), .Z(n9748) );
  XNOR U10626 ( .A(n9735), .B(n9738), .Z(n9756) );
  NAND U10627 ( .A(A[2]), .B(B[592]), .Z(n9738) );
  NANDN U10628 ( .A(n9757), .B(n9758), .Z(n9735) );
  AND U10629 ( .A(A[0]), .B(B[593]), .Z(n9758) );
  XOR U10630 ( .A(n9740), .B(n9759), .Z(n9737) );
  NAND U10631 ( .A(A[0]), .B(B[594]), .Z(n9759) );
  NAND U10632 ( .A(B[593]), .B(A[1]), .Z(n9740) );
  NAND U10633 ( .A(n9760), .B(n9761), .Z(n935) );
  NANDN U10634 ( .A(n9762), .B(n9763), .Z(n9761) );
  OR U10635 ( .A(n9764), .B(n9765), .Z(n9763) );
  NAND U10636 ( .A(n9765), .B(n9764), .Z(n9760) );
  XOR U10637 ( .A(n937), .B(n936), .Z(\A1[591] ) );
  XOR U10638 ( .A(n9765), .B(n9766), .Z(n936) );
  XNOR U10639 ( .A(n9764), .B(n9762), .Z(n9766) );
  AND U10640 ( .A(n9767), .B(n9768), .Z(n9762) );
  NANDN U10641 ( .A(n9769), .B(n9770), .Z(n9768) );
  NANDN U10642 ( .A(n9771), .B(n9772), .Z(n9770) );
  AND U10643 ( .A(B[590]), .B(A[3]), .Z(n9764) );
  XNOR U10644 ( .A(n9754), .B(n9773), .Z(n9765) );
  XNOR U10645 ( .A(n9752), .B(n9755), .Z(n9773) );
  NAND U10646 ( .A(A[2]), .B(B[591]), .Z(n9755) );
  NANDN U10647 ( .A(n9774), .B(n9775), .Z(n9752) );
  AND U10648 ( .A(A[0]), .B(B[592]), .Z(n9775) );
  XOR U10649 ( .A(n9757), .B(n9776), .Z(n9754) );
  NAND U10650 ( .A(A[0]), .B(B[593]), .Z(n9776) );
  NAND U10651 ( .A(B[592]), .B(A[1]), .Z(n9757) );
  NAND U10652 ( .A(n9777), .B(n9778), .Z(n937) );
  NANDN U10653 ( .A(n9779), .B(n9780), .Z(n9778) );
  OR U10654 ( .A(n9781), .B(n9782), .Z(n9780) );
  NAND U10655 ( .A(n9782), .B(n9781), .Z(n9777) );
  XOR U10656 ( .A(n939), .B(n938), .Z(\A1[590] ) );
  XOR U10657 ( .A(n9782), .B(n9783), .Z(n938) );
  XNOR U10658 ( .A(n9781), .B(n9779), .Z(n9783) );
  AND U10659 ( .A(n9784), .B(n9785), .Z(n9779) );
  NANDN U10660 ( .A(n9786), .B(n9787), .Z(n9785) );
  NANDN U10661 ( .A(n9788), .B(n9789), .Z(n9787) );
  AND U10662 ( .A(B[589]), .B(A[3]), .Z(n9781) );
  XNOR U10663 ( .A(n9771), .B(n9790), .Z(n9782) );
  XNOR U10664 ( .A(n9769), .B(n9772), .Z(n9790) );
  NAND U10665 ( .A(A[2]), .B(B[590]), .Z(n9772) );
  NANDN U10666 ( .A(n9791), .B(n9792), .Z(n9769) );
  AND U10667 ( .A(A[0]), .B(B[591]), .Z(n9792) );
  XOR U10668 ( .A(n9774), .B(n9793), .Z(n9771) );
  NAND U10669 ( .A(A[0]), .B(B[592]), .Z(n9793) );
  NAND U10670 ( .A(B[591]), .B(A[1]), .Z(n9774) );
  NAND U10671 ( .A(n9794), .B(n9795), .Z(n939) );
  NANDN U10672 ( .A(n9796), .B(n9797), .Z(n9795) );
  OR U10673 ( .A(n9798), .B(n9799), .Z(n9797) );
  NAND U10674 ( .A(n9799), .B(n9798), .Z(n9794) );
  XOR U10675 ( .A(n921), .B(n920), .Z(\A1[58] ) );
  XOR U10676 ( .A(n9629), .B(n9800), .Z(n920) );
  XNOR U10677 ( .A(n9628), .B(n9626), .Z(n9800) );
  AND U10678 ( .A(n9801), .B(n9802), .Z(n9626) );
  NANDN U10679 ( .A(n9803), .B(n9804), .Z(n9802) );
  NANDN U10680 ( .A(n9805), .B(n9806), .Z(n9804) );
  AND U10681 ( .A(B[57]), .B(A[3]), .Z(n9628) );
  XNOR U10682 ( .A(n9618), .B(n9807), .Z(n9629) );
  XNOR U10683 ( .A(n9616), .B(n9619), .Z(n9807) );
  NAND U10684 ( .A(A[2]), .B(B[58]), .Z(n9619) );
  NANDN U10685 ( .A(n9808), .B(n9809), .Z(n9616) );
  AND U10686 ( .A(A[0]), .B(B[59]), .Z(n9809) );
  XOR U10687 ( .A(n9621), .B(n9810), .Z(n9618) );
  NAND U10688 ( .A(A[0]), .B(B[60]), .Z(n9810) );
  NAND U10689 ( .A(B[59]), .B(A[1]), .Z(n9621) );
  NAND U10690 ( .A(n9811), .B(n9812), .Z(n921) );
  NANDN U10691 ( .A(n9813), .B(n9814), .Z(n9812) );
  OR U10692 ( .A(n9815), .B(n9816), .Z(n9814) );
  NAND U10693 ( .A(n9816), .B(n9815), .Z(n9811) );
  XOR U10694 ( .A(n941), .B(n940), .Z(\A1[589] ) );
  XOR U10695 ( .A(n9799), .B(n9817), .Z(n940) );
  XNOR U10696 ( .A(n9798), .B(n9796), .Z(n9817) );
  AND U10697 ( .A(n9818), .B(n9819), .Z(n9796) );
  NANDN U10698 ( .A(n9820), .B(n9821), .Z(n9819) );
  NANDN U10699 ( .A(n9822), .B(n9823), .Z(n9821) );
  AND U10700 ( .A(B[588]), .B(A[3]), .Z(n9798) );
  XNOR U10701 ( .A(n9788), .B(n9824), .Z(n9799) );
  XNOR U10702 ( .A(n9786), .B(n9789), .Z(n9824) );
  NAND U10703 ( .A(A[2]), .B(B[589]), .Z(n9789) );
  NANDN U10704 ( .A(n9825), .B(n9826), .Z(n9786) );
  AND U10705 ( .A(A[0]), .B(B[590]), .Z(n9826) );
  XOR U10706 ( .A(n9791), .B(n9827), .Z(n9788) );
  NAND U10707 ( .A(A[0]), .B(B[591]), .Z(n9827) );
  NAND U10708 ( .A(B[590]), .B(A[1]), .Z(n9791) );
  NAND U10709 ( .A(n9828), .B(n9829), .Z(n941) );
  NANDN U10710 ( .A(n9830), .B(n9831), .Z(n9829) );
  OR U10711 ( .A(n9832), .B(n9833), .Z(n9831) );
  NAND U10712 ( .A(n9833), .B(n9832), .Z(n9828) );
  XOR U10713 ( .A(n945), .B(n944), .Z(\A1[588] ) );
  XOR U10714 ( .A(n9833), .B(n9834), .Z(n944) );
  XNOR U10715 ( .A(n9832), .B(n9830), .Z(n9834) );
  AND U10716 ( .A(n9835), .B(n9836), .Z(n9830) );
  NANDN U10717 ( .A(n9837), .B(n9838), .Z(n9836) );
  NANDN U10718 ( .A(n9839), .B(n9840), .Z(n9838) );
  AND U10719 ( .A(B[587]), .B(A[3]), .Z(n9832) );
  XNOR U10720 ( .A(n9822), .B(n9841), .Z(n9833) );
  XNOR U10721 ( .A(n9820), .B(n9823), .Z(n9841) );
  NAND U10722 ( .A(A[2]), .B(B[588]), .Z(n9823) );
  NANDN U10723 ( .A(n9842), .B(n9843), .Z(n9820) );
  AND U10724 ( .A(A[0]), .B(B[589]), .Z(n9843) );
  XOR U10725 ( .A(n9825), .B(n9844), .Z(n9822) );
  NAND U10726 ( .A(A[0]), .B(B[590]), .Z(n9844) );
  NAND U10727 ( .A(B[589]), .B(A[1]), .Z(n9825) );
  NAND U10728 ( .A(n9845), .B(n9846), .Z(n945) );
  NANDN U10729 ( .A(n9847), .B(n9848), .Z(n9846) );
  OR U10730 ( .A(n9849), .B(n9850), .Z(n9848) );
  NAND U10731 ( .A(n9850), .B(n9849), .Z(n9845) );
  XOR U10732 ( .A(n947), .B(n946), .Z(\A1[587] ) );
  XOR U10733 ( .A(n9850), .B(n9851), .Z(n946) );
  XNOR U10734 ( .A(n9849), .B(n9847), .Z(n9851) );
  AND U10735 ( .A(n9852), .B(n9853), .Z(n9847) );
  NANDN U10736 ( .A(n9854), .B(n9855), .Z(n9853) );
  NANDN U10737 ( .A(n9856), .B(n9857), .Z(n9855) );
  AND U10738 ( .A(B[586]), .B(A[3]), .Z(n9849) );
  XNOR U10739 ( .A(n9839), .B(n9858), .Z(n9850) );
  XNOR U10740 ( .A(n9837), .B(n9840), .Z(n9858) );
  NAND U10741 ( .A(A[2]), .B(B[587]), .Z(n9840) );
  NANDN U10742 ( .A(n9859), .B(n9860), .Z(n9837) );
  AND U10743 ( .A(A[0]), .B(B[588]), .Z(n9860) );
  XOR U10744 ( .A(n9842), .B(n9861), .Z(n9839) );
  NAND U10745 ( .A(A[0]), .B(B[589]), .Z(n9861) );
  NAND U10746 ( .A(B[588]), .B(A[1]), .Z(n9842) );
  NAND U10747 ( .A(n9862), .B(n9863), .Z(n947) );
  NANDN U10748 ( .A(n9864), .B(n9865), .Z(n9863) );
  OR U10749 ( .A(n9866), .B(n9867), .Z(n9865) );
  NAND U10750 ( .A(n9867), .B(n9866), .Z(n9862) );
  XOR U10751 ( .A(n949), .B(n948), .Z(\A1[586] ) );
  XOR U10752 ( .A(n9867), .B(n9868), .Z(n948) );
  XNOR U10753 ( .A(n9866), .B(n9864), .Z(n9868) );
  AND U10754 ( .A(n9869), .B(n9870), .Z(n9864) );
  NANDN U10755 ( .A(n9871), .B(n9872), .Z(n9870) );
  NANDN U10756 ( .A(n9873), .B(n9874), .Z(n9872) );
  AND U10757 ( .A(B[585]), .B(A[3]), .Z(n9866) );
  XNOR U10758 ( .A(n9856), .B(n9875), .Z(n9867) );
  XNOR U10759 ( .A(n9854), .B(n9857), .Z(n9875) );
  NAND U10760 ( .A(A[2]), .B(B[586]), .Z(n9857) );
  NANDN U10761 ( .A(n9876), .B(n9877), .Z(n9854) );
  AND U10762 ( .A(A[0]), .B(B[587]), .Z(n9877) );
  XOR U10763 ( .A(n9859), .B(n9878), .Z(n9856) );
  NAND U10764 ( .A(A[0]), .B(B[588]), .Z(n9878) );
  NAND U10765 ( .A(B[587]), .B(A[1]), .Z(n9859) );
  NAND U10766 ( .A(n9879), .B(n9880), .Z(n949) );
  NANDN U10767 ( .A(n9881), .B(n9882), .Z(n9880) );
  OR U10768 ( .A(n9883), .B(n9884), .Z(n9882) );
  NAND U10769 ( .A(n9884), .B(n9883), .Z(n9879) );
  XOR U10770 ( .A(n951), .B(n950), .Z(\A1[585] ) );
  XOR U10771 ( .A(n9884), .B(n9885), .Z(n950) );
  XNOR U10772 ( .A(n9883), .B(n9881), .Z(n9885) );
  AND U10773 ( .A(n9886), .B(n9887), .Z(n9881) );
  NANDN U10774 ( .A(n9888), .B(n9889), .Z(n9887) );
  NANDN U10775 ( .A(n9890), .B(n9891), .Z(n9889) );
  AND U10776 ( .A(B[584]), .B(A[3]), .Z(n9883) );
  XNOR U10777 ( .A(n9873), .B(n9892), .Z(n9884) );
  XNOR U10778 ( .A(n9871), .B(n9874), .Z(n9892) );
  NAND U10779 ( .A(A[2]), .B(B[585]), .Z(n9874) );
  NANDN U10780 ( .A(n9893), .B(n9894), .Z(n9871) );
  AND U10781 ( .A(A[0]), .B(B[586]), .Z(n9894) );
  XOR U10782 ( .A(n9876), .B(n9895), .Z(n9873) );
  NAND U10783 ( .A(A[0]), .B(B[587]), .Z(n9895) );
  NAND U10784 ( .A(B[586]), .B(A[1]), .Z(n9876) );
  NAND U10785 ( .A(n9896), .B(n9897), .Z(n951) );
  NANDN U10786 ( .A(n9898), .B(n9899), .Z(n9897) );
  OR U10787 ( .A(n9900), .B(n9901), .Z(n9899) );
  NAND U10788 ( .A(n9901), .B(n9900), .Z(n9896) );
  XOR U10789 ( .A(n953), .B(n952), .Z(\A1[584] ) );
  XOR U10790 ( .A(n9901), .B(n9902), .Z(n952) );
  XNOR U10791 ( .A(n9900), .B(n9898), .Z(n9902) );
  AND U10792 ( .A(n9903), .B(n9904), .Z(n9898) );
  NANDN U10793 ( .A(n9905), .B(n9906), .Z(n9904) );
  NANDN U10794 ( .A(n9907), .B(n9908), .Z(n9906) );
  AND U10795 ( .A(B[583]), .B(A[3]), .Z(n9900) );
  XNOR U10796 ( .A(n9890), .B(n9909), .Z(n9901) );
  XNOR U10797 ( .A(n9888), .B(n9891), .Z(n9909) );
  NAND U10798 ( .A(A[2]), .B(B[584]), .Z(n9891) );
  NANDN U10799 ( .A(n9910), .B(n9911), .Z(n9888) );
  AND U10800 ( .A(A[0]), .B(B[585]), .Z(n9911) );
  XOR U10801 ( .A(n9893), .B(n9912), .Z(n9890) );
  NAND U10802 ( .A(A[0]), .B(B[586]), .Z(n9912) );
  NAND U10803 ( .A(B[585]), .B(A[1]), .Z(n9893) );
  NAND U10804 ( .A(n9913), .B(n9914), .Z(n953) );
  NANDN U10805 ( .A(n9915), .B(n9916), .Z(n9914) );
  OR U10806 ( .A(n9917), .B(n9918), .Z(n9916) );
  NAND U10807 ( .A(n9918), .B(n9917), .Z(n9913) );
  XOR U10808 ( .A(n955), .B(n954), .Z(\A1[583] ) );
  XOR U10809 ( .A(n9918), .B(n9919), .Z(n954) );
  XNOR U10810 ( .A(n9917), .B(n9915), .Z(n9919) );
  AND U10811 ( .A(n9920), .B(n9921), .Z(n9915) );
  NANDN U10812 ( .A(n9922), .B(n9923), .Z(n9921) );
  NANDN U10813 ( .A(n9924), .B(n9925), .Z(n9923) );
  AND U10814 ( .A(B[582]), .B(A[3]), .Z(n9917) );
  XNOR U10815 ( .A(n9907), .B(n9926), .Z(n9918) );
  XNOR U10816 ( .A(n9905), .B(n9908), .Z(n9926) );
  NAND U10817 ( .A(A[2]), .B(B[583]), .Z(n9908) );
  NANDN U10818 ( .A(n9927), .B(n9928), .Z(n9905) );
  AND U10819 ( .A(A[0]), .B(B[584]), .Z(n9928) );
  XOR U10820 ( .A(n9910), .B(n9929), .Z(n9907) );
  NAND U10821 ( .A(A[0]), .B(B[585]), .Z(n9929) );
  NAND U10822 ( .A(B[584]), .B(A[1]), .Z(n9910) );
  NAND U10823 ( .A(n9930), .B(n9931), .Z(n955) );
  NANDN U10824 ( .A(n9932), .B(n9933), .Z(n9931) );
  OR U10825 ( .A(n9934), .B(n9935), .Z(n9933) );
  NAND U10826 ( .A(n9935), .B(n9934), .Z(n9930) );
  XOR U10827 ( .A(n957), .B(n956), .Z(\A1[582] ) );
  XOR U10828 ( .A(n9935), .B(n9936), .Z(n956) );
  XNOR U10829 ( .A(n9934), .B(n9932), .Z(n9936) );
  AND U10830 ( .A(n9937), .B(n9938), .Z(n9932) );
  NANDN U10831 ( .A(n9939), .B(n9940), .Z(n9938) );
  NANDN U10832 ( .A(n9941), .B(n9942), .Z(n9940) );
  AND U10833 ( .A(B[581]), .B(A[3]), .Z(n9934) );
  XNOR U10834 ( .A(n9924), .B(n9943), .Z(n9935) );
  XNOR U10835 ( .A(n9922), .B(n9925), .Z(n9943) );
  NAND U10836 ( .A(A[2]), .B(B[582]), .Z(n9925) );
  NANDN U10837 ( .A(n9944), .B(n9945), .Z(n9922) );
  AND U10838 ( .A(A[0]), .B(B[583]), .Z(n9945) );
  XOR U10839 ( .A(n9927), .B(n9946), .Z(n9924) );
  NAND U10840 ( .A(A[0]), .B(B[584]), .Z(n9946) );
  NAND U10841 ( .A(B[583]), .B(A[1]), .Z(n9927) );
  NAND U10842 ( .A(n9947), .B(n9948), .Z(n957) );
  NANDN U10843 ( .A(n9949), .B(n9950), .Z(n9948) );
  OR U10844 ( .A(n9951), .B(n9952), .Z(n9950) );
  NAND U10845 ( .A(n9952), .B(n9951), .Z(n9947) );
  XOR U10846 ( .A(n959), .B(n958), .Z(\A1[581] ) );
  XOR U10847 ( .A(n9952), .B(n9953), .Z(n958) );
  XNOR U10848 ( .A(n9951), .B(n9949), .Z(n9953) );
  AND U10849 ( .A(n9954), .B(n9955), .Z(n9949) );
  NANDN U10850 ( .A(n9956), .B(n9957), .Z(n9955) );
  NANDN U10851 ( .A(n9958), .B(n9959), .Z(n9957) );
  AND U10852 ( .A(B[580]), .B(A[3]), .Z(n9951) );
  XNOR U10853 ( .A(n9941), .B(n9960), .Z(n9952) );
  XNOR U10854 ( .A(n9939), .B(n9942), .Z(n9960) );
  NAND U10855 ( .A(A[2]), .B(B[581]), .Z(n9942) );
  NANDN U10856 ( .A(n9961), .B(n9962), .Z(n9939) );
  AND U10857 ( .A(A[0]), .B(B[582]), .Z(n9962) );
  XOR U10858 ( .A(n9944), .B(n9963), .Z(n9941) );
  NAND U10859 ( .A(A[0]), .B(B[583]), .Z(n9963) );
  NAND U10860 ( .A(B[582]), .B(A[1]), .Z(n9944) );
  NAND U10861 ( .A(n9964), .B(n9965), .Z(n959) );
  NANDN U10862 ( .A(n9966), .B(n9967), .Z(n9965) );
  OR U10863 ( .A(n9968), .B(n9969), .Z(n9967) );
  NAND U10864 ( .A(n9969), .B(n9968), .Z(n9964) );
  XOR U10865 ( .A(n961), .B(n960), .Z(\A1[580] ) );
  XOR U10866 ( .A(n9969), .B(n9970), .Z(n960) );
  XNOR U10867 ( .A(n9968), .B(n9966), .Z(n9970) );
  AND U10868 ( .A(n9971), .B(n9972), .Z(n9966) );
  NANDN U10869 ( .A(n9973), .B(n9974), .Z(n9972) );
  NANDN U10870 ( .A(n9975), .B(n9976), .Z(n9974) );
  AND U10871 ( .A(B[579]), .B(A[3]), .Z(n9968) );
  XNOR U10872 ( .A(n9958), .B(n9977), .Z(n9969) );
  XNOR U10873 ( .A(n9956), .B(n9959), .Z(n9977) );
  NAND U10874 ( .A(A[2]), .B(B[580]), .Z(n9959) );
  NANDN U10875 ( .A(n9978), .B(n9979), .Z(n9956) );
  AND U10876 ( .A(A[0]), .B(B[581]), .Z(n9979) );
  XOR U10877 ( .A(n9961), .B(n9980), .Z(n9958) );
  NAND U10878 ( .A(A[0]), .B(B[582]), .Z(n9980) );
  NAND U10879 ( .A(B[581]), .B(A[1]), .Z(n9961) );
  NAND U10880 ( .A(n9981), .B(n9982), .Z(n961) );
  NANDN U10881 ( .A(n9983), .B(n9984), .Z(n9982) );
  OR U10882 ( .A(n9985), .B(n9986), .Z(n9984) );
  NAND U10883 ( .A(n9986), .B(n9985), .Z(n9981) );
  XOR U10884 ( .A(n943), .B(n942), .Z(\A1[57] ) );
  XOR U10885 ( .A(n9816), .B(n9987), .Z(n942) );
  XNOR U10886 ( .A(n9815), .B(n9813), .Z(n9987) );
  AND U10887 ( .A(n9988), .B(n9989), .Z(n9813) );
  NANDN U10888 ( .A(n9990), .B(n9991), .Z(n9989) );
  NANDN U10889 ( .A(n9992), .B(n9993), .Z(n9991) );
  AND U10890 ( .A(B[56]), .B(A[3]), .Z(n9815) );
  XNOR U10891 ( .A(n9805), .B(n9994), .Z(n9816) );
  XNOR U10892 ( .A(n9803), .B(n9806), .Z(n9994) );
  NAND U10893 ( .A(A[2]), .B(B[57]), .Z(n9806) );
  NANDN U10894 ( .A(n9995), .B(n9996), .Z(n9803) );
  AND U10895 ( .A(A[0]), .B(B[58]), .Z(n9996) );
  XOR U10896 ( .A(n9808), .B(n9997), .Z(n9805) );
  NAND U10897 ( .A(A[0]), .B(B[59]), .Z(n9997) );
  NAND U10898 ( .A(B[58]), .B(A[1]), .Z(n9808) );
  NAND U10899 ( .A(n9998), .B(n9999), .Z(n943) );
  NANDN U10900 ( .A(n10000), .B(n10001), .Z(n9999) );
  OR U10901 ( .A(n10002), .B(n10003), .Z(n10001) );
  NAND U10902 ( .A(n10003), .B(n10002), .Z(n9998) );
  XOR U10903 ( .A(n963), .B(n962), .Z(\A1[579] ) );
  XOR U10904 ( .A(n9986), .B(n10004), .Z(n962) );
  XNOR U10905 ( .A(n9985), .B(n9983), .Z(n10004) );
  AND U10906 ( .A(n10005), .B(n10006), .Z(n9983) );
  NANDN U10907 ( .A(n10007), .B(n10008), .Z(n10006) );
  NANDN U10908 ( .A(n10009), .B(n10010), .Z(n10008) );
  AND U10909 ( .A(B[578]), .B(A[3]), .Z(n9985) );
  XNOR U10910 ( .A(n9975), .B(n10011), .Z(n9986) );
  XNOR U10911 ( .A(n9973), .B(n9976), .Z(n10011) );
  NAND U10912 ( .A(A[2]), .B(B[579]), .Z(n9976) );
  NANDN U10913 ( .A(n10012), .B(n10013), .Z(n9973) );
  AND U10914 ( .A(A[0]), .B(B[580]), .Z(n10013) );
  XOR U10915 ( .A(n9978), .B(n10014), .Z(n9975) );
  NAND U10916 ( .A(A[0]), .B(B[581]), .Z(n10014) );
  NAND U10917 ( .A(B[580]), .B(A[1]), .Z(n9978) );
  NAND U10918 ( .A(n10015), .B(n10016), .Z(n963) );
  NANDN U10919 ( .A(n10017), .B(n10018), .Z(n10016) );
  OR U10920 ( .A(n10019), .B(n10020), .Z(n10018) );
  NAND U10921 ( .A(n10020), .B(n10019), .Z(n10015) );
  XOR U10922 ( .A(n967), .B(n966), .Z(\A1[578] ) );
  XOR U10923 ( .A(n10020), .B(n10021), .Z(n966) );
  XNOR U10924 ( .A(n10019), .B(n10017), .Z(n10021) );
  AND U10925 ( .A(n10022), .B(n10023), .Z(n10017) );
  NANDN U10926 ( .A(n10024), .B(n10025), .Z(n10023) );
  NANDN U10927 ( .A(n10026), .B(n10027), .Z(n10025) );
  AND U10928 ( .A(B[577]), .B(A[3]), .Z(n10019) );
  XNOR U10929 ( .A(n10009), .B(n10028), .Z(n10020) );
  XNOR U10930 ( .A(n10007), .B(n10010), .Z(n10028) );
  NAND U10931 ( .A(A[2]), .B(B[578]), .Z(n10010) );
  NANDN U10932 ( .A(n10029), .B(n10030), .Z(n10007) );
  AND U10933 ( .A(A[0]), .B(B[579]), .Z(n10030) );
  XOR U10934 ( .A(n10012), .B(n10031), .Z(n10009) );
  NAND U10935 ( .A(A[0]), .B(B[580]), .Z(n10031) );
  NAND U10936 ( .A(B[579]), .B(A[1]), .Z(n10012) );
  NAND U10937 ( .A(n10032), .B(n10033), .Z(n967) );
  NANDN U10938 ( .A(n10034), .B(n10035), .Z(n10033) );
  OR U10939 ( .A(n10036), .B(n10037), .Z(n10035) );
  NAND U10940 ( .A(n10037), .B(n10036), .Z(n10032) );
  XOR U10941 ( .A(n969), .B(n968), .Z(\A1[577] ) );
  XOR U10942 ( .A(n10037), .B(n10038), .Z(n968) );
  XNOR U10943 ( .A(n10036), .B(n10034), .Z(n10038) );
  AND U10944 ( .A(n10039), .B(n10040), .Z(n10034) );
  NANDN U10945 ( .A(n10041), .B(n10042), .Z(n10040) );
  NANDN U10946 ( .A(n10043), .B(n10044), .Z(n10042) );
  AND U10947 ( .A(B[576]), .B(A[3]), .Z(n10036) );
  XNOR U10948 ( .A(n10026), .B(n10045), .Z(n10037) );
  XNOR U10949 ( .A(n10024), .B(n10027), .Z(n10045) );
  NAND U10950 ( .A(A[2]), .B(B[577]), .Z(n10027) );
  NANDN U10951 ( .A(n10046), .B(n10047), .Z(n10024) );
  AND U10952 ( .A(A[0]), .B(B[578]), .Z(n10047) );
  XOR U10953 ( .A(n10029), .B(n10048), .Z(n10026) );
  NAND U10954 ( .A(A[0]), .B(B[579]), .Z(n10048) );
  NAND U10955 ( .A(B[578]), .B(A[1]), .Z(n10029) );
  NAND U10956 ( .A(n10049), .B(n10050), .Z(n969) );
  NANDN U10957 ( .A(n10051), .B(n10052), .Z(n10050) );
  OR U10958 ( .A(n10053), .B(n10054), .Z(n10052) );
  NAND U10959 ( .A(n10054), .B(n10053), .Z(n10049) );
  XOR U10960 ( .A(n971), .B(n970), .Z(\A1[576] ) );
  XOR U10961 ( .A(n10054), .B(n10055), .Z(n970) );
  XNOR U10962 ( .A(n10053), .B(n10051), .Z(n10055) );
  AND U10963 ( .A(n10056), .B(n10057), .Z(n10051) );
  NANDN U10964 ( .A(n10058), .B(n10059), .Z(n10057) );
  NANDN U10965 ( .A(n10060), .B(n10061), .Z(n10059) );
  AND U10966 ( .A(B[575]), .B(A[3]), .Z(n10053) );
  XNOR U10967 ( .A(n10043), .B(n10062), .Z(n10054) );
  XNOR U10968 ( .A(n10041), .B(n10044), .Z(n10062) );
  NAND U10969 ( .A(A[2]), .B(B[576]), .Z(n10044) );
  NANDN U10970 ( .A(n10063), .B(n10064), .Z(n10041) );
  AND U10971 ( .A(A[0]), .B(B[577]), .Z(n10064) );
  XOR U10972 ( .A(n10046), .B(n10065), .Z(n10043) );
  NAND U10973 ( .A(A[0]), .B(B[578]), .Z(n10065) );
  NAND U10974 ( .A(B[577]), .B(A[1]), .Z(n10046) );
  NAND U10975 ( .A(n10066), .B(n10067), .Z(n971) );
  NANDN U10976 ( .A(n10068), .B(n10069), .Z(n10067) );
  OR U10977 ( .A(n10070), .B(n10071), .Z(n10069) );
  NAND U10978 ( .A(n10071), .B(n10070), .Z(n10066) );
  XOR U10979 ( .A(n973), .B(n972), .Z(\A1[575] ) );
  XOR U10980 ( .A(n10071), .B(n10072), .Z(n972) );
  XNOR U10981 ( .A(n10070), .B(n10068), .Z(n10072) );
  AND U10982 ( .A(n10073), .B(n10074), .Z(n10068) );
  NANDN U10983 ( .A(n10075), .B(n10076), .Z(n10074) );
  NANDN U10984 ( .A(n10077), .B(n10078), .Z(n10076) );
  AND U10985 ( .A(B[574]), .B(A[3]), .Z(n10070) );
  XNOR U10986 ( .A(n10060), .B(n10079), .Z(n10071) );
  XNOR U10987 ( .A(n10058), .B(n10061), .Z(n10079) );
  NAND U10988 ( .A(A[2]), .B(B[575]), .Z(n10061) );
  NANDN U10989 ( .A(n10080), .B(n10081), .Z(n10058) );
  AND U10990 ( .A(A[0]), .B(B[576]), .Z(n10081) );
  XOR U10991 ( .A(n10063), .B(n10082), .Z(n10060) );
  NAND U10992 ( .A(A[0]), .B(B[577]), .Z(n10082) );
  NAND U10993 ( .A(B[576]), .B(A[1]), .Z(n10063) );
  NAND U10994 ( .A(n10083), .B(n10084), .Z(n973) );
  NANDN U10995 ( .A(n10085), .B(n10086), .Z(n10084) );
  OR U10996 ( .A(n10087), .B(n10088), .Z(n10086) );
  NAND U10997 ( .A(n10088), .B(n10087), .Z(n10083) );
  XOR U10998 ( .A(n975), .B(n974), .Z(\A1[574] ) );
  XOR U10999 ( .A(n10088), .B(n10089), .Z(n974) );
  XNOR U11000 ( .A(n10087), .B(n10085), .Z(n10089) );
  AND U11001 ( .A(n10090), .B(n10091), .Z(n10085) );
  NANDN U11002 ( .A(n10092), .B(n10093), .Z(n10091) );
  NANDN U11003 ( .A(n10094), .B(n10095), .Z(n10093) );
  AND U11004 ( .A(B[573]), .B(A[3]), .Z(n10087) );
  XNOR U11005 ( .A(n10077), .B(n10096), .Z(n10088) );
  XNOR U11006 ( .A(n10075), .B(n10078), .Z(n10096) );
  NAND U11007 ( .A(A[2]), .B(B[574]), .Z(n10078) );
  NANDN U11008 ( .A(n10097), .B(n10098), .Z(n10075) );
  AND U11009 ( .A(A[0]), .B(B[575]), .Z(n10098) );
  XOR U11010 ( .A(n10080), .B(n10099), .Z(n10077) );
  NAND U11011 ( .A(A[0]), .B(B[576]), .Z(n10099) );
  NAND U11012 ( .A(B[575]), .B(A[1]), .Z(n10080) );
  NAND U11013 ( .A(n10100), .B(n10101), .Z(n975) );
  NANDN U11014 ( .A(n10102), .B(n10103), .Z(n10101) );
  OR U11015 ( .A(n10104), .B(n10105), .Z(n10103) );
  NAND U11016 ( .A(n10105), .B(n10104), .Z(n10100) );
  XOR U11017 ( .A(n977), .B(n976), .Z(\A1[573] ) );
  XOR U11018 ( .A(n10105), .B(n10106), .Z(n976) );
  XNOR U11019 ( .A(n10104), .B(n10102), .Z(n10106) );
  AND U11020 ( .A(n10107), .B(n10108), .Z(n10102) );
  NANDN U11021 ( .A(n10109), .B(n10110), .Z(n10108) );
  NANDN U11022 ( .A(n10111), .B(n10112), .Z(n10110) );
  AND U11023 ( .A(B[572]), .B(A[3]), .Z(n10104) );
  XNOR U11024 ( .A(n10094), .B(n10113), .Z(n10105) );
  XNOR U11025 ( .A(n10092), .B(n10095), .Z(n10113) );
  NAND U11026 ( .A(A[2]), .B(B[573]), .Z(n10095) );
  NANDN U11027 ( .A(n10114), .B(n10115), .Z(n10092) );
  AND U11028 ( .A(A[0]), .B(B[574]), .Z(n10115) );
  XOR U11029 ( .A(n10097), .B(n10116), .Z(n10094) );
  NAND U11030 ( .A(A[0]), .B(B[575]), .Z(n10116) );
  NAND U11031 ( .A(B[574]), .B(A[1]), .Z(n10097) );
  NAND U11032 ( .A(n10117), .B(n10118), .Z(n977) );
  NANDN U11033 ( .A(n10119), .B(n10120), .Z(n10118) );
  OR U11034 ( .A(n10121), .B(n10122), .Z(n10120) );
  NAND U11035 ( .A(n10122), .B(n10121), .Z(n10117) );
  XOR U11036 ( .A(n979), .B(n978), .Z(\A1[572] ) );
  XOR U11037 ( .A(n10122), .B(n10123), .Z(n978) );
  XNOR U11038 ( .A(n10121), .B(n10119), .Z(n10123) );
  AND U11039 ( .A(n10124), .B(n10125), .Z(n10119) );
  NANDN U11040 ( .A(n10126), .B(n10127), .Z(n10125) );
  NANDN U11041 ( .A(n10128), .B(n10129), .Z(n10127) );
  AND U11042 ( .A(B[571]), .B(A[3]), .Z(n10121) );
  XNOR U11043 ( .A(n10111), .B(n10130), .Z(n10122) );
  XNOR U11044 ( .A(n10109), .B(n10112), .Z(n10130) );
  NAND U11045 ( .A(A[2]), .B(B[572]), .Z(n10112) );
  NANDN U11046 ( .A(n10131), .B(n10132), .Z(n10109) );
  AND U11047 ( .A(A[0]), .B(B[573]), .Z(n10132) );
  XOR U11048 ( .A(n10114), .B(n10133), .Z(n10111) );
  NAND U11049 ( .A(A[0]), .B(B[574]), .Z(n10133) );
  NAND U11050 ( .A(B[573]), .B(A[1]), .Z(n10114) );
  NAND U11051 ( .A(n10134), .B(n10135), .Z(n979) );
  NANDN U11052 ( .A(n10136), .B(n10137), .Z(n10135) );
  OR U11053 ( .A(n10138), .B(n10139), .Z(n10137) );
  NAND U11054 ( .A(n10139), .B(n10138), .Z(n10134) );
  XOR U11055 ( .A(n981), .B(n980), .Z(\A1[571] ) );
  XOR U11056 ( .A(n10139), .B(n10140), .Z(n980) );
  XNOR U11057 ( .A(n10138), .B(n10136), .Z(n10140) );
  AND U11058 ( .A(n10141), .B(n10142), .Z(n10136) );
  NANDN U11059 ( .A(n10143), .B(n10144), .Z(n10142) );
  NANDN U11060 ( .A(n10145), .B(n10146), .Z(n10144) );
  AND U11061 ( .A(B[570]), .B(A[3]), .Z(n10138) );
  XNOR U11062 ( .A(n10128), .B(n10147), .Z(n10139) );
  XNOR U11063 ( .A(n10126), .B(n10129), .Z(n10147) );
  NAND U11064 ( .A(A[2]), .B(B[571]), .Z(n10129) );
  NANDN U11065 ( .A(n10148), .B(n10149), .Z(n10126) );
  AND U11066 ( .A(A[0]), .B(B[572]), .Z(n10149) );
  XOR U11067 ( .A(n10131), .B(n10150), .Z(n10128) );
  NAND U11068 ( .A(A[0]), .B(B[573]), .Z(n10150) );
  NAND U11069 ( .A(B[572]), .B(A[1]), .Z(n10131) );
  NAND U11070 ( .A(n10151), .B(n10152), .Z(n981) );
  NANDN U11071 ( .A(n10153), .B(n10154), .Z(n10152) );
  OR U11072 ( .A(n10155), .B(n10156), .Z(n10154) );
  NAND U11073 ( .A(n10156), .B(n10155), .Z(n10151) );
  XOR U11074 ( .A(n983), .B(n982), .Z(\A1[570] ) );
  XOR U11075 ( .A(n10156), .B(n10157), .Z(n982) );
  XNOR U11076 ( .A(n10155), .B(n10153), .Z(n10157) );
  AND U11077 ( .A(n10158), .B(n10159), .Z(n10153) );
  NANDN U11078 ( .A(n10160), .B(n10161), .Z(n10159) );
  NANDN U11079 ( .A(n10162), .B(n10163), .Z(n10161) );
  AND U11080 ( .A(B[569]), .B(A[3]), .Z(n10155) );
  XNOR U11081 ( .A(n10145), .B(n10164), .Z(n10156) );
  XNOR U11082 ( .A(n10143), .B(n10146), .Z(n10164) );
  NAND U11083 ( .A(A[2]), .B(B[570]), .Z(n10146) );
  NANDN U11084 ( .A(n10165), .B(n10166), .Z(n10143) );
  AND U11085 ( .A(A[0]), .B(B[571]), .Z(n10166) );
  XOR U11086 ( .A(n10148), .B(n10167), .Z(n10145) );
  NAND U11087 ( .A(A[0]), .B(B[572]), .Z(n10167) );
  NAND U11088 ( .A(B[571]), .B(A[1]), .Z(n10148) );
  NAND U11089 ( .A(n10168), .B(n10169), .Z(n983) );
  NANDN U11090 ( .A(n10170), .B(n10171), .Z(n10169) );
  OR U11091 ( .A(n10172), .B(n10173), .Z(n10171) );
  NAND U11092 ( .A(n10173), .B(n10172), .Z(n10168) );
  XOR U11093 ( .A(n965), .B(n964), .Z(\A1[56] ) );
  XOR U11094 ( .A(n10003), .B(n10174), .Z(n964) );
  XNOR U11095 ( .A(n10002), .B(n10000), .Z(n10174) );
  AND U11096 ( .A(n10175), .B(n10176), .Z(n10000) );
  NANDN U11097 ( .A(n10177), .B(n10178), .Z(n10176) );
  NANDN U11098 ( .A(n10179), .B(n10180), .Z(n10178) );
  AND U11099 ( .A(B[55]), .B(A[3]), .Z(n10002) );
  XNOR U11100 ( .A(n9992), .B(n10181), .Z(n10003) );
  XNOR U11101 ( .A(n9990), .B(n9993), .Z(n10181) );
  NAND U11102 ( .A(A[2]), .B(B[56]), .Z(n9993) );
  NANDN U11103 ( .A(n10182), .B(n10183), .Z(n9990) );
  AND U11104 ( .A(A[0]), .B(B[57]), .Z(n10183) );
  XOR U11105 ( .A(n9995), .B(n10184), .Z(n9992) );
  NAND U11106 ( .A(A[0]), .B(B[58]), .Z(n10184) );
  NAND U11107 ( .A(B[57]), .B(A[1]), .Z(n9995) );
  NAND U11108 ( .A(n10185), .B(n10186), .Z(n965) );
  NANDN U11109 ( .A(n10187), .B(n10188), .Z(n10186) );
  OR U11110 ( .A(n10189), .B(n10190), .Z(n10188) );
  NAND U11111 ( .A(n10190), .B(n10189), .Z(n10185) );
  XOR U11112 ( .A(n985), .B(n984), .Z(\A1[569] ) );
  XOR U11113 ( .A(n10173), .B(n10191), .Z(n984) );
  XNOR U11114 ( .A(n10172), .B(n10170), .Z(n10191) );
  AND U11115 ( .A(n10192), .B(n10193), .Z(n10170) );
  NANDN U11116 ( .A(n10194), .B(n10195), .Z(n10193) );
  NANDN U11117 ( .A(n10196), .B(n10197), .Z(n10195) );
  AND U11118 ( .A(B[568]), .B(A[3]), .Z(n10172) );
  XNOR U11119 ( .A(n10162), .B(n10198), .Z(n10173) );
  XNOR U11120 ( .A(n10160), .B(n10163), .Z(n10198) );
  NAND U11121 ( .A(A[2]), .B(B[569]), .Z(n10163) );
  NANDN U11122 ( .A(n10199), .B(n10200), .Z(n10160) );
  AND U11123 ( .A(A[0]), .B(B[570]), .Z(n10200) );
  XOR U11124 ( .A(n10165), .B(n10201), .Z(n10162) );
  NAND U11125 ( .A(A[0]), .B(B[571]), .Z(n10201) );
  NAND U11126 ( .A(B[570]), .B(A[1]), .Z(n10165) );
  NAND U11127 ( .A(n10202), .B(n10203), .Z(n985) );
  NANDN U11128 ( .A(n10204), .B(n10205), .Z(n10203) );
  OR U11129 ( .A(n10206), .B(n10207), .Z(n10205) );
  NAND U11130 ( .A(n10207), .B(n10206), .Z(n10202) );
  XOR U11131 ( .A(n989), .B(n988), .Z(\A1[568] ) );
  XOR U11132 ( .A(n10207), .B(n10208), .Z(n988) );
  XNOR U11133 ( .A(n10206), .B(n10204), .Z(n10208) );
  AND U11134 ( .A(n10209), .B(n10210), .Z(n10204) );
  NANDN U11135 ( .A(n10211), .B(n10212), .Z(n10210) );
  NANDN U11136 ( .A(n10213), .B(n10214), .Z(n10212) );
  AND U11137 ( .A(B[567]), .B(A[3]), .Z(n10206) );
  XNOR U11138 ( .A(n10196), .B(n10215), .Z(n10207) );
  XNOR U11139 ( .A(n10194), .B(n10197), .Z(n10215) );
  NAND U11140 ( .A(A[2]), .B(B[568]), .Z(n10197) );
  NANDN U11141 ( .A(n10216), .B(n10217), .Z(n10194) );
  AND U11142 ( .A(A[0]), .B(B[569]), .Z(n10217) );
  XOR U11143 ( .A(n10199), .B(n10218), .Z(n10196) );
  NAND U11144 ( .A(A[0]), .B(B[570]), .Z(n10218) );
  NAND U11145 ( .A(B[569]), .B(A[1]), .Z(n10199) );
  NAND U11146 ( .A(n10219), .B(n10220), .Z(n989) );
  NANDN U11147 ( .A(n10221), .B(n10222), .Z(n10220) );
  OR U11148 ( .A(n10223), .B(n10224), .Z(n10222) );
  NAND U11149 ( .A(n10224), .B(n10223), .Z(n10219) );
  XOR U11150 ( .A(n991), .B(n990), .Z(\A1[567] ) );
  XOR U11151 ( .A(n10224), .B(n10225), .Z(n990) );
  XNOR U11152 ( .A(n10223), .B(n10221), .Z(n10225) );
  AND U11153 ( .A(n10226), .B(n10227), .Z(n10221) );
  NANDN U11154 ( .A(n10228), .B(n10229), .Z(n10227) );
  NANDN U11155 ( .A(n10230), .B(n10231), .Z(n10229) );
  AND U11156 ( .A(B[566]), .B(A[3]), .Z(n10223) );
  XNOR U11157 ( .A(n10213), .B(n10232), .Z(n10224) );
  XNOR U11158 ( .A(n10211), .B(n10214), .Z(n10232) );
  NAND U11159 ( .A(A[2]), .B(B[567]), .Z(n10214) );
  NANDN U11160 ( .A(n10233), .B(n10234), .Z(n10211) );
  AND U11161 ( .A(A[0]), .B(B[568]), .Z(n10234) );
  XOR U11162 ( .A(n10216), .B(n10235), .Z(n10213) );
  NAND U11163 ( .A(A[0]), .B(B[569]), .Z(n10235) );
  NAND U11164 ( .A(B[568]), .B(A[1]), .Z(n10216) );
  NAND U11165 ( .A(n10236), .B(n10237), .Z(n991) );
  NANDN U11166 ( .A(n10238), .B(n10239), .Z(n10237) );
  OR U11167 ( .A(n10240), .B(n10241), .Z(n10239) );
  NAND U11168 ( .A(n10241), .B(n10240), .Z(n10236) );
  XOR U11169 ( .A(n993), .B(n992), .Z(\A1[566] ) );
  XOR U11170 ( .A(n10241), .B(n10242), .Z(n992) );
  XNOR U11171 ( .A(n10240), .B(n10238), .Z(n10242) );
  AND U11172 ( .A(n10243), .B(n10244), .Z(n10238) );
  NANDN U11173 ( .A(n10245), .B(n10246), .Z(n10244) );
  NANDN U11174 ( .A(n10247), .B(n10248), .Z(n10246) );
  AND U11175 ( .A(B[565]), .B(A[3]), .Z(n10240) );
  XNOR U11176 ( .A(n10230), .B(n10249), .Z(n10241) );
  XNOR U11177 ( .A(n10228), .B(n10231), .Z(n10249) );
  NAND U11178 ( .A(A[2]), .B(B[566]), .Z(n10231) );
  NANDN U11179 ( .A(n10250), .B(n10251), .Z(n10228) );
  AND U11180 ( .A(A[0]), .B(B[567]), .Z(n10251) );
  XOR U11181 ( .A(n10233), .B(n10252), .Z(n10230) );
  NAND U11182 ( .A(A[0]), .B(B[568]), .Z(n10252) );
  NAND U11183 ( .A(B[567]), .B(A[1]), .Z(n10233) );
  NAND U11184 ( .A(n10253), .B(n10254), .Z(n993) );
  NANDN U11185 ( .A(n10255), .B(n10256), .Z(n10254) );
  OR U11186 ( .A(n10257), .B(n10258), .Z(n10256) );
  NAND U11187 ( .A(n10258), .B(n10257), .Z(n10253) );
  XOR U11188 ( .A(n995), .B(n994), .Z(\A1[565] ) );
  XOR U11189 ( .A(n10258), .B(n10259), .Z(n994) );
  XNOR U11190 ( .A(n10257), .B(n10255), .Z(n10259) );
  AND U11191 ( .A(n10260), .B(n10261), .Z(n10255) );
  NANDN U11192 ( .A(n10262), .B(n10263), .Z(n10261) );
  NANDN U11193 ( .A(n10264), .B(n10265), .Z(n10263) );
  AND U11194 ( .A(B[564]), .B(A[3]), .Z(n10257) );
  XNOR U11195 ( .A(n10247), .B(n10266), .Z(n10258) );
  XNOR U11196 ( .A(n10245), .B(n10248), .Z(n10266) );
  NAND U11197 ( .A(A[2]), .B(B[565]), .Z(n10248) );
  NANDN U11198 ( .A(n10267), .B(n10268), .Z(n10245) );
  AND U11199 ( .A(A[0]), .B(B[566]), .Z(n10268) );
  XOR U11200 ( .A(n10250), .B(n10269), .Z(n10247) );
  NAND U11201 ( .A(A[0]), .B(B[567]), .Z(n10269) );
  NAND U11202 ( .A(B[566]), .B(A[1]), .Z(n10250) );
  NAND U11203 ( .A(n10270), .B(n10271), .Z(n995) );
  NANDN U11204 ( .A(n10272), .B(n10273), .Z(n10271) );
  OR U11205 ( .A(n10274), .B(n10275), .Z(n10273) );
  NAND U11206 ( .A(n10275), .B(n10274), .Z(n10270) );
  XOR U11207 ( .A(n997), .B(n996), .Z(\A1[564] ) );
  XOR U11208 ( .A(n10275), .B(n10276), .Z(n996) );
  XNOR U11209 ( .A(n10274), .B(n10272), .Z(n10276) );
  AND U11210 ( .A(n10277), .B(n10278), .Z(n10272) );
  NANDN U11211 ( .A(n10279), .B(n10280), .Z(n10278) );
  NANDN U11212 ( .A(n10281), .B(n10282), .Z(n10280) );
  AND U11213 ( .A(B[563]), .B(A[3]), .Z(n10274) );
  XNOR U11214 ( .A(n10264), .B(n10283), .Z(n10275) );
  XNOR U11215 ( .A(n10262), .B(n10265), .Z(n10283) );
  NAND U11216 ( .A(A[2]), .B(B[564]), .Z(n10265) );
  NANDN U11217 ( .A(n10284), .B(n10285), .Z(n10262) );
  AND U11218 ( .A(A[0]), .B(B[565]), .Z(n10285) );
  XOR U11219 ( .A(n10267), .B(n10286), .Z(n10264) );
  NAND U11220 ( .A(A[0]), .B(B[566]), .Z(n10286) );
  NAND U11221 ( .A(B[565]), .B(A[1]), .Z(n10267) );
  NAND U11222 ( .A(n10287), .B(n10288), .Z(n997) );
  NANDN U11223 ( .A(n10289), .B(n10290), .Z(n10288) );
  OR U11224 ( .A(n10291), .B(n10292), .Z(n10290) );
  NAND U11225 ( .A(n10292), .B(n10291), .Z(n10287) );
  XOR U11226 ( .A(n999), .B(n998), .Z(\A1[563] ) );
  XOR U11227 ( .A(n10292), .B(n10293), .Z(n998) );
  XNOR U11228 ( .A(n10291), .B(n10289), .Z(n10293) );
  AND U11229 ( .A(n10294), .B(n10295), .Z(n10289) );
  NANDN U11230 ( .A(n10296), .B(n10297), .Z(n10295) );
  NANDN U11231 ( .A(n10298), .B(n10299), .Z(n10297) );
  AND U11232 ( .A(B[562]), .B(A[3]), .Z(n10291) );
  XNOR U11233 ( .A(n10281), .B(n10300), .Z(n10292) );
  XNOR U11234 ( .A(n10279), .B(n10282), .Z(n10300) );
  NAND U11235 ( .A(A[2]), .B(B[563]), .Z(n10282) );
  NANDN U11236 ( .A(n10301), .B(n10302), .Z(n10279) );
  AND U11237 ( .A(A[0]), .B(B[564]), .Z(n10302) );
  XOR U11238 ( .A(n10284), .B(n10303), .Z(n10281) );
  NAND U11239 ( .A(A[0]), .B(B[565]), .Z(n10303) );
  NAND U11240 ( .A(B[564]), .B(A[1]), .Z(n10284) );
  NAND U11241 ( .A(n10304), .B(n10305), .Z(n999) );
  NANDN U11242 ( .A(n10306), .B(n10307), .Z(n10305) );
  OR U11243 ( .A(n10308), .B(n10309), .Z(n10307) );
  NAND U11244 ( .A(n10309), .B(n10308), .Z(n10304) );
  XOR U11245 ( .A(n1001), .B(n1000), .Z(\A1[562] ) );
  XOR U11246 ( .A(n10309), .B(n10310), .Z(n1000) );
  XNOR U11247 ( .A(n10308), .B(n10306), .Z(n10310) );
  AND U11248 ( .A(n10311), .B(n10312), .Z(n10306) );
  NANDN U11249 ( .A(n10313), .B(n10314), .Z(n10312) );
  NANDN U11250 ( .A(n10315), .B(n10316), .Z(n10314) );
  AND U11251 ( .A(B[561]), .B(A[3]), .Z(n10308) );
  XNOR U11252 ( .A(n10298), .B(n10317), .Z(n10309) );
  XNOR U11253 ( .A(n10296), .B(n10299), .Z(n10317) );
  NAND U11254 ( .A(A[2]), .B(B[562]), .Z(n10299) );
  NANDN U11255 ( .A(n10318), .B(n10319), .Z(n10296) );
  AND U11256 ( .A(A[0]), .B(B[563]), .Z(n10319) );
  XOR U11257 ( .A(n10301), .B(n10320), .Z(n10298) );
  NAND U11258 ( .A(A[0]), .B(B[564]), .Z(n10320) );
  NAND U11259 ( .A(B[563]), .B(A[1]), .Z(n10301) );
  NAND U11260 ( .A(n10321), .B(n10322), .Z(n1001) );
  NANDN U11261 ( .A(n10323), .B(n10324), .Z(n10322) );
  OR U11262 ( .A(n10325), .B(n10326), .Z(n10324) );
  NAND U11263 ( .A(n10326), .B(n10325), .Z(n10321) );
  XOR U11264 ( .A(n1003), .B(n1002), .Z(\A1[561] ) );
  XOR U11265 ( .A(n10326), .B(n10327), .Z(n1002) );
  XNOR U11266 ( .A(n10325), .B(n10323), .Z(n10327) );
  AND U11267 ( .A(n10328), .B(n10329), .Z(n10323) );
  NANDN U11268 ( .A(n10330), .B(n10331), .Z(n10329) );
  NANDN U11269 ( .A(n10332), .B(n10333), .Z(n10331) );
  AND U11270 ( .A(B[560]), .B(A[3]), .Z(n10325) );
  XNOR U11271 ( .A(n10315), .B(n10334), .Z(n10326) );
  XNOR U11272 ( .A(n10313), .B(n10316), .Z(n10334) );
  NAND U11273 ( .A(A[2]), .B(B[561]), .Z(n10316) );
  NANDN U11274 ( .A(n10335), .B(n10336), .Z(n10313) );
  AND U11275 ( .A(A[0]), .B(B[562]), .Z(n10336) );
  XOR U11276 ( .A(n10318), .B(n10337), .Z(n10315) );
  NAND U11277 ( .A(A[0]), .B(B[563]), .Z(n10337) );
  NAND U11278 ( .A(B[562]), .B(A[1]), .Z(n10318) );
  NAND U11279 ( .A(n10338), .B(n10339), .Z(n1003) );
  NANDN U11280 ( .A(n10340), .B(n10341), .Z(n10339) );
  OR U11281 ( .A(n10342), .B(n10343), .Z(n10341) );
  NAND U11282 ( .A(n10343), .B(n10342), .Z(n10338) );
  XOR U11283 ( .A(n1005), .B(n1004), .Z(\A1[560] ) );
  XOR U11284 ( .A(n10343), .B(n10344), .Z(n1004) );
  XNOR U11285 ( .A(n10342), .B(n10340), .Z(n10344) );
  AND U11286 ( .A(n10345), .B(n10346), .Z(n10340) );
  NANDN U11287 ( .A(n10347), .B(n10348), .Z(n10346) );
  NANDN U11288 ( .A(n10349), .B(n10350), .Z(n10348) );
  AND U11289 ( .A(B[559]), .B(A[3]), .Z(n10342) );
  XNOR U11290 ( .A(n10332), .B(n10351), .Z(n10343) );
  XNOR U11291 ( .A(n10330), .B(n10333), .Z(n10351) );
  NAND U11292 ( .A(A[2]), .B(B[560]), .Z(n10333) );
  NANDN U11293 ( .A(n10352), .B(n10353), .Z(n10330) );
  AND U11294 ( .A(A[0]), .B(B[561]), .Z(n10353) );
  XOR U11295 ( .A(n10335), .B(n10354), .Z(n10332) );
  NAND U11296 ( .A(A[0]), .B(B[562]), .Z(n10354) );
  NAND U11297 ( .A(B[561]), .B(A[1]), .Z(n10335) );
  NAND U11298 ( .A(n10355), .B(n10356), .Z(n1005) );
  NANDN U11299 ( .A(n10357), .B(n10358), .Z(n10356) );
  OR U11300 ( .A(n10359), .B(n10360), .Z(n10358) );
  NAND U11301 ( .A(n10360), .B(n10359), .Z(n10355) );
  XOR U11302 ( .A(n987), .B(n986), .Z(\A1[55] ) );
  XOR U11303 ( .A(n10190), .B(n10361), .Z(n986) );
  XNOR U11304 ( .A(n10189), .B(n10187), .Z(n10361) );
  AND U11305 ( .A(n10362), .B(n10363), .Z(n10187) );
  NANDN U11306 ( .A(n10364), .B(n10365), .Z(n10363) );
  NANDN U11307 ( .A(n10366), .B(n10367), .Z(n10365) );
  AND U11308 ( .A(B[54]), .B(A[3]), .Z(n10189) );
  XNOR U11309 ( .A(n10179), .B(n10368), .Z(n10190) );
  XNOR U11310 ( .A(n10177), .B(n10180), .Z(n10368) );
  NAND U11311 ( .A(A[2]), .B(B[55]), .Z(n10180) );
  NANDN U11312 ( .A(n10369), .B(n10370), .Z(n10177) );
  AND U11313 ( .A(A[0]), .B(B[56]), .Z(n10370) );
  XOR U11314 ( .A(n10182), .B(n10371), .Z(n10179) );
  NAND U11315 ( .A(A[0]), .B(B[57]), .Z(n10371) );
  NAND U11316 ( .A(B[56]), .B(A[1]), .Z(n10182) );
  NAND U11317 ( .A(n10372), .B(n10373), .Z(n987) );
  NANDN U11318 ( .A(n10374), .B(n10375), .Z(n10373) );
  OR U11319 ( .A(n10376), .B(n10377), .Z(n10375) );
  NAND U11320 ( .A(n10377), .B(n10376), .Z(n10372) );
  XOR U11321 ( .A(n1007), .B(n1006), .Z(\A1[559] ) );
  XOR U11322 ( .A(n10360), .B(n10378), .Z(n1006) );
  XNOR U11323 ( .A(n10359), .B(n10357), .Z(n10378) );
  AND U11324 ( .A(n10379), .B(n10380), .Z(n10357) );
  NANDN U11325 ( .A(n10381), .B(n10382), .Z(n10380) );
  NANDN U11326 ( .A(n10383), .B(n10384), .Z(n10382) );
  AND U11327 ( .A(B[558]), .B(A[3]), .Z(n10359) );
  XNOR U11328 ( .A(n10349), .B(n10385), .Z(n10360) );
  XNOR U11329 ( .A(n10347), .B(n10350), .Z(n10385) );
  NAND U11330 ( .A(A[2]), .B(B[559]), .Z(n10350) );
  NANDN U11331 ( .A(n10386), .B(n10387), .Z(n10347) );
  AND U11332 ( .A(A[0]), .B(B[560]), .Z(n10387) );
  XOR U11333 ( .A(n10352), .B(n10388), .Z(n10349) );
  NAND U11334 ( .A(A[0]), .B(B[561]), .Z(n10388) );
  NAND U11335 ( .A(B[560]), .B(A[1]), .Z(n10352) );
  NAND U11336 ( .A(n10389), .B(n10390), .Z(n1007) );
  NANDN U11337 ( .A(n10391), .B(n10392), .Z(n10390) );
  OR U11338 ( .A(n10393), .B(n10394), .Z(n10392) );
  NAND U11339 ( .A(n10394), .B(n10393), .Z(n10389) );
  XOR U11340 ( .A(n1011), .B(n1010), .Z(\A1[558] ) );
  XOR U11341 ( .A(n10394), .B(n10395), .Z(n1010) );
  XNOR U11342 ( .A(n10393), .B(n10391), .Z(n10395) );
  AND U11343 ( .A(n10396), .B(n10397), .Z(n10391) );
  NANDN U11344 ( .A(n10398), .B(n10399), .Z(n10397) );
  NANDN U11345 ( .A(n10400), .B(n10401), .Z(n10399) );
  AND U11346 ( .A(B[557]), .B(A[3]), .Z(n10393) );
  XNOR U11347 ( .A(n10383), .B(n10402), .Z(n10394) );
  XNOR U11348 ( .A(n10381), .B(n10384), .Z(n10402) );
  NAND U11349 ( .A(A[2]), .B(B[558]), .Z(n10384) );
  NANDN U11350 ( .A(n10403), .B(n10404), .Z(n10381) );
  AND U11351 ( .A(A[0]), .B(B[559]), .Z(n10404) );
  XOR U11352 ( .A(n10386), .B(n10405), .Z(n10383) );
  NAND U11353 ( .A(A[0]), .B(B[560]), .Z(n10405) );
  NAND U11354 ( .A(B[559]), .B(A[1]), .Z(n10386) );
  NAND U11355 ( .A(n10406), .B(n10407), .Z(n1011) );
  NANDN U11356 ( .A(n10408), .B(n10409), .Z(n10407) );
  OR U11357 ( .A(n10410), .B(n10411), .Z(n10409) );
  NAND U11358 ( .A(n10411), .B(n10410), .Z(n10406) );
  XOR U11359 ( .A(n1013), .B(n1012), .Z(\A1[557] ) );
  XOR U11360 ( .A(n10411), .B(n10412), .Z(n1012) );
  XNOR U11361 ( .A(n10410), .B(n10408), .Z(n10412) );
  AND U11362 ( .A(n10413), .B(n10414), .Z(n10408) );
  NANDN U11363 ( .A(n10415), .B(n10416), .Z(n10414) );
  NANDN U11364 ( .A(n10417), .B(n10418), .Z(n10416) );
  AND U11365 ( .A(B[556]), .B(A[3]), .Z(n10410) );
  XNOR U11366 ( .A(n10400), .B(n10419), .Z(n10411) );
  XNOR U11367 ( .A(n10398), .B(n10401), .Z(n10419) );
  NAND U11368 ( .A(A[2]), .B(B[557]), .Z(n10401) );
  NANDN U11369 ( .A(n10420), .B(n10421), .Z(n10398) );
  AND U11370 ( .A(A[0]), .B(B[558]), .Z(n10421) );
  XOR U11371 ( .A(n10403), .B(n10422), .Z(n10400) );
  NAND U11372 ( .A(A[0]), .B(B[559]), .Z(n10422) );
  NAND U11373 ( .A(B[558]), .B(A[1]), .Z(n10403) );
  NAND U11374 ( .A(n10423), .B(n10424), .Z(n1013) );
  NANDN U11375 ( .A(n10425), .B(n10426), .Z(n10424) );
  OR U11376 ( .A(n10427), .B(n10428), .Z(n10426) );
  NAND U11377 ( .A(n10428), .B(n10427), .Z(n10423) );
  XOR U11378 ( .A(n1015), .B(n1014), .Z(\A1[556] ) );
  XOR U11379 ( .A(n10428), .B(n10429), .Z(n1014) );
  XNOR U11380 ( .A(n10427), .B(n10425), .Z(n10429) );
  AND U11381 ( .A(n10430), .B(n10431), .Z(n10425) );
  NANDN U11382 ( .A(n10432), .B(n10433), .Z(n10431) );
  NANDN U11383 ( .A(n10434), .B(n10435), .Z(n10433) );
  AND U11384 ( .A(B[555]), .B(A[3]), .Z(n10427) );
  XNOR U11385 ( .A(n10417), .B(n10436), .Z(n10428) );
  XNOR U11386 ( .A(n10415), .B(n10418), .Z(n10436) );
  NAND U11387 ( .A(A[2]), .B(B[556]), .Z(n10418) );
  NANDN U11388 ( .A(n10437), .B(n10438), .Z(n10415) );
  AND U11389 ( .A(A[0]), .B(B[557]), .Z(n10438) );
  XOR U11390 ( .A(n10420), .B(n10439), .Z(n10417) );
  NAND U11391 ( .A(A[0]), .B(B[558]), .Z(n10439) );
  NAND U11392 ( .A(B[557]), .B(A[1]), .Z(n10420) );
  NAND U11393 ( .A(n10440), .B(n10441), .Z(n1015) );
  NANDN U11394 ( .A(n10442), .B(n10443), .Z(n10441) );
  OR U11395 ( .A(n10444), .B(n10445), .Z(n10443) );
  NAND U11396 ( .A(n10445), .B(n10444), .Z(n10440) );
  XOR U11397 ( .A(n1017), .B(n1016), .Z(\A1[555] ) );
  XOR U11398 ( .A(n10445), .B(n10446), .Z(n1016) );
  XNOR U11399 ( .A(n10444), .B(n10442), .Z(n10446) );
  AND U11400 ( .A(n10447), .B(n10448), .Z(n10442) );
  NANDN U11401 ( .A(n10449), .B(n10450), .Z(n10448) );
  NANDN U11402 ( .A(n10451), .B(n10452), .Z(n10450) );
  AND U11403 ( .A(B[554]), .B(A[3]), .Z(n10444) );
  XNOR U11404 ( .A(n10434), .B(n10453), .Z(n10445) );
  XNOR U11405 ( .A(n10432), .B(n10435), .Z(n10453) );
  NAND U11406 ( .A(A[2]), .B(B[555]), .Z(n10435) );
  NANDN U11407 ( .A(n10454), .B(n10455), .Z(n10432) );
  AND U11408 ( .A(A[0]), .B(B[556]), .Z(n10455) );
  XOR U11409 ( .A(n10437), .B(n10456), .Z(n10434) );
  NAND U11410 ( .A(A[0]), .B(B[557]), .Z(n10456) );
  NAND U11411 ( .A(B[556]), .B(A[1]), .Z(n10437) );
  NAND U11412 ( .A(n10457), .B(n10458), .Z(n1017) );
  NANDN U11413 ( .A(n10459), .B(n10460), .Z(n10458) );
  OR U11414 ( .A(n10461), .B(n10462), .Z(n10460) );
  NAND U11415 ( .A(n10462), .B(n10461), .Z(n10457) );
  XOR U11416 ( .A(n1019), .B(n1018), .Z(\A1[554] ) );
  XOR U11417 ( .A(n10462), .B(n10463), .Z(n1018) );
  XNOR U11418 ( .A(n10461), .B(n10459), .Z(n10463) );
  AND U11419 ( .A(n10464), .B(n10465), .Z(n10459) );
  NANDN U11420 ( .A(n10466), .B(n10467), .Z(n10465) );
  NANDN U11421 ( .A(n10468), .B(n10469), .Z(n10467) );
  AND U11422 ( .A(B[553]), .B(A[3]), .Z(n10461) );
  XNOR U11423 ( .A(n10451), .B(n10470), .Z(n10462) );
  XNOR U11424 ( .A(n10449), .B(n10452), .Z(n10470) );
  NAND U11425 ( .A(A[2]), .B(B[554]), .Z(n10452) );
  NANDN U11426 ( .A(n10471), .B(n10472), .Z(n10449) );
  AND U11427 ( .A(A[0]), .B(B[555]), .Z(n10472) );
  XOR U11428 ( .A(n10454), .B(n10473), .Z(n10451) );
  NAND U11429 ( .A(A[0]), .B(B[556]), .Z(n10473) );
  NAND U11430 ( .A(B[555]), .B(A[1]), .Z(n10454) );
  NAND U11431 ( .A(n10474), .B(n10475), .Z(n1019) );
  NANDN U11432 ( .A(n10476), .B(n10477), .Z(n10475) );
  OR U11433 ( .A(n10478), .B(n10479), .Z(n10477) );
  NAND U11434 ( .A(n10479), .B(n10478), .Z(n10474) );
  XOR U11435 ( .A(n1021), .B(n1020), .Z(\A1[553] ) );
  XOR U11436 ( .A(n10479), .B(n10480), .Z(n1020) );
  XNOR U11437 ( .A(n10478), .B(n10476), .Z(n10480) );
  AND U11438 ( .A(n10481), .B(n10482), .Z(n10476) );
  NANDN U11439 ( .A(n10483), .B(n10484), .Z(n10482) );
  NANDN U11440 ( .A(n10485), .B(n10486), .Z(n10484) );
  AND U11441 ( .A(B[552]), .B(A[3]), .Z(n10478) );
  XNOR U11442 ( .A(n10468), .B(n10487), .Z(n10479) );
  XNOR U11443 ( .A(n10466), .B(n10469), .Z(n10487) );
  NAND U11444 ( .A(A[2]), .B(B[553]), .Z(n10469) );
  NANDN U11445 ( .A(n10488), .B(n10489), .Z(n10466) );
  AND U11446 ( .A(A[0]), .B(B[554]), .Z(n10489) );
  XOR U11447 ( .A(n10471), .B(n10490), .Z(n10468) );
  NAND U11448 ( .A(A[0]), .B(B[555]), .Z(n10490) );
  NAND U11449 ( .A(B[554]), .B(A[1]), .Z(n10471) );
  NAND U11450 ( .A(n10491), .B(n10492), .Z(n1021) );
  NANDN U11451 ( .A(n10493), .B(n10494), .Z(n10492) );
  OR U11452 ( .A(n10495), .B(n10496), .Z(n10494) );
  NAND U11453 ( .A(n10496), .B(n10495), .Z(n10491) );
  XOR U11454 ( .A(n1023), .B(n1022), .Z(\A1[552] ) );
  XOR U11455 ( .A(n10496), .B(n10497), .Z(n1022) );
  XNOR U11456 ( .A(n10495), .B(n10493), .Z(n10497) );
  AND U11457 ( .A(n10498), .B(n10499), .Z(n10493) );
  NANDN U11458 ( .A(n10500), .B(n10501), .Z(n10499) );
  NANDN U11459 ( .A(n10502), .B(n10503), .Z(n10501) );
  AND U11460 ( .A(B[551]), .B(A[3]), .Z(n10495) );
  XNOR U11461 ( .A(n10485), .B(n10504), .Z(n10496) );
  XNOR U11462 ( .A(n10483), .B(n10486), .Z(n10504) );
  NAND U11463 ( .A(A[2]), .B(B[552]), .Z(n10486) );
  NANDN U11464 ( .A(n10505), .B(n10506), .Z(n10483) );
  AND U11465 ( .A(A[0]), .B(B[553]), .Z(n10506) );
  XOR U11466 ( .A(n10488), .B(n10507), .Z(n10485) );
  NAND U11467 ( .A(A[0]), .B(B[554]), .Z(n10507) );
  NAND U11468 ( .A(B[553]), .B(A[1]), .Z(n10488) );
  NAND U11469 ( .A(n10508), .B(n10509), .Z(n1023) );
  NANDN U11470 ( .A(n10510), .B(n10511), .Z(n10509) );
  OR U11471 ( .A(n10512), .B(n10513), .Z(n10511) );
  NAND U11472 ( .A(n10513), .B(n10512), .Z(n10508) );
  XOR U11473 ( .A(n1025), .B(n1024), .Z(\A1[551] ) );
  XOR U11474 ( .A(n10513), .B(n10514), .Z(n1024) );
  XNOR U11475 ( .A(n10512), .B(n10510), .Z(n10514) );
  AND U11476 ( .A(n10515), .B(n10516), .Z(n10510) );
  NANDN U11477 ( .A(n10517), .B(n10518), .Z(n10516) );
  NANDN U11478 ( .A(n10519), .B(n10520), .Z(n10518) );
  AND U11479 ( .A(B[550]), .B(A[3]), .Z(n10512) );
  XNOR U11480 ( .A(n10502), .B(n10521), .Z(n10513) );
  XNOR U11481 ( .A(n10500), .B(n10503), .Z(n10521) );
  NAND U11482 ( .A(A[2]), .B(B[551]), .Z(n10503) );
  NANDN U11483 ( .A(n10522), .B(n10523), .Z(n10500) );
  AND U11484 ( .A(A[0]), .B(B[552]), .Z(n10523) );
  XOR U11485 ( .A(n10505), .B(n10524), .Z(n10502) );
  NAND U11486 ( .A(A[0]), .B(B[553]), .Z(n10524) );
  NAND U11487 ( .A(B[552]), .B(A[1]), .Z(n10505) );
  NAND U11488 ( .A(n10525), .B(n10526), .Z(n1025) );
  NANDN U11489 ( .A(n10527), .B(n10528), .Z(n10526) );
  OR U11490 ( .A(n10529), .B(n10530), .Z(n10528) );
  NAND U11491 ( .A(n10530), .B(n10529), .Z(n10525) );
  XOR U11492 ( .A(n1027), .B(n1026), .Z(\A1[550] ) );
  XOR U11493 ( .A(n10530), .B(n10531), .Z(n1026) );
  XNOR U11494 ( .A(n10529), .B(n10527), .Z(n10531) );
  AND U11495 ( .A(n10532), .B(n10533), .Z(n10527) );
  NANDN U11496 ( .A(n10534), .B(n10535), .Z(n10533) );
  NANDN U11497 ( .A(n10536), .B(n10537), .Z(n10535) );
  AND U11498 ( .A(B[549]), .B(A[3]), .Z(n10529) );
  XNOR U11499 ( .A(n10519), .B(n10538), .Z(n10530) );
  XNOR U11500 ( .A(n10517), .B(n10520), .Z(n10538) );
  NAND U11501 ( .A(A[2]), .B(B[550]), .Z(n10520) );
  NANDN U11502 ( .A(n10539), .B(n10540), .Z(n10517) );
  AND U11503 ( .A(A[0]), .B(B[551]), .Z(n10540) );
  XOR U11504 ( .A(n10522), .B(n10541), .Z(n10519) );
  NAND U11505 ( .A(A[0]), .B(B[552]), .Z(n10541) );
  NAND U11506 ( .A(B[551]), .B(A[1]), .Z(n10522) );
  NAND U11507 ( .A(n10542), .B(n10543), .Z(n1027) );
  NANDN U11508 ( .A(n10544), .B(n10545), .Z(n10543) );
  OR U11509 ( .A(n10546), .B(n10547), .Z(n10545) );
  NAND U11510 ( .A(n10547), .B(n10546), .Z(n10542) );
  XOR U11511 ( .A(n1009), .B(n1008), .Z(\A1[54] ) );
  XOR U11512 ( .A(n10377), .B(n10548), .Z(n1008) );
  XNOR U11513 ( .A(n10376), .B(n10374), .Z(n10548) );
  AND U11514 ( .A(n10549), .B(n10550), .Z(n10374) );
  NANDN U11515 ( .A(n10551), .B(n10552), .Z(n10550) );
  NANDN U11516 ( .A(n10553), .B(n10554), .Z(n10552) );
  AND U11517 ( .A(B[53]), .B(A[3]), .Z(n10376) );
  XNOR U11518 ( .A(n10366), .B(n10555), .Z(n10377) );
  XNOR U11519 ( .A(n10364), .B(n10367), .Z(n10555) );
  NAND U11520 ( .A(A[2]), .B(B[54]), .Z(n10367) );
  NANDN U11521 ( .A(n10556), .B(n10557), .Z(n10364) );
  AND U11522 ( .A(A[0]), .B(B[55]), .Z(n10557) );
  XOR U11523 ( .A(n10369), .B(n10558), .Z(n10366) );
  NAND U11524 ( .A(A[0]), .B(B[56]), .Z(n10558) );
  NAND U11525 ( .A(B[55]), .B(A[1]), .Z(n10369) );
  NAND U11526 ( .A(n10559), .B(n10560), .Z(n1009) );
  NANDN U11527 ( .A(n10561), .B(n10562), .Z(n10560) );
  OR U11528 ( .A(n10563), .B(n10564), .Z(n10562) );
  NAND U11529 ( .A(n10564), .B(n10563), .Z(n10559) );
  XOR U11530 ( .A(n1029), .B(n1028), .Z(\A1[549] ) );
  XOR U11531 ( .A(n10547), .B(n10565), .Z(n1028) );
  XNOR U11532 ( .A(n10546), .B(n10544), .Z(n10565) );
  AND U11533 ( .A(n10566), .B(n10567), .Z(n10544) );
  NANDN U11534 ( .A(n10568), .B(n10569), .Z(n10567) );
  NANDN U11535 ( .A(n10570), .B(n10571), .Z(n10569) );
  AND U11536 ( .A(B[548]), .B(A[3]), .Z(n10546) );
  XNOR U11537 ( .A(n10536), .B(n10572), .Z(n10547) );
  XNOR U11538 ( .A(n10534), .B(n10537), .Z(n10572) );
  NAND U11539 ( .A(A[2]), .B(B[549]), .Z(n10537) );
  NANDN U11540 ( .A(n10573), .B(n10574), .Z(n10534) );
  AND U11541 ( .A(A[0]), .B(B[550]), .Z(n10574) );
  XOR U11542 ( .A(n10539), .B(n10575), .Z(n10536) );
  NAND U11543 ( .A(A[0]), .B(B[551]), .Z(n10575) );
  NAND U11544 ( .A(B[550]), .B(A[1]), .Z(n10539) );
  NAND U11545 ( .A(n10576), .B(n10577), .Z(n1029) );
  NANDN U11546 ( .A(n10578), .B(n10579), .Z(n10577) );
  OR U11547 ( .A(n10580), .B(n10581), .Z(n10579) );
  NAND U11548 ( .A(n10581), .B(n10580), .Z(n10576) );
  XOR U11549 ( .A(n1033), .B(n1032), .Z(\A1[548] ) );
  XOR U11550 ( .A(n10581), .B(n10582), .Z(n1032) );
  XNOR U11551 ( .A(n10580), .B(n10578), .Z(n10582) );
  AND U11552 ( .A(n10583), .B(n10584), .Z(n10578) );
  NANDN U11553 ( .A(n10585), .B(n10586), .Z(n10584) );
  NANDN U11554 ( .A(n10587), .B(n10588), .Z(n10586) );
  AND U11555 ( .A(B[547]), .B(A[3]), .Z(n10580) );
  XNOR U11556 ( .A(n10570), .B(n10589), .Z(n10581) );
  XNOR U11557 ( .A(n10568), .B(n10571), .Z(n10589) );
  NAND U11558 ( .A(A[2]), .B(B[548]), .Z(n10571) );
  NANDN U11559 ( .A(n10590), .B(n10591), .Z(n10568) );
  AND U11560 ( .A(A[0]), .B(B[549]), .Z(n10591) );
  XOR U11561 ( .A(n10573), .B(n10592), .Z(n10570) );
  NAND U11562 ( .A(A[0]), .B(B[550]), .Z(n10592) );
  NAND U11563 ( .A(B[549]), .B(A[1]), .Z(n10573) );
  NAND U11564 ( .A(n10593), .B(n10594), .Z(n1033) );
  NANDN U11565 ( .A(n10595), .B(n10596), .Z(n10594) );
  OR U11566 ( .A(n10597), .B(n10598), .Z(n10596) );
  NAND U11567 ( .A(n10598), .B(n10597), .Z(n10593) );
  XOR U11568 ( .A(n1035), .B(n1034), .Z(\A1[547] ) );
  XOR U11569 ( .A(n10598), .B(n10599), .Z(n1034) );
  XNOR U11570 ( .A(n10597), .B(n10595), .Z(n10599) );
  AND U11571 ( .A(n10600), .B(n10601), .Z(n10595) );
  NANDN U11572 ( .A(n10602), .B(n10603), .Z(n10601) );
  NANDN U11573 ( .A(n10604), .B(n10605), .Z(n10603) );
  AND U11574 ( .A(B[546]), .B(A[3]), .Z(n10597) );
  XNOR U11575 ( .A(n10587), .B(n10606), .Z(n10598) );
  XNOR U11576 ( .A(n10585), .B(n10588), .Z(n10606) );
  NAND U11577 ( .A(A[2]), .B(B[547]), .Z(n10588) );
  NANDN U11578 ( .A(n10607), .B(n10608), .Z(n10585) );
  AND U11579 ( .A(A[0]), .B(B[548]), .Z(n10608) );
  XOR U11580 ( .A(n10590), .B(n10609), .Z(n10587) );
  NAND U11581 ( .A(A[0]), .B(B[549]), .Z(n10609) );
  NAND U11582 ( .A(B[548]), .B(A[1]), .Z(n10590) );
  NAND U11583 ( .A(n10610), .B(n10611), .Z(n1035) );
  NANDN U11584 ( .A(n10612), .B(n10613), .Z(n10611) );
  OR U11585 ( .A(n10614), .B(n10615), .Z(n10613) );
  NAND U11586 ( .A(n10615), .B(n10614), .Z(n10610) );
  XOR U11587 ( .A(n1037), .B(n1036), .Z(\A1[546] ) );
  XOR U11588 ( .A(n10615), .B(n10616), .Z(n1036) );
  XNOR U11589 ( .A(n10614), .B(n10612), .Z(n10616) );
  AND U11590 ( .A(n10617), .B(n10618), .Z(n10612) );
  NANDN U11591 ( .A(n10619), .B(n10620), .Z(n10618) );
  NANDN U11592 ( .A(n10621), .B(n10622), .Z(n10620) );
  AND U11593 ( .A(B[545]), .B(A[3]), .Z(n10614) );
  XNOR U11594 ( .A(n10604), .B(n10623), .Z(n10615) );
  XNOR U11595 ( .A(n10602), .B(n10605), .Z(n10623) );
  NAND U11596 ( .A(A[2]), .B(B[546]), .Z(n10605) );
  NANDN U11597 ( .A(n10624), .B(n10625), .Z(n10602) );
  AND U11598 ( .A(A[0]), .B(B[547]), .Z(n10625) );
  XOR U11599 ( .A(n10607), .B(n10626), .Z(n10604) );
  NAND U11600 ( .A(A[0]), .B(B[548]), .Z(n10626) );
  NAND U11601 ( .A(B[547]), .B(A[1]), .Z(n10607) );
  NAND U11602 ( .A(n10627), .B(n10628), .Z(n1037) );
  NANDN U11603 ( .A(n10629), .B(n10630), .Z(n10628) );
  OR U11604 ( .A(n10631), .B(n10632), .Z(n10630) );
  NAND U11605 ( .A(n10632), .B(n10631), .Z(n10627) );
  XOR U11606 ( .A(n1039), .B(n1038), .Z(\A1[545] ) );
  XOR U11607 ( .A(n10632), .B(n10633), .Z(n1038) );
  XNOR U11608 ( .A(n10631), .B(n10629), .Z(n10633) );
  AND U11609 ( .A(n10634), .B(n10635), .Z(n10629) );
  NANDN U11610 ( .A(n10636), .B(n10637), .Z(n10635) );
  NANDN U11611 ( .A(n10638), .B(n10639), .Z(n10637) );
  AND U11612 ( .A(B[544]), .B(A[3]), .Z(n10631) );
  XNOR U11613 ( .A(n10621), .B(n10640), .Z(n10632) );
  XNOR U11614 ( .A(n10619), .B(n10622), .Z(n10640) );
  NAND U11615 ( .A(A[2]), .B(B[545]), .Z(n10622) );
  NANDN U11616 ( .A(n10641), .B(n10642), .Z(n10619) );
  AND U11617 ( .A(A[0]), .B(B[546]), .Z(n10642) );
  XOR U11618 ( .A(n10624), .B(n10643), .Z(n10621) );
  NAND U11619 ( .A(A[0]), .B(B[547]), .Z(n10643) );
  NAND U11620 ( .A(B[546]), .B(A[1]), .Z(n10624) );
  NAND U11621 ( .A(n10644), .B(n10645), .Z(n1039) );
  NANDN U11622 ( .A(n10646), .B(n10647), .Z(n10645) );
  OR U11623 ( .A(n10648), .B(n10649), .Z(n10647) );
  NAND U11624 ( .A(n10649), .B(n10648), .Z(n10644) );
  XOR U11625 ( .A(n1041), .B(n1040), .Z(\A1[544] ) );
  XOR U11626 ( .A(n10649), .B(n10650), .Z(n1040) );
  XNOR U11627 ( .A(n10648), .B(n10646), .Z(n10650) );
  AND U11628 ( .A(n10651), .B(n10652), .Z(n10646) );
  NANDN U11629 ( .A(n10653), .B(n10654), .Z(n10652) );
  NANDN U11630 ( .A(n10655), .B(n10656), .Z(n10654) );
  AND U11631 ( .A(B[543]), .B(A[3]), .Z(n10648) );
  XNOR U11632 ( .A(n10638), .B(n10657), .Z(n10649) );
  XNOR U11633 ( .A(n10636), .B(n10639), .Z(n10657) );
  NAND U11634 ( .A(A[2]), .B(B[544]), .Z(n10639) );
  NANDN U11635 ( .A(n10658), .B(n10659), .Z(n10636) );
  AND U11636 ( .A(A[0]), .B(B[545]), .Z(n10659) );
  XOR U11637 ( .A(n10641), .B(n10660), .Z(n10638) );
  NAND U11638 ( .A(A[0]), .B(B[546]), .Z(n10660) );
  NAND U11639 ( .A(B[545]), .B(A[1]), .Z(n10641) );
  NAND U11640 ( .A(n10661), .B(n10662), .Z(n1041) );
  NANDN U11641 ( .A(n10663), .B(n10664), .Z(n10662) );
  OR U11642 ( .A(n10665), .B(n10666), .Z(n10664) );
  NAND U11643 ( .A(n10666), .B(n10665), .Z(n10661) );
  XOR U11644 ( .A(n1043), .B(n1042), .Z(\A1[543] ) );
  XOR U11645 ( .A(n10666), .B(n10667), .Z(n1042) );
  XNOR U11646 ( .A(n10665), .B(n10663), .Z(n10667) );
  AND U11647 ( .A(n10668), .B(n10669), .Z(n10663) );
  NANDN U11648 ( .A(n10670), .B(n10671), .Z(n10669) );
  NANDN U11649 ( .A(n10672), .B(n10673), .Z(n10671) );
  AND U11650 ( .A(B[542]), .B(A[3]), .Z(n10665) );
  XNOR U11651 ( .A(n10655), .B(n10674), .Z(n10666) );
  XNOR U11652 ( .A(n10653), .B(n10656), .Z(n10674) );
  NAND U11653 ( .A(A[2]), .B(B[543]), .Z(n10656) );
  NANDN U11654 ( .A(n10675), .B(n10676), .Z(n10653) );
  AND U11655 ( .A(A[0]), .B(B[544]), .Z(n10676) );
  XOR U11656 ( .A(n10658), .B(n10677), .Z(n10655) );
  NAND U11657 ( .A(A[0]), .B(B[545]), .Z(n10677) );
  NAND U11658 ( .A(B[544]), .B(A[1]), .Z(n10658) );
  NAND U11659 ( .A(n10678), .B(n10679), .Z(n1043) );
  NANDN U11660 ( .A(n10680), .B(n10681), .Z(n10679) );
  OR U11661 ( .A(n10682), .B(n10683), .Z(n10681) );
  NAND U11662 ( .A(n10683), .B(n10682), .Z(n10678) );
  XOR U11663 ( .A(n1045), .B(n1044), .Z(\A1[542] ) );
  XOR U11664 ( .A(n10683), .B(n10684), .Z(n1044) );
  XNOR U11665 ( .A(n10682), .B(n10680), .Z(n10684) );
  AND U11666 ( .A(n10685), .B(n10686), .Z(n10680) );
  NANDN U11667 ( .A(n10687), .B(n10688), .Z(n10686) );
  NANDN U11668 ( .A(n10689), .B(n10690), .Z(n10688) );
  AND U11669 ( .A(B[541]), .B(A[3]), .Z(n10682) );
  XNOR U11670 ( .A(n10672), .B(n10691), .Z(n10683) );
  XNOR U11671 ( .A(n10670), .B(n10673), .Z(n10691) );
  NAND U11672 ( .A(A[2]), .B(B[542]), .Z(n10673) );
  NANDN U11673 ( .A(n10692), .B(n10693), .Z(n10670) );
  AND U11674 ( .A(A[0]), .B(B[543]), .Z(n10693) );
  XOR U11675 ( .A(n10675), .B(n10694), .Z(n10672) );
  NAND U11676 ( .A(A[0]), .B(B[544]), .Z(n10694) );
  NAND U11677 ( .A(B[543]), .B(A[1]), .Z(n10675) );
  NAND U11678 ( .A(n10695), .B(n10696), .Z(n1045) );
  NANDN U11679 ( .A(n10697), .B(n10698), .Z(n10696) );
  OR U11680 ( .A(n10699), .B(n10700), .Z(n10698) );
  NAND U11681 ( .A(n10700), .B(n10699), .Z(n10695) );
  XOR U11682 ( .A(n1047), .B(n1046), .Z(\A1[541] ) );
  XOR U11683 ( .A(n10700), .B(n10701), .Z(n1046) );
  XNOR U11684 ( .A(n10699), .B(n10697), .Z(n10701) );
  AND U11685 ( .A(n10702), .B(n10703), .Z(n10697) );
  NANDN U11686 ( .A(n10704), .B(n10705), .Z(n10703) );
  NANDN U11687 ( .A(n10706), .B(n10707), .Z(n10705) );
  AND U11688 ( .A(B[540]), .B(A[3]), .Z(n10699) );
  XNOR U11689 ( .A(n10689), .B(n10708), .Z(n10700) );
  XNOR U11690 ( .A(n10687), .B(n10690), .Z(n10708) );
  NAND U11691 ( .A(A[2]), .B(B[541]), .Z(n10690) );
  NANDN U11692 ( .A(n10709), .B(n10710), .Z(n10687) );
  AND U11693 ( .A(A[0]), .B(B[542]), .Z(n10710) );
  XOR U11694 ( .A(n10692), .B(n10711), .Z(n10689) );
  NAND U11695 ( .A(A[0]), .B(B[543]), .Z(n10711) );
  NAND U11696 ( .A(B[542]), .B(A[1]), .Z(n10692) );
  NAND U11697 ( .A(n10712), .B(n10713), .Z(n1047) );
  NANDN U11698 ( .A(n10714), .B(n10715), .Z(n10713) );
  OR U11699 ( .A(n10716), .B(n10717), .Z(n10715) );
  NAND U11700 ( .A(n10717), .B(n10716), .Z(n10712) );
  XOR U11701 ( .A(n1049), .B(n1048), .Z(\A1[540] ) );
  XOR U11702 ( .A(n10717), .B(n10718), .Z(n1048) );
  XNOR U11703 ( .A(n10716), .B(n10714), .Z(n10718) );
  AND U11704 ( .A(n10719), .B(n10720), .Z(n10714) );
  NANDN U11705 ( .A(n10721), .B(n10722), .Z(n10720) );
  NANDN U11706 ( .A(n10723), .B(n10724), .Z(n10722) );
  AND U11707 ( .A(B[539]), .B(A[3]), .Z(n10716) );
  XNOR U11708 ( .A(n10706), .B(n10725), .Z(n10717) );
  XNOR U11709 ( .A(n10704), .B(n10707), .Z(n10725) );
  NAND U11710 ( .A(A[2]), .B(B[540]), .Z(n10707) );
  NANDN U11711 ( .A(n10726), .B(n10727), .Z(n10704) );
  AND U11712 ( .A(A[0]), .B(B[541]), .Z(n10727) );
  XOR U11713 ( .A(n10709), .B(n10728), .Z(n10706) );
  NAND U11714 ( .A(A[0]), .B(B[542]), .Z(n10728) );
  NAND U11715 ( .A(B[541]), .B(A[1]), .Z(n10709) );
  NAND U11716 ( .A(n10729), .B(n10730), .Z(n1049) );
  NANDN U11717 ( .A(n10731), .B(n10732), .Z(n10730) );
  OR U11718 ( .A(n10733), .B(n10734), .Z(n10732) );
  NAND U11719 ( .A(n10734), .B(n10733), .Z(n10729) );
  XOR U11720 ( .A(n1031), .B(n1030), .Z(\A1[53] ) );
  XOR U11721 ( .A(n10564), .B(n10735), .Z(n1030) );
  XNOR U11722 ( .A(n10563), .B(n10561), .Z(n10735) );
  AND U11723 ( .A(n10736), .B(n10737), .Z(n10561) );
  NANDN U11724 ( .A(n10738), .B(n10739), .Z(n10737) );
  NANDN U11725 ( .A(n10740), .B(n10741), .Z(n10739) );
  AND U11726 ( .A(B[52]), .B(A[3]), .Z(n10563) );
  XNOR U11727 ( .A(n10553), .B(n10742), .Z(n10564) );
  XNOR U11728 ( .A(n10551), .B(n10554), .Z(n10742) );
  NAND U11729 ( .A(A[2]), .B(B[53]), .Z(n10554) );
  NANDN U11730 ( .A(n10743), .B(n10744), .Z(n10551) );
  AND U11731 ( .A(A[0]), .B(B[54]), .Z(n10744) );
  XOR U11732 ( .A(n10556), .B(n10745), .Z(n10553) );
  NAND U11733 ( .A(A[0]), .B(B[55]), .Z(n10745) );
  NAND U11734 ( .A(B[54]), .B(A[1]), .Z(n10556) );
  NAND U11735 ( .A(n10746), .B(n10747), .Z(n1031) );
  NANDN U11736 ( .A(n10748), .B(n10749), .Z(n10747) );
  OR U11737 ( .A(n10750), .B(n10751), .Z(n10749) );
  NAND U11738 ( .A(n10751), .B(n10750), .Z(n10746) );
  XOR U11739 ( .A(n1051), .B(n1050), .Z(\A1[539] ) );
  XOR U11740 ( .A(n10734), .B(n10752), .Z(n1050) );
  XNOR U11741 ( .A(n10733), .B(n10731), .Z(n10752) );
  AND U11742 ( .A(n10753), .B(n10754), .Z(n10731) );
  NANDN U11743 ( .A(n10755), .B(n10756), .Z(n10754) );
  NANDN U11744 ( .A(n10757), .B(n10758), .Z(n10756) );
  AND U11745 ( .A(B[538]), .B(A[3]), .Z(n10733) );
  XNOR U11746 ( .A(n10723), .B(n10759), .Z(n10734) );
  XNOR U11747 ( .A(n10721), .B(n10724), .Z(n10759) );
  NAND U11748 ( .A(A[2]), .B(B[539]), .Z(n10724) );
  NANDN U11749 ( .A(n10760), .B(n10761), .Z(n10721) );
  AND U11750 ( .A(A[0]), .B(B[540]), .Z(n10761) );
  XOR U11751 ( .A(n10726), .B(n10762), .Z(n10723) );
  NAND U11752 ( .A(A[0]), .B(B[541]), .Z(n10762) );
  NAND U11753 ( .A(B[540]), .B(A[1]), .Z(n10726) );
  NAND U11754 ( .A(n10763), .B(n10764), .Z(n1051) );
  NANDN U11755 ( .A(n10765), .B(n10766), .Z(n10764) );
  OR U11756 ( .A(n10767), .B(n10768), .Z(n10766) );
  NAND U11757 ( .A(n10768), .B(n10767), .Z(n10763) );
  XOR U11758 ( .A(n1055), .B(n1054), .Z(\A1[538] ) );
  XOR U11759 ( .A(n10768), .B(n10769), .Z(n1054) );
  XNOR U11760 ( .A(n10767), .B(n10765), .Z(n10769) );
  AND U11761 ( .A(n10770), .B(n10771), .Z(n10765) );
  NANDN U11762 ( .A(n10772), .B(n10773), .Z(n10771) );
  NANDN U11763 ( .A(n10774), .B(n10775), .Z(n10773) );
  AND U11764 ( .A(B[537]), .B(A[3]), .Z(n10767) );
  XNOR U11765 ( .A(n10757), .B(n10776), .Z(n10768) );
  XNOR U11766 ( .A(n10755), .B(n10758), .Z(n10776) );
  NAND U11767 ( .A(A[2]), .B(B[538]), .Z(n10758) );
  NANDN U11768 ( .A(n10777), .B(n10778), .Z(n10755) );
  AND U11769 ( .A(A[0]), .B(B[539]), .Z(n10778) );
  XOR U11770 ( .A(n10760), .B(n10779), .Z(n10757) );
  NAND U11771 ( .A(A[0]), .B(B[540]), .Z(n10779) );
  NAND U11772 ( .A(B[539]), .B(A[1]), .Z(n10760) );
  NAND U11773 ( .A(n10780), .B(n10781), .Z(n1055) );
  NANDN U11774 ( .A(n10782), .B(n10783), .Z(n10781) );
  OR U11775 ( .A(n10784), .B(n10785), .Z(n10783) );
  NAND U11776 ( .A(n10785), .B(n10784), .Z(n10780) );
  XOR U11777 ( .A(n1057), .B(n1056), .Z(\A1[537] ) );
  XOR U11778 ( .A(n10785), .B(n10786), .Z(n1056) );
  XNOR U11779 ( .A(n10784), .B(n10782), .Z(n10786) );
  AND U11780 ( .A(n10787), .B(n10788), .Z(n10782) );
  NANDN U11781 ( .A(n10789), .B(n10790), .Z(n10788) );
  NANDN U11782 ( .A(n10791), .B(n10792), .Z(n10790) );
  AND U11783 ( .A(B[536]), .B(A[3]), .Z(n10784) );
  XNOR U11784 ( .A(n10774), .B(n10793), .Z(n10785) );
  XNOR U11785 ( .A(n10772), .B(n10775), .Z(n10793) );
  NAND U11786 ( .A(A[2]), .B(B[537]), .Z(n10775) );
  NANDN U11787 ( .A(n10794), .B(n10795), .Z(n10772) );
  AND U11788 ( .A(A[0]), .B(B[538]), .Z(n10795) );
  XOR U11789 ( .A(n10777), .B(n10796), .Z(n10774) );
  NAND U11790 ( .A(A[0]), .B(B[539]), .Z(n10796) );
  NAND U11791 ( .A(B[538]), .B(A[1]), .Z(n10777) );
  NAND U11792 ( .A(n10797), .B(n10798), .Z(n1057) );
  NANDN U11793 ( .A(n10799), .B(n10800), .Z(n10798) );
  OR U11794 ( .A(n10801), .B(n10802), .Z(n10800) );
  NAND U11795 ( .A(n10802), .B(n10801), .Z(n10797) );
  XOR U11796 ( .A(n1059), .B(n1058), .Z(\A1[536] ) );
  XOR U11797 ( .A(n10802), .B(n10803), .Z(n1058) );
  XNOR U11798 ( .A(n10801), .B(n10799), .Z(n10803) );
  AND U11799 ( .A(n10804), .B(n10805), .Z(n10799) );
  NANDN U11800 ( .A(n10806), .B(n10807), .Z(n10805) );
  NANDN U11801 ( .A(n10808), .B(n10809), .Z(n10807) );
  AND U11802 ( .A(B[535]), .B(A[3]), .Z(n10801) );
  XNOR U11803 ( .A(n10791), .B(n10810), .Z(n10802) );
  XNOR U11804 ( .A(n10789), .B(n10792), .Z(n10810) );
  NAND U11805 ( .A(A[2]), .B(B[536]), .Z(n10792) );
  NANDN U11806 ( .A(n10811), .B(n10812), .Z(n10789) );
  AND U11807 ( .A(A[0]), .B(B[537]), .Z(n10812) );
  XOR U11808 ( .A(n10794), .B(n10813), .Z(n10791) );
  NAND U11809 ( .A(A[0]), .B(B[538]), .Z(n10813) );
  NAND U11810 ( .A(B[537]), .B(A[1]), .Z(n10794) );
  NAND U11811 ( .A(n10814), .B(n10815), .Z(n1059) );
  NANDN U11812 ( .A(n10816), .B(n10817), .Z(n10815) );
  OR U11813 ( .A(n10818), .B(n10819), .Z(n10817) );
  NAND U11814 ( .A(n10819), .B(n10818), .Z(n10814) );
  XOR U11815 ( .A(n1061), .B(n1060), .Z(\A1[535] ) );
  XOR U11816 ( .A(n10819), .B(n10820), .Z(n1060) );
  XNOR U11817 ( .A(n10818), .B(n10816), .Z(n10820) );
  AND U11818 ( .A(n10821), .B(n10822), .Z(n10816) );
  NANDN U11819 ( .A(n10823), .B(n10824), .Z(n10822) );
  NANDN U11820 ( .A(n10825), .B(n10826), .Z(n10824) );
  AND U11821 ( .A(B[534]), .B(A[3]), .Z(n10818) );
  XNOR U11822 ( .A(n10808), .B(n10827), .Z(n10819) );
  XNOR U11823 ( .A(n10806), .B(n10809), .Z(n10827) );
  NAND U11824 ( .A(A[2]), .B(B[535]), .Z(n10809) );
  NANDN U11825 ( .A(n10828), .B(n10829), .Z(n10806) );
  AND U11826 ( .A(A[0]), .B(B[536]), .Z(n10829) );
  XOR U11827 ( .A(n10811), .B(n10830), .Z(n10808) );
  NAND U11828 ( .A(A[0]), .B(B[537]), .Z(n10830) );
  NAND U11829 ( .A(B[536]), .B(A[1]), .Z(n10811) );
  NAND U11830 ( .A(n10831), .B(n10832), .Z(n1061) );
  NANDN U11831 ( .A(n10833), .B(n10834), .Z(n10832) );
  OR U11832 ( .A(n10835), .B(n10836), .Z(n10834) );
  NAND U11833 ( .A(n10836), .B(n10835), .Z(n10831) );
  XOR U11834 ( .A(n1063), .B(n1062), .Z(\A1[534] ) );
  XOR U11835 ( .A(n10836), .B(n10837), .Z(n1062) );
  XNOR U11836 ( .A(n10835), .B(n10833), .Z(n10837) );
  AND U11837 ( .A(n10838), .B(n10839), .Z(n10833) );
  NANDN U11838 ( .A(n10840), .B(n10841), .Z(n10839) );
  NANDN U11839 ( .A(n10842), .B(n10843), .Z(n10841) );
  AND U11840 ( .A(B[533]), .B(A[3]), .Z(n10835) );
  XNOR U11841 ( .A(n10825), .B(n10844), .Z(n10836) );
  XNOR U11842 ( .A(n10823), .B(n10826), .Z(n10844) );
  NAND U11843 ( .A(A[2]), .B(B[534]), .Z(n10826) );
  NANDN U11844 ( .A(n10845), .B(n10846), .Z(n10823) );
  AND U11845 ( .A(A[0]), .B(B[535]), .Z(n10846) );
  XOR U11846 ( .A(n10828), .B(n10847), .Z(n10825) );
  NAND U11847 ( .A(A[0]), .B(B[536]), .Z(n10847) );
  NAND U11848 ( .A(B[535]), .B(A[1]), .Z(n10828) );
  NAND U11849 ( .A(n10848), .B(n10849), .Z(n1063) );
  NANDN U11850 ( .A(n10850), .B(n10851), .Z(n10849) );
  OR U11851 ( .A(n10852), .B(n10853), .Z(n10851) );
  NAND U11852 ( .A(n10853), .B(n10852), .Z(n10848) );
  XOR U11853 ( .A(n1065), .B(n1064), .Z(\A1[533] ) );
  XOR U11854 ( .A(n10853), .B(n10854), .Z(n1064) );
  XNOR U11855 ( .A(n10852), .B(n10850), .Z(n10854) );
  AND U11856 ( .A(n10855), .B(n10856), .Z(n10850) );
  NANDN U11857 ( .A(n10857), .B(n10858), .Z(n10856) );
  NANDN U11858 ( .A(n10859), .B(n10860), .Z(n10858) );
  AND U11859 ( .A(B[532]), .B(A[3]), .Z(n10852) );
  XNOR U11860 ( .A(n10842), .B(n10861), .Z(n10853) );
  XNOR U11861 ( .A(n10840), .B(n10843), .Z(n10861) );
  NAND U11862 ( .A(A[2]), .B(B[533]), .Z(n10843) );
  NANDN U11863 ( .A(n10862), .B(n10863), .Z(n10840) );
  AND U11864 ( .A(A[0]), .B(B[534]), .Z(n10863) );
  XOR U11865 ( .A(n10845), .B(n10864), .Z(n10842) );
  NAND U11866 ( .A(A[0]), .B(B[535]), .Z(n10864) );
  NAND U11867 ( .A(B[534]), .B(A[1]), .Z(n10845) );
  NAND U11868 ( .A(n10865), .B(n10866), .Z(n1065) );
  NANDN U11869 ( .A(n10867), .B(n10868), .Z(n10866) );
  OR U11870 ( .A(n10869), .B(n10870), .Z(n10868) );
  NAND U11871 ( .A(n10870), .B(n10869), .Z(n10865) );
  XOR U11872 ( .A(n1067), .B(n1066), .Z(\A1[532] ) );
  XOR U11873 ( .A(n10870), .B(n10871), .Z(n1066) );
  XNOR U11874 ( .A(n10869), .B(n10867), .Z(n10871) );
  AND U11875 ( .A(n10872), .B(n10873), .Z(n10867) );
  NANDN U11876 ( .A(n10874), .B(n10875), .Z(n10873) );
  NANDN U11877 ( .A(n10876), .B(n10877), .Z(n10875) );
  AND U11878 ( .A(B[531]), .B(A[3]), .Z(n10869) );
  XNOR U11879 ( .A(n10859), .B(n10878), .Z(n10870) );
  XNOR U11880 ( .A(n10857), .B(n10860), .Z(n10878) );
  NAND U11881 ( .A(A[2]), .B(B[532]), .Z(n10860) );
  NANDN U11882 ( .A(n10879), .B(n10880), .Z(n10857) );
  AND U11883 ( .A(A[0]), .B(B[533]), .Z(n10880) );
  XOR U11884 ( .A(n10862), .B(n10881), .Z(n10859) );
  NAND U11885 ( .A(A[0]), .B(B[534]), .Z(n10881) );
  NAND U11886 ( .A(B[533]), .B(A[1]), .Z(n10862) );
  NAND U11887 ( .A(n10882), .B(n10883), .Z(n1067) );
  NANDN U11888 ( .A(n10884), .B(n10885), .Z(n10883) );
  OR U11889 ( .A(n10886), .B(n10887), .Z(n10885) );
  NAND U11890 ( .A(n10887), .B(n10886), .Z(n10882) );
  XOR U11891 ( .A(n1069), .B(n1068), .Z(\A1[531] ) );
  XOR U11892 ( .A(n10887), .B(n10888), .Z(n1068) );
  XNOR U11893 ( .A(n10886), .B(n10884), .Z(n10888) );
  AND U11894 ( .A(n10889), .B(n10890), .Z(n10884) );
  NANDN U11895 ( .A(n10891), .B(n10892), .Z(n10890) );
  NANDN U11896 ( .A(n10893), .B(n10894), .Z(n10892) );
  AND U11897 ( .A(B[530]), .B(A[3]), .Z(n10886) );
  XNOR U11898 ( .A(n10876), .B(n10895), .Z(n10887) );
  XNOR U11899 ( .A(n10874), .B(n10877), .Z(n10895) );
  NAND U11900 ( .A(A[2]), .B(B[531]), .Z(n10877) );
  NANDN U11901 ( .A(n10896), .B(n10897), .Z(n10874) );
  AND U11902 ( .A(A[0]), .B(B[532]), .Z(n10897) );
  XOR U11903 ( .A(n10879), .B(n10898), .Z(n10876) );
  NAND U11904 ( .A(A[0]), .B(B[533]), .Z(n10898) );
  NAND U11905 ( .A(B[532]), .B(A[1]), .Z(n10879) );
  NAND U11906 ( .A(n10899), .B(n10900), .Z(n1069) );
  NANDN U11907 ( .A(n10901), .B(n10902), .Z(n10900) );
  OR U11908 ( .A(n10903), .B(n10904), .Z(n10902) );
  NAND U11909 ( .A(n10904), .B(n10903), .Z(n10899) );
  XOR U11910 ( .A(n1071), .B(n1070), .Z(\A1[530] ) );
  XOR U11911 ( .A(n10904), .B(n10905), .Z(n1070) );
  XNOR U11912 ( .A(n10903), .B(n10901), .Z(n10905) );
  AND U11913 ( .A(n10906), .B(n10907), .Z(n10901) );
  NANDN U11914 ( .A(n10908), .B(n10909), .Z(n10907) );
  NANDN U11915 ( .A(n10910), .B(n10911), .Z(n10909) );
  AND U11916 ( .A(B[529]), .B(A[3]), .Z(n10903) );
  XNOR U11917 ( .A(n10893), .B(n10912), .Z(n10904) );
  XNOR U11918 ( .A(n10891), .B(n10894), .Z(n10912) );
  NAND U11919 ( .A(A[2]), .B(B[530]), .Z(n10894) );
  NANDN U11920 ( .A(n10913), .B(n10914), .Z(n10891) );
  AND U11921 ( .A(A[0]), .B(B[531]), .Z(n10914) );
  XOR U11922 ( .A(n10896), .B(n10915), .Z(n10893) );
  NAND U11923 ( .A(A[0]), .B(B[532]), .Z(n10915) );
  NAND U11924 ( .A(B[531]), .B(A[1]), .Z(n10896) );
  NAND U11925 ( .A(n10916), .B(n10917), .Z(n1071) );
  NANDN U11926 ( .A(n10918), .B(n10919), .Z(n10917) );
  OR U11927 ( .A(n10920), .B(n10921), .Z(n10919) );
  NAND U11928 ( .A(n10921), .B(n10920), .Z(n10916) );
  XOR U11929 ( .A(n1053), .B(n1052), .Z(\A1[52] ) );
  XOR U11930 ( .A(n10751), .B(n10922), .Z(n1052) );
  XNOR U11931 ( .A(n10750), .B(n10748), .Z(n10922) );
  AND U11932 ( .A(n10923), .B(n10924), .Z(n10748) );
  NANDN U11933 ( .A(n10925), .B(n10926), .Z(n10924) );
  NANDN U11934 ( .A(n10927), .B(n10928), .Z(n10926) );
  AND U11935 ( .A(B[51]), .B(A[3]), .Z(n10750) );
  XNOR U11936 ( .A(n10740), .B(n10929), .Z(n10751) );
  XNOR U11937 ( .A(n10738), .B(n10741), .Z(n10929) );
  NAND U11938 ( .A(A[2]), .B(B[52]), .Z(n10741) );
  NANDN U11939 ( .A(n10930), .B(n10931), .Z(n10738) );
  AND U11940 ( .A(A[0]), .B(B[53]), .Z(n10931) );
  XOR U11941 ( .A(n10743), .B(n10932), .Z(n10740) );
  NAND U11942 ( .A(A[0]), .B(B[54]), .Z(n10932) );
  NAND U11943 ( .A(B[53]), .B(A[1]), .Z(n10743) );
  NAND U11944 ( .A(n10933), .B(n10934), .Z(n1053) );
  NANDN U11945 ( .A(n10935), .B(n10936), .Z(n10934) );
  OR U11946 ( .A(n10937), .B(n10938), .Z(n10936) );
  NAND U11947 ( .A(n10938), .B(n10937), .Z(n10933) );
  XOR U11948 ( .A(n1073), .B(n1072), .Z(\A1[529] ) );
  XOR U11949 ( .A(n10921), .B(n10939), .Z(n1072) );
  XNOR U11950 ( .A(n10920), .B(n10918), .Z(n10939) );
  AND U11951 ( .A(n10940), .B(n10941), .Z(n10918) );
  NANDN U11952 ( .A(n10942), .B(n10943), .Z(n10941) );
  NANDN U11953 ( .A(n10944), .B(n10945), .Z(n10943) );
  AND U11954 ( .A(B[528]), .B(A[3]), .Z(n10920) );
  XNOR U11955 ( .A(n10910), .B(n10946), .Z(n10921) );
  XNOR U11956 ( .A(n10908), .B(n10911), .Z(n10946) );
  NAND U11957 ( .A(A[2]), .B(B[529]), .Z(n10911) );
  NANDN U11958 ( .A(n10947), .B(n10948), .Z(n10908) );
  AND U11959 ( .A(A[0]), .B(B[530]), .Z(n10948) );
  XOR U11960 ( .A(n10913), .B(n10949), .Z(n10910) );
  NAND U11961 ( .A(A[0]), .B(B[531]), .Z(n10949) );
  NAND U11962 ( .A(B[530]), .B(A[1]), .Z(n10913) );
  NAND U11963 ( .A(n10950), .B(n10951), .Z(n1073) );
  NANDN U11964 ( .A(n10952), .B(n10953), .Z(n10951) );
  OR U11965 ( .A(n10954), .B(n10955), .Z(n10953) );
  NAND U11966 ( .A(n10955), .B(n10954), .Z(n10950) );
  XOR U11967 ( .A(n1077), .B(n1076), .Z(\A1[528] ) );
  XOR U11968 ( .A(n10955), .B(n10956), .Z(n1076) );
  XNOR U11969 ( .A(n10954), .B(n10952), .Z(n10956) );
  AND U11970 ( .A(n10957), .B(n10958), .Z(n10952) );
  NANDN U11971 ( .A(n10959), .B(n10960), .Z(n10958) );
  NANDN U11972 ( .A(n10961), .B(n10962), .Z(n10960) );
  AND U11973 ( .A(B[527]), .B(A[3]), .Z(n10954) );
  XNOR U11974 ( .A(n10944), .B(n10963), .Z(n10955) );
  XNOR U11975 ( .A(n10942), .B(n10945), .Z(n10963) );
  NAND U11976 ( .A(A[2]), .B(B[528]), .Z(n10945) );
  NANDN U11977 ( .A(n10964), .B(n10965), .Z(n10942) );
  AND U11978 ( .A(A[0]), .B(B[529]), .Z(n10965) );
  XOR U11979 ( .A(n10947), .B(n10966), .Z(n10944) );
  NAND U11980 ( .A(A[0]), .B(B[530]), .Z(n10966) );
  NAND U11981 ( .A(B[529]), .B(A[1]), .Z(n10947) );
  NAND U11982 ( .A(n10967), .B(n10968), .Z(n1077) );
  NANDN U11983 ( .A(n10969), .B(n10970), .Z(n10968) );
  OR U11984 ( .A(n10971), .B(n10972), .Z(n10970) );
  NAND U11985 ( .A(n10972), .B(n10971), .Z(n10967) );
  XOR U11986 ( .A(n1079), .B(n1078), .Z(\A1[527] ) );
  XOR U11987 ( .A(n10972), .B(n10973), .Z(n1078) );
  XNOR U11988 ( .A(n10971), .B(n10969), .Z(n10973) );
  AND U11989 ( .A(n10974), .B(n10975), .Z(n10969) );
  NANDN U11990 ( .A(n10976), .B(n10977), .Z(n10975) );
  NANDN U11991 ( .A(n10978), .B(n10979), .Z(n10977) );
  AND U11992 ( .A(B[526]), .B(A[3]), .Z(n10971) );
  XNOR U11993 ( .A(n10961), .B(n10980), .Z(n10972) );
  XNOR U11994 ( .A(n10959), .B(n10962), .Z(n10980) );
  NAND U11995 ( .A(A[2]), .B(B[527]), .Z(n10962) );
  NANDN U11996 ( .A(n10981), .B(n10982), .Z(n10959) );
  AND U11997 ( .A(A[0]), .B(B[528]), .Z(n10982) );
  XOR U11998 ( .A(n10964), .B(n10983), .Z(n10961) );
  NAND U11999 ( .A(A[0]), .B(B[529]), .Z(n10983) );
  NAND U12000 ( .A(B[528]), .B(A[1]), .Z(n10964) );
  NAND U12001 ( .A(n10984), .B(n10985), .Z(n1079) );
  NANDN U12002 ( .A(n10986), .B(n10987), .Z(n10985) );
  OR U12003 ( .A(n10988), .B(n10989), .Z(n10987) );
  NAND U12004 ( .A(n10989), .B(n10988), .Z(n10984) );
  XOR U12005 ( .A(n1081), .B(n1080), .Z(\A1[526] ) );
  XOR U12006 ( .A(n10989), .B(n10990), .Z(n1080) );
  XNOR U12007 ( .A(n10988), .B(n10986), .Z(n10990) );
  AND U12008 ( .A(n10991), .B(n10992), .Z(n10986) );
  NANDN U12009 ( .A(n10993), .B(n10994), .Z(n10992) );
  NANDN U12010 ( .A(n10995), .B(n10996), .Z(n10994) );
  AND U12011 ( .A(B[525]), .B(A[3]), .Z(n10988) );
  XNOR U12012 ( .A(n10978), .B(n10997), .Z(n10989) );
  XNOR U12013 ( .A(n10976), .B(n10979), .Z(n10997) );
  NAND U12014 ( .A(A[2]), .B(B[526]), .Z(n10979) );
  NANDN U12015 ( .A(n10998), .B(n10999), .Z(n10976) );
  AND U12016 ( .A(A[0]), .B(B[527]), .Z(n10999) );
  XOR U12017 ( .A(n10981), .B(n11000), .Z(n10978) );
  NAND U12018 ( .A(A[0]), .B(B[528]), .Z(n11000) );
  NAND U12019 ( .A(B[527]), .B(A[1]), .Z(n10981) );
  NAND U12020 ( .A(n11001), .B(n11002), .Z(n1081) );
  NANDN U12021 ( .A(n11003), .B(n11004), .Z(n11002) );
  OR U12022 ( .A(n11005), .B(n11006), .Z(n11004) );
  NAND U12023 ( .A(n11006), .B(n11005), .Z(n11001) );
  XOR U12024 ( .A(n1083), .B(n1082), .Z(\A1[525] ) );
  XOR U12025 ( .A(n11006), .B(n11007), .Z(n1082) );
  XNOR U12026 ( .A(n11005), .B(n11003), .Z(n11007) );
  AND U12027 ( .A(n11008), .B(n11009), .Z(n11003) );
  NANDN U12028 ( .A(n11010), .B(n11011), .Z(n11009) );
  NANDN U12029 ( .A(n11012), .B(n11013), .Z(n11011) );
  AND U12030 ( .A(B[524]), .B(A[3]), .Z(n11005) );
  XNOR U12031 ( .A(n10995), .B(n11014), .Z(n11006) );
  XNOR U12032 ( .A(n10993), .B(n10996), .Z(n11014) );
  NAND U12033 ( .A(A[2]), .B(B[525]), .Z(n10996) );
  NANDN U12034 ( .A(n11015), .B(n11016), .Z(n10993) );
  AND U12035 ( .A(A[0]), .B(B[526]), .Z(n11016) );
  XOR U12036 ( .A(n10998), .B(n11017), .Z(n10995) );
  NAND U12037 ( .A(A[0]), .B(B[527]), .Z(n11017) );
  NAND U12038 ( .A(B[526]), .B(A[1]), .Z(n10998) );
  NAND U12039 ( .A(n11018), .B(n11019), .Z(n1083) );
  NANDN U12040 ( .A(n11020), .B(n11021), .Z(n11019) );
  OR U12041 ( .A(n11022), .B(n11023), .Z(n11021) );
  NAND U12042 ( .A(n11023), .B(n11022), .Z(n11018) );
  XOR U12043 ( .A(n1085), .B(n1084), .Z(\A1[524] ) );
  XOR U12044 ( .A(n11023), .B(n11024), .Z(n1084) );
  XNOR U12045 ( .A(n11022), .B(n11020), .Z(n11024) );
  AND U12046 ( .A(n11025), .B(n11026), .Z(n11020) );
  NANDN U12047 ( .A(n11027), .B(n11028), .Z(n11026) );
  NANDN U12048 ( .A(n11029), .B(n11030), .Z(n11028) );
  AND U12049 ( .A(B[523]), .B(A[3]), .Z(n11022) );
  XNOR U12050 ( .A(n11012), .B(n11031), .Z(n11023) );
  XNOR U12051 ( .A(n11010), .B(n11013), .Z(n11031) );
  NAND U12052 ( .A(A[2]), .B(B[524]), .Z(n11013) );
  NANDN U12053 ( .A(n11032), .B(n11033), .Z(n11010) );
  AND U12054 ( .A(A[0]), .B(B[525]), .Z(n11033) );
  XOR U12055 ( .A(n11015), .B(n11034), .Z(n11012) );
  NAND U12056 ( .A(A[0]), .B(B[526]), .Z(n11034) );
  NAND U12057 ( .A(B[525]), .B(A[1]), .Z(n11015) );
  NAND U12058 ( .A(n11035), .B(n11036), .Z(n1085) );
  NANDN U12059 ( .A(n11037), .B(n11038), .Z(n11036) );
  OR U12060 ( .A(n11039), .B(n11040), .Z(n11038) );
  NAND U12061 ( .A(n11040), .B(n11039), .Z(n11035) );
  XOR U12062 ( .A(n1087), .B(n1086), .Z(\A1[523] ) );
  XOR U12063 ( .A(n11040), .B(n11041), .Z(n1086) );
  XNOR U12064 ( .A(n11039), .B(n11037), .Z(n11041) );
  AND U12065 ( .A(n11042), .B(n11043), .Z(n11037) );
  NANDN U12066 ( .A(n11044), .B(n11045), .Z(n11043) );
  NANDN U12067 ( .A(n11046), .B(n11047), .Z(n11045) );
  AND U12068 ( .A(B[522]), .B(A[3]), .Z(n11039) );
  XNOR U12069 ( .A(n11029), .B(n11048), .Z(n11040) );
  XNOR U12070 ( .A(n11027), .B(n11030), .Z(n11048) );
  NAND U12071 ( .A(A[2]), .B(B[523]), .Z(n11030) );
  NANDN U12072 ( .A(n11049), .B(n11050), .Z(n11027) );
  AND U12073 ( .A(A[0]), .B(B[524]), .Z(n11050) );
  XOR U12074 ( .A(n11032), .B(n11051), .Z(n11029) );
  NAND U12075 ( .A(A[0]), .B(B[525]), .Z(n11051) );
  NAND U12076 ( .A(B[524]), .B(A[1]), .Z(n11032) );
  NAND U12077 ( .A(n11052), .B(n11053), .Z(n1087) );
  NANDN U12078 ( .A(n11054), .B(n11055), .Z(n11053) );
  OR U12079 ( .A(n11056), .B(n11057), .Z(n11055) );
  NAND U12080 ( .A(n11057), .B(n11056), .Z(n11052) );
  XOR U12081 ( .A(n1089), .B(n1088), .Z(\A1[522] ) );
  XOR U12082 ( .A(n11057), .B(n11058), .Z(n1088) );
  XNOR U12083 ( .A(n11056), .B(n11054), .Z(n11058) );
  AND U12084 ( .A(n11059), .B(n11060), .Z(n11054) );
  NANDN U12085 ( .A(n11061), .B(n11062), .Z(n11060) );
  NANDN U12086 ( .A(n11063), .B(n11064), .Z(n11062) );
  AND U12087 ( .A(B[521]), .B(A[3]), .Z(n11056) );
  XNOR U12088 ( .A(n11046), .B(n11065), .Z(n11057) );
  XNOR U12089 ( .A(n11044), .B(n11047), .Z(n11065) );
  NAND U12090 ( .A(A[2]), .B(B[522]), .Z(n11047) );
  NANDN U12091 ( .A(n11066), .B(n11067), .Z(n11044) );
  AND U12092 ( .A(A[0]), .B(B[523]), .Z(n11067) );
  XOR U12093 ( .A(n11049), .B(n11068), .Z(n11046) );
  NAND U12094 ( .A(A[0]), .B(B[524]), .Z(n11068) );
  NAND U12095 ( .A(B[523]), .B(A[1]), .Z(n11049) );
  NAND U12096 ( .A(n11069), .B(n11070), .Z(n1089) );
  NANDN U12097 ( .A(n11071), .B(n11072), .Z(n11070) );
  OR U12098 ( .A(n11073), .B(n11074), .Z(n11072) );
  NAND U12099 ( .A(n11074), .B(n11073), .Z(n11069) );
  XOR U12100 ( .A(n1091), .B(n1090), .Z(\A1[521] ) );
  XOR U12101 ( .A(n11074), .B(n11075), .Z(n1090) );
  XNOR U12102 ( .A(n11073), .B(n11071), .Z(n11075) );
  AND U12103 ( .A(n11076), .B(n11077), .Z(n11071) );
  NANDN U12104 ( .A(n11078), .B(n11079), .Z(n11077) );
  NANDN U12105 ( .A(n11080), .B(n11081), .Z(n11079) );
  AND U12106 ( .A(B[520]), .B(A[3]), .Z(n11073) );
  XNOR U12107 ( .A(n11063), .B(n11082), .Z(n11074) );
  XNOR U12108 ( .A(n11061), .B(n11064), .Z(n11082) );
  NAND U12109 ( .A(A[2]), .B(B[521]), .Z(n11064) );
  NANDN U12110 ( .A(n11083), .B(n11084), .Z(n11061) );
  AND U12111 ( .A(A[0]), .B(B[522]), .Z(n11084) );
  XOR U12112 ( .A(n11066), .B(n11085), .Z(n11063) );
  NAND U12113 ( .A(A[0]), .B(B[523]), .Z(n11085) );
  NAND U12114 ( .A(B[522]), .B(A[1]), .Z(n11066) );
  NAND U12115 ( .A(n11086), .B(n11087), .Z(n1091) );
  NANDN U12116 ( .A(n11088), .B(n11089), .Z(n11087) );
  OR U12117 ( .A(n11090), .B(n11091), .Z(n11089) );
  NAND U12118 ( .A(n11091), .B(n11090), .Z(n11086) );
  XOR U12119 ( .A(n1093), .B(n1092), .Z(\A1[520] ) );
  XOR U12120 ( .A(n11091), .B(n11092), .Z(n1092) );
  XNOR U12121 ( .A(n11090), .B(n11088), .Z(n11092) );
  AND U12122 ( .A(n11093), .B(n11094), .Z(n11088) );
  NANDN U12123 ( .A(n11095), .B(n11096), .Z(n11094) );
  NANDN U12124 ( .A(n11097), .B(n11098), .Z(n11096) );
  AND U12125 ( .A(B[519]), .B(A[3]), .Z(n11090) );
  XNOR U12126 ( .A(n11080), .B(n11099), .Z(n11091) );
  XNOR U12127 ( .A(n11078), .B(n11081), .Z(n11099) );
  NAND U12128 ( .A(A[2]), .B(B[520]), .Z(n11081) );
  NANDN U12129 ( .A(n11100), .B(n11101), .Z(n11078) );
  AND U12130 ( .A(A[0]), .B(B[521]), .Z(n11101) );
  XOR U12131 ( .A(n11083), .B(n11102), .Z(n11080) );
  NAND U12132 ( .A(A[0]), .B(B[522]), .Z(n11102) );
  NAND U12133 ( .A(B[521]), .B(A[1]), .Z(n11083) );
  NAND U12134 ( .A(n11103), .B(n11104), .Z(n1093) );
  NANDN U12135 ( .A(n11105), .B(n11106), .Z(n11104) );
  OR U12136 ( .A(n11107), .B(n11108), .Z(n11106) );
  NAND U12137 ( .A(n11108), .B(n11107), .Z(n11103) );
  XOR U12138 ( .A(n1075), .B(n1074), .Z(\A1[51] ) );
  XOR U12139 ( .A(n10938), .B(n11109), .Z(n1074) );
  XNOR U12140 ( .A(n10937), .B(n10935), .Z(n11109) );
  AND U12141 ( .A(n11110), .B(n11111), .Z(n10935) );
  NANDN U12142 ( .A(n11112), .B(n11113), .Z(n11111) );
  NANDN U12143 ( .A(n11114), .B(n11115), .Z(n11113) );
  AND U12144 ( .A(B[50]), .B(A[3]), .Z(n10937) );
  XNOR U12145 ( .A(n10927), .B(n11116), .Z(n10938) );
  XNOR U12146 ( .A(n10925), .B(n10928), .Z(n11116) );
  NAND U12147 ( .A(A[2]), .B(B[51]), .Z(n10928) );
  NANDN U12148 ( .A(n11117), .B(n11118), .Z(n10925) );
  AND U12149 ( .A(A[0]), .B(B[52]), .Z(n11118) );
  XOR U12150 ( .A(n10930), .B(n11119), .Z(n10927) );
  NAND U12151 ( .A(A[0]), .B(B[53]), .Z(n11119) );
  NAND U12152 ( .A(B[52]), .B(A[1]), .Z(n10930) );
  NAND U12153 ( .A(n11120), .B(n11121), .Z(n1075) );
  NANDN U12154 ( .A(n11122), .B(n11123), .Z(n11121) );
  OR U12155 ( .A(n11124), .B(n11125), .Z(n11123) );
  NAND U12156 ( .A(n11125), .B(n11124), .Z(n11120) );
  XOR U12157 ( .A(n1095), .B(n1094), .Z(\A1[519] ) );
  XOR U12158 ( .A(n11108), .B(n11126), .Z(n1094) );
  XNOR U12159 ( .A(n11107), .B(n11105), .Z(n11126) );
  AND U12160 ( .A(n11127), .B(n11128), .Z(n11105) );
  NANDN U12161 ( .A(n11129), .B(n11130), .Z(n11128) );
  NANDN U12162 ( .A(n11131), .B(n11132), .Z(n11130) );
  AND U12163 ( .A(B[518]), .B(A[3]), .Z(n11107) );
  XNOR U12164 ( .A(n11097), .B(n11133), .Z(n11108) );
  XNOR U12165 ( .A(n11095), .B(n11098), .Z(n11133) );
  NAND U12166 ( .A(A[2]), .B(B[519]), .Z(n11098) );
  NANDN U12167 ( .A(n11134), .B(n11135), .Z(n11095) );
  AND U12168 ( .A(A[0]), .B(B[520]), .Z(n11135) );
  XOR U12169 ( .A(n11100), .B(n11136), .Z(n11097) );
  NAND U12170 ( .A(A[0]), .B(B[521]), .Z(n11136) );
  NAND U12171 ( .A(B[520]), .B(A[1]), .Z(n11100) );
  NAND U12172 ( .A(n11137), .B(n11138), .Z(n1095) );
  NANDN U12173 ( .A(n11139), .B(n11140), .Z(n11138) );
  OR U12174 ( .A(n11141), .B(n11142), .Z(n11140) );
  NAND U12175 ( .A(n11142), .B(n11141), .Z(n11137) );
  XOR U12176 ( .A(n1099), .B(n1098), .Z(\A1[518] ) );
  XOR U12177 ( .A(n11142), .B(n11143), .Z(n1098) );
  XNOR U12178 ( .A(n11141), .B(n11139), .Z(n11143) );
  AND U12179 ( .A(n11144), .B(n11145), .Z(n11139) );
  NANDN U12180 ( .A(n11146), .B(n11147), .Z(n11145) );
  NANDN U12181 ( .A(n11148), .B(n11149), .Z(n11147) );
  AND U12182 ( .A(B[517]), .B(A[3]), .Z(n11141) );
  XNOR U12183 ( .A(n11131), .B(n11150), .Z(n11142) );
  XNOR U12184 ( .A(n11129), .B(n11132), .Z(n11150) );
  NAND U12185 ( .A(A[2]), .B(B[518]), .Z(n11132) );
  NANDN U12186 ( .A(n11151), .B(n11152), .Z(n11129) );
  AND U12187 ( .A(A[0]), .B(B[519]), .Z(n11152) );
  XOR U12188 ( .A(n11134), .B(n11153), .Z(n11131) );
  NAND U12189 ( .A(A[0]), .B(B[520]), .Z(n11153) );
  NAND U12190 ( .A(B[519]), .B(A[1]), .Z(n11134) );
  NAND U12191 ( .A(n11154), .B(n11155), .Z(n1099) );
  NANDN U12192 ( .A(n11156), .B(n11157), .Z(n11155) );
  OR U12193 ( .A(n11158), .B(n11159), .Z(n11157) );
  NAND U12194 ( .A(n11159), .B(n11158), .Z(n11154) );
  XOR U12195 ( .A(n1101), .B(n1100), .Z(\A1[517] ) );
  XOR U12196 ( .A(n11159), .B(n11160), .Z(n1100) );
  XNOR U12197 ( .A(n11158), .B(n11156), .Z(n11160) );
  AND U12198 ( .A(n11161), .B(n11162), .Z(n11156) );
  NANDN U12199 ( .A(n11163), .B(n11164), .Z(n11162) );
  NANDN U12200 ( .A(n11165), .B(n11166), .Z(n11164) );
  AND U12201 ( .A(B[516]), .B(A[3]), .Z(n11158) );
  XNOR U12202 ( .A(n11148), .B(n11167), .Z(n11159) );
  XNOR U12203 ( .A(n11146), .B(n11149), .Z(n11167) );
  NAND U12204 ( .A(A[2]), .B(B[517]), .Z(n11149) );
  NANDN U12205 ( .A(n11168), .B(n11169), .Z(n11146) );
  AND U12206 ( .A(A[0]), .B(B[518]), .Z(n11169) );
  XOR U12207 ( .A(n11151), .B(n11170), .Z(n11148) );
  NAND U12208 ( .A(A[0]), .B(B[519]), .Z(n11170) );
  NAND U12209 ( .A(B[518]), .B(A[1]), .Z(n11151) );
  NAND U12210 ( .A(n11171), .B(n11172), .Z(n1101) );
  NANDN U12211 ( .A(n11173), .B(n11174), .Z(n11172) );
  OR U12212 ( .A(n11175), .B(n11176), .Z(n11174) );
  NAND U12213 ( .A(n11176), .B(n11175), .Z(n11171) );
  XOR U12214 ( .A(n1103), .B(n1102), .Z(\A1[516] ) );
  XOR U12215 ( .A(n11176), .B(n11177), .Z(n1102) );
  XNOR U12216 ( .A(n11175), .B(n11173), .Z(n11177) );
  AND U12217 ( .A(n11178), .B(n11179), .Z(n11173) );
  NANDN U12218 ( .A(n11180), .B(n11181), .Z(n11179) );
  NANDN U12219 ( .A(n11182), .B(n11183), .Z(n11181) );
  AND U12220 ( .A(B[515]), .B(A[3]), .Z(n11175) );
  XNOR U12221 ( .A(n11165), .B(n11184), .Z(n11176) );
  XNOR U12222 ( .A(n11163), .B(n11166), .Z(n11184) );
  NAND U12223 ( .A(A[2]), .B(B[516]), .Z(n11166) );
  NANDN U12224 ( .A(n11185), .B(n11186), .Z(n11163) );
  AND U12225 ( .A(A[0]), .B(B[517]), .Z(n11186) );
  XOR U12226 ( .A(n11168), .B(n11187), .Z(n11165) );
  NAND U12227 ( .A(A[0]), .B(B[518]), .Z(n11187) );
  NAND U12228 ( .A(B[517]), .B(A[1]), .Z(n11168) );
  NAND U12229 ( .A(n11188), .B(n11189), .Z(n1103) );
  NANDN U12230 ( .A(n11190), .B(n11191), .Z(n11189) );
  OR U12231 ( .A(n11192), .B(n11193), .Z(n11191) );
  NAND U12232 ( .A(n11193), .B(n11192), .Z(n11188) );
  XOR U12233 ( .A(n1105), .B(n1104), .Z(\A1[515] ) );
  XOR U12234 ( .A(n11193), .B(n11194), .Z(n1104) );
  XNOR U12235 ( .A(n11192), .B(n11190), .Z(n11194) );
  AND U12236 ( .A(n11195), .B(n11196), .Z(n11190) );
  NANDN U12237 ( .A(n11197), .B(n11198), .Z(n11196) );
  NANDN U12238 ( .A(n11199), .B(n11200), .Z(n11198) );
  AND U12239 ( .A(B[514]), .B(A[3]), .Z(n11192) );
  XNOR U12240 ( .A(n11182), .B(n11201), .Z(n11193) );
  XNOR U12241 ( .A(n11180), .B(n11183), .Z(n11201) );
  NAND U12242 ( .A(A[2]), .B(B[515]), .Z(n11183) );
  NANDN U12243 ( .A(n11202), .B(n11203), .Z(n11180) );
  AND U12244 ( .A(A[0]), .B(B[516]), .Z(n11203) );
  XOR U12245 ( .A(n11185), .B(n11204), .Z(n11182) );
  NAND U12246 ( .A(A[0]), .B(B[517]), .Z(n11204) );
  NAND U12247 ( .A(B[516]), .B(A[1]), .Z(n11185) );
  NAND U12248 ( .A(n11205), .B(n11206), .Z(n1105) );
  NANDN U12249 ( .A(n11207), .B(n11208), .Z(n11206) );
  OR U12250 ( .A(n11209), .B(n11210), .Z(n11208) );
  NAND U12251 ( .A(n11210), .B(n11209), .Z(n11205) );
  XOR U12252 ( .A(n1107), .B(n1106), .Z(\A1[514] ) );
  XOR U12253 ( .A(n11210), .B(n11211), .Z(n1106) );
  XNOR U12254 ( .A(n11209), .B(n11207), .Z(n11211) );
  AND U12255 ( .A(n11212), .B(n11213), .Z(n11207) );
  NANDN U12256 ( .A(n11214), .B(n11215), .Z(n11213) );
  NANDN U12257 ( .A(n11216), .B(n11217), .Z(n11215) );
  AND U12258 ( .A(B[513]), .B(A[3]), .Z(n11209) );
  XNOR U12259 ( .A(n11199), .B(n11218), .Z(n11210) );
  XNOR U12260 ( .A(n11197), .B(n11200), .Z(n11218) );
  NAND U12261 ( .A(A[2]), .B(B[514]), .Z(n11200) );
  NANDN U12262 ( .A(n11219), .B(n11220), .Z(n11197) );
  AND U12263 ( .A(A[0]), .B(B[515]), .Z(n11220) );
  XOR U12264 ( .A(n11202), .B(n11221), .Z(n11199) );
  NAND U12265 ( .A(A[0]), .B(B[516]), .Z(n11221) );
  NAND U12266 ( .A(B[515]), .B(A[1]), .Z(n11202) );
  NAND U12267 ( .A(n11222), .B(n11223), .Z(n1107) );
  NANDN U12268 ( .A(n11224), .B(n11225), .Z(n11223) );
  OR U12269 ( .A(n11226), .B(n11227), .Z(n11225) );
  NAND U12270 ( .A(n11227), .B(n11226), .Z(n11222) );
  XOR U12271 ( .A(n1109), .B(n1108), .Z(\A1[513] ) );
  XOR U12272 ( .A(n11227), .B(n11228), .Z(n1108) );
  XNOR U12273 ( .A(n11226), .B(n11224), .Z(n11228) );
  AND U12274 ( .A(n11229), .B(n11230), .Z(n11224) );
  NANDN U12275 ( .A(n11231), .B(n11232), .Z(n11230) );
  NANDN U12276 ( .A(n11233), .B(n11234), .Z(n11232) );
  AND U12277 ( .A(B[512]), .B(A[3]), .Z(n11226) );
  XNOR U12278 ( .A(n11216), .B(n11235), .Z(n11227) );
  XNOR U12279 ( .A(n11214), .B(n11217), .Z(n11235) );
  NAND U12280 ( .A(A[2]), .B(B[513]), .Z(n11217) );
  NANDN U12281 ( .A(n11236), .B(n11237), .Z(n11214) );
  AND U12282 ( .A(A[0]), .B(B[514]), .Z(n11237) );
  XOR U12283 ( .A(n11219), .B(n11238), .Z(n11216) );
  NAND U12284 ( .A(A[0]), .B(B[515]), .Z(n11238) );
  NAND U12285 ( .A(B[514]), .B(A[1]), .Z(n11219) );
  NAND U12286 ( .A(n11239), .B(n11240), .Z(n1109) );
  NANDN U12287 ( .A(n11241), .B(n11242), .Z(n11240) );
  OR U12288 ( .A(n11243), .B(n11244), .Z(n11242) );
  NAND U12289 ( .A(n11244), .B(n11243), .Z(n11239) );
  XOR U12290 ( .A(n1111), .B(n1110), .Z(\A1[512] ) );
  XOR U12291 ( .A(n11244), .B(n11245), .Z(n1110) );
  XNOR U12292 ( .A(n11243), .B(n11241), .Z(n11245) );
  AND U12293 ( .A(n11246), .B(n11247), .Z(n11241) );
  NANDN U12294 ( .A(n11248), .B(n11249), .Z(n11247) );
  NANDN U12295 ( .A(n11250), .B(n11251), .Z(n11249) );
  AND U12296 ( .A(B[511]), .B(A[3]), .Z(n11243) );
  XNOR U12297 ( .A(n11233), .B(n11252), .Z(n11244) );
  XNOR U12298 ( .A(n11231), .B(n11234), .Z(n11252) );
  NAND U12299 ( .A(A[2]), .B(B[512]), .Z(n11234) );
  NANDN U12300 ( .A(n11253), .B(n11254), .Z(n11231) );
  AND U12301 ( .A(A[0]), .B(B[513]), .Z(n11254) );
  XOR U12302 ( .A(n11236), .B(n11255), .Z(n11233) );
  NAND U12303 ( .A(A[0]), .B(B[514]), .Z(n11255) );
  NAND U12304 ( .A(B[513]), .B(A[1]), .Z(n11236) );
  NAND U12305 ( .A(n11256), .B(n11257), .Z(n1111) );
  NANDN U12306 ( .A(n11258), .B(n11259), .Z(n11257) );
  OR U12307 ( .A(n11260), .B(n11261), .Z(n11259) );
  NAND U12308 ( .A(n11261), .B(n11260), .Z(n11256) );
  XOR U12309 ( .A(n1113), .B(n1112), .Z(\A1[511] ) );
  XOR U12310 ( .A(n11261), .B(n11262), .Z(n1112) );
  XNOR U12311 ( .A(n11260), .B(n11258), .Z(n11262) );
  AND U12312 ( .A(n11263), .B(n11264), .Z(n11258) );
  NANDN U12313 ( .A(n11265), .B(n11266), .Z(n11264) );
  NANDN U12314 ( .A(n11267), .B(n11268), .Z(n11266) );
  AND U12315 ( .A(B[510]), .B(A[3]), .Z(n11260) );
  XNOR U12316 ( .A(n11250), .B(n11269), .Z(n11261) );
  XNOR U12317 ( .A(n11248), .B(n11251), .Z(n11269) );
  NAND U12318 ( .A(A[2]), .B(B[511]), .Z(n11251) );
  NANDN U12319 ( .A(n11270), .B(n11271), .Z(n11248) );
  AND U12320 ( .A(A[0]), .B(B[512]), .Z(n11271) );
  XOR U12321 ( .A(n11253), .B(n11272), .Z(n11250) );
  NAND U12322 ( .A(A[0]), .B(B[513]), .Z(n11272) );
  NAND U12323 ( .A(B[512]), .B(A[1]), .Z(n11253) );
  NAND U12324 ( .A(n11273), .B(n11274), .Z(n1113) );
  NANDN U12325 ( .A(n11275), .B(n11276), .Z(n11274) );
  OR U12326 ( .A(n11277), .B(n11278), .Z(n11276) );
  NAND U12327 ( .A(n11278), .B(n11277), .Z(n11273) );
  XOR U12328 ( .A(n1115), .B(n1114), .Z(\A1[510] ) );
  XOR U12329 ( .A(n11278), .B(n11279), .Z(n1114) );
  XNOR U12330 ( .A(n11277), .B(n11275), .Z(n11279) );
  AND U12331 ( .A(n11280), .B(n11281), .Z(n11275) );
  NANDN U12332 ( .A(n11282), .B(n11283), .Z(n11281) );
  NANDN U12333 ( .A(n11284), .B(n11285), .Z(n11283) );
  AND U12334 ( .A(B[509]), .B(A[3]), .Z(n11277) );
  XNOR U12335 ( .A(n11267), .B(n11286), .Z(n11278) );
  XNOR U12336 ( .A(n11265), .B(n11268), .Z(n11286) );
  NAND U12337 ( .A(A[2]), .B(B[510]), .Z(n11268) );
  NANDN U12338 ( .A(n11287), .B(n11288), .Z(n11265) );
  AND U12339 ( .A(A[0]), .B(B[511]), .Z(n11288) );
  XOR U12340 ( .A(n11270), .B(n11289), .Z(n11267) );
  NAND U12341 ( .A(A[0]), .B(B[512]), .Z(n11289) );
  NAND U12342 ( .A(B[511]), .B(A[1]), .Z(n11270) );
  NAND U12343 ( .A(n11290), .B(n11291), .Z(n1115) );
  NANDN U12344 ( .A(n11292), .B(n11293), .Z(n11291) );
  OR U12345 ( .A(n11294), .B(n11295), .Z(n11293) );
  NAND U12346 ( .A(n11295), .B(n11294), .Z(n11290) );
  XOR U12347 ( .A(n1097), .B(n1096), .Z(\A1[50] ) );
  XOR U12348 ( .A(n11125), .B(n11296), .Z(n1096) );
  XNOR U12349 ( .A(n11124), .B(n11122), .Z(n11296) );
  AND U12350 ( .A(n11297), .B(n11298), .Z(n11122) );
  NANDN U12351 ( .A(n11299), .B(n11300), .Z(n11298) );
  NANDN U12352 ( .A(n11301), .B(n11302), .Z(n11300) );
  AND U12353 ( .A(B[49]), .B(A[3]), .Z(n11124) );
  XNOR U12354 ( .A(n11114), .B(n11303), .Z(n11125) );
  XNOR U12355 ( .A(n11112), .B(n11115), .Z(n11303) );
  NAND U12356 ( .A(A[2]), .B(B[50]), .Z(n11115) );
  NANDN U12357 ( .A(n11304), .B(n11305), .Z(n11112) );
  AND U12358 ( .A(A[0]), .B(B[51]), .Z(n11305) );
  XOR U12359 ( .A(n11117), .B(n11306), .Z(n11114) );
  NAND U12360 ( .A(A[0]), .B(B[52]), .Z(n11306) );
  NAND U12361 ( .A(B[51]), .B(A[1]), .Z(n11117) );
  NAND U12362 ( .A(n11307), .B(n11308), .Z(n1097) );
  NANDN U12363 ( .A(n11309), .B(n11310), .Z(n11308) );
  OR U12364 ( .A(n11311), .B(n11312), .Z(n11310) );
  NAND U12365 ( .A(n11312), .B(n11311), .Z(n11307) );
  XOR U12366 ( .A(n1117), .B(n1116), .Z(\A1[509] ) );
  XOR U12367 ( .A(n11295), .B(n11313), .Z(n1116) );
  XNOR U12368 ( .A(n11294), .B(n11292), .Z(n11313) );
  AND U12369 ( .A(n11314), .B(n11315), .Z(n11292) );
  NANDN U12370 ( .A(n11316), .B(n11317), .Z(n11315) );
  NANDN U12371 ( .A(n11318), .B(n11319), .Z(n11317) );
  AND U12372 ( .A(B[508]), .B(A[3]), .Z(n11294) );
  XNOR U12373 ( .A(n11284), .B(n11320), .Z(n11295) );
  XNOR U12374 ( .A(n11282), .B(n11285), .Z(n11320) );
  NAND U12375 ( .A(A[2]), .B(B[509]), .Z(n11285) );
  NANDN U12376 ( .A(n11321), .B(n11322), .Z(n11282) );
  AND U12377 ( .A(A[0]), .B(B[510]), .Z(n11322) );
  XOR U12378 ( .A(n11287), .B(n11323), .Z(n11284) );
  NAND U12379 ( .A(A[0]), .B(B[511]), .Z(n11323) );
  NAND U12380 ( .A(B[510]), .B(A[1]), .Z(n11287) );
  NAND U12381 ( .A(n11324), .B(n11325), .Z(n1117) );
  NANDN U12382 ( .A(n11326), .B(n11327), .Z(n11325) );
  OR U12383 ( .A(n11328), .B(n11329), .Z(n11327) );
  NAND U12384 ( .A(n11329), .B(n11328), .Z(n11324) );
  XOR U12385 ( .A(n1121), .B(n1120), .Z(\A1[508] ) );
  XOR U12386 ( .A(n11329), .B(n11330), .Z(n1120) );
  XNOR U12387 ( .A(n11328), .B(n11326), .Z(n11330) );
  AND U12388 ( .A(n11331), .B(n11332), .Z(n11326) );
  NANDN U12389 ( .A(n11333), .B(n11334), .Z(n11332) );
  NANDN U12390 ( .A(n11335), .B(n11336), .Z(n11334) );
  AND U12391 ( .A(B[507]), .B(A[3]), .Z(n11328) );
  XNOR U12392 ( .A(n11318), .B(n11337), .Z(n11329) );
  XNOR U12393 ( .A(n11316), .B(n11319), .Z(n11337) );
  NAND U12394 ( .A(A[2]), .B(B[508]), .Z(n11319) );
  NANDN U12395 ( .A(n11338), .B(n11339), .Z(n11316) );
  AND U12396 ( .A(A[0]), .B(B[509]), .Z(n11339) );
  XOR U12397 ( .A(n11321), .B(n11340), .Z(n11318) );
  NAND U12398 ( .A(A[0]), .B(B[510]), .Z(n11340) );
  NAND U12399 ( .A(B[509]), .B(A[1]), .Z(n11321) );
  NAND U12400 ( .A(n11341), .B(n11342), .Z(n1121) );
  NANDN U12401 ( .A(n11343), .B(n11344), .Z(n11342) );
  OR U12402 ( .A(n11345), .B(n11346), .Z(n11344) );
  NAND U12403 ( .A(n11346), .B(n11345), .Z(n11341) );
  XOR U12404 ( .A(n1123), .B(n1122), .Z(\A1[507] ) );
  XOR U12405 ( .A(n11346), .B(n11347), .Z(n1122) );
  XNOR U12406 ( .A(n11345), .B(n11343), .Z(n11347) );
  AND U12407 ( .A(n11348), .B(n11349), .Z(n11343) );
  NANDN U12408 ( .A(n11350), .B(n11351), .Z(n11349) );
  NANDN U12409 ( .A(n11352), .B(n11353), .Z(n11351) );
  AND U12410 ( .A(B[506]), .B(A[3]), .Z(n11345) );
  XNOR U12411 ( .A(n11335), .B(n11354), .Z(n11346) );
  XNOR U12412 ( .A(n11333), .B(n11336), .Z(n11354) );
  NAND U12413 ( .A(A[2]), .B(B[507]), .Z(n11336) );
  NANDN U12414 ( .A(n11355), .B(n11356), .Z(n11333) );
  AND U12415 ( .A(A[0]), .B(B[508]), .Z(n11356) );
  XOR U12416 ( .A(n11338), .B(n11357), .Z(n11335) );
  NAND U12417 ( .A(A[0]), .B(B[509]), .Z(n11357) );
  NAND U12418 ( .A(B[508]), .B(A[1]), .Z(n11338) );
  NAND U12419 ( .A(n11358), .B(n11359), .Z(n1123) );
  NANDN U12420 ( .A(n11360), .B(n11361), .Z(n11359) );
  OR U12421 ( .A(n11362), .B(n11363), .Z(n11361) );
  NAND U12422 ( .A(n11363), .B(n11362), .Z(n11358) );
  XOR U12423 ( .A(n1125), .B(n1124), .Z(\A1[506] ) );
  XOR U12424 ( .A(n11363), .B(n11364), .Z(n1124) );
  XNOR U12425 ( .A(n11362), .B(n11360), .Z(n11364) );
  AND U12426 ( .A(n11365), .B(n11366), .Z(n11360) );
  NANDN U12427 ( .A(n11367), .B(n11368), .Z(n11366) );
  NANDN U12428 ( .A(n11369), .B(n11370), .Z(n11368) );
  AND U12429 ( .A(B[505]), .B(A[3]), .Z(n11362) );
  XNOR U12430 ( .A(n11352), .B(n11371), .Z(n11363) );
  XNOR U12431 ( .A(n11350), .B(n11353), .Z(n11371) );
  NAND U12432 ( .A(A[2]), .B(B[506]), .Z(n11353) );
  NANDN U12433 ( .A(n11372), .B(n11373), .Z(n11350) );
  AND U12434 ( .A(A[0]), .B(B[507]), .Z(n11373) );
  XOR U12435 ( .A(n11355), .B(n11374), .Z(n11352) );
  NAND U12436 ( .A(A[0]), .B(B[508]), .Z(n11374) );
  NAND U12437 ( .A(B[507]), .B(A[1]), .Z(n11355) );
  NAND U12438 ( .A(n11375), .B(n11376), .Z(n1125) );
  NANDN U12439 ( .A(n11377), .B(n11378), .Z(n11376) );
  OR U12440 ( .A(n11379), .B(n11380), .Z(n11378) );
  NAND U12441 ( .A(n11380), .B(n11379), .Z(n11375) );
  XOR U12442 ( .A(n1127), .B(n1126), .Z(\A1[505] ) );
  XOR U12443 ( .A(n11380), .B(n11381), .Z(n1126) );
  XNOR U12444 ( .A(n11379), .B(n11377), .Z(n11381) );
  AND U12445 ( .A(n11382), .B(n11383), .Z(n11377) );
  NANDN U12446 ( .A(n11384), .B(n11385), .Z(n11383) );
  NANDN U12447 ( .A(n11386), .B(n11387), .Z(n11385) );
  AND U12448 ( .A(B[504]), .B(A[3]), .Z(n11379) );
  XNOR U12449 ( .A(n11369), .B(n11388), .Z(n11380) );
  XNOR U12450 ( .A(n11367), .B(n11370), .Z(n11388) );
  NAND U12451 ( .A(A[2]), .B(B[505]), .Z(n11370) );
  NANDN U12452 ( .A(n11389), .B(n11390), .Z(n11367) );
  AND U12453 ( .A(A[0]), .B(B[506]), .Z(n11390) );
  XOR U12454 ( .A(n11372), .B(n11391), .Z(n11369) );
  NAND U12455 ( .A(A[0]), .B(B[507]), .Z(n11391) );
  NAND U12456 ( .A(B[506]), .B(A[1]), .Z(n11372) );
  NAND U12457 ( .A(n11392), .B(n11393), .Z(n1127) );
  NANDN U12458 ( .A(n11394), .B(n11395), .Z(n11393) );
  OR U12459 ( .A(n11396), .B(n11397), .Z(n11395) );
  NAND U12460 ( .A(n11397), .B(n11396), .Z(n11392) );
  XOR U12461 ( .A(n1129), .B(n1128), .Z(\A1[504] ) );
  XOR U12462 ( .A(n11397), .B(n11398), .Z(n1128) );
  XNOR U12463 ( .A(n11396), .B(n11394), .Z(n11398) );
  AND U12464 ( .A(n11399), .B(n11400), .Z(n11394) );
  NANDN U12465 ( .A(n11401), .B(n11402), .Z(n11400) );
  NANDN U12466 ( .A(n11403), .B(n11404), .Z(n11402) );
  AND U12467 ( .A(B[503]), .B(A[3]), .Z(n11396) );
  XNOR U12468 ( .A(n11386), .B(n11405), .Z(n11397) );
  XNOR U12469 ( .A(n11384), .B(n11387), .Z(n11405) );
  NAND U12470 ( .A(A[2]), .B(B[504]), .Z(n11387) );
  NANDN U12471 ( .A(n11406), .B(n11407), .Z(n11384) );
  AND U12472 ( .A(A[0]), .B(B[505]), .Z(n11407) );
  XOR U12473 ( .A(n11389), .B(n11408), .Z(n11386) );
  NAND U12474 ( .A(A[0]), .B(B[506]), .Z(n11408) );
  NAND U12475 ( .A(B[505]), .B(A[1]), .Z(n11389) );
  NAND U12476 ( .A(n11409), .B(n11410), .Z(n1129) );
  NANDN U12477 ( .A(n11411), .B(n11412), .Z(n11410) );
  OR U12478 ( .A(n11413), .B(n11414), .Z(n11412) );
  NAND U12479 ( .A(n11414), .B(n11413), .Z(n11409) );
  XOR U12480 ( .A(n1131), .B(n1130), .Z(\A1[503] ) );
  XOR U12481 ( .A(n11414), .B(n11415), .Z(n1130) );
  XNOR U12482 ( .A(n11413), .B(n11411), .Z(n11415) );
  AND U12483 ( .A(n11416), .B(n11417), .Z(n11411) );
  NANDN U12484 ( .A(n11418), .B(n11419), .Z(n11417) );
  NANDN U12485 ( .A(n11420), .B(n11421), .Z(n11419) );
  AND U12486 ( .A(B[502]), .B(A[3]), .Z(n11413) );
  XNOR U12487 ( .A(n11403), .B(n11422), .Z(n11414) );
  XNOR U12488 ( .A(n11401), .B(n11404), .Z(n11422) );
  NAND U12489 ( .A(A[2]), .B(B[503]), .Z(n11404) );
  NANDN U12490 ( .A(n11423), .B(n11424), .Z(n11401) );
  AND U12491 ( .A(A[0]), .B(B[504]), .Z(n11424) );
  XOR U12492 ( .A(n11406), .B(n11425), .Z(n11403) );
  NAND U12493 ( .A(A[0]), .B(B[505]), .Z(n11425) );
  NAND U12494 ( .A(B[504]), .B(A[1]), .Z(n11406) );
  NAND U12495 ( .A(n11426), .B(n11427), .Z(n1131) );
  NANDN U12496 ( .A(n11428), .B(n11429), .Z(n11427) );
  OR U12497 ( .A(n11430), .B(n11431), .Z(n11429) );
  NAND U12498 ( .A(n11431), .B(n11430), .Z(n11426) );
  XOR U12499 ( .A(n1133), .B(n1132), .Z(\A1[502] ) );
  XOR U12500 ( .A(n11431), .B(n11432), .Z(n1132) );
  XNOR U12501 ( .A(n11430), .B(n11428), .Z(n11432) );
  AND U12502 ( .A(n11433), .B(n11434), .Z(n11428) );
  NANDN U12503 ( .A(n11435), .B(n11436), .Z(n11434) );
  NANDN U12504 ( .A(n11437), .B(n11438), .Z(n11436) );
  AND U12505 ( .A(B[501]), .B(A[3]), .Z(n11430) );
  XNOR U12506 ( .A(n11420), .B(n11439), .Z(n11431) );
  XNOR U12507 ( .A(n11418), .B(n11421), .Z(n11439) );
  NAND U12508 ( .A(A[2]), .B(B[502]), .Z(n11421) );
  NANDN U12509 ( .A(n11440), .B(n11441), .Z(n11418) );
  AND U12510 ( .A(A[0]), .B(B[503]), .Z(n11441) );
  XOR U12511 ( .A(n11423), .B(n11442), .Z(n11420) );
  NAND U12512 ( .A(A[0]), .B(B[504]), .Z(n11442) );
  NAND U12513 ( .A(B[503]), .B(A[1]), .Z(n11423) );
  NAND U12514 ( .A(n11443), .B(n11444), .Z(n1133) );
  NANDN U12515 ( .A(n11445), .B(n11446), .Z(n11444) );
  OR U12516 ( .A(n11447), .B(n11448), .Z(n11446) );
  NAND U12517 ( .A(n11448), .B(n11447), .Z(n11443) );
  XOR U12518 ( .A(n1135), .B(n1134), .Z(\A1[501] ) );
  XOR U12519 ( .A(n11448), .B(n11449), .Z(n1134) );
  XNOR U12520 ( .A(n11447), .B(n11445), .Z(n11449) );
  AND U12521 ( .A(n11450), .B(n11451), .Z(n11445) );
  NANDN U12522 ( .A(n11452), .B(n11453), .Z(n11451) );
  NANDN U12523 ( .A(n11454), .B(n11455), .Z(n11453) );
  AND U12524 ( .A(B[500]), .B(A[3]), .Z(n11447) );
  XNOR U12525 ( .A(n11437), .B(n11456), .Z(n11448) );
  XNOR U12526 ( .A(n11435), .B(n11438), .Z(n11456) );
  NAND U12527 ( .A(A[2]), .B(B[501]), .Z(n11438) );
  NANDN U12528 ( .A(n11457), .B(n11458), .Z(n11435) );
  AND U12529 ( .A(A[0]), .B(B[502]), .Z(n11458) );
  XOR U12530 ( .A(n11440), .B(n11459), .Z(n11437) );
  NAND U12531 ( .A(A[0]), .B(B[503]), .Z(n11459) );
  NAND U12532 ( .A(B[502]), .B(A[1]), .Z(n11440) );
  NAND U12533 ( .A(n11460), .B(n11461), .Z(n1135) );
  NANDN U12534 ( .A(n11462), .B(n11463), .Z(n11461) );
  OR U12535 ( .A(n11464), .B(n11465), .Z(n11463) );
  NAND U12536 ( .A(n11465), .B(n11464), .Z(n11460) );
  XOR U12537 ( .A(n1137), .B(n1136), .Z(\A1[500] ) );
  XOR U12538 ( .A(n11465), .B(n11466), .Z(n1136) );
  XNOR U12539 ( .A(n11464), .B(n11462), .Z(n11466) );
  AND U12540 ( .A(n11467), .B(n11468), .Z(n11462) );
  NANDN U12541 ( .A(n11469), .B(n11470), .Z(n11468) );
  NANDN U12542 ( .A(n11471), .B(n11472), .Z(n11470) );
  AND U12543 ( .A(B[499]), .B(A[3]), .Z(n11464) );
  XNOR U12544 ( .A(n11454), .B(n11473), .Z(n11465) );
  XNOR U12545 ( .A(n11452), .B(n11455), .Z(n11473) );
  NAND U12546 ( .A(A[2]), .B(B[500]), .Z(n11455) );
  NANDN U12547 ( .A(n11474), .B(n11475), .Z(n11452) );
  AND U12548 ( .A(A[0]), .B(B[501]), .Z(n11475) );
  XOR U12549 ( .A(n11457), .B(n11476), .Z(n11454) );
  NAND U12550 ( .A(A[0]), .B(B[502]), .Z(n11476) );
  NAND U12551 ( .A(B[501]), .B(A[1]), .Z(n11457) );
  NAND U12552 ( .A(n11477), .B(n11478), .Z(n1137) );
  NANDN U12553 ( .A(n11479), .B(n11480), .Z(n11478) );
  OR U12554 ( .A(n11481), .B(n11482), .Z(n11480) );
  NAND U12555 ( .A(n11482), .B(n11481), .Z(n11477) );
  XOR U12556 ( .A(n919), .B(n918), .Z(\A1[4] ) );
  XOR U12557 ( .A(n9612), .B(n11483), .Z(n918) );
  XNOR U12558 ( .A(n9611), .B(n9609), .Z(n11483) );
  AND U12559 ( .A(n11484), .B(n11485), .Z(n9609) );
  NANDN U12560 ( .A(n11486), .B(n11487), .Z(n11485) );
  NANDN U12561 ( .A(n11488), .B(n11489), .Z(n11487) );
  AND U12562 ( .A(B[3]), .B(A[3]), .Z(n9611) );
  XNOR U12563 ( .A(n9601), .B(n11490), .Z(n9612) );
  XNOR U12564 ( .A(n9599), .B(n9602), .Z(n11490) );
  NAND U12565 ( .A(A[2]), .B(B[4]), .Z(n9602) );
  NANDN U12566 ( .A(n11491), .B(n11492), .Z(n9599) );
  AND U12567 ( .A(A[0]), .B(B[5]), .Z(n11492) );
  XOR U12568 ( .A(n9604), .B(n11493), .Z(n9601) );
  NAND U12569 ( .A(A[0]), .B(B[6]), .Z(n11493) );
  NAND U12570 ( .A(B[5]), .B(A[1]), .Z(n9604) );
  NAND U12571 ( .A(n11494), .B(n11495), .Z(n919) );
  NANDN U12572 ( .A(n11496), .B(n11497), .Z(n11495) );
  OR U12573 ( .A(n11498), .B(n11499), .Z(n11497) );
  NAND U12574 ( .A(n11499), .B(n11498), .Z(n11494) );
  XOR U12575 ( .A(n1119), .B(n1118), .Z(\A1[49] ) );
  XOR U12576 ( .A(n11312), .B(n11500), .Z(n1118) );
  XNOR U12577 ( .A(n11311), .B(n11309), .Z(n11500) );
  AND U12578 ( .A(n11501), .B(n11502), .Z(n11309) );
  NANDN U12579 ( .A(n11503), .B(n11504), .Z(n11502) );
  NANDN U12580 ( .A(n11505), .B(n11506), .Z(n11504) );
  AND U12581 ( .A(B[48]), .B(A[3]), .Z(n11311) );
  XNOR U12582 ( .A(n11301), .B(n11507), .Z(n11312) );
  XNOR U12583 ( .A(n11299), .B(n11302), .Z(n11507) );
  NAND U12584 ( .A(A[2]), .B(B[49]), .Z(n11302) );
  NANDN U12585 ( .A(n11508), .B(n11509), .Z(n11299) );
  AND U12586 ( .A(A[0]), .B(B[50]), .Z(n11509) );
  XOR U12587 ( .A(n11304), .B(n11510), .Z(n11301) );
  NAND U12588 ( .A(A[0]), .B(B[51]), .Z(n11510) );
  NAND U12589 ( .A(B[50]), .B(A[1]), .Z(n11304) );
  NAND U12590 ( .A(n11511), .B(n11512), .Z(n1119) );
  NANDN U12591 ( .A(n11513), .B(n11514), .Z(n11512) );
  OR U12592 ( .A(n11515), .B(n11516), .Z(n11514) );
  NAND U12593 ( .A(n11516), .B(n11515), .Z(n11511) );
  XOR U12594 ( .A(n1139), .B(n1138), .Z(\A1[499] ) );
  XOR U12595 ( .A(n11482), .B(n11517), .Z(n1138) );
  XNOR U12596 ( .A(n11481), .B(n11479), .Z(n11517) );
  AND U12597 ( .A(n11518), .B(n11519), .Z(n11479) );
  NANDN U12598 ( .A(n11520), .B(n11521), .Z(n11519) );
  NANDN U12599 ( .A(n11522), .B(n11523), .Z(n11521) );
  AND U12600 ( .A(B[498]), .B(A[3]), .Z(n11481) );
  XNOR U12601 ( .A(n11471), .B(n11524), .Z(n11482) );
  XNOR U12602 ( .A(n11469), .B(n11472), .Z(n11524) );
  NAND U12603 ( .A(A[2]), .B(B[499]), .Z(n11472) );
  NANDN U12604 ( .A(n11525), .B(n11526), .Z(n11469) );
  AND U12605 ( .A(A[0]), .B(B[500]), .Z(n11526) );
  XOR U12606 ( .A(n11474), .B(n11527), .Z(n11471) );
  NAND U12607 ( .A(A[0]), .B(B[501]), .Z(n11527) );
  NAND U12608 ( .A(B[500]), .B(A[1]), .Z(n11474) );
  NAND U12609 ( .A(n11528), .B(n11529), .Z(n1139) );
  NANDN U12610 ( .A(n11530), .B(n11531), .Z(n11529) );
  OR U12611 ( .A(n11532), .B(n11533), .Z(n11531) );
  NAND U12612 ( .A(n11533), .B(n11532), .Z(n11528) );
  XOR U12613 ( .A(n1145), .B(n1144), .Z(\A1[498] ) );
  XOR U12614 ( .A(n11533), .B(n11534), .Z(n1144) );
  XNOR U12615 ( .A(n11532), .B(n11530), .Z(n11534) );
  AND U12616 ( .A(n11535), .B(n11536), .Z(n11530) );
  NANDN U12617 ( .A(n11537), .B(n11538), .Z(n11536) );
  NANDN U12618 ( .A(n11539), .B(n11540), .Z(n11538) );
  AND U12619 ( .A(B[497]), .B(A[3]), .Z(n11532) );
  XNOR U12620 ( .A(n11522), .B(n11541), .Z(n11533) );
  XNOR U12621 ( .A(n11520), .B(n11523), .Z(n11541) );
  NAND U12622 ( .A(A[2]), .B(B[498]), .Z(n11523) );
  NANDN U12623 ( .A(n11542), .B(n11543), .Z(n11520) );
  AND U12624 ( .A(A[0]), .B(B[499]), .Z(n11543) );
  XOR U12625 ( .A(n11525), .B(n11544), .Z(n11522) );
  NAND U12626 ( .A(A[0]), .B(B[500]), .Z(n11544) );
  NAND U12627 ( .A(B[499]), .B(A[1]), .Z(n11525) );
  NAND U12628 ( .A(n11545), .B(n11546), .Z(n1145) );
  NANDN U12629 ( .A(n11547), .B(n11548), .Z(n11546) );
  OR U12630 ( .A(n11549), .B(n11550), .Z(n11548) );
  NAND U12631 ( .A(n11550), .B(n11549), .Z(n11545) );
  XOR U12632 ( .A(n1147), .B(n1146), .Z(\A1[497] ) );
  XOR U12633 ( .A(n11550), .B(n11551), .Z(n1146) );
  XNOR U12634 ( .A(n11549), .B(n11547), .Z(n11551) );
  AND U12635 ( .A(n11552), .B(n11553), .Z(n11547) );
  NANDN U12636 ( .A(n11554), .B(n11555), .Z(n11553) );
  NANDN U12637 ( .A(n11556), .B(n11557), .Z(n11555) );
  AND U12638 ( .A(B[496]), .B(A[3]), .Z(n11549) );
  XNOR U12639 ( .A(n11539), .B(n11558), .Z(n11550) );
  XNOR U12640 ( .A(n11537), .B(n11540), .Z(n11558) );
  NAND U12641 ( .A(A[2]), .B(B[497]), .Z(n11540) );
  NANDN U12642 ( .A(n11559), .B(n11560), .Z(n11537) );
  AND U12643 ( .A(A[0]), .B(B[498]), .Z(n11560) );
  XOR U12644 ( .A(n11542), .B(n11561), .Z(n11539) );
  NAND U12645 ( .A(A[0]), .B(B[499]), .Z(n11561) );
  NAND U12646 ( .A(B[498]), .B(A[1]), .Z(n11542) );
  NAND U12647 ( .A(n11562), .B(n11563), .Z(n1147) );
  NANDN U12648 ( .A(n11564), .B(n11565), .Z(n11563) );
  OR U12649 ( .A(n11566), .B(n11567), .Z(n11565) );
  NAND U12650 ( .A(n11567), .B(n11566), .Z(n11562) );
  XOR U12651 ( .A(n1149), .B(n1148), .Z(\A1[496] ) );
  XOR U12652 ( .A(n11567), .B(n11568), .Z(n1148) );
  XNOR U12653 ( .A(n11566), .B(n11564), .Z(n11568) );
  AND U12654 ( .A(n11569), .B(n11570), .Z(n11564) );
  NANDN U12655 ( .A(n11571), .B(n11572), .Z(n11570) );
  NANDN U12656 ( .A(n11573), .B(n11574), .Z(n11572) );
  AND U12657 ( .A(B[495]), .B(A[3]), .Z(n11566) );
  XNOR U12658 ( .A(n11556), .B(n11575), .Z(n11567) );
  XNOR U12659 ( .A(n11554), .B(n11557), .Z(n11575) );
  NAND U12660 ( .A(A[2]), .B(B[496]), .Z(n11557) );
  NANDN U12661 ( .A(n11576), .B(n11577), .Z(n11554) );
  AND U12662 ( .A(A[0]), .B(B[497]), .Z(n11577) );
  XOR U12663 ( .A(n11559), .B(n11578), .Z(n11556) );
  NAND U12664 ( .A(A[0]), .B(B[498]), .Z(n11578) );
  NAND U12665 ( .A(B[497]), .B(A[1]), .Z(n11559) );
  NAND U12666 ( .A(n11579), .B(n11580), .Z(n1149) );
  NANDN U12667 ( .A(n11581), .B(n11582), .Z(n11580) );
  OR U12668 ( .A(n11583), .B(n11584), .Z(n11582) );
  NAND U12669 ( .A(n11584), .B(n11583), .Z(n11579) );
  XOR U12670 ( .A(n1151), .B(n1150), .Z(\A1[495] ) );
  XOR U12671 ( .A(n11584), .B(n11585), .Z(n1150) );
  XNOR U12672 ( .A(n11583), .B(n11581), .Z(n11585) );
  AND U12673 ( .A(n11586), .B(n11587), .Z(n11581) );
  NANDN U12674 ( .A(n11588), .B(n11589), .Z(n11587) );
  NANDN U12675 ( .A(n11590), .B(n11591), .Z(n11589) );
  AND U12676 ( .A(B[494]), .B(A[3]), .Z(n11583) );
  XNOR U12677 ( .A(n11573), .B(n11592), .Z(n11584) );
  XNOR U12678 ( .A(n11571), .B(n11574), .Z(n11592) );
  NAND U12679 ( .A(A[2]), .B(B[495]), .Z(n11574) );
  NANDN U12680 ( .A(n11593), .B(n11594), .Z(n11571) );
  AND U12681 ( .A(A[0]), .B(B[496]), .Z(n11594) );
  XOR U12682 ( .A(n11576), .B(n11595), .Z(n11573) );
  NAND U12683 ( .A(A[0]), .B(B[497]), .Z(n11595) );
  NAND U12684 ( .A(B[496]), .B(A[1]), .Z(n11576) );
  NAND U12685 ( .A(n11596), .B(n11597), .Z(n1151) );
  NANDN U12686 ( .A(n11598), .B(n11599), .Z(n11597) );
  OR U12687 ( .A(n11600), .B(n11601), .Z(n11599) );
  NAND U12688 ( .A(n11601), .B(n11600), .Z(n11596) );
  XOR U12689 ( .A(n1153), .B(n1152), .Z(\A1[494] ) );
  XOR U12690 ( .A(n11601), .B(n11602), .Z(n1152) );
  XNOR U12691 ( .A(n11600), .B(n11598), .Z(n11602) );
  AND U12692 ( .A(n11603), .B(n11604), .Z(n11598) );
  NANDN U12693 ( .A(n11605), .B(n11606), .Z(n11604) );
  NANDN U12694 ( .A(n11607), .B(n11608), .Z(n11606) );
  AND U12695 ( .A(B[493]), .B(A[3]), .Z(n11600) );
  XNOR U12696 ( .A(n11590), .B(n11609), .Z(n11601) );
  XNOR U12697 ( .A(n11588), .B(n11591), .Z(n11609) );
  NAND U12698 ( .A(A[2]), .B(B[494]), .Z(n11591) );
  NANDN U12699 ( .A(n11610), .B(n11611), .Z(n11588) );
  AND U12700 ( .A(A[0]), .B(B[495]), .Z(n11611) );
  XOR U12701 ( .A(n11593), .B(n11612), .Z(n11590) );
  NAND U12702 ( .A(A[0]), .B(B[496]), .Z(n11612) );
  NAND U12703 ( .A(B[495]), .B(A[1]), .Z(n11593) );
  NAND U12704 ( .A(n11613), .B(n11614), .Z(n1153) );
  NANDN U12705 ( .A(n11615), .B(n11616), .Z(n11614) );
  OR U12706 ( .A(n11617), .B(n11618), .Z(n11616) );
  NAND U12707 ( .A(n11618), .B(n11617), .Z(n11613) );
  XOR U12708 ( .A(n1155), .B(n1154), .Z(\A1[493] ) );
  XOR U12709 ( .A(n11618), .B(n11619), .Z(n1154) );
  XNOR U12710 ( .A(n11617), .B(n11615), .Z(n11619) );
  AND U12711 ( .A(n11620), .B(n11621), .Z(n11615) );
  NANDN U12712 ( .A(n11622), .B(n11623), .Z(n11621) );
  NANDN U12713 ( .A(n11624), .B(n11625), .Z(n11623) );
  AND U12714 ( .A(B[492]), .B(A[3]), .Z(n11617) );
  XNOR U12715 ( .A(n11607), .B(n11626), .Z(n11618) );
  XNOR U12716 ( .A(n11605), .B(n11608), .Z(n11626) );
  NAND U12717 ( .A(A[2]), .B(B[493]), .Z(n11608) );
  NANDN U12718 ( .A(n11627), .B(n11628), .Z(n11605) );
  AND U12719 ( .A(A[0]), .B(B[494]), .Z(n11628) );
  XOR U12720 ( .A(n11610), .B(n11629), .Z(n11607) );
  NAND U12721 ( .A(A[0]), .B(B[495]), .Z(n11629) );
  NAND U12722 ( .A(B[494]), .B(A[1]), .Z(n11610) );
  NAND U12723 ( .A(n11630), .B(n11631), .Z(n1155) );
  NANDN U12724 ( .A(n11632), .B(n11633), .Z(n11631) );
  OR U12725 ( .A(n11634), .B(n11635), .Z(n11633) );
  NAND U12726 ( .A(n11635), .B(n11634), .Z(n11630) );
  XOR U12727 ( .A(n1157), .B(n1156), .Z(\A1[492] ) );
  XOR U12728 ( .A(n11635), .B(n11636), .Z(n1156) );
  XNOR U12729 ( .A(n11634), .B(n11632), .Z(n11636) );
  AND U12730 ( .A(n11637), .B(n11638), .Z(n11632) );
  NANDN U12731 ( .A(n11639), .B(n11640), .Z(n11638) );
  NANDN U12732 ( .A(n11641), .B(n11642), .Z(n11640) );
  AND U12733 ( .A(B[491]), .B(A[3]), .Z(n11634) );
  XNOR U12734 ( .A(n11624), .B(n11643), .Z(n11635) );
  XNOR U12735 ( .A(n11622), .B(n11625), .Z(n11643) );
  NAND U12736 ( .A(A[2]), .B(B[492]), .Z(n11625) );
  NANDN U12737 ( .A(n11644), .B(n11645), .Z(n11622) );
  AND U12738 ( .A(A[0]), .B(B[493]), .Z(n11645) );
  XOR U12739 ( .A(n11627), .B(n11646), .Z(n11624) );
  NAND U12740 ( .A(A[0]), .B(B[494]), .Z(n11646) );
  NAND U12741 ( .A(B[493]), .B(A[1]), .Z(n11627) );
  NAND U12742 ( .A(n11647), .B(n11648), .Z(n1157) );
  NANDN U12743 ( .A(n11649), .B(n11650), .Z(n11648) );
  OR U12744 ( .A(n11651), .B(n11652), .Z(n11650) );
  NAND U12745 ( .A(n11652), .B(n11651), .Z(n11647) );
  XOR U12746 ( .A(n1159), .B(n1158), .Z(\A1[491] ) );
  XOR U12747 ( .A(n11652), .B(n11653), .Z(n1158) );
  XNOR U12748 ( .A(n11651), .B(n11649), .Z(n11653) );
  AND U12749 ( .A(n11654), .B(n11655), .Z(n11649) );
  NANDN U12750 ( .A(n11656), .B(n11657), .Z(n11655) );
  NANDN U12751 ( .A(n11658), .B(n11659), .Z(n11657) );
  AND U12752 ( .A(B[490]), .B(A[3]), .Z(n11651) );
  XNOR U12753 ( .A(n11641), .B(n11660), .Z(n11652) );
  XNOR U12754 ( .A(n11639), .B(n11642), .Z(n11660) );
  NAND U12755 ( .A(A[2]), .B(B[491]), .Z(n11642) );
  NANDN U12756 ( .A(n11661), .B(n11662), .Z(n11639) );
  AND U12757 ( .A(A[0]), .B(B[492]), .Z(n11662) );
  XOR U12758 ( .A(n11644), .B(n11663), .Z(n11641) );
  NAND U12759 ( .A(A[0]), .B(B[493]), .Z(n11663) );
  NAND U12760 ( .A(B[492]), .B(A[1]), .Z(n11644) );
  NAND U12761 ( .A(n11664), .B(n11665), .Z(n1159) );
  NANDN U12762 ( .A(n11666), .B(n11667), .Z(n11665) );
  OR U12763 ( .A(n11668), .B(n11669), .Z(n11667) );
  NAND U12764 ( .A(n11669), .B(n11668), .Z(n11664) );
  XOR U12765 ( .A(n1161), .B(n1160), .Z(\A1[490] ) );
  XOR U12766 ( .A(n11669), .B(n11670), .Z(n1160) );
  XNOR U12767 ( .A(n11668), .B(n11666), .Z(n11670) );
  AND U12768 ( .A(n11671), .B(n11672), .Z(n11666) );
  NANDN U12769 ( .A(n11673), .B(n11674), .Z(n11672) );
  NANDN U12770 ( .A(n11675), .B(n11676), .Z(n11674) );
  AND U12771 ( .A(B[489]), .B(A[3]), .Z(n11668) );
  XNOR U12772 ( .A(n11658), .B(n11677), .Z(n11669) );
  XNOR U12773 ( .A(n11656), .B(n11659), .Z(n11677) );
  NAND U12774 ( .A(A[2]), .B(B[490]), .Z(n11659) );
  NANDN U12775 ( .A(n11678), .B(n11679), .Z(n11656) );
  AND U12776 ( .A(A[0]), .B(B[491]), .Z(n11679) );
  XOR U12777 ( .A(n11661), .B(n11680), .Z(n11658) );
  NAND U12778 ( .A(A[0]), .B(B[492]), .Z(n11680) );
  NAND U12779 ( .A(B[491]), .B(A[1]), .Z(n11661) );
  NAND U12780 ( .A(n11681), .B(n11682), .Z(n1161) );
  NANDN U12781 ( .A(n11683), .B(n11684), .Z(n11682) );
  OR U12782 ( .A(n11685), .B(n11686), .Z(n11684) );
  NAND U12783 ( .A(n11686), .B(n11685), .Z(n11681) );
  XOR U12784 ( .A(n1143), .B(n1142), .Z(\A1[48] ) );
  XOR U12785 ( .A(n11516), .B(n11687), .Z(n1142) );
  XNOR U12786 ( .A(n11515), .B(n11513), .Z(n11687) );
  AND U12787 ( .A(n11688), .B(n11689), .Z(n11513) );
  NANDN U12788 ( .A(n11690), .B(n11691), .Z(n11689) );
  NANDN U12789 ( .A(n11692), .B(n11693), .Z(n11691) );
  AND U12790 ( .A(B[47]), .B(A[3]), .Z(n11515) );
  XNOR U12791 ( .A(n11505), .B(n11694), .Z(n11516) );
  XNOR U12792 ( .A(n11503), .B(n11506), .Z(n11694) );
  NAND U12793 ( .A(A[2]), .B(B[48]), .Z(n11506) );
  NANDN U12794 ( .A(n11695), .B(n11696), .Z(n11503) );
  AND U12795 ( .A(A[0]), .B(B[49]), .Z(n11696) );
  XOR U12796 ( .A(n11508), .B(n11697), .Z(n11505) );
  NAND U12797 ( .A(A[0]), .B(B[50]), .Z(n11697) );
  NAND U12798 ( .A(B[49]), .B(A[1]), .Z(n11508) );
  NAND U12799 ( .A(n11698), .B(n11699), .Z(n1143) );
  NANDN U12800 ( .A(n11700), .B(n11701), .Z(n11699) );
  OR U12801 ( .A(n11702), .B(n11703), .Z(n11701) );
  NAND U12802 ( .A(n11703), .B(n11702), .Z(n11698) );
  XOR U12803 ( .A(n1163), .B(n1162), .Z(\A1[489] ) );
  XOR U12804 ( .A(n11686), .B(n11704), .Z(n1162) );
  XNOR U12805 ( .A(n11685), .B(n11683), .Z(n11704) );
  AND U12806 ( .A(n11705), .B(n11706), .Z(n11683) );
  NANDN U12807 ( .A(n11707), .B(n11708), .Z(n11706) );
  NANDN U12808 ( .A(n11709), .B(n11710), .Z(n11708) );
  AND U12809 ( .A(B[488]), .B(A[3]), .Z(n11685) );
  XNOR U12810 ( .A(n11675), .B(n11711), .Z(n11686) );
  XNOR U12811 ( .A(n11673), .B(n11676), .Z(n11711) );
  NAND U12812 ( .A(A[2]), .B(B[489]), .Z(n11676) );
  NANDN U12813 ( .A(n11712), .B(n11713), .Z(n11673) );
  AND U12814 ( .A(A[0]), .B(B[490]), .Z(n11713) );
  XOR U12815 ( .A(n11678), .B(n11714), .Z(n11675) );
  NAND U12816 ( .A(A[0]), .B(B[491]), .Z(n11714) );
  NAND U12817 ( .A(B[490]), .B(A[1]), .Z(n11678) );
  NAND U12818 ( .A(n11715), .B(n11716), .Z(n1163) );
  NANDN U12819 ( .A(n11717), .B(n11718), .Z(n11716) );
  OR U12820 ( .A(n11719), .B(n11720), .Z(n11718) );
  NAND U12821 ( .A(n11720), .B(n11719), .Z(n11715) );
  XOR U12822 ( .A(n1167), .B(n1166), .Z(\A1[488] ) );
  XOR U12823 ( .A(n11720), .B(n11721), .Z(n1166) );
  XNOR U12824 ( .A(n11719), .B(n11717), .Z(n11721) );
  AND U12825 ( .A(n11722), .B(n11723), .Z(n11717) );
  NANDN U12826 ( .A(n11724), .B(n11725), .Z(n11723) );
  NANDN U12827 ( .A(n11726), .B(n11727), .Z(n11725) );
  AND U12828 ( .A(B[487]), .B(A[3]), .Z(n11719) );
  XNOR U12829 ( .A(n11709), .B(n11728), .Z(n11720) );
  XNOR U12830 ( .A(n11707), .B(n11710), .Z(n11728) );
  NAND U12831 ( .A(A[2]), .B(B[488]), .Z(n11710) );
  NANDN U12832 ( .A(n11729), .B(n11730), .Z(n11707) );
  AND U12833 ( .A(A[0]), .B(B[489]), .Z(n11730) );
  XOR U12834 ( .A(n11712), .B(n11731), .Z(n11709) );
  NAND U12835 ( .A(A[0]), .B(B[490]), .Z(n11731) );
  NAND U12836 ( .A(B[489]), .B(A[1]), .Z(n11712) );
  NAND U12837 ( .A(n11732), .B(n11733), .Z(n1167) );
  NANDN U12838 ( .A(n11734), .B(n11735), .Z(n11733) );
  OR U12839 ( .A(n11736), .B(n11737), .Z(n11735) );
  NAND U12840 ( .A(n11737), .B(n11736), .Z(n11732) );
  XOR U12841 ( .A(n1169), .B(n1168), .Z(\A1[487] ) );
  XOR U12842 ( .A(n11737), .B(n11738), .Z(n1168) );
  XNOR U12843 ( .A(n11736), .B(n11734), .Z(n11738) );
  AND U12844 ( .A(n11739), .B(n11740), .Z(n11734) );
  NANDN U12845 ( .A(n11741), .B(n11742), .Z(n11740) );
  NANDN U12846 ( .A(n11743), .B(n11744), .Z(n11742) );
  AND U12847 ( .A(B[486]), .B(A[3]), .Z(n11736) );
  XNOR U12848 ( .A(n11726), .B(n11745), .Z(n11737) );
  XNOR U12849 ( .A(n11724), .B(n11727), .Z(n11745) );
  NAND U12850 ( .A(A[2]), .B(B[487]), .Z(n11727) );
  NANDN U12851 ( .A(n11746), .B(n11747), .Z(n11724) );
  AND U12852 ( .A(A[0]), .B(B[488]), .Z(n11747) );
  XOR U12853 ( .A(n11729), .B(n11748), .Z(n11726) );
  NAND U12854 ( .A(A[0]), .B(B[489]), .Z(n11748) );
  NAND U12855 ( .A(B[488]), .B(A[1]), .Z(n11729) );
  NAND U12856 ( .A(n11749), .B(n11750), .Z(n1169) );
  NANDN U12857 ( .A(n11751), .B(n11752), .Z(n11750) );
  OR U12858 ( .A(n11753), .B(n11754), .Z(n11752) );
  NAND U12859 ( .A(n11754), .B(n11753), .Z(n11749) );
  XOR U12860 ( .A(n1171), .B(n1170), .Z(\A1[486] ) );
  XOR U12861 ( .A(n11754), .B(n11755), .Z(n1170) );
  XNOR U12862 ( .A(n11753), .B(n11751), .Z(n11755) );
  AND U12863 ( .A(n11756), .B(n11757), .Z(n11751) );
  NANDN U12864 ( .A(n11758), .B(n11759), .Z(n11757) );
  NANDN U12865 ( .A(n11760), .B(n11761), .Z(n11759) );
  AND U12866 ( .A(B[485]), .B(A[3]), .Z(n11753) );
  XNOR U12867 ( .A(n11743), .B(n11762), .Z(n11754) );
  XNOR U12868 ( .A(n11741), .B(n11744), .Z(n11762) );
  NAND U12869 ( .A(A[2]), .B(B[486]), .Z(n11744) );
  NANDN U12870 ( .A(n11763), .B(n11764), .Z(n11741) );
  AND U12871 ( .A(A[0]), .B(B[487]), .Z(n11764) );
  XOR U12872 ( .A(n11746), .B(n11765), .Z(n11743) );
  NAND U12873 ( .A(A[0]), .B(B[488]), .Z(n11765) );
  NAND U12874 ( .A(B[487]), .B(A[1]), .Z(n11746) );
  NAND U12875 ( .A(n11766), .B(n11767), .Z(n1171) );
  NANDN U12876 ( .A(n11768), .B(n11769), .Z(n11767) );
  OR U12877 ( .A(n11770), .B(n11771), .Z(n11769) );
  NAND U12878 ( .A(n11771), .B(n11770), .Z(n11766) );
  XOR U12879 ( .A(n1173), .B(n1172), .Z(\A1[485] ) );
  XOR U12880 ( .A(n11771), .B(n11772), .Z(n1172) );
  XNOR U12881 ( .A(n11770), .B(n11768), .Z(n11772) );
  AND U12882 ( .A(n11773), .B(n11774), .Z(n11768) );
  NANDN U12883 ( .A(n11775), .B(n11776), .Z(n11774) );
  NANDN U12884 ( .A(n11777), .B(n11778), .Z(n11776) );
  AND U12885 ( .A(B[484]), .B(A[3]), .Z(n11770) );
  XNOR U12886 ( .A(n11760), .B(n11779), .Z(n11771) );
  XNOR U12887 ( .A(n11758), .B(n11761), .Z(n11779) );
  NAND U12888 ( .A(A[2]), .B(B[485]), .Z(n11761) );
  NANDN U12889 ( .A(n11780), .B(n11781), .Z(n11758) );
  AND U12890 ( .A(A[0]), .B(B[486]), .Z(n11781) );
  XOR U12891 ( .A(n11763), .B(n11782), .Z(n11760) );
  NAND U12892 ( .A(A[0]), .B(B[487]), .Z(n11782) );
  NAND U12893 ( .A(B[486]), .B(A[1]), .Z(n11763) );
  NAND U12894 ( .A(n11783), .B(n11784), .Z(n1173) );
  NANDN U12895 ( .A(n11785), .B(n11786), .Z(n11784) );
  OR U12896 ( .A(n11787), .B(n11788), .Z(n11786) );
  NAND U12897 ( .A(n11788), .B(n11787), .Z(n11783) );
  XOR U12898 ( .A(n1175), .B(n1174), .Z(\A1[484] ) );
  XOR U12899 ( .A(n11788), .B(n11789), .Z(n1174) );
  XNOR U12900 ( .A(n11787), .B(n11785), .Z(n11789) );
  AND U12901 ( .A(n11790), .B(n11791), .Z(n11785) );
  NANDN U12902 ( .A(n11792), .B(n11793), .Z(n11791) );
  NANDN U12903 ( .A(n11794), .B(n11795), .Z(n11793) );
  AND U12904 ( .A(B[483]), .B(A[3]), .Z(n11787) );
  XNOR U12905 ( .A(n11777), .B(n11796), .Z(n11788) );
  XNOR U12906 ( .A(n11775), .B(n11778), .Z(n11796) );
  NAND U12907 ( .A(A[2]), .B(B[484]), .Z(n11778) );
  NANDN U12908 ( .A(n11797), .B(n11798), .Z(n11775) );
  AND U12909 ( .A(A[0]), .B(B[485]), .Z(n11798) );
  XOR U12910 ( .A(n11780), .B(n11799), .Z(n11777) );
  NAND U12911 ( .A(A[0]), .B(B[486]), .Z(n11799) );
  NAND U12912 ( .A(B[485]), .B(A[1]), .Z(n11780) );
  NAND U12913 ( .A(n11800), .B(n11801), .Z(n1175) );
  NANDN U12914 ( .A(n11802), .B(n11803), .Z(n11801) );
  OR U12915 ( .A(n11804), .B(n11805), .Z(n11803) );
  NAND U12916 ( .A(n11805), .B(n11804), .Z(n11800) );
  XOR U12917 ( .A(n1177), .B(n1176), .Z(\A1[483] ) );
  XOR U12918 ( .A(n11805), .B(n11806), .Z(n1176) );
  XNOR U12919 ( .A(n11804), .B(n11802), .Z(n11806) );
  AND U12920 ( .A(n11807), .B(n11808), .Z(n11802) );
  NANDN U12921 ( .A(n11809), .B(n11810), .Z(n11808) );
  NANDN U12922 ( .A(n11811), .B(n11812), .Z(n11810) );
  AND U12923 ( .A(B[482]), .B(A[3]), .Z(n11804) );
  XNOR U12924 ( .A(n11794), .B(n11813), .Z(n11805) );
  XNOR U12925 ( .A(n11792), .B(n11795), .Z(n11813) );
  NAND U12926 ( .A(A[2]), .B(B[483]), .Z(n11795) );
  NANDN U12927 ( .A(n11814), .B(n11815), .Z(n11792) );
  AND U12928 ( .A(A[0]), .B(B[484]), .Z(n11815) );
  XOR U12929 ( .A(n11797), .B(n11816), .Z(n11794) );
  NAND U12930 ( .A(A[0]), .B(B[485]), .Z(n11816) );
  NAND U12931 ( .A(B[484]), .B(A[1]), .Z(n11797) );
  NAND U12932 ( .A(n11817), .B(n11818), .Z(n1177) );
  NANDN U12933 ( .A(n11819), .B(n11820), .Z(n11818) );
  OR U12934 ( .A(n11821), .B(n11822), .Z(n11820) );
  NAND U12935 ( .A(n11822), .B(n11821), .Z(n11817) );
  XOR U12936 ( .A(n1179), .B(n1178), .Z(\A1[482] ) );
  XOR U12937 ( .A(n11822), .B(n11823), .Z(n1178) );
  XNOR U12938 ( .A(n11821), .B(n11819), .Z(n11823) );
  AND U12939 ( .A(n11824), .B(n11825), .Z(n11819) );
  NANDN U12940 ( .A(n11826), .B(n11827), .Z(n11825) );
  NANDN U12941 ( .A(n11828), .B(n11829), .Z(n11827) );
  AND U12942 ( .A(B[481]), .B(A[3]), .Z(n11821) );
  XNOR U12943 ( .A(n11811), .B(n11830), .Z(n11822) );
  XNOR U12944 ( .A(n11809), .B(n11812), .Z(n11830) );
  NAND U12945 ( .A(A[2]), .B(B[482]), .Z(n11812) );
  NANDN U12946 ( .A(n11831), .B(n11832), .Z(n11809) );
  AND U12947 ( .A(A[0]), .B(B[483]), .Z(n11832) );
  XOR U12948 ( .A(n11814), .B(n11833), .Z(n11811) );
  NAND U12949 ( .A(A[0]), .B(B[484]), .Z(n11833) );
  NAND U12950 ( .A(B[483]), .B(A[1]), .Z(n11814) );
  NAND U12951 ( .A(n11834), .B(n11835), .Z(n1179) );
  NANDN U12952 ( .A(n11836), .B(n11837), .Z(n11835) );
  OR U12953 ( .A(n11838), .B(n11839), .Z(n11837) );
  NAND U12954 ( .A(n11839), .B(n11838), .Z(n11834) );
  XOR U12955 ( .A(n1181), .B(n1180), .Z(\A1[481] ) );
  XOR U12956 ( .A(n11839), .B(n11840), .Z(n1180) );
  XNOR U12957 ( .A(n11838), .B(n11836), .Z(n11840) );
  AND U12958 ( .A(n11841), .B(n11842), .Z(n11836) );
  NANDN U12959 ( .A(n11843), .B(n11844), .Z(n11842) );
  NANDN U12960 ( .A(n11845), .B(n11846), .Z(n11844) );
  AND U12961 ( .A(B[480]), .B(A[3]), .Z(n11838) );
  XNOR U12962 ( .A(n11828), .B(n11847), .Z(n11839) );
  XNOR U12963 ( .A(n11826), .B(n11829), .Z(n11847) );
  NAND U12964 ( .A(A[2]), .B(B[481]), .Z(n11829) );
  NANDN U12965 ( .A(n11848), .B(n11849), .Z(n11826) );
  AND U12966 ( .A(A[0]), .B(B[482]), .Z(n11849) );
  XOR U12967 ( .A(n11831), .B(n11850), .Z(n11828) );
  NAND U12968 ( .A(A[0]), .B(B[483]), .Z(n11850) );
  NAND U12969 ( .A(B[482]), .B(A[1]), .Z(n11831) );
  NAND U12970 ( .A(n11851), .B(n11852), .Z(n1181) );
  NANDN U12971 ( .A(n11853), .B(n11854), .Z(n11852) );
  OR U12972 ( .A(n11855), .B(n11856), .Z(n11854) );
  NAND U12973 ( .A(n11856), .B(n11855), .Z(n11851) );
  XOR U12974 ( .A(n1183), .B(n1182), .Z(\A1[480] ) );
  XOR U12975 ( .A(n11856), .B(n11857), .Z(n1182) );
  XNOR U12976 ( .A(n11855), .B(n11853), .Z(n11857) );
  AND U12977 ( .A(n11858), .B(n11859), .Z(n11853) );
  NANDN U12978 ( .A(n11860), .B(n11861), .Z(n11859) );
  NANDN U12979 ( .A(n11862), .B(n11863), .Z(n11861) );
  AND U12980 ( .A(B[479]), .B(A[3]), .Z(n11855) );
  XNOR U12981 ( .A(n11845), .B(n11864), .Z(n11856) );
  XNOR U12982 ( .A(n11843), .B(n11846), .Z(n11864) );
  NAND U12983 ( .A(A[2]), .B(B[480]), .Z(n11846) );
  NANDN U12984 ( .A(n11865), .B(n11866), .Z(n11843) );
  AND U12985 ( .A(A[0]), .B(B[481]), .Z(n11866) );
  XOR U12986 ( .A(n11848), .B(n11867), .Z(n11845) );
  NAND U12987 ( .A(A[0]), .B(B[482]), .Z(n11867) );
  NAND U12988 ( .A(B[481]), .B(A[1]), .Z(n11848) );
  NAND U12989 ( .A(n11868), .B(n11869), .Z(n1183) );
  NANDN U12990 ( .A(n11870), .B(n11871), .Z(n11869) );
  OR U12991 ( .A(n11872), .B(n11873), .Z(n11871) );
  NAND U12992 ( .A(n11873), .B(n11872), .Z(n11868) );
  XOR U12993 ( .A(n1165), .B(n1164), .Z(\A1[47] ) );
  XOR U12994 ( .A(n11703), .B(n11874), .Z(n1164) );
  XNOR U12995 ( .A(n11702), .B(n11700), .Z(n11874) );
  AND U12996 ( .A(n11875), .B(n11876), .Z(n11700) );
  NANDN U12997 ( .A(n11877), .B(n11878), .Z(n11876) );
  NANDN U12998 ( .A(n11879), .B(n11880), .Z(n11878) );
  AND U12999 ( .A(B[46]), .B(A[3]), .Z(n11702) );
  XNOR U13000 ( .A(n11692), .B(n11881), .Z(n11703) );
  XNOR U13001 ( .A(n11690), .B(n11693), .Z(n11881) );
  NAND U13002 ( .A(A[2]), .B(B[47]), .Z(n11693) );
  NANDN U13003 ( .A(n11882), .B(n11883), .Z(n11690) );
  AND U13004 ( .A(A[0]), .B(B[48]), .Z(n11883) );
  XOR U13005 ( .A(n11695), .B(n11884), .Z(n11692) );
  NAND U13006 ( .A(A[0]), .B(B[49]), .Z(n11884) );
  NAND U13007 ( .A(B[48]), .B(A[1]), .Z(n11695) );
  NAND U13008 ( .A(n11885), .B(n11886), .Z(n1165) );
  NANDN U13009 ( .A(n11887), .B(n11888), .Z(n11886) );
  OR U13010 ( .A(n11889), .B(n11890), .Z(n11888) );
  NAND U13011 ( .A(n11890), .B(n11889), .Z(n11885) );
  XOR U13012 ( .A(n1185), .B(n1184), .Z(\A1[479] ) );
  XOR U13013 ( .A(n11873), .B(n11891), .Z(n1184) );
  XNOR U13014 ( .A(n11872), .B(n11870), .Z(n11891) );
  AND U13015 ( .A(n11892), .B(n11893), .Z(n11870) );
  NANDN U13016 ( .A(n11894), .B(n11895), .Z(n11893) );
  NANDN U13017 ( .A(n11896), .B(n11897), .Z(n11895) );
  AND U13018 ( .A(B[478]), .B(A[3]), .Z(n11872) );
  XNOR U13019 ( .A(n11862), .B(n11898), .Z(n11873) );
  XNOR U13020 ( .A(n11860), .B(n11863), .Z(n11898) );
  NAND U13021 ( .A(A[2]), .B(B[479]), .Z(n11863) );
  NANDN U13022 ( .A(n11899), .B(n11900), .Z(n11860) );
  AND U13023 ( .A(A[0]), .B(B[480]), .Z(n11900) );
  XOR U13024 ( .A(n11865), .B(n11901), .Z(n11862) );
  NAND U13025 ( .A(A[0]), .B(B[481]), .Z(n11901) );
  NAND U13026 ( .A(B[480]), .B(A[1]), .Z(n11865) );
  NAND U13027 ( .A(n11902), .B(n11903), .Z(n1185) );
  NANDN U13028 ( .A(n11904), .B(n11905), .Z(n11903) );
  OR U13029 ( .A(n11906), .B(n11907), .Z(n11905) );
  NAND U13030 ( .A(n11907), .B(n11906), .Z(n11902) );
  XOR U13031 ( .A(n1189), .B(n1188), .Z(\A1[478] ) );
  XOR U13032 ( .A(n11907), .B(n11908), .Z(n1188) );
  XNOR U13033 ( .A(n11906), .B(n11904), .Z(n11908) );
  AND U13034 ( .A(n11909), .B(n11910), .Z(n11904) );
  NANDN U13035 ( .A(n11911), .B(n11912), .Z(n11910) );
  NANDN U13036 ( .A(n11913), .B(n11914), .Z(n11912) );
  AND U13037 ( .A(B[477]), .B(A[3]), .Z(n11906) );
  XNOR U13038 ( .A(n11896), .B(n11915), .Z(n11907) );
  XNOR U13039 ( .A(n11894), .B(n11897), .Z(n11915) );
  NAND U13040 ( .A(A[2]), .B(B[478]), .Z(n11897) );
  NANDN U13041 ( .A(n11916), .B(n11917), .Z(n11894) );
  AND U13042 ( .A(A[0]), .B(B[479]), .Z(n11917) );
  XOR U13043 ( .A(n11899), .B(n11918), .Z(n11896) );
  NAND U13044 ( .A(A[0]), .B(B[480]), .Z(n11918) );
  NAND U13045 ( .A(B[479]), .B(A[1]), .Z(n11899) );
  NAND U13046 ( .A(n11919), .B(n11920), .Z(n1189) );
  NANDN U13047 ( .A(n11921), .B(n11922), .Z(n11920) );
  OR U13048 ( .A(n11923), .B(n11924), .Z(n11922) );
  NAND U13049 ( .A(n11924), .B(n11923), .Z(n11919) );
  XOR U13050 ( .A(n1191), .B(n1190), .Z(\A1[477] ) );
  XOR U13051 ( .A(n11924), .B(n11925), .Z(n1190) );
  XNOR U13052 ( .A(n11923), .B(n11921), .Z(n11925) );
  AND U13053 ( .A(n11926), .B(n11927), .Z(n11921) );
  NANDN U13054 ( .A(n11928), .B(n11929), .Z(n11927) );
  NANDN U13055 ( .A(n11930), .B(n11931), .Z(n11929) );
  AND U13056 ( .A(B[476]), .B(A[3]), .Z(n11923) );
  XNOR U13057 ( .A(n11913), .B(n11932), .Z(n11924) );
  XNOR U13058 ( .A(n11911), .B(n11914), .Z(n11932) );
  NAND U13059 ( .A(A[2]), .B(B[477]), .Z(n11914) );
  NANDN U13060 ( .A(n11933), .B(n11934), .Z(n11911) );
  AND U13061 ( .A(A[0]), .B(B[478]), .Z(n11934) );
  XOR U13062 ( .A(n11916), .B(n11935), .Z(n11913) );
  NAND U13063 ( .A(A[0]), .B(B[479]), .Z(n11935) );
  NAND U13064 ( .A(B[478]), .B(A[1]), .Z(n11916) );
  NAND U13065 ( .A(n11936), .B(n11937), .Z(n1191) );
  NANDN U13066 ( .A(n11938), .B(n11939), .Z(n11937) );
  OR U13067 ( .A(n11940), .B(n11941), .Z(n11939) );
  NAND U13068 ( .A(n11941), .B(n11940), .Z(n11936) );
  XOR U13069 ( .A(n1193), .B(n1192), .Z(\A1[476] ) );
  XOR U13070 ( .A(n11941), .B(n11942), .Z(n1192) );
  XNOR U13071 ( .A(n11940), .B(n11938), .Z(n11942) );
  AND U13072 ( .A(n11943), .B(n11944), .Z(n11938) );
  NANDN U13073 ( .A(n11945), .B(n11946), .Z(n11944) );
  NANDN U13074 ( .A(n11947), .B(n11948), .Z(n11946) );
  AND U13075 ( .A(B[475]), .B(A[3]), .Z(n11940) );
  XNOR U13076 ( .A(n11930), .B(n11949), .Z(n11941) );
  XNOR U13077 ( .A(n11928), .B(n11931), .Z(n11949) );
  NAND U13078 ( .A(A[2]), .B(B[476]), .Z(n11931) );
  NANDN U13079 ( .A(n11950), .B(n11951), .Z(n11928) );
  AND U13080 ( .A(A[0]), .B(B[477]), .Z(n11951) );
  XOR U13081 ( .A(n11933), .B(n11952), .Z(n11930) );
  NAND U13082 ( .A(A[0]), .B(B[478]), .Z(n11952) );
  NAND U13083 ( .A(B[477]), .B(A[1]), .Z(n11933) );
  NAND U13084 ( .A(n11953), .B(n11954), .Z(n1193) );
  NANDN U13085 ( .A(n11955), .B(n11956), .Z(n11954) );
  OR U13086 ( .A(n11957), .B(n11958), .Z(n11956) );
  NAND U13087 ( .A(n11958), .B(n11957), .Z(n11953) );
  XOR U13088 ( .A(n1195), .B(n1194), .Z(\A1[475] ) );
  XOR U13089 ( .A(n11958), .B(n11959), .Z(n1194) );
  XNOR U13090 ( .A(n11957), .B(n11955), .Z(n11959) );
  AND U13091 ( .A(n11960), .B(n11961), .Z(n11955) );
  NANDN U13092 ( .A(n11962), .B(n11963), .Z(n11961) );
  NANDN U13093 ( .A(n11964), .B(n11965), .Z(n11963) );
  AND U13094 ( .A(B[474]), .B(A[3]), .Z(n11957) );
  XNOR U13095 ( .A(n11947), .B(n11966), .Z(n11958) );
  XNOR U13096 ( .A(n11945), .B(n11948), .Z(n11966) );
  NAND U13097 ( .A(A[2]), .B(B[475]), .Z(n11948) );
  NANDN U13098 ( .A(n11967), .B(n11968), .Z(n11945) );
  AND U13099 ( .A(A[0]), .B(B[476]), .Z(n11968) );
  XOR U13100 ( .A(n11950), .B(n11969), .Z(n11947) );
  NAND U13101 ( .A(A[0]), .B(B[477]), .Z(n11969) );
  NAND U13102 ( .A(B[476]), .B(A[1]), .Z(n11950) );
  NAND U13103 ( .A(n11970), .B(n11971), .Z(n1195) );
  NANDN U13104 ( .A(n11972), .B(n11973), .Z(n11971) );
  OR U13105 ( .A(n11974), .B(n11975), .Z(n11973) );
  NAND U13106 ( .A(n11975), .B(n11974), .Z(n11970) );
  XOR U13107 ( .A(n1197), .B(n1196), .Z(\A1[474] ) );
  XOR U13108 ( .A(n11975), .B(n11976), .Z(n1196) );
  XNOR U13109 ( .A(n11974), .B(n11972), .Z(n11976) );
  AND U13110 ( .A(n11977), .B(n11978), .Z(n11972) );
  NANDN U13111 ( .A(n11979), .B(n11980), .Z(n11978) );
  NANDN U13112 ( .A(n11981), .B(n11982), .Z(n11980) );
  AND U13113 ( .A(B[473]), .B(A[3]), .Z(n11974) );
  XNOR U13114 ( .A(n11964), .B(n11983), .Z(n11975) );
  XNOR U13115 ( .A(n11962), .B(n11965), .Z(n11983) );
  NAND U13116 ( .A(A[2]), .B(B[474]), .Z(n11965) );
  NANDN U13117 ( .A(n11984), .B(n11985), .Z(n11962) );
  AND U13118 ( .A(A[0]), .B(B[475]), .Z(n11985) );
  XOR U13119 ( .A(n11967), .B(n11986), .Z(n11964) );
  NAND U13120 ( .A(A[0]), .B(B[476]), .Z(n11986) );
  NAND U13121 ( .A(B[475]), .B(A[1]), .Z(n11967) );
  NAND U13122 ( .A(n11987), .B(n11988), .Z(n1197) );
  NANDN U13123 ( .A(n11989), .B(n11990), .Z(n11988) );
  OR U13124 ( .A(n11991), .B(n11992), .Z(n11990) );
  NAND U13125 ( .A(n11992), .B(n11991), .Z(n11987) );
  XOR U13126 ( .A(n1199), .B(n1198), .Z(\A1[473] ) );
  XOR U13127 ( .A(n11992), .B(n11993), .Z(n1198) );
  XNOR U13128 ( .A(n11991), .B(n11989), .Z(n11993) );
  AND U13129 ( .A(n11994), .B(n11995), .Z(n11989) );
  NANDN U13130 ( .A(n11996), .B(n11997), .Z(n11995) );
  NANDN U13131 ( .A(n11998), .B(n11999), .Z(n11997) );
  AND U13132 ( .A(B[472]), .B(A[3]), .Z(n11991) );
  XNOR U13133 ( .A(n11981), .B(n12000), .Z(n11992) );
  XNOR U13134 ( .A(n11979), .B(n11982), .Z(n12000) );
  NAND U13135 ( .A(A[2]), .B(B[473]), .Z(n11982) );
  NANDN U13136 ( .A(n12001), .B(n12002), .Z(n11979) );
  AND U13137 ( .A(A[0]), .B(B[474]), .Z(n12002) );
  XOR U13138 ( .A(n11984), .B(n12003), .Z(n11981) );
  NAND U13139 ( .A(A[0]), .B(B[475]), .Z(n12003) );
  NAND U13140 ( .A(B[474]), .B(A[1]), .Z(n11984) );
  NAND U13141 ( .A(n12004), .B(n12005), .Z(n1199) );
  NANDN U13142 ( .A(n12006), .B(n12007), .Z(n12005) );
  OR U13143 ( .A(n12008), .B(n12009), .Z(n12007) );
  NAND U13144 ( .A(n12009), .B(n12008), .Z(n12004) );
  XOR U13145 ( .A(n1201), .B(n1200), .Z(\A1[472] ) );
  XOR U13146 ( .A(n12009), .B(n12010), .Z(n1200) );
  XNOR U13147 ( .A(n12008), .B(n12006), .Z(n12010) );
  AND U13148 ( .A(n12011), .B(n12012), .Z(n12006) );
  NANDN U13149 ( .A(n12013), .B(n12014), .Z(n12012) );
  NANDN U13150 ( .A(n12015), .B(n12016), .Z(n12014) );
  AND U13151 ( .A(B[471]), .B(A[3]), .Z(n12008) );
  XNOR U13152 ( .A(n11998), .B(n12017), .Z(n12009) );
  XNOR U13153 ( .A(n11996), .B(n11999), .Z(n12017) );
  NAND U13154 ( .A(A[2]), .B(B[472]), .Z(n11999) );
  NANDN U13155 ( .A(n12018), .B(n12019), .Z(n11996) );
  AND U13156 ( .A(A[0]), .B(B[473]), .Z(n12019) );
  XOR U13157 ( .A(n12001), .B(n12020), .Z(n11998) );
  NAND U13158 ( .A(A[0]), .B(B[474]), .Z(n12020) );
  NAND U13159 ( .A(B[473]), .B(A[1]), .Z(n12001) );
  NAND U13160 ( .A(n12021), .B(n12022), .Z(n1201) );
  NANDN U13161 ( .A(n12023), .B(n12024), .Z(n12022) );
  OR U13162 ( .A(n12025), .B(n12026), .Z(n12024) );
  NAND U13163 ( .A(n12026), .B(n12025), .Z(n12021) );
  XOR U13164 ( .A(n1203), .B(n1202), .Z(\A1[471] ) );
  XOR U13165 ( .A(n12026), .B(n12027), .Z(n1202) );
  XNOR U13166 ( .A(n12025), .B(n12023), .Z(n12027) );
  AND U13167 ( .A(n12028), .B(n12029), .Z(n12023) );
  NANDN U13168 ( .A(n12030), .B(n12031), .Z(n12029) );
  NANDN U13169 ( .A(n12032), .B(n12033), .Z(n12031) );
  AND U13170 ( .A(B[470]), .B(A[3]), .Z(n12025) );
  XNOR U13171 ( .A(n12015), .B(n12034), .Z(n12026) );
  XNOR U13172 ( .A(n12013), .B(n12016), .Z(n12034) );
  NAND U13173 ( .A(A[2]), .B(B[471]), .Z(n12016) );
  NANDN U13174 ( .A(n12035), .B(n12036), .Z(n12013) );
  AND U13175 ( .A(A[0]), .B(B[472]), .Z(n12036) );
  XOR U13176 ( .A(n12018), .B(n12037), .Z(n12015) );
  NAND U13177 ( .A(A[0]), .B(B[473]), .Z(n12037) );
  NAND U13178 ( .A(B[472]), .B(A[1]), .Z(n12018) );
  NAND U13179 ( .A(n12038), .B(n12039), .Z(n1203) );
  NANDN U13180 ( .A(n12040), .B(n12041), .Z(n12039) );
  OR U13181 ( .A(n12042), .B(n12043), .Z(n12041) );
  NAND U13182 ( .A(n12043), .B(n12042), .Z(n12038) );
  XOR U13183 ( .A(n1205), .B(n1204), .Z(\A1[470] ) );
  XOR U13184 ( .A(n12043), .B(n12044), .Z(n1204) );
  XNOR U13185 ( .A(n12042), .B(n12040), .Z(n12044) );
  AND U13186 ( .A(n12045), .B(n12046), .Z(n12040) );
  NANDN U13187 ( .A(n12047), .B(n12048), .Z(n12046) );
  NANDN U13188 ( .A(n12049), .B(n12050), .Z(n12048) );
  AND U13189 ( .A(B[469]), .B(A[3]), .Z(n12042) );
  XNOR U13190 ( .A(n12032), .B(n12051), .Z(n12043) );
  XNOR U13191 ( .A(n12030), .B(n12033), .Z(n12051) );
  NAND U13192 ( .A(A[2]), .B(B[470]), .Z(n12033) );
  NANDN U13193 ( .A(n12052), .B(n12053), .Z(n12030) );
  AND U13194 ( .A(A[0]), .B(B[471]), .Z(n12053) );
  XOR U13195 ( .A(n12035), .B(n12054), .Z(n12032) );
  NAND U13196 ( .A(A[0]), .B(B[472]), .Z(n12054) );
  NAND U13197 ( .A(B[471]), .B(A[1]), .Z(n12035) );
  NAND U13198 ( .A(n12055), .B(n12056), .Z(n1205) );
  NANDN U13199 ( .A(n12057), .B(n12058), .Z(n12056) );
  OR U13200 ( .A(n12059), .B(n12060), .Z(n12058) );
  NAND U13201 ( .A(n12060), .B(n12059), .Z(n12055) );
  XOR U13202 ( .A(n1187), .B(n1186), .Z(\A1[46] ) );
  XOR U13203 ( .A(n11890), .B(n12061), .Z(n1186) );
  XNOR U13204 ( .A(n11889), .B(n11887), .Z(n12061) );
  AND U13205 ( .A(n12062), .B(n12063), .Z(n11887) );
  NANDN U13206 ( .A(n12064), .B(n12065), .Z(n12063) );
  NANDN U13207 ( .A(n12066), .B(n12067), .Z(n12065) );
  AND U13208 ( .A(B[45]), .B(A[3]), .Z(n11889) );
  XNOR U13209 ( .A(n11879), .B(n12068), .Z(n11890) );
  XNOR U13210 ( .A(n11877), .B(n11880), .Z(n12068) );
  NAND U13211 ( .A(A[2]), .B(B[46]), .Z(n11880) );
  NANDN U13212 ( .A(n12069), .B(n12070), .Z(n11877) );
  AND U13213 ( .A(A[0]), .B(B[47]), .Z(n12070) );
  XOR U13214 ( .A(n11882), .B(n12071), .Z(n11879) );
  NAND U13215 ( .A(A[0]), .B(B[48]), .Z(n12071) );
  NAND U13216 ( .A(B[47]), .B(A[1]), .Z(n11882) );
  NAND U13217 ( .A(n12072), .B(n12073), .Z(n1187) );
  NANDN U13218 ( .A(n12074), .B(n12075), .Z(n12073) );
  OR U13219 ( .A(n12076), .B(n12077), .Z(n12075) );
  NAND U13220 ( .A(n12077), .B(n12076), .Z(n12072) );
  XOR U13221 ( .A(n1207), .B(n1206), .Z(\A1[469] ) );
  XOR U13222 ( .A(n12060), .B(n12078), .Z(n1206) );
  XNOR U13223 ( .A(n12059), .B(n12057), .Z(n12078) );
  AND U13224 ( .A(n12079), .B(n12080), .Z(n12057) );
  NANDN U13225 ( .A(n12081), .B(n12082), .Z(n12080) );
  NANDN U13226 ( .A(n12083), .B(n12084), .Z(n12082) );
  AND U13227 ( .A(B[468]), .B(A[3]), .Z(n12059) );
  XNOR U13228 ( .A(n12049), .B(n12085), .Z(n12060) );
  XNOR U13229 ( .A(n12047), .B(n12050), .Z(n12085) );
  NAND U13230 ( .A(A[2]), .B(B[469]), .Z(n12050) );
  NANDN U13231 ( .A(n12086), .B(n12087), .Z(n12047) );
  AND U13232 ( .A(A[0]), .B(B[470]), .Z(n12087) );
  XOR U13233 ( .A(n12052), .B(n12088), .Z(n12049) );
  NAND U13234 ( .A(A[0]), .B(B[471]), .Z(n12088) );
  NAND U13235 ( .A(B[470]), .B(A[1]), .Z(n12052) );
  NAND U13236 ( .A(n12089), .B(n12090), .Z(n1207) );
  NANDN U13237 ( .A(n12091), .B(n12092), .Z(n12090) );
  OR U13238 ( .A(n12093), .B(n12094), .Z(n12092) );
  NAND U13239 ( .A(n12094), .B(n12093), .Z(n12089) );
  XOR U13240 ( .A(n1211), .B(n1210), .Z(\A1[468] ) );
  XOR U13241 ( .A(n12094), .B(n12095), .Z(n1210) );
  XNOR U13242 ( .A(n12093), .B(n12091), .Z(n12095) );
  AND U13243 ( .A(n12096), .B(n12097), .Z(n12091) );
  NANDN U13244 ( .A(n12098), .B(n12099), .Z(n12097) );
  NANDN U13245 ( .A(n12100), .B(n12101), .Z(n12099) );
  AND U13246 ( .A(B[467]), .B(A[3]), .Z(n12093) );
  XNOR U13247 ( .A(n12083), .B(n12102), .Z(n12094) );
  XNOR U13248 ( .A(n12081), .B(n12084), .Z(n12102) );
  NAND U13249 ( .A(A[2]), .B(B[468]), .Z(n12084) );
  NANDN U13250 ( .A(n12103), .B(n12104), .Z(n12081) );
  AND U13251 ( .A(A[0]), .B(B[469]), .Z(n12104) );
  XOR U13252 ( .A(n12086), .B(n12105), .Z(n12083) );
  NAND U13253 ( .A(A[0]), .B(B[470]), .Z(n12105) );
  NAND U13254 ( .A(B[469]), .B(A[1]), .Z(n12086) );
  NAND U13255 ( .A(n12106), .B(n12107), .Z(n1211) );
  NANDN U13256 ( .A(n12108), .B(n12109), .Z(n12107) );
  OR U13257 ( .A(n12110), .B(n12111), .Z(n12109) );
  NAND U13258 ( .A(n12111), .B(n12110), .Z(n12106) );
  XOR U13259 ( .A(n1213), .B(n1212), .Z(\A1[467] ) );
  XOR U13260 ( .A(n12111), .B(n12112), .Z(n1212) );
  XNOR U13261 ( .A(n12110), .B(n12108), .Z(n12112) );
  AND U13262 ( .A(n12113), .B(n12114), .Z(n12108) );
  NANDN U13263 ( .A(n12115), .B(n12116), .Z(n12114) );
  NANDN U13264 ( .A(n12117), .B(n12118), .Z(n12116) );
  AND U13265 ( .A(B[466]), .B(A[3]), .Z(n12110) );
  XNOR U13266 ( .A(n12100), .B(n12119), .Z(n12111) );
  XNOR U13267 ( .A(n12098), .B(n12101), .Z(n12119) );
  NAND U13268 ( .A(A[2]), .B(B[467]), .Z(n12101) );
  NANDN U13269 ( .A(n12120), .B(n12121), .Z(n12098) );
  AND U13270 ( .A(A[0]), .B(B[468]), .Z(n12121) );
  XOR U13271 ( .A(n12103), .B(n12122), .Z(n12100) );
  NAND U13272 ( .A(A[0]), .B(B[469]), .Z(n12122) );
  NAND U13273 ( .A(B[468]), .B(A[1]), .Z(n12103) );
  NAND U13274 ( .A(n12123), .B(n12124), .Z(n1213) );
  NANDN U13275 ( .A(n12125), .B(n12126), .Z(n12124) );
  OR U13276 ( .A(n12127), .B(n12128), .Z(n12126) );
  NAND U13277 ( .A(n12128), .B(n12127), .Z(n12123) );
  XOR U13278 ( .A(n1215), .B(n1214), .Z(\A1[466] ) );
  XOR U13279 ( .A(n12128), .B(n12129), .Z(n1214) );
  XNOR U13280 ( .A(n12127), .B(n12125), .Z(n12129) );
  AND U13281 ( .A(n12130), .B(n12131), .Z(n12125) );
  NANDN U13282 ( .A(n12132), .B(n12133), .Z(n12131) );
  NANDN U13283 ( .A(n12134), .B(n12135), .Z(n12133) );
  AND U13284 ( .A(B[465]), .B(A[3]), .Z(n12127) );
  XNOR U13285 ( .A(n12117), .B(n12136), .Z(n12128) );
  XNOR U13286 ( .A(n12115), .B(n12118), .Z(n12136) );
  NAND U13287 ( .A(A[2]), .B(B[466]), .Z(n12118) );
  NANDN U13288 ( .A(n12137), .B(n12138), .Z(n12115) );
  AND U13289 ( .A(A[0]), .B(B[467]), .Z(n12138) );
  XOR U13290 ( .A(n12120), .B(n12139), .Z(n12117) );
  NAND U13291 ( .A(A[0]), .B(B[468]), .Z(n12139) );
  NAND U13292 ( .A(B[467]), .B(A[1]), .Z(n12120) );
  NAND U13293 ( .A(n12140), .B(n12141), .Z(n1215) );
  NANDN U13294 ( .A(n12142), .B(n12143), .Z(n12141) );
  OR U13295 ( .A(n12144), .B(n12145), .Z(n12143) );
  NAND U13296 ( .A(n12145), .B(n12144), .Z(n12140) );
  XOR U13297 ( .A(n1217), .B(n1216), .Z(\A1[465] ) );
  XOR U13298 ( .A(n12145), .B(n12146), .Z(n1216) );
  XNOR U13299 ( .A(n12144), .B(n12142), .Z(n12146) );
  AND U13300 ( .A(n12147), .B(n12148), .Z(n12142) );
  NANDN U13301 ( .A(n12149), .B(n12150), .Z(n12148) );
  NANDN U13302 ( .A(n12151), .B(n12152), .Z(n12150) );
  AND U13303 ( .A(B[464]), .B(A[3]), .Z(n12144) );
  XNOR U13304 ( .A(n12134), .B(n12153), .Z(n12145) );
  XNOR U13305 ( .A(n12132), .B(n12135), .Z(n12153) );
  NAND U13306 ( .A(A[2]), .B(B[465]), .Z(n12135) );
  NANDN U13307 ( .A(n12154), .B(n12155), .Z(n12132) );
  AND U13308 ( .A(A[0]), .B(B[466]), .Z(n12155) );
  XOR U13309 ( .A(n12137), .B(n12156), .Z(n12134) );
  NAND U13310 ( .A(A[0]), .B(B[467]), .Z(n12156) );
  NAND U13311 ( .A(B[466]), .B(A[1]), .Z(n12137) );
  NAND U13312 ( .A(n12157), .B(n12158), .Z(n1217) );
  NANDN U13313 ( .A(n12159), .B(n12160), .Z(n12158) );
  OR U13314 ( .A(n12161), .B(n12162), .Z(n12160) );
  NAND U13315 ( .A(n12162), .B(n12161), .Z(n12157) );
  XOR U13316 ( .A(n1219), .B(n1218), .Z(\A1[464] ) );
  XOR U13317 ( .A(n12162), .B(n12163), .Z(n1218) );
  XNOR U13318 ( .A(n12161), .B(n12159), .Z(n12163) );
  AND U13319 ( .A(n12164), .B(n12165), .Z(n12159) );
  NANDN U13320 ( .A(n12166), .B(n12167), .Z(n12165) );
  NANDN U13321 ( .A(n12168), .B(n12169), .Z(n12167) );
  AND U13322 ( .A(B[463]), .B(A[3]), .Z(n12161) );
  XNOR U13323 ( .A(n12151), .B(n12170), .Z(n12162) );
  XNOR U13324 ( .A(n12149), .B(n12152), .Z(n12170) );
  NAND U13325 ( .A(A[2]), .B(B[464]), .Z(n12152) );
  NANDN U13326 ( .A(n12171), .B(n12172), .Z(n12149) );
  AND U13327 ( .A(A[0]), .B(B[465]), .Z(n12172) );
  XOR U13328 ( .A(n12154), .B(n12173), .Z(n12151) );
  NAND U13329 ( .A(A[0]), .B(B[466]), .Z(n12173) );
  NAND U13330 ( .A(B[465]), .B(A[1]), .Z(n12154) );
  NAND U13331 ( .A(n12174), .B(n12175), .Z(n1219) );
  NANDN U13332 ( .A(n12176), .B(n12177), .Z(n12175) );
  OR U13333 ( .A(n12178), .B(n12179), .Z(n12177) );
  NAND U13334 ( .A(n12179), .B(n12178), .Z(n12174) );
  XOR U13335 ( .A(n1221), .B(n1220), .Z(\A1[463] ) );
  XOR U13336 ( .A(n12179), .B(n12180), .Z(n1220) );
  XNOR U13337 ( .A(n12178), .B(n12176), .Z(n12180) );
  AND U13338 ( .A(n12181), .B(n12182), .Z(n12176) );
  NANDN U13339 ( .A(n12183), .B(n12184), .Z(n12182) );
  NANDN U13340 ( .A(n12185), .B(n12186), .Z(n12184) );
  AND U13341 ( .A(B[462]), .B(A[3]), .Z(n12178) );
  XNOR U13342 ( .A(n12168), .B(n12187), .Z(n12179) );
  XNOR U13343 ( .A(n12166), .B(n12169), .Z(n12187) );
  NAND U13344 ( .A(A[2]), .B(B[463]), .Z(n12169) );
  NANDN U13345 ( .A(n12188), .B(n12189), .Z(n12166) );
  AND U13346 ( .A(A[0]), .B(B[464]), .Z(n12189) );
  XOR U13347 ( .A(n12171), .B(n12190), .Z(n12168) );
  NAND U13348 ( .A(A[0]), .B(B[465]), .Z(n12190) );
  NAND U13349 ( .A(B[464]), .B(A[1]), .Z(n12171) );
  NAND U13350 ( .A(n12191), .B(n12192), .Z(n1221) );
  NANDN U13351 ( .A(n12193), .B(n12194), .Z(n12192) );
  OR U13352 ( .A(n12195), .B(n12196), .Z(n12194) );
  NAND U13353 ( .A(n12196), .B(n12195), .Z(n12191) );
  XOR U13354 ( .A(n1223), .B(n1222), .Z(\A1[462] ) );
  XOR U13355 ( .A(n12196), .B(n12197), .Z(n1222) );
  XNOR U13356 ( .A(n12195), .B(n12193), .Z(n12197) );
  AND U13357 ( .A(n12198), .B(n12199), .Z(n12193) );
  NANDN U13358 ( .A(n12200), .B(n12201), .Z(n12199) );
  NANDN U13359 ( .A(n12202), .B(n12203), .Z(n12201) );
  AND U13360 ( .A(B[461]), .B(A[3]), .Z(n12195) );
  XNOR U13361 ( .A(n12185), .B(n12204), .Z(n12196) );
  XNOR U13362 ( .A(n12183), .B(n12186), .Z(n12204) );
  NAND U13363 ( .A(A[2]), .B(B[462]), .Z(n12186) );
  NANDN U13364 ( .A(n12205), .B(n12206), .Z(n12183) );
  AND U13365 ( .A(A[0]), .B(B[463]), .Z(n12206) );
  XOR U13366 ( .A(n12188), .B(n12207), .Z(n12185) );
  NAND U13367 ( .A(A[0]), .B(B[464]), .Z(n12207) );
  NAND U13368 ( .A(B[463]), .B(A[1]), .Z(n12188) );
  NAND U13369 ( .A(n12208), .B(n12209), .Z(n1223) );
  NANDN U13370 ( .A(n12210), .B(n12211), .Z(n12209) );
  OR U13371 ( .A(n12212), .B(n12213), .Z(n12211) );
  NAND U13372 ( .A(n12213), .B(n12212), .Z(n12208) );
  XOR U13373 ( .A(n1225), .B(n1224), .Z(\A1[461] ) );
  XOR U13374 ( .A(n12213), .B(n12214), .Z(n1224) );
  XNOR U13375 ( .A(n12212), .B(n12210), .Z(n12214) );
  AND U13376 ( .A(n12215), .B(n12216), .Z(n12210) );
  NANDN U13377 ( .A(n12217), .B(n12218), .Z(n12216) );
  NANDN U13378 ( .A(n12219), .B(n12220), .Z(n12218) );
  AND U13379 ( .A(B[460]), .B(A[3]), .Z(n12212) );
  XNOR U13380 ( .A(n12202), .B(n12221), .Z(n12213) );
  XNOR U13381 ( .A(n12200), .B(n12203), .Z(n12221) );
  NAND U13382 ( .A(A[2]), .B(B[461]), .Z(n12203) );
  NANDN U13383 ( .A(n12222), .B(n12223), .Z(n12200) );
  AND U13384 ( .A(A[0]), .B(B[462]), .Z(n12223) );
  XOR U13385 ( .A(n12205), .B(n12224), .Z(n12202) );
  NAND U13386 ( .A(A[0]), .B(B[463]), .Z(n12224) );
  NAND U13387 ( .A(B[462]), .B(A[1]), .Z(n12205) );
  NAND U13388 ( .A(n12225), .B(n12226), .Z(n1225) );
  NANDN U13389 ( .A(n12227), .B(n12228), .Z(n12226) );
  OR U13390 ( .A(n12229), .B(n12230), .Z(n12228) );
  NAND U13391 ( .A(n12230), .B(n12229), .Z(n12225) );
  XOR U13392 ( .A(n1227), .B(n1226), .Z(\A1[460] ) );
  XOR U13393 ( .A(n12230), .B(n12231), .Z(n1226) );
  XNOR U13394 ( .A(n12229), .B(n12227), .Z(n12231) );
  AND U13395 ( .A(n12232), .B(n12233), .Z(n12227) );
  NANDN U13396 ( .A(n12234), .B(n12235), .Z(n12233) );
  NANDN U13397 ( .A(n12236), .B(n12237), .Z(n12235) );
  AND U13398 ( .A(B[459]), .B(A[3]), .Z(n12229) );
  XNOR U13399 ( .A(n12219), .B(n12238), .Z(n12230) );
  XNOR U13400 ( .A(n12217), .B(n12220), .Z(n12238) );
  NAND U13401 ( .A(A[2]), .B(B[460]), .Z(n12220) );
  NANDN U13402 ( .A(n12239), .B(n12240), .Z(n12217) );
  AND U13403 ( .A(A[0]), .B(B[461]), .Z(n12240) );
  XOR U13404 ( .A(n12222), .B(n12241), .Z(n12219) );
  NAND U13405 ( .A(A[0]), .B(B[462]), .Z(n12241) );
  NAND U13406 ( .A(B[461]), .B(A[1]), .Z(n12222) );
  NAND U13407 ( .A(n12242), .B(n12243), .Z(n1227) );
  NANDN U13408 ( .A(n12244), .B(n12245), .Z(n12243) );
  OR U13409 ( .A(n12246), .B(n12247), .Z(n12245) );
  NAND U13410 ( .A(n12247), .B(n12246), .Z(n12242) );
  XOR U13411 ( .A(n1209), .B(n1208), .Z(\A1[45] ) );
  XOR U13412 ( .A(n12077), .B(n12248), .Z(n1208) );
  XNOR U13413 ( .A(n12076), .B(n12074), .Z(n12248) );
  AND U13414 ( .A(n12249), .B(n12250), .Z(n12074) );
  NANDN U13415 ( .A(n12251), .B(n12252), .Z(n12250) );
  NANDN U13416 ( .A(n12253), .B(n12254), .Z(n12252) );
  AND U13417 ( .A(B[44]), .B(A[3]), .Z(n12076) );
  XNOR U13418 ( .A(n12066), .B(n12255), .Z(n12077) );
  XNOR U13419 ( .A(n12064), .B(n12067), .Z(n12255) );
  NAND U13420 ( .A(A[2]), .B(B[45]), .Z(n12067) );
  NANDN U13421 ( .A(n12256), .B(n12257), .Z(n12064) );
  AND U13422 ( .A(A[0]), .B(B[46]), .Z(n12257) );
  XOR U13423 ( .A(n12069), .B(n12258), .Z(n12066) );
  NAND U13424 ( .A(A[0]), .B(B[47]), .Z(n12258) );
  NAND U13425 ( .A(B[46]), .B(A[1]), .Z(n12069) );
  NAND U13426 ( .A(n12259), .B(n12260), .Z(n1209) );
  NANDN U13427 ( .A(n12261), .B(n12262), .Z(n12260) );
  OR U13428 ( .A(n12263), .B(n12264), .Z(n12262) );
  NAND U13429 ( .A(n12264), .B(n12263), .Z(n12259) );
  XOR U13430 ( .A(n1229), .B(n1228), .Z(\A1[459] ) );
  XOR U13431 ( .A(n12247), .B(n12265), .Z(n1228) );
  XNOR U13432 ( .A(n12246), .B(n12244), .Z(n12265) );
  AND U13433 ( .A(n12266), .B(n12267), .Z(n12244) );
  NANDN U13434 ( .A(n12268), .B(n12269), .Z(n12267) );
  NANDN U13435 ( .A(n12270), .B(n12271), .Z(n12269) );
  AND U13436 ( .A(B[458]), .B(A[3]), .Z(n12246) );
  XNOR U13437 ( .A(n12236), .B(n12272), .Z(n12247) );
  XNOR U13438 ( .A(n12234), .B(n12237), .Z(n12272) );
  NAND U13439 ( .A(A[2]), .B(B[459]), .Z(n12237) );
  NANDN U13440 ( .A(n12273), .B(n12274), .Z(n12234) );
  AND U13441 ( .A(A[0]), .B(B[460]), .Z(n12274) );
  XOR U13442 ( .A(n12239), .B(n12275), .Z(n12236) );
  NAND U13443 ( .A(A[0]), .B(B[461]), .Z(n12275) );
  NAND U13444 ( .A(B[460]), .B(A[1]), .Z(n12239) );
  NAND U13445 ( .A(n12276), .B(n12277), .Z(n1229) );
  NANDN U13446 ( .A(n12278), .B(n12279), .Z(n12277) );
  OR U13447 ( .A(n12280), .B(n12281), .Z(n12279) );
  NAND U13448 ( .A(n12281), .B(n12280), .Z(n12276) );
  XOR U13449 ( .A(n1233), .B(n1232), .Z(\A1[458] ) );
  XOR U13450 ( .A(n12281), .B(n12282), .Z(n1232) );
  XNOR U13451 ( .A(n12280), .B(n12278), .Z(n12282) );
  AND U13452 ( .A(n12283), .B(n12284), .Z(n12278) );
  NANDN U13453 ( .A(n12285), .B(n12286), .Z(n12284) );
  NANDN U13454 ( .A(n12287), .B(n12288), .Z(n12286) );
  AND U13455 ( .A(B[457]), .B(A[3]), .Z(n12280) );
  XNOR U13456 ( .A(n12270), .B(n12289), .Z(n12281) );
  XNOR U13457 ( .A(n12268), .B(n12271), .Z(n12289) );
  NAND U13458 ( .A(A[2]), .B(B[458]), .Z(n12271) );
  NANDN U13459 ( .A(n12290), .B(n12291), .Z(n12268) );
  AND U13460 ( .A(A[0]), .B(B[459]), .Z(n12291) );
  XOR U13461 ( .A(n12273), .B(n12292), .Z(n12270) );
  NAND U13462 ( .A(A[0]), .B(B[460]), .Z(n12292) );
  NAND U13463 ( .A(B[459]), .B(A[1]), .Z(n12273) );
  NAND U13464 ( .A(n12293), .B(n12294), .Z(n1233) );
  NANDN U13465 ( .A(n12295), .B(n12296), .Z(n12294) );
  OR U13466 ( .A(n12297), .B(n12298), .Z(n12296) );
  NAND U13467 ( .A(n12298), .B(n12297), .Z(n12293) );
  XOR U13468 ( .A(n1235), .B(n1234), .Z(\A1[457] ) );
  XOR U13469 ( .A(n12298), .B(n12299), .Z(n1234) );
  XNOR U13470 ( .A(n12297), .B(n12295), .Z(n12299) );
  AND U13471 ( .A(n12300), .B(n12301), .Z(n12295) );
  NANDN U13472 ( .A(n12302), .B(n12303), .Z(n12301) );
  NANDN U13473 ( .A(n12304), .B(n12305), .Z(n12303) );
  AND U13474 ( .A(B[456]), .B(A[3]), .Z(n12297) );
  XNOR U13475 ( .A(n12287), .B(n12306), .Z(n12298) );
  XNOR U13476 ( .A(n12285), .B(n12288), .Z(n12306) );
  NAND U13477 ( .A(A[2]), .B(B[457]), .Z(n12288) );
  NANDN U13478 ( .A(n12307), .B(n12308), .Z(n12285) );
  AND U13479 ( .A(A[0]), .B(B[458]), .Z(n12308) );
  XOR U13480 ( .A(n12290), .B(n12309), .Z(n12287) );
  NAND U13481 ( .A(A[0]), .B(B[459]), .Z(n12309) );
  NAND U13482 ( .A(B[458]), .B(A[1]), .Z(n12290) );
  NAND U13483 ( .A(n12310), .B(n12311), .Z(n1235) );
  NANDN U13484 ( .A(n12312), .B(n12313), .Z(n12311) );
  OR U13485 ( .A(n12314), .B(n12315), .Z(n12313) );
  NAND U13486 ( .A(n12315), .B(n12314), .Z(n12310) );
  XOR U13487 ( .A(n1237), .B(n1236), .Z(\A1[456] ) );
  XOR U13488 ( .A(n12315), .B(n12316), .Z(n1236) );
  XNOR U13489 ( .A(n12314), .B(n12312), .Z(n12316) );
  AND U13490 ( .A(n12317), .B(n12318), .Z(n12312) );
  NANDN U13491 ( .A(n12319), .B(n12320), .Z(n12318) );
  NANDN U13492 ( .A(n12321), .B(n12322), .Z(n12320) );
  AND U13493 ( .A(B[455]), .B(A[3]), .Z(n12314) );
  XNOR U13494 ( .A(n12304), .B(n12323), .Z(n12315) );
  XNOR U13495 ( .A(n12302), .B(n12305), .Z(n12323) );
  NAND U13496 ( .A(A[2]), .B(B[456]), .Z(n12305) );
  NANDN U13497 ( .A(n12324), .B(n12325), .Z(n12302) );
  AND U13498 ( .A(A[0]), .B(B[457]), .Z(n12325) );
  XOR U13499 ( .A(n12307), .B(n12326), .Z(n12304) );
  NAND U13500 ( .A(A[0]), .B(B[458]), .Z(n12326) );
  NAND U13501 ( .A(B[457]), .B(A[1]), .Z(n12307) );
  NAND U13502 ( .A(n12327), .B(n12328), .Z(n1237) );
  NANDN U13503 ( .A(n12329), .B(n12330), .Z(n12328) );
  OR U13504 ( .A(n12331), .B(n12332), .Z(n12330) );
  NAND U13505 ( .A(n12332), .B(n12331), .Z(n12327) );
  XOR U13506 ( .A(n1239), .B(n1238), .Z(\A1[455] ) );
  XOR U13507 ( .A(n12332), .B(n12333), .Z(n1238) );
  XNOR U13508 ( .A(n12331), .B(n12329), .Z(n12333) );
  AND U13509 ( .A(n12334), .B(n12335), .Z(n12329) );
  NANDN U13510 ( .A(n12336), .B(n12337), .Z(n12335) );
  NANDN U13511 ( .A(n12338), .B(n12339), .Z(n12337) );
  AND U13512 ( .A(B[454]), .B(A[3]), .Z(n12331) );
  XNOR U13513 ( .A(n12321), .B(n12340), .Z(n12332) );
  XNOR U13514 ( .A(n12319), .B(n12322), .Z(n12340) );
  NAND U13515 ( .A(A[2]), .B(B[455]), .Z(n12322) );
  NANDN U13516 ( .A(n12341), .B(n12342), .Z(n12319) );
  AND U13517 ( .A(A[0]), .B(B[456]), .Z(n12342) );
  XOR U13518 ( .A(n12324), .B(n12343), .Z(n12321) );
  NAND U13519 ( .A(A[0]), .B(B[457]), .Z(n12343) );
  NAND U13520 ( .A(B[456]), .B(A[1]), .Z(n12324) );
  NAND U13521 ( .A(n12344), .B(n12345), .Z(n1239) );
  NANDN U13522 ( .A(n12346), .B(n12347), .Z(n12345) );
  OR U13523 ( .A(n12348), .B(n12349), .Z(n12347) );
  NAND U13524 ( .A(n12349), .B(n12348), .Z(n12344) );
  XOR U13525 ( .A(n1241), .B(n1240), .Z(\A1[454] ) );
  XOR U13526 ( .A(n12349), .B(n12350), .Z(n1240) );
  XNOR U13527 ( .A(n12348), .B(n12346), .Z(n12350) );
  AND U13528 ( .A(n12351), .B(n12352), .Z(n12346) );
  NANDN U13529 ( .A(n12353), .B(n12354), .Z(n12352) );
  NANDN U13530 ( .A(n12355), .B(n12356), .Z(n12354) );
  AND U13531 ( .A(B[453]), .B(A[3]), .Z(n12348) );
  XNOR U13532 ( .A(n12338), .B(n12357), .Z(n12349) );
  XNOR U13533 ( .A(n12336), .B(n12339), .Z(n12357) );
  NAND U13534 ( .A(A[2]), .B(B[454]), .Z(n12339) );
  NANDN U13535 ( .A(n12358), .B(n12359), .Z(n12336) );
  AND U13536 ( .A(A[0]), .B(B[455]), .Z(n12359) );
  XOR U13537 ( .A(n12341), .B(n12360), .Z(n12338) );
  NAND U13538 ( .A(A[0]), .B(B[456]), .Z(n12360) );
  NAND U13539 ( .A(B[455]), .B(A[1]), .Z(n12341) );
  NAND U13540 ( .A(n12361), .B(n12362), .Z(n1241) );
  NANDN U13541 ( .A(n12363), .B(n12364), .Z(n12362) );
  OR U13542 ( .A(n12365), .B(n12366), .Z(n12364) );
  NAND U13543 ( .A(n12366), .B(n12365), .Z(n12361) );
  XOR U13544 ( .A(n1243), .B(n1242), .Z(\A1[453] ) );
  XOR U13545 ( .A(n12366), .B(n12367), .Z(n1242) );
  XNOR U13546 ( .A(n12365), .B(n12363), .Z(n12367) );
  AND U13547 ( .A(n12368), .B(n12369), .Z(n12363) );
  NANDN U13548 ( .A(n12370), .B(n12371), .Z(n12369) );
  NANDN U13549 ( .A(n12372), .B(n12373), .Z(n12371) );
  AND U13550 ( .A(B[452]), .B(A[3]), .Z(n12365) );
  XNOR U13551 ( .A(n12355), .B(n12374), .Z(n12366) );
  XNOR U13552 ( .A(n12353), .B(n12356), .Z(n12374) );
  NAND U13553 ( .A(A[2]), .B(B[453]), .Z(n12356) );
  NANDN U13554 ( .A(n12375), .B(n12376), .Z(n12353) );
  AND U13555 ( .A(A[0]), .B(B[454]), .Z(n12376) );
  XOR U13556 ( .A(n12358), .B(n12377), .Z(n12355) );
  NAND U13557 ( .A(A[0]), .B(B[455]), .Z(n12377) );
  NAND U13558 ( .A(B[454]), .B(A[1]), .Z(n12358) );
  NAND U13559 ( .A(n12378), .B(n12379), .Z(n1243) );
  NANDN U13560 ( .A(n12380), .B(n12381), .Z(n12379) );
  OR U13561 ( .A(n12382), .B(n12383), .Z(n12381) );
  NAND U13562 ( .A(n12383), .B(n12382), .Z(n12378) );
  XOR U13563 ( .A(n1245), .B(n1244), .Z(\A1[452] ) );
  XOR U13564 ( .A(n12383), .B(n12384), .Z(n1244) );
  XNOR U13565 ( .A(n12382), .B(n12380), .Z(n12384) );
  AND U13566 ( .A(n12385), .B(n12386), .Z(n12380) );
  NANDN U13567 ( .A(n12387), .B(n12388), .Z(n12386) );
  NANDN U13568 ( .A(n12389), .B(n12390), .Z(n12388) );
  AND U13569 ( .A(B[451]), .B(A[3]), .Z(n12382) );
  XNOR U13570 ( .A(n12372), .B(n12391), .Z(n12383) );
  XNOR U13571 ( .A(n12370), .B(n12373), .Z(n12391) );
  NAND U13572 ( .A(A[2]), .B(B[452]), .Z(n12373) );
  NANDN U13573 ( .A(n12392), .B(n12393), .Z(n12370) );
  AND U13574 ( .A(A[0]), .B(B[453]), .Z(n12393) );
  XOR U13575 ( .A(n12375), .B(n12394), .Z(n12372) );
  NAND U13576 ( .A(A[0]), .B(B[454]), .Z(n12394) );
  NAND U13577 ( .A(B[453]), .B(A[1]), .Z(n12375) );
  NAND U13578 ( .A(n12395), .B(n12396), .Z(n1245) );
  NANDN U13579 ( .A(n12397), .B(n12398), .Z(n12396) );
  OR U13580 ( .A(n12399), .B(n12400), .Z(n12398) );
  NAND U13581 ( .A(n12400), .B(n12399), .Z(n12395) );
  XOR U13582 ( .A(n1247), .B(n1246), .Z(\A1[451] ) );
  XOR U13583 ( .A(n12400), .B(n12401), .Z(n1246) );
  XNOR U13584 ( .A(n12399), .B(n12397), .Z(n12401) );
  AND U13585 ( .A(n12402), .B(n12403), .Z(n12397) );
  NANDN U13586 ( .A(n12404), .B(n12405), .Z(n12403) );
  NANDN U13587 ( .A(n12406), .B(n12407), .Z(n12405) );
  AND U13588 ( .A(B[450]), .B(A[3]), .Z(n12399) );
  XNOR U13589 ( .A(n12389), .B(n12408), .Z(n12400) );
  XNOR U13590 ( .A(n12387), .B(n12390), .Z(n12408) );
  NAND U13591 ( .A(A[2]), .B(B[451]), .Z(n12390) );
  NANDN U13592 ( .A(n12409), .B(n12410), .Z(n12387) );
  AND U13593 ( .A(A[0]), .B(B[452]), .Z(n12410) );
  XOR U13594 ( .A(n12392), .B(n12411), .Z(n12389) );
  NAND U13595 ( .A(A[0]), .B(B[453]), .Z(n12411) );
  NAND U13596 ( .A(B[452]), .B(A[1]), .Z(n12392) );
  NAND U13597 ( .A(n12412), .B(n12413), .Z(n1247) );
  NANDN U13598 ( .A(n12414), .B(n12415), .Z(n12413) );
  OR U13599 ( .A(n12416), .B(n12417), .Z(n12415) );
  NAND U13600 ( .A(n12417), .B(n12416), .Z(n12412) );
  XOR U13601 ( .A(n1249), .B(n1248), .Z(\A1[450] ) );
  XOR U13602 ( .A(n12417), .B(n12418), .Z(n1248) );
  XNOR U13603 ( .A(n12416), .B(n12414), .Z(n12418) );
  AND U13604 ( .A(n12419), .B(n12420), .Z(n12414) );
  NANDN U13605 ( .A(n12421), .B(n12422), .Z(n12420) );
  NANDN U13606 ( .A(n12423), .B(n12424), .Z(n12422) );
  AND U13607 ( .A(B[449]), .B(A[3]), .Z(n12416) );
  XNOR U13608 ( .A(n12406), .B(n12425), .Z(n12417) );
  XNOR U13609 ( .A(n12404), .B(n12407), .Z(n12425) );
  NAND U13610 ( .A(A[2]), .B(B[450]), .Z(n12407) );
  NANDN U13611 ( .A(n12426), .B(n12427), .Z(n12404) );
  AND U13612 ( .A(A[0]), .B(B[451]), .Z(n12427) );
  XOR U13613 ( .A(n12409), .B(n12428), .Z(n12406) );
  NAND U13614 ( .A(A[0]), .B(B[452]), .Z(n12428) );
  NAND U13615 ( .A(B[451]), .B(A[1]), .Z(n12409) );
  NAND U13616 ( .A(n12429), .B(n12430), .Z(n1249) );
  NANDN U13617 ( .A(n12431), .B(n12432), .Z(n12430) );
  OR U13618 ( .A(n12433), .B(n12434), .Z(n12432) );
  NAND U13619 ( .A(n12434), .B(n12433), .Z(n12429) );
  XOR U13620 ( .A(n1231), .B(n1230), .Z(\A1[44] ) );
  XOR U13621 ( .A(n12264), .B(n12435), .Z(n1230) );
  XNOR U13622 ( .A(n12263), .B(n12261), .Z(n12435) );
  AND U13623 ( .A(n12436), .B(n12437), .Z(n12261) );
  NANDN U13624 ( .A(n12438), .B(n12439), .Z(n12437) );
  NANDN U13625 ( .A(n12440), .B(n12441), .Z(n12439) );
  AND U13626 ( .A(B[43]), .B(A[3]), .Z(n12263) );
  XNOR U13627 ( .A(n12253), .B(n12442), .Z(n12264) );
  XNOR U13628 ( .A(n12251), .B(n12254), .Z(n12442) );
  NAND U13629 ( .A(A[2]), .B(B[44]), .Z(n12254) );
  NANDN U13630 ( .A(n12443), .B(n12444), .Z(n12251) );
  AND U13631 ( .A(A[0]), .B(B[45]), .Z(n12444) );
  XOR U13632 ( .A(n12256), .B(n12445), .Z(n12253) );
  NAND U13633 ( .A(A[0]), .B(B[46]), .Z(n12445) );
  NAND U13634 ( .A(B[45]), .B(A[1]), .Z(n12256) );
  NAND U13635 ( .A(n12446), .B(n12447), .Z(n1231) );
  NANDN U13636 ( .A(n12448), .B(n12449), .Z(n12447) );
  OR U13637 ( .A(n12450), .B(n12451), .Z(n12449) );
  NAND U13638 ( .A(n12451), .B(n12450), .Z(n12446) );
  XOR U13639 ( .A(n1251), .B(n1250), .Z(\A1[449] ) );
  XOR U13640 ( .A(n12434), .B(n12452), .Z(n1250) );
  XNOR U13641 ( .A(n12433), .B(n12431), .Z(n12452) );
  AND U13642 ( .A(n12453), .B(n12454), .Z(n12431) );
  NANDN U13643 ( .A(n12455), .B(n12456), .Z(n12454) );
  NANDN U13644 ( .A(n12457), .B(n12458), .Z(n12456) );
  AND U13645 ( .A(B[448]), .B(A[3]), .Z(n12433) );
  XNOR U13646 ( .A(n12423), .B(n12459), .Z(n12434) );
  XNOR U13647 ( .A(n12421), .B(n12424), .Z(n12459) );
  NAND U13648 ( .A(A[2]), .B(B[449]), .Z(n12424) );
  NANDN U13649 ( .A(n12460), .B(n12461), .Z(n12421) );
  AND U13650 ( .A(A[0]), .B(B[450]), .Z(n12461) );
  XOR U13651 ( .A(n12426), .B(n12462), .Z(n12423) );
  NAND U13652 ( .A(A[0]), .B(B[451]), .Z(n12462) );
  NAND U13653 ( .A(B[450]), .B(A[1]), .Z(n12426) );
  NAND U13654 ( .A(n12463), .B(n12464), .Z(n1251) );
  NANDN U13655 ( .A(n12465), .B(n12466), .Z(n12464) );
  OR U13656 ( .A(n12467), .B(n12468), .Z(n12466) );
  NAND U13657 ( .A(n12468), .B(n12467), .Z(n12463) );
  XOR U13658 ( .A(n1255), .B(n1254), .Z(\A1[448] ) );
  XOR U13659 ( .A(n12468), .B(n12469), .Z(n1254) );
  XNOR U13660 ( .A(n12467), .B(n12465), .Z(n12469) );
  AND U13661 ( .A(n12470), .B(n12471), .Z(n12465) );
  NANDN U13662 ( .A(n12472), .B(n12473), .Z(n12471) );
  NANDN U13663 ( .A(n12474), .B(n12475), .Z(n12473) );
  AND U13664 ( .A(B[447]), .B(A[3]), .Z(n12467) );
  XNOR U13665 ( .A(n12457), .B(n12476), .Z(n12468) );
  XNOR U13666 ( .A(n12455), .B(n12458), .Z(n12476) );
  NAND U13667 ( .A(A[2]), .B(B[448]), .Z(n12458) );
  NANDN U13668 ( .A(n12477), .B(n12478), .Z(n12455) );
  AND U13669 ( .A(A[0]), .B(B[449]), .Z(n12478) );
  XOR U13670 ( .A(n12460), .B(n12479), .Z(n12457) );
  NAND U13671 ( .A(A[0]), .B(B[450]), .Z(n12479) );
  NAND U13672 ( .A(B[449]), .B(A[1]), .Z(n12460) );
  NAND U13673 ( .A(n12480), .B(n12481), .Z(n1255) );
  NANDN U13674 ( .A(n12482), .B(n12483), .Z(n12481) );
  OR U13675 ( .A(n12484), .B(n12485), .Z(n12483) );
  NAND U13676 ( .A(n12485), .B(n12484), .Z(n12480) );
  XOR U13677 ( .A(n1257), .B(n1256), .Z(\A1[447] ) );
  XOR U13678 ( .A(n12485), .B(n12486), .Z(n1256) );
  XNOR U13679 ( .A(n12484), .B(n12482), .Z(n12486) );
  AND U13680 ( .A(n12487), .B(n12488), .Z(n12482) );
  NANDN U13681 ( .A(n12489), .B(n12490), .Z(n12488) );
  NANDN U13682 ( .A(n12491), .B(n12492), .Z(n12490) );
  AND U13683 ( .A(B[446]), .B(A[3]), .Z(n12484) );
  XNOR U13684 ( .A(n12474), .B(n12493), .Z(n12485) );
  XNOR U13685 ( .A(n12472), .B(n12475), .Z(n12493) );
  NAND U13686 ( .A(A[2]), .B(B[447]), .Z(n12475) );
  NANDN U13687 ( .A(n12494), .B(n12495), .Z(n12472) );
  AND U13688 ( .A(A[0]), .B(B[448]), .Z(n12495) );
  XOR U13689 ( .A(n12477), .B(n12496), .Z(n12474) );
  NAND U13690 ( .A(A[0]), .B(B[449]), .Z(n12496) );
  NAND U13691 ( .A(B[448]), .B(A[1]), .Z(n12477) );
  NAND U13692 ( .A(n12497), .B(n12498), .Z(n1257) );
  NANDN U13693 ( .A(n12499), .B(n12500), .Z(n12498) );
  OR U13694 ( .A(n12501), .B(n12502), .Z(n12500) );
  NAND U13695 ( .A(n12502), .B(n12501), .Z(n12497) );
  XOR U13696 ( .A(n1259), .B(n1258), .Z(\A1[446] ) );
  XOR U13697 ( .A(n12502), .B(n12503), .Z(n1258) );
  XNOR U13698 ( .A(n12501), .B(n12499), .Z(n12503) );
  AND U13699 ( .A(n12504), .B(n12505), .Z(n12499) );
  NANDN U13700 ( .A(n12506), .B(n12507), .Z(n12505) );
  NANDN U13701 ( .A(n12508), .B(n12509), .Z(n12507) );
  AND U13702 ( .A(B[445]), .B(A[3]), .Z(n12501) );
  XNOR U13703 ( .A(n12491), .B(n12510), .Z(n12502) );
  XNOR U13704 ( .A(n12489), .B(n12492), .Z(n12510) );
  NAND U13705 ( .A(A[2]), .B(B[446]), .Z(n12492) );
  NANDN U13706 ( .A(n12511), .B(n12512), .Z(n12489) );
  AND U13707 ( .A(A[0]), .B(B[447]), .Z(n12512) );
  XOR U13708 ( .A(n12494), .B(n12513), .Z(n12491) );
  NAND U13709 ( .A(A[0]), .B(B[448]), .Z(n12513) );
  NAND U13710 ( .A(B[447]), .B(A[1]), .Z(n12494) );
  NAND U13711 ( .A(n12514), .B(n12515), .Z(n1259) );
  NANDN U13712 ( .A(n12516), .B(n12517), .Z(n12515) );
  OR U13713 ( .A(n12518), .B(n12519), .Z(n12517) );
  NAND U13714 ( .A(n12519), .B(n12518), .Z(n12514) );
  XOR U13715 ( .A(n1261), .B(n1260), .Z(\A1[445] ) );
  XOR U13716 ( .A(n12519), .B(n12520), .Z(n1260) );
  XNOR U13717 ( .A(n12518), .B(n12516), .Z(n12520) );
  AND U13718 ( .A(n12521), .B(n12522), .Z(n12516) );
  NANDN U13719 ( .A(n12523), .B(n12524), .Z(n12522) );
  NANDN U13720 ( .A(n12525), .B(n12526), .Z(n12524) );
  AND U13721 ( .A(B[444]), .B(A[3]), .Z(n12518) );
  XNOR U13722 ( .A(n12508), .B(n12527), .Z(n12519) );
  XNOR U13723 ( .A(n12506), .B(n12509), .Z(n12527) );
  NAND U13724 ( .A(A[2]), .B(B[445]), .Z(n12509) );
  NANDN U13725 ( .A(n12528), .B(n12529), .Z(n12506) );
  AND U13726 ( .A(A[0]), .B(B[446]), .Z(n12529) );
  XOR U13727 ( .A(n12511), .B(n12530), .Z(n12508) );
  NAND U13728 ( .A(A[0]), .B(B[447]), .Z(n12530) );
  NAND U13729 ( .A(B[446]), .B(A[1]), .Z(n12511) );
  NAND U13730 ( .A(n12531), .B(n12532), .Z(n1261) );
  NANDN U13731 ( .A(n12533), .B(n12534), .Z(n12532) );
  OR U13732 ( .A(n12535), .B(n12536), .Z(n12534) );
  NAND U13733 ( .A(n12536), .B(n12535), .Z(n12531) );
  XOR U13734 ( .A(n1263), .B(n1262), .Z(\A1[444] ) );
  XOR U13735 ( .A(n12536), .B(n12537), .Z(n1262) );
  XNOR U13736 ( .A(n12535), .B(n12533), .Z(n12537) );
  AND U13737 ( .A(n12538), .B(n12539), .Z(n12533) );
  NANDN U13738 ( .A(n12540), .B(n12541), .Z(n12539) );
  NANDN U13739 ( .A(n12542), .B(n12543), .Z(n12541) );
  AND U13740 ( .A(B[443]), .B(A[3]), .Z(n12535) );
  XNOR U13741 ( .A(n12525), .B(n12544), .Z(n12536) );
  XNOR U13742 ( .A(n12523), .B(n12526), .Z(n12544) );
  NAND U13743 ( .A(A[2]), .B(B[444]), .Z(n12526) );
  NANDN U13744 ( .A(n12545), .B(n12546), .Z(n12523) );
  AND U13745 ( .A(A[0]), .B(B[445]), .Z(n12546) );
  XOR U13746 ( .A(n12528), .B(n12547), .Z(n12525) );
  NAND U13747 ( .A(A[0]), .B(B[446]), .Z(n12547) );
  NAND U13748 ( .A(B[445]), .B(A[1]), .Z(n12528) );
  NAND U13749 ( .A(n12548), .B(n12549), .Z(n1263) );
  NANDN U13750 ( .A(n12550), .B(n12551), .Z(n12549) );
  OR U13751 ( .A(n12552), .B(n12553), .Z(n12551) );
  NAND U13752 ( .A(n12553), .B(n12552), .Z(n12548) );
  XOR U13753 ( .A(n1265), .B(n1264), .Z(\A1[443] ) );
  XOR U13754 ( .A(n12553), .B(n12554), .Z(n1264) );
  XNOR U13755 ( .A(n12552), .B(n12550), .Z(n12554) );
  AND U13756 ( .A(n12555), .B(n12556), .Z(n12550) );
  NANDN U13757 ( .A(n12557), .B(n12558), .Z(n12556) );
  NANDN U13758 ( .A(n12559), .B(n12560), .Z(n12558) );
  AND U13759 ( .A(B[442]), .B(A[3]), .Z(n12552) );
  XNOR U13760 ( .A(n12542), .B(n12561), .Z(n12553) );
  XNOR U13761 ( .A(n12540), .B(n12543), .Z(n12561) );
  NAND U13762 ( .A(A[2]), .B(B[443]), .Z(n12543) );
  NANDN U13763 ( .A(n12562), .B(n12563), .Z(n12540) );
  AND U13764 ( .A(A[0]), .B(B[444]), .Z(n12563) );
  XOR U13765 ( .A(n12545), .B(n12564), .Z(n12542) );
  NAND U13766 ( .A(A[0]), .B(B[445]), .Z(n12564) );
  NAND U13767 ( .A(B[444]), .B(A[1]), .Z(n12545) );
  NAND U13768 ( .A(n12565), .B(n12566), .Z(n1265) );
  NANDN U13769 ( .A(n12567), .B(n12568), .Z(n12566) );
  OR U13770 ( .A(n12569), .B(n12570), .Z(n12568) );
  NAND U13771 ( .A(n12570), .B(n12569), .Z(n12565) );
  XOR U13772 ( .A(n1267), .B(n1266), .Z(\A1[442] ) );
  XOR U13773 ( .A(n12570), .B(n12571), .Z(n1266) );
  XNOR U13774 ( .A(n12569), .B(n12567), .Z(n12571) );
  AND U13775 ( .A(n12572), .B(n12573), .Z(n12567) );
  NANDN U13776 ( .A(n12574), .B(n12575), .Z(n12573) );
  NANDN U13777 ( .A(n12576), .B(n12577), .Z(n12575) );
  AND U13778 ( .A(B[441]), .B(A[3]), .Z(n12569) );
  XNOR U13779 ( .A(n12559), .B(n12578), .Z(n12570) );
  XNOR U13780 ( .A(n12557), .B(n12560), .Z(n12578) );
  NAND U13781 ( .A(A[2]), .B(B[442]), .Z(n12560) );
  NANDN U13782 ( .A(n12579), .B(n12580), .Z(n12557) );
  AND U13783 ( .A(A[0]), .B(B[443]), .Z(n12580) );
  XOR U13784 ( .A(n12562), .B(n12581), .Z(n12559) );
  NAND U13785 ( .A(A[0]), .B(B[444]), .Z(n12581) );
  NAND U13786 ( .A(B[443]), .B(A[1]), .Z(n12562) );
  NAND U13787 ( .A(n12582), .B(n12583), .Z(n1267) );
  NANDN U13788 ( .A(n12584), .B(n12585), .Z(n12583) );
  OR U13789 ( .A(n12586), .B(n12587), .Z(n12585) );
  NAND U13790 ( .A(n12587), .B(n12586), .Z(n12582) );
  XOR U13791 ( .A(n1269), .B(n1268), .Z(\A1[441] ) );
  XOR U13792 ( .A(n12587), .B(n12588), .Z(n1268) );
  XNOR U13793 ( .A(n12586), .B(n12584), .Z(n12588) );
  AND U13794 ( .A(n12589), .B(n12590), .Z(n12584) );
  NANDN U13795 ( .A(n12591), .B(n12592), .Z(n12590) );
  NANDN U13796 ( .A(n12593), .B(n12594), .Z(n12592) );
  AND U13797 ( .A(B[440]), .B(A[3]), .Z(n12586) );
  XNOR U13798 ( .A(n12576), .B(n12595), .Z(n12587) );
  XNOR U13799 ( .A(n12574), .B(n12577), .Z(n12595) );
  NAND U13800 ( .A(A[2]), .B(B[441]), .Z(n12577) );
  NANDN U13801 ( .A(n12596), .B(n12597), .Z(n12574) );
  AND U13802 ( .A(A[0]), .B(B[442]), .Z(n12597) );
  XOR U13803 ( .A(n12579), .B(n12598), .Z(n12576) );
  NAND U13804 ( .A(A[0]), .B(B[443]), .Z(n12598) );
  NAND U13805 ( .A(B[442]), .B(A[1]), .Z(n12579) );
  NAND U13806 ( .A(n12599), .B(n12600), .Z(n1269) );
  NANDN U13807 ( .A(n12601), .B(n12602), .Z(n12600) );
  OR U13808 ( .A(n12603), .B(n12604), .Z(n12602) );
  NAND U13809 ( .A(n12604), .B(n12603), .Z(n12599) );
  XOR U13810 ( .A(n1271), .B(n1270), .Z(\A1[440] ) );
  XOR U13811 ( .A(n12604), .B(n12605), .Z(n1270) );
  XNOR U13812 ( .A(n12603), .B(n12601), .Z(n12605) );
  AND U13813 ( .A(n12606), .B(n12607), .Z(n12601) );
  NANDN U13814 ( .A(n12608), .B(n12609), .Z(n12607) );
  NANDN U13815 ( .A(n12610), .B(n12611), .Z(n12609) );
  AND U13816 ( .A(B[439]), .B(A[3]), .Z(n12603) );
  XNOR U13817 ( .A(n12593), .B(n12612), .Z(n12604) );
  XNOR U13818 ( .A(n12591), .B(n12594), .Z(n12612) );
  NAND U13819 ( .A(A[2]), .B(B[440]), .Z(n12594) );
  NANDN U13820 ( .A(n12613), .B(n12614), .Z(n12591) );
  AND U13821 ( .A(A[0]), .B(B[441]), .Z(n12614) );
  XOR U13822 ( .A(n12596), .B(n12615), .Z(n12593) );
  NAND U13823 ( .A(A[0]), .B(B[442]), .Z(n12615) );
  NAND U13824 ( .A(B[441]), .B(A[1]), .Z(n12596) );
  NAND U13825 ( .A(n12616), .B(n12617), .Z(n1271) );
  NANDN U13826 ( .A(n12618), .B(n12619), .Z(n12617) );
  OR U13827 ( .A(n12620), .B(n12621), .Z(n12619) );
  NAND U13828 ( .A(n12621), .B(n12620), .Z(n12616) );
  XOR U13829 ( .A(n1253), .B(n1252), .Z(\A1[43] ) );
  XOR U13830 ( .A(n12451), .B(n12622), .Z(n1252) );
  XNOR U13831 ( .A(n12450), .B(n12448), .Z(n12622) );
  AND U13832 ( .A(n12623), .B(n12624), .Z(n12448) );
  NANDN U13833 ( .A(n12625), .B(n12626), .Z(n12624) );
  NANDN U13834 ( .A(n12627), .B(n12628), .Z(n12626) );
  AND U13835 ( .A(B[42]), .B(A[3]), .Z(n12450) );
  XNOR U13836 ( .A(n12440), .B(n12629), .Z(n12451) );
  XNOR U13837 ( .A(n12438), .B(n12441), .Z(n12629) );
  NAND U13838 ( .A(A[2]), .B(B[43]), .Z(n12441) );
  NANDN U13839 ( .A(n12630), .B(n12631), .Z(n12438) );
  AND U13840 ( .A(A[0]), .B(B[44]), .Z(n12631) );
  XOR U13841 ( .A(n12443), .B(n12632), .Z(n12440) );
  NAND U13842 ( .A(A[0]), .B(B[45]), .Z(n12632) );
  NAND U13843 ( .A(B[44]), .B(A[1]), .Z(n12443) );
  NAND U13844 ( .A(n12633), .B(n12634), .Z(n1253) );
  NANDN U13845 ( .A(n12635), .B(n12636), .Z(n12634) );
  OR U13846 ( .A(n12637), .B(n12638), .Z(n12636) );
  NAND U13847 ( .A(n12638), .B(n12637), .Z(n12633) );
  XOR U13848 ( .A(n1273), .B(n1272), .Z(\A1[439] ) );
  XOR U13849 ( .A(n12621), .B(n12639), .Z(n1272) );
  XNOR U13850 ( .A(n12620), .B(n12618), .Z(n12639) );
  AND U13851 ( .A(n12640), .B(n12641), .Z(n12618) );
  NANDN U13852 ( .A(n12642), .B(n12643), .Z(n12641) );
  NANDN U13853 ( .A(n12644), .B(n12645), .Z(n12643) );
  AND U13854 ( .A(B[438]), .B(A[3]), .Z(n12620) );
  XNOR U13855 ( .A(n12610), .B(n12646), .Z(n12621) );
  XNOR U13856 ( .A(n12608), .B(n12611), .Z(n12646) );
  NAND U13857 ( .A(A[2]), .B(B[439]), .Z(n12611) );
  NANDN U13858 ( .A(n12647), .B(n12648), .Z(n12608) );
  AND U13859 ( .A(A[0]), .B(B[440]), .Z(n12648) );
  XOR U13860 ( .A(n12613), .B(n12649), .Z(n12610) );
  NAND U13861 ( .A(A[0]), .B(B[441]), .Z(n12649) );
  NAND U13862 ( .A(B[440]), .B(A[1]), .Z(n12613) );
  NAND U13863 ( .A(n12650), .B(n12651), .Z(n1273) );
  NANDN U13864 ( .A(n12652), .B(n12653), .Z(n12651) );
  OR U13865 ( .A(n12654), .B(n12655), .Z(n12653) );
  NAND U13866 ( .A(n12655), .B(n12654), .Z(n12650) );
  XOR U13867 ( .A(n1277), .B(n1276), .Z(\A1[438] ) );
  XOR U13868 ( .A(n12655), .B(n12656), .Z(n1276) );
  XNOR U13869 ( .A(n12654), .B(n12652), .Z(n12656) );
  AND U13870 ( .A(n12657), .B(n12658), .Z(n12652) );
  NANDN U13871 ( .A(n12659), .B(n12660), .Z(n12658) );
  NANDN U13872 ( .A(n12661), .B(n12662), .Z(n12660) );
  AND U13873 ( .A(B[437]), .B(A[3]), .Z(n12654) );
  XNOR U13874 ( .A(n12644), .B(n12663), .Z(n12655) );
  XNOR U13875 ( .A(n12642), .B(n12645), .Z(n12663) );
  NAND U13876 ( .A(A[2]), .B(B[438]), .Z(n12645) );
  NANDN U13877 ( .A(n12664), .B(n12665), .Z(n12642) );
  AND U13878 ( .A(A[0]), .B(B[439]), .Z(n12665) );
  XOR U13879 ( .A(n12647), .B(n12666), .Z(n12644) );
  NAND U13880 ( .A(A[0]), .B(B[440]), .Z(n12666) );
  NAND U13881 ( .A(B[439]), .B(A[1]), .Z(n12647) );
  NAND U13882 ( .A(n12667), .B(n12668), .Z(n1277) );
  NANDN U13883 ( .A(n12669), .B(n12670), .Z(n12668) );
  OR U13884 ( .A(n12671), .B(n12672), .Z(n12670) );
  NAND U13885 ( .A(n12672), .B(n12671), .Z(n12667) );
  XOR U13886 ( .A(n1279), .B(n1278), .Z(\A1[437] ) );
  XOR U13887 ( .A(n12672), .B(n12673), .Z(n1278) );
  XNOR U13888 ( .A(n12671), .B(n12669), .Z(n12673) );
  AND U13889 ( .A(n12674), .B(n12675), .Z(n12669) );
  NANDN U13890 ( .A(n12676), .B(n12677), .Z(n12675) );
  NANDN U13891 ( .A(n12678), .B(n12679), .Z(n12677) );
  AND U13892 ( .A(B[436]), .B(A[3]), .Z(n12671) );
  XNOR U13893 ( .A(n12661), .B(n12680), .Z(n12672) );
  XNOR U13894 ( .A(n12659), .B(n12662), .Z(n12680) );
  NAND U13895 ( .A(A[2]), .B(B[437]), .Z(n12662) );
  NANDN U13896 ( .A(n12681), .B(n12682), .Z(n12659) );
  AND U13897 ( .A(A[0]), .B(B[438]), .Z(n12682) );
  XOR U13898 ( .A(n12664), .B(n12683), .Z(n12661) );
  NAND U13899 ( .A(A[0]), .B(B[439]), .Z(n12683) );
  NAND U13900 ( .A(B[438]), .B(A[1]), .Z(n12664) );
  NAND U13901 ( .A(n12684), .B(n12685), .Z(n1279) );
  NANDN U13902 ( .A(n12686), .B(n12687), .Z(n12685) );
  OR U13903 ( .A(n12688), .B(n12689), .Z(n12687) );
  NAND U13904 ( .A(n12689), .B(n12688), .Z(n12684) );
  XOR U13905 ( .A(n1281), .B(n1280), .Z(\A1[436] ) );
  XOR U13906 ( .A(n12689), .B(n12690), .Z(n1280) );
  XNOR U13907 ( .A(n12688), .B(n12686), .Z(n12690) );
  AND U13908 ( .A(n12691), .B(n12692), .Z(n12686) );
  NANDN U13909 ( .A(n12693), .B(n12694), .Z(n12692) );
  NANDN U13910 ( .A(n12695), .B(n12696), .Z(n12694) );
  AND U13911 ( .A(B[435]), .B(A[3]), .Z(n12688) );
  XNOR U13912 ( .A(n12678), .B(n12697), .Z(n12689) );
  XNOR U13913 ( .A(n12676), .B(n12679), .Z(n12697) );
  NAND U13914 ( .A(A[2]), .B(B[436]), .Z(n12679) );
  NANDN U13915 ( .A(n12698), .B(n12699), .Z(n12676) );
  AND U13916 ( .A(A[0]), .B(B[437]), .Z(n12699) );
  XOR U13917 ( .A(n12681), .B(n12700), .Z(n12678) );
  NAND U13918 ( .A(A[0]), .B(B[438]), .Z(n12700) );
  NAND U13919 ( .A(B[437]), .B(A[1]), .Z(n12681) );
  NAND U13920 ( .A(n12701), .B(n12702), .Z(n1281) );
  NANDN U13921 ( .A(n12703), .B(n12704), .Z(n12702) );
  OR U13922 ( .A(n12705), .B(n12706), .Z(n12704) );
  NAND U13923 ( .A(n12706), .B(n12705), .Z(n12701) );
  XOR U13924 ( .A(n1283), .B(n1282), .Z(\A1[435] ) );
  XOR U13925 ( .A(n12706), .B(n12707), .Z(n1282) );
  XNOR U13926 ( .A(n12705), .B(n12703), .Z(n12707) );
  AND U13927 ( .A(n12708), .B(n12709), .Z(n12703) );
  NANDN U13928 ( .A(n12710), .B(n12711), .Z(n12709) );
  NANDN U13929 ( .A(n12712), .B(n12713), .Z(n12711) );
  AND U13930 ( .A(B[434]), .B(A[3]), .Z(n12705) );
  XNOR U13931 ( .A(n12695), .B(n12714), .Z(n12706) );
  XNOR U13932 ( .A(n12693), .B(n12696), .Z(n12714) );
  NAND U13933 ( .A(A[2]), .B(B[435]), .Z(n12696) );
  NANDN U13934 ( .A(n12715), .B(n12716), .Z(n12693) );
  AND U13935 ( .A(A[0]), .B(B[436]), .Z(n12716) );
  XOR U13936 ( .A(n12698), .B(n12717), .Z(n12695) );
  NAND U13937 ( .A(A[0]), .B(B[437]), .Z(n12717) );
  NAND U13938 ( .A(B[436]), .B(A[1]), .Z(n12698) );
  NAND U13939 ( .A(n12718), .B(n12719), .Z(n1283) );
  NANDN U13940 ( .A(n12720), .B(n12721), .Z(n12719) );
  OR U13941 ( .A(n12722), .B(n12723), .Z(n12721) );
  NAND U13942 ( .A(n12723), .B(n12722), .Z(n12718) );
  XOR U13943 ( .A(n1285), .B(n1284), .Z(\A1[434] ) );
  XOR U13944 ( .A(n12723), .B(n12724), .Z(n1284) );
  XNOR U13945 ( .A(n12722), .B(n12720), .Z(n12724) );
  AND U13946 ( .A(n12725), .B(n12726), .Z(n12720) );
  NANDN U13947 ( .A(n12727), .B(n12728), .Z(n12726) );
  NANDN U13948 ( .A(n12729), .B(n12730), .Z(n12728) );
  AND U13949 ( .A(B[433]), .B(A[3]), .Z(n12722) );
  XNOR U13950 ( .A(n12712), .B(n12731), .Z(n12723) );
  XNOR U13951 ( .A(n12710), .B(n12713), .Z(n12731) );
  NAND U13952 ( .A(A[2]), .B(B[434]), .Z(n12713) );
  NANDN U13953 ( .A(n12732), .B(n12733), .Z(n12710) );
  AND U13954 ( .A(A[0]), .B(B[435]), .Z(n12733) );
  XOR U13955 ( .A(n12715), .B(n12734), .Z(n12712) );
  NAND U13956 ( .A(A[0]), .B(B[436]), .Z(n12734) );
  NAND U13957 ( .A(B[435]), .B(A[1]), .Z(n12715) );
  NAND U13958 ( .A(n12735), .B(n12736), .Z(n1285) );
  NANDN U13959 ( .A(n12737), .B(n12738), .Z(n12736) );
  OR U13960 ( .A(n12739), .B(n12740), .Z(n12738) );
  NAND U13961 ( .A(n12740), .B(n12739), .Z(n12735) );
  XOR U13962 ( .A(n1287), .B(n1286), .Z(\A1[433] ) );
  XOR U13963 ( .A(n12740), .B(n12741), .Z(n1286) );
  XNOR U13964 ( .A(n12739), .B(n12737), .Z(n12741) );
  AND U13965 ( .A(n12742), .B(n12743), .Z(n12737) );
  NANDN U13966 ( .A(n12744), .B(n12745), .Z(n12743) );
  NANDN U13967 ( .A(n12746), .B(n12747), .Z(n12745) );
  AND U13968 ( .A(B[432]), .B(A[3]), .Z(n12739) );
  XNOR U13969 ( .A(n12729), .B(n12748), .Z(n12740) );
  XNOR U13970 ( .A(n12727), .B(n12730), .Z(n12748) );
  NAND U13971 ( .A(A[2]), .B(B[433]), .Z(n12730) );
  NANDN U13972 ( .A(n12749), .B(n12750), .Z(n12727) );
  AND U13973 ( .A(A[0]), .B(B[434]), .Z(n12750) );
  XOR U13974 ( .A(n12732), .B(n12751), .Z(n12729) );
  NAND U13975 ( .A(A[0]), .B(B[435]), .Z(n12751) );
  NAND U13976 ( .A(B[434]), .B(A[1]), .Z(n12732) );
  NAND U13977 ( .A(n12752), .B(n12753), .Z(n1287) );
  NANDN U13978 ( .A(n12754), .B(n12755), .Z(n12753) );
  OR U13979 ( .A(n12756), .B(n12757), .Z(n12755) );
  NAND U13980 ( .A(n12757), .B(n12756), .Z(n12752) );
  XOR U13981 ( .A(n1289), .B(n1288), .Z(\A1[432] ) );
  XOR U13982 ( .A(n12757), .B(n12758), .Z(n1288) );
  XNOR U13983 ( .A(n12756), .B(n12754), .Z(n12758) );
  AND U13984 ( .A(n12759), .B(n12760), .Z(n12754) );
  NANDN U13985 ( .A(n12761), .B(n12762), .Z(n12760) );
  NANDN U13986 ( .A(n12763), .B(n12764), .Z(n12762) );
  AND U13987 ( .A(B[431]), .B(A[3]), .Z(n12756) );
  XNOR U13988 ( .A(n12746), .B(n12765), .Z(n12757) );
  XNOR U13989 ( .A(n12744), .B(n12747), .Z(n12765) );
  NAND U13990 ( .A(A[2]), .B(B[432]), .Z(n12747) );
  NANDN U13991 ( .A(n12766), .B(n12767), .Z(n12744) );
  AND U13992 ( .A(A[0]), .B(B[433]), .Z(n12767) );
  XOR U13993 ( .A(n12749), .B(n12768), .Z(n12746) );
  NAND U13994 ( .A(A[0]), .B(B[434]), .Z(n12768) );
  NAND U13995 ( .A(B[433]), .B(A[1]), .Z(n12749) );
  NAND U13996 ( .A(n12769), .B(n12770), .Z(n1289) );
  NANDN U13997 ( .A(n12771), .B(n12772), .Z(n12770) );
  OR U13998 ( .A(n12773), .B(n12774), .Z(n12772) );
  NAND U13999 ( .A(n12774), .B(n12773), .Z(n12769) );
  XOR U14000 ( .A(n1291), .B(n1290), .Z(\A1[431] ) );
  XOR U14001 ( .A(n12774), .B(n12775), .Z(n1290) );
  XNOR U14002 ( .A(n12773), .B(n12771), .Z(n12775) );
  AND U14003 ( .A(n12776), .B(n12777), .Z(n12771) );
  NANDN U14004 ( .A(n12778), .B(n12779), .Z(n12777) );
  NANDN U14005 ( .A(n12780), .B(n12781), .Z(n12779) );
  AND U14006 ( .A(B[430]), .B(A[3]), .Z(n12773) );
  XNOR U14007 ( .A(n12763), .B(n12782), .Z(n12774) );
  XNOR U14008 ( .A(n12761), .B(n12764), .Z(n12782) );
  NAND U14009 ( .A(A[2]), .B(B[431]), .Z(n12764) );
  NANDN U14010 ( .A(n12783), .B(n12784), .Z(n12761) );
  AND U14011 ( .A(A[0]), .B(B[432]), .Z(n12784) );
  XOR U14012 ( .A(n12766), .B(n12785), .Z(n12763) );
  NAND U14013 ( .A(A[0]), .B(B[433]), .Z(n12785) );
  NAND U14014 ( .A(B[432]), .B(A[1]), .Z(n12766) );
  NAND U14015 ( .A(n12786), .B(n12787), .Z(n1291) );
  NANDN U14016 ( .A(n12788), .B(n12789), .Z(n12787) );
  OR U14017 ( .A(n12790), .B(n12791), .Z(n12789) );
  NAND U14018 ( .A(n12791), .B(n12790), .Z(n12786) );
  XOR U14019 ( .A(n1293), .B(n1292), .Z(\A1[430] ) );
  XOR U14020 ( .A(n12791), .B(n12792), .Z(n1292) );
  XNOR U14021 ( .A(n12790), .B(n12788), .Z(n12792) );
  AND U14022 ( .A(n12793), .B(n12794), .Z(n12788) );
  NANDN U14023 ( .A(n12795), .B(n12796), .Z(n12794) );
  NANDN U14024 ( .A(n12797), .B(n12798), .Z(n12796) );
  AND U14025 ( .A(B[429]), .B(A[3]), .Z(n12790) );
  XNOR U14026 ( .A(n12780), .B(n12799), .Z(n12791) );
  XNOR U14027 ( .A(n12778), .B(n12781), .Z(n12799) );
  NAND U14028 ( .A(A[2]), .B(B[430]), .Z(n12781) );
  NANDN U14029 ( .A(n12800), .B(n12801), .Z(n12778) );
  AND U14030 ( .A(A[0]), .B(B[431]), .Z(n12801) );
  XOR U14031 ( .A(n12783), .B(n12802), .Z(n12780) );
  NAND U14032 ( .A(A[0]), .B(B[432]), .Z(n12802) );
  NAND U14033 ( .A(B[431]), .B(A[1]), .Z(n12783) );
  NAND U14034 ( .A(n12803), .B(n12804), .Z(n1293) );
  NANDN U14035 ( .A(n12805), .B(n12806), .Z(n12804) );
  OR U14036 ( .A(n12807), .B(n12808), .Z(n12806) );
  NAND U14037 ( .A(n12808), .B(n12807), .Z(n12803) );
  XOR U14038 ( .A(n1275), .B(n1274), .Z(\A1[42] ) );
  XOR U14039 ( .A(n12638), .B(n12809), .Z(n1274) );
  XNOR U14040 ( .A(n12637), .B(n12635), .Z(n12809) );
  AND U14041 ( .A(n12810), .B(n12811), .Z(n12635) );
  NANDN U14042 ( .A(n12812), .B(n12813), .Z(n12811) );
  NANDN U14043 ( .A(n12814), .B(n12815), .Z(n12813) );
  AND U14044 ( .A(B[41]), .B(A[3]), .Z(n12637) );
  XNOR U14045 ( .A(n12627), .B(n12816), .Z(n12638) );
  XNOR U14046 ( .A(n12625), .B(n12628), .Z(n12816) );
  NAND U14047 ( .A(A[2]), .B(B[42]), .Z(n12628) );
  NANDN U14048 ( .A(n12817), .B(n12818), .Z(n12625) );
  AND U14049 ( .A(A[0]), .B(B[43]), .Z(n12818) );
  XOR U14050 ( .A(n12630), .B(n12819), .Z(n12627) );
  NAND U14051 ( .A(A[0]), .B(B[44]), .Z(n12819) );
  NAND U14052 ( .A(B[43]), .B(A[1]), .Z(n12630) );
  NAND U14053 ( .A(n12820), .B(n12821), .Z(n1275) );
  NANDN U14054 ( .A(n12822), .B(n12823), .Z(n12821) );
  OR U14055 ( .A(n12824), .B(n12825), .Z(n12823) );
  NAND U14056 ( .A(n12825), .B(n12824), .Z(n12820) );
  XOR U14057 ( .A(n1295), .B(n1294), .Z(\A1[429] ) );
  XOR U14058 ( .A(n12808), .B(n12826), .Z(n1294) );
  XNOR U14059 ( .A(n12807), .B(n12805), .Z(n12826) );
  AND U14060 ( .A(n12827), .B(n12828), .Z(n12805) );
  NANDN U14061 ( .A(n12829), .B(n12830), .Z(n12828) );
  NANDN U14062 ( .A(n12831), .B(n12832), .Z(n12830) );
  AND U14063 ( .A(B[428]), .B(A[3]), .Z(n12807) );
  XNOR U14064 ( .A(n12797), .B(n12833), .Z(n12808) );
  XNOR U14065 ( .A(n12795), .B(n12798), .Z(n12833) );
  NAND U14066 ( .A(A[2]), .B(B[429]), .Z(n12798) );
  NANDN U14067 ( .A(n12834), .B(n12835), .Z(n12795) );
  AND U14068 ( .A(A[0]), .B(B[430]), .Z(n12835) );
  XOR U14069 ( .A(n12800), .B(n12836), .Z(n12797) );
  NAND U14070 ( .A(A[0]), .B(B[431]), .Z(n12836) );
  NAND U14071 ( .A(B[430]), .B(A[1]), .Z(n12800) );
  NAND U14072 ( .A(n12837), .B(n12838), .Z(n1295) );
  NANDN U14073 ( .A(n12839), .B(n12840), .Z(n12838) );
  OR U14074 ( .A(n12841), .B(n12842), .Z(n12840) );
  NAND U14075 ( .A(n12842), .B(n12841), .Z(n12837) );
  XOR U14076 ( .A(n1299), .B(n1298), .Z(\A1[428] ) );
  XOR U14077 ( .A(n12842), .B(n12843), .Z(n1298) );
  XNOR U14078 ( .A(n12841), .B(n12839), .Z(n12843) );
  AND U14079 ( .A(n12844), .B(n12845), .Z(n12839) );
  NANDN U14080 ( .A(n12846), .B(n12847), .Z(n12845) );
  NANDN U14081 ( .A(n12848), .B(n12849), .Z(n12847) );
  AND U14082 ( .A(B[427]), .B(A[3]), .Z(n12841) );
  XNOR U14083 ( .A(n12831), .B(n12850), .Z(n12842) );
  XNOR U14084 ( .A(n12829), .B(n12832), .Z(n12850) );
  NAND U14085 ( .A(A[2]), .B(B[428]), .Z(n12832) );
  NANDN U14086 ( .A(n12851), .B(n12852), .Z(n12829) );
  AND U14087 ( .A(A[0]), .B(B[429]), .Z(n12852) );
  XOR U14088 ( .A(n12834), .B(n12853), .Z(n12831) );
  NAND U14089 ( .A(A[0]), .B(B[430]), .Z(n12853) );
  NAND U14090 ( .A(B[429]), .B(A[1]), .Z(n12834) );
  NAND U14091 ( .A(n12854), .B(n12855), .Z(n1299) );
  NANDN U14092 ( .A(n12856), .B(n12857), .Z(n12855) );
  OR U14093 ( .A(n12858), .B(n12859), .Z(n12857) );
  NAND U14094 ( .A(n12859), .B(n12858), .Z(n12854) );
  XOR U14095 ( .A(n1301), .B(n1300), .Z(\A1[427] ) );
  XOR U14096 ( .A(n12859), .B(n12860), .Z(n1300) );
  XNOR U14097 ( .A(n12858), .B(n12856), .Z(n12860) );
  AND U14098 ( .A(n12861), .B(n12862), .Z(n12856) );
  NANDN U14099 ( .A(n12863), .B(n12864), .Z(n12862) );
  NANDN U14100 ( .A(n12865), .B(n12866), .Z(n12864) );
  AND U14101 ( .A(B[426]), .B(A[3]), .Z(n12858) );
  XNOR U14102 ( .A(n12848), .B(n12867), .Z(n12859) );
  XNOR U14103 ( .A(n12846), .B(n12849), .Z(n12867) );
  NAND U14104 ( .A(A[2]), .B(B[427]), .Z(n12849) );
  NANDN U14105 ( .A(n12868), .B(n12869), .Z(n12846) );
  AND U14106 ( .A(A[0]), .B(B[428]), .Z(n12869) );
  XOR U14107 ( .A(n12851), .B(n12870), .Z(n12848) );
  NAND U14108 ( .A(A[0]), .B(B[429]), .Z(n12870) );
  NAND U14109 ( .A(B[428]), .B(A[1]), .Z(n12851) );
  NAND U14110 ( .A(n12871), .B(n12872), .Z(n1301) );
  NANDN U14111 ( .A(n12873), .B(n12874), .Z(n12872) );
  OR U14112 ( .A(n12875), .B(n12876), .Z(n12874) );
  NAND U14113 ( .A(n12876), .B(n12875), .Z(n12871) );
  XOR U14114 ( .A(n1303), .B(n1302), .Z(\A1[426] ) );
  XOR U14115 ( .A(n12876), .B(n12877), .Z(n1302) );
  XNOR U14116 ( .A(n12875), .B(n12873), .Z(n12877) );
  AND U14117 ( .A(n12878), .B(n12879), .Z(n12873) );
  NANDN U14118 ( .A(n12880), .B(n12881), .Z(n12879) );
  NANDN U14119 ( .A(n12882), .B(n12883), .Z(n12881) );
  AND U14120 ( .A(B[425]), .B(A[3]), .Z(n12875) );
  XNOR U14121 ( .A(n12865), .B(n12884), .Z(n12876) );
  XNOR U14122 ( .A(n12863), .B(n12866), .Z(n12884) );
  NAND U14123 ( .A(A[2]), .B(B[426]), .Z(n12866) );
  NANDN U14124 ( .A(n12885), .B(n12886), .Z(n12863) );
  AND U14125 ( .A(A[0]), .B(B[427]), .Z(n12886) );
  XOR U14126 ( .A(n12868), .B(n12887), .Z(n12865) );
  NAND U14127 ( .A(A[0]), .B(B[428]), .Z(n12887) );
  NAND U14128 ( .A(B[427]), .B(A[1]), .Z(n12868) );
  NAND U14129 ( .A(n12888), .B(n12889), .Z(n1303) );
  NANDN U14130 ( .A(n12890), .B(n12891), .Z(n12889) );
  OR U14131 ( .A(n12892), .B(n12893), .Z(n12891) );
  NAND U14132 ( .A(n12893), .B(n12892), .Z(n12888) );
  XOR U14133 ( .A(n1305), .B(n1304), .Z(\A1[425] ) );
  XOR U14134 ( .A(n12893), .B(n12894), .Z(n1304) );
  XNOR U14135 ( .A(n12892), .B(n12890), .Z(n12894) );
  AND U14136 ( .A(n12895), .B(n12896), .Z(n12890) );
  NANDN U14137 ( .A(n12897), .B(n12898), .Z(n12896) );
  NANDN U14138 ( .A(n12899), .B(n12900), .Z(n12898) );
  AND U14139 ( .A(B[424]), .B(A[3]), .Z(n12892) );
  XNOR U14140 ( .A(n12882), .B(n12901), .Z(n12893) );
  XNOR U14141 ( .A(n12880), .B(n12883), .Z(n12901) );
  NAND U14142 ( .A(A[2]), .B(B[425]), .Z(n12883) );
  NANDN U14143 ( .A(n12902), .B(n12903), .Z(n12880) );
  AND U14144 ( .A(A[0]), .B(B[426]), .Z(n12903) );
  XOR U14145 ( .A(n12885), .B(n12904), .Z(n12882) );
  NAND U14146 ( .A(A[0]), .B(B[427]), .Z(n12904) );
  NAND U14147 ( .A(B[426]), .B(A[1]), .Z(n12885) );
  NAND U14148 ( .A(n12905), .B(n12906), .Z(n1305) );
  NANDN U14149 ( .A(n12907), .B(n12908), .Z(n12906) );
  OR U14150 ( .A(n12909), .B(n12910), .Z(n12908) );
  NAND U14151 ( .A(n12910), .B(n12909), .Z(n12905) );
  XOR U14152 ( .A(n1307), .B(n1306), .Z(\A1[424] ) );
  XOR U14153 ( .A(n12910), .B(n12911), .Z(n1306) );
  XNOR U14154 ( .A(n12909), .B(n12907), .Z(n12911) );
  AND U14155 ( .A(n12912), .B(n12913), .Z(n12907) );
  NANDN U14156 ( .A(n12914), .B(n12915), .Z(n12913) );
  NANDN U14157 ( .A(n12916), .B(n12917), .Z(n12915) );
  AND U14158 ( .A(B[423]), .B(A[3]), .Z(n12909) );
  XNOR U14159 ( .A(n12899), .B(n12918), .Z(n12910) );
  XNOR U14160 ( .A(n12897), .B(n12900), .Z(n12918) );
  NAND U14161 ( .A(A[2]), .B(B[424]), .Z(n12900) );
  NANDN U14162 ( .A(n12919), .B(n12920), .Z(n12897) );
  AND U14163 ( .A(A[0]), .B(B[425]), .Z(n12920) );
  XOR U14164 ( .A(n12902), .B(n12921), .Z(n12899) );
  NAND U14165 ( .A(A[0]), .B(B[426]), .Z(n12921) );
  NAND U14166 ( .A(B[425]), .B(A[1]), .Z(n12902) );
  NAND U14167 ( .A(n12922), .B(n12923), .Z(n1307) );
  NANDN U14168 ( .A(n12924), .B(n12925), .Z(n12923) );
  OR U14169 ( .A(n12926), .B(n12927), .Z(n12925) );
  NAND U14170 ( .A(n12927), .B(n12926), .Z(n12922) );
  XOR U14171 ( .A(n1309), .B(n1308), .Z(\A1[423] ) );
  XOR U14172 ( .A(n12927), .B(n12928), .Z(n1308) );
  XNOR U14173 ( .A(n12926), .B(n12924), .Z(n12928) );
  AND U14174 ( .A(n12929), .B(n12930), .Z(n12924) );
  NANDN U14175 ( .A(n12931), .B(n12932), .Z(n12930) );
  NANDN U14176 ( .A(n12933), .B(n12934), .Z(n12932) );
  AND U14177 ( .A(B[422]), .B(A[3]), .Z(n12926) );
  XNOR U14178 ( .A(n12916), .B(n12935), .Z(n12927) );
  XNOR U14179 ( .A(n12914), .B(n12917), .Z(n12935) );
  NAND U14180 ( .A(A[2]), .B(B[423]), .Z(n12917) );
  NANDN U14181 ( .A(n12936), .B(n12937), .Z(n12914) );
  AND U14182 ( .A(A[0]), .B(B[424]), .Z(n12937) );
  XOR U14183 ( .A(n12919), .B(n12938), .Z(n12916) );
  NAND U14184 ( .A(A[0]), .B(B[425]), .Z(n12938) );
  NAND U14185 ( .A(B[424]), .B(A[1]), .Z(n12919) );
  NAND U14186 ( .A(n12939), .B(n12940), .Z(n1309) );
  NANDN U14187 ( .A(n12941), .B(n12942), .Z(n12940) );
  OR U14188 ( .A(n12943), .B(n12944), .Z(n12942) );
  NAND U14189 ( .A(n12944), .B(n12943), .Z(n12939) );
  XOR U14190 ( .A(n1311), .B(n1310), .Z(\A1[422] ) );
  XOR U14191 ( .A(n12944), .B(n12945), .Z(n1310) );
  XNOR U14192 ( .A(n12943), .B(n12941), .Z(n12945) );
  AND U14193 ( .A(n12946), .B(n12947), .Z(n12941) );
  NANDN U14194 ( .A(n12948), .B(n12949), .Z(n12947) );
  NANDN U14195 ( .A(n12950), .B(n12951), .Z(n12949) );
  AND U14196 ( .A(B[421]), .B(A[3]), .Z(n12943) );
  XNOR U14197 ( .A(n12933), .B(n12952), .Z(n12944) );
  XNOR U14198 ( .A(n12931), .B(n12934), .Z(n12952) );
  NAND U14199 ( .A(A[2]), .B(B[422]), .Z(n12934) );
  NANDN U14200 ( .A(n12953), .B(n12954), .Z(n12931) );
  AND U14201 ( .A(A[0]), .B(B[423]), .Z(n12954) );
  XOR U14202 ( .A(n12936), .B(n12955), .Z(n12933) );
  NAND U14203 ( .A(A[0]), .B(B[424]), .Z(n12955) );
  NAND U14204 ( .A(B[423]), .B(A[1]), .Z(n12936) );
  NAND U14205 ( .A(n12956), .B(n12957), .Z(n1311) );
  NANDN U14206 ( .A(n12958), .B(n12959), .Z(n12957) );
  OR U14207 ( .A(n12960), .B(n12961), .Z(n12959) );
  NAND U14208 ( .A(n12961), .B(n12960), .Z(n12956) );
  XOR U14209 ( .A(n1313), .B(n1312), .Z(\A1[421] ) );
  XOR U14210 ( .A(n12961), .B(n12962), .Z(n1312) );
  XNOR U14211 ( .A(n12960), .B(n12958), .Z(n12962) );
  AND U14212 ( .A(n12963), .B(n12964), .Z(n12958) );
  NANDN U14213 ( .A(n12965), .B(n12966), .Z(n12964) );
  NANDN U14214 ( .A(n12967), .B(n12968), .Z(n12966) );
  AND U14215 ( .A(B[420]), .B(A[3]), .Z(n12960) );
  XNOR U14216 ( .A(n12950), .B(n12969), .Z(n12961) );
  XNOR U14217 ( .A(n12948), .B(n12951), .Z(n12969) );
  NAND U14218 ( .A(A[2]), .B(B[421]), .Z(n12951) );
  NANDN U14219 ( .A(n12970), .B(n12971), .Z(n12948) );
  AND U14220 ( .A(A[0]), .B(B[422]), .Z(n12971) );
  XOR U14221 ( .A(n12953), .B(n12972), .Z(n12950) );
  NAND U14222 ( .A(A[0]), .B(B[423]), .Z(n12972) );
  NAND U14223 ( .A(B[422]), .B(A[1]), .Z(n12953) );
  NAND U14224 ( .A(n12973), .B(n12974), .Z(n1313) );
  NANDN U14225 ( .A(n12975), .B(n12976), .Z(n12974) );
  OR U14226 ( .A(n12977), .B(n12978), .Z(n12976) );
  NAND U14227 ( .A(n12978), .B(n12977), .Z(n12973) );
  XOR U14228 ( .A(n1315), .B(n1314), .Z(\A1[420] ) );
  XOR U14229 ( .A(n12978), .B(n12979), .Z(n1314) );
  XNOR U14230 ( .A(n12977), .B(n12975), .Z(n12979) );
  AND U14231 ( .A(n12980), .B(n12981), .Z(n12975) );
  NANDN U14232 ( .A(n12982), .B(n12983), .Z(n12981) );
  NANDN U14233 ( .A(n12984), .B(n12985), .Z(n12983) );
  AND U14234 ( .A(B[419]), .B(A[3]), .Z(n12977) );
  XNOR U14235 ( .A(n12967), .B(n12986), .Z(n12978) );
  XNOR U14236 ( .A(n12965), .B(n12968), .Z(n12986) );
  NAND U14237 ( .A(A[2]), .B(B[420]), .Z(n12968) );
  NANDN U14238 ( .A(n12987), .B(n12988), .Z(n12965) );
  AND U14239 ( .A(A[0]), .B(B[421]), .Z(n12988) );
  XOR U14240 ( .A(n12970), .B(n12989), .Z(n12967) );
  NAND U14241 ( .A(A[0]), .B(B[422]), .Z(n12989) );
  NAND U14242 ( .A(B[421]), .B(A[1]), .Z(n12970) );
  NAND U14243 ( .A(n12990), .B(n12991), .Z(n1315) );
  NANDN U14244 ( .A(n12992), .B(n12993), .Z(n12991) );
  OR U14245 ( .A(n12994), .B(n12995), .Z(n12993) );
  NAND U14246 ( .A(n12995), .B(n12994), .Z(n12990) );
  XOR U14247 ( .A(n1297), .B(n1296), .Z(\A1[41] ) );
  XOR U14248 ( .A(n12825), .B(n12996), .Z(n1296) );
  XNOR U14249 ( .A(n12824), .B(n12822), .Z(n12996) );
  AND U14250 ( .A(n12997), .B(n12998), .Z(n12822) );
  NANDN U14251 ( .A(n12999), .B(n13000), .Z(n12998) );
  NANDN U14252 ( .A(n13001), .B(n13002), .Z(n13000) );
  AND U14253 ( .A(B[40]), .B(A[3]), .Z(n12824) );
  XNOR U14254 ( .A(n12814), .B(n13003), .Z(n12825) );
  XNOR U14255 ( .A(n12812), .B(n12815), .Z(n13003) );
  NAND U14256 ( .A(A[2]), .B(B[41]), .Z(n12815) );
  NANDN U14257 ( .A(n13004), .B(n13005), .Z(n12812) );
  AND U14258 ( .A(A[0]), .B(B[42]), .Z(n13005) );
  XOR U14259 ( .A(n12817), .B(n13006), .Z(n12814) );
  NAND U14260 ( .A(A[0]), .B(B[43]), .Z(n13006) );
  NAND U14261 ( .A(B[42]), .B(A[1]), .Z(n12817) );
  NAND U14262 ( .A(n13007), .B(n13008), .Z(n1297) );
  NANDN U14263 ( .A(n13009), .B(n13010), .Z(n13008) );
  OR U14264 ( .A(n13011), .B(n13012), .Z(n13010) );
  NAND U14265 ( .A(n13012), .B(n13011), .Z(n13007) );
  XOR U14266 ( .A(n1317), .B(n1316), .Z(\A1[419] ) );
  XOR U14267 ( .A(n12995), .B(n13013), .Z(n1316) );
  XNOR U14268 ( .A(n12994), .B(n12992), .Z(n13013) );
  AND U14269 ( .A(n13014), .B(n13015), .Z(n12992) );
  NANDN U14270 ( .A(n13016), .B(n13017), .Z(n13015) );
  NANDN U14271 ( .A(n13018), .B(n13019), .Z(n13017) );
  AND U14272 ( .A(B[418]), .B(A[3]), .Z(n12994) );
  XNOR U14273 ( .A(n12984), .B(n13020), .Z(n12995) );
  XNOR U14274 ( .A(n12982), .B(n12985), .Z(n13020) );
  NAND U14275 ( .A(A[2]), .B(B[419]), .Z(n12985) );
  NANDN U14276 ( .A(n13021), .B(n13022), .Z(n12982) );
  AND U14277 ( .A(A[0]), .B(B[420]), .Z(n13022) );
  XOR U14278 ( .A(n12987), .B(n13023), .Z(n12984) );
  NAND U14279 ( .A(A[0]), .B(B[421]), .Z(n13023) );
  NAND U14280 ( .A(B[420]), .B(A[1]), .Z(n12987) );
  NAND U14281 ( .A(n13024), .B(n13025), .Z(n1317) );
  NANDN U14282 ( .A(n13026), .B(n13027), .Z(n13025) );
  OR U14283 ( .A(n13028), .B(n13029), .Z(n13027) );
  NAND U14284 ( .A(n13029), .B(n13028), .Z(n13024) );
  XOR U14285 ( .A(n1321), .B(n1320), .Z(\A1[418] ) );
  XOR U14286 ( .A(n13029), .B(n13030), .Z(n1320) );
  XNOR U14287 ( .A(n13028), .B(n13026), .Z(n13030) );
  AND U14288 ( .A(n13031), .B(n13032), .Z(n13026) );
  NANDN U14289 ( .A(n13033), .B(n13034), .Z(n13032) );
  NANDN U14290 ( .A(n13035), .B(n13036), .Z(n13034) );
  AND U14291 ( .A(B[417]), .B(A[3]), .Z(n13028) );
  XNOR U14292 ( .A(n13018), .B(n13037), .Z(n13029) );
  XNOR U14293 ( .A(n13016), .B(n13019), .Z(n13037) );
  NAND U14294 ( .A(A[2]), .B(B[418]), .Z(n13019) );
  NANDN U14295 ( .A(n13038), .B(n13039), .Z(n13016) );
  AND U14296 ( .A(A[0]), .B(B[419]), .Z(n13039) );
  XOR U14297 ( .A(n13021), .B(n13040), .Z(n13018) );
  NAND U14298 ( .A(A[0]), .B(B[420]), .Z(n13040) );
  NAND U14299 ( .A(B[419]), .B(A[1]), .Z(n13021) );
  NAND U14300 ( .A(n13041), .B(n13042), .Z(n1321) );
  NANDN U14301 ( .A(n13043), .B(n13044), .Z(n13042) );
  OR U14302 ( .A(n13045), .B(n13046), .Z(n13044) );
  NAND U14303 ( .A(n13046), .B(n13045), .Z(n13041) );
  XOR U14304 ( .A(n1323), .B(n1322), .Z(\A1[417] ) );
  XOR U14305 ( .A(n13046), .B(n13047), .Z(n1322) );
  XNOR U14306 ( .A(n13045), .B(n13043), .Z(n13047) );
  AND U14307 ( .A(n13048), .B(n13049), .Z(n13043) );
  NANDN U14308 ( .A(n13050), .B(n13051), .Z(n13049) );
  NANDN U14309 ( .A(n13052), .B(n13053), .Z(n13051) );
  AND U14310 ( .A(B[416]), .B(A[3]), .Z(n13045) );
  XNOR U14311 ( .A(n13035), .B(n13054), .Z(n13046) );
  XNOR U14312 ( .A(n13033), .B(n13036), .Z(n13054) );
  NAND U14313 ( .A(A[2]), .B(B[417]), .Z(n13036) );
  NANDN U14314 ( .A(n13055), .B(n13056), .Z(n13033) );
  AND U14315 ( .A(A[0]), .B(B[418]), .Z(n13056) );
  XOR U14316 ( .A(n13038), .B(n13057), .Z(n13035) );
  NAND U14317 ( .A(A[0]), .B(B[419]), .Z(n13057) );
  NAND U14318 ( .A(B[418]), .B(A[1]), .Z(n13038) );
  NAND U14319 ( .A(n13058), .B(n13059), .Z(n1323) );
  NANDN U14320 ( .A(n13060), .B(n13061), .Z(n13059) );
  OR U14321 ( .A(n13062), .B(n13063), .Z(n13061) );
  NAND U14322 ( .A(n13063), .B(n13062), .Z(n13058) );
  XOR U14323 ( .A(n1325), .B(n1324), .Z(\A1[416] ) );
  XOR U14324 ( .A(n13063), .B(n13064), .Z(n1324) );
  XNOR U14325 ( .A(n13062), .B(n13060), .Z(n13064) );
  AND U14326 ( .A(n13065), .B(n13066), .Z(n13060) );
  NANDN U14327 ( .A(n13067), .B(n13068), .Z(n13066) );
  NANDN U14328 ( .A(n13069), .B(n13070), .Z(n13068) );
  AND U14329 ( .A(B[415]), .B(A[3]), .Z(n13062) );
  XNOR U14330 ( .A(n13052), .B(n13071), .Z(n13063) );
  XNOR U14331 ( .A(n13050), .B(n13053), .Z(n13071) );
  NAND U14332 ( .A(A[2]), .B(B[416]), .Z(n13053) );
  NANDN U14333 ( .A(n13072), .B(n13073), .Z(n13050) );
  AND U14334 ( .A(A[0]), .B(B[417]), .Z(n13073) );
  XOR U14335 ( .A(n13055), .B(n13074), .Z(n13052) );
  NAND U14336 ( .A(A[0]), .B(B[418]), .Z(n13074) );
  NAND U14337 ( .A(B[417]), .B(A[1]), .Z(n13055) );
  NAND U14338 ( .A(n13075), .B(n13076), .Z(n1325) );
  NANDN U14339 ( .A(n13077), .B(n13078), .Z(n13076) );
  OR U14340 ( .A(n13079), .B(n13080), .Z(n13078) );
  NAND U14341 ( .A(n13080), .B(n13079), .Z(n13075) );
  XOR U14342 ( .A(n1327), .B(n1326), .Z(\A1[415] ) );
  XOR U14343 ( .A(n13080), .B(n13081), .Z(n1326) );
  XNOR U14344 ( .A(n13079), .B(n13077), .Z(n13081) );
  AND U14345 ( .A(n13082), .B(n13083), .Z(n13077) );
  NANDN U14346 ( .A(n13084), .B(n13085), .Z(n13083) );
  NANDN U14347 ( .A(n13086), .B(n13087), .Z(n13085) );
  AND U14348 ( .A(B[414]), .B(A[3]), .Z(n13079) );
  XNOR U14349 ( .A(n13069), .B(n13088), .Z(n13080) );
  XNOR U14350 ( .A(n13067), .B(n13070), .Z(n13088) );
  NAND U14351 ( .A(A[2]), .B(B[415]), .Z(n13070) );
  NANDN U14352 ( .A(n13089), .B(n13090), .Z(n13067) );
  AND U14353 ( .A(A[0]), .B(B[416]), .Z(n13090) );
  XOR U14354 ( .A(n13072), .B(n13091), .Z(n13069) );
  NAND U14355 ( .A(A[0]), .B(B[417]), .Z(n13091) );
  NAND U14356 ( .A(B[416]), .B(A[1]), .Z(n13072) );
  NAND U14357 ( .A(n13092), .B(n13093), .Z(n1327) );
  NANDN U14358 ( .A(n13094), .B(n13095), .Z(n13093) );
  OR U14359 ( .A(n13096), .B(n13097), .Z(n13095) );
  NAND U14360 ( .A(n13097), .B(n13096), .Z(n13092) );
  XOR U14361 ( .A(n1329), .B(n1328), .Z(\A1[414] ) );
  XOR U14362 ( .A(n13097), .B(n13098), .Z(n1328) );
  XNOR U14363 ( .A(n13096), .B(n13094), .Z(n13098) );
  AND U14364 ( .A(n13099), .B(n13100), .Z(n13094) );
  NANDN U14365 ( .A(n13101), .B(n13102), .Z(n13100) );
  NANDN U14366 ( .A(n13103), .B(n13104), .Z(n13102) );
  AND U14367 ( .A(B[413]), .B(A[3]), .Z(n13096) );
  XNOR U14368 ( .A(n13086), .B(n13105), .Z(n13097) );
  XNOR U14369 ( .A(n13084), .B(n13087), .Z(n13105) );
  NAND U14370 ( .A(A[2]), .B(B[414]), .Z(n13087) );
  NANDN U14371 ( .A(n13106), .B(n13107), .Z(n13084) );
  AND U14372 ( .A(A[0]), .B(B[415]), .Z(n13107) );
  XOR U14373 ( .A(n13089), .B(n13108), .Z(n13086) );
  NAND U14374 ( .A(A[0]), .B(B[416]), .Z(n13108) );
  NAND U14375 ( .A(B[415]), .B(A[1]), .Z(n13089) );
  NAND U14376 ( .A(n13109), .B(n13110), .Z(n1329) );
  NANDN U14377 ( .A(n13111), .B(n13112), .Z(n13110) );
  OR U14378 ( .A(n13113), .B(n13114), .Z(n13112) );
  NAND U14379 ( .A(n13114), .B(n13113), .Z(n13109) );
  XOR U14380 ( .A(n1331), .B(n1330), .Z(\A1[413] ) );
  XOR U14381 ( .A(n13114), .B(n13115), .Z(n1330) );
  XNOR U14382 ( .A(n13113), .B(n13111), .Z(n13115) );
  AND U14383 ( .A(n13116), .B(n13117), .Z(n13111) );
  NANDN U14384 ( .A(n13118), .B(n13119), .Z(n13117) );
  NANDN U14385 ( .A(n13120), .B(n13121), .Z(n13119) );
  AND U14386 ( .A(B[412]), .B(A[3]), .Z(n13113) );
  XNOR U14387 ( .A(n13103), .B(n13122), .Z(n13114) );
  XNOR U14388 ( .A(n13101), .B(n13104), .Z(n13122) );
  NAND U14389 ( .A(A[2]), .B(B[413]), .Z(n13104) );
  NANDN U14390 ( .A(n13123), .B(n13124), .Z(n13101) );
  AND U14391 ( .A(A[0]), .B(B[414]), .Z(n13124) );
  XOR U14392 ( .A(n13106), .B(n13125), .Z(n13103) );
  NAND U14393 ( .A(A[0]), .B(B[415]), .Z(n13125) );
  NAND U14394 ( .A(B[414]), .B(A[1]), .Z(n13106) );
  NAND U14395 ( .A(n13126), .B(n13127), .Z(n1331) );
  NANDN U14396 ( .A(n13128), .B(n13129), .Z(n13127) );
  OR U14397 ( .A(n13130), .B(n13131), .Z(n13129) );
  NAND U14398 ( .A(n13131), .B(n13130), .Z(n13126) );
  XOR U14399 ( .A(n1333), .B(n1332), .Z(\A1[412] ) );
  XOR U14400 ( .A(n13131), .B(n13132), .Z(n1332) );
  XNOR U14401 ( .A(n13130), .B(n13128), .Z(n13132) );
  AND U14402 ( .A(n13133), .B(n13134), .Z(n13128) );
  NANDN U14403 ( .A(n13135), .B(n13136), .Z(n13134) );
  NANDN U14404 ( .A(n13137), .B(n13138), .Z(n13136) );
  AND U14405 ( .A(B[411]), .B(A[3]), .Z(n13130) );
  XNOR U14406 ( .A(n13120), .B(n13139), .Z(n13131) );
  XNOR U14407 ( .A(n13118), .B(n13121), .Z(n13139) );
  NAND U14408 ( .A(A[2]), .B(B[412]), .Z(n13121) );
  NANDN U14409 ( .A(n13140), .B(n13141), .Z(n13118) );
  AND U14410 ( .A(A[0]), .B(B[413]), .Z(n13141) );
  XOR U14411 ( .A(n13123), .B(n13142), .Z(n13120) );
  NAND U14412 ( .A(A[0]), .B(B[414]), .Z(n13142) );
  NAND U14413 ( .A(B[413]), .B(A[1]), .Z(n13123) );
  NAND U14414 ( .A(n13143), .B(n13144), .Z(n1333) );
  NANDN U14415 ( .A(n13145), .B(n13146), .Z(n13144) );
  OR U14416 ( .A(n13147), .B(n13148), .Z(n13146) );
  NAND U14417 ( .A(n13148), .B(n13147), .Z(n13143) );
  XOR U14418 ( .A(n1335), .B(n1334), .Z(\A1[411] ) );
  XOR U14419 ( .A(n13148), .B(n13149), .Z(n1334) );
  XNOR U14420 ( .A(n13147), .B(n13145), .Z(n13149) );
  AND U14421 ( .A(n13150), .B(n13151), .Z(n13145) );
  NANDN U14422 ( .A(n13152), .B(n13153), .Z(n13151) );
  NANDN U14423 ( .A(n13154), .B(n13155), .Z(n13153) );
  AND U14424 ( .A(B[410]), .B(A[3]), .Z(n13147) );
  XNOR U14425 ( .A(n13137), .B(n13156), .Z(n13148) );
  XNOR U14426 ( .A(n13135), .B(n13138), .Z(n13156) );
  NAND U14427 ( .A(A[2]), .B(B[411]), .Z(n13138) );
  NANDN U14428 ( .A(n13157), .B(n13158), .Z(n13135) );
  AND U14429 ( .A(A[0]), .B(B[412]), .Z(n13158) );
  XOR U14430 ( .A(n13140), .B(n13159), .Z(n13137) );
  NAND U14431 ( .A(A[0]), .B(B[413]), .Z(n13159) );
  NAND U14432 ( .A(B[412]), .B(A[1]), .Z(n13140) );
  NAND U14433 ( .A(n13160), .B(n13161), .Z(n1335) );
  NANDN U14434 ( .A(n13162), .B(n13163), .Z(n13161) );
  OR U14435 ( .A(n13164), .B(n13165), .Z(n13163) );
  NAND U14436 ( .A(n13165), .B(n13164), .Z(n13160) );
  XOR U14437 ( .A(n1337), .B(n1336), .Z(\A1[410] ) );
  XOR U14438 ( .A(n13165), .B(n13166), .Z(n1336) );
  XNOR U14439 ( .A(n13164), .B(n13162), .Z(n13166) );
  AND U14440 ( .A(n13167), .B(n13168), .Z(n13162) );
  NANDN U14441 ( .A(n13169), .B(n13170), .Z(n13168) );
  NANDN U14442 ( .A(n13171), .B(n13172), .Z(n13170) );
  AND U14443 ( .A(B[409]), .B(A[3]), .Z(n13164) );
  XNOR U14444 ( .A(n13154), .B(n13173), .Z(n13165) );
  XNOR U14445 ( .A(n13152), .B(n13155), .Z(n13173) );
  NAND U14446 ( .A(A[2]), .B(B[410]), .Z(n13155) );
  NANDN U14447 ( .A(n13174), .B(n13175), .Z(n13152) );
  AND U14448 ( .A(A[0]), .B(B[411]), .Z(n13175) );
  XOR U14449 ( .A(n13157), .B(n13176), .Z(n13154) );
  NAND U14450 ( .A(A[0]), .B(B[412]), .Z(n13176) );
  NAND U14451 ( .A(B[411]), .B(A[1]), .Z(n13157) );
  NAND U14452 ( .A(n13177), .B(n13178), .Z(n1337) );
  NANDN U14453 ( .A(n13179), .B(n13180), .Z(n13178) );
  OR U14454 ( .A(n13181), .B(n13182), .Z(n13180) );
  NAND U14455 ( .A(n13182), .B(n13181), .Z(n13177) );
  XOR U14456 ( .A(n1319), .B(n1318), .Z(\A1[40] ) );
  XOR U14457 ( .A(n13012), .B(n13183), .Z(n1318) );
  XNOR U14458 ( .A(n13011), .B(n13009), .Z(n13183) );
  AND U14459 ( .A(n13184), .B(n13185), .Z(n13009) );
  NANDN U14460 ( .A(n13186), .B(n13187), .Z(n13185) );
  NANDN U14461 ( .A(n13188), .B(n13189), .Z(n13187) );
  AND U14462 ( .A(B[39]), .B(A[3]), .Z(n13011) );
  XNOR U14463 ( .A(n13001), .B(n13190), .Z(n13012) );
  XNOR U14464 ( .A(n12999), .B(n13002), .Z(n13190) );
  NAND U14465 ( .A(A[2]), .B(B[40]), .Z(n13002) );
  NANDN U14466 ( .A(n13191), .B(n13192), .Z(n12999) );
  AND U14467 ( .A(A[0]), .B(B[41]), .Z(n13192) );
  XOR U14468 ( .A(n13004), .B(n13193), .Z(n13001) );
  NAND U14469 ( .A(A[0]), .B(B[42]), .Z(n13193) );
  NAND U14470 ( .A(B[41]), .B(A[1]), .Z(n13004) );
  NAND U14471 ( .A(n13194), .B(n13195), .Z(n1319) );
  NANDN U14472 ( .A(n13196), .B(n13197), .Z(n13195) );
  OR U14473 ( .A(n13198), .B(n13199), .Z(n13197) );
  NAND U14474 ( .A(n13199), .B(n13198), .Z(n13194) );
  XOR U14475 ( .A(n1339), .B(n1338), .Z(\A1[409] ) );
  XOR U14476 ( .A(n13182), .B(n13200), .Z(n1338) );
  XNOR U14477 ( .A(n13181), .B(n13179), .Z(n13200) );
  AND U14478 ( .A(n13201), .B(n13202), .Z(n13179) );
  NANDN U14479 ( .A(n13203), .B(n13204), .Z(n13202) );
  NANDN U14480 ( .A(n13205), .B(n13206), .Z(n13204) );
  AND U14481 ( .A(B[408]), .B(A[3]), .Z(n13181) );
  XNOR U14482 ( .A(n13171), .B(n13207), .Z(n13182) );
  XNOR U14483 ( .A(n13169), .B(n13172), .Z(n13207) );
  NAND U14484 ( .A(A[2]), .B(B[409]), .Z(n13172) );
  NANDN U14485 ( .A(n13208), .B(n13209), .Z(n13169) );
  AND U14486 ( .A(A[0]), .B(B[410]), .Z(n13209) );
  XOR U14487 ( .A(n13174), .B(n13210), .Z(n13171) );
  NAND U14488 ( .A(A[0]), .B(B[411]), .Z(n13210) );
  NAND U14489 ( .A(B[410]), .B(A[1]), .Z(n13174) );
  NAND U14490 ( .A(n13211), .B(n13212), .Z(n1339) );
  NANDN U14491 ( .A(n13213), .B(n13214), .Z(n13212) );
  OR U14492 ( .A(n13215), .B(n13216), .Z(n13214) );
  NAND U14493 ( .A(n13216), .B(n13215), .Z(n13211) );
  XOR U14494 ( .A(n1343), .B(n1342), .Z(\A1[408] ) );
  XOR U14495 ( .A(n13216), .B(n13217), .Z(n1342) );
  XNOR U14496 ( .A(n13215), .B(n13213), .Z(n13217) );
  AND U14497 ( .A(n13218), .B(n13219), .Z(n13213) );
  NANDN U14498 ( .A(n13220), .B(n13221), .Z(n13219) );
  NANDN U14499 ( .A(n13222), .B(n13223), .Z(n13221) );
  AND U14500 ( .A(B[407]), .B(A[3]), .Z(n13215) );
  XNOR U14501 ( .A(n13205), .B(n13224), .Z(n13216) );
  XNOR U14502 ( .A(n13203), .B(n13206), .Z(n13224) );
  NAND U14503 ( .A(A[2]), .B(B[408]), .Z(n13206) );
  NANDN U14504 ( .A(n13225), .B(n13226), .Z(n13203) );
  AND U14505 ( .A(A[0]), .B(B[409]), .Z(n13226) );
  XOR U14506 ( .A(n13208), .B(n13227), .Z(n13205) );
  NAND U14507 ( .A(A[0]), .B(B[410]), .Z(n13227) );
  NAND U14508 ( .A(B[409]), .B(A[1]), .Z(n13208) );
  NAND U14509 ( .A(n13228), .B(n13229), .Z(n1343) );
  NANDN U14510 ( .A(n13230), .B(n13231), .Z(n13229) );
  OR U14511 ( .A(n13232), .B(n13233), .Z(n13231) );
  NAND U14512 ( .A(n13233), .B(n13232), .Z(n13228) );
  XOR U14513 ( .A(n1345), .B(n1344), .Z(\A1[407] ) );
  XOR U14514 ( .A(n13233), .B(n13234), .Z(n1344) );
  XNOR U14515 ( .A(n13232), .B(n13230), .Z(n13234) );
  AND U14516 ( .A(n13235), .B(n13236), .Z(n13230) );
  NANDN U14517 ( .A(n13237), .B(n13238), .Z(n13236) );
  NANDN U14518 ( .A(n13239), .B(n13240), .Z(n13238) );
  AND U14519 ( .A(B[406]), .B(A[3]), .Z(n13232) );
  XNOR U14520 ( .A(n13222), .B(n13241), .Z(n13233) );
  XNOR U14521 ( .A(n13220), .B(n13223), .Z(n13241) );
  NAND U14522 ( .A(A[2]), .B(B[407]), .Z(n13223) );
  NANDN U14523 ( .A(n13242), .B(n13243), .Z(n13220) );
  AND U14524 ( .A(A[0]), .B(B[408]), .Z(n13243) );
  XOR U14525 ( .A(n13225), .B(n13244), .Z(n13222) );
  NAND U14526 ( .A(A[0]), .B(B[409]), .Z(n13244) );
  NAND U14527 ( .A(B[408]), .B(A[1]), .Z(n13225) );
  NAND U14528 ( .A(n13245), .B(n13246), .Z(n1345) );
  NANDN U14529 ( .A(n13247), .B(n13248), .Z(n13246) );
  OR U14530 ( .A(n13249), .B(n13250), .Z(n13248) );
  NAND U14531 ( .A(n13250), .B(n13249), .Z(n13245) );
  XOR U14532 ( .A(n1347), .B(n1346), .Z(\A1[406] ) );
  XOR U14533 ( .A(n13250), .B(n13251), .Z(n1346) );
  XNOR U14534 ( .A(n13249), .B(n13247), .Z(n13251) );
  AND U14535 ( .A(n13252), .B(n13253), .Z(n13247) );
  NANDN U14536 ( .A(n13254), .B(n13255), .Z(n13253) );
  NANDN U14537 ( .A(n13256), .B(n13257), .Z(n13255) );
  AND U14538 ( .A(B[405]), .B(A[3]), .Z(n13249) );
  XNOR U14539 ( .A(n13239), .B(n13258), .Z(n13250) );
  XNOR U14540 ( .A(n13237), .B(n13240), .Z(n13258) );
  NAND U14541 ( .A(A[2]), .B(B[406]), .Z(n13240) );
  NANDN U14542 ( .A(n13259), .B(n13260), .Z(n13237) );
  AND U14543 ( .A(A[0]), .B(B[407]), .Z(n13260) );
  XOR U14544 ( .A(n13242), .B(n13261), .Z(n13239) );
  NAND U14545 ( .A(A[0]), .B(B[408]), .Z(n13261) );
  NAND U14546 ( .A(B[407]), .B(A[1]), .Z(n13242) );
  NAND U14547 ( .A(n13262), .B(n13263), .Z(n1347) );
  NANDN U14548 ( .A(n13264), .B(n13265), .Z(n13263) );
  OR U14549 ( .A(n13266), .B(n13267), .Z(n13265) );
  NAND U14550 ( .A(n13267), .B(n13266), .Z(n13262) );
  XOR U14551 ( .A(n1349), .B(n1348), .Z(\A1[405] ) );
  XOR U14552 ( .A(n13267), .B(n13268), .Z(n1348) );
  XNOR U14553 ( .A(n13266), .B(n13264), .Z(n13268) );
  AND U14554 ( .A(n13269), .B(n13270), .Z(n13264) );
  NANDN U14555 ( .A(n13271), .B(n13272), .Z(n13270) );
  NANDN U14556 ( .A(n13273), .B(n13274), .Z(n13272) );
  AND U14557 ( .A(B[404]), .B(A[3]), .Z(n13266) );
  XNOR U14558 ( .A(n13256), .B(n13275), .Z(n13267) );
  XNOR U14559 ( .A(n13254), .B(n13257), .Z(n13275) );
  NAND U14560 ( .A(A[2]), .B(B[405]), .Z(n13257) );
  NANDN U14561 ( .A(n13276), .B(n13277), .Z(n13254) );
  AND U14562 ( .A(A[0]), .B(B[406]), .Z(n13277) );
  XOR U14563 ( .A(n13259), .B(n13278), .Z(n13256) );
  NAND U14564 ( .A(A[0]), .B(B[407]), .Z(n13278) );
  NAND U14565 ( .A(B[406]), .B(A[1]), .Z(n13259) );
  NAND U14566 ( .A(n13279), .B(n13280), .Z(n1349) );
  NANDN U14567 ( .A(n13281), .B(n13282), .Z(n13280) );
  OR U14568 ( .A(n13283), .B(n13284), .Z(n13282) );
  NAND U14569 ( .A(n13284), .B(n13283), .Z(n13279) );
  XOR U14570 ( .A(n1351), .B(n1350), .Z(\A1[404] ) );
  XOR U14571 ( .A(n13284), .B(n13285), .Z(n1350) );
  XNOR U14572 ( .A(n13283), .B(n13281), .Z(n13285) );
  AND U14573 ( .A(n13286), .B(n13287), .Z(n13281) );
  NANDN U14574 ( .A(n13288), .B(n13289), .Z(n13287) );
  NANDN U14575 ( .A(n13290), .B(n13291), .Z(n13289) );
  AND U14576 ( .A(B[403]), .B(A[3]), .Z(n13283) );
  XNOR U14577 ( .A(n13273), .B(n13292), .Z(n13284) );
  XNOR U14578 ( .A(n13271), .B(n13274), .Z(n13292) );
  NAND U14579 ( .A(A[2]), .B(B[404]), .Z(n13274) );
  NANDN U14580 ( .A(n13293), .B(n13294), .Z(n13271) );
  AND U14581 ( .A(A[0]), .B(B[405]), .Z(n13294) );
  XOR U14582 ( .A(n13276), .B(n13295), .Z(n13273) );
  NAND U14583 ( .A(A[0]), .B(B[406]), .Z(n13295) );
  NAND U14584 ( .A(B[405]), .B(A[1]), .Z(n13276) );
  NAND U14585 ( .A(n13296), .B(n13297), .Z(n1351) );
  NANDN U14586 ( .A(n13298), .B(n13299), .Z(n13297) );
  OR U14587 ( .A(n13300), .B(n13301), .Z(n13299) );
  NAND U14588 ( .A(n13301), .B(n13300), .Z(n13296) );
  XOR U14589 ( .A(n1353), .B(n1352), .Z(\A1[403] ) );
  XOR U14590 ( .A(n13301), .B(n13302), .Z(n1352) );
  XNOR U14591 ( .A(n13300), .B(n13298), .Z(n13302) );
  AND U14592 ( .A(n13303), .B(n13304), .Z(n13298) );
  NANDN U14593 ( .A(n13305), .B(n13306), .Z(n13304) );
  NANDN U14594 ( .A(n13307), .B(n13308), .Z(n13306) );
  AND U14595 ( .A(B[402]), .B(A[3]), .Z(n13300) );
  XNOR U14596 ( .A(n13290), .B(n13309), .Z(n13301) );
  XNOR U14597 ( .A(n13288), .B(n13291), .Z(n13309) );
  NAND U14598 ( .A(A[2]), .B(B[403]), .Z(n13291) );
  NANDN U14599 ( .A(n13310), .B(n13311), .Z(n13288) );
  AND U14600 ( .A(A[0]), .B(B[404]), .Z(n13311) );
  XOR U14601 ( .A(n13293), .B(n13312), .Z(n13290) );
  NAND U14602 ( .A(A[0]), .B(B[405]), .Z(n13312) );
  NAND U14603 ( .A(B[404]), .B(A[1]), .Z(n13293) );
  NAND U14604 ( .A(n13313), .B(n13314), .Z(n1353) );
  NANDN U14605 ( .A(n13315), .B(n13316), .Z(n13314) );
  OR U14606 ( .A(n13317), .B(n13318), .Z(n13316) );
  NAND U14607 ( .A(n13318), .B(n13317), .Z(n13313) );
  XOR U14608 ( .A(n1355), .B(n1354), .Z(\A1[402] ) );
  XOR U14609 ( .A(n13318), .B(n13319), .Z(n1354) );
  XNOR U14610 ( .A(n13317), .B(n13315), .Z(n13319) );
  AND U14611 ( .A(n13320), .B(n13321), .Z(n13315) );
  NANDN U14612 ( .A(n13322), .B(n13323), .Z(n13321) );
  NANDN U14613 ( .A(n13324), .B(n13325), .Z(n13323) );
  AND U14614 ( .A(B[401]), .B(A[3]), .Z(n13317) );
  XNOR U14615 ( .A(n13307), .B(n13326), .Z(n13318) );
  XNOR U14616 ( .A(n13305), .B(n13308), .Z(n13326) );
  NAND U14617 ( .A(A[2]), .B(B[402]), .Z(n13308) );
  NANDN U14618 ( .A(n13327), .B(n13328), .Z(n13305) );
  AND U14619 ( .A(A[0]), .B(B[403]), .Z(n13328) );
  XOR U14620 ( .A(n13310), .B(n13329), .Z(n13307) );
  NAND U14621 ( .A(A[0]), .B(B[404]), .Z(n13329) );
  NAND U14622 ( .A(B[403]), .B(A[1]), .Z(n13310) );
  NAND U14623 ( .A(n13330), .B(n13331), .Z(n1355) );
  NANDN U14624 ( .A(n13332), .B(n13333), .Z(n13331) );
  OR U14625 ( .A(n13334), .B(n13335), .Z(n13333) );
  NAND U14626 ( .A(n13335), .B(n13334), .Z(n13330) );
  XOR U14627 ( .A(n1357), .B(n1356), .Z(\A1[401] ) );
  XOR U14628 ( .A(n13335), .B(n13336), .Z(n1356) );
  XNOR U14629 ( .A(n13334), .B(n13332), .Z(n13336) );
  AND U14630 ( .A(n13337), .B(n13338), .Z(n13332) );
  NANDN U14631 ( .A(n13339), .B(n13340), .Z(n13338) );
  NANDN U14632 ( .A(n13341), .B(n13342), .Z(n13340) );
  AND U14633 ( .A(B[400]), .B(A[3]), .Z(n13334) );
  XNOR U14634 ( .A(n13324), .B(n13343), .Z(n13335) );
  XNOR U14635 ( .A(n13322), .B(n13325), .Z(n13343) );
  NAND U14636 ( .A(A[2]), .B(B[401]), .Z(n13325) );
  NANDN U14637 ( .A(n13344), .B(n13345), .Z(n13322) );
  AND U14638 ( .A(A[0]), .B(B[402]), .Z(n13345) );
  XOR U14639 ( .A(n13327), .B(n13346), .Z(n13324) );
  NAND U14640 ( .A(A[0]), .B(B[403]), .Z(n13346) );
  NAND U14641 ( .A(B[402]), .B(A[1]), .Z(n13327) );
  NAND U14642 ( .A(n13347), .B(n13348), .Z(n1357) );
  NANDN U14643 ( .A(n13349), .B(n13350), .Z(n13348) );
  OR U14644 ( .A(n13351), .B(n13352), .Z(n13350) );
  NAND U14645 ( .A(n13352), .B(n13351), .Z(n13347) );
  XOR U14646 ( .A(n1359), .B(n1358), .Z(\A1[400] ) );
  XOR U14647 ( .A(n13352), .B(n13353), .Z(n1358) );
  XNOR U14648 ( .A(n13351), .B(n13349), .Z(n13353) );
  AND U14649 ( .A(n13354), .B(n13355), .Z(n13349) );
  NANDN U14650 ( .A(n13356), .B(n13357), .Z(n13355) );
  NANDN U14651 ( .A(n13358), .B(n13359), .Z(n13357) );
  AND U14652 ( .A(B[399]), .B(A[3]), .Z(n13351) );
  XNOR U14653 ( .A(n13341), .B(n13360), .Z(n13352) );
  XNOR U14654 ( .A(n13339), .B(n13342), .Z(n13360) );
  NAND U14655 ( .A(A[2]), .B(B[400]), .Z(n13342) );
  NANDN U14656 ( .A(n13361), .B(n13362), .Z(n13339) );
  AND U14657 ( .A(A[0]), .B(B[401]), .Z(n13362) );
  XOR U14658 ( .A(n13344), .B(n13363), .Z(n13341) );
  NAND U14659 ( .A(A[0]), .B(B[402]), .Z(n13363) );
  NAND U14660 ( .A(B[401]), .B(A[1]), .Z(n13344) );
  NAND U14661 ( .A(n13364), .B(n13365), .Z(n1359) );
  NANDN U14662 ( .A(n13366), .B(n13367), .Z(n13365) );
  OR U14663 ( .A(n13368), .B(n13369), .Z(n13367) );
  NAND U14664 ( .A(n13369), .B(n13368), .Z(n13364) );
  XOR U14665 ( .A(n1141), .B(n1140), .Z(\A1[3] ) );
  XOR U14666 ( .A(n11499), .B(n13370), .Z(n1140) );
  XNOR U14667 ( .A(n11498), .B(n11496), .Z(n13370) );
  AND U14668 ( .A(n13371), .B(n13372), .Z(n11496) );
  NANDN U14669 ( .A(n13373), .B(n13374), .Z(n13372) );
  NANDN U14670 ( .A(n13375), .B(n13376), .Z(n13374) );
  AND U14671 ( .A(B[2]), .B(A[3]), .Z(n11498) );
  XNOR U14672 ( .A(n11488), .B(n13377), .Z(n11499) );
  XNOR U14673 ( .A(n11486), .B(n11489), .Z(n13377) );
  NAND U14674 ( .A(A[2]), .B(B[3]), .Z(n11489) );
  NANDN U14675 ( .A(n13378), .B(n13379), .Z(n11486) );
  AND U14676 ( .A(A[0]), .B(B[4]), .Z(n13379) );
  XOR U14677 ( .A(n11491), .B(n13380), .Z(n11488) );
  NAND U14678 ( .A(A[0]), .B(B[5]), .Z(n13380) );
  NAND U14679 ( .A(B[4]), .B(A[1]), .Z(n11491) );
  NAND U14680 ( .A(n13381), .B(n13382), .Z(n1141) );
  NANDN U14681 ( .A(n13383), .B(n13384), .Z(n13382) );
  OR U14682 ( .A(n13385), .B(n13386), .Z(n13384) );
  NAND U14683 ( .A(n13386), .B(n13385), .Z(n13381) );
  XOR U14684 ( .A(n1341), .B(n1340), .Z(\A1[39] ) );
  XOR U14685 ( .A(n13199), .B(n13387), .Z(n1340) );
  XNOR U14686 ( .A(n13198), .B(n13196), .Z(n13387) );
  AND U14687 ( .A(n13388), .B(n13389), .Z(n13196) );
  NANDN U14688 ( .A(n13390), .B(n13391), .Z(n13389) );
  NANDN U14689 ( .A(n13392), .B(n13393), .Z(n13391) );
  AND U14690 ( .A(B[38]), .B(A[3]), .Z(n13198) );
  XNOR U14691 ( .A(n13188), .B(n13394), .Z(n13199) );
  XNOR U14692 ( .A(n13186), .B(n13189), .Z(n13394) );
  NAND U14693 ( .A(A[2]), .B(B[39]), .Z(n13189) );
  NANDN U14694 ( .A(n13395), .B(n13396), .Z(n13186) );
  AND U14695 ( .A(A[0]), .B(B[40]), .Z(n13396) );
  XOR U14696 ( .A(n13191), .B(n13397), .Z(n13188) );
  NAND U14697 ( .A(A[0]), .B(B[41]), .Z(n13397) );
  NAND U14698 ( .A(B[40]), .B(A[1]), .Z(n13191) );
  NAND U14699 ( .A(n13398), .B(n13399), .Z(n1341) );
  NANDN U14700 ( .A(n13400), .B(n13401), .Z(n13399) );
  OR U14701 ( .A(n13402), .B(n13403), .Z(n13401) );
  NAND U14702 ( .A(n13403), .B(n13402), .Z(n13398) );
  XOR U14703 ( .A(n1361), .B(n1360), .Z(\A1[399] ) );
  XOR U14704 ( .A(n13369), .B(n13404), .Z(n1360) );
  XNOR U14705 ( .A(n13368), .B(n13366), .Z(n13404) );
  AND U14706 ( .A(n13405), .B(n13406), .Z(n13366) );
  NANDN U14707 ( .A(n13407), .B(n13408), .Z(n13406) );
  NANDN U14708 ( .A(n13409), .B(n13410), .Z(n13408) );
  AND U14709 ( .A(B[398]), .B(A[3]), .Z(n13368) );
  XNOR U14710 ( .A(n13358), .B(n13411), .Z(n13369) );
  XNOR U14711 ( .A(n13356), .B(n13359), .Z(n13411) );
  NAND U14712 ( .A(A[2]), .B(B[399]), .Z(n13359) );
  NANDN U14713 ( .A(n13412), .B(n13413), .Z(n13356) );
  AND U14714 ( .A(A[0]), .B(B[400]), .Z(n13413) );
  XOR U14715 ( .A(n13361), .B(n13414), .Z(n13358) );
  NAND U14716 ( .A(A[0]), .B(B[401]), .Z(n13414) );
  NAND U14717 ( .A(B[400]), .B(A[1]), .Z(n13361) );
  NAND U14718 ( .A(n13415), .B(n13416), .Z(n1361) );
  NANDN U14719 ( .A(n13417), .B(n13418), .Z(n13416) );
  OR U14720 ( .A(n13419), .B(n13420), .Z(n13418) );
  NAND U14721 ( .A(n13420), .B(n13419), .Z(n13415) );
  XOR U14722 ( .A(n1367), .B(n1366), .Z(\A1[398] ) );
  XOR U14723 ( .A(n13420), .B(n13421), .Z(n1366) );
  XNOR U14724 ( .A(n13419), .B(n13417), .Z(n13421) );
  AND U14725 ( .A(n13422), .B(n13423), .Z(n13417) );
  NANDN U14726 ( .A(n13424), .B(n13425), .Z(n13423) );
  NANDN U14727 ( .A(n13426), .B(n13427), .Z(n13425) );
  AND U14728 ( .A(B[397]), .B(A[3]), .Z(n13419) );
  XNOR U14729 ( .A(n13409), .B(n13428), .Z(n13420) );
  XNOR U14730 ( .A(n13407), .B(n13410), .Z(n13428) );
  NAND U14731 ( .A(A[2]), .B(B[398]), .Z(n13410) );
  NANDN U14732 ( .A(n13429), .B(n13430), .Z(n13407) );
  AND U14733 ( .A(A[0]), .B(B[399]), .Z(n13430) );
  XOR U14734 ( .A(n13412), .B(n13431), .Z(n13409) );
  NAND U14735 ( .A(A[0]), .B(B[400]), .Z(n13431) );
  NAND U14736 ( .A(B[399]), .B(A[1]), .Z(n13412) );
  NAND U14737 ( .A(n13432), .B(n13433), .Z(n1367) );
  NANDN U14738 ( .A(n13434), .B(n13435), .Z(n13433) );
  OR U14739 ( .A(n13436), .B(n13437), .Z(n13435) );
  NAND U14740 ( .A(n13437), .B(n13436), .Z(n13432) );
  XOR U14741 ( .A(n1369), .B(n1368), .Z(\A1[397] ) );
  XOR U14742 ( .A(n13437), .B(n13438), .Z(n1368) );
  XNOR U14743 ( .A(n13436), .B(n13434), .Z(n13438) );
  AND U14744 ( .A(n13439), .B(n13440), .Z(n13434) );
  NANDN U14745 ( .A(n13441), .B(n13442), .Z(n13440) );
  NANDN U14746 ( .A(n13443), .B(n13444), .Z(n13442) );
  AND U14747 ( .A(B[396]), .B(A[3]), .Z(n13436) );
  XNOR U14748 ( .A(n13426), .B(n13445), .Z(n13437) );
  XNOR U14749 ( .A(n13424), .B(n13427), .Z(n13445) );
  NAND U14750 ( .A(A[2]), .B(B[397]), .Z(n13427) );
  NANDN U14751 ( .A(n13446), .B(n13447), .Z(n13424) );
  AND U14752 ( .A(A[0]), .B(B[398]), .Z(n13447) );
  XOR U14753 ( .A(n13429), .B(n13448), .Z(n13426) );
  NAND U14754 ( .A(A[0]), .B(B[399]), .Z(n13448) );
  NAND U14755 ( .A(B[398]), .B(A[1]), .Z(n13429) );
  NAND U14756 ( .A(n13449), .B(n13450), .Z(n1369) );
  NANDN U14757 ( .A(n13451), .B(n13452), .Z(n13450) );
  OR U14758 ( .A(n13453), .B(n13454), .Z(n13452) );
  NAND U14759 ( .A(n13454), .B(n13453), .Z(n13449) );
  XOR U14760 ( .A(n1371), .B(n1370), .Z(\A1[396] ) );
  XOR U14761 ( .A(n13454), .B(n13455), .Z(n1370) );
  XNOR U14762 ( .A(n13453), .B(n13451), .Z(n13455) );
  AND U14763 ( .A(n13456), .B(n13457), .Z(n13451) );
  NANDN U14764 ( .A(n13458), .B(n13459), .Z(n13457) );
  NANDN U14765 ( .A(n13460), .B(n13461), .Z(n13459) );
  AND U14766 ( .A(B[395]), .B(A[3]), .Z(n13453) );
  XNOR U14767 ( .A(n13443), .B(n13462), .Z(n13454) );
  XNOR U14768 ( .A(n13441), .B(n13444), .Z(n13462) );
  NAND U14769 ( .A(A[2]), .B(B[396]), .Z(n13444) );
  NANDN U14770 ( .A(n13463), .B(n13464), .Z(n13441) );
  AND U14771 ( .A(A[0]), .B(B[397]), .Z(n13464) );
  XOR U14772 ( .A(n13446), .B(n13465), .Z(n13443) );
  NAND U14773 ( .A(A[0]), .B(B[398]), .Z(n13465) );
  NAND U14774 ( .A(B[397]), .B(A[1]), .Z(n13446) );
  NAND U14775 ( .A(n13466), .B(n13467), .Z(n1371) );
  NANDN U14776 ( .A(n13468), .B(n13469), .Z(n13467) );
  OR U14777 ( .A(n13470), .B(n13471), .Z(n13469) );
  NAND U14778 ( .A(n13471), .B(n13470), .Z(n13466) );
  XOR U14779 ( .A(n1373), .B(n1372), .Z(\A1[395] ) );
  XOR U14780 ( .A(n13471), .B(n13472), .Z(n1372) );
  XNOR U14781 ( .A(n13470), .B(n13468), .Z(n13472) );
  AND U14782 ( .A(n13473), .B(n13474), .Z(n13468) );
  NANDN U14783 ( .A(n13475), .B(n13476), .Z(n13474) );
  NANDN U14784 ( .A(n13477), .B(n13478), .Z(n13476) );
  AND U14785 ( .A(B[394]), .B(A[3]), .Z(n13470) );
  XNOR U14786 ( .A(n13460), .B(n13479), .Z(n13471) );
  XNOR U14787 ( .A(n13458), .B(n13461), .Z(n13479) );
  NAND U14788 ( .A(A[2]), .B(B[395]), .Z(n13461) );
  NANDN U14789 ( .A(n13480), .B(n13481), .Z(n13458) );
  AND U14790 ( .A(A[0]), .B(B[396]), .Z(n13481) );
  XOR U14791 ( .A(n13463), .B(n13482), .Z(n13460) );
  NAND U14792 ( .A(A[0]), .B(B[397]), .Z(n13482) );
  NAND U14793 ( .A(B[396]), .B(A[1]), .Z(n13463) );
  NAND U14794 ( .A(n13483), .B(n13484), .Z(n1373) );
  NANDN U14795 ( .A(n13485), .B(n13486), .Z(n13484) );
  OR U14796 ( .A(n13487), .B(n13488), .Z(n13486) );
  NAND U14797 ( .A(n13488), .B(n13487), .Z(n13483) );
  XOR U14798 ( .A(n1375), .B(n1374), .Z(\A1[394] ) );
  XOR U14799 ( .A(n13488), .B(n13489), .Z(n1374) );
  XNOR U14800 ( .A(n13487), .B(n13485), .Z(n13489) );
  AND U14801 ( .A(n13490), .B(n13491), .Z(n13485) );
  NANDN U14802 ( .A(n13492), .B(n13493), .Z(n13491) );
  NANDN U14803 ( .A(n13494), .B(n13495), .Z(n13493) );
  AND U14804 ( .A(B[393]), .B(A[3]), .Z(n13487) );
  XNOR U14805 ( .A(n13477), .B(n13496), .Z(n13488) );
  XNOR U14806 ( .A(n13475), .B(n13478), .Z(n13496) );
  NAND U14807 ( .A(A[2]), .B(B[394]), .Z(n13478) );
  NANDN U14808 ( .A(n13497), .B(n13498), .Z(n13475) );
  AND U14809 ( .A(A[0]), .B(B[395]), .Z(n13498) );
  XOR U14810 ( .A(n13480), .B(n13499), .Z(n13477) );
  NAND U14811 ( .A(A[0]), .B(B[396]), .Z(n13499) );
  NAND U14812 ( .A(B[395]), .B(A[1]), .Z(n13480) );
  NAND U14813 ( .A(n13500), .B(n13501), .Z(n1375) );
  NANDN U14814 ( .A(n13502), .B(n13503), .Z(n13501) );
  OR U14815 ( .A(n13504), .B(n13505), .Z(n13503) );
  NAND U14816 ( .A(n13505), .B(n13504), .Z(n13500) );
  XOR U14817 ( .A(n1377), .B(n1376), .Z(\A1[393] ) );
  XOR U14818 ( .A(n13505), .B(n13506), .Z(n1376) );
  XNOR U14819 ( .A(n13504), .B(n13502), .Z(n13506) );
  AND U14820 ( .A(n13507), .B(n13508), .Z(n13502) );
  NANDN U14821 ( .A(n13509), .B(n13510), .Z(n13508) );
  NANDN U14822 ( .A(n13511), .B(n13512), .Z(n13510) );
  AND U14823 ( .A(B[392]), .B(A[3]), .Z(n13504) );
  XNOR U14824 ( .A(n13494), .B(n13513), .Z(n13505) );
  XNOR U14825 ( .A(n13492), .B(n13495), .Z(n13513) );
  NAND U14826 ( .A(A[2]), .B(B[393]), .Z(n13495) );
  NANDN U14827 ( .A(n13514), .B(n13515), .Z(n13492) );
  AND U14828 ( .A(A[0]), .B(B[394]), .Z(n13515) );
  XOR U14829 ( .A(n13497), .B(n13516), .Z(n13494) );
  NAND U14830 ( .A(A[0]), .B(B[395]), .Z(n13516) );
  NAND U14831 ( .A(B[394]), .B(A[1]), .Z(n13497) );
  NAND U14832 ( .A(n13517), .B(n13518), .Z(n1377) );
  NANDN U14833 ( .A(n13519), .B(n13520), .Z(n13518) );
  OR U14834 ( .A(n13521), .B(n13522), .Z(n13520) );
  NAND U14835 ( .A(n13522), .B(n13521), .Z(n13517) );
  XOR U14836 ( .A(n1379), .B(n1378), .Z(\A1[392] ) );
  XOR U14837 ( .A(n13522), .B(n13523), .Z(n1378) );
  XNOR U14838 ( .A(n13521), .B(n13519), .Z(n13523) );
  AND U14839 ( .A(n13524), .B(n13525), .Z(n13519) );
  NANDN U14840 ( .A(n13526), .B(n13527), .Z(n13525) );
  NANDN U14841 ( .A(n13528), .B(n13529), .Z(n13527) );
  AND U14842 ( .A(B[391]), .B(A[3]), .Z(n13521) );
  XNOR U14843 ( .A(n13511), .B(n13530), .Z(n13522) );
  XNOR U14844 ( .A(n13509), .B(n13512), .Z(n13530) );
  NAND U14845 ( .A(A[2]), .B(B[392]), .Z(n13512) );
  NANDN U14846 ( .A(n13531), .B(n13532), .Z(n13509) );
  AND U14847 ( .A(A[0]), .B(B[393]), .Z(n13532) );
  XOR U14848 ( .A(n13514), .B(n13533), .Z(n13511) );
  NAND U14849 ( .A(A[0]), .B(B[394]), .Z(n13533) );
  NAND U14850 ( .A(B[393]), .B(A[1]), .Z(n13514) );
  NAND U14851 ( .A(n13534), .B(n13535), .Z(n1379) );
  NANDN U14852 ( .A(n13536), .B(n13537), .Z(n13535) );
  OR U14853 ( .A(n13538), .B(n13539), .Z(n13537) );
  NAND U14854 ( .A(n13539), .B(n13538), .Z(n13534) );
  XOR U14855 ( .A(n1381), .B(n1380), .Z(\A1[391] ) );
  XOR U14856 ( .A(n13539), .B(n13540), .Z(n1380) );
  XNOR U14857 ( .A(n13538), .B(n13536), .Z(n13540) );
  AND U14858 ( .A(n13541), .B(n13542), .Z(n13536) );
  NANDN U14859 ( .A(n13543), .B(n13544), .Z(n13542) );
  NANDN U14860 ( .A(n13545), .B(n13546), .Z(n13544) );
  AND U14861 ( .A(B[390]), .B(A[3]), .Z(n13538) );
  XNOR U14862 ( .A(n13528), .B(n13547), .Z(n13539) );
  XNOR U14863 ( .A(n13526), .B(n13529), .Z(n13547) );
  NAND U14864 ( .A(A[2]), .B(B[391]), .Z(n13529) );
  NANDN U14865 ( .A(n13548), .B(n13549), .Z(n13526) );
  AND U14866 ( .A(A[0]), .B(B[392]), .Z(n13549) );
  XOR U14867 ( .A(n13531), .B(n13550), .Z(n13528) );
  NAND U14868 ( .A(A[0]), .B(B[393]), .Z(n13550) );
  NAND U14869 ( .A(B[392]), .B(A[1]), .Z(n13531) );
  NAND U14870 ( .A(n13551), .B(n13552), .Z(n1381) );
  NANDN U14871 ( .A(n13553), .B(n13554), .Z(n13552) );
  OR U14872 ( .A(n13555), .B(n13556), .Z(n13554) );
  NAND U14873 ( .A(n13556), .B(n13555), .Z(n13551) );
  XOR U14874 ( .A(n1383), .B(n1382), .Z(\A1[390] ) );
  XOR U14875 ( .A(n13556), .B(n13557), .Z(n1382) );
  XNOR U14876 ( .A(n13555), .B(n13553), .Z(n13557) );
  AND U14877 ( .A(n13558), .B(n13559), .Z(n13553) );
  NANDN U14878 ( .A(n13560), .B(n13561), .Z(n13559) );
  NANDN U14879 ( .A(n13562), .B(n13563), .Z(n13561) );
  AND U14880 ( .A(B[389]), .B(A[3]), .Z(n13555) );
  XNOR U14881 ( .A(n13545), .B(n13564), .Z(n13556) );
  XNOR U14882 ( .A(n13543), .B(n13546), .Z(n13564) );
  NAND U14883 ( .A(A[2]), .B(B[390]), .Z(n13546) );
  NANDN U14884 ( .A(n13565), .B(n13566), .Z(n13543) );
  AND U14885 ( .A(A[0]), .B(B[391]), .Z(n13566) );
  XOR U14886 ( .A(n13548), .B(n13567), .Z(n13545) );
  NAND U14887 ( .A(A[0]), .B(B[392]), .Z(n13567) );
  NAND U14888 ( .A(B[391]), .B(A[1]), .Z(n13548) );
  NAND U14889 ( .A(n13568), .B(n13569), .Z(n1383) );
  NANDN U14890 ( .A(n13570), .B(n13571), .Z(n13569) );
  OR U14891 ( .A(n13572), .B(n13573), .Z(n13571) );
  NAND U14892 ( .A(n13573), .B(n13572), .Z(n13568) );
  XOR U14893 ( .A(n1365), .B(n1364), .Z(\A1[38] ) );
  XOR U14894 ( .A(n13403), .B(n13574), .Z(n1364) );
  XNOR U14895 ( .A(n13402), .B(n13400), .Z(n13574) );
  AND U14896 ( .A(n13575), .B(n13576), .Z(n13400) );
  NANDN U14897 ( .A(n13577), .B(n13578), .Z(n13576) );
  NANDN U14898 ( .A(n13579), .B(n13580), .Z(n13578) );
  AND U14899 ( .A(B[37]), .B(A[3]), .Z(n13402) );
  XNOR U14900 ( .A(n13392), .B(n13581), .Z(n13403) );
  XNOR U14901 ( .A(n13390), .B(n13393), .Z(n13581) );
  NAND U14902 ( .A(A[2]), .B(B[38]), .Z(n13393) );
  NANDN U14903 ( .A(n13582), .B(n13583), .Z(n13390) );
  AND U14904 ( .A(A[0]), .B(B[39]), .Z(n13583) );
  XOR U14905 ( .A(n13395), .B(n13584), .Z(n13392) );
  NAND U14906 ( .A(A[0]), .B(B[40]), .Z(n13584) );
  NAND U14907 ( .A(B[39]), .B(A[1]), .Z(n13395) );
  NAND U14908 ( .A(n13585), .B(n13586), .Z(n1365) );
  NANDN U14909 ( .A(n13587), .B(n13588), .Z(n13586) );
  OR U14910 ( .A(n13589), .B(n13590), .Z(n13588) );
  NAND U14911 ( .A(n13590), .B(n13589), .Z(n13585) );
  XOR U14912 ( .A(n1385), .B(n1384), .Z(\A1[389] ) );
  XOR U14913 ( .A(n13573), .B(n13591), .Z(n1384) );
  XNOR U14914 ( .A(n13572), .B(n13570), .Z(n13591) );
  AND U14915 ( .A(n13592), .B(n13593), .Z(n13570) );
  NANDN U14916 ( .A(n13594), .B(n13595), .Z(n13593) );
  NANDN U14917 ( .A(n13596), .B(n13597), .Z(n13595) );
  AND U14918 ( .A(B[388]), .B(A[3]), .Z(n13572) );
  XNOR U14919 ( .A(n13562), .B(n13598), .Z(n13573) );
  XNOR U14920 ( .A(n13560), .B(n13563), .Z(n13598) );
  NAND U14921 ( .A(A[2]), .B(B[389]), .Z(n13563) );
  NANDN U14922 ( .A(n13599), .B(n13600), .Z(n13560) );
  AND U14923 ( .A(A[0]), .B(B[390]), .Z(n13600) );
  XOR U14924 ( .A(n13565), .B(n13601), .Z(n13562) );
  NAND U14925 ( .A(A[0]), .B(B[391]), .Z(n13601) );
  NAND U14926 ( .A(B[390]), .B(A[1]), .Z(n13565) );
  NAND U14927 ( .A(n13602), .B(n13603), .Z(n1385) );
  NANDN U14928 ( .A(n13604), .B(n13605), .Z(n13603) );
  OR U14929 ( .A(n13606), .B(n13607), .Z(n13605) );
  NAND U14930 ( .A(n13607), .B(n13606), .Z(n13602) );
  XOR U14931 ( .A(n1389), .B(n1388), .Z(\A1[388] ) );
  XOR U14932 ( .A(n13607), .B(n13608), .Z(n1388) );
  XNOR U14933 ( .A(n13606), .B(n13604), .Z(n13608) );
  AND U14934 ( .A(n13609), .B(n13610), .Z(n13604) );
  NANDN U14935 ( .A(n13611), .B(n13612), .Z(n13610) );
  NANDN U14936 ( .A(n13613), .B(n13614), .Z(n13612) );
  AND U14937 ( .A(B[387]), .B(A[3]), .Z(n13606) );
  XNOR U14938 ( .A(n13596), .B(n13615), .Z(n13607) );
  XNOR U14939 ( .A(n13594), .B(n13597), .Z(n13615) );
  NAND U14940 ( .A(A[2]), .B(B[388]), .Z(n13597) );
  NANDN U14941 ( .A(n13616), .B(n13617), .Z(n13594) );
  AND U14942 ( .A(A[0]), .B(B[389]), .Z(n13617) );
  XOR U14943 ( .A(n13599), .B(n13618), .Z(n13596) );
  NAND U14944 ( .A(A[0]), .B(B[390]), .Z(n13618) );
  NAND U14945 ( .A(B[389]), .B(A[1]), .Z(n13599) );
  NAND U14946 ( .A(n13619), .B(n13620), .Z(n1389) );
  NANDN U14947 ( .A(n13621), .B(n13622), .Z(n13620) );
  OR U14948 ( .A(n13623), .B(n13624), .Z(n13622) );
  NAND U14949 ( .A(n13624), .B(n13623), .Z(n13619) );
  XOR U14950 ( .A(n1391), .B(n1390), .Z(\A1[387] ) );
  XOR U14951 ( .A(n13624), .B(n13625), .Z(n1390) );
  XNOR U14952 ( .A(n13623), .B(n13621), .Z(n13625) );
  AND U14953 ( .A(n13626), .B(n13627), .Z(n13621) );
  NANDN U14954 ( .A(n13628), .B(n13629), .Z(n13627) );
  NANDN U14955 ( .A(n13630), .B(n13631), .Z(n13629) );
  AND U14956 ( .A(B[386]), .B(A[3]), .Z(n13623) );
  XNOR U14957 ( .A(n13613), .B(n13632), .Z(n13624) );
  XNOR U14958 ( .A(n13611), .B(n13614), .Z(n13632) );
  NAND U14959 ( .A(A[2]), .B(B[387]), .Z(n13614) );
  NANDN U14960 ( .A(n13633), .B(n13634), .Z(n13611) );
  AND U14961 ( .A(A[0]), .B(B[388]), .Z(n13634) );
  XOR U14962 ( .A(n13616), .B(n13635), .Z(n13613) );
  NAND U14963 ( .A(A[0]), .B(B[389]), .Z(n13635) );
  NAND U14964 ( .A(B[388]), .B(A[1]), .Z(n13616) );
  NAND U14965 ( .A(n13636), .B(n13637), .Z(n1391) );
  NANDN U14966 ( .A(n13638), .B(n13639), .Z(n13637) );
  OR U14967 ( .A(n13640), .B(n13641), .Z(n13639) );
  NAND U14968 ( .A(n13641), .B(n13640), .Z(n13636) );
  XOR U14969 ( .A(n1393), .B(n1392), .Z(\A1[386] ) );
  XOR U14970 ( .A(n13641), .B(n13642), .Z(n1392) );
  XNOR U14971 ( .A(n13640), .B(n13638), .Z(n13642) );
  AND U14972 ( .A(n13643), .B(n13644), .Z(n13638) );
  NANDN U14973 ( .A(n13645), .B(n13646), .Z(n13644) );
  NANDN U14974 ( .A(n13647), .B(n13648), .Z(n13646) );
  AND U14975 ( .A(B[385]), .B(A[3]), .Z(n13640) );
  XNOR U14976 ( .A(n13630), .B(n13649), .Z(n13641) );
  XNOR U14977 ( .A(n13628), .B(n13631), .Z(n13649) );
  NAND U14978 ( .A(A[2]), .B(B[386]), .Z(n13631) );
  NANDN U14979 ( .A(n13650), .B(n13651), .Z(n13628) );
  AND U14980 ( .A(A[0]), .B(B[387]), .Z(n13651) );
  XOR U14981 ( .A(n13633), .B(n13652), .Z(n13630) );
  NAND U14982 ( .A(A[0]), .B(B[388]), .Z(n13652) );
  NAND U14983 ( .A(B[387]), .B(A[1]), .Z(n13633) );
  NAND U14984 ( .A(n13653), .B(n13654), .Z(n1393) );
  NANDN U14985 ( .A(n13655), .B(n13656), .Z(n13654) );
  OR U14986 ( .A(n13657), .B(n13658), .Z(n13656) );
  NAND U14987 ( .A(n13658), .B(n13657), .Z(n13653) );
  XOR U14988 ( .A(n1395), .B(n1394), .Z(\A1[385] ) );
  XOR U14989 ( .A(n13658), .B(n13659), .Z(n1394) );
  XNOR U14990 ( .A(n13657), .B(n13655), .Z(n13659) );
  AND U14991 ( .A(n13660), .B(n13661), .Z(n13655) );
  NANDN U14992 ( .A(n13662), .B(n13663), .Z(n13661) );
  NANDN U14993 ( .A(n13664), .B(n13665), .Z(n13663) );
  AND U14994 ( .A(B[384]), .B(A[3]), .Z(n13657) );
  XNOR U14995 ( .A(n13647), .B(n13666), .Z(n13658) );
  XNOR U14996 ( .A(n13645), .B(n13648), .Z(n13666) );
  NAND U14997 ( .A(A[2]), .B(B[385]), .Z(n13648) );
  NANDN U14998 ( .A(n13667), .B(n13668), .Z(n13645) );
  AND U14999 ( .A(A[0]), .B(B[386]), .Z(n13668) );
  XOR U15000 ( .A(n13650), .B(n13669), .Z(n13647) );
  NAND U15001 ( .A(A[0]), .B(B[387]), .Z(n13669) );
  NAND U15002 ( .A(B[386]), .B(A[1]), .Z(n13650) );
  NAND U15003 ( .A(n13670), .B(n13671), .Z(n1395) );
  NANDN U15004 ( .A(n13672), .B(n13673), .Z(n13671) );
  OR U15005 ( .A(n13674), .B(n13675), .Z(n13673) );
  NAND U15006 ( .A(n13675), .B(n13674), .Z(n13670) );
  XOR U15007 ( .A(n1397), .B(n1396), .Z(\A1[384] ) );
  XOR U15008 ( .A(n13675), .B(n13676), .Z(n1396) );
  XNOR U15009 ( .A(n13674), .B(n13672), .Z(n13676) );
  AND U15010 ( .A(n13677), .B(n13678), .Z(n13672) );
  NANDN U15011 ( .A(n13679), .B(n13680), .Z(n13678) );
  NANDN U15012 ( .A(n13681), .B(n13682), .Z(n13680) );
  AND U15013 ( .A(B[383]), .B(A[3]), .Z(n13674) );
  XNOR U15014 ( .A(n13664), .B(n13683), .Z(n13675) );
  XNOR U15015 ( .A(n13662), .B(n13665), .Z(n13683) );
  NAND U15016 ( .A(A[2]), .B(B[384]), .Z(n13665) );
  NANDN U15017 ( .A(n13684), .B(n13685), .Z(n13662) );
  AND U15018 ( .A(A[0]), .B(B[385]), .Z(n13685) );
  XOR U15019 ( .A(n13667), .B(n13686), .Z(n13664) );
  NAND U15020 ( .A(A[0]), .B(B[386]), .Z(n13686) );
  NAND U15021 ( .A(B[385]), .B(A[1]), .Z(n13667) );
  NAND U15022 ( .A(n13687), .B(n13688), .Z(n1397) );
  NANDN U15023 ( .A(n13689), .B(n13690), .Z(n13688) );
  OR U15024 ( .A(n13691), .B(n13692), .Z(n13690) );
  NAND U15025 ( .A(n13692), .B(n13691), .Z(n13687) );
  XOR U15026 ( .A(n1399), .B(n1398), .Z(\A1[383] ) );
  XOR U15027 ( .A(n13692), .B(n13693), .Z(n1398) );
  XNOR U15028 ( .A(n13691), .B(n13689), .Z(n13693) );
  AND U15029 ( .A(n13694), .B(n13695), .Z(n13689) );
  NANDN U15030 ( .A(n13696), .B(n13697), .Z(n13695) );
  NANDN U15031 ( .A(n13698), .B(n13699), .Z(n13697) );
  AND U15032 ( .A(B[382]), .B(A[3]), .Z(n13691) );
  XNOR U15033 ( .A(n13681), .B(n13700), .Z(n13692) );
  XNOR U15034 ( .A(n13679), .B(n13682), .Z(n13700) );
  NAND U15035 ( .A(A[2]), .B(B[383]), .Z(n13682) );
  NANDN U15036 ( .A(n13701), .B(n13702), .Z(n13679) );
  AND U15037 ( .A(A[0]), .B(B[384]), .Z(n13702) );
  XOR U15038 ( .A(n13684), .B(n13703), .Z(n13681) );
  NAND U15039 ( .A(A[0]), .B(B[385]), .Z(n13703) );
  NAND U15040 ( .A(B[384]), .B(A[1]), .Z(n13684) );
  NAND U15041 ( .A(n13704), .B(n13705), .Z(n1399) );
  NANDN U15042 ( .A(n13706), .B(n13707), .Z(n13705) );
  OR U15043 ( .A(n13708), .B(n13709), .Z(n13707) );
  NAND U15044 ( .A(n13709), .B(n13708), .Z(n13704) );
  XOR U15045 ( .A(n1401), .B(n1400), .Z(\A1[382] ) );
  XOR U15046 ( .A(n13709), .B(n13710), .Z(n1400) );
  XNOR U15047 ( .A(n13708), .B(n13706), .Z(n13710) );
  AND U15048 ( .A(n13711), .B(n13712), .Z(n13706) );
  NANDN U15049 ( .A(n13713), .B(n13714), .Z(n13712) );
  NANDN U15050 ( .A(n13715), .B(n13716), .Z(n13714) );
  AND U15051 ( .A(B[381]), .B(A[3]), .Z(n13708) );
  XNOR U15052 ( .A(n13698), .B(n13717), .Z(n13709) );
  XNOR U15053 ( .A(n13696), .B(n13699), .Z(n13717) );
  NAND U15054 ( .A(A[2]), .B(B[382]), .Z(n13699) );
  NANDN U15055 ( .A(n13718), .B(n13719), .Z(n13696) );
  AND U15056 ( .A(A[0]), .B(B[383]), .Z(n13719) );
  XOR U15057 ( .A(n13701), .B(n13720), .Z(n13698) );
  NAND U15058 ( .A(A[0]), .B(B[384]), .Z(n13720) );
  NAND U15059 ( .A(B[383]), .B(A[1]), .Z(n13701) );
  NAND U15060 ( .A(n13721), .B(n13722), .Z(n1401) );
  NANDN U15061 ( .A(n13723), .B(n13724), .Z(n13722) );
  OR U15062 ( .A(n13725), .B(n13726), .Z(n13724) );
  NAND U15063 ( .A(n13726), .B(n13725), .Z(n13721) );
  XOR U15064 ( .A(n1403), .B(n1402), .Z(\A1[381] ) );
  XOR U15065 ( .A(n13726), .B(n13727), .Z(n1402) );
  XNOR U15066 ( .A(n13725), .B(n13723), .Z(n13727) );
  AND U15067 ( .A(n13728), .B(n13729), .Z(n13723) );
  NANDN U15068 ( .A(n13730), .B(n13731), .Z(n13729) );
  NANDN U15069 ( .A(n13732), .B(n13733), .Z(n13731) );
  AND U15070 ( .A(B[380]), .B(A[3]), .Z(n13725) );
  XNOR U15071 ( .A(n13715), .B(n13734), .Z(n13726) );
  XNOR U15072 ( .A(n13713), .B(n13716), .Z(n13734) );
  NAND U15073 ( .A(A[2]), .B(B[381]), .Z(n13716) );
  NANDN U15074 ( .A(n13735), .B(n13736), .Z(n13713) );
  AND U15075 ( .A(A[0]), .B(B[382]), .Z(n13736) );
  XOR U15076 ( .A(n13718), .B(n13737), .Z(n13715) );
  NAND U15077 ( .A(A[0]), .B(B[383]), .Z(n13737) );
  NAND U15078 ( .A(B[382]), .B(A[1]), .Z(n13718) );
  NAND U15079 ( .A(n13738), .B(n13739), .Z(n1403) );
  NANDN U15080 ( .A(n13740), .B(n13741), .Z(n13739) );
  OR U15081 ( .A(n13742), .B(n13743), .Z(n13741) );
  NAND U15082 ( .A(n13743), .B(n13742), .Z(n13738) );
  XOR U15083 ( .A(n1405), .B(n1404), .Z(\A1[380] ) );
  XOR U15084 ( .A(n13743), .B(n13744), .Z(n1404) );
  XNOR U15085 ( .A(n13742), .B(n13740), .Z(n13744) );
  AND U15086 ( .A(n13745), .B(n13746), .Z(n13740) );
  NANDN U15087 ( .A(n13747), .B(n13748), .Z(n13746) );
  NANDN U15088 ( .A(n13749), .B(n13750), .Z(n13748) );
  AND U15089 ( .A(B[379]), .B(A[3]), .Z(n13742) );
  XNOR U15090 ( .A(n13732), .B(n13751), .Z(n13743) );
  XNOR U15091 ( .A(n13730), .B(n13733), .Z(n13751) );
  NAND U15092 ( .A(A[2]), .B(B[380]), .Z(n13733) );
  NANDN U15093 ( .A(n13752), .B(n13753), .Z(n13730) );
  AND U15094 ( .A(A[0]), .B(B[381]), .Z(n13753) );
  XOR U15095 ( .A(n13735), .B(n13754), .Z(n13732) );
  NAND U15096 ( .A(A[0]), .B(B[382]), .Z(n13754) );
  NAND U15097 ( .A(B[381]), .B(A[1]), .Z(n13735) );
  NAND U15098 ( .A(n13755), .B(n13756), .Z(n1405) );
  NANDN U15099 ( .A(n13757), .B(n13758), .Z(n13756) );
  OR U15100 ( .A(n13759), .B(n13760), .Z(n13758) );
  NAND U15101 ( .A(n13760), .B(n13759), .Z(n13755) );
  XOR U15102 ( .A(n1387), .B(n1386), .Z(\A1[37] ) );
  XOR U15103 ( .A(n13590), .B(n13761), .Z(n1386) );
  XNOR U15104 ( .A(n13589), .B(n13587), .Z(n13761) );
  AND U15105 ( .A(n13762), .B(n13763), .Z(n13587) );
  NANDN U15106 ( .A(n13764), .B(n13765), .Z(n13763) );
  NANDN U15107 ( .A(n13766), .B(n13767), .Z(n13765) );
  AND U15108 ( .A(B[36]), .B(A[3]), .Z(n13589) );
  XNOR U15109 ( .A(n13579), .B(n13768), .Z(n13590) );
  XNOR U15110 ( .A(n13577), .B(n13580), .Z(n13768) );
  NAND U15111 ( .A(A[2]), .B(B[37]), .Z(n13580) );
  NANDN U15112 ( .A(n13769), .B(n13770), .Z(n13577) );
  AND U15113 ( .A(A[0]), .B(B[38]), .Z(n13770) );
  XOR U15114 ( .A(n13582), .B(n13771), .Z(n13579) );
  NAND U15115 ( .A(A[0]), .B(B[39]), .Z(n13771) );
  NAND U15116 ( .A(B[38]), .B(A[1]), .Z(n13582) );
  NAND U15117 ( .A(n13772), .B(n13773), .Z(n1387) );
  NANDN U15118 ( .A(n13774), .B(n13775), .Z(n13773) );
  OR U15119 ( .A(n13776), .B(n13777), .Z(n13775) );
  NAND U15120 ( .A(n13777), .B(n13776), .Z(n13772) );
  XOR U15121 ( .A(n1407), .B(n1406), .Z(\A1[379] ) );
  XOR U15122 ( .A(n13760), .B(n13778), .Z(n1406) );
  XNOR U15123 ( .A(n13759), .B(n13757), .Z(n13778) );
  AND U15124 ( .A(n13779), .B(n13780), .Z(n13757) );
  NANDN U15125 ( .A(n13781), .B(n13782), .Z(n13780) );
  NANDN U15126 ( .A(n13783), .B(n13784), .Z(n13782) );
  AND U15127 ( .A(B[378]), .B(A[3]), .Z(n13759) );
  XNOR U15128 ( .A(n13749), .B(n13785), .Z(n13760) );
  XNOR U15129 ( .A(n13747), .B(n13750), .Z(n13785) );
  NAND U15130 ( .A(A[2]), .B(B[379]), .Z(n13750) );
  NANDN U15131 ( .A(n13786), .B(n13787), .Z(n13747) );
  AND U15132 ( .A(A[0]), .B(B[380]), .Z(n13787) );
  XOR U15133 ( .A(n13752), .B(n13788), .Z(n13749) );
  NAND U15134 ( .A(A[0]), .B(B[381]), .Z(n13788) );
  NAND U15135 ( .A(B[380]), .B(A[1]), .Z(n13752) );
  NAND U15136 ( .A(n13789), .B(n13790), .Z(n1407) );
  NANDN U15137 ( .A(n13791), .B(n13792), .Z(n13790) );
  OR U15138 ( .A(n13793), .B(n13794), .Z(n13792) );
  NAND U15139 ( .A(n13794), .B(n13793), .Z(n13789) );
  XOR U15140 ( .A(n1411), .B(n1410), .Z(\A1[378] ) );
  XOR U15141 ( .A(n13794), .B(n13795), .Z(n1410) );
  XNOR U15142 ( .A(n13793), .B(n13791), .Z(n13795) );
  AND U15143 ( .A(n13796), .B(n13797), .Z(n13791) );
  NANDN U15144 ( .A(n13798), .B(n13799), .Z(n13797) );
  NANDN U15145 ( .A(n13800), .B(n13801), .Z(n13799) );
  AND U15146 ( .A(B[377]), .B(A[3]), .Z(n13793) );
  XNOR U15147 ( .A(n13783), .B(n13802), .Z(n13794) );
  XNOR U15148 ( .A(n13781), .B(n13784), .Z(n13802) );
  NAND U15149 ( .A(A[2]), .B(B[378]), .Z(n13784) );
  NANDN U15150 ( .A(n13803), .B(n13804), .Z(n13781) );
  AND U15151 ( .A(A[0]), .B(B[379]), .Z(n13804) );
  XOR U15152 ( .A(n13786), .B(n13805), .Z(n13783) );
  NAND U15153 ( .A(A[0]), .B(B[380]), .Z(n13805) );
  NAND U15154 ( .A(B[379]), .B(A[1]), .Z(n13786) );
  NAND U15155 ( .A(n13806), .B(n13807), .Z(n1411) );
  NANDN U15156 ( .A(n13808), .B(n13809), .Z(n13807) );
  OR U15157 ( .A(n13810), .B(n13811), .Z(n13809) );
  NAND U15158 ( .A(n13811), .B(n13810), .Z(n13806) );
  XOR U15159 ( .A(n1413), .B(n1412), .Z(\A1[377] ) );
  XOR U15160 ( .A(n13811), .B(n13812), .Z(n1412) );
  XNOR U15161 ( .A(n13810), .B(n13808), .Z(n13812) );
  AND U15162 ( .A(n13813), .B(n13814), .Z(n13808) );
  NANDN U15163 ( .A(n13815), .B(n13816), .Z(n13814) );
  NANDN U15164 ( .A(n13817), .B(n13818), .Z(n13816) );
  AND U15165 ( .A(B[376]), .B(A[3]), .Z(n13810) );
  XNOR U15166 ( .A(n13800), .B(n13819), .Z(n13811) );
  XNOR U15167 ( .A(n13798), .B(n13801), .Z(n13819) );
  NAND U15168 ( .A(A[2]), .B(B[377]), .Z(n13801) );
  NANDN U15169 ( .A(n13820), .B(n13821), .Z(n13798) );
  AND U15170 ( .A(A[0]), .B(B[378]), .Z(n13821) );
  XOR U15171 ( .A(n13803), .B(n13822), .Z(n13800) );
  NAND U15172 ( .A(A[0]), .B(B[379]), .Z(n13822) );
  NAND U15173 ( .A(B[378]), .B(A[1]), .Z(n13803) );
  NAND U15174 ( .A(n13823), .B(n13824), .Z(n1413) );
  NANDN U15175 ( .A(n13825), .B(n13826), .Z(n13824) );
  OR U15176 ( .A(n13827), .B(n13828), .Z(n13826) );
  NAND U15177 ( .A(n13828), .B(n13827), .Z(n13823) );
  XOR U15178 ( .A(n1415), .B(n1414), .Z(\A1[376] ) );
  XOR U15179 ( .A(n13828), .B(n13829), .Z(n1414) );
  XNOR U15180 ( .A(n13827), .B(n13825), .Z(n13829) );
  AND U15181 ( .A(n13830), .B(n13831), .Z(n13825) );
  NANDN U15182 ( .A(n13832), .B(n13833), .Z(n13831) );
  NANDN U15183 ( .A(n13834), .B(n13835), .Z(n13833) );
  AND U15184 ( .A(B[375]), .B(A[3]), .Z(n13827) );
  XNOR U15185 ( .A(n13817), .B(n13836), .Z(n13828) );
  XNOR U15186 ( .A(n13815), .B(n13818), .Z(n13836) );
  NAND U15187 ( .A(A[2]), .B(B[376]), .Z(n13818) );
  NANDN U15188 ( .A(n13837), .B(n13838), .Z(n13815) );
  AND U15189 ( .A(A[0]), .B(B[377]), .Z(n13838) );
  XOR U15190 ( .A(n13820), .B(n13839), .Z(n13817) );
  NAND U15191 ( .A(A[0]), .B(B[378]), .Z(n13839) );
  NAND U15192 ( .A(B[377]), .B(A[1]), .Z(n13820) );
  NAND U15193 ( .A(n13840), .B(n13841), .Z(n1415) );
  NANDN U15194 ( .A(n13842), .B(n13843), .Z(n13841) );
  OR U15195 ( .A(n13844), .B(n13845), .Z(n13843) );
  NAND U15196 ( .A(n13845), .B(n13844), .Z(n13840) );
  XOR U15197 ( .A(n1417), .B(n1416), .Z(\A1[375] ) );
  XOR U15198 ( .A(n13845), .B(n13846), .Z(n1416) );
  XNOR U15199 ( .A(n13844), .B(n13842), .Z(n13846) );
  AND U15200 ( .A(n13847), .B(n13848), .Z(n13842) );
  NANDN U15201 ( .A(n13849), .B(n13850), .Z(n13848) );
  NANDN U15202 ( .A(n13851), .B(n13852), .Z(n13850) );
  AND U15203 ( .A(B[374]), .B(A[3]), .Z(n13844) );
  XNOR U15204 ( .A(n13834), .B(n13853), .Z(n13845) );
  XNOR U15205 ( .A(n13832), .B(n13835), .Z(n13853) );
  NAND U15206 ( .A(A[2]), .B(B[375]), .Z(n13835) );
  NANDN U15207 ( .A(n13854), .B(n13855), .Z(n13832) );
  AND U15208 ( .A(A[0]), .B(B[376]), .Z(n13855) );
  XOR U15209 ( .A(n13837), .B(n13856), .Z(n13834) );
  NAND U15210 ( .A(A[0]), .B(B[377]), .Z(n13856) );
  NAND U15211 ( .A(B[376]), .B(A[1]), .Z(n13837) );
  NAND U15212 ( .A(n13857), .B(n13858), .Z(n1417) );
  NANDN U15213 ( .A(n13859), .B(n13860), .Z(n13858) );
  OR U15214 ( .A(n13861), .B(n13862), .Z(n13860) );
  NAND U15215 ( .A(n13862), .B(n13861), .Z(n13857) );
  XOR U15216 ( .A(n1419), .B(n1418), .Z(\A1[374] ) );
  XOR U15217 ( .A(n13862), .B(n13863), .Z(n1418) );
  XNOR U15218 ( .A(n13861), .B(n13859), .Z(n13863) );
  AND U15219 ( .A(n13864), .B(n13865), .Z(n13859) );
  NANDN U15220 ( .A(n13866), .B(n13867), .Z(n13865) );
  NANDN U15221 ( .A(n13868), .B(n13869), .Z(n13867) );
  AND U15222 ( .A(B[373]), .B(A[3]), .Z(n13861) );
  XNOR U15223 ( .A(n13851), .B(n13870), .Z(n13862) );
  XNOR U15224 ( .A(n13849), .B(n13852), .Z(n13870) );
  NAND U15225 ( .A(A[2]), .B(B[374]), .Z(n13852) );
  NANDN U15226 ( .A(n13871), .B(n13872), .Z(n13849) );
  AND U15227 ( .A(A[0]), .B(B[375]), .Z(n13872) );
  XOR U15228 ( .A(n13854), .B(n13873), .Z(n13851) );
  NAND U15229 ( .A(A[0]), .B(B[376]), .Z(n13873) );
  NAND U15230 ( .A(B[375]), .B(A[1]), .Z(n13854) );
  NAND U15231 ( .A(n13874), .B(n13875), .Z(n1419) );
  NANDN U15232 ( .A(n13876), .B(n13877), .Z(n13875) );
  OR U15233 ( .A(n13878), .B(n13879), .Z(n13877) );
  NAND U15234 ( .A(n13879), .B(n13878), .Z(n13874) );
  XOR U15235 ( .A(n1421), .B(n1420), .Z(\A1[373] ) );
  XOR U15236 ( .A(n13879), .B(n13880), .Z(n1420) );
  XNOR U15237 ( .A(n13878), .B(n13876), .Z(n13880) );
  AND U15238 ( .A(n13881), .B(n13882), .Z(n13876) );
  NANDN U15239 ( .A(n13883), .B(n13884), .Z(n13882) );
  NANDN U15240 ( .A(n13885), .B(n13886), .Z(n13884) );
  AND U15241 ( .A(B[372]), .B(A[3]), .Z(n13878) );
  XNOR U15242 ( .A(n13868), .B(n13887), .Z(n13879) );
  XNOR U15243 ( .A(n13866), .B(n13869), .Z(n13887) );
  NAND U15244 ( .A(A[2]), .B(B[373]), .Z(n13869) );
  NANDN U15245 ( .A(n13888), .B(n13889), .Z(n13866) );
  AND U15246 ( .A(A[0]), .B(B[374]), .Z(n13889) );
  XOR U15247 ( .A(n13871), .B(n13890), .Z(n13868) );
  NAND U15248 ( .A(A[0]), .B(B[375]), .Z(n13890) );
  NAND U15249 ( .A(B[374]), .B(A[1]), .Z(n13871) );
  NAND U15250 ( .A(n13891), .B(n13892), .Z(n1421) );
  NANDN U15251 ( .A(n13893), .B(n13894), .Z(n13892) );
  OR U15252 ( .A(n13895), .B(n13896), .Z(n13894) );
  NAND U15253 ( .A(n13896), .B(n13895), .Z(n13891) );
  XOR U15254 ( .A(n1423), .B(n1422), .Z(\A1[372] ) );
  XOR U15255 ( .A(n13896), .B(n13897), .Z(n1422) );
  XNOR U15256 ( .A(n13895), .B(n13893), .Z(n13897) );
  AND U15257 ( .A(n13898), .B(n13899), .Z(n13893) );
  NANDN U15258 ( .A(n13900), .B(n13901), .Z(n13899) );
  NANDN U15259 ( .A(n13902), .B(n13903), .Z(n13901) );
  AND U15260 ( .A(B[371]), .B(A[3]), .Z(n13895) );
  XNOR U15261 ( .A(n13885), .B(n13904), .Z(n13896) );
  XNOR U15262 ( .A(n13883), .B(n13886), .Z(n13904) );
  NAND U15263 ( .A(A[2]), .B(B[372]), .Z(n13886) );
  NANDN U15264 ( .A(n13905), .B(n13906), .Z(n13883) );
  AND U15265 ( .A(A[0]), .B(B[373]), .Z(n13906) );
  XOR U15266 ( .A(n13888), .B(n13907), .Z(n13885) );
  NAND U15267 ( .A(A[0]), .B(B[374]), .Z(n13907) );
  NAND U15268 ( .A(B[373]), .B(A[1]), .Z(n13888) );
  NAND U15269 ( .A(n13908), .B(n13909), .Z(n1423) );
  NANDN U15270 ( .A(n13910), .B(n13911), .Z(n13909) );
  OR U15271 ( .A(n13912), .B(n13913), .Z(n13911) );
  NAND U15272 ( .A(n13913), .B(n13912), .Z(n13908) );
  XOR U15273 ( .A(n1425), .B(n1424), .Z(\A1[371] ) );
  XOR U15274 ( .A(n13913), .B(n13914), .Z(n1424) );
  XNOR U15275 ( .A(n13912), .B(n13910), .Z(n13914) );
  AND U15276 ( .A(n13915), .B(n13916), .Z(n13910) );
  NANDN U15277 ( .A(n13917), .B(n13918), .Z(n13916) );
  NANDN U15278 ( .A(n13919), .B(n13920), .Z(n13918) );
  AND U15279 ( .A(B[370]), .B(A[3]), .Z(n13912) );
  XNOR U15280 ( .A(n13902), .B(n13921), .Z(n13913) );
  XNOR U15281 ( .A(n13900), .B(n13903), .Z(n13921) );
  NAND U15282 ( .A(A[2]), .B(B[371]), .Z(n13903) );
  NANDN U15283 ( .A(n13922), .B(n13923), .Z(n13900) );
  AND U15284 ( .A(A[0]), .B(B[372]), .Z(n13923) );
  XOR U15285 ( .A(n13905), .B(n13924), .Z(n13902) );
  NAND U15286 ( .A(A[0]), .B(B[373]), .Z(n13924) );
  NAND U15287 ( .A(B[372]), .B(A[1]), .Z(n13905) );
  NAND U15288 ( .A(n13925), .B(n13926), .Z(n1425) );
  NANDN U15289 ( .A(n13927), .B(n13928), .Z(n13926) );
  OR U15290 ( .A(n13929), .B(n13930), .Z(n13928) );
  NAND U15291 ( .A(n13930), .B(n13929), .Z(n13925) );
  XOR U15292 ( .A(n1427), .B(n1426), .Z(\A1[370] ) );
  XOR U15293 ( .A(n13930), .B(n13931), .Z(n1426) );
  XNOR U15294 ( .A(n13929), .B(n13927), .Z(n13931) );
  AND U15295 ( .A(n13932), .B(n13933), .Z(n13927) );
  NANDN U15296 ( .A(n13934), .B(n13935), .Z(n13933) );
  NANDN U15297 ( .A(n13936), .B(n13937), .Z(n13935) );
  AND U15298 ( .A(B[369]), .B(A[3]), .Z(n13929) );
  XNOR U15299 ( .A(n13919), .B(n13938), .Z(n13930) );
  XNOR U15300 ( .A(n13917), .B(n13920), .Z(n13938) );
  NAND U15301 ( .A(A[2]), .B(B[370]), .Z(n13920) );
  NANDN U15302 ( .A(n13939), .B(n13940), .Z(n13917) );
  AND U15303 ( .A(A[0]), .B(B[371]), .Z(n13940) );
  XOR U15304 ( .A(n13922), .B(n13941), .Z(n13919) );
  NAND U15305 ( .A(A[0]), .B(B[372]), .Z(n13941) );
  NAND U15306 ( .A(B[371]), .B(A[1]), .Z(n13922) );
  NAND U15307 ( .A(n13942), .B(n13943), .Z(n1427) );
  NANDN U15308 ( .A(n13944), .B(n13945), .Z(n13943) );
  OR U15309 ( .A(n13946), .B(n13947), .Z(n13945) );
  NAND U15310 ( .A(n13947), .B(n13946), .Z(n13942) );
  XOR U15311 ( .A(n1409), .B(n1408), .Z(\A1[36] ) );
  XOR U15312 ( .A(n13777), .B(n13948), .Z(n1408) );
  XNOR U15313 ( .A(n13776), .B(n13774), .Z(n13948) );
  AND U15314 ( .A(n13949), .B(n13950), .Z(n13774) );
  NANDN U15315 ( .A(n13951), .B(n13952), .Z(n13950) );
  NANDN U15316 ( .A(n13953), .B(n13954), .Z(n13952) );
  AND U15317 ( .A(B[35]), .B(A[3]), .Z(n13776) );
  XNOR U15318 ( .A(n13766), .B(n13955), .Z(n13777) );
  XNOR U15319 ( .A(n13764), .B(n13767), .Z(n13955) );
  NAND U15320 ( .A(A[2]), .B(B[36]), .Z(n13767) );
  NANDN U15321 ( .A(n13956), .B(n13957), .Z(n13764) );
  AND U15322 ( .A(A[0]), .B(B[37]), .Z(n13957) );
  XOR U15323 ( .A(n13769), .B(n13958), .Z(n13766) );
  NAND U15324 ( .A(A[0]), .B(B[38]), .Z(n13958) );
  NAND U15325 ( .A(B[37]), .B(A[1]), .Z(n13769) );
  NAND U15326 ( .A(n13959), .B(n13960), .Z(n1409) );
  NANDN U15327 ( .A(n13961), .B(n13962), .Z(n13960) );
  OR U15328 ( .A(n13963), .B(n13964), .Z(n13962) );
  NAND U15329 ( .A(n13964), .B(n13963), .Z(n13959) );
  XOR U15330 ( .A(n1429), .B(n1428), .Z(\A1[369] ) );
  XOR U15331 ( .A(n13947), .B(n13965), .Z(n1428) );
  XNOR U15332 ( .A(n13946), .B(n13944), .Z(n13965) );
  AND U15333 ( .A(n13966), .B(n13967), .Z(n13944) );
  NANDN U15334 ( .A(n13968), .B(n13969), .Z(n13967) );
  NANDN U15335 ( .A(n13970), .B(n13971), .Z(n13969) );
  AND U15336 ( .A(B[368]), .B(A[3]), .Z(n13946) );
  XNOR U15337 ( .A(n13936), .B(n13972), .Z(n13947) );
  XNOR U15338 ( .A(n13934), .B(n13937), .Z(n13972) );
  NAND U15339 ( .A(A[2]), .B(B[369]), .Z(n13937) );
  NANDN U15340 ( .A(n13973), .B(n13974), .Z(n13934) );
  AND U15341 ( .A(A[0]), .B(B[370]), .Z(n13974) );
  XOR U15342 ( .A(n13939), .B(n13975), .Z(n13936) );
  NAND U15343 ( .A(A[0]), .B(B[371]), .Z(n13975) );
  NAND U15344 ( .A(B[370]), .B(A[1]), .Z(n13939) );
  NAND U15345 ( .A(n13976), .B(n13977), .Z(n1429) );
  NANDN U15346 ( .A(n13978), .B(n13979), .Z(n13977) );
  OR U15347 ( .A(n13980), .B(n13981), .Z(n13979) );
  NAND U15348 ( .A(n13981), .B(n13980), .Z(n13976) );
  XOR U15349 ( .A(n1433), .B(n1432), .Z(\A1[368] ) );
  XOR U15350 ( .A(n13981), .B(n13982), .Z(n1432) );
  XNOR U15351 ( .A(n13980), .B(n13978), .Z(n13982) );
  AND U15352 ( .A(n13983), .B(n13984), .Z(n13978) );
  NANDN U15353 ( .A(n13985), .B(n13986), .Z(n13984) );
  NANDN U15354 ( .A(n13987), .B(n13988), .Z(n13986) );
  AND U15355 ( .A(B[367]), .B(A[3]), .Z(n13980) );
  XNOR U15356 ( .A(n13970), .B(n13989), .Z(n13981) );
  XNOR U15357 ( .A(n13968), .B(n13971), .Z(n13989) );
  NAND U15358 ( .A(A[2]), .B(B[368]), .Z(n13971) );
  NANDN U15359 ( .A(n13990), .B(n13991), .Z(n13968) );
  AND U15360 ( .A(A[0]), .B(B[369]), .Z(n13991) );
  XOR U15361 ( .A(n13973), .B(n13992), .Z(n13970) );
  NAND U15362 ( .A(A[0]), .B(B[370]), .Z(n13992) );
  NAND U15363 ( .A(B[369]), .B(A[1]), .Z(n13973) );
  NAND U15364 ( .A(n13993), .B(n13994), .Z(n1433) );
  NANDN U15365 ( .A(n13995), .B(n13996), .Z(n13994) );
  OR U15366 ( .A(n13997), .B(n13998), .Z(n13996) );
  NAND U15367 ( .A(n13998), .B(n13997), .Z(n13993) );
  XOR U15368 ( .A(n1435), .B(n1434), .Z(\A1[367] ) );
  XOR U15369 ( .A(n13998), .B(n13999), .Z(n1434) );
  XNOR U15370 ( .A(n13997), .B(n13995), .Z(n13999) );
  AND U15371 ( .A(n14000), .B(n14001), .Z(n13995) );
  NANDN U15372 ( .A(n14002), .B(n14003), .Z(n14001) );
  NANDN U15373 ( .A(n14004), .B(n14005), .Z(n14003) );
  AND U15374 ( .A(B[366]), .B(A[3]), .Z(n13997) );
  XNOR U15375 ( .A(n13987), .B(n14006), .Z(n13998) );
  XNOR U15376 ( .A(n13985), .B(n13988), .Z(n14006) );
  NAND U15377 ( .A(A[2]), .B(B[367]), .Z(n13988) );
  NANDN U15378 ( .A(n14007), .B(n14008), .Z(n13985) );
  AND U15379 ( .A(A[0]), .B(B[368]), .Z(n14008) );
  XOR U15380 ( .A(n13990), .B(n14009), .Z(n13987) );
  NAND U15381 ( .A(A[0]), .B(B[369]), .Z(n14009) );
  NAND U15382 ( .A(B[368]), .B(A[1]), .Z(n13990) );
  NAND U15383 ( .A(n14010), .B(n14011), .Z(n1435) );
  NANDN U15384 ( .A(n14012), .B(n14013), .Z(n14011) );
  OR U15385 ( .A(n14014), .B(n14015), .Z(n14013) );
  NAND U15386 ( .A(n14015), .B(n14014), .Z(n14010) );
  XOR U15387 ( .A(n1437), .B(n1436), .Z(\A1[366] ) );
  XOR U15388 ( .A(n14015), .B(n14016), .Z(n1436) );
  XNOR U15389 ( .A(n14014), .B(n14012), .Z(n14016) );
  AND U15390 ( .A(n14017), .B(n14018), .Z(n14012) );
  NANDN U15391 ( .A(n14019), .B(n14020), .Z(n14018) );
  NANDN U15392 ( .A(n14021), .B(n14022), .Z(n14020) );
  AND U15393 ( .A(B[365]), .B(A[3]), .Z(n14014) );
  XNOR U15394 ( .A(n14004), .B(n14023), .Z(n14015) );
  XNOR U15395 ( .A(n14002), .B(n14005), .Z(n14023) );
  NAND U15396 ( .A(A[2]), .B(B[366]), .Z(n14005) );
  NANDN U15397 ( .A(n14024), .B(n14025), .Z(n14002) );
  AND U15398 ( .A(A[0]), .B(B[367]), .Z(n14025) );
  XOR U15399 ( .A(n14007), .B(n14026), .Z(n14004) );
  NAND U15400 ( .A(A[0]), .B(B[368]), .Z(n14026) );
  NAND U15401 ( .A(B[367]), .B(A[1]), .Z(n14007) );
  NAND U15402 ( .A(n14027), .B(n14028), .Z(n1437) );
  NANDN U15403 ( .A(n14029), .B(n14030), .Z(n14028) );
  OR U15404 ( .A(n14031), .B(n14032), .Z(n14030) );
  NAND U15405 ( .A(n14032), .B(n14031), .Z(n14027) );
  XOR U15406 ( .A(n1439), .B(n1438), .Z(\A1[365] ) );
  XOR U15407 ( .A(n14032), .B(n14033), .Z(n1438) );
  XNOR U15408 ( .A(n14031), .B(n14029), .Z(n14033) );
  AND U15409 ( .A(n14034), .B(n14035), .Z(n14029) );
  NANDN U15410 ( .A(n14036), .B(n14037), .Z(n14035) );
  NANDN U15411 ( .A(n14038), .B(n14039), .Z(n14037) );
  AND U15412 ( .A(B[364]), .B(A[3]), .Z(n14031) );
  XNOR U15413 ( .A(n14021), .B(n14040), .Z(n14032) );
  XNOR U15414 ( .A(n14019), .B(n14022), .Z(n14040) );
  NAND U15415 ( .A(A[2]), .B(B[365]), .Z(n14022) );
  NANDN U15416 ( .A(n14041), .B(n14042), .Z(n14019) );
  AND U15417 ( .A(A[0]), .B(B[366]), .Z(n14042) );
  XOR U15418 ( .A(n14024), .B(n14043), .Z(n14021) );
  NAND U15419 ( .A(A[0]), .B(B[367]), .Z(n14043) );
  NAND U15420 ( .A(B[366]), .B(A[1]), .Z(n14024) );
  NAND U15421 ( .A(n14044), .B(n14045), .Z(n1439) );
  NANDN U15422 ( .A(n14046), .B(n14047), .Z(n14045) );
  OR U15423 ( .A(n14048), .B(n14049), .Z(n14047) );
  NAND U15424 ( .A(n14049), .B(n14048), .Z(n14044) );
  XOR U15425 ( .A(n1441), .B(n1440), .Z(\A1[364] ) );
  XOR U15426 ( .A(n14049), .B(n14050), .Z(n1440) );
  XNOR U15427 ( .A(n14048), .B(n14046), .Z(n14050) );
  AND U15428 ( .A(n14051), .B(n14052), .Z(n14046) );
  NANDN U15429 ( .A(n14053), .B(n14054), .Z(n14052) );
  NANDN U15430 ( .A(n14055), .B(n14056), .Z(n14054) );
  AND U15431 ( .A(B[363]), .B(A[3]), .Z(n14048) );
  XNOR U15432 ( .A(n14038), .B(n14057), .Z(n14049) );
  XNOR U15433 ( .A(n14036), .B(n14039), .Z(n14057) );
  NAND U15434 ( .A(A[2]), .B(B[364]), .Z(n14039) );
  NANDN U15435 ( .A(n14058), .B(n14059), .Z(n14036) );
  AND U15436 ( .A(A[0]), .B(B[365]), .Z(n14059) );
  XOR U15437 ( .A(n14041), .B(n14060), .Z(n14038) );
  NAND U15438 ( .A(A[0]), .B(B[366]), .Z(n14060) );
  NAND U15439 ( .A(B[365]), .B(A[1]), .Z(n14041) );
  NAND U15440 ( .A(n14061), .B(n14062), .Z(n1441) );
  NANDN U15441 ( .A(n14063), .B(n14064), .Z(n14062) );
  OR U15442 ( .A(n14065), .B(n14066), .Z(n14064) );
  NAND U15443 ( .A(n14066), .B(n14065), .Z(n14061) );
  XOR U15444 ( .A(n1443), .B(n1442), .Z(\A1[363] ) );
  XOR U15445 ( .A(n14066), .B(n14067), .Z(n1442) );
  XNOR U15446 ( .A(n14065), .B(n14063), .Z(n14067) );
  AND U15447 ( .A(n14068), .B(n14069), .Z(n14063) );
  NANDN U15448 ( .A(n14070), .B(n14071), .Z(n14069) );
  NANDN U15449 ( .A(n14072), .B(n14073), .Z(n14071) );
  AND U15450 ( .A(B[362]), .B(A[3]), .Z(n14065) );
  XNOR U15451 ( .A(n14055), .B(n14074), .Z(n14066) );
  XNOR U15452 ( .A(n14053), .B(n14056), .Z(n14074) );
  NAND U15453 ( .A(A[2]), .B(B[363]), .Z(n14056) );
  NANDN U15454 ( .A(n14075), .B(n14076), .Z(n14053) );
  AND U15455 ( .A(A[0]), .B(B[364]), .Z(n14076) );
  XOR U15456 ( .A(n14058), .B(n14077), .Z(n14055) );
  NAND U15457 ( .A(A[0]), .B(B[365]), .Z(n14077) );
  NAND U15458 ( .A(B[364]), .B(A[1]), .Z(n14058) );
  NAND U15459 ( .A(n14078), .B(n14079), .Z(n1443) );
  NANDN U15460 ( .A(n14080), .B(n14081), .Z(n14079) );
  OR U15461 ( .A(n14082), .B(n14083), .Z(n14081) );
  NAND U15462 ( .A(n14083), .B(n14082), .Z(n14078) );
  XOR U15463 ( .A(n1445), .B(n1444), .Z(\A1[362] ) );
  XOR U15464 ( .A(n14083), .B(n14084), .Z(n1444) );
  XNOR U15465 ( .A(n14082), .B(n14080), .Z(n14084) );
  AND U15466 ( .A(n14085), .B(n14086), .Z(n14080) );
  NANDN U15467 ( .A(n14087), .B(n14088), .Z(n14086) );
  NANDN U15468 ( .A(n14089), .B(n14090), .Z(n14088) );
  AND U15469 ( .A(B[361]), .B(A[3]), .Z(n14082) );
  XNOR U15470 ( .A(n14072), .B(n14091), .Z(n14083) );
  XNOR U15471 ( .A(n14070), .B(n14073), .Z(n14091) );
  NAND U15472 ( .A(A[2]), .B(B[362]), .Z(n14073) );
  NANDN U15473 ( .A(n14092), .B(n14093), .Z(n14070) );
  AND U15474 ( .A(A[0]), .B(B[363]), .Z(n14093) );
  XOR U15475 ( .A(n14075), .B(n14094), .Z(n14072) );
  NAND U15476 ( .A(A[0]), .B(B[364]), .Z(n14094) );
  NAND U15477 ( .A(B[363]), .B(A[1]), .Z(n14075) );
  NAND U15478 ( .A(n14095), .B(n14096), .Z(n1445) );
  NANDN U15479 ( .A(n14097), .B(n14098), .Z(n14096) );
  OR U15480 ( .A(n14099), .B(n14100), .Z(n14098) );
  NAND U15481 ( .A(n14100), .B(n14099), .Z(n14095) );
  XOR U15482 ( .A(n1447), .B(n1446), .Z(\A1[361] ) );
  XOR U15483 ( .A(n14100), .B(n14101), .Z(n1446) );
  XNOR U15484 ( .A(n14099), .B(n14097), .Z(n14101) );
  AND U15485 ( .A(n14102), .B(n14103), .Z(n14097) );
  NANDN U15486 ( .A(n14104), .B(n14105), .Z(n14103) );
  NANDN U15487 ( .A(n14106), .B(n14107), .Z(n14105) );
  AND U15488 ( .A(B[360]), .B(A[3]), .Z(n14099) );
  XNOR U15489 ( .A(n14089), .B(n14108), .Z(n14100) );
  XNOR U15490 ( .A(n14087), .B(n14090), .Z(n14108) );
  NAND U15491 ( .A(A[2]), .B(B[361]), .Z(n14090) );
  NANDN U15492 ( .A(n14109), .B(n14110), .Z(n14087) );
  AND U15493 ( .A(A[0]), .B(B[362]), .Z(n14110) );
  XOR U15494 ( .A(n14092), .B(n14111), .Z(n14089) );
  NAND U15495 ( .A(A[0]), .B(B[363]), .Z(n14111) );
  NAND U15496 ( .A(B[362]), .B(A[1]), .Z(n14092) );
  NAND U15497 ( .A(n14112), .B(n14113), .Z(n1447) );
  NANDN U15498 ( .A(n14114), .B(n14115), .Z(n14113) );
  OR U15499 ( .A(n14116), .B(n14117), .Z(n14115) );
  NAND U15500 ( .A(n14117), .B(n14116), .Z(n14112) );
  XOR U15501 ( .A(n1449), .B(n1448), .Z(\A1[360] ) );
  XOR U15502 ( .A(n14117), .B(n14118), .Z(n1448) );
  XNOR U15503 ( .A(n14116), .B(n14114), .Z(n14118) );
  AND U15504 ( .A(n14119), .B(n14120), .Z(n14114) );
  NANDN U15505 ( .A(n14121), .B(n14122), .Z(n14120) );
  NANDN U15506 ( .A(n14123), .B(n14124), .Z(n14122) );
  AND U15507 ( .A(B[359]), .B(A[3]), .Z(n14116) );
  XNOR U15508 ( .A(n14106), .B(n14125), .Z(n14117) );
  XNOR U15509 ( .A(n14104), .B(n14107), .Z(n14125) );
  NAND U15510 ( .A(A[2]), .B(B[360]), .Z(n14107) );
  NANDN U15511 ( .A(n14126), .B(n14127), .Z(n14104) );
  AND U15512 ( .A(A[0]), .B(B[361]), .Z(n14127) );
  XOR U15513 ( .A(n14109), .B(n14128), .Z(n14106) );
  NAND U15514 ( .A(A[0]), .B(B[362]), .Z(n14128) );
  NAND U15515 ( .A(B[361]), .B(A[1]), .Z(n14109) );
  NAND U15516 ( .A(n14129), .B(n14130), .Z(n1449) );
  NANDN U15517 ( .A(n14131), .B(n14132), .Z(n14130) );
  OR U15518 ( .A(n14133), .B(n14134), .Z(n14132) );
  NAND U15519 ( .A(n14134), .B(n14133), .Z(n14129) );
  XOR U15520 ( .A(n1431), .B(n1430), .Z(\A1[35] ) );
  XOR U15521 ( .A(n13964), .B(n14135), .Z(n1430) );
  XNOR U15522 ( .A(n13963), .B(n13961), .Z(n14135) );
  AND U15523 ( .A(n14136), .B(n14137), .Z(n13961) );
  NANDN U15524 ( .A(n14138), .B(n14139), .Z(n14137) );
  NANDN U15525 ( .A(n14140), .B(n14141), .Z(n14139) );
  AND U15526 ( .A(B[34]), .B(A[3]), .Z(n13963) );
  XNOR U15527 ( .A(n13953), .B(n14142), .Z(n13964) );
  XNOR U15528 ( .A(n13951), .B(n13954), .Z(n14142) );
  NAND U15529 ( .A(A[2]), .B(B[35]), .Z(n13954) );
  NANDN U15530 ( .A(n14143), .B(n14144), .Z(n13951) );
  AND U15531 ( .A(A[0]), .B(B[36]), .Z(n14144) );
  XOR U15532 ( .A(n13956), .B(n14145), .Z(n13953) );
  NAND U15533 ( .A(A[0]), .B(B[37]), .Z(n14145) );
  NAND U15534 ( .A(B[36]), .B(A[1]), .Z(n13956) );
  NAND U15535 ( .A(n14146), .B(n14147), .Z(n1431) );
  NANDN U15536 ( .A(n14148), .B(n14149), .Z(n14147) );
  OR U15537 ( .A(n14150), .B(n14151), .Z(n14149) );
  NAND U15538 ( .A(n14151), .B(n14150), .Z(n14146) );
  XOR U15539 ( .A(n1451), .B(n1450), .Z(\A1[359] ) );
  XOR U15540 ( .A(n14134), .B(n14152), .Z(n1450) );
  XNOR U15541 ( .A(n14133), .B(n14131), .Z(n14152) );
  AND U15542 ( .A(n14153), .B(n14154), .Z(n14131) );
  NANDN U15543 ( .A(n14155), .B(n14156), .Z(n14154) );
  NANDN U15544 ( .A(n14157), .B(n14158), .Z(n14156) );
  AND U15545 ( .A(B[358]), .B(A[3]), .Z(n14133) );
  XNOR U15546 ( .A(n14123), .B(n14159), .Z(n14134) );
  XNOR U15547 ( .A(n14121), .B(n14124), .Z(n14159) );
  NAND U15548 ( .A(A[2]), .B(B[359]), .Z(n14124) );
  NANDN U15549 ( .A(n14160), .B(n14161), .Z(n14121) );
  AND U15550 ( .A(A[0]), .B(B[360]), .Z(n14161) );
  XOR U15551 ( .A(n14126), .B(n14162), .Z(n14123) );
  NAND U15552 ( .A(A[0]), .B(B[361]), .Z(n14162) );
  NAND U15553 ( .A(B[360]), .B(A[1]), .Z(n14126) );
  NAND U15554 ( .A(n14163), .B(n14164), .Z(n1451) );
  NANDN U15555 ( .A(n14165), .B(n14166), .Z(n14164) );
  OR U15556 ( .A(n14167), .B(n14168), .Z(n14166) );
  NAND U15557 ( .A(n14168), .B(n14167), .Z(n14163) );
  XOR U15558 ( .A(n1455), .B(n1454), .Z(\A1[358] ) );
  XOR U15559 ( .A(n14168), .B(n14169), .Z(n1454) );
  XNOR U15560 ( .A(n14167), .B(n14165), .Z(n14169) );
  AND U15561 ( .A(n14170), .B(n14171), .Z(n14165) );
  NANDN U15562 ( .A(n14172), .B(n14173), .Z(n14171) );
  NANDN U15563 ( .A(n14174), .B(n14175), .Z(n14173) );
  AND U15564 ( .A(B[357]), .B(A[3]), .Z(n14167) );
  XNOR U15565 ( .A(n14157), .B(n14176), .Z(n14168) );
  XNOR U15566 ( .A(n14155), .B(n14158), .Z(n14176) );
  NAND U15567 ( .A(A[2]), .B(B[358]), .Z(n14158) );
  NANDN U15568 ( .A(n14177), .B(n14178), .Z(n14155) );
  AND U15569 ( .A(A[0]), .B(B[359]), .Z(n14178) );
  XOR U15570 ( .A(n14160), .B(n14179), .Z(n14157) );
  NAND U15571 ( .A(A[0]), .B(B[360]), .Z(n14179) );
  NAND U15572 ( .A(B[359]), .B(A[1]), .Z(n14160) );
  NAND U15573 ( .A(n14180), .B(n14181), .Z(n1455) );
  NANDN U15574 ( .A(n14182), .B(n14183), .Z(n14181) );
  OR U15575 ( .A(n14184), .B(n14185), .Z(n14183) );
  NAND U15576 ( .A(n14185), .B(n14184), .Z(n14180) );
  XOR U15577 ( .A(n1457), .B(n1456), .Z(\A1[357] ) );
  XOR U15578 ( .A(n14185), .B(n14186), .Z(n1456) );
  XNOR U15579 ( .A(n14184), .B(n14182), .Z(n14186) );
  AND U15580 ( .A(n14187), .B(n14188), .Z(n14182) );
  NANDN U15581 ( .A(n14189), .B(n14190), .Z(n14188) );
  NANDN U15582 ( .A(n14191), .B(n14192), .Z(n14190) );
  AND U15583 ( .A(B[356]), .B(A[3]), .Z(n14184) );
  XNOR U15584 ( .A(n14174), .B(n14193), .Z(n14185) );
  XNOR U15585 ( .A(n14172), .B(n14175), .Z(n14193) );
  NAND U15586 ( .A(A[2]), .B(B[357]), .Z(n14175) );
  NANDN U15587 ( .A(n14194), .B(n14195), .Z(n14172) );
  AND U15588 ( .A(A[0]), .B(B[358]), .Z(n14195) );
  XOR U15589 ( .A(n14177), .B(n14196), .Z(n14174) );
  NAND U15590 ( .A(A[0]), .B(B[359]), .Z(n14196) );
  NAND U15591 ( .A(B[358]), .B(A[1]), .Z(n14177) );
  NAND U15592 ( .A(n14197), .B(n14198), .Z(n1457) );
  NANDN U15593 ( .A(n14199), .B(n14200), .Z(n14198) );
  OR U15594 ( .A(n14201), .B(n14202), .Z(n14200) );
  NAND U15595 ( .A(n14202), .B(n14201), .Z(n14197) );
  XOR U15596 ( .A(n1459), .B(n1458), .Z(\A1[356] ) );
  XOR U15597 ( .A(n14202), .B(n14203), .Z(n1458) );
  XNOR U15598 ( .A(n14201), .B(n14199), .Z(n14203) );
  AND U15599 ( .A(n14204), .B(n14205), .Z(n14199) );
  NANDN U15600 ( .A(n14206), .B(n14207), .Z(n14205) );
  NANDN U15601 ( .A(n14208), .B(n14209), .Z(n14207) );
  AND U15602 ( .A(B[355]), .B(A[3]), .Z(n14201) );
  XNOR U15603 ( .A(n14191), .B(n14210), .Z(n14202) );
  XNOR U15604 ( .A(n14189), .B(n14192), .Z(n14210) );
  NAND U15605 ( .A(A[2]), .B(B[356]), .Z(n14192) );
  NANDN U15606 ( .A(n14211), .B(n14212), .Z(n14189) );
  AND U15607 ( .A(A[0]), .B(B[357]), .Z(n14212) );
  XOR U15608 ( .A(n14194), .B(n14213), .Z(n14191) );
  NAND U15609 ( .A(A[0]), .B(B[358]), .Z(n14213) );
  NAND U15610 ( .A(B[357]), .B(A[1]), .Z(n14194) );
  NAND U15611 ( .A(n14214), .B(n14215), .Z(n1459) );
  NANDN U15612 ( .A(n14216), .B(n14217), .Z(n14215) );
  OR U15613 ( .A(n14218), .B(n14219), .Z(n14217) );
  NAND U15614 ( .A(n14219), .B(n14218), .Z(n14214) );
  XOR U15615 ( .A(n1461), .B(n1460), .Z(\A1[355] ) );
  XOR U15616 ( .A(n14219), .B(n14220), .Z(n1460) );
  XNOR U15617 ( .A(n14218), .B(n14216), .Z(n14220) );
  AND U15618 ( .A(n14221), .B(n14222), .Z(n14216) );
  NANDN U15619 ( .A(n14223), .B(n14224), .Z(n14222) );
  NANDN U15620 ( .A(n14225), .B(n14226), .Z(n14224) );
  AND U15621 ( .A(B[354]), .B(A[3]), .Z(n14218) );
  XNOR U15622 ( .A(n14208), .B(n14227), .Z(n14219) );
  XNOR U15623 ( .A(n14206), .B(n14209), .Z(n14227) );
  NAND U15624 ( .A(A[2]), .B(B[355]), .Z(n14209) );
  NANDN U15625 ( .A(n14228), .B(n14229), .Z(n14206) );
  AND U15626 ( .A(A[0]), .B(B[356]), .Z(n14229) );
  XOR U15627 ( .A(n14211), .B(n14230), .Z(n14208) );
  NAND U15628 ( .A(A[0]), .B(B[357]), .Z(n14230) );
  NAND U15629 ( .A(B[356]), .B(A[1]), .Z(n14211) );
  NAND U15630 ( .A(n14231), .B(n14232), .Z(n1461) );
  NANDN U15631 ( .A(n14233), .B(n14234), .Z(n14232) );
  OR U15632 ( .A(n14235), .B(n14236), .Z(n14234) );
  NAND U15633 ( .A(n14236), .B(n14235), .Z(n14231) );
  XOR U15634 ( .A(n1463), .B(n1462), .Z(\A1[354] ) );
  XOR U15635 ( .A(n14236), .B(n14237), .Z(n1462) );
  XNOR U15636 ( .A(n14235), .B(n14233), .Z(n14237) );
  AND U15637 ( .A(n14238), .B(n14239), .Z(n14233) );
  NANDN U15638 ( .A(n14240), .B(n14241), .Z(n14239) );
  NANDN U15639 ( .A(n14242), .B(n14243), .Z(n14241) );
  AND U15640 ( .A(B[353]), .B(A[3]), .Z(n14235) );
  XNOR U15641 ( .A(n14225), .B(n14244), .Z(n14236) );
  XNOR U15642 ( .A(n14223), .B(n14226), .Z(n14244) );
  NAND U15643 ( .A(A[2]), .B(B[354]), .Z(n14226) );
  NANDN U15644 ( .A(n14245), .B(n14246), .Z(n14223) );
  AND U15645 ( .A(A[0]), .B(B[355]), .Z(n14246) );
  XOR U15646 ( .A(n14228), .B(n14247), .Z(n14225) );
  NAND U15647 ( .A(A[0]), .B(B[356]), .Z(n14247) );
  NAND U15648 ( .A(B[355]), .B(A[1]), .Z(n14228) );
  NAND U15649 ( .A(n14248), .B(n14249), .Z(n1463) );
  NANDN U15650 ( .A(n14250), .B(n14251), .Z(n14249) );
  OR U15651 ( .A(n14252), .B(n14253), .Z(n14251) );
  NAND U15652 ( .A(n14253), .B(n14252), .Z(n14248) );
  XOR U15653 ( .A(n1465), .B(n1464), .Z(\A1[353] ) );
  XOR U15654 ( .A(n14253), .B(n14254), .Z(n1464) );
  XNOR U15655 ( .A(n14252), .B(n14250), .Z(n14254) );
  AND U15656 ( .A(n14255), .B(n14256), .Z(n14250) );
  NANDN U15657 ( .A(n14257), .B(n14258), .Z(n14256) );
  NANDN U15658 ( .A(n14259), .B(n14260), .Z(n14258) );
  AND U15659 ( .A(B[352]), .B(A[3]), .Z(n14252) );
  XNOR U15660 ( .A(n14242), .B(n14261), .Z(n14253) );
  XNOR U15661 ( .A(n14240), .B(n14243), .Z(n14261) );
  NAND U15662 ( .A(A[2]), .B(B[353]), .Z(n14243) );
  NANDN U15663 ( .A(n14262), .B(n14263), .Z(n14240) );
  AND U15664 ( .A(A[0]), .B(B[354]), .Z(n14263) );
  XOR U15665 ( .A(n14245), .B(n14264), .Z(n14242) );
  NAND U15666 ( .A(A[0]), .B(B[355]), .Z(n14264) );
  NAND U15667 ( .A(B[354]), .B(A[1]), .Z(n14245) );
  NAND U15668 ( .A(n14265), .B(n14266), .Z(n1465) );
  NANDN U15669 ( .A(n14267), .B(n14268), .Z(n14266) );
  OR U15670 ( .A(n14269), .B(n14270), .Z(n14268) );
  NAND U15671 ( .A(n14270), .B(n14269), .Z(n14265) );
  XOR U15672 ( .A(n1467), .B(n1466), .Z(\A1[352] ) );
  XOR U15673 ( .A(n14270), .B(n14271), .Z(n1466) );
  XNOR U15674 ( .A(n14269), .B(n14267), .Z(n14271) );
  AND U15675 ( .A(n14272), .B(n14273), .Z(n14267) );
  NANDN U15676 ( .A(n14274), .B(n14275), .Z(n14273) );
  NANDN U15677 ( .A(n14276), .B(n14277), .Z(n14275) );
  AND U15678 ( .A(B[351]), .B(A[3]), .Z(n14269) );
  XNOR U15679 ( .A(n14259), .B(n14278), .Z(n14270) );
  XNOR U15680 ( .A(n14257), .B(n14260), .Z(n14278) );
  NAND U15681 ( .A(A[2]), .B(B[352]), .Z(n14260) );
  NANDN U15682 ( .A(n14279), .B(n14280), .Z(n14257) );
  AND U15683 ( .A(A[0]), .B(B[353]), .Z(n14280) );
  XOR U15684 ( .A(n14262), .B(n14281), .Z(n14259) );
  NAND U15685 ( .A(A[0]), .B(B[354]), .Z(n14281) );
  NAND U15686 ( .A(B[353]), .B(A[1]), .Z(n14262) );
  NAND U15687 ( .A(n14282), .B(n14283), .Z(n1467) );
  NANDN U15688 ( .A(n14284), .B(n14285), .Z(n14283) );
  OR U15689 ( .A(n14286), .B(n14287), .Z(n14285) );
  NAND U15690 ( .A(n14287), .B(n14286), .Z(n14282) );
  XOR U15691 ( .A(n1469), .B(n1468), .Z(\A1[351] ) );
  XOR U15692 ( .A(n14287), .B(n14288), .Z(n1468) );
  XNOR U15693 ( .A(n14286), .B(n14284), .Z(n14288) );
  AND U15694 ( .A(n14289), .B(n14290), .Z(n14284) );
  NANDN U15695 ( .A(n14291), .B(n14292), .Z(n14290) );
  NANDN U15696 ( .A(n14293), .B(n14294), .Z(n14292) );
  AND U15697 ( .A(B[350]), .B(A[3]), .Z(n14286) );
  XNOR U15698 ( .A(n14276), .B(n14295), .Z(n14287) );
  XNOR U15699 ( .A(n14274), .B(n14277), .Z(n14295) );
  NAND U15700 ( .A(A[2]), .B(B[351]), .Z(n14277) );
  NANDN U15701 ( .A(n14296), .B(n14297), .Z(n14274) );
  AND U15702 ( .A(A[0]), .B(B[352]), .Z(n14297) );
  XOR U15703 ( .A(n14279), .B(n14298), .Z(n14276) );
  NAND U15704 ( .A(A[0]), .B(B[353]), .Z(n14298) );
  NAND U15705 ( .A(B[352]), .B(A[1]), .Z(n14279) );
  NAND U15706 ( .A(n14299), .B(n14300), .Z(n1469) );
  NANDN U15707 ( .A(n14301), .B(n14302), .Z(n14300) );
  OR U15708 ( .A(n14303), .B(n14304), .Z(n14302) );
  NAND U15709 ( .A(n14304), .B(n14303), .Z(n14299) );
  XOR U15710 ( .A(n1471), .B(n1470), .Z(\A1[350] ) );
  XOR U15711 ( .A(n14304), .B(n14305), .Z(n1470) );
  XNOR U15712 ( .A(n14303), .B(n14301), .Z(n14305) );
  AND U15713 ( .A(n14306), .B(n14307), .Z(n14301) );
  NANDN U15714 ( .A(n14308), .B(n14309), .Z(n14307) );
  NANDN U15715 ( .A(n14310), .B(n14311), .Z(n14309) );
  AND U15716 ( .A(B[349]), .B(A[3]), .Z(n14303) );
  XNOR U15717 ( .A(n14293), .B(n14312), .Z(n14304) );
  XNOR U15718 ( .A(n14291), .B(n14294), .Z(n14312) );
  NAND U15719 ( .A(A[2]), .B(B[350]), .Z(n14294) );
  NANDN U15720 ( .A(n14313), .B(n14314), .Z(n14291) );
  AND U15721 ( .A(A[0]), .B(B[351]), .Z(n14314) );
  XOR U15722 ( .A(n14296), .B(n14315), .Z(n14293) );
  NAND U15723 ( .A(A[0]), .B(B[352]), .Z(n14315) );
  NAND U15724 ( .A(B[351]), .B(A[1]), .Z(n14296) );
  NAND U15725 ( .A(n14316), .B(n14317), .Z(n1471) );
  NANDN U15726 ( .A(n14318), .B(n14319), .Z(n14317) );
  OR U15727 ( .A(n14320), .B(n14321), .Z(n14319) );
  NAND U15728 ( .A(n14321), .B(n14320), .Z(n14316) );
  XOR U15729 ( .A(n1453), .B(n1452), .Z(\A1[34] ) );
  XOR U15730 ( .A(n14151), .B(n14322), .Z(n1452) );
  XNOR U15731 ( .A(n14150), .B(n14148), .Z(n14322) );
  AND U15732 ( .A(n14323), .B(n14324), .Z(n14148) );
  NANDN U15733 ( .A(n14325), .B(n14326), .Z(n14324) );
  NANDN U15734 ( .A(n14327), .B(n14328), .Z(n14326) );
  AND U15735 ( .A(B[33]), .B(A[3]), .Z(n14150) );
  XNOR U15736 ( .A(n14140), .B(n14329), .Z(n14151) );
  XNOR U15737 ( .A(n14138), .B(n14141), .Z(n14329) );
  NAND U15738 ( .A(A[2]), .B(B[34]), .Z(n14141) );
  NANDN U15739 ( .A(n14330), .B(n14331), .Z(n14138) );
  AND U15740 ( .A(A[0]), .B(B[35]), .Z(n14331) );
  XOR U15741 ( .A(n14143), .B(n14332), .Z(n14140) );
  NAND U15742 ( .A(A[0]), .B(B[36]), .Z(n14332) );
  NAND U15743 ( .A(B[35]), .B(A[1]), .Z(n14143) );
  NAND U15744 ( .A(n14333), .B(n14334), .Z(n1453) );
  NANDN U15745 ( .A(n14335), .B(n14336), .Z(n14334) );
  OR U15746 ( .A(n14337), .B(n14338), .Z(n14336) );
  NAND U15747 ( .A(n14338), .B(n14337), .Z(n14333) );
  XOR U15748 ( .A(n1473), .B(n1472), .Z(\A1[349] ) );
  XOR U15749 ( .A(n14321), .B(n14339), .Z(n1472) );
  XNOR U15750 ( .A(n14320), .B(n14318), .Z(n14339) );
  AND U15751 ( .A(n14340), .B(n14341), .Z(n14318) );
  NANDN U15752 ( .A(n14342), .B(n14343), .Z(n14341) );
  NANDN U15753 ( .A(n14344), .B(n14345), .Z(n14343) );
  AND U15754 ( .A(B[348]), .B(A[3]), .Z(n14320) );
  XNOR U15755 ( .A(n14310), .B(n14346), .Z(n14321) );
  XNOR U15756 ( .A(n14308), .B(n14311), .Z(n14346) );
  NAND U15757 ( .A(A[2]), .B(B[349]), .Z(n14311) );
  NANDN U15758 ( .A(n14347), .B(n14348), .Z(n14308) );
  AND U15759 ( .A(A[0]), .B(B[350]), .Z(n14348) );
  XOR U15760 ( .A(n14313), .B(n14349), .Z(n14310) );
  NAND U15761 ( .A(A[0]), .B(B[351]), .Z(n14349) );
  NAND U15762 ( .A(B[350]), .B(A[1]), .Z(n14313) );
  NAND U15763 ( .A(n14350), .B(n14351), .Z(n1473) );
  NANDN U15764 ( .A(n14352), .B(n14353), .Z(n14351) );
  OR U15765 ( .A(n14354), .B(n14355), .Z(n14353) );
  NAND U15766 ( .A(n14355), .B(n14354), .Z(n14350) );
  XOR U15767 ( .A(n1477), .B(n1476), .Z(\A1[348] ) );
  XOR U15768 ( .A(n14355), .B(n14356), .Z(n1476) );
  XNOR U15769 ( .A(n14354), .B(n14352), .Z(n14356) );
  AND U15770 ( .A(n14357), .B(n14358), .Z(n14352) );
  NANDN U15771 ( .A(n14359), .B(n14360), .Z(n14358) );
  NANDN U15772 ( .A(n14361), .B(n14362), .Z(n14360) );
  AND U15773 ( .A(B[347]), .B(A[3]), .Z(n14354) );
  XNOR U15774 ( .A(n14344), .B(n14363), .Z(n14355) );
  XNOR U15775 ( .A(n14342), .B(n14345), .Z(n14363) );
  NAND U15776 ( .A(A[2]), .B(B[348]), .Z(n14345) );
  NANDN U15777 ( .A(n14364), .B(n14365), .Z(n14342) );
  AND U15778 ( .A(A[0]), .B(B[349]), .Z(n14365) );
  XOR U15779 ( .A(n14347), .B(n14366), .Z(n14344) );
  NAND U15780 ( .A(A[0]), .B(B[350]), .Z(n14366) );
  NAND U15781 ( .A(B[349]), .B(A[1]), .Z(n14347) );
  NAND U15782 ( .A(n14367), .B(n14368), .Z(n1477) );
  NANDN U15783 ( .A(n14369), .B(n14370), .Z(n14368) );
  OR U15784 ( .A(n14371), .B(n14372), .Z(n14370) );
  NAND U15785 ( .A(n14372), .B(n14371), .Z(n14367) );
  XOR U15786 ( .A(n1479), .B(n1478), .Z(\A1[347] ) );
  XOR U15787 ( .A(n14372), .B(n14373), .Z(n1478) );
  XNOR U15788 ( .A(n14371), .B(n14369), .Z(n14373) );
  AND U15789 ( .A(n14374), .B(n14375), .Z(n14369) );
  NANDN U15790 ( .A(n14376), .B(n14377), .Z(n14375) );
  NANDN U15791 ( .A(n14378), .B(n14379), .Z(n14377) );
  AND U15792 ( .A(B[346]), .B(A[3]), .Z(n14371) );
  XNOR U15793 ( .A(n14361), .B(n14380), .Z(n14372) );
  XNOR U15794 ( .A(n14359), .B(n14362), .Z(n14380) );
  NAND U15795 ( .A(A[2]), .B(B[347]), .Z(n14362) );
  NANDN U15796 ( .A(n14381), .B(n14382), .Z(n14359) );
  AND U15797 ( .A(A[0]), .B(B[348]), .Z(n14382) );
  XOR U15798 ( .A(n14364), .B(n14383), .Z(n14361) );
  NAND U15799 ( .A(A[0]), .B(B[349]), .Z(n14383) );
  NAND U15800 ( .A(B[348]), .B(A[1]), .Z(n14364) );
  NAND U15801 ( .A(n14384), .B(n14385), .Z(n1479) );
  NANDN U15802 ( .A(n14386), .B(n14387), .Z(n14385) );
  OR U15803 ( .A(n14388), .B(n14389), .Z(n14387) );
  NAND U15804 ( .A(n14389), .B(n14388), .Z(n14384) );
  XOR U15805 ( .A(n1481), .B(n1480), .Z(\A1[346] ) );
  XOR U15806 ( .A(n14389), .B(n14390), .Z(n1480) );
  XNOR U15807 ( .A(n14388), .B(n14386), .Z(n14390) );
  AND U15808 ( .A(n14391), .B(n14392), .Z(n14386) );
  NANDN U15809 ( .A(n14393), .B(n14394), .Z(n14392) );
  NANDN U15810 ( .A(n14395), .B(n14396), .Z(n14394) );
  AND U15811 ( .A(B[345]), .B(A[3]), .Z(n14388) );
  XNOR U15812 ( .A(n14378), .B(n14397), .Z(n14389) );
  XNOR U15813 ( .A(n14376), .B(n14379), .Z(n14397) );
  NAND U15814 ( .A(A[2]), .B(B[346]), .Z(n14379) );
  NANDN U15815 ( .A(n14398), .B(n14399), .Z(n14376) );
  AND U15816 ( .A(A[0]), .B(B[347]), .Z(n14399) );
  XOR U15817 ( .A(n14381), .B(n14400), .Z(n14378) );
  NAND U15818 ( .A(A[0]), .B(B[348]), .Z(n14400) );
  NAND U15819 ( .A(B[347]), .B(A[1]), .Z(n14381) );
  NAND U15820 ( .A(n14401), .B(n14402), .Z(n1481) );
  NANDN U15821 ( .A(n14403), .B(n14404), .Z(n14402) );
  OR U15822 ( .A(n14405), .B(n14406), .Z(n14404) );
  NAND U15823 ( .A(n14406), .B(n14405), .Z(n14401) );
  XOR U15824 ( .A(n1483), .B(n1482), .Z(\A1[345] ) );
  XOR U15825 ( .A(n14406), .B(n14407), .Z(n1482) );
  XNOR U15826 ( .A(n14405), .B(n14403), .Z(n14407) );
  AND U15827 ( .A(n14408), .B(n14409), .Z(n14403) );
  NANDN U15828 ( .A(n14410), .B(n14411), .Z(n14409) );
  NANDN U15829 ( .A(n14412), .B(n14413), .Z(n14411) );
  AND U15830 ( .A(B[344]), .B(A[3]), .Z(n14405) );
  XNOR U15831 ( .A(n14395), .B(n14414), .Z(n14406) );
  XNOR U15832 ( .A(n14393), .B(n14396), .Z(n14414) );
  NAND U15833 ( .A(A[2]), .B(B[345]), .Z(n14396) );
  NANDN U15834 ( .A(n14415), .B(n14416), .Z(n14393) );
  AND U15835 ( .A(A[0]), .B(B[346]), .Z(n14416) );
  XOR U15836 ( .A(n14398), .B(n14417), .Z(n14395) );
  NAND U15837 ( .A(A[0]), .B(B[347]), .Z(n14417) );
  NAND U15838 ( .A(B[346]), .B(A[1]), .Z(n14398) );
  NAND U15839 ( .A(n14418), .B(n14419), .Z(n1483) );
  NANDN U15840 ( .A(n14420), .B(n14421), .Z(n14419) );
  OR U15841 ( .A(n14422), .B(n14423), .Z(n14421) );
  NAND U15842 ( .A(n14423), .B(n14422), .Z(n14418) );
  XOR U15843 ( .A(n1485), .B(n1484), .Z(\A1[344] ) );
  XOR U15844 ( .A(n14423), .B(n14424), .Z(n1484) );
  XNOR U15845 ( .A(n14422), .B(n14420), .Z(n14424) );
  AND U15846 ( .A(n14425), .B(n14426), .Z(n14420) );
  NANDN U15847 ( .A(n14427), .B(n14428), .Z(n14426) );
  NANDN U15848 ( .A(n14429), .B(n14430), .Z(n14428) );
  AND U15849 ( .A(B[343]), .B(A[3]), .Z(n14422) );
  XNOR U15850 ( .A(n14412), .B(n14431), .Z(n14423) );
  XNOR U15851 ( .A(n14410), .B(n14413), .Z(n14431) );
  NAND U15852 ( .A(A[2]), .B(B[344]), .Z(n14413) );
  NANDN U15853 ( .A(n14432), .B(n14433), .Z(n14410) );
  AND U15854 ( .A(A[0]), .B(B[345]), .Z(n14433) );
  XOR U15855 ( .A(n14415), .B(n14434), .Z(n14412) );
  NAND U15856 ( .A(A[0]), .B(B[346]), .Z(n14434) );
  NAND U15857 ( .A(B[345]), .B(A[1]), .Z(n14415) );
  NAND U15858 ( .A(n14435), .B(n14436), .Z(n1485) );
  NANDN U15859 ( .A(n14437), .B(n14438), .Z(n14436) );
  OR U15860 ( .A(n14439), .B(n14440), .Z(n14438) );
  NAND U15861 ( .A(n14440), .B(n14439), .Z(n14435) );
  XOR U15862 ( .A(n1487), .B(n1486), .Z(\A1[343] ) );
  XOR U15863 ( .A(n14440), .B(n14441), .Z(n1486) );
  XNOR U15864 ( .A(n14439), .B(n14437), .Z(n14441) );
  AND U15865 ( .A(n14442), .B(n14443), .Z(n14437) );
  NANDN U15866 ( .A(n14444), .B(n14445), .Z(n14443) );
  NANDN U15867 ( .A(n14446), .B(n14447), .Z(n14445) );
  AND U15868 ( .A(B[342]), .B(A[3]), .Z(n14439) );
  XNOR U15869 ( .A(n14429), .B(n14448), .Z(n14440) );
  XNOR U15870 ( .A(n14427), .B(n14430), .Z(n14448) );
  NAND U15871 ( .A(A[2]), .B(B[343]), .Z(n14430) );
  NANDN U15872 ( .A(n14449), .B(n14450), .Z(n14427) );
  AND U15873 ( .A(A[0]), .B(B[344]), .Z(n14450) );
  XOR U15874 ( .A(n14432), .B(n14451), .Z(n14429) );
  NAND U15875 ( .A(A[0]), .B(B[345]), .Z(n14451) );
  NAND U15876 ( .A(B[344]), .B(A[1]), .Z(n14432) );
  NAND U15877 ( .A(n14452), .B(n14453), .Z(n1487) );
  NANDN U15878 ( .A(n14454), .B(n14455), .Z(n14453) );
  OR U15879 ( .A(n14456), .B(n14457), .Z(n14455) );
  NAND U15880 ( .A(n14457), .B(n14456), .Z(n14452) );
  XOR U15881 ( .A(n1489), .B(n1488), .Z(\A1[342] ) );
  XOR U15882 ( .A(n14457), .B(n14458), .Z(n1488) );
  XNOR U15883 ( .A(n14456), .B(n14454), .Z(n14458) );
  AND U15884 ( .A(n14459), .B(n14460), .Z(n14454) );
  NANDN U15885 ( .A(n14461), .B(n14462), .Z(n14460) );
  NANDN U15886 ( .A(n14463), .B(n14464), .Z(n14462) );
  AND U15887 ( .A(B[341]), .B(A[3]), .Z(n14456) );
  XNOR U15888 ( .A(n14446), .B(n14465), .Z(n14457) );
  XNOR U15889 ( .A(n14444), .B(n14447), .Z(n14465) );
  NAND U15890 ( .A(A[2]), .B(B[342]), .Z(n14447) );
  NANDN U15891 ( .A(n14466), .B(n14467), .Z(n14444) );
  AND U15892 ( .A(A[0]), .B(B[343]), .Z(n14467) );
  XOR U15893 ( .A(n14449), .B(n14468), .Z(n14446) );
  NAND U15894 ( .A(A[0]), .B(B[344]), .Z(n14468) );
  NAND U15895 ( .A(B[343]), .B(A[1]), .Z(n14449) );
  NAND U15896 ( .A(n14469), .B(n14470), .Z(n1489) );
  NANDN U15897 ( .A(n14471), .B(n14472), .Z(n14470) );
  OR U15898 ( .A(n14473), .B(n14474), .Z(n14472) );
  NAND U15899 ( .A(n14474), .B(n14473), .Z(n14469) );
  XOR U15900 ( .A(n1491), .B(n1490), .Z(\A1[341] ) );
  XOR U15901 ( .A(n14474), .B(n14475), .Z(n1490) );
  XNOR U15902 ( .A(n14473), .B(n14471), .Z(n14475) );
  AND U15903 ( .A(n14476), .B(n14477), .Z(n14471) );
  NANDN U15904 ( .A(n14478), .B(n14479), .Z(n14477) );
  NANDN U15905 ( .A(n14480), .B(n14481), .Z(n14479) );
  AND U15906 ( .A(B[340]), .B(A[3]), .Z(n14473) );
  XNOR U15907 ( .A(n14463), .B(n14482), .Z(n14474) );
  XNOR U15908 ( .A(n14461), .B(n14464), .Z(n14482) );
  NAND U15909 ( .A(A[2]), .B(B[341]), .Z(n14464) );
  NANDN U15910 ( .A(n14483), .B(n14484), .Z(n14461) );
  AND U15911 ( .A(A[0]), .B(B[342]), .Z(n14484) );
  XOR U15912 ( .A(n14466), .B(n14485), .Z(n14463) );
  NAND U15913 ( .A(A[0]), .B(B[343]), .Z(n14485) );
  NAND U15914 ( .A(B[342]), .B(A[1]), .Z(n14466) );
  NAND U15915 ( .A(n14486), .B(n14487), .Z(n1491) );
  NANDN U15916 ( .A(n14488), .B(n14489), .Z(n14487) );
  OR U15917 ( .A(n14490), .B(n14491), .Z(n14489) );
  NAND U15918 ( .A(n14491), .B(n14490), .Z(n14486) );
  XOR U15919 ( .A(n1493), .B(n1492), .Z(\A1[340] ) );
  XOR U15920 ( .A(n14491), .B(n14492), .Z(n1492) );
  XNOR U15921 ( .A(n14490), .B(n14488), .Z(n14492) );
  AND U15922 ( .A(n14493), .B(n14494), .Z(n14488) );
  NANDN U15923 ( .A(n14495), .B(n14496), .Z(n14494) );
  NANDN U15924 ( .A(n14497), .B(n14498), .Z(n14496) );
  AND U15925 ( .A(B[339]), .B(A[3]), .Z(n14490) );
  XNOR U15926 ( .A(n14480), .B(n14499), .Z(n14491) );
  XNOR U15927 ( .A(n14478), .B(n14481), .Z(n14499) );
  NAND U15928 ( .A(A[2]), .B(B[340]), .Z(n14481) );
  NANDN U15929 ( .A(n14500), .B(n14501), .Z(n14478) );
  AND U15930 ( .A(A[0]), .B(B[341]), .Z(n14501) );
  XOR U15931 ( .A(n14483), .B(n14502), .Z(n14480) );
  NAND U15932 ( .A(A[0]), .B(B[342]), .Z(n14502) );
  NAND U15933 ( .A(B[341]), .B(A[1]), .Z(n14483) );
  NAND U15934 ( .A(n14503), .B(n14504), .Z(n1493) );
  NANDN U15935 ( .A(n14505), .B(n14506), .Z(n14504) );
  OR U15936 ( .A(n14507), .B(n14508), .Z(n14506) );
  NAND U15937 ( .A(n14508), .B(n14507), .Z(n14503) );
  XOR U15938 ( .A(n1475), .B(n1474), .Z(\A1[33] ) );
  XOR U15939 ( .A(n14338), .B(n14509), .Z(n1474) );
  XNOR U15940 ( .A(n14337), .B(n14335), .Z(n14509) );
  AND U15941 ( .A(n14510), .B(n14511), .Z(n14335) );
  NANDN U15942 ( .A(n14512), .B(n14513), .Z(n14511) );
  NANDN U15943 ( .A(n14514), .B(n14515), .Z(n14513) );
  AND U15944 ( .A(B[32]), .B(A[3]), .Z(n14337) );
  XNOR U15945 ( .A(n14327), .B(n14516), .Z(n14338) );
  XNOR U15946 ( .A(n14325), .B(n14328), .Z(n14516) );
  NAND U15947 ( .A(A[2]), .B(B[33]), .Z(n14328) );
  NANDN U15948 ( .A(n14517), .B(n14518), .Z(n14325) );
  AND U15949 ( .A(A[0]), .B(B[34]), .Z(n14518) );
  XOR U15950 ( .A(n14330), .B(n14519), .Z(n14327) );
  NAND U15951 ( .A(A[0]), .B(B[35]), .Z(n14519) );
  NAND U15952 ( .A(B[34]), .B(A[1]), .Z(n14330) );
  NAND U15953 ( .A(n14520), .B(n14521), .Z(n1475) );
  NANDN U15954 ( .A(n14522), .B(n14523), .Z(n14521) );
  OR U15955 ( .A(n14524), .B(n14525), .Z(n14523) );
  NAND U15956 ( .A(n14525), .B(n14524), .Z(n14520) );
  XOR U15957 ( .A(n1495), .B(n1494), .Z(\A1[339] ) );
  XOR U15958 ( .A(n14508), .B(n14526), .Z(n1494) );
  XNOR U15959 ( .A(n14507), .B(n14505), .Z(n14526) );
  AND U15960 ( .A(n14527), .B(n14528), .Z(n14505) );
  NANDN U15961 ( .A(n14529), .B(n14530), .Z(n14528) );
  NANDN U15962 ( .A(n14531), .B(n14532), .Z(n14530) );
  AND U15963 ( .A(B[338]), .B(A[3]), .Z(n14507) );
  XNOR U15964 ( .A(n14497), .B(n14533), .Z(n14508) );
  XNOR U15965 ( .A(n14495), .B(n14498), .Z(n14533) );
  NAND U15966 ( .A(A[2]), .B(B[339]), .Z(n14498) );
  NANDN U15967 ( .A(n14534), .B(n14535), .Z(n14495) );
  AND U15968 ( .A(A[0]), .B(B[340]), .Z(n14535) );
  XOR U15969 ( .A(n14500), .B(n14536), .Z(n14497) );
  NAND U15970 ( .A(A[0]), .B(B[341]), .Z(n14536) );
  NAND U15971 ( .A(B[340]), .B(A[1]), .Z(n14500) );
  NAND U15972 ( .A(n14537), .B(n14538), .Z(n1495) );
  NANDN U15973 ( .A(n14539), .B(n14540), .Z(n14538) );
  OR U15974 ( .A(n14541), .B(n14542), .Z(n14540) );
  NAND U15975 ( .A(n14542), .B(n14541), .Z(n14537) );
  XOR U15976 ( .A(n1499), .B(n1498), .Z(\A1[338] ) );
  XOR U15977 ( .A(n14542), .B(n14543), .Z(n1498) );
  XNOR U15978 ( .A(n14541), .B(n14539), .Z(n14543) );
  AND U15979 ( .A(n14544), .B(n14545), .Z(n14539) );
  NANDN U15980 ( .A(n14546), .B(n14547), .Z(n14545) );
  NANDN U15981 ( .A(n14548), .B(n14549), .Z(n14547) );
  AND U15982 ( .A(B[337]), .B(A[3]), .Z(n14541) );
  XNOR U15983 ( .A(n14531), .B(n14550), .Z(n14542) );
  XNOR U15984 ( .A(n14529), .B(n14532), .Z(n14550) );
  NAND U15985 ( .A(A[2]), .B(B[338]), .Z(n14532) );
  NANDN U15986 ( .A(n14551), .B(n14552), .Z(n14529) );
  AND U15987 ( .A(A[0]), .B(B[339]), .Z(n14552) );
  XOR U15988 ( .A(n14534), .B(n14553), .Z(n14531) );
  NAND U15989 ( .A(A[0]), .B(B[340]), .Z(n14553) );
  NAND U15990 ( .A(B[339]), .B(A[1]), .Z(n14534) );
  NAND U15991 ( .A(n14554), .B(n14555), .Z(n1499) );
  NANDN U15992 ( .A(n14556), .B(n14557), .Z(n14555) );
  OR U15993 ( .A(n14558), .B(n14559), .Z(n14557) );
  NAND U15994 ( .A(n14559), .B(n14558), .Z(n14554) );
  XOR U15995 ( .A(n1501), .B(n1500), .Z(\A1[337] ) );
  XOR U15996 ( .A(n14559), .B(n14560), .Z(n1500) );
  XNOR U15997 ( .A(n14558), .B(n14556), .Z(n14560) );
  AND U15998 ( .A(n14561), .B(n14562), .Z(n14556) );
  NANDN U15999 ( .A(n14563), .B(n14564), .Z(n14562) );
  NANDN U16000 ( .A(n14565), .B(n14566), .Z(n14564) );
  AND U16001 ( .A(B[336]), .B(A[3]), .Z(n14558) );
  XNOR U16002 ( .A(n14548), .B(n14567), .Z(n14559) );
  XNOR U16003 ( .A(n14546), .B(n14549), .Z(n14567) );
  NAND U16004 ( .A(A[2]), .B(B[337]), .Z(n14549) );
  NANDN U16005 ( .A(n14568), .B(n14569), .Z(n14546) );
  AND U16006 ( .A(A[0]), .B(B[338]), .Z(n14569) );
  XOR U16007 ( .A(n14551), .B(n14570), .Z(n14548) );
  NAND U16008 ( .A(A[0]), .B(B[339]), .Z(n14570) );
  NAND U16009 ( .A(B[338]), .B(A[1]), .Z(n14551) );
  NAND U16010 ( .A(n14571), .B(n14572), .Z(n1501) );
  NANDN U16011 ( .A(n14573), .B(n14574), .Z(n14572) );
  OR U16012 ( .A(n14575), .B(n14576), .Z(n14574) );
  NAND U16013 ( .A(n14576), .B(n14575), .Z(n14571) );
  XOR U16014 ( .A(n1503), .B(n1502), .Z(\A1[336] ) );
  XOR U16015 ( .A(n14576), .B(n14577), .Z(n1502) );
  XNOR U16016 ( .A(n14575), .B(n14573), .Z(n14577) );
  AND U16017 ( .A(n14578), .B(n14579), .Z(n14573) );
  NANDN U16018 ( .A(n14580), .B(n14581), .Z(n14579) );
  NANDN U16019 ( .A(n14582), .B(n14583), .Z(n14581) );
  AND U16020 ( .A(B[335]), .B(A[3]), .Z(n14575) );
  XNOR U16021 ( .A(n14565), .B(n14584), .Z(n14576) );
  XNOR U16022 ( .A(n14563), .B(n14566), .Z(n14584) );
  NAND U16023 ( .A(A[2]), .B(B[336]), .Z(n14566) );
  NANDN U16024 ( .A(n14585), .B(n14586), .Z(n14563) );
  AND U16025 ( .A(A[0]), .B(B[337]), .Z(n14586) );
  XOR U16026 ( .A(n14568), .B(n14587), .Z(n14565) );
  NAND U16027 ( .A(A[0]), .B(B[338]), .Z(n14587) );
  NAND U16028 ( .A(B[337]), .B(A[1]), .Z(n14568) );
  NAND U16029 ( .A(n14588), .B(n14589), .Z(n1503) );
  NANDN U16030 ( .A(n14590), .B(n14591), .Z(n14589) );
  OR U16031 ( .A(n14592), .B(n14593), .Z(n14591) );
  NAND U16032 ( .A(n14593), .B(n14592), .Z(n14588) );
  XOR U16033 ( .A(n1505), .B(n1504), .Z(\A1[335] ) );
  XOR U16034 ( .A(n14593), .B(n14594), .Z(n1504) );
  XNOR U16035 ( .A(n14592), .B(n14590), .Z(n14594) );
  AND U16036 ( .A(n14595), .B(n14596), .Z(n14590) );
  NANDN U16037 ( .A(n14597), .B(n14598), .Z(n14596) );
  NANDN U16038 ( .A(n14599), .B(n14600), .Z(n14598) );
  AND U16039 ( .A(B[334]), .B(A[3]), .Z(n14592) );
  XNOR U16040 ( .A(n14582), .B(n14601), .Z(n14593) );
  XNOR U16041 ( .A(n14580), .B(n14583), .Z(n14601) );
  NAND U16042 ( .A(A[2]), .B(B[335]), .Z(n14583) );
  NANDN U16043 ( .A(n14602), .B(n14603), .Z(n14580) );
  AND U16044 ( .A(A[0]), .B(B[336]), .Z(n14603) );
  XOR U16045 ( .A(n14585), .B(n14604), .Z(n14582) );
  NAND U16046 ( .A(A[0]), .B(B[337]), .Z(n14604) );
  NAND U16047 ( .A(B[336]), .B(A[1]), .Z(n14585) );
  NAND U16048 ( .A(n14605), .B(n14606), .Z(n1505) );
  NANDN U16049 ( .A(n14607), .B(n14608), .Z(n14606) );
  OR U16050 ( .A(n14609), .B(n14610), .Z(n14608) );
  NAND U16051 ( .A(n14610), .B(n14609), .Z(n14605) );
  XOR U16052 ( .A(n1507), .B(n1506), .Z(\A1[334] ) );
  XOR U16053 ( .A(n14610), .B(n14611), .Z(n1506) );
  XNOR U16054 ( .A(n14609), .B(n14607), .Z(n14611) );
  AND U16055 ( .A(n14612), .B(n14613), .Z(n14607) );
  NANDN U16056 ( .A(n14614), .B(n14615), .Z(n14613) );
  NANDN U16057 ( .A(n14616), .B(n14617), .Z(n14615) );
  AND U16058 ( .A(B[333]), .B(A[3]), .Z(n14609) );
  XNOR U16059 ( .A(n14599), .B(n14618), .Z(n14610) );
  XNOR U16060 ( .A(n14597), .B(n14600), .Z(n14618) );
  NAND U16061 ( .A(A[2]), .B(B[334]), .Z(n14600) );
  NANDN U16062 ( .A(n14619), .B(n14620), .Z(n14597) );
  AND U16063 ( .A(A[0]), .B(B[335]), .Z(n14620) );
  XOR U16064 ( .A(n14602), .B(n14621), .Z(n14599) );
  NAND U16065 ( .A(A[0]), .B(B[336]), .Z(n14621) );
  NAND U16066 ( .A(B[335]), .B(A[1]), .Z(n14602) );
  NAND U16067 ( .A(n14622), .B(n14623), .Z(n1507) );
  NANDN U16068 ( .A(n14624), .B(n14625), .Z(n14623) );
  OR U16069 ( .A(n14626), .B(n14627), .Z(n14625) );
  NAND U16070 ( .A(n14627), .B(n14626), .Z(n14622) );
  XOR U16071 ( .A(n1509), .B(n1508), .Z(\A1[333] ) );
  XOR U16072 ( .A(n14627), .B(n14628), .Z(n1508) );
  XNOR U16073 ( .A(n14626), .B(n14624), .Z(n14628) );
  AND U16074 ( .A(n14629), .B(n14630), .Z(n14624) );
  NANDN U16075 ( .A(n14631), .B(n14632), .Z(n14630) );
  NANDN U16076 ( .A(n14633), .B(n14634), .Z(n14632) );
  AND U16077 ( .A(B[332]), .B(A[3]), .Z(n14626) );
  XNOR U16078 ( .A(n14616), .B(n14635), .Z(n14627) );
  XNOR U16079 ( .A(n14614), .B(n14617), .Z(n14635) );
  NAND U16080 ( .A(A[2]), .B(B[333]), .Z(n14617) );
  NANDN U16081 ( .A(n14636), .B(n14637), .Z(n14614) );
  AND U16082 ( .A(A[0]), .B(B[334]), .Z(n14637) );
  XOR U16083 ( .A(n14619), .B(n14638), .Z(n14616) );
  NAND U16084 ( .A(A[0]), .B(B[335]), .Z(n14638) );
  NAND U16085 ( .A(B[334]), .B(A[1]), .Z(n14619) );
  NAND U16086 ( .A(n14639), .B(n14640), .Z(n1509) );
  NANDN U16087 ( .A(n14641), .B(n14642), .Z(n14640) );
  OR U16088 ( .A(n14643), .B(n14644), .Z(n14642) );
  NAND U16089 ( .A(n14644), .B(n14643), .Z(n14639) );
  XOR U16090 ( .A(n1511), .B(n1510), .Z(\A1[332] ) );
  XOR U16091 ( .A(n14644), .B(n14645), .Z(n1510) );
  XNOR U16092 ( .A(n14643), .B(n14641), .Z(n14645) );
  AND U16093 ( .A(n14646), .B(n14647), .Z(n14641) );
  NANDN U16094 ( .A(n14648), .B(n14649), .Z(n14647) );
  NANDN U16095 ( .A(n14650), .B(n14651), .Z(n14649) );
  AND U16096 ( .A(B[331]), .B(A[3]), .Z(n14643) );
  XNOR U16097 ( .A(n14633), .B(n14652), .Z(n14644) );
  XNOR U16098 ( .A(n14631), .B(n14634), .Z(n14652) );
  NAND U16099 ( .A(A[2]), .B(B[332]), .Z(n14634) );
  NANDN U16100 ( .A(n14653), .B(n14654), .Z(n14631) );
  AND U16101 ( .A(A[0]), .B(B[333]), .Z(n14654) );
  XOR U16102 ( .A(n14636), .B(n14655), .Z(n14633) );
  NAND U16103 ( .A(A[0]), .B(B[334]), .Z(n14655) );
  NAND U16104 ( .A(B[333]), .B(A[1]), .Z(n14636) );
  NAND U16105 ( .A(n14656), .B(n14657), .Z(n1511) );
  NANDN U16106 ( .A(n14658), .B(n14659), .Z(n14657) );
  OR U16107 ( .A(n14660), .B(n14661), .Z(n14659) );
  NAND U16108 ( .A(n14661), .B(n14660), .Z(n14656) );
  XOR U16109 ( .A(n1513), .B(n1512), .Z(\A1[331] ) );
  XOR U16110 ( .A(n14661), .B(n14662), .Z(n1512) );
  XNOR U16111 ( .A(n14660), .B(n14658), .Z(n14662) );
  AND U16112 ( .A(n14663), .B(n14664), .Z(n14658) );
  NANDN U16113 ( .A(n14665), .B(n14666), .Z(n14664) );
  NANDN U16114 ( .A(n14667), .B(n14668), .Z(n14666) );
  AND U16115 ( .A(B[330]), .B(A[3]), .Z(n14660) );
  XNOR U16116 ( .A(n14650), .B(n14669), .Z(n14661) );
  XNOR U16117 ( .A(n14648), .B(n14651), .Z(n14669) );
  NAND U16118 ( .A(A[2]), .B(B[331]), .Z(n14651) );
  NANDN U16119 ( .A(n14670), .B(n14671), .Z(n14648) );
  AND U16120 ( .A(A[0]), .B(B[332]), .Z(n14671) );
  XOR U16121 ( .A(n14653), .B(n14672), .Z(n14650) );
  NAND U16122 ( .A(A[0]), .B(B[333]), .Z(n14672) );
  NAND U16123 ( .A(B[332]), .B(A[1]), .Z(n14653) );
  NAND U16124 ( .A(n14673), .B(n14674), .Z(n1513) );
  NANDN U16125 ( .A(n14675), .B(n14676), .Z(n14674) );
  OR U16126 ( .A(n14677), .B(n14678), .Z(n14676) );
  NAND U16127 ( .A(n14678), .B(n14677), .Z(n14673) );
  XOR U16128 ( .A(n1515), .B(n1514), .Z(\A1[330] ) );
  XOR U16129 ( .A(n14678), .B(n14679), .Z(n1514) );
  XNOR U16130 ( .A(n14677), .B(n14675), .Z(n14679) );
  AND U16131 ( .A(n14680), .B(n14681), .Z(n14675) );
  NANDN U16132 ( .A(n14682), .B(n14683), .Z(n14681) );
  NANDN U16133 ( .A(n14684), .B(n14685), .Z(n14683) );
  AND U16134 ( .A(B[329]), .B(A[3]), .Z(n14677) );
  XNOR U16135 ( .A(n14667), .B(n14686), .Z(n14678) );
  XNOR U16136 ( .A(n14665), .B(n14668), .Z(n14686) );
  NAND U16137 ( .A(A[2]), .B(B[330]), .Z(n14668) );
  NANDN U16138 ( .A(n14687), .B(n14688), .Z(n14665) );
  AND U16139 ( .A(A[0]), .B(B[331]), .Z(n14688) );
  XOR U16140 ( .A(n14670), .B(n14689), .Z(n14667) );
  NAND U16141 ( .A(A[0]), .B(B[332]), .Z(n14689) );
  NAND U16142 ( .A(B[331]), .B(A[1]), .Z(n14670) );
  NAND U16143 ( .A(n14690), .B(n14691), .Z(n1515) );
  NANDN U16144 ( .A(n14692), .B(n14693), .Z(n14691) );
  OR U16145 ( .A(n14694), .B(n14695), .Z(n14693) );
  NAND U16146 ( .A(n14695), .B(n14694), .Z(n14690) );
  XOR U16147 ( .A(n1497), .B(n1496), .Z(\A1[32] ) );
  XOR U16148 ( .A(n14525), .B(n14696), .Z(n1496) );
  XNOR U16149 ( .A(n14524), .B(n14522), .Z(n14696) );
  AND U16150 ( .A(n14697), .B(n14698), .Z(n14522) );
  NANDN U16151 ( .A(n14699), .B(n14700), .Z(n14698) );
  NANDN U16152 ( .A(n14701), .B(n14702), .Z(n14700) );
  AND U16153 ( .A(B[31]), .B(A[3]), .Z(n14524) );
  XNOR U16154 ( .A(n14514), .B(n14703), .Z(n14525) );
  XNOR U16155 ( .A(n14512), .B(n14515), .Z(n14703) );
  NAND U16156 ( .A(A[2]), .B(B[32]), .Z(n14515) );
  NANDN U16157 ( .A(n14704), .B(n14705), .Z(n14512) );
  AND U16158 ( .A(A[0]), .B(B[33]), .Z(n14705) );
  XOR U16159 ( .A(n14517), .B(n14706), .Z(n14514) );
  NAND U16160 ( .A(A[0]), .B(B[34]), .Z(n14706) );
  NAND U16161 ( .A(B[33]), .B(A[1]), .Z(n14517) );
  NAND U16162 ( .A(n14707), .B(n14708), .Z(n1497) );
  NANDN U16163 ( .A(n14709), .B(n14710), .Z(n14708) );
  OR U16164 ( .A(n14711), .B(n14712), .Z(n14710) );
  NAND U16165 ( .A(n14712), .B(n14711), .Z(n14707) );
  XOR U16166 ( .A(n1517), .B(n1516), .Z(\A1[329] ) );
  XOR U16167 ( .A(n14695), .B(n14713), .Z(n1516) );
  XNOR U16168 ( .A(n14694), .B(n14692), .Z(n14713) );
  AND U16169 ( .A(n14714), .B(n14715), .Z(n14692) );
  NANDN U16170 ( .A(n14716), .B(n14717), .Z(n14715) );
  NANDN U16171 ( .A(n14718), .B(n14719), .Z(n14717) );
  AND U16172 ( .A(B[328]), .B(A[3]), .Z(n14694) );
  XNOR U16173 ( .A(n14684), .B(n14720), .Z(n14695) );
  XNOR U16174 ( .A(n14682), .B(n14685), .Z(n14720) );
  NAND U16175 ( .A(A[2]), .B(B[329]), .Z(n14685) );
  NANDN U16176 ( .A(n14721), .B(n14722), .Z(n14682) );
  AND U16177 ( .A(A[0]), .B(B[330]), .Z(n14722) );
  XOR U16178 ( .A(n14687), .B(n14723), .Z(n14684) );
  NAND U16179 ( .A(A[0]), .B(B[331]), .Z(n14723) );
  NAND U16180 ( .A(B[330]), .B(A[1]), .Z(n14687) );
  NAND U16181 ( .A(n14724), .B(n14725), .Z(n1517) );
  NANDN U16182 ( .A(n14726), .B(n14727), .Z(n14725) );
  OR U16183 ( .A(n14728), .B(n14729), .Z(n14727) );
  NAND U16184 ( .A(n14729), .B(n14728), .Z(n14724) );
  XOR U16185 ( .A(n1521), .B(n1520), .Z(\A1[328] ) );
  XOR U16186 ( .A(n14729), .B(n14730), .Z(n1520) );
  XNOR U16187 ( .A(n14728), .B(n14726), .Z(n14730) );
  AND U16188 ( .A(n14731), .B(n14732), .Z(n14726) );
  NANDN U16189 ( .A(n14733), .B(n14734), .Z(n14732) );
  NANDN U16190 ( .A(n14735), .B(n14736), .Z(n14734) );
  AND U16191 ( .A(B[327]), .B(A[3]), .Z(n14728) );
  XNOR U16192 ( .A(n14718), .B(n14737), .Z(n14729) );
  XNOR U16193 ( .A(n14716), .B(n14719), .Z(n14737) );
  NAND U16194 ( .A(A[2]), .B(B[328]), .Z(n14719) );
  NANDN U16195 ( .A(n14738), .B(n14739), .Z(n14716) );
  AND U16196 ( .A(A[0]), .B(B[329]), .Z(n14739) );
  XOR U16197 ( .A(n14721), .B(n14740), .Z(n14718) );
  NAND U16198 ( .A(A[0]), .B(B[330]), .Z(n14740) );
  NAND U16199 ( .A(B[329]), .B(A[1]), .Z(n14721) );
  NAND U16200 ( .A(n14741), .B(n14742), .Z(n1521) );
  NANDN U16201 ( .A(n14743), .B(n14744), .Z(n14742) );
  OR U16202 ( .A(n14745), .B(n14746), .Z(n14744) );
  NAND U16203 ( .A(n14746), .B(n14745), .Z(n14741) );
  XOR U16204 ( .A(n1523), .B(n1522), .Z(\A1[327] ) );
  XOR U16205 ( .A(n14746), .B(n14747), .Z(n1522) );
  XNOR U16206 ( .A(n14745), .B(n14743), .Z(n14747) );
  AND U16207 ( .A(n14748), .B(n14749), .Z(n14743) );
  NANDN U16208 ( .A(n14750), .B(n14751), .Z(n14749) );
  NANDN U16209 ( .A(n14752), .B(n14753), .Z(n14751) );
  AND U16210 ( .A(B[326]), .B(A[3]), .Z(n14745) );
  XNOR U16211 ( .A(n14735), .B(n14754), .Z(n14746) );
  XNOR U16212 ( .A(n14733), .B(n14736), .Z(n14754) );
  NAND U16213 ( .A(A[2]), .B(B[327]), .Z(n14736) );
  NANDN U16214 ( .A(n14755), .B(n14756), .Z(n14733) );
  AND U16215 ( .A(A[0]), .B(B[328]), .Z(n14756) );
  XOR U16216 ( .A(n14738), .B(n14757), .Z(n14735) );
  NAND U16217 ( .A(A[0]), .B(B[329]), .Z(n14757) );
  NAND U16218 ( .A(B[328]), .B(A[1]), .Z(n14738) );
  NAND U16219 ( .A(n14758), .B(n14759), .Z(n1523) );
  NANDN U16220 ( .A(n14760), .B(n14761), .Z(n14759) );
  OR U16221 ( .A(n14762), .B(n14763), .Z(n14761) );
  NAND U16222 ( .A(n14763), .B(n14762), .Z(n14758) );
  XOR U16223 ( .A(n1525), .B(n1524), .Z(\A1[326] ) );
  XOR U16224 ( .A(n14763), .B(n14764), .Z(n1524) );
  XNOR U16225 ( .A(n14762), .B(n14760), .Z(n14764) );
  AND U16226 ( .A(n14765), .B(n14766), .Z(n14760) );
  NANDN U16227 ( .A(n14767), .B(n14768), .Z(n14766) );
  NANDN U16228 ( .A(n14769), .B(n14770), .Z(n14768) );
  AND U16229 ( .A(B[325]), .B(A[3]), .Z(n14762) );
  XNOR U16230 ( .A(n14752), .B(n14771), .Z(n14763) );
  XNOR U16231 ( .A(n14750), .B(n14753), .Z(n14771) );
  NAND U16232 ( .A(A[2]), .B(B[326]), .Z(n14753) );
  NANDN U16233 ( .A(n14772), .B(n14773), .Z(n14750) );
  AND U16234 ( .A(A[0]), .B(B[327]), .Z(n14773) );
  XOR U16235 ( .A(n14755), .B(n14774), .Z(n14752) );
  NAND U16236 ( .A(A[0]), .B(B[328]), .Z(n14774) );
  NAND U16237 ( .A(B[327]), .B(A[1]), .Z(n14755) );
  NAND U16238 ( .A(n14775), .B(n14776), .Z(n1525) );
  NANDN U16239 ( .A(n14777), .B(n14778), .Z(n14776) );
  OR U16240 ( .A(n14779), .B(n14780), .Z(n14778) );
  NAND U16241 ( .A(n14780), .B(n14779), .Z(n14775) );
  XOR U16242 ( .A(n1527), .B(n1526), .Z(\A1[325] ) );
  XOR U16243 ( .A(n14780), .B(n14781), .Z(n1526) );
  XNOR U16244 ( .A(n14779), .B(n14777), .Z(n14781) );
  AND U16245 ( .A(n14782), .B(n14783), .Z(n14777) );
  NANDN U16246 ( .A(n14784), .B(n14785), .Z(n14783) );
  NANDN U16247 ( .A(n14786), .B(n14787), .Z(n14785) );
  AND U16248 ( .A(B[324]), .B(A[3]), .Z(n14779) );
  XNOR U16249 ( .A(n14769), .B(n14788), .Z(n14780) );
  XNOR U16250 ( .A(n14767), .B(n14770), .Z(n14788) );
  NAND U16251 ( .A(A[2]), .B(B[325]), .Z(n14770) );
  NANDN U16252 ( .A(n14789), .B(n14790), .Z(n14767) );
  AND U16253 ( .A(A[0]), .B(B[326]), .Z(n14790) );
  XOR U16254 ( .A(n14772), .B(n14791), .Z(n14769) );
  NAND U16255 ( .A(A[0]), .B(B[327]), .Z(n14791) );
  NAND U16256 ( .A(B[326]), .B(A[1]), .Z(n14772) );
  NAND U16257 ( .A(n14792), .B(n14793), .Z(n1527) );
  NANDN U16258 ( .A(n14794), .B(n14795), .Z(n14793) );
  OR U16259 ( .A(n14796), .B(n14797), .Z(n14795) );
  NAND U16260 ( .A(n14797), .B(n14796), .Z(n14792) );
  XOR U16261 ( .A(n1529), .B(n1528), .Z(\A1[324] ) );
  XOR U16262 ( .A(n14797), .B(n14798), .Z(n1528) );
  XNOR U16263 ( .A(n14796), .B(n14794), .Z(n14798) );
  AND U16264 ( .A(n14799), .B(n14800), .Z(n14794) );
  NANDN U16265 ( .A(n14801), .B(n14802), .Z(n14800) );
  NANDN U16266 ( .A(n14803), .B(n14804), .Z(n14802) );
  AND U16267 ( .A(B[323]), .B(A[3]), .Z(n14796) );
  XNOR U16268 ( .A(n14786), .B(n14805), .Z(n14797) );
  XNOR U16269 ( .A(n14784), .B(n14787), .Z(n14805) );
  NAND U16270 ( .A(A[2]), .B(B[324]), .Z(n14787) );
  NANDN U16271 ( .A(n14806), .B(n14807), .Z(n14784) );
  AND U16272 ( .A(A[0]), .B(B[325]), .Z(n14807) );
  XOR U16273 ( .A(n14789), .B(n14808), .Z(n14786) );
  NAND U16274 ( .A(A[0]), .B(B[326]), .Z(n14808) );
  NAND U16275 ( .A(B[325]), .B(A[1]), .Z(n14789) );
  NAND U16276 ( .A(n14809), .B(n14810), .Z(n1529) );
  NANDN U16277 ( .A(n14811), .B(n14812), .Z(n14810) );
  OR U16278 ( .A(n14813), .B(n14814), .Z(n14812) );
  NAND U16279 ( .A(n14814), .B(n14813), .Z(n14809) );
  XOR U16280 ( .A(n1531), .B(n1530), .Z(\A1[323] ) );
  XOR U16281 ( .A(n14814), .B(n14815), .Z(n1530) );
  XNOR U16282 ( .A(n14813), .B(n14811), .Z(n14815) );
  AND U16283 ( .A(n14816), .B(n14817), .Z(n14811) );
  NANDN U16284 ( .A(n14818), .B(n14819), .Z(n14817) );
  NANDN U16285 ( .A(n14820), .B(n14821), .Z(n14819) );
  AND U16286 ( .A(B[322]), .B(A[3]), .Z(n14813) );
  XNOR U16287 ( .A(n14803), .B(n14822), .Z(n14814) );
  XNOR U16288 ( .A(n14801), .B(n14804), .Z(n14822) );
  NAND U16289 ( .A(A[2]), .B(B[323]), .Z(n14804) );
  NANDN U16290 ( .A(n14823), .B(n14824), .Z(n14801) );
  AND U16291 ( .A(A[0]), .B(B[324]), .Z(n14824) );
  XOR U16292 ( .A(n14806), .B(n14825), .Z(n14803) );
  NAND U16293 ( .A(A[0]), .B(B[325]), .Z(n14825) );
  NAND U16294 ( .A(B[324]), .B(A[1]), .Z(n14806) );
  NAND U16295 ( .A(n14826), .B(n14827), .Z(n1531) );
  NANDN U16296 ( .A(n14828), .B(n14829), .Z(n14827) );
  OR U16297 ( .A(n14830), .B(n14831), .Z(n14829) );
  NAND U16298 ( .A(n14831), .B(n14830), .Z(n14826) );
  XOR U16299 ( .A(n1533), .B(n1532), .Z(\A1[322] ) );
  XOR U16300 ( .A(n14831), .B(n14832), .Z(n1532) );
  XNOR U16301 ( .A(n14830), .B(n14828), .Z(n14832) );
  AND U16302 ( .A(n14833), .B(n14834), .Z(n14828) );
  NANDN U16303 ( .A(n14835), .B(n14836), .Z(n14834) );
  NANDN U16304 ( .A(n14837), .B(n14838), .Z(n14836) );
  AND U16305 ( .A(B[321]), .B(A[3]), .Z(n14830) );
  XNOR U16306 ( .A(n14820), .B(n14839), .Z(n14831) );
  XNOR U16307 ( .A(n14818), .B(n14821), .Z(n14839) );
  NAND U16308 ( .A(A[2]), .B(B[322]), .Z(n14821) );
  NANDN U16309 ( .A(n14840), .B(n14841), .Z(n14818) );
  AND U16310 ( .A(A[0]), .B(B[323]), .Z(n14841) );
  XOR U16311 ( .A(n14823), .B(n14842), .Z(n14820) );
  NAND U16312 ( .A(A[0]), .B(B[324]), .Z(n14842) );
  NAND U16313 ( .A(B[323]), .B(A[1]), .Z(n14823) );
  NAND U16314 ( .A(n14843), .B(n14844), .Z(n1533) );
  NANDN U16315 ( .A(n14845), .B(n14846), .Z(n14844) );
  OR U16316 ( .A(n14847), .B(n14848), .Z(n14846) );
  NAND U16317 ( .A(n14848), .B(n14847), .Z(n14843) );
  XOR U16318 ( .A(n1535), .B(n1534), .Z(\A1[321] ) );
  XOR U16319 ( .A(n14848), .B(n14849), .Z(n1534) );
  XNOR U16320 ( .A(n14847), .B(n14845), .Z(n14849) );
  AND U16321 ( .A(n14850), .B(n14851), .Z(n14845) );
  NANDN U16322 ( .A(n14852), .B(n14853), .Z(n14851) );
  NANDN U16323 ( .A(n14854), .B(n14855), .Z(n14853) );
  AND U16324 ( .A(B[320]), .B(A[3]), .Z(n14847) );
  XNOR U16325 ( .A(n14837), .B(n14856), .Z(n14848) );
  XNOR U16326 ( .A(n14835), .B(n14838), .Z(n14856) );
  NAND U16327 ( .A(A[2]), .B(B[321]), .Z(n14838) );
  NANDN U16328 ( .A(n14857), .B(n14858), .Z(n14835) );
  AND U16329 ( .A(A[0]), .B(B[322]), .Z(n14858) );
  XOR U16330 ( .A(n14840), .B(n14859), .Z(n14837) );
  NAND U16331 ( .A(A[0]), .B(B[323]), .Z(n14859) );
  NAND U16332 ( .A(B[322]), .B(A[1]), .Z(n14840) );
  NAND U16333 ( .A(n14860), .B(n14861), .Z(n1535) );
  NANDN U16334 ( .A(n14862), .B(n14863), .Z(n14861) );
  OR U16335 ( .A(n14864), .B(n14865), .Z(n14863) );
  NAND U16336 ( .A(n14865), .B(n14864), .Z(n14860) );
  XOR U16337 ( .A(n1537), .B(n1536), .Z(\A1[320] ) );
  XOR U16338 ( .A(n14865), .B(n14866), .Z(n1536) );
  XNOR U16339 ( .A(n14864), .B(n14862), .Z(n14866) );
  AND U16340 ( .A(n14867), .B(n14868), .Z(n14862) );
  NANDN U16341 ( .A(n14869), .B(n14870), .Z(n14868) );
  NANDN U16342 ( .A(n14871), .B(n14872), .Z(n14870) );
  AND U16343 ( .A(B[319]), .B(A[3]), .Z(n14864) );
  XNOR U16344 ( .A(n14854), .B(n14873), .Z(n14865) );
  XNOR U16345 ( .A(n14852), .B(n14855), .Z(n14873) );
  NAND U16346 ( .A(A[2]), .B(B[320]), .Z(n14855) );
  NANDN U16347 ( .A(n14874), .B(n14875), .Z(n14852) );
  AND U16348 ( .A(A[0]), .B(B[321]), .Z(n14875) );
  XOR U16349 ( .A(n14857), .B(n14876), .Z(n14854) );
  NAND U16350 ( .A(A[0]), .B(B[322]), .Z(n14876) );
  NAND U16351 ( .A(B[321]), .B(A[1]), .Z(n14857) );
  NAND U16352 ( .A(n14877), .B(n14878), .Z(n1537) );
  NANDN U16353 ( .A(n14879), .B(n14880), .Z(n14878) );
  OR U16354 ( .A(n14881), .B(n14882), .Z(n14880) );
  NAND U16355 ( .A(n14882), .B(n14881), .Z(n14877) );
  XOR U16356 ( .A(n1519), .B(n1518), .Z(\A1[31] ) );
  XOR U16357 ( .A(n14712), .B(n14883), .Z(n1518) );
  XNOR U16358 ( .A(n14711), .B(n14709), .Z(n14883) );
  AND U16359 ( .A(n14884), .B(n14885), .Z(n14709) );
  NANDN U16360 ( .A(n14886), .B(n14887), .Z(n14885) );
  NANDN U16361 ( .A(n14888), .B(n14889), .Z(n14887) );
  AND U16362 ( .A(B[30]), .B(A[3]), .Z(n14711) );
  XNOR U16363 ( .A(n14701), .B(n14890), .Z(n14712) );
  XNOR U16364 ( .A(n14699), .B(n14702), .Z(n14890) );
  NAND U16365 ( .A(A[2]), .B(B[31]), .Z(n14702) );
  NANDN U16366 ( .A(n14891), .B(n14892), .Z(n14699) );
  AND U16367 ( .A(A[0]), .B(B[32]), .Z(n14892) );
  XOR U16368 ( .A(n14704), .B(n14893), .Z(n14701) );
  NAND U16369 ( .A(A[0]), .B(B[33]), .Z(n14893) );
  NAND U16370 ( .A(B[32]), .B(A[1]), .Z(n14704) );
  NAND U16371 ( .A(n14894), .B(n14895), .Z(n1519) );
  NANDN U16372 ( .A(n14896), .B(n14897), .Z(n14895) );
  OR U16373 ( .A(n14898), .B(n14899), .Z(n14897) );
  NAND U16374 ( .A(n14899), .B(n14898), .Z(n14894) );
  XOR U16375 ( .A(n1539), .B(n1538), .Z(\A1[319] ) );
  XOR U16376 ( .A(n14882), .B(n14900), .Z(n1538) );
  XNOR U16377 ( .A(n14881), .B(n14879), .Z(n14900) );
  AND U16378 ( .A(n14901), .B(n14902), .Z(n14879) );
  NANDN U16379 ( .A(n14903), .B(n14904), .Z(n14902) );
  NANDN U16380 ( .A(n14905), .B(n14906), .Z(n14904) );
  AND U16381 ( .A(B[318]), .B(A[3]), .Z(n14881) );
  XNOR U16382 ( .A(n14871), .B(n14907), .Z(n14882) );
  XNOR U16383 ( .A(n14869), .B(n14872), .Z(n14907) );
  NAND U16384 ( .A(A[2]), .B(B[319]), .Z(n14872) );
  NANDN U16385 ( .A(n14908), .B(n14909), .Z(n14869) );
  AND U16386 ( .A(A[0]), .B(B[320]), .Z(n14909) );
  XOR U16387 ( .A(n14874), .B(n14910), .Z(n14871) );
  NAND U16388 ( .A(A[0]), .B(B[321]), .Z(n14910) );
  NAND U16389 ( .A(B[320]), .B(A[1]), .Z(n14874) );
  NAND U16390 ( .A(n14911), .B(n14912), .Z(n1539) );
  NANDN U16391 ( .A(n14913), .B(n14914), .Z(n14912) );
  OR U16392 ( .A(n14915), .B(n14916), .Z(n14914) );
  NAND U16393 ( .A(n14916), .B(n14915), .Z(n14911) );
  XOR U16394 ( .A(n1543), .B(n1542), .Z(\A1[318] ) );
  XOR U16395 ( .A(n14916), .B(n14917), .Z(n1542) );
  XNOR U16396 ( .A(n14915), .B(n14913), .Z(n14917) );
  AND U16397 ( .A(n14918), .B(n14919), .Z(n14913) );
  NANDN U16398 ( .A(n14920), .B(n14921), .Z(n14919) );
  NANDN U16399 ( .A(n14922), .B(n14923), .Z(n14921) );
  AND U16400 ( .A(B[317]), .B(A[3]), .Z(n14915) );
  XNOR U16401 ( .A(n14905), .B(n14924), .Z(n14916) );
  XNOR U16402 ( .A(n14903), .B(n14906), .Z(n14924) );
  NAND U16403 ( .A(A[2]), .B(B[318]), .Z(n14906) );
  NANDN U16404 ( .A(n14925), .B(n14926), .Z(n14903) );
  AND U16405 ( .A(A[0]), .B(B[319]), .Z(n14926) );
  XOR U16406 ( .A(n14908), .B(n14927), .Z(n14905) );
  NAND U16407 ( .A(A[0]), .B(B[320]), .Z(n14927) );
  NAND U16408 ( .A(B[319]), .B(A[1]), .Z(n14908) );
  NAND U16409 ( .A(n14928), .B(n14929), .Z(n1543) );
  NANDN U16410 ( .A(n14930), .B(n14931), .Z(n14929) );
  OR U16411 ( .A(n14932), .B(n14933), .Z(n14931) );
  NAND U16412 ( .A(n14933), .B(n14932), .Z(n14928) );
  XOR U16413 ( .A(n1545), .B(n1544), .Z(\A1[317] ) );
  XOR U16414 ( .A(n14933), .B(n14934), .Z(n1544) );
  XNOR U16415 ( .A(n14932), .B(n14930), .Z(n14934) );
  AND U16416 ( .A(n14935), .B(n14936), .Z(n14930) );
  NANDN U16417 ( .A(n14937), .B(n14938), .Z(n14936) );
  NANDN U16418 ( .A(n14939), .B(n14940), .Z(n14938) );
  AND U16419 ( .A(B[316]), .B(A[3]), .Z(n14932) );
  XNOR U16420 ( .A(n14922), .B(n14941), .Z(n14933) );
  XNOR U16421 ( .A(n14920), .B(n14923), .Z(n14941) );
  NAND U16422 ( .A(A[2]), .B(B[317]), .Z(n14923) );
  NANDN U16423 ( .A(n14942), .B(n14943), .Z(n14920) );
  AND U16424 ( .A(A[0]), .B(B[318]), .Z(n14943) );
  XOR U16425 ( .A(n14925), .B(n14944), .Z(n14922) );
  NAND U16426 ( .A(A[0]), .B(B[319]), .Z(n14944) );
  NAND U16427 ( .A(B[318]), .B(A[1]), .Z(n14925) );
  NAND U16428 ( .A(n14945), .B(n14946), .Z(n1545) );
  NANDN U16429 ( .A(n14947), .B(n14948), .Z(n14946) );
  OR U16430 ( .A(n14949), .B(n14950), .Z(n14948) );
  NAND U16431 ( .A(n14950), .B(n14949), .Z(n14945) );
  XOR U16432 ( .A(n1547), .B(n1546), .Z(\A1[316] ) );
  XOR U16433 ( .A(n14950), .B(n14951), .Z(n1546) );
  XNOR U16434 ( .A(n14949), .B(n14947), .Z(n14951) );
  AND U16435 ( .A(n14952), .B(n14953), .Z(n14947) );
  NANDN U16436 ( .A(n14954), .B(n14955), .Z(n14953) );
  NANDN U16437 ( .A(n14956), .B(n14957), .Z(n14955) );
  AND U16438 ( .A(B[315]), .B(A[3]), .Z(n14949) );
  XNOR U16439 ( .A(n14939), .B(n14958), .Z(n14950) );
  XNOR U16440 ( .A(n14937), .B(n14940), .Z(n14958) );
  NAND U16441 ( .A(A[2]), .B(B[316]), .Z(n14940) );
  NANDN U16442 ( .A(n14959), .B(n14960), .Z(n14937) );
  AND U16443 ( .A(A[0]), .B(B[317]), .Z(n14960) );
  XOR U16444 ( .A(n14942), .B(n14961), .Z(n14939) );
  NAND U16445 ( .A(A[0]), .B(B[318]), .Z(n14961) );
  NAND U16446 ( .A(B[317]), .B(A[1]), .Z(n14942) );
  NAND U16447 ( .A(n14962), .B(n14963), .Z(n1547) );
  NANDN U16448 ( .A(n14964), .B(n14965), .Z(n14963) );
  OR U16449 ( .A(n14966), .B(n14967), .Z(n14965) );
  NAND U16450 ( .A(n14967), .B(n14966), .Z(n14962) );
  XOR U16451 ( .A(n1549), .B(n1548), .Z(\A1[315] ) );
  XOR U16452 ( .A(n14967), .B(n14968), .Z(n1548) );
  XNOR U16453 ( .A(n14966), .B(n14964), .Z(n14968) );
  AND U16454 ( .A(n14969), .B(n14970), .Z(n14964) );
  NANDN U16455 ( .A(n14971), .B(n14972), .Z(n14970) );
  NANDN U16456 ( .A(n14973), .B(n14974), .Z(n14972) );
  AND U16457 ( .A(B[314]), .B(A[3]), .Z(n14966) );
  XNOR U16458 ( .A(n14956), .B(n14975), .Z(n14967) );
  XNOR U16459 ( .A(n14954), .B(n14957), .Z(n14975) );
  NAND U16460 ( .A(A[2]), .B(B[315]), .Z(n14957) );
  NANDN U16461 ( .A(n14976), .B(n14977), .Z(n14954) );
  AND U16462 ( .A(A[0]), .B(B[316]), .Z(n14977) );
  XOR U16463 ( .A(n14959), .B(n14978), .Z(n14956) );
  NAND U16464 ( .A(A[0]), .B(B[317]), .Z(n14978) );
  NAND U16465 ( .A(B[316]), .B(A[1]), .Z(n14959) );
  NAND U16466 ( .A(n14979), .B(n14980), .Z(n1549) );
  NANDN U16467 ( .A(n14981), .B(n14982), .Z(n14980) );
  OR U16468 ( .A(n14983), .B(n14984), .Z(n14982) );
  NAND U16469 ( .A(n14984), .B(n14983), .Z(n14979) );
  XOR U16470 ( .A(n1551), .B(n1550), .Z(\A1[314] ) );
  XOR U16471 ( .A(n14984), .B(n14985), .Z(n1550) );
  XNOR U16472 ( .A(n14983), .B(n14981), .Z(n14985) );
  AND U16473 ( .A(n14986), .B(n14987), .Z(n14981) );
  NANDN U16474 ( .A(n14988), .B(n14989), .Z(n14987) );
  NANDN U16475 ( .A(n14990), .B(n14991), .Z(n14989) );
  AND U16476 ( .A(B[313]), .B(A[3]), .Z(n14983) );
  XNOR U16477 ( .A(n14973), .B(n14992), .Z(n14984) );
  XNOR U16478 ( .A(n14971), .B(n14974), .Z(n14992) );
  NAND U16479 ( .A(A[2]), .B(B[314]), .Z(n14974) );
  NANDN U16480 ( .A(n14993), .B(n14994), .Z(n14971) );
  AND U16481 ( .A(A[0]), .B(B[315]), .Z(n14994) );
  XOR U16482 ( .A(n14976), .B(n14995), .Z(n14973) );
  NAND U16483 ( .A(A[0]), .B(B[316]), .Z(n14995) );
  NAND U16484 ( .A(B[315]), .B(A[1]), .Z(n14976) );
  NAND U16485 ( .A(n14996), .B(n14997), .Z(n1551) );
  NANDN U16486 ( .A(n14998), .B(n14999), .Z(n14997) );
  OR U16487 ( .A(n15000), .B(n15001), .Z(n14999) );
  NAND U16488 ( .A(n15001), .B(n15000), .Z(n14996) );
  XOR U16489 ( .A(n1553), .B(n1552), .Z(\A1[313] ) );
  XOR U16490 ( .A(n15001), .B(n15002), .Z(n1552) );
  XNOR U16491 ( .A(n15000), .B(n14998), .Z(n15002) );
  AND U16492 ( .A(n15003), .B(n15004), .Z(n14998) );
  NANDN U16493 ( .A(n15005), .B(n15006), .Z(n15004) );
  NANDN U16494 ( .A(n15007), .B(n15008), .Z(n15006) );
  AND U16495 ( .A(B[312]), .B(A[3]), .Z(n15000) );
  XNOR U16496 ( .A(n14990), .B(n15009), .Z(n15001) );
  XNOR U16497 ( .A(n14988), .B(n14991), .Z(n15009) );
  NAND U16498 ( .A(A[2]), .B(B[313]), .Z(n14991) );
  NANDN U16499 ( .A(n15010), .B(n15011), .Z(n14988) );
  AND U16500 ( .A(A[0]), .B(B[314]), .Z(n15011) );
  XOR U16501 ( .A(n14993), .B(n15012), .Z(n14990) );
  NAND U16502 ( .A(A[0]), .B(B[315]), .Z(n15012) );
  NAND U16503 ( .A(B[314]), .B(A[1]), .Z(n14993) );
  NAND U16504 ( .A(n15013), .B(n15014), .Z(n1553) );
  NANDN U16505 ( .A(n15015), .B(n15016), .Z(n15014) );
  OR U16506 ( .A(n15017), .B(n15018), .Z(n15016) );
  NAND U16507 ( .A(n15018), .B(n15017), .Z(n15013) );
  XOR U16508 ( .A(n1555), .B(n1554), .Z(\A1[312] ) );
  XOR U16509 ( .A(n15018), .B(n15019), .Z(n1554) );
  XNOR U16510 ( .A(n15017), .B(n15015), .Z(n15019) );
  AND U16511 ( .A(n15020), .B(n15021), .Z(n15015) );
  NANDN U16512 ( .A(n15022), .B(n15023), .Z(n15021) );
  NANDN U16513 ( .A(n15024), .B(n15025), .Z(n15023) );
  AND U16514 ( .A(B[311]), .B(A[3]), .Z(n15017) );
  XNOR U16515 ( .A(n15007), .B(n15026), .Z(n15018) );
  XNOR U16516 ( .A(n15005), .B(n15008), .Z(n15026) );
  NAND U16517 ( .A(A[2]), .B(B[312]), .Z(n15008) );
  NANDN U16518 ( .A(n15027), .B(n15028), .Z(n15005) );
  AND U16519 ( .A(A[0]), .B(B[313]), .Z(n15028) );
  XOR U16520 ( .A(n15010), .B(n15029), .Z(n15007) );
  NAND U16521 ( .A(A[0]), .B(B[314]), .Z(n15029) );
  NAND U16522 ( .A(B[313]), .B(A[1]), .Z(n15010) );
  NAND U16523 ( .A(n15030), .B(n15031), .Z(n1555) );
  NANDN U16524 ( .A(n15032), .B(n15033), .Z(n15031) );
  OR U16525 ( .A(n15034), .B(n15035), .Z(n15033) );
  NAND U16526 ( .A(n15035), .B(n15034), .Z(n15030) );
  XOR U16527 ( .A(n1557), .B(n1556), .Z(\A1[311] ) );
  XOR U16528 ( .A(n15035), .B(n15036), .Z(n1556) );
  XNOR U16529 ( .A(n15034), .B(n15032), .Z(n15036) );
  AND U16530 ( .A(n15037), .B(n15038), .Z(n15032) );
  NANDN U16531 ( .A(n15039), .B(n15040), .Z(n15038) );
  NANDN U16532 ( .A(n15041), .B(n15042), .Z(n15040) );
  AND U16533 ( .A(B[310]), .B(A[3]), .Z(n15034) );
  XNOR U16534 ( .A(n15024), .B(n15043), .Z(n15035) );
  XNOR U16535 ( .A(n15022), .B(n15025), .Z(n15043) );
  NAND U16536 ( .A(A[2]), .B(B[311]), .Z(n15025) );
  NANDN U16537 ( .A(n15044), .B(n15045), .Z(n15022) );
  AND U16538 ( .A(A[0]), .B(B[312]), .Z(n15045) );
  XOR U16539 ( .A(n15027), .B(n15046), .Z(n15024) );
  NAND U16540 ( .A(A[0]), .B(B[313]), .Z(n15046) );
  NAND U16541 ( .A(B[312]), .B(A[1]), .Z(n15027) );
  NAND U16542 ( .A(n15047), .B(n15048), .Z(n1557) );
  NANDN U16543 ( .A(n15049), .B(n15050), .Z(n15048) );
  OR U16544 ( .A(n15051), .B(n15052), .Z(n15050) );
  NAND U16545 ( .A(n15052), .B(n15051), .Z(n15047) );
  XOR U16546 ( .A(n1559), .B(n1558), .Z(\A1[310] ) );
  XOR U16547 ( .A(n15052), .B(n15053), .Z(n1558) );
  XNOR U16548 ( .A(n15051), .B(n15049), .Z(n15053) );
  AND U16549 ( .A(n15054), .B(n15055), .Z(n15049) );
  NANDN U16550 ( .A(n15056), .B(n15057), .Z(n15055) );
  NANDN U16551 ( .A(n15058), .B(n15059), .Z(n15057) );
  AND U16552 ( .A(B[309]), .B(A[3]), .Z(n15051) );
  XNOR U16553 ( .A(n15041), .B(n15060), .Z(n15052) );
  XNOR U16554 ( .A(n15039), .B(n15042), .Z(n15060) );
  NAND U16555 ( .A(A[2]), .B(B[310]), .Z(n15042) );
  NANDN U16556 ( .A(n15061), .B(n15062), .Z(n15039) );
  AND U16557 ( .A(A[0]), .B(B[311]), .Z(n15062) );
  XOR U16558 ( .A(n15044), .B(n15063), .Z(n15041) );
  NAND U16559 ( .A(A[0]), .B(B[312]), .Z(n15063) );
  NAND U16560 ( .A(B[311]), .B(A[1]), .Z(n15044) );
  NAND U16561 ( .A(n15064), .B(n15065), .Z(n1559) );
  NANDN U16562 ( .A(n15066), .B(n15067), .Z(n15065) );
  OR U16563 ( .A(n15068), .B(n15069), .Z(n15067) );
  NAND U16564 ( .A(n15069), .B(n15068), .Z(n15064) );
  XOR U16565 ( .A(n1541), .B(n1540), .Z(\A1[30] ) );
  XOR U16566 ( .A(n14899), .B(n15070), .Z(n1540) );
  XNOR U16567 ( .A(n14898), .B(n14896), .Z(n15070) );
  AND U16568 ( .A(n15071), .B(n15072), .Z(n14896) );
  NANDN U16569 ( .A(n15073), .B(n15074), .Z(n15072) );
  NANDN U16570 ( .A(n15075), .B(n15076), .Z(n15074) );
  AND U16571 ( .A(B[29]), .B(A[3]), .Z(n14898) );
  XNOR U16572 ( .A(n14888), .B(n15077), .Z(n14899) );
  XNOR U16573 ( .A(n14886), .B(n14889), .Z(n15077) );
  NAND U16574 ( .A(A[2]), .B(B[30]), .Z(n14889) );
  NANDN U16575 ( .A(n15078), .B(n15079), .Z(n14886) );
  AND U16576 ( .A(A[0]), .B(B[31]), .Z(n15079) );
  XOR U16577 ( .A(n14891), .B(n15080), .Z(n14888) );
  NAND U16578 ( .A(A[0]), .B(B[32]), .Z(n15080) );
  NAND U16579 ( .A(B[31]), .B(A[1]), .Z(n14891) );
  NAND U16580 ( .A(n15081), .B(n15082), .Z(n1541) );
  NANDN U16581 ( .A(n15083), .B(n15084), .Z(n15082) );
  OR U16582 ( .A(n15085), .B(n15086), .Z(n15084) );
  NAND U16583 ( .A(n15086), .B(n15085), .Z(n15081) );
  XOR U16584 ( .A(n1561), .B(n1560), .Z(\A1[309] ) );
  XOR U16585 ( .A(n15069), .B(n15087), .Z(n1560) );
  XNOR U16586 ( .A(n15068), .B(n15066), .Z(n15087) );
  AND U16587 ( .A(n15088), .B(n15089), .Z(n15066) );
  NANDN U16588 ( .A(n15090), .B(n15091), .Z(n15089) );
  NANDN U16589 ( .A(n15092), .B(n15093), .Z(n15091) );
  AND U16590 ( .A(B[308]), .B(A[3]), .Z(n15068) );
  XNOR U16591 ( .A(n15058), .B(n15094), .Z(n15069) );
  XNOR U16592 ( .A(n15056), .B(n15059), .Z(n15094) );
  NAND U16593 ( .A(A[2]), .B(B[309]), .Z(n15059) );
  NANDN U16594 ( .A(n15095), .B(n15096), .Z(n15056) );
  AND U16595 ( .A(A[0]), .B(B[310]), .Z(n15096) );
  XOR U16596 ( .A(n15061), .B(n15097), .Z(n15058) );
  NAND U16597 ( .A(A[0]), .B(B[311]), .Z(n15097) );
  NAND U16598 ( .A(B[310]), .B(A[1]), .Z(n15061) );
  NAND U16599 ( .A(n15098), .B(n15099), .Z(n1561) );
  NANDN U16600 ( .A(n15100), .B(n15101), .Z(n15099) );
  OR U16601 ( .A(n15102), .B(n15103), .Z(n15101) );
  NAND U16602 ( .A(n15103), .B(n15102), .Z(n15098) );
  XOR U16603 ( .A(n1565), .B(n1564), .Z(\A1[308] ) );
  XOR U16604 ( .A(n15103), .B(n15104), .Z(n1564) );
  XNOR U16605 ( .A(n15102), .B(n15100), .Z(n15104) );
  AND U16606 ( .A(n15105), .B(n15106), .Z(n15100) );
  NANDN U16607 ( .A(n15107), .B(n15108), .Z(n15106) );
  NANDN U16608 ( .A(n15109), .B(n15110), .Z(n15108) );
  AND U16609 ( .A(B[307]), .B(A[3]), .Z(n15102) );
  XNOR U16610 ( .A(n15092), .B(n15111), .Z(n15103) );
  XNOR U16611 ( .A(n15090), .B(n15093), .Z(n15111) );
  NAND U16612 ( .A(A[2]), .B(B[308]), .Z(n15093) );
  NANDN U16613 ( .A(n15112), .B(n15113), .Z(n15090) );
  AND U16614 ( .A(A[0]), .B(B[309]), .Z(n15113) );
  XOR U16615 ( .A(n15095), .B(n15114), .Z(n15092) );
  NAND U16616 ( .A(A[0]), .B(B[310]), .Z(n15114) );
  NAND U16617 ( .A(B[309]), .B(A[1]), .Z(n15095) );
  NAND U16618 ( .A(n15115), .B(n15116), .Z(n1565) );
  NANDN U16619 ( .A(n15117), .B(n15118), .Z(n15116) );
  OR U16620 ( .A(n15119), .B(n15120), .Z(n15118) );
  NAND U16621 ( .A(n15120), .B(n15119), .Z(n15115) );
  XOR U16622 ( .A(n1567), .B(n1566), .Z(\A1[307] ) );
  XOR U16623 ( .A(n15120), .B(n15121), .Z(n1566) );
  XNOR U16624 ( .A(n15119), .B(n15117), .Z(n15121) );
  AND U16625 ( .A(n15122), .B(n15123), .Z(n15117) );
  NANDN U16626 ( .A(n15124), .B(n15125), .Z(n15123) );
  NANDN U16627 ( .A(n15126), .B(n15127), .Z(n15125) );
  AND U16628 ( .A(B[306]), .B(A[3]), .Z(n15119) );
  XNOR U16629 ( .A(n15109), .B(n15128), .Z(n15120) );
  XNOR U16630 ( .A(n15107), .B(n15110), .Z(n15128) );
  NAND U16631 ( .A(A[2]), .B(B[307]), .Z(n15110) );
  NANDN U16632 ( .A(n15129), .B(n15130), .Z(n15107) );
  AND U16633 ( .A(A[0]), .B(B[308]), .Z(n15130) );
  XOR U16634 ( .A(n15112), .B(n15131), .Z(n15109) );
  NAND U16635 ( .A(A[0]), .B(B[309]), .Z(n15131) );
  NAND U16636 ( .A(B[308]), .B(A[1]), .Z(n15112) );
  NAND U16637 ( .A(n15132), .B(n15133), .Z(n1567) );
  NANDN U16638 ( .A(n15134), .B(n15135), .Z(n15133) );
  OR U16639 ( .A(n15136), .B(n15137), .Z(n15135) );
  NAND U16640 ( .A(n15137), .B(n15136), .Z(n15132) );
  XOR U16641 ( .A(n1569), .B(n1568), .Z(\A1[306] ) );
  XOR U16642 ( .A(n15137), .B(n15138), .Z(n1568) );
  XNOR U16643 ( .A(n15136), .B(n15134), .Z(n15138) );
  AND U16644 ( .A(n15139), .B(n15140), .Z(n15134) );
  NANDN U16645 ( .A(n15141), .B(n15142), .Z(n15140) );
  NANDN U16646 ( .A(n15143), .B(n15144), .Z(n15142) );
  AND U16647 ( .A(B[305]), .B(A[3]), .Z(n15136) );
  XNOR U16648 ( .A(n15126), .B(n15145), .Z(n15137) );
  XNOR U16649 ( .A(n15124), .B(n15127), .Z(n15145) );
  NAND U16650 ( .A(A[2]), .B(B[306]), .Z(n15127) );
  NANDN U16651 ( .A(n15146), .B(n15147), .Z(n15124) );
  AND U16652 ( .A(A[0]), .B(B[307]), .Z(n15147) );
  XOR U16653 ( .A(n15129), .B(n15148), .Z(n15126) );
  NAND U16654 ( .A(A[0]), .B(B[308]), .Z(n15148) );
  NAND U16655 ( .A(B[307]), .B(A[1]), .Z(n15129) );
  NAND U16656 ( .A(n15149), .B(n15150), .Z(n1569) );
  NANDN U16657 ( .A(n15151), .B(n15152), .Z(n15150) );
  OR U16658 ( .A(n15153), .B(n15154), .Z(n15152) );
  NAND U16659 ( .A(n15154), .B(n15153), .Z(n15149) );
  XOR U16660 ( .A(n1571), .B(n1570), .Z(\A1[305] ) );
  XOR U16661 ( .A(n15154), .B(n15155), .Z(n1570) );
  XNOR U16662 ( .A(n15153), .B(n15151), .Z(n15155) );
  AND U16663 ( .A(n15156), .B(n15157), .Z(n15151) );
  NANDN U16664 ( .A(n15158), .B(n15159), .Z(n15157) );
  NANDN U16665 ( .A(n15160), .B(n15161), .Z(n15159) );
  AND U16666 ( .A(B[304]), .B(A[3]), .Z(n15153) );
  XNOR U16667 ( .A(n15143), .B(n15162), .Z(n15154) );
  XNOR U16668 ( .A(n15141), .B(n15144), .Z(n15162) );
  NAND U16669 ( .A(A[2]), .B(B[305]), .Z(n15144) );
  NANDN U16670 ( .A(n15163), .B(n15164), .Z(n15141) );
  AND U16671 ( .A(A[0]), .B(B[306]), .Z(n15164) );
  XOR U16672 ( .A(n15146), .B(n15165), .Z(n15143) );
  NAND U16673 ( .A(A[0]), .B(B[307]), .Z(n15165) );
  NAND U16674 ( .A(B[306]), .B(A[1]), .Z(n15146) );
  NAND U16675 ( .A(n15166), .B(n15167), .Z(n1571) );
  NANDN U16676 ( .A(n15168), .B(n15169), .Z(n15167) );
  OR U16677 ( .A(n15170), .B(n15171), .Z(n15169) );
  NAND U16678 ( .A(n15171), .B(n15170), .Z(n15166) );
  XOR U16679 ( .A(n1573), .B(n1572), .Z(\A1[304] ) );
  XOR U16680 ( .A(n15171), .B(n15172), .Z(n1572) );
  XNOR U16681 ( .A(n15170), .B(n15168), .Z(n15172) );
  AND U16682 ( .A(n15173), .B(n15174), .Z(n15168) );
  NANDN U16683 ( .A(n15175), .B(n15176), .Z(n15174) );
  NANDN U16684 ( .A(n15177), .B(n15178), .Z(n15176) );
  AND U16685 ( .A(B[303]), .B(A[3]), .Z(n15170) );
  XNOR U16686 ( .A(n15160), .B(n15179), .Z(n15171) );
  XNOR U16687 ( .A(n15158), .B(n15161), .Z(n15179) );
  NAND U16688 ( .A(A[2]), .B(B[304]), .Z(n15161) );
  NANDN U16689 ( .A(n15180), .B(n15181), .Z(n15158) );
  AND U16690 ( .A(A[0]), .B(B[305]), .Z(n15181) );
  XOR U16691 ( .A(n15163), .B(n15182), .Z(n15160) );
  NAND U16692 ( .A(A[0]), .B(B[306]), .Z(n15182) );
  NAND U16693 ( .A(B[305]), .B(A[1]), .Z(n15163) );
  NAND U16694 ( .A(n15183), .B(n15184), .Z(n1573) );
  NANDN U16695 ( .A(n15185), .B(n15186), .Z(n15184) );
  OR U16696 ( .A(n15187), .B(n15188), .Z(n15186) );
  NAND U16697 ( .A(n15188), .B(n15187), .Z(n15183) );
  XOR U16698 ( .A(n1575), .B(n1574), .Z(\A1[303] ) );
  XOR U16699 ( .A(n15188), .B(n15189), .Z(n1574) );
  XNOR U16700 ( .A(n15187), .B(n15185), .Z(n15189) );
  AND U16701 ( .A(n15190), .B(n15191), .Z(n15185) );
  NANDN U16702 ( .A(n15192), .B(n15193), .Z(n15191) );
  NANDN U16703 ( .A(n15194), .B(n15195), .Z(n15193) );
  AND U16704 ( .A(B[302]), .B(A[3]), .Z(n15187) );
  XNOR U16705 ( .A(n15177), .B(n15196), .Z(n15188) );
  XNOR U16706 ( .A(n15175), .B(n15178), .Z(n15196) );
  NAND U16707 ( .A(A[2]), .B(B[303]), .Z(n15178) );
  NANDN U16708 ( .A(n15197), .B(n15198), .Z(n15175) );
  AND U16709 ( .A(A[0]), .B(B[304]), .Z(n15198) );
  XOR U16710 ( .A(n15180), .B(n15199), .Z(n15177) );
  NAND U16711 ( .A(A[0]), .B(B[305]), .Z(n15199) );
  NAND U16712 ( .A(B[304]), .B(A[1]), .Z(n15180) );
  NAND U16713 ( .A(n15200), .B(n15201), .Z(n1575) );
  NANDN U16714 ( .A(n15202), .B(n15203), .Z(n15201) );
  OR U16715 ( .A(n15204), .B(n15205), .Z(n15203) );
  NAND U16716 ( .A(n15205), .B(n15204), .Z(n15200) );
  XOR U16717 ( .A(n1577), .B(n1576), .Z(\A1[302] ) );
  XOR U16718 ( .A(n15205), .B(n15206), .Z(n1576) );
  XNOR U16719 ( .A(n15204), .B(n15202), .Z(n15206) );
  AND U16720 ( .A(n15207), .B(n15208), .Z(n15202) );
  NANDN U16721 ( .A(n15209), .B(n15210), .Z(n15208) );
  NANDN U16722 ( .A(n15211), .B(n15212), .Z(n15210) );
  AND U16723 ( .A(B[301]), .B(A[3]), .Z(n15204) );
  XNOR U16724 ( .A(n15194), .B(n15213), .Z(n15205) );
  XNOR U16725 ( .A(n15192), .B(n15195), .Z(n15213) );
  NAND U16726 ( .A(A[2]), .B(B[302]), .Z(n15195) );
  NANDN U16727 ( .A(n15214), .B(n15215), .Z(n15192) );
  AND U16728 ( .A(A[0]), .B(B[303]), .Z(n15215) );
  XOR U16729 ( .A(n15197), .B(n15216), .Z(n15194) );
  NAND U16730 ( .A(A[0]), .B(B[304]), .Z(n15216) );
  NAND U16731 ( .A(B[303]), .B(A[1]), .Z(n15197) );
  NAND U16732 ( .A(n15217), .B(n15218), .Z(n1577) );
  NANDN U16733 ( .A(n15219), .B(n15220), .Z(n15218) );
  OR U16734 ( .A(n15221), .B(n15222), .Z(n15220) );
  NAND U16735 ( .A(n15222), .B(n15221), .Z(n15217) );
  XOR U16736 ( .A(n1579), .B(n1578), .Z(\A1[301] ) );
  XOR U16737 ( .A(n15222), .B(n15223), .Z(n1578) );
  XNOR U16738 ( .A(n15221), .B(n15219), .Z(n15223) );
  AND U16739 ( .A(n15224), .B(n15225), .Z(n15219) );
  NANDN U16740 ( .A(n15226), .B(n15227), .Z(n15225) );
  NANDN U16741 ( .A(n15228), .B(n15229), .Z(n15227) );
  AND U16742 ( .A(B[300]), .B(A[3]), .Z(n15221) );
  XNOR U16743 ( .A(n15211), .B(n15230), .Z(n15222) );
  XNOR U16744 ( .A(n15209), .B(n15212), .Z(n15230) );
  NAND U16745 ( .A(A[2]), .B(B[301]), .Z(n15212) );
  NANDN U16746 ( .A(n15231), .B(n15232), .Z(n15209) );
  AND U16747 ( .A(A[0]), .B(B[302]), .Z(n15232) );
  XOR U16748 ( .A(n15214), .B(n15233), .Z(n15211) );
  NAND U16749 ( .A(A[0]), .B(B[303]), .Z(n15233) );
  NAND U16750 ( .A(B[302]), .B(A[1]), .Z(n15214) );
  NAND U16751 ( .A(n15234), .B(n15235), .Z(n1579) );
  NANDN U16752 ( .A(n15236), .B(n15237), .Z(n15235) );
  OR U16753 ( .A(n15238), .B(n15239), .Z(n15237) );
  NAND U16754 ( .A(n15239), .B(n15238), .Z(n15234) );
  XOR U16755 ( .A(n1581), .B(n1580), .Z(\A1[300] ) );
  XOR U16756 ( .A(n15239), .B(n15240), .Z(n1580) );
  XNOR U16757 ( .A(n15238), .B(n15236), .Z(n15240) );
  AND U16758 ( .A(n15241), .B(n15242), .Z(n15236) );
  NANDN U16759 ( .A(n15243), .B(n15244), .Z(n15242) );
  NANDN U16760 ( .A(n15245), .B(n15246), .Z(n15244) );
  AND U16761 ( .A(B[299]), .B(A[3]), .Z(n15238) );
  XNOR U16762 ( .A(n15228), .B(n15247), .Z(n15239) );
  XNOR U16763 ( .A(n15226), .B(n15229), .Z(n15247) );
  NAND U16764 ( .A(A[2]), .B(B[300]), .Z(n15229) );
  NANDN U16765 ( .A(n15248), .B(n15249), .Z(n15226) );
  AND U16766 ( .A(A[0]), .B(B[301]), .Z(n15249) );
  XOR U16767 ( .A(n15231), .B(n15250), .Z(n15228) );
  NAND U16768 ( .A(A[0]), .B(B[302]), .Z(n15250) );
  NAND U16769 ( .A(B[301]), .B(A[1]), .Z(n15231) );
  NAND U16770 ( .A(n15251), .B(n15252), .Z(n1581) );
  NANDN U16771 ( .A(n15253), .B(n15254), .Z(n15252) );
  OR U16772 ( .A(n15255), .B(n15256), .Z(n15254) );
  NAND U16773 ( .A(n15256), .B(n15255), .Z(n15251) );
  XOR U16774 ( .A(n1363), .B(n1362), .Z(\A1[2] ) );
  XOR U16775 ( .A(n13386), .B(n15257), .Z(n1362) );
  XNOR U16776 ( .A(n13385), .B(n13383), .Z(n15257) );
  AND U16777 ( .A(n15258), .B(n15259), .Z(n13383) );
  NANDN U16778 ( .A(n15260), .B(n15261), .Z(n15259) );
  NANDN U16779 ( .A(n15262), .B(n15263), .Z(n15261) );
  AND U16780 ( .A(B[1]), .B(A[3]), .Z(n13385) );
  XNOR U16781 ( .A(n13375), .B(n15264), .Z(n13386) );
  XNOR U16782 ( .A(n13373), .B(n13376), .Z(n15264) );
  NAND U16783 ( .A(A[2]), .B(B[2]), .Z(n13376) );
  NANDN U16784 ( .A(n15265), .B(n15266), .Z(n13373) );
  AND U16785 ( .A(A[0]), .B(B[3]), .Z(n15266) );
  XOR U16786 ( .A(n13378), .B(n15267), .Z(n13375) );
  NAND U16787 ( .A(A[0]), .B(B[4]), .Z(n15267) );
  NAND U16788 ( .A(B[3]), .B(A[1]), .Z(n13378) );
  NAND U16789 ( .A(n15268), .B(n15269), .Z(n1363) );
  NANDN U16790 ( .A(n15270), .B(n15271), .Z(n15269) );
  OR U16791 ( .A(n15272), .B(n15273), .Z(n15271) );
  NAND U16792 ( .A(n15273), .B(n15272), .Z(n15268) );
  XOR U16793 ( .A(n1563), .B(n1562), .Z(\A1[29] ) );
  XOR U16794 ( .A(n15086), .B(n15274), .Z(n1562) );
  XNOR U16795 ( .A(n15085), .B(n15083), .Z(n15274) );
  AND U16796 ( .A(n15275), .B(n15276), .Z(n15083) );
  NANDN U16797 ( .A(n15277), .B(n15278), .Z(n15276) );
  NANDN U16798 ( .A(n15279), .B(n15280), .Z(n15278) );
  AND U16799 ( .A(B[28]), .B(A[3]), .Z(n15085) );
  XNOR U16800 ( .A(n15075), .B(n15281), .Z(n15086) );
  XNOR U16801 ( .A(n15073), .B(n15076), .Z(n15281) );
  NAND U16802 ( .A(A[2]), .B(B[29]), .Z(n15076) );
  NANDN U16803 ( .A(n15282), .B(n15283), .Z(n15073) );
  AND U16804 ( .A(A[0]), .B(B[30]), .Z(n15283) );
  XOR U16805 ( .A(n15078), .B(n15284), .Z(n15075) );
  NAND U16806 ( .A(A[0]), .B(B[31]), .Z(n15284) );
  NAND U16807 ( .A(B[30]), .B(A[1]), .Z(n15078) );
  NAND U16808 ( .A(n15285), .B(n15286), .Z(n1563) );
  NANDN U16809 ( .A(n15287), .B(n15288), .Z(n15286) );
  OR U16810 ( .A(n15289), .B(n15290), .Z(n15288) );
  NAND U16811 ( .A(n15290), .B(n15289), .Z(n15285) );
  XOR U16812 ( .A(n1583), .B(n1582), .Z(\A1[299] ) );
  XOR U16813 ( .A(n15256), .B(n15291), .Z(n1582) );
  XNOR U16814 ( .A(n15255), .B(n15253), .Z(n15291) );
  AND U16815 ( .A(n15292), .B(n15293), .Z(n15253) );
  NANDN U16816 ( .A(n15294), .B(n15295), .Z(n15293) );
  NANDN U16817 ( .A(n15296), .B(n15297), .Z(n15295) );
  AND U16818 ( .A(B[298]), .B(A[3]), .Z(n15255) );
  XNOR U16819 ( .A(n15245), .B(n15298), .Z(n15256) );
  XNOR U16820 ( .A(n15243), .B(n15246), .Z(n15298) );
  NAND U16821 ( .A(A[2]), .B(B[299]), .Z(n15246) );
  NANDN U16822 ( .A(n15299), .B(n15300), .Z(n15243) );
  AND U16823 ( .A(A[0]), .B(B[300]), .Z(n15300) );
  XOR U16824 ( .A(n15248), .B(n15301), .Z(n15245) );
  NAND U16825 ( .A(A[0]), .B(B[301]), .Z(n15301) );
  NAND U16826 ( .A(B[300]), .B(A[1]), .Z(n15248) );
  NAND U16827 ( .A(n15302), .B(n15303), .Z(n1583) );
  NANDN U16828 ( .A(n15304), .B(n15305), .Z(n15303) );
  OR U16829 ( .A(n15306), .B(n15307), .Z(n15305) );
  NAND U16830 ( .A(n15307), .B(n15306), .Z(n15302) );
  XOR U16831 ( .A(n1587), .B(n1586), .Z(\A1[298] ) );
  XOR U16832 ( .A(n15307), .B(n15308), .Z(n1586) );
  XNOR U16833 ( .A(n15306), .B(n15304), .Z(n15308) );
  AND U16834 ( .A(n15309), .B(n15310), .Z(n15304) );
  NANDN U16835 ( .A(n15311), .B(n15312), .Z(n15310) );
  NANDN U16836 ( .A(n15313), .B(n15314), .Z(n15312) );
  AND U16837 ( .A(B[297]), .B(A[3]), .Z(n15306) );
  XNOR U16838 ( .A(n15296), .B(n15315), .Z(n15307) );
  XNOR U16839 ( .A(n15294), .B(n15297), .Z(n15315) );
  NAND U16840 ( .A(A[2]), .B(B[298]), .Z(n15297) );
  NANDN U16841 ( .A(n15316), .B(n15317), .Z(n15294) );
  AND U16842 ( .A(A[0]), .B(B[299]), .Z(n15317) );
  XOR U16843 ( .A(n15299), .B(n15318), .Z(n15296) );
  NAND U16844 ( .A(A[0]), .B(B[300]), .Z(n15318) );
  NAND U16845 ( .A(B[299]), .B(A[1]), .Z(n15299) );
  NAND U16846 ( .A(n15319), .B(n15320), .Z(n1587) );
  NANDN U16847 ( .A(n15321), .B(n15322), .Z(n15320) );
  OR U16848 ( .A(n15323), .B(n15324), .Z(n15322) );
  NAND U16849 ( .A(n15324), .B(n15323), .Z(n15319) );
  XOR U16850 ( .A(n1589), .B(n1588), .Z(\A1[297] ) );
  XOR U16851 ( .A(n15324), .B(n15325), .Z(n1588) );
  XNOR U16852 ( .A(n15323), .B(n15321), .Z(n15325) );
  AND U16853 ( .A(n15326), .B(n15327), .Z(n15321) );
  NANDN U16854 ( .A(n15328), .B(n15329), .Z(n15327) );
  NANDN U16855 ( .A(n15330), .B(n15331), .Z(n15329) );
  AND U16856 ( .A(B[296]), .B(A[3]), .Z(n15323) );
  XNOR U16857 ( .A(n15313), .B(n15332), .Z(n15324) );
  XNOR U16858 ( .A(n15311), .B(n15314), .Z(n15332) );
  NAND U16859 ( .A(A[2]), .B(B[297]), .Z(n15314) );
  NANDN U16860 ( .A(n15333), .B(n15334), .Z(n15311) );
  AND U16861 ( .A(A[0]), .B(B[298]), .Z(n15334) );
  XOR U16862 ( .A(n15316), .B(n15335), .Z(n15313) );
  NAND U16863 ( .A(A[0]), .B(B[299]), .Z(n15335) );
  NAND U16864 ( .A(B[298]), .B(A[1]), .Z(n15316) );
  NAND U16865 ( .A(n15336), .B(n15337), .Z(n1589) );
  NANDN U16866 ( .A(n15338), .B(n15339), .Z(n15337) );
  OR U16867 ( .A(n15340), .B(n15341), .Z(n15339) );
  NAND U16868 ( .A(n15341), .B(n15340), .Z(n15336) );
  XOR U16869 ( .A(n1591), .B(n1590), .Z(\A1[296] ) );
  XOR U16870 ( .A(n15341), .B(n15342), .Z(n1590) );
  XNOR U16871 ( .A(n15340), .B(n15338), .Z(n15342) );
  AND U16872 ( .A(n15343), .B(n15344), .Z(n15338) );
  NANDN U16873 ( .A(n15345), .B(n15346), .Z(n15344) );
  NANDN U16874 ( .A(n15347), .B(n15348), .Z(n15346) );
  AND U16875 ( .A(B[295]), .B(A[3]), .Z(n15340) );
  XNOR U16876 ( .A(n15330), .B(n15349), .Z(n15341) );
  XNOR U16877 ( .A(n15328), .B(n15331), .Z(n15349) );
  NAND U16878 ( .A(A[2]), .B(B[296]), .Z(n15331) );
  NANDN U16879 ( .A(n15350), .B(n15351), .Z(n15328) );
  AND U16880 ( .A(A[0]), .B(B[297]), .Z(n15351) );
  XOR U16881 ( .A(n15333), .B(n15352), .Z(n15330) );
  NAND U16882 ( .A(A[0]), .B(B[298]), .Z(n15352) );
  NAND U16883 ( .A(B[297]), .B(A[1]), .Z(n15333) );
  NAND U16884 ( .A(n15353), .B(n15354), .Z(n1591) );
  NANDN U16885 ( .A(n15355), .B(n15356), .Z(n15354) );
  OR U16886 ( .A(n15357), .B(n15358), .Z(n15356) );
  NAND U16887 ( .A(n15358), .B(n15357), .Z(n15353) );
  XOR U16888 ( .A(n1593), .B(n1592), .Z(\A1[295] ) );
  XOR U16889 ( .A(n15358), .B(n15359), .Z(n1592) );
  XNOR U16890 ( .A(n15357), .B(n15355), .Z(n15359) );
  AND U16891 ( .A(n15360), .B(n15361), .Z(n15355) );
  NANDN U16892 ( .A(n15362), .B(n15363), .Z(n15361) );
  NANDN U16893 ( .A(n15364), .B(n15365), .Z(n15363) );
  AND U16894 ( .A(B[294]), .B(A[3]), .Z(n15357) );
  XNOR U16895 ( .A(n15347), .B(n15366), .Z(n15358) );
  XNOR U16896 ( .A(n15345), .B(n15348), .Z(n15366) );
  NAND U16897 ( .A(A[2]), .B(B[295]), .Z(n15348) );
  NANDN U16898 ( .A(n15367), .B(n15368), .Z(n15345) );
  AND U16899 ( .A(A[0]), .B(B[296]), .Z(n15368) );
  XOR U16900 ( .A(n15350), .B(n15369), .Z(n15347) );
  NAND U16901 ( .A(A[0]), .B(B[297]), .Z(n15369) );
  NAND U16902 ( .A(B[296]), .B(A[1]), .Z(n15350) );
  NAND U16903 ( .A(n15370), .B(n15371), .Z(n1593) );
  NANDN U16904 ( .A(n15372), .B(n15373), .Z(n15371) );
  OR U16905 ( .A(n15374), .B(n15375), .Z(n15373) );
  NAND U16906 ( .A(n15375), .B(n15374), .Z(n15370) );
  XOR U16907 ( .A(n1595), .B(n1594), .Z(\A1[294] ) );
  XOR U16908 ( .A(n15375), .B(n15376), .Z(n1594) );
  XNOR U16909 ( .A(n15374), .B(n15372), .Z(n15376) );
  AND U16910 ( .A(n15377), .B(n15378), .Z(n15372) );
  NANDN U16911 ( .A(n15379), .B(n15380), .Z(n15378) );
  NANDN U16912 ( .A(n15381), .B(n15382), .Z(n15380) );
  AND U16913 ( .A(B[293]), .B(A[3]), .Z(n15374) );
  XNOR U16914 ( .A(n15364), .B(n15383), .Z(n15375) );
  XNOR U16915 ( .A(n15362), .B(n15365), .Z(n15383) );
  NAND U16916 ( .A(A[2]), .B(B[294]), .Z(n15365) );
  NANDN U16917 ( .A(n15384), .B(n15385), .Z(n15362) );
  AND U16918 ( .A(A[0]), .B(B[295]), .Z(n15385) );
  XOR U16919 ( .A(n15367), .B(n15386), .Z(n15364) );
  NAND U16920 ( .A(A[0]), .B(B[296]), .Z(n15386) );
  NAND U16921 ( .A(B[295]), .B(A[1]), .Z(n15367) );
  NAND U16922 ( .A(n15387), .B(n15388), .Z(n1595) );
  NANDN U16923 ( .A(n15389), .B(n15390), .Z(n15388) );
  OR U16924 ( .A(n15391), .B(n15392), .Z(n15390) );
  NAND U16925 ( .A(n15392), .B(n15391), .Z(n15387) );
  XOR U16926 ( .A(n1597), .B(n1596), .Z(\A1[293] ) );
  XOR U16927 ( .A(n15392), .B(n15393), .Z(n1596) );
  XNOR U16928 ( .A(n15391), .B(n15389), .Z(n15393) );
  AND U16929 ( .A(n15394), .B(n15395), .Z(n15389) );
  NANDN U16930 ( .A(n15396), .B(n15397), .Z(n15395) );
  NANDN U16931 ( .A(n15398), .B(n15399), .Z(n15397) );
  AND U16932 ( .A(B[292]), .B(A[3]), .Z(n15391) );
  XNOR U16933 ( .A(n15381), .B(n15400), .Z(n15392) );
  XNOR U16934 ( .A(n15379), .B(n15382), .Z(n15400) );
  NAND U16935 ( .A(A[2]), .B(B[293]), .Z(n15382) );
  NANDN U16936 ( .A(n15401), .B(n15402), .Z(n15379) );
  AND U16937 ( .A(A[0]), .B(B[294]), .Z(n15402) );
  XOR U16938 ( .A(n15384), .B(n15403), .Z(n15381) );
  NAND U16939 ( .A(A[0]), .B(B[295]), .Z(n15403) );
  NAND U16940 ( .A(B[294]), .B(A[1]), .Z(n15384) );
  NAND U16941 ( .A(n15404), .B(n15405), .Z(n1597) );
  NANDN U16942 ( .A(n15406), .B(n15407), .Z(n15405) );
  OR U16943 ( .A(n15408), .B(n15409), .Z(n15407) );
  NAND U16944 ( .A(n15409), .B(n15408), .Z(n15404) );
  XOR U16945 ( .A(n1599), .B(n1598), .Z(\A1[292] ) );
  XOR U16946 ( .A(n15409), .B(n15410), .Z(n1598) );
  XNOR U16947 ( .A(n15408), .B(n15406), .Z(n15410) );
  AND U16948 ( .A(n15411), .B(n15412), .Z(n15406) );
  NANDN U16949 ( .A(n15413), .B(n15414), .Z(n15412) );
  NANDN U16950 ( .A(n15415), .B(n15416), .Z(n15414) );
  AND U16951 ( .A(B[291]), .B(A[3]), .Z(n15408) );
  XNOR U16952 ( .A(n15398), .B(n15417), .Z(n15409) );
  XNOR U16953 ( .A(n15396), .B(n15399), .Z(n15417) );
  NAND U16954 ( .A(A[2]), .B(B[292]), .Z(n15399) );
  NANDN U16955 ( .A(n15418), .B(n15419), .Z(n15396) );
  AND U16956 ( .A(A[0]), .B(B[293]), .Z(n15419) );
  XOR U16957 ( .A(n15401), .B(n15420), .Z(n15398) );
  NAND U16958 ( .A(A[0]), .B(B[294]), .Z(n15420) );
  NAND U16959 ( .A(B[293]), .B(A[1]), .Z(n15401) );
  NAND U16960 ( .A(n15421), .B(n15422), .Z(n1599) );
  NANDN U16961 ( .A(n15423), .B(n15424), .Z(n15422) );
  OR U16962 ( .A(n15425), .B(n15426), .Z(n15424) );
  NAND U16963 ( .A(n15426), .B(n15425), .Z(n15421) );
  XOR U16964 ( .A(n1601), .B(n1600), .Z(\A1[291] ) );
  XOR U16965 ( .A(n15426), .B(n15427), .Z(n1600) );
  XNOR U16966 ( .A(n15425), .B(n15423), .Z(n15427) );
  AND U16967 ( .A(n15428), .B(n15429), .Z(n15423) );
  NANDN U16968 ( .A(n15430), .B(n15431), .Z(n15429) );
  NANDN U16969 ( .A(n15432), .B(n15433), .Z(n15431) );
  AND U16970 ( .A(B[290]), .B(A[3]), .Z(n15425) );
  XNOR U16971 ( .A(n15415), .B(n15434), .Z(n15426) );
  XNOR U16972 ( .A(n15413), .B(n15416), .Z(n15434) );
  NAND U16973 ( .A(A[2]), .B(B[291]), .Z(n15416) );
  NANDN U16974 ( .A(n15435), .B(n15436), .Z(n15413) );
  AND U16975 ( .A(A[0]), .B(B[292]), .Z(n15436) );
  XOR U16976 ( .A(n15418), .B(n15437), .Z(n15415) );
  NAND U16977 ( .A(A[0]), .B(B[293]), .Z(n15437) );
  NAND U16978 ( .A(B[292]), .B(A[1]), .Z(n15418) );
  NAND U16979 ( .A(n15438), .B(n15439), .Z(n1601) );
  NANDN U16980 ( .A(n15440), .B(n15441), .Z(n15439) );
  OR U16981 ( .A(n15442), .B(n15443), .Z(n15441) );
  NAND U16982 ( .A(n15443), .B(n15442), .Z(n15438) );
  XOR U16983 ( .A(n1603), .B(n1602), .Z(\A1[290] ) );
  XOR U16984 ( .A(n15443), .B(n15444), .Z(n1602) );
  XNOR U16985 ( .A(n15442), .B(n15440), .Z(n15444) );
  AND U16986 ( .A(n15445), .B(n15446), .Z(n15440) );
  NANDN U16987 ( .A(n15447), .B(n15448), .Z(n15446) );
  NANDN U16988 ( .A(n15449), .B(n15450), .Z(n15448) );
  AND U16989 ( .A(B[289]), .B(A[3]), .Z(n15442) );
  XNOR U16990 ( .A(n15432), .B(n15451), .Z(n15443) );
  XNOR U16991 ( .A(n15430), .B(n15433), .Z(n15451) );
  NAND U16992 ( .A(A[2]), .B(B[290]), .Z(n15433) );
  NANDN U16993 ( .A(n15452), .B(n15453), .Z(n15430) );
  AND U16994 ( .A(A[0]), .B(B[291]), .Z(n15453) );
  XOR U16995 ( .A(n15435), .B(n15454), .Z(n15432) );
  NAND U16996 ( .A(A[0]), .B(B[292]), .Z(n15454) );
  NAND U16997 ( .A(B[291]), .B(A[1]), .Z(n15435) );
  NAND U16998 ( .A(n15455), .B(n15456), .Z(n1603) );
  NANDN U16999 ( .A(n15457), .B(n15458), .Z(n15456) );
  OR U17000 ( .A(n15459), .B(n15460), .Z(n15458) );
  NAND U17001 ( .A(n15460), .B(n15459), .Z(n15455) );
  XOR U17002 ( .A(n1585), .B(n1584), .Z(\A1[28] ) );
  XOR U17003 ( .A(n15290), .B(n15461), .Z(n1584) );
  XNOR U17004 ( .A(n15289), .B(n15287), .Z(n15461) );
  AND U17005 ( .A(n15462), .B(n15463), .Z(n15287) );
  NANDN U17006 ( .A(n15464), .B(n15465), .Z(n15463) );
  NANDN U17007 ( .A(n15466), .B(n15467), .Z(n15465) );
  AND U17008 ( .A(B[27]), .B(A[3]), .Z(n15289) );
  XNOR U17009 ( .A(n15279), .B(n15468), .Z(n15290) );
  XNOR U17010 ( .A(n15277), .B(n15280), .Z(n15468) );
  NAND U17011 ( .A(A[2]), .B(B[28]), .Z(n15280) );
  NANDN U17012 ( .A(n15469), .B(n15470), .Z(n15277) );
  AND U17013 ( .A(A[0]), .B(B[29]), .Z(n15470) );
  XOR U17014 ( .A(n15282), .B(n15471), .Z(n15279) );
  NAND U17015 ( .A(A[0]), .B(B[30]), .Z(n15471) );
  NAND U17016 ( .A(B[29]), .B(A[1]), .Z(n15282) );
  NAND U17017 ( .A(n15472), .B(n15473), .Z(n1585) );
  NANDN U17018 ( .A(n15474), .B(n15475), .Z(n15473) );
  OR U17019 ( .A(n15476), .B(n15477), .Z(n15475) );
  NAND U17020 ( .A(n15477), .B(n15476), .Z(n15472) );
  XOR U17021 ( .A(n1605), .B(n1604), .Z(\A1[289] ) );
  XOR U17022 ( .A(n15460), .B(n15478), .Z(n1604) );
  XNOR U17023 ( .A(n15459), .B(n15457), .Z(n15478) );
  AND U17024 ( .A(n15479), .B(n15480), .Z(n15457) );
  NANDN U17025 ( .A(n15481), .B(n15482), .Z(n15480) );
  NANDN U17026 ( .A(n15483), .B(n15484), .Z(n15482) );
  AND U17027 ( .A(B[288]), .B(A[3]), .Z(n15459) );
  XNOR U17028 ( .A(n15449), .B(n15485), .Z(n15460) );
  XNOR U17029 ( .A(n15447), .B(n15450), .Z(n15485) );
  NAND U17030 ( .A(A[2]), .B(B[289]), .Z(n15450) );
  NANDN U17031 ( .A(n15486), .B(n15487), .Z(n15447) );
  AND U17032 ( .A(A[0]), .B(B[290]), .Z(n15487) );
  XOR U17033 ( .A(n15452), .B(n15488), .Z(n15449) );
  NAND U17034 ( .A(A[0]), .B(B[291]), .Z(n15488) );
  NAND U17035 ( .A(B[290]), .B(A[1]), .Z(n15452) );
  NAND U17036 ( .A(n15489), .B(n15490), .Z(n1605) );
  NANDN U17037 ( .A(n15491), .B(n15492), .Z(n15490) );
  OR U17038 ( .A(n15493), .B(n15494), .Z(n15492) );
  NAND U17039 ( .A(n15494), .B(n15493), .Z(n15489) );
  XOR U17040 ( .A(n1609), .B(n1608), .Z(\A1[288] ) );
  XOR U17041 ( .A(n15494), .B(n15495), .Z(n1608) );
  XNOR U17042 ( .A(n15493), .B(n15491), .Z(n15495) );
  AND U17043 ( .A(n15496), .B(n15497), .Z(n15491) );
  NANDN U17044 ( .A(n15498), .B(n15499), .Z(n15497) );
  NANDN U17045 ( .A(n15500), .B(n15501), .Z(n15499) );
  AND U17046 ( .A(B[287]), .B(A[3]), .Z(n15493) );
  XNOR U17047 ( .A(n15483), .B(n15502), .Z(n15494) );
  XNOR U17048 ( .A(n15481), .B(n15484), .Z(n15502) );
  NAND U17049 ( .A(A[2]), .B(B[288]), .Z(n15484) );
  NANDN U17050 ( .A(n15503), .B(n15504), .Z(n15481) );
  AND U17051 ( .A(A[0]), .B(B[289]), .Z(n15504) );
  XOR U17052 ( .A(n15486), .B(n15505), .Z(n15483) );
  NAND U17053 ( .A(A[0]), .B(B[290]), .Z(n15505) );
  NAND U17054 ( .A(B[289]), .B(A[1]), .Z(n15486) );
  NAND U17055 ( .A(n15506), .B(n15507), .Z(n1609) );
  NANDN U17056 ( .A(n15508), .B(n15509), .Z(n15507) );
  OR U17057 ( .A(n15510), .B(n15511), .Z(n15509) );
  NAND U17058 ( .A(n15511), .B(n15510), .Z(n15506) );
  XOR U17059 ( .A(n1611), .B(n1610), .Z(\A1[287] ) );
  XOR U17060 ( .A(n15511), .B(n15512), .Z(n1610) );
  XNOR U17061 ( .A(n15510), .B(n15508), .Z(n15512) );
  AND U17062 ( .A(n15513), .B(n15514), .Z(n15508) );
  NANDN U17063 ( .A(n15515), .B(n15516), .Z(n15514) );
  NANDN U17064 ( .A(n15517), .B(n15518), .Z(n15516) );
  AND U17065 ( .A(B[286]), .B(A[3]), .Z(n15510) );
  XNOR U17066 ( .A(n15500), .B(n15519), .Z(n15511) );
  XNOR U17067 ( .A(n15498), .B(n15501), .Z(n15519) );
  NAND U17068 ( .A(A[2]), .B(B[287]), .Z(n15501) );
  NANDN U17069 ( .A(n15520), .B(n15521), .Z(n15498) );
  AND U17070 ( .A(A[0]), .B(B[288]), .Z(n15521) );
  XOR U17071 ( .A(n15503), .B(n15522), .Z(n15500) );
  NAND U17072 ( .A(A[0]), .B(B[289]), .Z(n15522) );
  NAND U17073 ( .A(B[288]), .B(A[1]), .Z(n15503) );
  NAND U17074 ( .A(n15523), .B(n15524), .Z(n1611) );
  NANDN U17075 ( .A(n15525), .B(n15526), .Z(n15524) );
  OR U17076 ( .A(n15527), .B(n15528), .Z(n15526) );
  NAND U17077 ( .A(n15528), .B(n15527), .Z(n15523) );
  XOR U17078 ( .A(n1613), .B(n1612), .Z(\A1[286] ) );
  XOR U17079 ( .A(n15528), .B(n15529), .Z(n1612) );
  XNOR U17080 ( .A(n15527), .B(n15525), .Z(n15529) );
  AND U17081 ( .A(n15530), .B(n15531), .Z(n15525) );
  NANDN U17082 ( .A(n15532), .B(n15533), .Z(n15531) );
  NANDN U17083 ( .A(n15534), .B(n15535), .Z(n15533) );
  AND U17084 ( .A(B[285]), .B(A[3]), .Z(n15527) );
  XNOR U17085 ( .A(n15517), .B(n15536), .Z(n15528) );
  XNOR U17086 ( .A(n15515), .B(n15518), .Z(n15536) );
  NAND U17087 ( .A(A[2]), .B(B[286]), .Z(n15518) );
  NANDN U17088 ( .A(n15537), .B(n15538), .Z(n15515) );
  AND U17089 ( .A(A[0]), .B(B[287]), .Z(n15538) );
  XOR U17090 ( .A(n15520), .B(n15539), .Z(n15517) );
  NAND U17091 ( .A(A[0]), .B(B[288]), .Z(n15539) );
  NAND U17092 ( .A(B[287]), .B(A[1]), .Z(n15520) );
  NAND U17093 ( .A(n15540), .B(n15541), .Z(n1613) );
  NANDN U17094 ( .A(n15542), .B(n15543), .Z(n15541) );
  OR U17095 ( .A(n15544), .B(n15545), .Z(n15543) );
  NAND U17096 ( .A(n15545), .B(n15544), .Z(n15540) );
  XOR U17097 ( .A(n1615), .B(n1614), .Z(\A1[285] ) );
  XOR U17098 ( .A(n15545), .B(n15546), .Z(n1614) );
  XNOR U17099 ( .A(n15544), .B(n15542), .Z(n15546) );
  AND U17100 ( .A(n15547), .B(n15548), .Z(n15542) );
  NANDN U17101 ( .A(n15549), .B(n15550), .Z(n15548) );
  NANDN U17102 ( .A(n15551), .B(n15552), .Z(n15550) );
  AND U17103 ( .A(B[284]), .B(A[3]), .Z(n15544) );
  XNOR U17104 ( .A(n15534), .B(n15553), .Z(n15545) );
  XNOR U17105 ( .A(n15532), .B(n15535), .Z(n15553) );
  NAND U17106 ( .A(A[2]), .B(B[285]), .Z(n15535) );
  NANDN U17107 ( .A(n15554), .B(n15555), .Z(n15532) );
  AND U17108 ( .A(A[0]), .B(B[286]), .Z(n15555) );
  XOR U17109 ( .A(n15537), .B(n15556), .Z(n15534) );
  NAND U17110 ( .A(A[0]), .B(B[287]), .Z(n15556) );
  NAND U17111 ( .A(B[286]), .B(A[1]), .Z(n15537) );
  NAND U17112 ( .A(n15557), .B(n15558), .Z(n1615) );
  NANDN U17113 ( .A(n15559), .B(n15560), .Z(n15558) );
  OR U17114 ( .A(n15561), .B(n15562), .Z(n15560) );
  NAND U17115 ( .A(n15562), .B(n15561), .Z(n15557) );
  XOR U17116 ( .A(n1617), .B(n1616), .Z(\A1[284] ) );
  XOR U17117 ( .A(n15562), .B(n15563), .Z(n1616) );
  XNOR U17118 ( .A(n15561), .B(n15559), .Z(n15563) );
  AND U17119 ( .A(n15564), .B(n15565), .Z(n15559) );
  NANDN U17120 ( .A(n15566), .B(n15567), .Z(n15565) );
  NANDN U17121 ( .A(n15568), .B(n15569), .Z(n15567) );
  AND U17122 ( .A(B[283]), .B(A[3]), .Z(n15561) );
  XNOR U17123 ( .A(n15551), .B(n15570), .Z(n15562) );
  XNOR U17124 ( .A(n15549), .B(n15552), .Z(n15570) );
  NAND U17125 ( .A(A[2]), .B(B[284]), .Z(n15552) );
  NANDN U17126 ( .A(n15571), .B(n15572), .Z(n15549) );
  AND U17127 ( .A(A[0]), .B(B[285]), .Z(n15572) );
  XOR U17128 ( .A(n15554), .B(n15573), .Z(n15551) );
  NAND U17129 ( .A(A[0]), .B(B[286]), .Z(n15573) );
  NAND U17130 ( .A(B[285]), .B(A[1]), .Z(n15554) );
  NAND U17131 ( .A(n15574), .B(n15575), .Z(n1617) );
  NANDN U17132 ( .A(n15576), .B(n15577), .Z(n15575) );
  OR U17133 ( .A(n15578), .B(n15579), .Z(n15577) );
  NAND U17134 ( .A(n15579), .B(n15578), .Z(n15574) );
  XOR U17135 ( .A(n1619), .B(n1618), .Z(\A1[283] ) );
  XOR U17136 ( .A(n15579), .B(n15580), .Z(n1618) );
  XNOR U17137 ( .A(n15578), .B(n15576), .Z(n15580) );
  AND U17138 ( .A(n15581), .B(n15582), .Z(n15576) );
  NANDN U17139 ( .A(n15583), .B(n15584), .Z(n15582) );
  NANDN U17140 ( .A(n15585), .B(n15586), .Z(n15584) );
  AND U17141 ( .A(B[282]), .B(A[3]), .Z(n15578) );
  XNOR U17142 ( .A(n15568), .B(n15587), .Z(n15579) );
  XNOR U17143 ( .A(n15566), .B(n15569), .Z(n15587) );
  NAND U17144 ( .A(A[2]), .B(B[283]), .Z(n15569) );
  NANDN U17145 ( .A(n15588), .B(n15589), .Z(n15566) );
  AND U17146 ( .A(A[0]), .B(B[284]), .Z(n15589) );
  XOR U17147 ( .A(n15571), .B(n15590), .Z(n15568) );
  NAND U17148 ( .A(A[0]), .B(B[285]), .Z(n15590) );
  NAND U17149 ( .A(B[284]), .B(A[1]), .Z(n15571) );
  NAND U17150 ( .A(n15591), .B(n15592), .Z(n1619) );
  NANDN U17151 ( .A(n15593), .B(n15594), .Z(n15592) );
  OR U17152 ( .A(n15595), .B(n15596), .Z(n15594) );
  NAND U17153 ( .A(n15596), .B(n15595), .Z(n15591) );
  XOR U17154 ( .A(n1621), .B(n1620), .Z(\A1[282] ) );
  XOR U17155 ( .A(n15596), .B(n15597), .Z(n1620) );
  XNOR U17156 ( .A(n15595), .B(n15593), .Z(n15597) );
  AND U17157 ( .A(n15598), .B(n15599), .Z(n15593) );
  NANDN U17158 ( .A(n15600), .B(n15601), .Z(n15599) );
  NANDN U17159 ( .A(n15602), .B(n15603), .Z(n15601) );
  AND U17160 ( .A(B[281]), .B(A[3]), .Z(n15595) );
  XNOR U17161 ( .A(n15585), .B(n15604), .Z(n15596) );
  XNOR U17162 ( .A(n15583), .B(n15586), .Z(n15604) );
  NAND U17163 ( .A(A[2]), .B(B[282]), .Z(n15586) );
  NANDN U17164 ( .A(n15605), .B(n15606), .Z(n15583) );
  AND U17165 ( .A(A[0]), .B(B[283]), .Z(n15606) );
  XOR U17166 ( .A(n15588), .B(n15607), .Z(n15585) );
  NAND U17167 ( .A(A[0]), .B(B[284]), .Z(n15607) );
  NAND U17168 ( .A(B[283]), .B(A[1]), .Z(n15588) );
  NAND U17169 ( .A(n15608), .B(n15609), .Z(n1621) );
  NANDN U17170 ( .A(n15610), .B(n15611), .Z(n15609) );
  OR U17171 ( .A(n15612), .B(n15613), .Z(n15611) );
  NAND U17172 ( .A(n15613), .B(n15612), .Z(n15608) );
  XOR U17173 ( .A(n1623), .B(n1622), .Z(\A1[281] ) );
  XOR U17174 ( .A(n15613), .B(n15614), .Z(n1622) );
  XNOR U17175 ( .A(n15612), .B(n15610), .Z(n15614) );
  AND U17176 ( .A(n15615), .B(n15616), .Z(n15610) );
  NANDN U17177 ( .A(n15617), .B(n15618), .Z(n15616) );
  NANDN U17178 ( .A(n15619), .B(n15620), .Z(n15618) );
  AND U17179 ( .A(B[280]), .B(A[3]), .Z(n15612) );
  XNOR U17180 ( .A(n15602), .B(n15621), .Z(n15613) );
  XNOR U17181 ( .A(n15600), .B(n15603), .Z(n15621) );
  NAND U17182 ( .A(A[2]), .B(B[281]), .Z(n15603) );
  NANDN U17183 ( .A(n15622), .B(n15623), .Z(n15600) );
  AND U17184 ( .A(A[0]), .B(B[282]), .Z(n15623) );
  XOR U17185 ( .A(n15605), .B(n15624), .Z(n15602) );
  NAND U17186 ( .A(A[0]), .B(B[283]), .Z(n15624) );
  NAND U17187 ( .A(B[282]), .B(A[1]), .Z(n15605) );
  NAND U17188 ( .A(n15625), .B(n15626), .Z(n1623) );
  NANDN U17189 ( .A(n15627), .B(n15628), .Z(n15626) );
  OR U17190 ( .A(n15629), .B(n15630), .Z(n15628) );
  NAND U17191 ( .A(n15630), .B(n15629), .Z(n15625) );
  XOR U17192 ( .A(n1625), .B(n1624), .Z(\A1[280] ) );
  XOR U17193 ( .A(n15630), .B(n15631), .Z(n1624) );
  XNOR U17194 ( .A(n15629), .B(n15627), .Z(n15631) );
  AND U17195 ( .A(n15632), .B(n15633), .Z(n15627) );
  NANDN U17196 ( .A(n15634), .B(n15635), .Z(n15633) );
  NANDN U17197 ( .A(n15636), .B(n15637), .Z(n15635) );
  AND U17198 ( .A(B[279]), .B(A[3]), .Z(n15629) );
  XNOR U17199 ( .A(n15619), .B(n15638), .Z(n15630) );
  XNOR U17200 ( .A(n15617), .B(n15620), .Z(n15638) );
  NAND U17201 ( .A(A[2]), .B(B[280]), .Z(n15620) );
  NANDN U17202 ( .A(n15639), .B(n15640), .Z(n15617) );
  AND U17203 ( .A(A[0]), .B(B[281]), .Z(n15640) );
  XOR U17204 ( .A(n15622), .B(n15641), .Z(n15619) );
  NAND U17205 ( .A(A[0]), .B(B[282]), .Z(n15641) );
  NAND U17206 ( .A(B[281]), .B(A[1]), .Z(n15622) );
  NAND U17207 ( .A(n15642), .B(n15643), .Z(n1625) );
  NANDN U17208 ( .A(n15644), .B(n15645), .Z(n15643) );
  OR U17209 ( .A(n15646), .B(n15647), .Z(n15645) );
  NAND U17210 ( .A(n15647), .B(n15646), .Z(n15642) );
  XOR U17211 ( .A(n1607), .B(n1606), .Z(\A1[27] ) );
  XOR U17212 ( .A(n15477), .B(n15648), .Z(n1606) );
  XNOR U17213 ( .A(n15476), .B(n15474), .Z(n15648) );
  AND U17214 ( .A(n15649), .B(n15650), .Z(n15474) );
  NANDN U17215 ( .A(n15651), .B(n15652), .Z(n15650) );
  NANDN U17216 ( .A(n15653), .B(n15654), .Z(n15652) );
  AND U17217 ( .A(B[26]), .B(A[3]), .Z(n15476) );
  XNOR U17218 ( .A(n15466), .B(n15655), .Z(n15477) );
  XNOR U17219 ( .A(n15464), .B(n15467), .Z(n15655) );
  NAND U17220 ( .A(A[2]), .B(B[27]), .Z(n15467) );
  NANDN U17221 ( .A(n15656), .B(n15657), .Z(n15464) );
  AND U17222 ( .A(A[0]), .B(B[28]), .Z(n15657) );
  XOR U17223 ( .A(n15469), .B(n15658), .Z(n15466) );
  NAND U17224 ( .A(A[0]), .B(B[29]), .Z(n15658) );
  NAND U17225 ( .A(B[28]), .B(A[1]), .Z(n15469) );
  NAND U17226 ( .A(n15659), .B(n15660), .Z(n1607) );
  NANDN U17227 ( .A(n15661), .B(n15662), .Z(n15660) );
  OR U17228 ( .A(n15663), .B(n15664), .Z(n15662) );
  NAND U17229 ( .A(n15664), .B(n15663), .Z(n15659) );
  XOR U17230 ( .A(n1627), .B(n1626), .Z(\A1[279] ) );
  XOR U17231 ( .A(n15647), .B(n15665), .Z(n1626) );
  XNOR U17232 ( .A(n15646), .B(n15644), .Z(n15665) );
  AND U17233 ( .A(n15666), .B(n15667), .Z(n15644) );
  NANDN U17234 ( .A(n15668), .B(n15669), .Z(n15667) );
  NANDN U17235 ( .A(n15670), .B(n15671), .Z(n15669) );
  AND U17236 ( .A(B[278]), .B(A[3]), .Z(n15646) );
  XNOR U17237 ( .A(n15636), .B(n15672), .Z(n15647) );
  XNOR U17238 ( .A(n15634), .B(n15637), .Z(n15672) );
  NAND U17239 ( .A(A[2]), .B(B[279]), .Z(n15637) );
  NANDN U17240 ( .A(n15673), .B(n15674), .Z(n15634) );
  AND U17241 ( .A(A[0]), .B(B[280]), .Z(n15674) );
  XOR U17242 ( .A(n15639), .B(n15675), .Z(n15636) );
  NAND U17243 ( .A(A[0]), .B(B[281]), .Z(n15675) );
  NAND U17244 ( .A(B[280]), .B(A[1]), .Z(n15639) );
  NAND U17245 ( .A(n15676), .B(n15677), .Z(n1627) );
  NANDN U17246 ( .A(n15678), .B(n15679), .Z(n15677) );
  OR U17247 ( .A(n15680), .B(n15681), .Z(n15679) );
  NAND U17248 ( .A(n15681), .B(n15680), .Z(n15676) );
  XOR U17249 ( .A(n1631), .B(n1630), .Z(\A1[278] ) );
  XOR U17250 ( .A(n15681), .B(n15682), .Z(n1630) );
  XNOR U17251 ( .A(n15680), .B(n15678), .Z(n15682) );
  AND U17252 ( .A(n15683), .B(n15684), .Z(n15678) );
  NANDN U17253 ( .A(n15685), .B(n15686), .Z(n15684) );
  NANDN U17254 ( .A(n15687), .B(n15688), .Z(n15686) );
  AND U17255 ( .A(B[277]), .B(A[3]), .Z(n15680) );
  XNOR U17256 ( .A(n15670), .B(n15689), .Z(n15681) );
  XNOR U17257 ( .A(n15668), .B(n15671), .Z(n15689) );
  NAND U17258 ( .A(A[2]), .B(B[278]), .Z(n15671) );
  NANDN U17259 ( .A(n15690), .B(n15691), .Z(n15668) );
  AND U17260 ( .A(A[0]), .B(B[279]), .Z(n15691) );
  XOR U17261 ( .A(n15673), .B(n15692), .Z(n15670) );
  NAND U17262 ( .A(A[0]), .B(B[280]), .Z(n15692) );
  NAND U17263 ( .A(B[279]), .B(A[1]), .Z(n15673) );
  NAND U17264 ( .A(n15693), .B(n15694), .Z(n1631) );
  NANDN U17265 ( .A(n15695), .B(n15696), .Z(n15694) );
  OR U17266 ( .A(n15697), .B(n15698), .Z(n15696) );
  NAND U17267 ( .A(n15698), .B(n15697), .Z(n15693) );
  XOR U17268 ( .A(n1633), .B(n1632), .Z(\A1[277] ) );
  XOR U17269 ( .A(n15698), .B(n15699), .Z(n1632) );
  XNOR U17270 ( .A(n15697), .B(n15695), .Z(n15699) );
  AND U17271 ( .A(n15700), .B(n15701), .Z(n15695) );
  NANDN U17272 ( .A(n15702), .B(n15703), .Z(n15701) );
  NANDN U17273 ( .A(n15704), .B(n15705), .Z(n15703) );
  AND U17274 ( .A(B[276]), .B(A[3]), .Z(n15697) );
  XNOR U17275 ( .A(n15687), .B(n15706), .Z(n15698) );
  XNOR U17276 ( .A(n15685), .B(n15688), .Z(n15706) );
  NAND U17277 ( .A(A[2]), .B(B[277]), .Z(n15688) );
  NANDN U17278 ( .A(n15707), .B(n15708), .Z(n15685) );
  AND U17279 ( .A(A[0]), .B(B[278]), .Z(n15708) );
  XOR U17280 ( .A(n15690), .B(n15709), .Z(n15687) );
  NAND U17281 ( .A(A[0]), .B(B[279]), .Z(n15709) );
  NAND U17282 ( .A(B[278]), .B(A[1]), .Z(n15690) );
  NAND U17283 ( .A(n15710), .B(n15711), .Z(n1633) );
  NANDN U17284 ( .A(n15712), .B(n15713), .Z(n15711) );
  OR U17285 ( .A(n15714), .B(n15715), .Z(n15713) );
  NAND U17286 ( .A(n15715), .B(n15714), .Z(n15710) );
  XOR U17287 ( .A(n1635), .B(n1634), .Z(\A1[276] ) );
  XOR U17288 ( .A(n15715), .B(n15716), .Z(n1634) );
  XNOR U17289 ( .A(n15714), .B(n15712), .Z(n15716) );
  AND U17290 ( .A(n15717), .B(n15718), .Z(n15712) );
  NANDN U17291 ( .A(n15719), .B(n15720), .Z(n15718) );
  NANDN U17292 ( .A(n15721), .B(n15722), .Z(n15720) );
  AND U17293 ( .A(B[275]), .B(A[3]), .Z(n15714) );
  XNOR U17294 ( .A(n15704), .B(n15723), .Z(n15715) );
  XNOR U17295 ( .A(n15702), .B(n15705), .Z(n15723) );
  NAND U17296 ( .A(A[2]), .B(B[276]), .Z(n15705) );
  NANDN U17297 ( .A(n15724), .B(n15725), .Z(n15702) );
  AND U17298 ( .A(A[0]), .B(B[277]), .Z(n15725) );
  XOR U17299 ( .A(n15707), .B(n15726), .Z(n15704) );
  NAND U17300 ( .A(A[0]), .B(B[278]), .Z(n15726) );
  NAND U17301 ( .A(B[277]), .B(A[1]), .Z(n15707) );
  NAND U17302 ( .A(n15727), .B(n15728), .Z(n1635) );
  NANDN U17303 ( .A(n15729), .B(n15730), .Z(n15728) );
  OR U17304 ( .A(n15731), .B(n15732), .Z(n15730) );
  NAND U17305 ( .A(n15732), .B(n15731), .Z(n15727) );
  XOR U17306 ( .A(n1637), .B(n1636), .Z(\A1[275] ) );
  XOR U17307 ( .A(n15732), .B(n15733), .Z(n1636) );
  XNOR U17308 ( .A(n15731), .B(n15729), .Z(n15733) );
  AND U17309 ( .A(n15734), .B(n15735), .Z(n15729) );
  NANDN U17310 ( .A(n15736), .B(n15737), .Z(n15735) );
  NANDN U17311 ( .A(n15738), .B(n15739), .Z(n15737) );
  AND U17312 ( .A(B[274]), .B(A[3]), .Z(n15731) );
  XNOR U17313 ( .A(n15721), .B(n15740), .Z(n15732) );
  XNOR U17314 ( .A(n15719), .B(n15722), .Z(n15740) );
  NAND U17315 ( .A(A[2]), .B(B[275]), .Z(n15722) );
  NANDN U17316 ( .A(n15741), .B(n15742), .Z(n15719) );
  AND U17317 ( .A(A[0]), .B(B[276]), .Z(n15742) );
  XOR U17318 ( .A(n15724), .B(n15743), .Z(n15721) );
  NAND U17319 ( .A(A[0]), .B(B[277]), .Z(n15743) );
  NAND U17320 ( .A(B[276]), .B(A[1]), .Z(n15724) );
  NAND U17321 ( .A(n15744), .B(n15745), .Z(n1637) );
  NANDN U17322 ( .A(n15746), .B(n15747), .Z(n15745) );
  OR U17323 ( .A(n15748), .B(n15749), .Z(n15747) );
  NAND U17324 ( .A(n15749), .B(n15748), .Z(n15744) );
  XOR U17325 ( .A(n1639), .B(n1638), .Z(\A1[274] ) );
  XOR U17326 ( .A(n15749), .B(n15750), .Z(n1638) );
  XNOR U17327 ( .A(n15748), .B(n15746), .Z(n15750) );
  AND U17328 ( .A(n15751), .B(n15752), .Z(n15746) );
  NANDN U17329 ( .A(n15753), .B(n15754), .Z(n15752) );
  NANDN U17330 ( .A(n15755), .B(n15756), .Z(n15754) );
  AND U17331 ( .A(B[273]), .B(A[3]), .Z(n15748) );
  XNOR U17332 ( .A(n15738), .B(n15757), .Z(n15749) );
  XNOR U17333 ( .A(n15736), .B(n15739), .Z(n15757) );
  NAND U17334 ( .A(A[2]), .B(B[274]), .Z(n15739) );
  NANDN U17335 ( .A(n15758), .B(n15759), .Z(n15736) );
  AND U17336 ( .A(A[0]), .B(B[275]), .Z(n15759) );
  XOR U17337 ( .A(n15741), .B(n15760), .Z(n15738) );
  NAND U17338 ( .A(A[0]), .B(B[276]), .Z(n15760) );
  NAND U17339 ( .A(B[275]), .B(A[1]), .Z(n15741) );
  NAND U17340 ( .A(n15761), .B(n15762), .Z(n1639) );
  NANDN U17341 ( .A(n15763), .B(n15764), .Z(n15762) );
  OR U17342 ( .A(n15765), .B(n15766), .Z(n15764) );
  NAND U17343 ( .A(n15766), .B(n15765), .Z(n15761) );
  XOR U17344 ( .A(n1641), .B(n1640), .Z(\A1[273] ) );
  XOR U17345 ( .A(n15766), .B(n15767), .Z(n1640) );
  XNOR U17346 ( .A(n15765), .B(n15763), .Z(n15767) );
  AND U17347 ( .A(n15768), .B(n15769), .Z(n15763) );
  NANDN U17348 ( .A(n15770), .B(n15771), .Z(n15769) );
  NANDN U17349 ( .A(n15772), .B(n15773), .Z(n15771) );
  AND U17350 ( .A(B[272]), .B(A[3]), .Z(n15765) );
  XNOR U17351 ( .A(n15755), .B(n15774), .Z(n15766) );
  XNOR U17352 ( .A(n15753), .B(n15756), .Z(n15774) );
  NAND U17353 ( .A(A[2]), .B(B[273]), .Z(n15756) );
  NANDN U17354 ( .A(n15775), .B(n15776), .Z(n15753) );
  AND U17355 ( .A(A[0]), .B(B[274]), .Z(n15776) );
  XOR U17356 ( .A(n15758), .B(n15777), .Z(n15755) );
  NAND U17357 ( .A(A[0]), .B(B[275]), .Z(n15777) );
  NAND U17358 ( .A(B[274]), .B(A[1]), .Z(n15758) );
  NAND U17359 ( .A(n15778), .B(n15779), .Z(n1641) );
  NANDN U17360 ( .A(n15780), .B(n15781), .Z(n15779) );
  OR U17361 ( .A(n15782), .B(n15783), .Z(n15781) );
  NAND U17362 ( .A(n15783), .B(n15782), .Z(n15778) );
  XOR U17363 ( .A(n1643), .B(n1642), .Z(\A1[272] ) );
  XOR U17364 ( .A(n15783), .B(n15784), .Z(n1642) );
  XNOR U17365 ( .A(n15782), .B(n15780), .Z(n15784) );
  AND U17366 ( .A(n15785), .B(n15786), .Z(n15780) );
  NANDN U17367 ( .A(n15787), .B(n15788), .Z(n15786) );
  NANDN U17368 ( .A(n15789), .B(n15790), .Z(n15788) );
  AND U17369 ( .A(B[271]), .B(A[3]), .Z(n15782) );
  XNOR U17370 ( .A(n15772), .B(n15791), .Z(n15783) );
  XNOR U17371 ( .A(n15770), .B(n15773), .Z(n15791) );
  NAND U17372 ( .A(A[2]), .B(B[272]), .Z(n15773) );
  NANDN U17373 ( .A(n15792), .B(n15793), .Z(n15770) );
  AND U17374 ( .A(A[0]), .B(B[273]), .Z(n15793) );
  XOR U17375 ( .A(n15775), .B(n15794), .Z(n15772) );
  NAND U17376 ( .A(A[0]), .B(B[274]), .Z(n15794) );
  NAND U17377 ( .A(B[273]), .B(A[1]), .Z(n15775) );
  NAND U17378 ( .A(n15795), .B(n15796), .Z(n1643) );
  NANDN U17379 ( .A(n15797), .B(n15798), .Z(n15796) );
  OR U17380 ( .A(n15799), .B(n15800), .Z(n15798) );
  NAND U17381 ( .A(n15800), .B(n15799), .Z(n15795) );
  XOR U17382 ( .A(n1645), .B(n1644), .Z(\A1[271] ) );
  XOR U17383 ( .A(n15800), .B(n15801), .Z(n1644) );
  XNOR U17384 ( .A(n15799), .B(n15797), .Z(n15801) );
  AND U17385 ( .A(n15802), .B(n15803), .Z(n15797) );
  NANDN U17386 ( .A(n15804), .B(n15805), .Z(n15803) );
  NANDN U17387 ( .A(n15806), .B(n15807), .Z(n15805) );
  AND U17388 ( .A(B[270]), .B(A[3]), .Z(n15799) );
  XNOR U17389 ( .A(n15789), .B(n15808), .Z(n15800) );
  XNOR U17390 ( .A(n15787), .B(n15790), .Z(n15808) );
  NAND U17391 ( .A(A[2]), .B(B[271]), .Z(n15790) );
  NANDN U17392 ( .A(n15809), .B(n15810), .Z(n15787) );
  AND U17393 ( .A(A[0]), .B(B[272]), .Z(n15810) );
  XOR U17394 ( .A(n15792), .B(n15811), .Z(n15789) );
  NAND U17395 ( .A(A[0]), .B(B[273]), .Z(n15811) );
  NAND U17396 ( .A(B[272]), .B(A[1]), .Z(n15792) );
  NAND U17397 ( .A(n15812), .B(n15813), .Z(n1645) );
  NANDN U17398 ( .A(n15814), .B(n15815), .Z(n15813) );
  OR U17399 ( .A(n15816), .B(n15817), .Z(n15815) );
  NAND U17400 ( .A(n15817), .B(n15816), .Z(n15812) );
  XOR U17401 ( .A(n1647), .B(n1646), .Z(\A1[270] ) );
  XOR U17402 ( .A(n15817), .B(n15818), .Z(n1646) );
  XNOR U17403 ( .A(n15816), .B(n15814), .Z(n15818) );
  AND U17404 ( .A(n15819), .B(n15820), .Z(n15814) );
  NANDN U17405 ( .A(n15821), .B(n15822), .Z(n15820) );
  NANDN U17406 ( .A(n15823), .B(n15824), .Z(n15822) );
  AND U17407 ( .A(B[269]), .B(A[3]), .Z(n15816) );
  XNOR U17408 ( .A(n15806), .B(n15825), .Z(n15817) );
  XNOR U17409 ( .A(n15804), .B(n15807), .Z(n15825) );
  NAND U17410 ( .A(A[2]), .B(B[270]), .Z(n15807) );
  NANDN U17411 ( .A(n15826), .B(n15827), .Z(n15804) );
  AND U17412 ( .A(A[0]), .B(B[271]), .Z(n15827) );
  XOR U17413 ( .A(n15809), .B(n15828), .Z(n15806) );
  NAND U17414 ( .A(A[0]), .B(B[272]), .Z(n15828) );
  NAND U17415 ( .A(B[271]), .B(A[1]), .Z(n15809) );
  NAND U17416 ( .A(n15829), .B(n15830), .Z(n1647) );
  NANDN U17417 ( .A(n15831), .B(n15832), .Z(n15830) );
  OR U17418 ( .A(n15833), .B(n15834), .Z(n15832) );
  NAND U17419 ( .A(n15834), .B(n15833), .Z(n15829) );
  XOR U17420 ( .A(n1629), .B(n1628), .Z(\A1[26] ) );
  XOR U17421 ( .A(n15664), .B(n15835), .Z(n1628) );
  XNOR U17422 ( .A(n15663), .B(n15661), .Z(n15835) );
  AND U17423 ( .A(n15836), .B(n15837), .Z(n15661) );
  NANDN U17424 ( .A(n15838), .B(n15839), .Z(n15837) );
  NANDN U17425 ( .A(n15840), .B(n15841), .Z(n15839) );
  AND U17426 ( .A(B[25]), .B(A[3]), .Z(n15663) );
  XNOR U17427 ( .A(n15653), .B(n15842), .Z(n15664) );
  XNOR U17428 ( .A(n15651), .B(n15654), .Z(n15842) );
  NAND U17429 ( .A(A[2]), .B(B[26]), .Z(n15654) );
  NANDN U17430 ( .A(n15843), .B(n15844), .Z(n15651) );
  AND U17431 ( .A(A[0]), .B(B[27]), .Z(n15844) );
  XOR U17432 ( .A(n15656), .B(n15845), .Z(n15653) );
  NAND U17433 ( .A(A[0]), .B(B[28]), .Z(n15845) );
  NAND U17434 ( .A(B[27]), .B(A[1]), .Z(n15656) );
  NAND U17435 ( .A(n15846), .B(n15847), .Z(n1629) );
  NANDN U17436 ( .A(n15848), .B(n15849), .Z(n15847) );
  OR U17437 ( .A(n15850), .B(n15851), .Z(n15849) );
  NAND U17438 ( .A(n15851), .B(n15850), .Z(n15846) );
  XOR U17439 ( .A(n1649), .B(n1648), .Z(\A1[269] ) );
  XOR U17440 ( .A(n15834), .B(n15852), .Z(n1648) );
  XNOR U17441 ( .A(n15833), .B(n15831), .Z(n15852) );
  AND U17442 ( .A(n15853), .B(n15854), .Z(n15831) );
  NANDN U17443 ( .A(n15855), .B(n15856), .Z(n15854) );
  NANDN U17444 ( .A(n15857), .B(n15858), .Z(n15856) );
  AND U17445 ( .A(B[268]), .B(A[3]), .Z(n15833) );
  XNOR U17446 ( .A(n15823), .B(n15859), .Z(n15834) );
  XNOR U17447 ( .A(n15821), .B(n15824), .Z(n15859) );
  NAND U17448 ( .A(A[2]), .B(B[269]), .Z(n15824) );
  NANDN U17449 ( .A(n15860), .B(n15861), .Z(n15821) );
  AND U17450 ( .A(A[0]), .B(B[270]), .Z(n15861) );
  XOR U17451 ( .A(n15826), .B(n15862), .Z(n15823) );
  NAND U17452 ( .A(A[0]), .B(B[271]), .Z(n15862) );
  NAND U17453 ( .A(B[270]), .B(A[1]), .Z(n15826) );
  NAND U17454 ( .A(n15863), .B(n15864), .Z(n1649) );
  NANDN U17455 ( .A(n15865), .B(n15866), .Z(n15864) );
  OR U17456 ( .A(n15867), .B(n15868), .Z(n15866) );
  NAND U17457 ( .A(n15868), .B(n15867), .Z(n15863) );
  XOR U17458 ( .A(n1653), .B(n1652), .Z(\A1[268] ) );
  XOR U17459 ( .A(n15868), .B(n15869), .Z(n1652) );
  XNOR U17460 ( .A(n15867), .B(n15865), .Z(n15869) );
  AND U17461 ( .A(n15870), .B(n15871), .Z(n15865) );
  NANDN U17462 ( .A(n15872), .B(n15873), .Z(n15871) );
  NANDN U17463 ( .A(n15874), .B(n15875), .Z(n15873) );
  AND U17464 ( .A(B[267]), .B(A[3]), .Z(n15867) );
  XNOR U17465 ( .A(n15857), .B(n15876), .Z(n15868) );
  XNOR U17466 ( .A(n15855), .B(n15858), .Z(n15876) );
  NAND U17467 ( .A(A[2]), .B(B[268]), .Z(n15858) );
  NANDN U17468 ( .A(n15877), .B(n15878), .Z(n15855) );
  AND U17469 ( .A(A[0]), .B(B[269]), .Z(n15878) );
  XOR U17470 ( .A(n15860), .B(n15879), .Z(n15857) );
  NAND U17471 ( .A(A[0]), .B(B[270]), .Z(n15879) );
  NAND U17472 ( .A(B[269]), .B(A[1]), .Z(n15860) );
  NAND U17473 ( .A(n15880), .B(n15881), .Z(n1653) );
  NANDN U17474 ( .A(n15882), .B(n15883), .Z(n15881) );
  OR U17475 ( .A(n15884), .B(n15885), .Z(n15883) );
  NAND U17476 ( .A(n15885), .B(n15884), .Z(n15880) );
  XOR U17477 ( .A(n1655), .B(n1654), .Z(\A1[267] ) );
  XOR U17478 ( .A(n15885), .B(n15886), .Z(n1654) );
  XNOR U17479 ( .A(n15884), .B(n15882), .Z(n15886) );
  AND U17480 ( .A(n15887), .B(n15888), .Z(n15882) );
  NANDN U17481 ( .A(n15889), .B(n15890), .Z(n15888) );
  NANDN U17482 ( .A(n15891), .B(n15892), .Z(n15890) );
  AND U17483 ( .A(B[266]), .B(A[3]), .Z(n15884) );
  XNOR U17484 ( .A(n15874), .B(n15893), .Z(n15885) );
  XNOR U17485 ( .A(n15872), .B(n15875), .Z(n15893) );
  NAND U17486 ( .A(A[2]), .B(B[267]), .Z(n15875) );
  NANDN U17487 ( .A(n15894), .B(n15895), .Z(n15872) );
  AND U17488 ( .A(A[0]), .B(B[268]), .Z(n15895) );
  XOR U17489 ( .A(n15877), .B(n15896), .Z(n15874) );
  NAND U17490 ( .A(A[0]), .B(B[269]), .Z(n15896) );
  NAND U17491 ( .A(B[268]), .B(A[1]), .Z(n15877) );
  NAND U17492 ( .A(n15897), .B(n15898), .Z(n1655) );
  NANDN U17493 ( .A(n15899), .B(n15900), .Z(n15898) );
  OR U17494 ( .A(n15901), .B(n15902), .Z(n15900) );
  NAND U17495 ( .A(n15902), .B(n15901), .Z(n15897) );
  XOR U17496 ( .A(n1657), .B(n1656), .Z(\A1[266] ) );
  XOR U17497 ( .A(n15902), .B(n15903), .Z(n1656) );
  XNOR U17498 ( .A(n15901), .B(n15899), .Z(n15903) );
  AND U17499 ( .A(n15904), .B(n15905), .Z(n15899) );
  NANDN U17500 ( .A(n15906), .B(n15907), .Z(n15905) );
  NANDN U17501 ( .A(n15908), .B(n15909), .Z(n15907) );
  AND U17502 ( .A(B[265]), .B(A[3]), .Z(n15901) );
  XNOR U17503 ( .A(n15891), .B(n15910), .Z(n15902) );
  XNOR U17504 ( .A(n15889), .B(n15892), .Z(n15910) );
  NAND U17505 ( .A(A[2]), .B(B[266]), .Z(n15892) );
  NANDN U17506 ( .A(n15911), .B(n15912), .Z(n15889) );
  AND U17507 ( .A(A[0]), .B(B[267]), .Z(n15912) );
  XOR U17508 ( .A(n15894), .B(n15913), .Z(n15891) );
  NAND U17509 ( .A(A[0]), .B(B[268]), .Z(n15913) );
  NAND U17510 ( .A(B[267]), .B(A[1]), .Z(n15894) );
  NAND U17511 ( .A(n15914), .B(n15915), .Z(n1657) );
  NANDN U17512 ( .A(n15916), .B(n15917), .Z(n15915) );
  OR U17513 ( .A(n15918), .B(n15919), .Z(n15917) );
  NAND U17514 ( .A(n15919), .B(n15918), .Z(n15914) );
  XOR U17515 ( .A(n1659), .B(n1658), .Z(\A1[265] ) );
  XOR U17516 ( .A(n15919), .B(n15920), .Z(n1658) );
  XNOR U17517 ( .A(n15918), .B(n15916), .Z(n15920) );
  AND U17518 ( .A(n15921), .B(n15922), .Z(n15916) );
  NANDN U17519 ( .A(n15923), .B(n15924), .Z(n15922) );
  NANDN U17520 ( .A(n15925), .B(n15926), .Z(n15924) );
  AND U17521 ( .A(B[264]), .B(A[3]), .Z(n15918) );
  XNOR U17522 ( .A(n15908), .B(n15927), .Z(n15919) );
  XNOR U17523 ( .A(n15906), .B(n15909), .Z(n15927) );
  NAND U17524 ( .A(A[2]), .B(B[265]), .Z(n15909) );
  NANDN U17525 ( .A(n15928), .B(n15929), .Z(n15906) );
  AND U17526 ( .A(A[0]), .B(B[266]), .Z(n15929) );
  XOR U17527 ( .A(n15911), .B(n15930), .Z(n15908) );
  NAND U17528 ( .A(A[0]), .B(B[267]), .Z(n15930) );
  NAND U17529 ( .A(B[266]), .B(A[1]), .Z(n15911) );
  NAND U17530 ( .A(n15931), .B(n15932), .Z(n1659) );
  NANDN U17531 ( .A(n15933), .B(n15934), .Z(n15932) );
  OR U17532 ( .A(n15935), .B(n15936), .Z(n15934) );
  NAND U17533 ( .A(n15936), .B(n15935), .Z(n15931) );
  XOR U17534 ( .A(n1661), .B(n1660), .Z(\A1[264] ) );
  XOR U17535 ( .A(n15936), .B(n15937), .Z(n1660) );
  XNOR U17536 ( .A(n15935), .B(n15933), .Z(n15937) );
  AND U17537 ( .A(n15938), .B(n15939), .Z(n15933) );
  NANDN U17538 ( .A(n15940), .B(n15941), .Z(n15939) );
  NANDN U17539 ( .A(n15942), .B(n15943), .Z(n15941) );
  AND U17540 ( .A(B[263]), .B(A[3]), .Z(n15935) );
  XNOR U17541 ( .A(n15925), .B(n15944), .Z(n15936) );
  XNOR U17542 ( .A(n15923), .B(n15926), .Z(n15944) );
  NAND U17543 ( .A(A[2]), .B(B[264]), .Z(n15926) );
  NANDN U17544 ( .A(n15945), .B(n15946), .Z(n15923) );
  AND U17545 ( .A(A[0]), .B(B[265]), .Z(n15946) );
  XOR U17546 ( .A(n15928), .B(n15947), .Z(n15925) );
  NAND U17547 ( .A(A[0]), .B(B[266]), .Z(n15947) );
  NAND U17548 ( .A(B[265]), .B(A[1]), .Z(n15928) );
  NAND U17549 ( .A(n15948), .B(n15949), .Z(n1661) );
  NANDN U17550 ( .A(n15950), .B(n15951), .Z(n15949) );
  OR U17551 ( .A(n15952), .B(n15953), .Z(n15951) );
  NAND U17552 ( .A(n15953), .B(n15952), .Z(n15948) );
  XOR U17553 ( .A(n1663), .B(n1662), .Z(\A1[263] ) );
  XOR U17554 ( .A(n15953), .B(n15954), .Z(n1662) );
  XNOR U17555 ( .A(n15952), .B(n15950), .Z(n15954) );
  AND U17556 ( .A(n15955), .B(n15956), .Z(n15950) );
  NANDN U17557 ( .A(n15957), .B(n15958), .Z(n15956) );
  NANDN U17558 ( .A(n15959), .B(n15960), .Z(n15958) );
  AND U17559 ( .A(B[262]), .B(A[3]), .Z(n15952) );
  XNOR U17560 ( .A(n15942), .B(n15961), .Z(n15953) );
  XNOR U17561 ( .A(n15940), .B(n15943), .Z(n15961) );
  NAND U17562 ( .A(A[2]), .B(B[263]), .Z(n15943) );
  NANDN U17563 ( .A(n15962), .B(n15963), .Z(n15940) );
  AND U17564 ( .A(A[0]), .B(B[264]), .Z(n15963) );
  XOR U17565 ( .A(n15945), .B(n15964), .Z(n15942) );
  NAND U17566 ( .A(A[0]), .B(B[265]), .Z(n15964) );
  NAND U17567 ( .A(B[264]), .B(A[1]), .Z(n15945) );
  NAND U17568 ( .A(n15965), .B(n15966), .Z(n1663) );
  NANDN U17569 ( .A(n15967), .B(n15968), .Z(n15966) );
  OR U17570 ( .A(n15969), .B(n15970), .Z(n15968) );
  NAND U17571 ( .A(n15970), .B(n15969), .Z(n15965) );
  XOR U17572 ( .A(n1665), .B(n1664), .Z(\A1[262] ) );
  XOR U17573 ( .A(n15970), .B(n15971), .Z(n1664) );
  XNOR U17574 ( .A(n15969), .B(n15967), .Z(n15971) );
  AND U17575 ( .A(n15972), .B(n15973), .Z(n15967) );
  NANDN U17576 ( .A(n15974), .B(n15975), .Z(n15973) );
  NANDN U17577 ( .A(n15976), .B(n15977), .Z(n15975) );
  AND U17578 ( .A(B[261]), .B(A[3]), .Z(n15969) );
  XNOR U17579 ( .A(n15959), .B(n15978), .Z(n15970) );
  XNOR U17580 ( .A(n15957), .B(n15960), .Z(n15978) );
  NAND U17581 ( .A(A[2]), .B(B[262]), .Z(n15960) );
  NANDN U17582 ( .A(n15979), .B(n15980), .Z(n15957) );
  AND U17583 ( .A(A[0]), .B(B[263]), .Z(n15980) );
  XOR U17584 ( .A(n15962), .B(n15981), .Z(n15959) );
  NAND U17585 ( .A(A[0]), .B(B[264]), .Z(n15981) );
  NAND U17586 ( .A(B[263]), .B(A[1]), .Z(n15962) );
  NAND U17587 ( .A(n15982), .B(n15983), .Z(n1665) );
  NANDN U17588 ( .A(n15984), .B(n15985), .Z(n15983) );
  OR U17589 ( .A(n15986), .B(n15987), .Z(n15985) );
  NAND U17590 ( .A(n15987), .B(n15986), .Z(n15982) );
  XOR U17591 ( .A(n1667), .B(n1666), .Z(\A1[261] ) );
  XOR U17592 ( .A(n15987), .B(n15988), .Z(n1666) );
  XNOR U17593 ( .A(n15986), .B(n15984), .Z(n15988) );
  AND U17594 ( .A(n15989), .B(n15990), .Z(n15984) );
  NANDN U17595 ( .A(n15991), .B(n15992), .Z(n15990) );
  NANDN U17596 ( .A(n15993), .B(n15994), .Z(n15992) );
  AND U17597 ( .A(B[260]), .B(A[3]), .Z(n15986) );
  XNOR U17598 ( .A(n15976), .B(n15995), .Z(n15987) );
  XNOR U17599 ( .A(n15974), .B(n15977), .Z(n15995) );
  NAND U17600 ( .A(A[2]), .B(B[261]), .Z(n15977) );
  NANDN U17601 ( .A(n15996), .B(n15997), .Z(n15974) );
  AND U17602 ( .A(A[0]), .B(B[262]), .Z(n15997) );
  XOR U17603 ( .A(n15979), .B(n15998), .Z(n15976) );
  NAND U17604 ( .A(A[0]), .B(B[263]), .Z(n15998) );
  NAND U17605 ( .A(B[262]), .B(A[1]), .Z(n15979) );
  NAND U17606 ( .A(n15999), .B(n16000), .Z(n1667) );
  NANDN U17607 ( .A(n16001), .B(n16002), .Z(n16000) );
  OR U17608 ( .A(n16003), .B(n16004), .Z(n16002) );
  NAND U17609 ( .A(n16004), .B(n16003), .Z(n15999) );
  XOR U17610 ( .A(n1669), .B(n1668), .Z(\A1[260] ) );
  XOR U17611 ( .A(n16004), .B(n16005), .Z(n1668) );
  XNOR U17612 ( .A(n16003), .B(n16001), .Z(n16005) );
  AND U17613 ( .A(n16006), .B(n16007), .Z(n16001) );
  NANDN U17614 ( .A(n16008), .B(n16009), .Z(n16007) );
  NANDN U17615 ( .A(n16010), .B(n16011), .Z(n16009) );
  AND U17616 ( .A(B[259]), .B(A[3]), .Z(n16003) );
  XNOR U17617 ( .A(n15993), .B(n16012), .Z(n16004) );
  XNOR U17618 ( .A(n15991), .B(n15994), .Z(n16012) );
  NAND U17619 ( .A(A[2]), .B(B[260]), .Z(n15994) );
  NANDN U17620 ( .A(n16013), .B(n16014), .Z(n15991) );
  AND U17621 ( .A(A[0]), .B(B[261]), .Z(n16014) );
  XOR U17622 ( .A(n15996), .B(n16015), .Z(n15993) );
  NAND U17623 ( .A(A[0]), .B(B[262]), .Z(n16015) );
  NAND U17624 ( .A(B[261]), .B(A[1]), .Z(n15996) );
  NAND U17625 ( .A(n16016), .B(n16017), .Z(n1669) );
  NANDN U17626 ( .A(n16018), .B(n16019), .Z(n16017) );
  OR U17627 ( .A(n16020), .B(n16021), .Z(n16019) );
  NAND U17628 ( .A(n16021), .B(n16020), .Z(n16016) );
  XOR U17629 ( .A(n1651), .B(n1650), .Z(\A1[25] ) );
  XOR U17630 ( .A(n15851), .B(n16022), .Z(n1650) );
  XNOR U17631 ( .A(n15850), .B(n15848), .Z(n16022) );
  AND U17632 ( .A(n16023), .B(n16024), .Z(n15848) );
  NANDN U17633 ( .A(n16025), .B(n16026), .Z(n16024) );
  NANDN U17634 ( .A(n16027), .B(n16028), .Z(n16026) );
  AND U17635 ( .A(B[24]), .B(A[3]), .Z(n15850) );
  XNOR U17636 ( .A(n15840), .B(n16029), .Z(n15851) );
  XNOR U17637 ( .A(n15838), .B(n15841), .Z(n16029) );
  NAND U17638 ( .A(A[2]), .B(B[25]), .Z(n15841) );
  NANDN U17639 ( .A(n16030), .B(n16031), .Z(n15838) );
  AND U17640 ( .A(A[0]), .B(B[26]), .Z(n16031) );
  XOR U17641 ( .A(n15843), .B(n16032), .Z(n15840) );
  NAND U17642 ( .A(A[0]), .B(B[27]), .Z(n16032) );
  NAND U17643 ( .A(B[26]), .B(A[1]), .Z(n15843) );
  NAND U17644 ( .A(n16033), .B(n16034), .Z(n1651) );
  NANDN U17645 ( .A(n16035), .B(n16036), .Z(n16034) );
  OR U17646 ( .A(n16037), .B(n16038), .Z(n16036) );
  NAND U17647 ( .A(n16038), .B(n16037), .Z(n16033) );
  XOR U17648 ( .A(n1671), .B(n1670), .Z(\A1[259] ) );
  XOR U17649 ( .A(n16021), .B(n16039), .Z(n1670) );
  XNOR U17650 ( .A(n16020), .B(n16018), .Z(n16039) );
  AND U17651 ( .A(n16040), .B(n16041), .Z(n16018) );
  NANDN U17652 ( .A(n16042), .B(n16043), .Z(n16041) );
  NANDN U17653 ( .A(n16044), .B(n16045), .Z(n16043) );
  AND U17654 ( .A(B[258]), .B(A[3]), .Z(n16020) );
  XNOR U17655 ( .A(n16010), .B(n16046), .Z(n16021) );
  XNOR U17656 ( .A(n16008), .B(n16011), .Z(n16046) );
  NAND U17657 ( .A(A[2]), .B(B[259]), .Z(n16011) );
  NANDN U17658 ( .A(n16047), .B(n16048), .Z(n16008) );
  AND U17659 ( .A(A[0]), .B(B[260]), .Z(n16048) );
  XOR U17660 ( .A(n16013), .B(n16049), .Z(n16010) );
  NAND U17661 ( .A(A[0]), .B(B[261]), .Z(n16049) );
  NAND U17662 ( .A(B[260]), .B(A[1]), .Z(n16013) );
  NAND U17663 ( .A(n16050), .B(n16051), .Z(n1671) );
  NANDN U17664 ( .A(n16052), .B(n16053), .Z(n16051) );
  OR U17665 ( .A(n16054), .B(n16055), .Z(n16053) );
  NAND U17666 ( .A(n16055), .B(n16054), .Z(n16050) );
  XOR U17667 ( .A(n1675), .B(n1674), .Z(\A1[258] ) );
  XOR U17668 ( .A(n16055), .B(n16056), .Z(n1674) );
  XNOR U17669 ( .A(n16054), .B(n16052), .Z(n16056) );
  AND U17670 ( .A(n16057), .B(n16058), .Z(n16052) );
  NANDN U17671 ( .A(n16059), .B(n16060), .Z(n16058) );
  NANDN U17672 ( .A(n16061), .B(n16062), .Z(n16060) );
  AND U17673 ( .A(B[257]), .B(A[3]), .Z(n16054) );
  XNOR U17674 ( .A(n16044), .B(n16063), .Z(n16055) );
  XNOR U17675 ( .A(n16042), .B(n16045), .Z(n16063) );
  NAND U17676 ( .A(A[2]), .B(B[258]), .Z(n16045) );
  NANDN U17677 ( .A(n16064), .B(n16065), .Z(n16042) );
  AND U17678 ( .A(A[0]), .B(B[259]), .Z(n16065) );
  XOR U17679 ( .A(n16047), .B(n16066), .Z(n16044) );
  NAND U17680 ( .A(A[0]), .B(B[260]), .Z(n16066) );
  NAND U17681 ( .A(B[259]), .B(A[1]), .Z(n16047) );
  NAND U17682 ( .A(n16067), .B(n16068), .Z(n1675) );
  NANDN U17683 ( .A(n16069), .B(n16070), .Z(n16068) );
  OR U17684 ( .A(n16071), .B(n16072), .Z(n16070) );
  NAND U17685 ( .A(n16072), .B(n16071), .Z(n16067) );
  XOR U17686 ( .A(n1677), .B(n1676), .Z(\A1[257] ) );
  XOR U17687 ( .A(n16072), .B(n16073), .Z(n1676) );
  XNOR U17688 ( .A(n16071), .B(n16069), .Z(n16073) );
  AND U17689 ( .A(n16074), .B(n16075), .Z(n16069) );
  NANDN U17690 ( .A(n16076), .B(n16077), .Z(n16075) );
  NANDN U17691 ( .A(n16078), .B(n16079), .Z(n16077) );
  AND U17692 ( .A(B[256]), .B(A[3]), .Z(n16071) );
  XNOR U17693 ( .A(n16061), .B(n16080), .Z(n16072) );
  XNOR U17694 ( .A(n16059), .B(n16062), .Z(n16080) );
  NAND U17695 ( .A(A[2]), .B(B[257]), .Z(n16062) );
  NANDN U17696 ( .A(n16081), .B(n16082), .Z(n16059) );
  AND U17697 ( .A(A[0]), .B(B[258]), .Z(n16082) );
  XOR U17698 ( .A(n16064), .B(n16083), .Z(n16061) );
  NAND U17699 ( .A(A[0]), .B(B[259]), .Z(n16083) );
  NAND U17700 ( .A(B[258]), .B(A[1]), .Z(n16064) );
  NAND U17701 ( .A(n16084), .B(n16085), .Z(n1677) );
  NANDN U17702 ( .A(n16086), .B(n16087), .Z(n16085) );
  OR U17703 ( .A(n16088), .B(n16089), .Z(n16087) );
  NAND U17704 ( .A(n16089), .B(n16088), .Z(n16084) );
  XOR U17705 ( .A(n1679), .B(n1678), .Z(\A1[256] ) );
  XOR U17706 ( .A(n16089), .B(n16090), .Z(n1678) );
  XNOR U17707 ( .A(n16088), .B(n16086), .Z(n16090) );
  AND U17708 ( .A(n16091), .B(n16092), .Z(n16086) );
  NANDN U17709 ( .A(n16093), .B(n16094), .Z(n16092) );
  NANDN U17710 ( .A(n16095), .B(n16096), .Z(n16094) );
  AND U17711 ( .A(B[255]), .B(A[3]), .Z(n16088) );
  XNOR U17712 ( .A(n16078), .B(n16097), .Z(n16089) );
  XNOR U17713 ( .A(n16076), .B(n16079), .Z(n16097) );
  NAND U17714 ( .A(A[2]), .B(B[256]), .Z(n16079) );
  NANDN U17715 ( .A(n16098), .B(n16099), .Z(n16076) );
  AND U17716 ( .A(A[0]), .B(B[257]), .Z(n16099) );
  XOR U17717 ( .A(n16081), .B(n16100), .Z(n16078) );
  NAND U17718 ( .A(A[0]), .B(B[258]), .Z(n16100) );
  NAND U17719 ( .A(B[257]), .B(A[1]), .Z(n16081) );
  NAND U17720 ( .A(n16101), .B(n16102), .Z(n1679) );
  NANDN U17721 ( .A(n16103), .B(n16104), .Z(n16102) );
  OR U17722 ( .A(n16105), .B(n16106), .Z(n16104) );
  NAND U17723 ( .A(n16106), .B(n16105), .Z(n16101) );
  XOR U17724 ( .A(n1681), .B(n1680), .Z(\A1[255] ) );
  XOR U17725 ( .A(n16106), .B(n16107), .Z(n1680) );
  XNOR U17726 ( .A(n16105), .B(n16103), .Z(n16107) );
  AND U17727 ( .A(n16108), .B(n16109), .Z(n16103) );
  NANDN U17728 ( .A(n16110), .B(n16111), .Z(n16109) );
  NANDN U17729 ( .A(n16112), .B(n16113), .Z(n16111) );
  AND U17730 ( .A(B[254]), .B(A[3]), .Z(n16105) );
  XNOR U17731 ( .A(n16095), .B(n16114), .Z(n16106) );
  XNOR U17732 ( .A(n16093), .B(n16096), .Z(n16114) );
  NAND U17733 ( .A(A[2]), .B(B[255]), .Z(n16096) );
  NANDN U17734 ( .A(n16115), .B(n16116), .Z(n16093) );
  AND U17735 ( .A(A[0]), .B(B[256]), .Z(n16116) );
  XOR U17736 ( .A(n16098), .B(n16117), .Z(n16095) );
  NAND U17737 ( .A(A[0]), .B(B[257]), .Z(n16117) );
  NAND U17738 ( .A(B[256]), .B(A[1]), .Z(n16098) );
  NAND U17739 ( .A(n16118), .B(n16119), .Z(n1681) );
  NANDN U17740 ( .A(n16120), .B(n16121), .Z(n16119) );
  OR U17741 ( .A(n16122), .B(n16123), .Z(n16121) );
  NAND U17742 ( .A(n16123), .B(n16122), .Z(n16118) );
  XOR U17743 ( .A(n1683), .B(n1682), .Z(\A1[254] ) );
  XOR U17744 ( .A(n16123), .B(n16124), .Z(n1682) );
  XNOR U17745 ( .A(n16122), .B(n16120), .Z(n16124) );
  AND U17746 ( .A(n16125), .B(n16126), .Z(n16120) );
  NANDN U17747 ( .A(n16127), .B(n16128), .Z(n16126) );
  NANDN U17748 ( .A(n16129), .B(n16130), .Z(n16128) );
  AND U17749 ( .A(B[253]), .B(A[3]), .Z(n16122) );
  XNOR U17750 ( .A(n16112), .B(n16131), .Z(n16123) );
  XNOR U17751 ( .A(n16110), .B(n16113), .Z(n16131) );
  NAND U17752 ( .A(A[2]), .B(B[254]), .Z(n16113) );
  NANDN U17753 ( .A(n16132), .B(n16133), .Z(n16110) );
  AND U17754 ( .A(A[0]), .B(B[255]), .Z(n16133) );
  XOR U17755 ( .A(n16115), .B(n16134), .Z(n16112) );
  NAND U17756 ( .A(A[0]), .B(B[256]), .Z(n16134) );
  NAND U17757 ( .A(B[255]), .B(A[1]), .Z(n16115) );
  NAND U17758 ( .A(n16135), .B(n16136), .Z(n1683) );
  NANDN U17759 ( .A(n16137), .B(n16138), .Z(n16136) );
  OR U17760 ( .A(n16139), .B(n16140), .Z(n16138) );
  NAND U17761 ( .A(n16140), .B(n16139), .Z(n16135) );
  XOR U17762 ( .A(n1685), .B(n1684), .Z(\A1[253] ) );
  XOR U17763 ( .A(n16140), .B(n16141), .Z(n1684) );
  XNOR U17764 ( .A(n16139), .B(n16137), .Z(n16141) );
  AND U17765 ( .A(n16142), .B(n16143), .Z(n16137) );
  NANDN U17766 ( .A(n16144), .B(n16145), .Z(n16143) );
  NANDN U17767 ( .A(n16146), .B(n16147), .Z(n16145) );
  AND U17768 ( .A(B[252]), .B(A[3]), .Z(n16139) );
  XNOR U17769 ( .A(n16129), .B(n16148), .Z(n16140) );
  XNOR U17770 ( .A(n16127), .B(n16130), .Z(n16148) );
  NAND U17771 ( .A(A[2]), .B(B[253]), .Z(n16130) );
  NANDN U17772 ( .A(n16149), .B(n16150), .Z(n16127) );
  AND U17773 ( .A(A[0]), .B(B[254]), .Z(n16150) );
  XOR U17774 ( .A(n16132), .B(n16151), .Z(n16129) );
  NAND U17775 ( .A(A[0]), .B(B[255]), .Z(n16151) );
  NAND U17776 ( .A(B[254]), .B(A[1]), .Z(n16132) );
  NAND U17777 ( .A(n16152), .B(n16153), .Z(n1685) );
  NANDN U17778 ( .A(n16154), .B(n16155), .Z(n16153) );
  OR U17779 ( .A(n16156), .B(n16157), .Z(n16155) );
  NAND U17780 ( .A(n16157), .B(n16156), .Z(n16152) );
  XOR U17781 ( .A(n1687), .B(n1686), .Z(\A1[252] ) );
  XOR U17782 ( .A(n16157), .B(n16158), .Z(n1686) );
  XNOR U17783 ( .A(n16156), .B(n16154), .Z(n16158) );
  AND U17784 ( .A(n16159), .B(n16160), .Z(n16154) );
  NANDN U17785 ( .A(n16161), .B(n16162), .Z(n16160) );
  NANDN U17786 ( .A(n16163), .B(n16164), .Z(n16162) );
  AND U17787 ( .A(B[251]), .B(A[3]), .Z(n16156) );
  XNOR U17788 ( .A(n16146), .B(n16165), .Z(n16157) );
  XNOR U17789 ( .A(n16144), .B(n16147), .Z(n16165) );
  NAND U17790 ( .A(A[2]), .B(B[252]), .Z(n16147) );
  NANDN U17791 ( .A(n16166), .B(n16167), .Z(n16144) );
  AND U17792 ( .A(A[0]), .B(B[253]), .Z(n16167) );
  XOR U17793 ( .A(n16149), .B(n16168), .Z(n16146) );
  NAND U17794 ( .A(A[0]), .B(B[254]), .Z(n16168) );
  NAND U17795 ( .A(B[253]), .B(A[1]), .Z(n16149) );
  NAND U17796 ( .A(n16169), .B(n16170), .Z(n1687) );
  NANDN U17797 ( .A(n16171), .B(n16172), .Z(n16170) );
  OR U17798 ( .A(n16173), .B(n16174), .Z(n16172) );
  NAND U17799 ( .A(n16174), .B(n16173), .Z(n16169) );
  XOR U17800 ( .A(n1689), .B(n1688), .Z(\A1[251] ) );
  XOR U17801 ( .A(n16174), .B(n16175), .Z(n1688) );
  XNOR U17802 ( .A(n16173), .B(n16171), .Z(n16175) );
  AND U17803 ( .A(n16176), .B(n16177), .Z(n16171) );
  NANDN U17804 ( .A(n16178), .B(n16179), .Z(n16177) );
  NANDN U17805 ( .A(n16180), .B(n16181), .Z(n16179) );
  AND U17806 ( .A(B[250]), .B(A[3]), .Z(n16173) );
  XNOR U17807 ( .A(n16163), .B(n16182), .Z(n16174) );
  XNOR U17808 ( .A(n16161), .B(n16164), .Z(n16182) );
  NAND U17809 ( .A(A[2]), .B(B[251]), .Z(n16164) );
  NANDN U17810 ( .A(n16183), .B(n16184), .Z(n16161) );
  AND U17811 ( .A(A[0]), .B(B[252]), .Z(n16184) );
  XOR U17812 ( .A(n16166), .B(n16185), .Z(n16163) );
  NAND U17813 ( .A(A[0]), .B(B[253]), .Z(n16185) );
  NAND U17814 ( .A(B[252]), .B(A[1]), .Z(n16166) );
  NAND U17815 ( .A(n16186), .B(n16187), .Z(n1689) );
  NANDN U17816 ( .A(n16188), .B(n16189), .Z(n16187) );
  OR U17817 ( .A(n16190), .B(n16191), .Z(n16189) );
  NAND U17818 ( .A(n16191), .B(n16190), .Z(n16186) );
  XOR U17819 ( .A(n1691), .B(n1690), .Z(\A1[250] ) );
  XOR U17820 ( .A(n16191), .B(n16192), .Z(n1690) );
  XNOR U17821 ( .A(n16190), .B(n16188), .Z(n16192) );
  AND U17822 ( .A(n16193), .B(n16194), .Z(n16188) );
  NANDN U17823 ( .A(n16195), .B(n16196), .Z(n16194) );
  NANDN U17824 ( .A(n16197), .B(n16198), .Z(n16196) );
  AND U17825 ( .A(B[249]), .B(A[3]), .Z(n16190) );
  XNOR U17826 ( .A(n16180), .B(n16199), .Z(n16191) );
  XNOR U17827 ( .A(n16178), .B(n16181), .Z(n16199) );
  NAND U17828 ( .A(A[2]), .B(B[250]), .Z(n16181) );
  NANDN U17829 ( .A(n16200), .B(n16201), .Z(n16178) );
  AND U17830 ( .A(A[0]), .B(B[251]), .Z(n16201) );
  XOR U17831 ( .A(n16183), .B(n16202), .Z(n16180) );
  NAND U17832 ( .A(A[0]), .B(B[252]), .Z(n16202) );
  NAND U17833 ( .A(B[251]), .B(A[1]), .Z(n16183) );
  NAND U17834 ( .A(n16203), .B(n16204), .Z(n1691) );
  NANDN U17835 ( .A(n16205), .B(n16206), .Z(n16204) );
  OR U17836 ( .A(n16207), .B(n16208), .Z(n16206) );
  NAND U17837 ( .A(n16208), .B(n16207), .Z(n16203) );
  XOR U17838 ( .A(n1673), .B(n1672), .Z(\A1[24] ) );
  XOR U17839 ( .A(n16038), .B(n16209), .Z(n1672) );
  XNOR U17840 ( .A(n16037), .B(n16035), .Z(n16209) );
  AND U17841 ( .A(n16210), .B(n16211), .Z(n16035) );
  NANDN U17842 ( .A(n16212), .B(n16213), .Z(n16211) );
  NANDN U17843 ( .A(n16214), .B(n16215), .Z(n16213) );
  AND U17844 ( .A(B[23]), .B(A[3]), .Z(n16037) );
  XNOR U17845 ( .A(n16027), .B(n16216), .Z(n16038) );
  XNOR U17846 ( .A(n16025), .B(n16028), .Z(n16216) );
  NAND U17847 ( .A(A[2]), .B(B[24]), .Z(n16028) );
  NANDN U17848 ( .A(n16217), .B(n16218), .Z(n16025) );
  AND U17849 ( .A(A[0]), .B(B[25]), .Z(n16218) );
  XOR U17850 ( .A(n16030), .B(n16219), .Z(n16027) );
  NAND U17851 ( .A(A[0]), .B(B[26]), .Z(n16219) );
  NAND U17852 ( .A(B[25]), .B(A[1]), .Z(n16030) );
  NAND U17853 ( .A(n16220), .B(n16221), .Z(n1673) );
  NANDN U17854 ( .A(n16222), .B(n16223), .Z(n16221) );
  OR U17855 ( .A(n16224), .B(n16225), .Z(n16223) );
  NAND U17856 ( .A(n16225), .B(n16224), .Z(n16220) );
  XOR U17857 ( .A(n1693), .B(n1692), .Z(\A1[249] ) );
  XOR U17858 ( .A(n16208), .B(n16226), .Z(n1692) );
  XNOR U17859 ( .A(n16207), .B(n16205), .Z(n16226) );
  AND U17860 ( .A(n16227), .B(n16228), .Z(n16205) );
  NANDN U17861 ( .A(n16229), .B(n16230), .Z(n16228) );
  NANDN U17862 ( .A(n16231), .B(n16232), .Z(n16230) );
  AND U17863 ( .A(B[248]), .B(A[3]), .Z(n16207) );
  XNOR U17864 ( .A(n16197), .B(n16233), .Z(n16208) );
  XNOR U17865 ( .A(n16195), .B(n16198), .Z(n16233) );
  NAND U17866 ( .A(A[2]), .B(B[249]), .Z(n16198) );
  NANDN U17867 ( .A(n16234), .B(n16235), .Z(n16195) );
  AND U17868 ( .A(A[0]), .B(B[250]), .Z(n16235) );
  XOR U17869 ( .A(n16200), .B(n16236), .Z(n16197) );
  NAND U17870 ( .A(A[0]), .B(B[251]), .Z(n16236) );
  NAND U17871 ( .A(B[250]), .B(A[1]), .Z(n16200) );
  NAND U17872 ( .A(n16237), .B(n16238), .Z(n1693) );
  NANDN U17873 ( .A(n16239), .B(n16240), .Z(n16238) );
  OR U17874 ( .A(n16241), .B(n16242), .Z(n16240) );
  NAND U17875 ( .A(n16242), .B(n16241), .Z(n16237) );
  XOR U17876 ( .A(n1697), .B(n1696), .Z(\A1[248] ) );
  XOR U17877 ( .A(n16242), .B(n16243), .Z(n1696) );
  XNOR U17878 ( .A(n16241), .B(n16239), .Z(n16243) );
  AND U17879 ( .A(n16244), .B(n16245), .Z(n16239) );
  NANDN U17880 ( .A(n16246), .B(n16247), .Z(n16245) );
  NANDN U17881 ( .A(n16248), .B(n16249), .Z(n16247) );
  AND U17882 ( .A(B[247]), .B(A[3]), .Z(n16241) );
  XNOR U17883 ( .A(n16231), .B(n16250), .Z(n16242) );
  XNOR U17884 ( .A(n16229), .B(n16232), .Z(n16250) );
  NAND U17885 ( .A(A[2]), .B(B[248]), .Z(n16232) );
  NANDN U17886 ( .A(n16251), .B(n16252), .Z(n16229) );
  AND U17887 ( .A(A[0]), .B(B[249]), .Z(n16252) );
  XOR U17888 ( .A(n16234), .B(n16253), .Z(n16231) );
  NAND U17889 ( .A(A[0]), .B(B[250]), .Z(n16253) );
  NAND U17890 ( .A(B[249]), .B(A[1]), .Z(n16234) );
  NAND U17891 ( .A(n16254), .B(n16255), .Z(n1697) );
  NANDN U17892 ( .A(n16256), .B(n16257), .Z(n16255) );
  OR U17893 ( .A(n16258), .B(n16259), .Z(n16257) );
  NAND U17894 ( .A(n16259), .B(n16258), .Z(n16254) );
  XOR U17895 ( .A(n1699), .B(n1698), .Z(\A1[247] ) );
  XOR U17896 ( .A(n16259), .B(n16260), .Z(n1698) );
  XNOR U17897 ( .A(n16258), .B(n16256), .Z(n16260) );
  AND U17898 ( .A(n16261), .B(n16262), .Z(n16256) );
  NANDN U17899 ( .A(n16263), .B(n16264), .Z(n16262) );
  NANDN U17900 ( .A(n16265), .B(n16266), .Z(n16264) );
  AND U17901 ( .A(B[246]), .B(A[3]), .Z(n16258) );
  XNOR U17902 ( .A(n16248), .B(n16267), .Z(n16259) );
  XNOR U17903 ( .A(n16246), .B(n16249), .Z(n16267) );
  NAND U17904 ( .A(A[2]), .B(B[247]), .Z(n16249) );
  NANDN U17905 ( .A(n16268), .B(n16269), .Z(n16246) );
  AND U17906 ( .A(A[0]), .B(B[248]), .Z(n16269) );
  XOR U17907 ( .A(n16251), .B(n16270), .Z(n16248) );
  NAND U17908 ( .A(A[0]), .B(B[249]), .Z(n16270) );
  NAND U17909 ( .A(B[248]), .B(A[1]), .Z(n16251) );
  NAND U17910 ( .A(n16271), .B(n16272), .Z(n1699) );
  NANDN U17911 ( .A(n16273), .B(n16274), .Z(n16272) );
  OR U17912 ( .A(n16275), .B(n16276), .Z(n16274) );
  NAND U17913 ( .A(n16276), .B(n16275), .Z(n16271) );
  XOR U17914 ( .A(n1701), .B(n1700), .Z(\A1[246] ) );
  XOR U17915 ( .A(n16276), .B(n16277), .Z(n1700) );
  XNOR U17916 ( .A(n16275), .B(n16273), .Z(n16277) );
  AND U17917 ( .A(n16278), .B(n16279), .Z(n16273) );
  NANDN U17918 ( .A(n16280), .B(n16281), .Z(n16279) );
  NANDN U17919 ( .A(n16282), .B(n16283), .Z(n16281) );
  AND U17920 ( .A(B[245]), .B(A[3]), .Z(n16275) );
  XNOR U17921 ( .A(n16265), .B(n16284), .Z(n16276) );
  XNOR U17922 ( .A(n16263), .B(n16266), .Z(n16284) );
  NAND U17923 ( .A(A[2]), .B(B[246]), .Z(n16266) );
  NANDN U17924 ( .A(n16285), .B(n16286), .Z(n16263) );
  AND U17925 ( .A(A[0]), .B(B[247]), .Z(n16286) );
  XOR U17926 ( .A(n16268), .B(n16287), .Z(n16265) );
  NAND U17927 ( .A(A[0]), .B(B[248]), .Z(n16287) );
  NAND U17928 ( .A(B[247]), .B(A[1]), .Z(n16268) );
  NAND U17929 ( .A(n16288), .B(n16289), .Z(n1701) );
  NANDN U17930 ( .A(n16290), .B(n16291), .Z(n16289) );
  OR U17931 ( .A(n16292), .B(n16293), .Z(n16291) );
  NAND U17932 ( .A(n16293), .B(n16292), .Z(n16288) );
  XOR U17933 ( .A(n1703), .B(n1702), .Z(\A1[245] ) );
  XOR U17934 ( .A(n16293), .B(n16294), .Z(n1702) );
  XNOR U17935 ( .A(n16292), .B(n16290), .Z(n16294) );
  AND U17936 ( .A(n16295), .B(n16296), .Z(n16290) );
  NANDN U17937 ( .A(n16297), .B(n16298), .Z(n16296) );
  NANDN U17938 ( .A(n16299), .B(n16300), .Z(n16298) );
  AND U17939 ( .A(B[244]), .B(A[3]), .Z(n16292) );
  XNOR U17940 ( .A(n16282), .B(n16301), .Z(n16293) );
  XNOR U17941 ( .A(n16280), .B(n16283), .Z(n16301) );
  NAND U17942 ( .A(A[2]), .B(B[245]), .Z(n16283) );
  NANDN U17943 ( .A(n16302), .B(n16303), .Z(n16280) );
  AND U17944 ( .A(A[0]), .B(B[246]), .Z(n16303) );
  XOR U17945 ( .A(n16285), .B(n16304), .Z(n16282) );
  NAND U17946 ( .A(A[0]), .B(B[247]), .Z(n16304) );
  NAND U17947 ( .A(B[246]), .B(A[1]), .Z(n16285) );
  NAND U17948 ( .A(n16305), .B(n16306), .Z(n1703) );
  NANDN U17949 ( .A(n16307), .B(n16308), .Z(n16306) );
  OR U17950 ( .A(n16309), .B(n16310), .Z(n16308) );
  NAND U17951 ( .A(n16310), .B(n16309), .Z(n16305) );
  XOR U17952 ( .A(n1705), .B(n1704), .Z(\A1[244] ) );
  XOR U17953 ( .A(n16310), .B(n16311), .Z(n1704) );
  XNOR U17954 ( .A(n16309), .B(n16307), .Z(n16311) );
  AND U17955 ( .A(n16312), .B(n16313), .Z(n16307) );
  NANDN U17956 ( .A(n16314), .B(n16315), .Z(n16313) );
  NANDN U17957 ( .A(n16316), .B(n16317), .Z(n16315) );
  AND U17958 ( .A(B[243]), .B(A[3]), .Z(n16309) );
  XNOR U17959 ( .A(n16299), .B(n16318), .Z(n16310) );
  XNOR U17960 ( .A(n16297), .B(n16300), .Z(n16318) );
  NAND U17961 ( .A(A[2]), .B(B[244]), .Z(n16300) );
  NANDN U17962 ( .A(n16319), .B(n16320), .Z(n16297) );
  AND U17963 ( .A(A[0]), .B(B[245]), .Z(n16320) );
  XOR U17964 ( .A(n16302), .B(n16321), .Z(n16299) );
  NAND U17965 ( .A(A[0]), .B(B[246]), .Z(n16321) );
  NAND U17966 ( .A(B[245]), .B(A[1]), .Z(n16302) );
  NAND U17967 ( .A(n16322), .B(n16323), .Z(n1705) );
  NANDN U17968 ( .A(n16324), .B(n16325), .Z(n16323) );
  OR U17969 ( .A(n16326), .B(n16327), .Z(n16325) );
  NAND U17970 ( .A(n16327), .B(n16326), .Z(n16322) );
  XOR U17971 ( .A(n1707), .B(n1706), .Z(\A1[243] ) );
  XOR U17972 ( .A(n16327), .B(n16328), .Z(n1706) );
  XNOR U17973 ( .A(n16326), .B(n16324), .Z(n16328) );
  AND U17974 ( .A(n16329), .B(n16330), .Z(n16324) );
  NANDN U17975 ( .A(n16331), .B(n16332), .Z(n16330) );
  NANDN U17976 ( .A(n16333), .B(n16334), .Z(n16332) );
  AND U17977 ( .A(B[242]), .B(A[3]), .Z(n16326) );
  XNOR U17978 ( .A(n16316), .B(n16335), .Z(n16327) );
  XNOR U17979 ( .A(n16314), .B(n16317), .Z(n16335) );
  NAND U17980 ( .A(A[2]), .B(B[243]), .Z(n16317) );
  NANDN U17981 ( .A(n16336), .B(n16337), .Z(n16314) );
  AND U17982 ( .A(A[0]), .B(B[244]), .Z(n16337) );
  XOR U17983 ( .A(n16319), .B(n16338), .Z(n16316) );
  NAND U17984 ( .A(A[0]), .B(B[245]), .Z(n16338) );
  NAND U17985 ( .A(B[244]), .B(A[1]), .Z(n16319) );
  NAND U17986 ( .A(n16339), .B(n16340), .Z(n1707) );
  NANDN U17987 ( .A(n16341), .B(n16342), .Z(n16340) );
  OR U17988 ( .A(n16343), .B(n16344), .Z(n16342) );
  NAND U17989 ( .A(n16344), .B(n16343), .Z(n16339) );
  XOR U17990 ( .A(n1709), .B(n1708), .Z(\A1[242] ) );
  XOR U17991 ( .A(n16344), .B(n16345), .Z(n1708) );
  XNOR U17992 ( .A(n16343), .B(n16341), .Z(n16345) );
  AND U17993 ( .A(n16346), .B(n16347), .Z(n16341) );
  NANDN U17994 ( .A(n16348), .B(n16349), .Z(n16347) );
  NANDN U17995 ( .A(n16350), .B(n16351), .Z(n16349) );
  AND U17996 ( .A(B[241]), .B(A[3]), .Z(n16343) );
  XNOR U17997 ( .A(n16333), .B(n16352), .Z(n16344) );
  XNOR U17998 ( .A(n16331), .B(n16334), .Z(n16352) );
  NAND U17999 ( .A(A[2]), .B(B[242]), .Z(n16334) );
  NANDN U18000 ( .A(n16353), .B(n16354), .Z(n16331) );
  AND U18001 ( .A(A[0]), .B(B[243]), .Z(n16354) );
  XOR U18002 ( .A(n16336), .B(n16355), .Z(n16333) );
  NAND U18003 ( .A(A[0]), .B(B[244]), .Z(n16355) );
  NAND U18004 ( .A(B[243]), .B(A[1]), .Z(n16336) );
  NAND U18005 ( .A(n16356), .B(n16357), .Z(n1709) );
  NANDN U18006 ( .A(n16358), .B(n16359), .Z(n16357) );
  OR U18007 ( .A(n16360), .B(n16361), .Z(n16359) );
  NAND U18008 ( .A(n16361), .B(n16360), .Z(n16356) );
  XOR U18009 ( .A(n1711), .B(n1710), .Z(\A1[241] ) );
  XOR U18010 ( .A(n16361), .B(n16362), .Z(n1710) );
  XNOR U18011 ( .A(n16360), .B(n16358), .Z(n16362) );
  AND U18012 ( .A(n16363), .B(n16364), .Z(n16358) );
  NANDN U18013 ( .A(n16365), .B(n16366), .Z(n16364) );
  NANDN U18014 ( .A(n16367), .B(n16368), .Z(n16366) );
  AND U18015 ( .A(B[240]), .B(A[3]), .Z(n16360) );
  XNOR U18016 ( .A(n16350), .B(n16369), .Z(n16361) );
  XNOR U18017 ( .A(n16348), .B(n16351), .Z(n16369) );
  NAND U18018 ( .A(A[2]), .B(B[241]), .Z(n16351) );
  NANDN U18019 ( .A(n16370), .B(n16371), .Z(n16348) );
  AND U18020 ( .A(A[0]), .B(B[242]), .Z(n16371) );
  XOR U18021 ( .A(n16353), .B(n16372), .Z(n16350) );
  NAND U18022 ( .A(A[0]), .B(B[243]), .Z(n16372) );
  NAND U18023 ( .A(B[242]), .B(A[1]), .Z(n16353) );
  NAND U18024 ( .A(n16373), .B(n16374), .Z(n1711) );
  NANDN U18025 ( .A(n16375), .B(n16376), .Z(n16374) );
  OR U18026 ( .A(n16377), .B(n16378), .Z(n16376) );
  NAND U18027 ( .A(n16378), .B(n16377), .Z(n16373) );
  XOR U18028 ( .A(n1713), .B(n1712), .Z(\A1[240] ) );
  XOR U18029 ( .A(n16378), .B(n16379), .Z(n1712) );
  XNOR U18030 ( .A(n16377), .B(n16375), .Z(n16379) );
  AND U18031 ( .A(n16380), .B(n16381), .Z(n16375) );
  NANDN U18032 ( .A(n16382), .B(n16383), .Z(n16381) );
  NANDN U18033 ( .A(n16384), .B(n16385), .Z(n16383) );
  AND U18034 ( .A(B[239]), .B(A[3]), .Z(n16377) );
  XNOR U18035 ( .A(n16367), .B(n16386), .Z(n16378) );
  XNOR U18036 ( .A(n16365), .B(n16368), .Z(n16386) );
  NAND U18037 ( .A(A[2]), .B(B[240]), .Z(n16368) );
  NANDN U18038 ( .A(n16387), .B(n16388), .Z(n16365) );
  AND U18039 ( .A(A[0]), .B(B[241]), .Z(n16388) );
  XOR U18040 ( .A(n16370), .B(n16389), .Z(n16367) );
  NAND U18041 ( .A(A[0]), .B(B[242]), .Z(n16389) );
  NAND U18042 ( .A(B[241]), .B(A[1]), .Z(n16370) );
  NAND U18043 ( .A(n16390), .B(n16391), .Z(n1713) );
  NANDN U18044 ( .A(n16392), .B(n16393), .Z(n16391) );
  OR U18045 ( .A(n16394), .B(n16395), .Z(n16393) );
  NAND U18046 ( .A(n16395), .B(n16394), .Z(n16390) );
  XOR U18047 ( .A(n1695), .B(n1694), .Z(\A1[23] ) );
  XOR U18048 ( .A(n16225), .B(n16396), .Z(n1694) );
  XNOR U18049 ( .A(n16224), .B(n16222), .Z(n16396) );
  AND U18050 ( .A(n16397), .B(n16398), .Z(n16222) );
  NANDN U18051 ( .A(n16399), .B(n16400), .Z(n16398) );
  NANDN U18052 ( .A(n16401), .B(n16402), .Z(n16400) );
  AND U18053 ( .A(B[22]), .B(A[3]), .Z(n16224) );
  XNOR U18054 ( .A(n16214), .B(n16403), .Z(n16225) );
  XNOR U18055 ( .A(n16212), .B(n16215), .Z(n16403) );
  NAND U18056 ( .A(A[2]), .B(B[23]), .Z(n16215) );
  NANDN U18057 ( .A(n16404), .B(n16405), .Z(n16212) );
  AND U18058 ( .A(A[0]), .B(B[24]), .Z(n16405) );
  XOR U18059 ( .A(n16217), .B(n16406), .Z(n16214) );
  NAND U18060 ( .A(A[0]), .B(B[25]), .Z(n16406) );
  NAND U18061 ( .A(B[24]), .B(A[1]), .Z(n16217) );
  NAND U18062 ( .A(n16407), .B(n16408), .Z(n1695) );
  NANDN U18063 ( .A(n16409), .B(n16410), .Z(n16408) );
  OR U18064 ( .A(n16411), .B(n16412), .Z(n16410) );
  NAND U18065 ( .A(n16412), .B(n16411), .Z(n16407) );
  XOR U18066 ( .A(n1715), .B(n1714), .Z(\A1[239] ) );
  XOR U18067 ( .A(n16395), .B(n16413), .Z(n1714) );
  XNOR U18068 ( .A(n16394), .B(n16392), .Z(n16413) );
  AND U18069 ( .A(n16414), .B(n16415), .Z(n16392) );
  NANDN U18070 ( .A(n16416), .B(n16417), .Z(n16415) );
  NANDN U18071 ( .A(n16418), .B(n16419), .Z(n16417) );
  AND U18072 ( .A(B[238]), .B(A[3]), .Z(n16394) );
  XNOR U18073 ( .A(n16384), .B(n16420), .Z(n16395) );
  XNOR U18074 ( .A(n16382), .B(n16385), .Z(n16420) );
  NAND U18075 ( .A(A[2]), .B(B[239]), .Z(n16385) );
  NANDN U18076 ( .A(n16421), .B(n16422), .Z(n16382) );
  AND U18077 ( .A(A[0]), .B(B[240]), .Z(n16422) );
  XOR U18078 ( .A(n16387), .B(n16423), .Z(n16384) );
  NAND U18079 ( .A(A[0]), .B(B[241]), .Z(n16423) );
  NAND U18080 ( .A(B[240]), .B(A[1]), .Z(n16387) );
  NAND U18081 ( .A(n16424), .B(n16425), .Z(n1715) );
  NANDN U18082 ( .A(n16426), .B(n16427), .Z(n16425) );
  OR U18083 ( .A(n16428), .B(n16429), .Z(n16427) );
  NAND U18084 ( .A(n16429), .B(n16428), .Z(n16424) );
  XOR U18085 ( .A(n1719), .B(n1718), .Z(\A1[238] ) );
  XOR U18086 ( .A(n16429), .B(n16430), .Z(n1718) );
  XNOR U18087 ( .A(n16428), .B(n16426), .Z(n16430) );
  AND U18088 ( .A(n16431), .B(n16432), .Z(n16426) );
  NANDN U18089 ( .A(n16433), .B(n16434), .Z(n16432) );
  NANDN U18090 ( .A(n16435), .B(n16436), .Z(n16434) );
  AND U18091 ( .A(B[237]), .B(A[3]), .Z(n16428) );
  XNOR U18092 ( .A(n16418), .B(n16437), .Z(n16429) );
  XNOR U18093 ( .A(n16416), .B(n16419), .Z(n16437) );
  NAND U18094 ( .A(A[2]), .B(B[238]), .Z(n16419) );
  NANDN U18095 ( .A(n16438), .B(n16439), .Z(n16416) );
  AND U18096 ( .A(A[0]), .B(B[239]), .Z(n16439) );
  XOR U18097 ( .A(n16421), .B(n16440), .Z(n16418) );
  NAND U18098 ( .A(A[0]), .B(B[240]), .Z(n16440) );
  NAND U18099 ( .A(B[239]), .B(A[1]), .Z(n16421) );
  NAND U18100 ( .A(n16441), .B(n16442), .Z(n1719) );
  NANDN U18101 ( .A(n16443), .B(n16444), .Z(n16442) );
  OR U18102 ( .A(n16445), .B(n16446), .Z(n16444) );
  NAND U18103 ( .A(n16446), .B(n16445), .Z(n16441) );
  XOR U18104 ( .A(n1721), .B(n1720), .Z(\A1[237] ) );
  XOR U18105 ( .A(n16446), .B(n16447), .Z(n1720) );
  XNOR U18106 ( .A(n16445), .B(n16443), .Z(n16447) );
  AND U18107 ( .A(n16448), .B(n16449), .Z(n16443) );
  NANDN U18108 ( .A(n16450), .B(n16451), .Z(n16449) );
  NANDN U18109 ( .A(n16452), .B(n16453), .Z(n16451) );
  AND U18110 ( .A(B[236]), .B(A[3]), .Z(n16445) );
  XNOR U18111 ( .A(n16435), .B(n16454), .Z(n16446) );
  XNOR U18112 ( .A(n16433), .B(n16436), .Z(n16454) );
  NAND U18113 ( .A(A[2]), .B(B[237]), .Z(n16436) );
  NANDN U18114 ( .A(n16455), .B(n16456), .Z(n16433) );
  AND U18115 ( .A(A[0]), .B(B[238]), .Z(n16456) );
  XOR U18116 ( .A(n16438), .B(n16457), .Z(n16435) );
  NAND U18117 ( .A(A[0]), .B(B[239]), .Z(n16457) );
  NAND U18118 ( .A(B[238]), .B(A[1]), .Z(n16438) );
  NAND U18119 ( .A(n16458), .B(n16459), .Z(n1721) );
  NANDN U18120 ( .A(n16460), .B(n16461), .Z(n16459) );
  OR U18121 ( .A(n16462), .B(n16463), .Z(n16461) );
  NAND U18122 ( .A(n16463), .B(n16462), .Z(n16458) );
  XOR U18123 ( .A(n1723), .B(n1722), .Z(\A1[236] ) );
  XOR U18124 ( .A(n16463), .B(n16464), .Z(n1722) );
  XNOR U18125 ( .A(n16462), .B(n16460), .Z(n16464) );
  AND U18126 ( .A(n16465), .B(n16466), .Z(n16460) );
  NANDN U18127 ( .A(n16467), .B(n16468), .Z(n16466) );
  NANDN U18128 ( .A(n16469), .B(n16470), .Z(n16468) );
  AND U18129 ( .A(B[235]), .B(A[3]), .Z(n16462) );
  XNOR U18130 ( .A(n16452), .B(n16471), .Z(n16463) );
  XNOR U18131 ( .A(n16450), .B(n16453), .Z(n16471) );
  NAND U18132 ( .A(A[2]), .B(B[236]), .Z(n16453) );
  NANDN U18133 ( .A(n16472), .B(n16473), .Z(n16450) );
  AND U18134 ( .A(A[0]), .B(B[237]), .Z(n16473) );
  XOR U18135 ( .A(n16455), .B(n16474), .Z(n16452) );
  NAND U18136 ( .A(A[0]), .B(B[238]), .Z(n16474) );
  NAND U18137 ( .A(B[237]), .B(A[1]), .Z(n16455) );
  NAND U18138 ( .A(n16475), .B(n16476), .Z(n1723) );
  NANDN U18139 ( .A(n16477), .B(n16478), .Z(n16476) );
  OR U18140 ( .A(n16479), .B(n16480), .Z(n16478) );
  NAND U18141 ( .A(n16480), .B(n16479), .Z(n16475) );
  XOR U18142 ( .A(n1725), .B(n1724), .Z(\A1[235] ) );
  XOR U18143 ( .A(n16480), .B(n16481), .Z(n1724) );
  XNOR U18144 ( .A(n16479), .B(n16477), .Z(n16481) );
  AND U18145 ( .A(n16482), .B(n16483), .Z(n16477) );
  NANDN U18146 ( .A(n16484), .B(n16485), .Z(n16483) );
  NANDN U18147 ( .A(n16486), .B(n16487), .Z(n16485) );
  AND U18148 ( .A(B[234]), .B(A[3]), .Z(n16479) );
  XNOR U18149 ( .A(n16469), .B(n16488), .Z(n16480) );
  XNOR U18150 ( .A(n16467), .B(n16470), .Z(n16488) );
  NAND U18151 ( .A(A[2]), .B(B[235]), .Z(n16470) );
  NANDN U18152 ( .A(n16489), .B(n16490), .Z(n16467) );
  AND U18153 ( .A(A[0]), .B(B[236]), .Z(n16490) );
  XOR U18154 ( .A(n16472), .B(n16491), .Z(n16469) );
  NAND U18155 ( .A(A[0]), .B(B[237]), .Z(n16491) );
  NAND U18156 ( .A(B[236]), .B(A[1]), .Z(n16472) );
  NAND U18157 ( .A(n16492), .B(n16493), .Z(n1725) );
  NANDN U18158 ( .A(n16494), .B(n16495), .Z(n16493) );
  OR U18159 ( .A(n16496), .B(n16497), .Z(n16495) );
  NAND U18160 ( .A(n16497), .B(n16496), .Z(n16492) );
  XOR U18161 ( .A(n1727), .B(n1726), .Z(\A1[234] ) );
  XOR U18162 ( .A(n16497), .B(n16498), .Z(n1726) );
  XNOR U18163 ( .A(n16496), .B(n16494), .Z(n16498) );
  AND U18164 ( .A(n16499), .B(n16500), .Z(n16494) );
  NANDN U18165 ( .A(n16501), .B(n16502), .Z(n16500) );
  NANDN U18166 ( .A(n16503), .B(n16504), .Z(n16502) );
  AND U18167 ( .A(B[233]), .B(A[3]), .Z(n16496) );
  XNOR U18168 ( .A(n16486), .B(n16505), .Z(n16497) );
  XNOR U18169 ( .A(n16484), .B(n16487), .Z(n16505) );
  NAND U18170 ( .A(A[2]), .B(B[234]), .Z(n16487) );
  NANDN U18171 ( .A(n16506), .B(n16507), .Z(n16484) );
  AND U18172 ( .A(A[0]), .B(B[235]), .Z(n16507) );
  XOR U18173 ( .A(n16489), .B(n16508), .Z(n16486) );
  NAND U18174 ( .A(A[0]), .B(B[236]), .Z(n16508) );
  NAND U18175 ( .A(B[235]), .B(A[1]), .Z(n16489) );
  NAND U18176 ( .A(n16509), .B(n16510), .Z(n1727) );
  NANDN U18177 ( .A(n16511), .B(n16512), .Z(n16510) );
  OR U18178 ( .A(n16513), .B(n16514), .Z(n16512) );
  NAND U18179 ( .A(n16514), .B(n16513), .Z(n16509) );
  XOR U18180 ( .A(n1729), .B(n1728), .Z(\A1[233] ) );
  XOR U18181 ( .A(n16514), .B(n16515), .Z(n1728) );
  XNOR U18182 ( .A(n16513), .B(n16511), .Z(n16515) );
  AND U18183 ( .A(n16516), .B(n16517), .Z(n16511) );
  NANDN U18184 ( .A(n16518), .B(n16519), .Z(n16517) );
  NANDN U18185 ( .A(n16520), .B(n16521), .Z(n16519) );
  AND U18186 ( .A(B[232]), .B(A[3]), .Z(n16513) );
  XNOR U18187 ( .A(n16503), .B(n16522), .Z(n16514) );
  XNOR U18188 ( .A(n16501), .B(n16504), .Z(n16522) );
  NAND U18189 ( .A(A[2]), .B(B[233]), .Z(n16504) );
  NANDN U18190 ( .A(n16523), .B(n16524), .Z(n16501) );
  AND U18191 ( .A(A[0]), .B(B[234]), .Z(n16524) );
  XOR U18192 ( .A(n16506), .B(n16525), .Z(n16503) );
  NAND U18193 ( .A(A[0]), .B(B[235]), .Z(n16525) );
  NAND U18194 ( .A(B[234]), .B(A[1]), .Z(n16506) );
  NAND U18195 ( .A(n16526), .B(n16527), .Z(n1729) );
  NANDN U18196 ( .A(n16528), .B(n16529), .Z(n16527) );
  OR U18197 ( .A(n16530), .B(n16531), .Z(n16529) );
  NAND U18198 ( .A(n16531), .B(n16530), .Z(n16526) );
  XOR U18199 ( .A(n1731), .B(n1730), .Z(\A1[232] ) );
  XOR U18200 ( .A(n16531), .B(n16532), .Z(n1730) );
  XNOR U18201 ( .A(n16530), .B(n16528), .Z(n16532) );
  AND U18202 ( .A(n16533), .B(n16534), .Z(n16528) );
  NANDN U18203 ( .A(n16535), .B(n16536), .Z(n16534) );
  NANDN U18204 ( .A(n16537), .B(n16538), .Z(n16536) );
  AND U18205 ( .A(B[231]), .B(A[3]), .Z(n16530) );
  XNOR U18206 ( .A(n16520), .B(n16539), .Z(n16531) );
  XNOR U18207 ( .A(n16518), .B(n16521), .Z(n16539) );
  NAND U18208 ( .A(A[2]), .B(B[232]), .Z(n16521) );
  NANDN U18209 ( .A(n16540), .B(n16541), .Z(n16518) );
  AND U18210 ( .A(A[0]), .B(B[233]), .Z(n16541) );
  XOR U18211 ( .A(n16523), .B(n16542), .Z(n16520) );
  NAND U18212 ( .A(A[0]), .B(B[234]), .Z(n16542) );
  NAND U18213 ( .A(B[233]), .B(A[1]), .Z(n16523) );
  NAND U18214 ( .A(n16543), .B(n16544), .Z(n1731) );
  NANDN U18215 ( .A(n16545), .B(n16546), .Z(n16544) );
  OR U18216 ( .A(n16547), .B(n16548), .Z(n16546) );
  NAND U18217 ( .A(n16548), .B(n16547), .Z(n16543) );
  XOR U18218 ( .A(n1733), .B(n1732), .Z(\A1[231] ) );
  XOR U18219 ( .A(n16548), .B(n16549), .Z(n1732) );
  XNOR U18220 ( .A(n16547), .B(n16545), .Z(n16549) );
  AND U18221 ( .A(n16550), .B(n16551), .Z(n16545) );
  NANDN U18222 ( .A(n16552), .B(n16553), .Z(n16551) );
  NANDN U18223 ( .A(n16554), .B(n16555), .Z(n16553) );
  AND U18224 ( .A(B[230]), .B(A[3]), .Z(n16547) );
  XNOR U18225 ( .A(n16537), .B(n16556), .Z(n16548) );
  XNOR U18226 ( .A(n16535), .B(n16538), .Z(n16556) );
  NAND U18227 ( .A(A[2]), .B(B[231]), .Z(n16538) );
  NANDN U18228 ( .A(n16557), .B(n16558), .Z(n16535) );
  AND U18229 ( .A(A[0]), .B(B[232]), .Z(n16558) );
  XOR U18230 ( .A(n16540), .B(n16559), .Z(n16537) );
  NAND U18231 ( .A(A[0]), .B(B[233]), .Z(n16559) );
  NAND U18232 ( .A(B[232]), .B(A[1]), .Z(n16540) );
  NAND U18233 ( .A(n16560), .B(n16561), .Z(n1733) );
  NANDN U18234 ( .A(n16562), .B(n16563), .Z(n16561) );
  OR U18235 ( .A(n16564), .B(n16565), .Z(n16563) );
  NAND U18236 ( .A(n16565), .B(n16564), .Z(n16560) );
  XOR U18237 ( .A(n1735), .B(n1734), .Z(\A1[230] ) );
  XOR U18238 ( .A(n16565), .B(n16566), .Z(n1734) );
  XNOR U18239 ( .A(n16564), .B(n16562), .Z(n16566) );
  AND U18240 ( .A(n16567), .B(n16568), .Z(n16562) );
  NANDN U18241 ( .A(n16569), .B(n16570), .Z(n16568) );
  NANDN U18242 ( .A(n16571), .B(n16572), .Z(n16570) );
  AND U18243 ( .A(B[229]), .B(A[3]), .Z(n16564) );
  XNOR U18244 ( .A(n16554), .B(n16573), .Z(n16565) );
  XNOR U18245 ( .A(n16552), .B(n16555), .Z(n16573) );
  NAND U18246 ( .A(A[2]), .B(B[230]), .Z(n16555) );
  NANDN U18247 ( .A(n16574), .B(n16575), .Z(n16552) );
  AND U18248 ( .A(A[0]), .B(B[231]), .Z(n16575) );
  XOR U18249 ( .A(n16557), .B(n16576), .Z(n16554) );
  NAND U18250 ( .A(A[0]), .B(B[232]), .Z(n16576) );
  NAND U18251 ( .A(B[231]), .B(A[1]), .Z(n16557) );
  NAND U18252 ( .A(n16577), .B(n16578), .Z(n1735) );
  NANDN U18253 ( .A(n16579), .B(n16580), .Z(n16578) );
  OR U18254 ( .A(n16581), .B(n16582), .Z(n16580) );
  NAND U18255 ( .A(n16582), .B(n16581), .Z(n16577) );
  XOR U18256 ( .A(n1717), .B(n1716), .Z(\A1[22] ) );
  XOR U18257 ( .A(n16412), .B(n16583), .Z(n1716) );
  XNOR U18258 ( .A(n16411), .B(n16409), .Z(n16583) );
  AND U18259 ( .A(n16584), .B(n16585), .Z(n16409) );
  NANDN U18260 ( .A(n16586), .B(n16587), .Z(n16585) );
  NANDN U18261 ( .A(n16588), .B(n16589), .Z(n16587) );
  AND U18262 ( .A(B[21]), .B(A[3]), .Z(n16411) );
  XNOR U18263 ( .A(n16401), .B(n16590), .Z(n16412) );
  XNOR U18264 ( .A(n16399), .B(n16402), .Z(n16590) );
  NAND U18265 ( .A(A[2]), .B(B[22]), .Z(n16402) );
  NANDN U18266 ( .A(n16591), .B(n16592), .Z(n16399) );
  AND U18267 ( .A(A[0]), .B(B[23]), .Z(n16592) );
  XOR U18268 ( .A(n16404), .B(n16593), .Z(n16401) );
  NAND U18269 ( .A(A[0]), .B(B[24]), .Z(n16593) );
  NAND U18270 ( .A(B[23]), .B(A[1]), .Z(n16404) );
  NAND U18271 ( .A(n16594), .B(n16595), .Z(n1717) );
  NANDN U18272 ( .A(n16596), .B(n16597), .Z(n16595) );
  OR U18273 ( .A(n16598), .B(n16599), .Z(n16597) );
  NAND U18274 ( .A(n16599), .B(n16598), .Z(n16594) );
  XOR U18275 ( .A(n1737), .B(n1736), .Z(\A1[229] ) );
  XOR U18276 ( .A(n16582), .B(n16600), .Z(n1736) );
  XNOR U18277 ( .A(n16581), .B(n16579), .Z(n16600) );
  AND U18278 ( .A(n16601), .B(n16602), .Z(n16579) );
  NANDN U18279 ( .A(n16603), .B(n16604), .Z(n16602) );
  NANDN U18280 ( .A(n16605), .B(n16606), .Z(n16604) );
  AND U18281 ( .A(B[228]), .B(A[3]), .Z(n16581) );
  XNOR U18282 ( .A(n16571), .B(n16607), .Z(n16582) );
  XNOR U18283 ( .A(n16569), .B(n16572), .Z(n16607) );
  NAND U18284 ( .A(A[2]), .B(B[229]), .Z(n16572) );
  NANDN U18285 ( .A(n16608), .B(n16609), .Z(n16569) );
  AND U18286 ( .A(A[0]), .B(B[230]), .Z(n16609) );
  XOR U18287 ( .A(n16574), .B(n16610), .Z(n16571) );
  NAND U18288 ( .A(A[0]), .B(B[231]), .Z(n16610) );
  NAND U18289 ( .A(B[230]), .B(A[1]), .Z(n16574) );
  NAND U18290 ( .A(n16611), .B(n16612), .Z(n1737) );
  NANDN U18291 ( .A(n16613), .B(n16614), .Z(n16612) );
  OR U18292 ( .A(n16615), .B(n16616), .Z(n16614) );
  NAND U18293 ( .A(n16616), .B(n16615), .Z(n16611) );
  XOR U18294 ( .A(n1741), .B(n1740), .Z(\A1[228] ) );
  XOR U18295 ( .A(n16616), .B(n16617), .Z(n1740) );
  XNOR U18296 ( .A(n16615), .B(n16613), .Z(n16617) );
  AND U18297 ( .A(n16618), .B(n16619), .Z(n16613) );
  NANDN U18298 ( .A(n16620), .B(n16621), .Z(n16619) );
  NANDN U18299 ( .A(n16622), .B(n16623), .Z(n16621) );
  AND U18300 ( .A(B[227]), .B(A[3]), .Z(n16615) );
  XNOR U18301 ( .A(n16605), .B(n16624), .Z(n16616) );
  XNOR U18302 ( .A(n16603), .B(n16606), .Z(n16624) );
  NAND U18303 ( .A(A[2]), .B(B[228]), .Z(n16606) );
  NANDN U18304 ( .A(n16625), .B(n16626), .Z(n16603) );
  AND U18305 ( .A(A[0]), .B(B[229]), .Z(n16626) );
  XOR U18306 ( .A(n16608), .B(n16627), .Z(n16605) );
  NAND U18307 ( .A(A[0]), .B(B[230]), .Z(n16627) );
  NAND U18308 ( .A(B[229]), .B(A[1]), .Z(n16608) );
  NAND U18309 ( .A(n16628), .B(n16629), .Z(n1741) );
  NANDN U18310 ( .A(n16630), .B(n16631), .Z(n16629) );
  OR U18311 ( .A(n16632), .B(n16633), .Z(n16631) );
  NAND U18312 ( .A(n16633), .B(n16632), .Z(n16628) );
  XOR U18313 ( .A(n1743), .B(n1742), .Z(\A1[227] ) );
  XOR U18314 ( .A(n16633), .B(n16634), .Z(n1742) );
  XNOR U18315 ( .A(n16632), .B(n16630), .Z(n16634) );
  AND U18316 ( .A(n16635), .B(n16636), .Z(n16630) );
  NANDN U18317 ( .A(n16637), .B(n16638), .Z(n16636) );
  NANDN U18318 ( .A(n16639), .B(n16640), .Z(n16638) );
  AND U18319 ( .A(B[226]), .B(A[3]), .Z(n16632) );
  XNOR U18320 ( .A(n16622), .B(n16641), .Z(n16633) );
  XNOR U18321 ( .A(n16620), .B(n16623), .Z(n16641) );
  NAND U18322 ( .A(A[2]), .B(B[227]), .Z(n16623) );
  NANDN U18323 ( .A(n16642), .B(n16643), .Z(n16620) );
  AND U18324 ( .A(A[0]), .B(B[228]), .Z(n16643) );
  XOR U18325 ( .A(n16625), .B(n16644), .Z(n16622) );
  NAND U18326 ( .A(A[0]), .B(B[229]), .Z(n16644) );
  NAND U18327 ( .A(B[228]), .B(A[1]), .Z(n16625) );
  NAND U18328 ( .A(n16645), .B(n16646), .Z(n1743) );
  NANDN U18329 ( .A(n16647), .B(n16648), .Z(n16646) );
  OR U18330 ( .A(n16649), .B(n16650), .Z(n16648) );
  NAND U18331 ( .A(n16650), .B(n16649), .Z(n16645) );
  XOR U18332 ( .A(n1745), .B(n1744), .Z(\A1[226] ) );
  XOR U18333 ( .A(n16650), .B(n16651), .Z(n1744) );
  XNOR U18334 ( .A(n16649), .B(n16647), .Z(n16651) );
  AND U18335 ( .A(n16652), .B(n16653), .Z(n16647) );
  NANDN U18336 ( .A(n16654), .B(n16655), .Z(n16653) );
  NANDN U18337 ( .A(n16656), .B(n16657), .Z(n16655) );
  AND U18338 ( .A(B[225]), .B(A[3]), .Z(n16649) );
  XNOR U18339 ( .A(n16639), .B(n16658), .Z(n16650) );
  XNOR U18340 ( .A(n16637), .B(n16640), .Z(n16658) );
  NAND U18341 ( .A(A[2]), .B(B[226]), .Z(n16640) );
  NANDN U18342 ( .A(n16659), .B(n16660), .Z(n16637) );
  AND U18343 ( .A(A[0]), .B(B[227]), .Z(n16660) );
  XOR U18344 ( .A(n16642), .B(n16661), .Z(n16639) );
  NAND U18345 ( .A(A[0]), .B(B[228]), .Z(n16661) );
  NAND U18346 ( .A(B[227]), .B(A[1]), .Z(n16642) );
  NAND U18347 ( .A(n16662), .B(n16663), .Z(n1745) );
  NANDN U18348 ( .A(n16664), .B(n16665), .Z(n16663) );
  OR U18349 ( .A(n16666), .B(n16667), .Z(n16665) );
  NAND U18350 ( .A(n16667), .B(n16666), .Z(n16662) );
  XOR U18351 ( .A(n1747), .B(n1746), .Z(\A1[225] ) );
  XOR U18352 ( .A(n16667), .B(n16668), .Z(n1746) );
  XNOR U18353 ( .A(n16666), .B(n16664), .Z(n16668) );
  AND U18354 ( .A(n16669), .B(n16670), .Z(n16664) );
  NANDN U18355 ( .A(n16671), .B(n16672), .Z(n16670) );
  NANDN U18356 ( .A(n16673), .B(n16674), .Z(n16672) );
  AND U18357 ( .A(B[224]), .B(A[3]), .Z(n16666) );
  XNOR U18358 ( .A(n16656), .B(n16675), .Z(n16667) );
  XNOR U18359 ( .A(n16654), .B(n16657), .Z(n16675) );
  NAND U18360 ( .A(A[2]), .B(B[225]), .Z(n16657) );
  NANDN U18361 ( .A(n16676), .B(n16677), .Z(n16654) );
  AND U18362 ( .A(A[0]), .B(B[226]), .Z(n16677) );
  XOR U18363 ( .A(n16659), .B(n16678), .Z(n16656) );
  NAND U18364 ( .A(A[0]), .B(B[227]), .Z(n16678) );
  NAND U18365 ( .A(B[226]), .B(A[1]), .Z(n16659) );
  NAND U18366 ( .A(n16679), .B(n16680), .Z(n1747) );
  NANDN U18367 ( .A(n16681), .B(n16682), .Z(n16680) );
  OR U18368 ( .A(n16683), .B(n16684), .Z(n16682) );
  NAND U18369 ( .A(n16684), .B(n16683), .Z(n16679) );
  XOR U18370 ( .A(n1749), .B(n1748), .Z(\A1[224] ) );
  XOR U18371 ( .A(n16684), .B(n16685), .Z(n1748) );
  XNOR U18372 ( .A(n16683), .B(n16681), .Z(n16685) );
  AND U18373 ( .A(n16686), .B(n16687), .Z(n16681) );
  NANDN U18374 ( .A(n16688), .B(n16689), .Z(n16687) );
  NANDN U18375 ( .A(n16690), .B(n16691), .Z(n16689) );
  AND U18376 ( .A(B[223]), .B(A[3]), .Z(n16683) );
  XNOR U18377 ( .A(n16673), .B(n16692), .Z(n16684) );
  XNOR U18378 ( .A(n16671), .B(n16674), .Z(n16692) );
  NAND U18379 ( .A(A[2]), .B(B[224]), .Z(n16674) );
  NANDN U18380 ( .A(n16693), .B(n16694), .Z(n16671) );
  AND U18381 ( .A(A[0]), .B(B[225]), .Z(n16694) );
  XOR U18382 ( .A(n16676), .B(n16695), .Z(n16673) );
  NAND U18383 ( .A(A[0]), .B(B[226]), .Z(n16695) );
  NAND U18384 ( .A(B[225]), .B(A[1]), .Z(n16676) );
  NAND U18385 ( .A(n16696), .B(n16697), .Z(n1749) );
  NANDN U18386 ( .A(n16698), .B(n16699), .Z(n16697) );
  OR U18387 ( .A(n16700), .B(n16701), .Z(n16699) );
  NAND U18388 ( .A(n16701), .B(n16700), .Z(n16696) );
  XOR U18389 ( .A(n1751), .B(n1750), .Z(\A1[223] ) );
  XOR U18390 ( .A(n16701), .B(n16702), .Z(n1750) );
  XNOR U18391 ( .A(n16700), .B(n16698), .Z(n16702) );
  AND U18392 ( .A(n16703), .B(n16704), .Z(n16698) );
  NANDN U18393 ( .A(n16705), .B(n16706), .Z(n16704) );
  NANDN U18394 ( .A(n16707), .B(n16708), .Z(n16706) );
  AND U18395 ( .A(B[222]), .B(A[3]), .Z(n16700) );
  XNOR U18396 ( .A(n16690), .B(n16709), .Z(n16701) );
  XNOR U18397 ( .A(n16688), .B(n16691), .Z(n16709) );
  NAND U18398 ( .A(A[2]), .B(B[223]), .Z(n16691) );
  NANDN U18399 ( .A(n16710), .B(n16711), .Z(n16688) );
  AND U18400 ( .A(A[0]), .B(B[224]), .Z(n16711) );
  XOR U18401 ( .A(n16693), .B(n16712), .Z(n16690) );
  NAND U18402 ( .A(A[0]), .B(B[225]), .Z(n16712) );
  NAND U18403 ( .A(B[224]), .B(A[1]), .Z(n16693) );
  NAND U18404 ( .A(n16713), .B(n16714), .Z(n1751) );
  NANDN U18405 ( .A(n16715), .B(n16716), .Z(n16714) );
  OR U18406 ( .A(n16717), .B(n16718), .Z(n16716) );
  NAND U18407 ( .A(n16718), .B(n16717), .Z(n16713) );
  XOR U18408 ( .A(n1753), .B(n1752), .Z(\A1[222] ) );
  XOR U18409 ( .A(n16718), .B(n16719), .Z(n1752) );
  XNOR U18410 ( .A(n16717), .B(n16715), .Z(n16719) );
  AND U18411 ( .A(n16720), .B(n16721), .Z(n16715) );
  NANDN U18412 ( .A(n16722), .B(n16723), .Z(n16721) );
  NANDN U18413 ( .A(n16724), .B(n16725), .Z(n16723) );
  AND U18414 ( .A(B[221]), .B(A[3]), .Z(n16717) );
  XNOR U18415 ( .A(n16707), .B(n16726), .Z(n16718) );
  XNOR U18416 ( .A(n16705), .B(n16708), .Z(n16726) );
  NAND U18417 ( .A(A[2]), .B(B[222]), .Z(n16708) );
  NANDN U18418 ( .A(n16727), .B(n16728), .Z(n16705) );
  AND U18419 ( .A(A[0]), .B(B[223]), .Z(n16728) );
  XOR U18420 ( .A(n16710), .B(n16729), .Z(n16707) );
  NAND U18421 ( .A(A[0]), .B(B[224]), .Z(n16729) );
  NAND U18422 ( .A(B[223]), .B(A[1]), .Z(n16710) );
  NAND U18423 ( .A(n16730), .B(n16731), .Z(n1753) );
  NANDN U18424 ( .A(n16732), .B(n16733), .Z(n16731) );
  OR U18425 ( .A(n16734), .B(n16735), .Z(n16733) );
  NAND U18426 ( .A(n16735), .B(n16734), .Z(n16730) );
  XOR U18427 ( .A(n1755), .B(n1754), .Z(\A1[221] ) );
  XOR U18428 ( .A(n16735), .B(n16736), .Z(n1754) );
  XNOR U18429 ( .A(n16734), .B(n16732), .Z(n16736) );
  AND U18430 ( .A(n16737), .B(n16738), .Z(n16732) );
  NANDN U18431 ( .A(n16739), .B(n16740), .Z(n16738) );
  NANDN U18432 ( .A(n16741), .B(n16742), .Z(n16740) );
  AND U18433 ( .A(B[220]), .B(A[3]), .Z(n16734) );
  XNOR U18434 ( .A(n16724), .B(n16743), .Z(n16735) );
  XNOR U18435 ( .A(n16722), .B(n16725), .Z(n16743) );
  NAND U18436 ( .A(A[2]), .B(B[221]), .Z(n16725) );
  NANDN U18437 ( .A(n16744), .B(n16745), .Z(n16722) );
  AND U18438 ( .A(A[0]), .B(B[222]), .Z(n16745) );
  XOR U18439 ( .A(n16727), .B(n16746), .Z(n16724) );
  NAND U18440 ( .A(A[0]), .B(B[223]), .Z(n16746) );
  NAND U18441 ( .A(B[222]), .B(A[1]), .Z(n16727) );
  NAND U18442 ( .A(n16747), .B(n16748), .Z(n1755) );
  NANDN U18443 ( .A(n16749), .B(n16750), .Z(n16748) );
  OR U18444 ( .A(n16751), .B(n16752), .Z(n16750) );
  NAND U18445 ( .A(n16752), .B(n16751), .Z(n16747) );
  XOR U18446 ( .A(n1757), .B(n1756), .Z(\A1[220] ) );
  XOR U18447 ( .A(n16752), .B(n16753), .Z(n1756) );
  XNOR U18448 ( .A(n16751), .B(n16749), .Z(n16753) );
  AND U18449 ( .A(n16754), .B(n16755), .Z(n16749) );
  NANDN U18450 ( .A(n16756), .B(n16757), .Z(n16755) );
  NANDN U18451 ( .A(n16758), .B(n16759), .Z(n16757) );
  AND U18452 ( .A(B[219]), .B(A[3]), .Z(n16751) );
  XNOR U18453 ( .A(n16741), .B(n16760), .Z(n16752) );
  XNOR U18454 ( .A(n16739), .B(n16742), .Z(n16760) );
  NAND U18455 ( .A(A[2]), .B(B[220]), .Z(n16742) );
  NANDN U18456 ( .A(n16761), .B(n16762), .Z(n16739) );
  AND U18457 ( .A(A[0]), .B(B[221]), .Z(n16762) );
  XOR U18458 ( .A(n16744), .B(n16763), .Z(n16741) );
  NAND U18459 ( .A(A[0]), .B(B[222]), .Z(n16763) );
  NAND U18460 ( .A(B[221]), .B(A[1]), .Z(n16744) );
  NAND U18461 ( .A(n16764), .B(n16765), .Z(n1757) );
  NANDN U18462 ( .A(n16766), .B(n16767), .Z(n16765) );
  OR U18463 ( .A(n16768), .B(n16769), .Z(n16767) );
  NAND U18464 ( .A(n16769), .B(n16768), .Z(n16764) );
  XOR U18465 ( .A(n1739), .B(n1738), .Z(\A1[21] ) );
  XOR U18466 ( .A(n16599), .B(n16770), .Z(n1738) );
  XNOR U18467 ( .A(n16598), .B(n16596), .Z(n16770) );
  AND U18468 ( .A(n16771), .B(n16772), .Z(n16596) );
  NANDN U18469 ( .A(n16773), .B(n16774), .Z(n16772) );
  NANDN U18470 ( .A(n16775), .B(n16776), .Z(n16774) );
  AND U18471 ( .A(B[20]), .B(A[3]), .Z(n16598) );
  XNOR U18472 ( .A(n16588), .B(n16777), .Z(n16599) );
  XNOR U18473 ( .A(n16586), .B(n16589), .Z(n16777) );
  NAND U18474 ( .A(A[2]), .B(B[21]), .Z(n16589) );
  NANDN U18475 ( .A(n16778), .B(n16779), .Z(n16586) );
  AND U18476 ( .A(A[0]), .B(B[22]), .Z(n16779) );
  XOR U18477 ( .A(n16591), .B(n16780), .Z(n16588) );
  NAND U18478 ( .A(A[0]), .B(B[23]), .Z(n16780) );
  NAND U18479 ( .A(B[22]), .B(A[1]), .Z(n16591) );
  NAND U18480 ( .A(n16781), .B(n16782), .Z(n1739) );
  NANDN U18481 ( .A(n16783), .B(n16784), .Z(n16782) );
  OR U18482 ( .A(n16785), .B(n16786), .Z(n16784) );
  NAND U18483 ( .A(n16786), .B(n16785), .Z(n16781) );
  XOR U18484 ( .A(n1759), .B(n1758), .Z(\A1[219] ) );
  XOR U18485 ( .A(n16769), .B(n16787), .Z(n1758) );
  XNOR U18486 ( .A(n16768), .B(n16766), .Z(n16787) );
  AND U18487 ( .A(n16788), .B(n16789), .Z(n16766) );
  NANDN U18488 ( .A(n16790), .B(n16791), .Z(n16789) );
  NANDN U18489 ( .A(n16792), .B(n16793), .Z(n16791) );
  AND U18490 ( .A(B[218]), .B(A[3]), .Z(n16768) );
  XNOR U18491 ( .A(n16758), .B(n16794), .Z(n16769) );
  XNOR U18492 ( .A(n16756), .B(n16759), .Z(n16794) );
  NAND U18493 ( .A(A[2]), .B(B[219]), .Z(n16759) );
  NANDN U18494 ( .A(n16795), .B(n16796), .Z(n16756) );
  AND U18495 ( .A(A[0]), .B(B[220]), .Z(n16796) );
  XOR U18496 ( .A(n16761), .B(n16797), .Z(n16758) );
  NAND U18497 ( .A(A[0]), .B(B[221]), .Z(n16797) );
  NAND U18498 ( .A(B[220]), .B(A[1]), .Z(n16761) );
  NAND U18499 ( .A(n16798), .B(n16799), .Z(n1759) );
  NANDN U18500 ( .A(n16800), .B(n16801), .Z(n16799) );
  OR U18501 ( .A(n16802), .B(n16803), .Z(n16801) );
  NAND U18502 ( .A(n16803), .B(n16802), .Z(n16798) );
  XOR U18503 ( .A(n1763), .B(n1762), .Z(\A1[218] ) );
  XOR U18504 ( .A(n16803), .B(n16804), .Z(n1762) );
  XNOR U18505 ( .A(n16802), .B(n16800), .Z(n16804) );
  AND U18506 ( .A(n16805), .B(n16806), .Z(n16800) );
  NANDN U18507 ( .A(n16807), .B(n16808), .Z(n16806) );
  NANDN U18508 ( .A(n16809), .B(n16810), .Z(n16808) );
  AND U18509 ( .A(B[217]), .B(A[3]), .Z(n16802) );
  XNOR U18510 ( .A(n16792), .B(n16811), .Z(n16803) );
  XNOR U18511 ( .A(n16790), .B(n16793), .Z(n16811) );
  NAND U18512 ( .A(A[2]), .B(B[218]), .Z(n16793) );
  NANDN U18513 ( .A(n16812), .B(n16813), .Z(n16790) );
  AND U18514 ( .A(A[0]), .B(B[219]), .Z(n16813) );
  XOR U18515 ( .A(n16795), .B(n16814), .Z(n16792) );
  NAND U18516 ( .A(A[0]), .B(B[220]), .Z(n16814) );
  NAND U18517 ( .A(B[219]), .B(A[1]), .Z(n16795) );
  NAND U18518 ( .A(n16815), .B(n16816), .Z(n1763) );
  NANDN U18519 ( .A(n16817), .B(n16818), .Z(n16816) );
  OR U18520 ( .A(n16819), .B(n16820), .Z(n16818) );
  NAND U18521 ( .A(n16820), .B(n16819), .Z(n16815) );
  XOR U18522 ( .A(n1765), .B(n1764), .Z(\A1[217] ) );
  XOR U18523 ( .A(n16820), .B(n16821), .Z(n1764) );
  XNOR U18524 ( .A(n16819), .B(n16817), .Z(n16821) );
  AND U18525 ( .A(n16822), .B(n16823), .Z(n16817) );
  NANDN U18526 ( .A(n16824), .B(n16825), .Z(n16823) );
  NANDN U18527 ( .A(n16826), .B(n16827), .Z(n16825) );
  AND U18528 ( .A(B[216]), .B(A[3]), .Z(n16819) );
  XNOR U18529 ( .A(n16809), .B(n16828), .Z(n16820) );
  XNOR U18530 ( .A(n16807), .B(n16810), .Z(n16828) );
  NAND U18531 ( .A(A[2]), .B(B[217]), .Z(n16810) );
  NANDN U18532 ( .A(n16829), .B(n16830), .Z(n16807) );
  AND U18533 ( .A(A[0]), .B(B[218]), .Z(n16830) );
  XOR U18534 ( .A(n16812), .B(n16831), .Z(n16809) );
  NAND U18535 ( .A(A[0]), .B(B[219]), .Z(n16831) );
  NAND U18536 ( .A(B[218]), .B(A[1]), .Z(n16812) );
  NAND U18537 ( .A(n16832), .B(n16833), .Z(n1765) );
  NANDN U18538 ( .A(n16834), .B(n16835), .Z(n16833) );
  OR U18539 ( .A(n16836), .B(n16837), .Z(n16835) );
  NAND U18540 ( .A(n16837), .B(n16836), .Z(n16832) );
  XOR U18541 ( .A(n1767), .B(n1766), .Z(\A1[216] ) );
  XOR U18542 ( .A(n16837), .B(n16838), .Z(n1766) );
  XNOR U18543 ( .A(n16836), .B(n16834), .Z(n16838) );
  AND U18544 ( .A(n16839), .B(n16840), .Z(n16834) );
  NANDN U18545 ( .A(n16841), .B(n16842), .Z(n16840) );
  NANDN U18546 ( .A(n16843), .B(n16844), .Z(n16842) );
  AND U18547 ( .A(B[215]), .B(A[3]), .Z(n16836) );
  XNOR U18548 ( .A(n16826), .B(n16845), .Z(n16837) );
  XNOR U18549 ( .A(n16824), .B(n16827), .Z(n16845) );
  NAND U18550 ( .A(A[2]), .B(B[216]), .Z(n16827) );
  NANDN U18551 ( .A(n16846), .B(n16847), .Z(n16824) );
  AND U18552 ( .A(A[0]), .B(B[217]), .Z(n16847) );
  XOR U18553 ( .A(n16829), .B(n16848), .Z(n16826) );
  NAND U18554 ( .A(A[0]), .B(B[218]), .Z(n16848) );
  NAND U18555 ( .A(B[217]), .B(A[1]), .Z(n16829) );
  NAND U18556 ( .A(n16849), .B(n16850), .Z(n1767) );
  NANDN U18557 ( .A(n16851), .B(n16852), .Z(n16850) );
  OR U18558 ( .A(n16853), .B(n16854), .Z(n16852) );
  NAND U18559 ( .A(n16854), .B(n16853), .Z(n16849) );
  XOR U18560 ( .A(n1769), .B(n1768), .Z(\A1[215] ) );
  XOR U18561 ( .A(n16854), .B(n16855), .Z(n1768) );
  XNOR U18562 ( .A(n16853), .B(n16851), .Z(n16855) );
  AND U18563 ( .A(n16856), .B(n16857), .Z(n16851) );
  NANDN U18564 ( .A(n16858), .B(n16859), .Z(n16857) );
  NANDN U18565 ( .A(n16860), .B(n16861), .Z(n16859) );
  AND U18566 ( .A(B[214]), .B(A[3]), .Z(n16853) );
  XNOR U18567 ( .A(n16843), .B(n16862), .Z(n16854) );
  XNOR U18568 ( .A(n16841), .B(n16844), .Z(n16862) );
  NAND U18569 ( .A(A[2]), .B(B[215]), .Z(n16844) );
  NANDN U18570 ( .A(n16863), .B(n16864), .Z(n16841) );
  AND U18571 ( .A(A[0]), .B(B[216]), .Z(n16864) );
  XOR U18572 ( .A(n16846), .B(n16865), .Z(n16843) );
  NAND U18573 ( .A(A[0]), .B(B[217]), .Z(n16865) );
  NAND U18574 ( .A(B[216]), .B(A[1]), .Z(n16846) );
  NAND U18575 ( .A(n16866), .B(n16867), .Z(n1769) );
  NANDN U18576 ( .A(n16868), .B(n16869), .Z(n16867) );
  OR U18577 ( .A(n16870), .B(n16871), .Z(n16869) );
  NAND U18578 ( .A(n16871), .B(n16870), .Z(n16866) );
  XOR U18579 ( .A(n1771), .B(n1770), .Z(\A1[214] ) );
  XOR U18580 ( .A(n16871), .B(n16872), .Z(n1770) );
  XNOR U18581 ( .A(n16870), .B(n16868), .Z(n16872) );
  AND U18582 ( .A(n16873), .B(n16874), .Z(n16868) );
  NANDN U18583 ( .A(n16875), .B(n16876), .Z(n16874) );
  NANDN U18584 ( .A(n16877), .B(n16878), .Z(n16876) );
  AND U18585 ( .A(B[213]), .B(A[3]), .Z(n16870) );
  XNOR U18586 ( .A(n16860), .B(n16879), .Z(n16871) );
  XNOR U18587 ( .A(n16858), .B(n16861), .Z(n16879) );
  NAND U18588 ( .A(A[2]), .B(B[214]), .Z(n16861) );
  NANDN U18589 ( .A(n16880), .B(n16881), .Z(n16858) );
  AND U18590 ( .A(A[0]), .B(B[215]), .Z(n16881) );
  XOR U18591 ( .A(n16863), .B(n16882), .Z(n16860) );
  NAND U18592 ( .A(A[0]), .B(B[216]), .Z(n16882) );
  NAND U18593 ( .A(B[215]), .B(A[1]), .Z(n16863) );
  NAND U18594 ( .A(n16883), .B(n16884), .Z(n1771) );
  NANDN U18595 ( .A(n16885), .B(n16886), .Z(n16884) );
  OR U18596 ( .A(n16887), .B(n16888), .Z(n16886) );
  NAND U18597 ( .A(n16888), .B(n16887), .Z(n16883) );
  XOR U18598 ( .A(n1773), .B(n1772), .Z(\A1[213] ) );
  XOR U18599 ( .A(n16888), .B(n16889), .Z(n1772) );
  XNOR U18600 ( .A(n16887), .B(n16885), .Z(n16889) );
  AND U18601 ( .A(n16890), .B(n16891), .Z(n16885) );
  NANDN U18602 ( .A(n16892), .B(n16893), .Z(n16891) );
  NANDN U18603 ( .A(n16894), .B(n16895), .Z(n16893) );
  AND U18604 ( .A(B[212]), .B(A[3]), .Z(n16887) );
  XNOR U18605 ( .A(n16877), .B(n16896), .Z(n16888) );
  XNOR U18606 ( .A(n16875), .B(n16878), .Z(n16896) );
  NAND U18607 ( .A(A[2]), .B(B[213]), .Z(n16878) );
  NANDN U18608 ( .A(n16897), .B(n16898), .Z(n16875) );
  AND U18609 ( .A(A[0]), .B(B[214]), .Z(n16898) );
  XOR U18610 ( .A(n16880), .B(n16899), .Z(n16877) );
  NAND U18611 ( .A(A[0]), .B(B[215]), .Z(n16899) );
  NAND U18612 ( .A(B[214]), .B(A[1]), .Z(n16880) );
  NAND U18613 ( .A(n16900), .B(n16901), .Z(n1773) );
  NANDN U18614 ( .A(n16902), .B(n16903), .Z(n16901) );
  OR U18615 ( .A(n16904), .B(n16905), .Z(n16903) );
  NAND U18616 ( .A(n16905), .B(n16904), .Z(n16900) );
  XOR U18617 ( .A(n1775), .B(n1774), .Z(\A1[212] ) );
  XOR U18618 ( .A(n16905), .B(n16906), .Z(n1774) );
  XNOR U18619 ( .A(n16904), .B(n16902), .Z(n16906) );
  AND U18620 ( .A(n16907), .B(n16908), .Z(n16902) );
  NANDN U18621 ( .A(n16909), .B(n16910), .Z(n16908) );
  NANDN U18622 ( .A(n16911), .B(n16912), .Z(n16910) );
  AND U18623 ( .A(B[211]), .B(A[3]), .Z(n16904) );
  XNOR U18624 ( .A(n16894), .B(n16913), .Z(n16905) );
  XNOR U18625 ( .A(n16892), .B(n16895), .Z(n16913) );
  NAND U18626 ( .A(A[2]), .B(B[212]), .Z(n16895) );
  NANDN U18627 ( .A(n16914), .B(n16915), .Z(n16892) );
  AND U18628 ( .A(A[0]), .B(B[213]), .Z(n16915) );
  XOR U18629 ( .A(n16897), .B(n16916), .Z(n16894) );
  NAND U18630 ( .A(A[0]), .B(B[214]), .Z(n16916) );
  NAND U18631 ( .A(B[213]), .B(A[1]), .Z(n16897) );
  NAND U18632 ( .A(n16917), .B(n16918), .Z(n1775) );
  NANDN U18633 ( .A(n16919), .B(n16920), .Z(n16918) );
  OR U18634 ( .A(n16921), .B(n16922), .Z(n16920) );
  NAND U18635 ( .A(n16922), .B(n16921), .Z(n16917) );
  XOR U18636 ( .A(n1777), .B(n1776), .Z(\A1[211] ) );
  XOR U18637 ( .A(n16922), .B(n16923), .Z(n1776) );
  XNOR U18638 ( .A(n16921), .B(n16919), .Z(n16923) );
  AND U18639 ( .A(n16924), .B(n16925), .Z(n16919) );
  NANDN U18640 ( .A(n16926), .B(n16927), .Z(n16925) );
  NANDN U18641 ( .A(n16928), .B(n16929), .Z(n16927) );
  AND U18642 ( .A(B[210]), .B(A[3]), .Z(n16921) );
  XNOR U18643 ( .A(n16911), .B(n16930), .Z(n16922) );
  XNOR U18644 ( .A(n16909), .B(n16912), .Z(n16930) );
  NAND U18645 ( .A(A[2]), .B(B[211]), .Z(n16912) );
  NANDN U18646 ( .A(n16931), .B(n16932), .Z(n16909) );
  AND U18647 ( .A(A[0]), .B(B[212]), .Z(n16932) );
  XOR U18648 ( .A(n16914), .B(n16933), .Z(n16911) );
  NAND U18649 ( .A(A[0]), .B(B[213]), .Z(n16933) );
  NAND U18650 ( .A(B[212]), .B(A[1]), .Z(n16914) );
  NAND U18651 ( .A(n16934), .B(n16935), .Z(n1777) );
  NANDN U18652 ( .A(n16936), .B(n16937), .Z(n16935) );
  OR U18653 ( .A(n16938), .B(n16939), .Z(n16937) );
  NAND U18654 ( .A(n16939), .B(n16938), .Z(n16934) );
  XOR U18655 ( .A(n1779), .B(n1778), .Z(\A1[210] ) );
  XOR U18656 ( .A(n16939), .B(n16940), .Z(n1778) );
  XNOR U18657 ( .A(n16938), .B(n16936), .Z(n16940) );
  AND U18658 ( .A(n16941), .B(n16942), .Z(n16936) );
  NANDN U18659 ( .A(n16943), .B(n16944), .Z(n16942) );
  NANDN U18660 ( .A(n16945), .B(n16946), .Z(n16944) );
  AND U18661 ( .A(B[209]), .B(A[3]), .Z(n16938) );
  XNOR U18662 ( .A(n16928), .B(n16947), .Z(n16939) );
  XNOR U18663 ( .A(n16926), .B(n16929), .Z(n16947) );
  NAND U18664 ( .A(A[2]), .B(B[210]), .Z(n16929) );
  NANDN U18665 ( .A(n16948), .B(n16949), .Z(n16926) );
  AND U18666 ( .A(A[0]), .B(B[211]), .Z(n16949) );
  XOR U18667 ( .A(n16931), .B(n16950), .Z(n16928) );
  NAND U18668 ( .A(A[0]), .B(B[212]), .Z(n16950) );
  NAND U18669 ( .A(B[211]), .B(A[1]), .Z(n16931) );
  NAND U18670 ( .A(n16951), .B(n16952), .Z(n1779) );
  NANDN U18671 ( .A(n16953), .B(n16954), .Z(n16952) );
  OR U18672 ( .A(n16955), .B(n16956), .Z(n16954) );
  NAND U18673 ( .A(n16956), .B(n16955), .Z(n16951) );
  XOR U18674 ( .A(n1761), .B(n1760), .Z(\A1[20] ) );
  XOR U18675 ( .A(n16786), .B(n16957), .Z(n1760) );
  XNOR U18676 ( .A(n16785), .B(n16783), .Z(n16957) );
  AND U18677 ( .A(n16958), .B(n16959), .Z(n16783) );
  NANDN U18678 ( .A(n16960), .B(n16961), .Z(n16959) );
  NANDN U18679 ( .A(n16962), .B(n16963), .Z(n16961) );
  AND U18680 ( .A(B[19]), .B(A[3]), .Z(n16785) );
  XNOR U18681 ( .A(n16775), .B(n16964), .Z(n16786) );
  XNOR U18682 ( .A(n16773), .B(n16776), .Z(n16964) );
  NAND U18683 ( .A(A[2]), .B(B[20]), .Z(n16776) );
  NANDN U18684 ( .A(n16965), .B(n16966), .Z(n16773) );
  AND U18685 ( .A(A[0]), .B(B[21]), .Z(n16966) );
  XOR U18686 ( .A(n16778), .B(n16967), .Z(n16775) );
  NAND U18687 ( .A(A[0]), .B(B[22]), .Z(n16967) );
  NAND U18688 ( .A(B[21]), .B(A[1]), .Z(n16778) );
  NAND U18689 ( .A(n16968), .B(n16969), .Z(n1761) );
  NANDN U18690 ( .A(n16970), .B(n16971), .Z(n16969) );
  OR U18691 ( .A(n16972), .B(n16973), .Z(n16971) );
  NAND U18692 ( .A(n16973), .B(n16972), .Z(n16968) );
  XOR U18693 ( .A(n1781), .B(n1780), .Z(\A1[209] ) );
  XOR U18694 ( .A(n16956), .B(n16974), .Z(n1780) );
  XNOR U18695 ( .A(n16955), .B(n16953), .Z(n16974) );
  AND U18696 ( .A(n16975), .B(n16976), .Z(n16953) );
  NANDN U18697 ( .A(n16977), .B(n16978), .Z(n16976) );
  NANDN U18698 ( .A(n16979), .B(n16980), .Z(n16978) );
  AND U18699 ( .A(B[208]), .B(A[3]), .Z(n16955) );
  XNOR U18700 ( .A(n16945), .B(n16981), .Z(n16956) );
  XNOR U18701 ( .A(n16943), .B(n16946), .Z(n16981) );
  NAND U18702 ( .A(A[2]), .B(B[209]), .Z(n16946) );
  NANDN U18703 ( .A(n16982), .B(n16983), .Z(n16943) );
  AND U18704 ( .A(A[0]), .B(B[210]), .Z(n16983) );
  XOR U18705 ( .A(n16948), .B(n16984), .Z(n16945) );
  NAND U18706 ( .A(A[0]), .B(B[211]), .Z(n16984) );
  NAND U18707 ( .A(B[210]), .B(A[1]), .Z(n16948) );
  NAND U18708 ( .A(n16985), .B(n16986), .Z(n1781) );
  NANDN U18709 ( .A(n16987), .B(n16988), .Z(n16986) );
  OR U18710 ( .A(n16989), .B(n16990), .Z(n16988) );
  NAND U18711 ( .A(n16990), .B(n16989), .Z(n16985) );
  XOR U18712 ( .A(n1785), .B(n1784), .Z(\A1[208] ) );
  XOR U18713 ( .A(n16990), .B(n16991), .Z(n1784) );
  XNOR U18714 ( .A(n16989), .B(n16987), .Z(n16991) );
  AND U18715 ( .A(n16992), .B(n16993), .Z(n16987) );
  NANDN U18716 ( .A(n16994), .B(n16995), .Z(n16993) );
  NANDN U18717 ( .A(n16996), .B(n16997), .Z(n16995) );
  AND U18718 ( .A(B[207]), .B(A[3]), .Z(n16989) );
  XNOR U18719 ( .A(n16979), .B(n16998), .Z(n16990) );
  XNOR U18720 ( .A(n16977), .B(n16980), .Z(n16998) );
  NAND U18721 ( .A(A[2]), .B(B[208]), .Z(n16980) );
  NANDN U18722 ( .A(n16999), .B(n17000), .Z(n16977) );
  AND U18723 ( .A(A[0]), .B(B[209]), .Z(n17000) );
  XOR U18724 ( .A(n16982), .B(n17001), .Z(n16979) );
  NAND U18725 ( .A(A[0]), .B(B[210]), .Z(n17001) );
  NAND U18726 ( .A(B[209]), .B(A[1]), .Z(n16982) );
  NAND U18727 ( .A(n17002), .B(n17003), .Z(n1785) );
  NANDN U18728 ( .A(n17004), .B(n17005), .Z(n17003) );
  OR U18729 ( .A(n17006), .B(n17007), .Z(n17005) );
  NAND U18730 ( .A(n17007), .B(n17006), .Z(n17002) );
  XOR U18731 ( .A(n1787), .B(n1786), .Z(\A1[207] ) );
  XOR U18732 ( .A(n17007), .B(n17008), .Z(n1786) );
  XNOR U18733 ( .A(n17006), .B(n17004), .Z(n17008) );
  AND U18734 ( .A(n17009), .B(n17010), .Z(n17004) );
  NANDN U18735 ( .A(n17011), .B(n17012), .Z(n17010) );
  NANDN U18736 ( .A(n17013), .B(n17014), .Z(n17012) );
  AND U18737 ( .A(B[206]), .B(A[3]), .Z(n17006) );
  XNOR U18738 ( .A(n16996), .B(n17015), .Z(n17007) );
  XNOR U18739 ( .A(n16994), .B(n16997), .Z(n17015) );
  NAND U18740 ( .A(A[2]), .B(B[207]), .Z(n16997) );
  NANDN U18741 ( .A(n17016), .B(n17017), .Z(n16994) );
  AND U18742 ( .A(A[0]), .B(B[208]), .Z(n17017) );
  XOR U18743 ( .A(n16999), .B(n17018), .Z(n16996) );
  NAND U18744 ( .A(A[0]), .B(B[209]), .Z(n17018) );
  NAND U18745 ( .A(B[208]), .B(A[1]), .Z(n16999) );
  NAND U18746 ( .A(n17019), .B(n17020), .Z(n1787) );
  NANDN U18747 ( .A(n17021), .B(n17022), .Z(n17020) );
  OR U18748 ( .A(n17023), .B(n17024), .Z(n17022) );
  NAND U18749 ( .A(n17024), .B(n17023), .Z(n17019) );
  XOR U18750 ( .A(n1789), .B(n1788), .Z(\A1[206] ) );
  XOR U18751 ( .A(n17024), .B(n17025), .Z(n1788) );
  XNOR U18752 ( .A(n17023), .B(n17021), .Z(n17025) );
  AND U18753 ( .A(n17026), .B(n17027), .Z(n17021) );
  NANDN U18754 ( .A(n17028), .B(n17029), .Z(n17027) );
  NANDN U18755 ( .A(n17030), .B(n17031), .Z(n17029) );
  AND U18756 ( .A(B[205]), .B(A[3]), .Z(n17023) );
  XNOR U18757 ( .A(n17013), .B(n17032), .Z(n17024) );
  XNOR U18758 ( .A(n17011), .B(n17014), .Z(n17032) );
  NAND U18759 ( .A(A[2]), .B(B[206]), .Z(n17014) );
  NANDN U18760 ( .A(n17033), .B(n17034), .Z(n17011) );
  AND U18761 ( .A(A[0]), .B(B[207]), .Z(n17034) );
  XOR U18762 ( .A(n17016), .B(n17035), .Z(n17013) );
  NAND U18763 ( .A(A[0]), .B(B[208]), .Z(n17035) );
  NAND U18764 ( .A(B[207]), .B(A[1]), .Z(n17016) );
  NAND U18765 ( .A(n17036), .B(n17037), .Z(n1789) );
  NANDN U18766 ( .A(n17038), .B(n17039), .Z(n17037) );
  OR U18767 ( .A(n17040), .B(n17041), .Z(n17039) );
  NAND U18768 ( .A(n17041), .B(n17040), .Z(n17036) );
  XOR U18769 ( .A(n1791), .B(n1790), .Z(\A1[205] ) );
  XOR U18770 ( .A(n17041), .B(n17042), .Z(n1790) );
  XNOR U18771 ( .A(n17040), .B(n17038), .Z(n17042) );
  AND U18772 ( .A(n17043), .B(n17044), .Z(n17038) );
  NANDN U18773 ( .A(n17045), .B(n17046), .Z(n17044) );
  NANDN U18774 ( .A(n17047), .B(n17048), .Z(n17046) );
  AND U18775 ( .A(B[204]), .B(A[3]), .Z(n17040) );
  XNOR U18776 ( .A(n17030), .B(n17049), .Z(n17041) );
  XNOR U18777 ( .A(n17028), .B(n17031), .Z(n17049) );
  NAND U18778 ( .A(A[2]), .B(B[205]), .Z(n17031) );
  NANDN U18779 ( .A(n17050), .B(n17051), .Z(n17028) );
  AND U18780 ( .A(A[0]), .B(B[206]), .Z(n17051) );
  XOR U18781 ( .A(n17033), .B(n17052), .Z(n17030) );
  NAND U18782 ( .A(A[0]), .B(B[207]), .Z(n17052) );
  NAND U18783 ( .A(B[206]), .B(A[1]), .Z(n17033) );
  NAND U18784 ( .A(n17053), .B(n17054), .Z(n1791) );
  NANDN U18785 ( .A(n17055), .B(n17056), .Z(n17054) );
  OR U18786 ( .A(n17057), .B(n17058), .Z(n17056) );
  NAND U18787 ( .A(n17058), .B(n17057), .Z(n17053) );
  XOR U18788 ( .A(n1793), .B(n1792), .Z(\A1[204] ) );
  XOR U18789 ( .A(n17058), .B(n17059), .Z(n1792) );
  XNOR U18790 ( .A(n17057), .B(n17055), .Z(n17059) );
  AND U18791 ( .A(n17060), .B(n17061), .Z(n17055) );
  NANDN U18792 ( .A(n17062), .B(n17063), .Z(n17061) );
  NANDN U18793 ( .A(n17064), .B(n17065), .Z(n17063) );
  AND U18794 ( .A(B[203]), .B(A[3]), .Z(n17057) );
  XNOR U18795 ( .A(n17047), .B(n17066), .Z(n17058) );
  XNOR U18796 ( .A(n17045), .B(n17048), .Z(n17066) );
  NAND U18797 ( .A(A[2]), .B(B[204]), .Z(n17048) );
  NANDN U18798 ( .A(n17067), .B(n17068), .Z(n17045) );
  AND U18799 ( .A(A[0]), .B(B[205]), .Z(n17068) );
  XOR U18800 ( .A(n17050), .B(n17069), .Z(n17047) );
  NAND U18801 ( .A(A[0]), .B(B[206]), .Z(n17069) );
  NAND U18802 ( .A(B[205]), .B(A[1]), .Z(n17050) );
  NAND U18803 ( .A(n17070), .B(n17071), .Z(n1793) );
  NANDN U18804 ( .A(n17072), .B(n17073), .Z(n17071) );
  OR U18805 ( .A(n17074), .B(n17075), .Z(n17073) );
  NAND U18806 ( .A(n17075), .B(n17074), .Z(n17070) );
  XOR U18807 ( .A(n1795), .B(n1794), .Z(\A1[203] ) );
  XOR U18808 ( .A(n17075), .B(n17076), .Z(n1794) );
  XNOR U18809 ( .A(n17074), .B(n17072), .Z(n17076) );
  AND U18810 ( .A(n17077), .B(n17078), .Z(n17072) );
  NANDN U18811 ( .A(n17079), .B(n17080), .Z(n17078) );
  NANDN U18812 ( .A(n17081), .B(n17082), .Z(n17080) );
  AND U18813 ( .A(B[202]), .B(A[3]), .Z(n17074) );
  XNOR U18814 ( .A(n17064), .B(n17083), .Z(n17075) );
  XNOR U18815 ( .A(n17062), .B(n17065), .Z(n17083) );
  NAND U18816 ( .A(A[2]), .B(B[203]), .Z(n17065) );
  NANDN U18817 ( .A(n17084), .B(n17085), .Z(n17062) );
  AND U18818 ( .A(A[0]), .B(B[204]), .Z(n17085) );
  XOR U18819 ( .A(n17067), .B(n17086), .Z(n17064) );
  NAND U18820 ( .A(A[0]), .B(B[205]), .Z(n17086) );
  NAND U18821 ( .A(B[204]), .B(A[1]), .Z(n17067) );
  NAND U18822 ( .A(n17087), .B(n17088), .Z(n1795) );
  NANDN U18823 ( .A(n17089), .B(n17090), .Z(n17088) );
  OR U18824 ( .A(n17091), .B(n17092), .Z(n17090) );
  NAND U18825 ( .A(n17092), .B(n17091), .Z(n17087) );
  XOR U18826 ( .A(n1797), .B(n1796), .Z(\A1[202] ) );
  XOR U18827 ( .A(n17092), .B(n17093), .Z(n1796) );
  XNOR U18828 ( .A(n17091), .B(n17089), .Z(n17093) );
  AND U18829 ( .A(n17094), .B(n17095), .Z(n17089) );
  NANDN U18830 ( .A(n17096), .B(n17097), .Z(n17095) );
  NANDN U18831 ( .A(n17098), .B(n17099), .Z(n17097) );
  AND U18832 ( .A(B[201]), .B(A[3]), .Z(n17091) );
  XNOR U18833 ( .A(n17081), .B(n17100), .Z(n17092) );
  XNOR U18834 ( .A(n17079), .B(n17082), .Z(n17100) );
  NAND U18835 ( .A(A[2]), .B(B[202]), .Z(n17082) );
  NANDN U18836 ( .A(n17101), .B(n17102), .Z(n17079) );
  AND U18837 ( .A(A[0]), .B(B[203]), .Z(n17102) );
  XOR U18838 ( .A(n17084), .B(n17103), .Z(n17081) );
  NAND U18839 ( .A(A[0]), .B(B[204]), .Z(n17103) );
  NAND U18840 ( .A(B[203]), .B(A[1]), .Z(n17084) );
  NAND U18841 ( .A(n17104), .B(n17105), .Z(n1797) );
  NANDN U18842 ( .A(n17106), .B(n17107), .Z(n17105) );
  OR U18843 ( .A(n17108), .B(n17109), .Z(n17107) );
  NAND U18844 ( .A(n17109), .B(n17108), .Z(n17104) );
  XOR U18845 ( .A(n1799), .B(n1798), .Z(\A1[201] ) );
  XOR U18846 ( .A(n17109), .B(n17110), .Z(n1798) );
  XNOR U18847 ( .A(n17108), .B(n17106), .Z(n17110) );
  AND U18848 ( .A(n17111), .B(n17112), .Z(n17106) );
  NANDN U18849 ( .A(n17113), .B(n17114), .Z(n17112) );
  NANDN U18850 ( .A(n17115), .B(n17116), .Z(n17114) );
  AND U18851 ( .A(B[200]), .B(A[3]), .Z(n17108) );
  XNOR U18852 ( .A(n17098), .B(n17117), .Z(n17109) );
  XNOR U18853 ( .A(n17096), .B(n17099), .Z(n17117) );
  NAND U18854 ( .A(A[2]), .B(B[201]), .Z(n17099) );
  NANDN U18855 ( .A(n17118), .B(n17119), .Z(n17096) );
  AND U18856 ( .A(A[0]), .B(B[202]), .Z(n17119) );
  XOR U18857 ( .A(n17101), .B(n17120), .Z(n17098) );
  NAND U18858 ( .A(A[0]), .B(B[203]), .Z(n17120) );
  NAND U18859 ( .A(B[202]), .B(A[1]), .Z(n17101) );
  NAND U18860 ( .A(n17121), .B(n17122), .Z(n1799) );
  NANDN U18861 ( .A(n17123), .B(n17124), .Z(n17122) );
  OR U18862 ( .A(n17125), .B(n17126), .Z(n17124) );
  NAND U18863 ( .A(n17126), .B(n17125), .Z(n17121) );
  XOR U18864 ( .A(n1801), .B(n1800), .Z(\A1[200] ) );
  XOR U18865 ( .A(n17126), .B(n17127), .Z(n1800) );
  XNOR U18866 ( .A(n17125), .B(n17123), .Z(n17127) );
  AND U18867 ( .A(n17128), .B(n17129), .Z(n17123) );
  NANDN U18868 ( .A(n17130), .B(n17131), .Z(n17129) );
  NANDN U18869 ( .A(n17132), .B(n17133), .Z(n17131) );
  AND U18870 ( .A(B[199]), .B(A[3]), .Z(n17125) );
  XNOR U18871 ( .A(n17115), .B(n17134), .Z(n17126) );
  XNOR U18872 ( .A(n17113), .B(n17116), .Z(n17134) );
  NAND U18873 ( .A(A[2]), .B(B[200]), .Z(n17116) );
  NANDN U18874 ( .A(n17135), .B(n17136), .Z(n17113) );
  AND U18875 ( .A(A[0]), .B(B[201]), .Z(n17136) );
  XOR U18876 ( .A(n17118), .B(n17137), .Z(n17115) );
  NAND U18877 ( .A(A[0]), .B(B[202]), .Z(n17137) );
  NAND U18878 ( .A(B[201]), .B(A[1]), .Z(n17118) );
  NAND U18879 ( .A(n17138), .B(n17139), .Z(n1801) );
  NANDN U18880 ( .A(n17140), .B(n17141), .Z(n17139) );
  OR U18881 ( .A(n17142), .B(n17143), .Z(n17141) );
  NAND U18882 ( .A(n17143), .B(n17142), .Z(n17138) );
  XOR U18883 ( .A(n15273), .B(n17144), .Z(\A1[1] ) );
  XNOR U18884 ( .A(n15272), .B(n15270), .Z(n17144) );
  AND U18885 ( .A(n17145), .B(n17146), .Z(n15270) );
  NANDN U18886 ( .A(n17147), .B(n17148), .Z(n17146) );
  NANDN U18887 ( .A(n17149), .B(n25), .Z(n17148) );
  NANDN U18888 ( .A(n25), .B(n17149), .Z(n17145) );
  AND U18889 ( .A(B[0]), .B(A[3]), .Z(n15272) );
  XNOR U18890 ( .A(n15262), .B(n17151), .Z(n15273) );
  XNOR U18891 ( .A(n15260), .B(n15263), .Z(n17151) );
  NAND U18892 ( .A(B[1]), .B(A[2]), .Z(n15263) );
  NANDN U18893 ( .A(n17152), .B(n17153), .Z(n15260) );
  AND U18894 ( .A(A[0]), .B(B[2]), .Z(n17153) );
  XOR U18895 ( .A(n15265), .B(n17154), .Z(n15262) );
  NAND U18896 ( .A(A[0]), .B(B[3]), .Z(n17154) );
  NAND U18897 ( .A(B[2]), .B(A[1]), .Z(n15265) );
  XOR U18898 ( .A(n1783), .B(n1782), .Z(\A1[19] ) );
  XOR U18899 ( .A(n16973), .B(n17155), .Z(n1782) );
  XNOR U18900 ( .A(n16972), .B(n16970), .Z(n17155) );
  AND U18901 ( .A(n17156), .B(n17157), .Z(n16970) );
  NANDN U18902 ( .A(n17158), .B(n17159), .Z(n17157) );
  NANDN U18903 ( .A(n17160), .B(n17161), .Z(n17159) );
  AND U18904 ( .A(B[18]), .B(A[3]), .Z(n16972) );
  XNOR U18905 ( .A(n16962), .B(n17162), .Z(n16973) );
  XNOR U18906 ( .A(n16960), .B(n16963), .Z(n17162) );
  NAND U18907 ( .A(A[2]), .B(B[19]), .Z(n16963) );
  NANDN U18908 ( .A(n17163), .B(n17164), .Z(n16960) );
  AND U18909 ( .A(A[0]), .B(B[20]), .Z(n17164) );
  XOR U18910 ( .A(n16965), .B(n17165), .Z(n16962) );
  NAND U18911 ( .A(A[0]), .B(B[21]), .Z(n17165) );
  NAND U18912 ( .A(B[20]), .B(A[1]), .Z(n16965) );
  NAND U18913 ( .A(n17166), .B(n17167), .Z(n1783) );
  NANDN U18914 ( .A(n17168), .B(n17169), .Z(n17167) );
  OR U18915 ( .A(n17170), .B(n17171), .Z(n17169) );
  NAND U18916 ( .A(n17171), .B(n17170), .Z(n17166) );
  XOR U18917 ( .A(n1803), .B(n1802), .Z(\A1[199] ) );
  XOR U18918 ( .A(n17143), .B(n17172), .Z(n1802) );
  XNOR U18919 ( .A(n17142), .B(n17140), .Z(n17172) );
  AND U18920 ( .A(n17173), .B(n17174), .Z(n17140) );
  NANDN U18921 ( .A(n17175), .B(n17176), .Z(n17174) );
  NANDN U18922 ( .A(n17177), .B(n17178), .Z(n17176) );
  AND U18923 ( .A(B[198]), .B(A[3]), .Z(n17142) );
  XNOR U18924 ( .A(n17132), .B(n17179), .Z(n17143) );
  XNOR U18925 ( .A(n17130), .B(n17133), .Z(n17179) );
  NAND U18926 ( .A(A[2]), .B(B[199]), .Z(n17133) );
  NANDN U18927 ( .A(n17180), .B(n17181), .Z(n17130) );
  AND U18928 ( .A(A[0]), .B(B[200]), .Z(n17181) );
  XOR U18929 ( .A(n17135), .B(n17182), .Z(n17132) );
  NAND U18930 ( .A(A[0]), .B(B[201]), .Z(n17182) );
  NAND U18931 ( .A(B[200]), .B(A[1]), .Z(n17135) );
  NAND U18932 ( .A(n17183), .B(n17184), .Z(n1803) );
  NANDN U18933 ( .A(n17185), .B(n17186), .Z(n17184) );
  OR U18934 ( .A(n17187), .B(n17188), .Z(n17186) );
  NAND U18935 ( .A(n17188), .B(n17187), .Z(n17183) );
  XOR U18936 ( .A(n1807), .B(n1806), .Z(\A1[198] ) );
  XOR U18937 ( .A(n17188), .B(n17189), .Z(n1806) );
  XNOR U18938 ( .A(n17187), .B(n17185), .Z(n17189) );
  AND U18939 ( .A(n17190), .B(n17191), .Z(n17185) );
  NANDN U18940 ( .A(n17192), .B(n17193), .Z(n17191) );
  NANDN U18941 ( .A(n17194), .B(n17195), .Z(n17193) );
  AND U18942 ( .A(B[197]), .B(A[3]), .Z(n17187) );
  XNOR U18943 ( .A(n17177), .B(n17196), .Z(n17188) );
  XNOR U18944 ( .A(n17175), .B(n17178), .Z(n17196) );
  NAND U18945 ( .A(A[2]), .B(B[198]), .Z(n17178) );
  NANDN U18946 ( .A(n17197), .B(n17198), .Z(n17175) );
  AND U18947 ( .A(A[0]), .B(B[199]), .Z(n17198) );
  XOR U18948 ( .A(n17180), .B(n17199), .Z(n17177) );
  NAND U18949 ( .A(A[0]), .B(B[200]), .Z(n17199) );
  NAND U18950 ( .A(B[199]), .B(A[1]), .Z(n17180) );
  NAND U18951 ( .A(n17200), .B(n17201), .Z(n1807) );
  NANDN U18952 ( .A(n17202), .B(n17203), .Z(n17201) );
  OR U18953 ( .A(n17204), .B(n17205), .Z(n17203) );
  NAND U18954 ( .A(n17205), .B(n17204), .Z(n17200) );
  XOR U18955 ( .A(n1809), .B(n1808), .Z(\A1[197] ) );
  XOR U18956 ( .A(n17205), .B(n17206), .Z(n1808) );
  XNOR U18957 ( .A(n17204), .B(n17202), .Z(n17206) );
  AND U18958 ( .A(n17207), .B(n17208), .Z(n17202) );
  NANDN U18959 ( .A(n17209), .B(n17210), .Z(n17208) );
  NANDN U18960 ( .A(n17211), .B(n17212), .Z(n17210) );
  AND U18961 ( .A(B[196]), .B(A[3]), .Z(n17204) );
  XNOR U18962 ( .A(n17194), .B(n17213), .Z(n17205) );
  XNOR U18963 ( .A(n17192), .B(n17195), .Z(n17213) );
  NAND U18964 ( .A(A[2]), .B(B[197]), .Z(n17195) );
  NANDN U18965 ( .A(n17214), .B(n17215), .Z(n17192) );
  AND U18966 ( .A(A[0]), .B(B[198]), .Z(n17215) );
  XOR U18967 ( .A(n17197), .B(n17216), .Z(n17194) );
  NAND U18968 ( .A(A[0]), .B(B[199]), .Z(n17216) );
  NAND U18969 ( .A(B[198]), .B(A[1]), .Z(n17197) );
  NAND U18970 ( .A(n17217), .B(n17218), .Z(n1809) );
  NANDN U18971 ( .A(n17219), .B(n17220), .Z(n17218) );
  OR U18972 ( .A(n17221), .B(n17222), .Z(n17220) );
  NAND U18973 ( .A(n17222), .B(n17221), .Z(n17217) );
  XOR U18974 ( .A(n1811), .B(n1810), .Z(\A1[196] ) );
  XOR U18975 ( .A(n17222), .B(n17223), .Z(n1810) );
  XNOR U18976 ( .A(n17221), .B(n17219), .Z(n17223) );
  AND U18977 ( .A(n17224), .B(n17225), .Z(n17219) );
  NANDN U18978 ( .A(n17226), .B(n17227), .Z(n17225) );
  NANDN U18979 ( .A(n17228), .B(n17229), .Z(n17227) );
  AND U18980 ( .A(B[195]), .B(A[3]), .Z(n17221) );
  XNOR U18981 ( .A(n17211), .B(n17230), .Z(n17222) );
  XNOR U18982 ( .A(n17209), .B(n17212), .Z(n17230) );
  NAND U18983 ( .A(A[2]), .B(B[196]), .Z(n17212) );
  NANDN U18984 ( .A(n17231), .B(n17232), .Z(n17209) );
  AND U18985 ( .A(A[0]), .B(B[197]), .Z(n17232) );
  XOR U18986 ( .A(n17214), .B(n17233), .Z(n17211) );
  NAND U18987 ( .A(A[0]), .B(B[198]), .Z(n17233) );
  NAND U18988 ( .A(B[197]), .B(A[1]), .Z(n17214) );
  NAND U18989 ( .A(n17234), .B(n17235), .Z(n1811) );
  NANDN U18990 ( .A(n17236), .B(n17237), .Z(n17235) );
  OR U18991 ( .A(n17238), .B(n17239), .Z(n17237) );
  NAND U18992 ( .A(n17239), .B(n17238), .Z(n17234) );
  XOR U18993 ( .A(n1813), .B(n1812), .Z(\A1[195] ) );
  XOR U18994 ( .A(n17239), .B(n17240), .Z(n1812) );
  XNOR U18995 ( .A(n17238), .B(n17236), .Z(n17240) );
  AND U18996 ( .A(n17241), .B(n17242), .Z(n17236) );
  NANDN U18997 ( .A(n17243), .B(n17244), .Z(n17242) );
  NANDN U18998 ( .A(n17245), .B(n17246), .Z(n17244) );
  AND U18999 ( .A(B[194]), .B(A[3]), .Z(n17238) );
  XNOR U19000 ( .A(n17228), .B(n17247), .Z(n17239) );
  XNOR U19001 ( .A(n17226), .B(n17229), .Z(n17247) );
  NAND U19002 ( .A(A[2]), .B(B[195]), .Z(n17229) );
  NANDN U19003 ( .A(n17248), .B(n17249), .Z(n17226) );
  AND U19004 ( .A(A[0]), .B(B[196]), .Z(n17249) );
  XOR U19005 ( .A(n17231), .B(n17250), .Z(n17228) );
  NAND U19006 ( .A(A[0]), .B(B[197]), .Z(n17250) );
  NAND U19007 ( .A(B[196]), .B(A[1]), .Z(n17231) );
  NAND U19008 ( .A(n17251), .B(n17252), .Z(n1813) );
  NANDN U19009 ( .A(n17253), .B(n17254), .Z(n17252) );
  OR U19010 ( .A(n17255), .B(n17256), .Z(n17254) );
  NAND U19011 ( .A(n17256), .B(n17255), .Z(n17251) );
  XOR U19012 ( .A(n1815), .B(n1814), .Z(\A1[194] ) );
  XOR U19013 ( .A(n17256), .B(n17257), .Z(n1814) );
  XNOR U19014 ( .A(n17255), .B(n17253), .Z(n17257) );
  AND U19015 ( .A(n17258), .B(n17259), .Z(n17253) );
  NANDN U19016 ( .A(n17260), .B(n17261), .Z(n17259) );
  NANDN U19017 ( .A(n17262), .B(n17263), .Z(n17261) );
  AND U19018 ( .A(B[193]), .B(A[3]), .Z(n17255) );
  XNOR U19019 ( .A(n17245), .B(n17264), .Z(n17256) );
  XNOR U19020 ( .A(n17243), .B(n17246), .Z(n17264) );
  NAND U19021 ( .A(A[2]), .B(B[194]), .Z(n17246) );
  NANDN U19022 ( .A(n17265), .B(n17266), .Z(n17243) );
  AND U19023 ( .A(A[0]), .B(B[195]), .Z(n17266) );
  XOR U19024 ( .A(n17248), .B(n17267), .Z(n17245) );
  NAND U19025 ( .A(A[0]), .B(B[196]), .Z(n17267) );
  NAND U19026 ( .A(B[195]), .B(A[1]), .Z(n17248) );
  NAND U19027 ( .A(n17268), .B(n17269), .Z(n1815) );
  NANDN U19028 ( .A(n17270), .B(n17271), .Z(n17269) );
  OR U19029 ( .A(n17272), .B(n17273), .Z(n17271) );
  NAND U19030 ( .A(n17273), .B(n17272), .Z(n17268) );
  XOR U19031 ( .A(n1817), .B(n1816), .Z(\A1[193] ) );
  XOR U19032 ( .A(n17273), .B(n17274), .Z(n1816) );
  XNOR U19033 ( .A(n17272), .B(n17270), .Z(n17274) );
  AND U19034 ( .A(n17275), .B(n17276), .Z(n17270) );
  NANDN U19035 ( .A(n17277), .B(n17278), .Z(n17276) );
  NANDN U19036 ( .A(n17279), .B(n17280), .Z(n17278) );
  AND U19037 ( .A(B[192]), .B(A[3]), .Z(n17272) );
  XNOR U19038 ( .A(n17262), .B(n17281), .Z(n17273) );
  XNOR U19039 ( .A(n17260), .B(n17263), .Z(n17281) );
  NAND U19040 ( .A(A[2]), .B(B[193]), .Z(n17263) );
  NANDN U19041 ( .A(n17282), .B(n17283), .Z(n17260) );
  AND U19042 ( .A(A[0]), .B(B[194]), .Z(n17283) );
  XOR U19043 ( .A(n17265), .B(n17284), .Z(n17262) );
  NAND U19044 ( .A(A[0]), .B(B[195]), .Z(n17284) );
  NAND U19045 ( .A(B[194]), .B(A[1]), .Z(n17265) );
  NAND U19046 ( .A(n17285), .B(n17286), .Z(n1817) );
  NANDN U19047 ( .A(n17287), .B(n17288), .Z(n17286) );
  OR U19048 ( .A(n17289), .B(n17290), .Z(n17288) );
  NAND U19049 ( .A(n17290), .B(n17289), .Z(n17285) );
  XOR U19050 ( .A(n1819), .B(n1818), .Z(\A1[192] ) );
  XOR U19051 ( .A(n17290), .B(n17291), .Z(n1818) );
  XNOR U19052 ( .A(n17289), .B(n17287), .Z(n17291) );
  AND U19053 ( .A(n17292), .B(n17293), .Z(n17287) );
  NANDN U19054 ( .A(n17294), .B(n17295), .Z(n17293) );
  NANDN U19055 ( .A(n17296), .B(n17297), .Z(n17295) );
  AND U19056 ( .A(B[191]), .B(A[3]), .Z(n17289) );
  XNOR U19057 ( .A(n17279), .B(n17298), .Z(n17290) );
  XNOR U19058 ( .A(n17277), .B(n17280), .Z(n17298) );
  NAND U19059 ( .A(A[2]), .B(B[192]), .Z(n17280) );
  NANDN U19060 ( .A(n17299), .B(n17300), .Z(n17277) );
  AND U19061 ( .A(A[0]), .B(B[193]), .Z(n17300) );
  XOR U19062 ( .A(n17282), .B(n17301), .Z(n17279) );
  NAND U19063 ( .A(A[0]), .B(B[194]), .Z(n17301) );
  NAND U19064 ( .A(B[193]), .B(A[1]), .Z(n17282) );
  NAND U19065 ( .A(n17302), .B(n17303), .Z(n1819) );
  NANDN U19066 ( .A(n17304), .B(n17305), .Z(n17303) );
  OR U19067 ( .A(n17306), .B(n17307), .Z(n17305) );
  NAND U19068 ( .A(n17307), .B(n17306), .Z(n17302) );
  XOR U19069 ( .A(n1821), .B(n1820), .Z(\A1[191] ) );
  XOR U19070 ( .A(n17307), .B(n17308), .Z(n1820) );
  XNOR U19071 ( .A(n17306), .B(n17304), .Z(n17308) );
  AND U19072 ( .A(n17309), .B(n17310), .Z(n17304) );
  NANDN U19073 ( .A(n17311), .B(n17312), .Z(n17310) );
  NANDN U19074 ( .A(n17313), .B(n17314), .Z(n17312) );
  AND U19075 ( .A(B[190]), .B(A[3]), .Z(n17306) );
  XNOR U19076 ( .A(n17296), .B(n17315), .Z(n17307) );
  XNOR U19077 ( .A(n17294), .B(n17297), .Z(n17315) );
  NAND U19078 ( .A(A[2]), .B(B[191]), .Z(n17297) );
  NANDN U19079 ( .A(n17316), .B(n17317), .Z(n17294) );
  AND U19080 ( .A(A[0]), .B(B[192]), .Z(n17317) );
  XOR U19081 ( .A(n17299), .B(n17318), .Z(n17296) );
  NAND U19082 ( .A(A[0]), .B(B[193]), .Z(n17318) );
  NAND U19083 ( .A(B[192]), .B(A[1]), .Z(n17299) );
  NAND U19084 ( .A(n17319), .B(n17320), .Z(n1821) );
  NANDN U19085 ( .A(n17321), .B(n17322), .Z(n17320) );
  OR U19086 ( .A(n17323), .B(n17324), .Z(n17322) );
  NAND U19087 ( .A(n17324), .B(n17323), .Z(n17319) );
  XOR U19088 ( .A(n1823), .B(n1822), .Z(\A1[190] ) );
  XOR U19089 ( .A(n17324), .B(n17325), .Z(n1822) );
  XNOR U19090 ( .A(n17323), .B(n17321), .Z(n17325) );
  AND U19091 ( .A(n17326), .B(n17327), .Z(n17321) );
  NANDN U19092 ( .A(n17328), .B(n17329), .Z(n17327) );
  NANDN U19093 ( .A(n17330), .B(n17331), .Z(n17329) );
  AND U19094 ( .A(B[189]), .B(A[3]), .Z(n17323) );
  XNOR U19095 ( .A(n17313), .B(n17332), .Z(n17324) );
  XNOR U19096 ( .A(n17311), .B(n17314), .Z(n17332) );
  NAND U19097 ( .A(A[2]), .B(B[190]), .Z(n17314) );
  NANDN U19098 ( .A(n17333), .B(n17334), .Z(n17311) );
  AND U19099 ( .A(A[0]), .B(B[191]), .Z(n17334) );
  XOR U19100 ( .A(n17316), .B(n17335), .Z(n17313) );
  NAND U19101 ( .A(A[0]), .B(B[192]), .Z(n17335) );
  NAND U19102 ( .A(B[191]), .B(A[1]), .Z(n17316) );
  NAND U19103 ( .A(n17336), .B(n17337), .Z(n1823) );
  NANDN U19104 ( .A(n17338), .B(n17339), .Z(n17337) );
  OR U19105 ( .A(n17340), .B(n17341), .Z(n17339) );
  NAND U19106 ( .A(n17341), .B(n17340), .Z(n17336) );
  XOR U19107 ( .A(n1805), .B(n1804), .Z(\A1[18] ) );
  XOR U19108 ( .A(n17171), .B(n17342), .Z(n1804) );
  XNOR U19109 ( .A(n17170), .B(n17168), .Z(n17342) );
  AND U19110 ( .A(n17343), .B(n17344), .Z(n17168) );
  NANDN U19111 ( .A(n17345), .B(n17346), .Z(n17344) );
  NANDN U19112 ( .A(n17347), .B(n17348), .Z(n17346) );
  AND U19113 ( .A(B[17]), .B(A[3]), .Z(n17170) );
  XNOR U19114 ( .A(n17160), .B(n17349), .Z(n17171) );
  XNOR U19115 ( .A(n17158), .B(n17161), .Z(n17349) );
  NAND U19116 ( .A(A[2]), .B(B[18]), .Z(n17161) );
  NANDN U19117 ( .A(n17350), .B(n17351), .Z(n17158) );
  AND U19118 ( .A(A[0]), .B(B[19]), .Z(n17351) );
  XOR U19119 ( .A(n17163), .B(n17352), .Z(n17160) );
  NAND U19120 ( .A(A[0]), .B(B[20]), .Z(n17352) );
  NAND U19121 ( .A(B[19]), .B(A[1]), .Z(n17163) );
  NAND U19122 ( .A(n17353), .B(n17354), .Z(n1805) );
  NANDN U19123 ( .A(n17355), .B(n17356), .Z(n17354) );
  OR U19124 ( .A(n17357), .B(n17358), .Z(n17356) );
  NAND U19125 ( .A(n17358), .B(n17357), .Z(n17353) );
  XOR U19126 ( .A(n1825), .B(n1824), .Z(\A1[189] ) );
  XOR U19127 ( .A(n17341), .B(n17359), .Z(n1824) );
  XNOR U19128 ( .A(n17340), .B(n17338), .Z(n17359) );
  AND U19129 ( .A(n17360), .B(n17361), .Z(n17338) );
  NANDN U19130 ( .A(n17362), .B(n17363), .Z(n17361) );
  NANDN U19131 ( .A(n17364), .B(n17365), .Z(n17363) );
  AND U19132 ( .A(B[188]), .B(A[3]), .Z(n17340) );
  XNOR U19133 ( .A(n17330), .B(n17366), .Z(n17341) );
  XNOR U19134 ( .A(n17328), .B(n17331), .Z(n17366) );
  NAND U19135 ( .A(A[2]), .B(B[189]), .Z(n17331) );
  NANDN U19136 ( .A(n17367), .B(n17368), .Z(n17328) );
  AND U19137 ( .A(A[0]), .B(B[190]), .Z(n17368) );
  XOR U19138 ( .A(n17333), .B(n17369), .Z(n17330) );
  NAND U19139 ( .A(A[0]), .B(B[191]), .Z(n17369) );
  NAND U19140 ( .A(B[190]), .B(A[1]), .Z(n17333) );
  NAND U19141 ( .A(n17370), .B(n17371), .Z(n1825) );
  NANDN U19142 ( .A(n17372), .B(n17373), .Z(n17371) );
  OR U19143 ( .A(n17374), .B(n17375), .Z(n17373) );
  NAND U19144 ( .A(n17375), .B(n17374), .Z(n17370) );
  XOR U19145 ( .A(n1829), .B(n1828), .Z(\A1[188] ) );
  XOR U19146 ( .A(n17375), .B(n17376), .Z(n1828) );
  XNOR U19147 ( .A(n17374), .B(n17372), .Z(n17376) );
  AND U19148 ( .A(n17377), .B(n17378), .Z(n17372) );
  NANDN U19149 ( .A(n17379), .B(n17380), .Z(n17378) );
  NANDN U19150 ( .A(n17381), .B(n17382), .Z(n17380) );
  AND U19151 ( .A(B[187]), .B(A[3]), .Z(n17374) );
  XNOR U19152 ( .A(n17364), .B(n17383), .Z(n17375) );
  XNOR U19153 ( .A(n17362), .B(n17365), .Z(n17383) );
  NAND U19154 ( .A(A[2]), .B(B[188]), .Z(n17365) );
  NANDN U19155 ( .A(n17384), .B(n17385), .Z(n17362) );
  AND U19156 ( .A(A[0]), .B(B[189]), .Z(n17385) );
  XOR U19157 ( .A(n17367), .B(n17386), .Z(n17364) );
  NAND U19158 ( .A(A[0]), .B(B[190]), .Z(n17386) );
  NAND U19159 ( .A(B[189]), .B(A[1]), .Z(n17367) );
  NAND U19160 ( .A(n17387), .B(n17388), .Z(n1829) );
  NANDN U19161 ( .A(n17389), .B(n17390), .Z(n17388) );
  OR U19162 ( .A(n17391), .B(n17392), .Z(n17390) );
  NAND U19163 ( .A(n17392), .B(n17391), .Z(n17387) );
  XOR U19164 ( .A(n1831), .B(n1830), .Z(\A1[187] ) );
  XOR U19165 ( .A(n17392), .B(n17393), .Z(n1830) );
  XNOR U19166 ( .A(n17391), .B(n17389), .Z(n17393) );
  AND U19167 ( .A(n17394), .B(n17395), .Z(n17389) );
  NANDN U19168 ( .A(n17396), .B(n17397), .Z(n17395) );
  NANDN U19169 ( .A(n17398), .B(n17399), .Z(n17397) );
  AND U19170 ( .A(B[186]), .B(A[3]), .Z(n17391) );
  XNOR U19171 ( .A(n17381), .B(n17400), .Z(n17392) );
  XNOR U19172 ( .A(n17379), .B(n17382), .Z(n17400) );
  NAND U19173 ( .A(A[2]), .B(B[187]), .Z(n17382) );
  NANDN U19174 ( .A(n17401), .B(n17402), .Z(n17379) );
  AND U19175 ( .A(A[0]), .B(B[188]), .Z(n17402) );
  XOR U19176 ( .A(n17384), .B(n17403), .Z(n17381) );
  NAND U19177 ( .A(A[0]), .B(B[189]), .Z(n17403) );
  NAND U19178 ( .A(B[188]), .B(A[1]), .Z(n17384) );
  NAND U19179 ( .A(n17404), .B(n17405), .Z(n1831) );
  NANDN U19180 ( .A(n17406), .B(n17407), .Z(n17405) );
  OR U19181 ( .A(n17408), .B(n17409), .Z(n17407) );
  NAND U19182 ( .A(n17409), .B(n17408), .Z(n17404) );
  XOR U19183 ( .A(n1833), .B(n1832), .Z(\A1[186] ) );
  XOR U19184 ( .A(n17409), .B(n17410), .Z(n1832) );
  XNOR U19185 ( .A(n17408), .B(n17406), .Z(n17410) );
  AND U19186 ( .A(n17411), .B(n17412), .Z(n17406) );
  NANDN U19187 ( .A(n17413), .B(n17414), .Z(n17412) );
  NANDN U19188 ( .A(n17415), .B(n17416), .Z(n17414) );
  AND U19189 ( .A(B[185]), .B(A[3]), .Z(n17408) );
  XNOR U19190 ( .A(n17398), .B(n17417), .Z(n17409) );
  XNOR U19191 ( .A(n17396), .B(n17399), .Z(n17417) );
  NAND U19192 ( .A(A[2]), .B(B[186]), .Z(n17399) );
  NANDN U19193 ( .A(n17418), .B(n17419), .Z(n17396) );
  AND U19194 ( .A(A[0]), .B(B[187]), .Z(n17419) );
  XOR U19195 ( .A(n17401), .B(n17420), .Z(n17398) );
  NAND U19196 ( .A(A[0]), .B(B[188]), .Z(n17420) );
  NAND U19197 ( .A(B[187]), .B(A[1]), .Z(n17401) );
  NAND U19198 ( .A(n17421), .B(n17422), .Z(n1833) );
  NANDN U19199 ( .A(n17423), .B(n17424), .Z(n17422) );
  OR U19200 ( .A(n17425), .B(n17426), .Z(n17424) );
  NAND U19201 ( .A(n17426), .B(n17425), .Z(n17421) );
  XOR U19202 ( .A(n1835), .B(n1834), .Z(\A1[185] ) );
  XOR U19203 ( .A(n17426), .B(n17427), .Z(n1834) );
  XNOR U19204 ( .A(n17425), .B(n17423), .Z(n17427) );
  AND U19205 ( .A(n17428), .B(n17429), .Z(n17423) );
  NANDN U19206 ( .A(n17430), .B(n17431), .Z(n17429) );
  NANDN U19207 ( .A(n17432), .B(n17433), .Z(n17431) );
  AND U19208 ( .A(B[184]), .B(A[3]), .Z(n17425) );
  XNOR U19209 ( .A(n17415), .B(n17434), .Z(n17426) );
  XNOR U19210 ( .A(n17413), .B(n17416), .Z(n17434) );
  NAND U19211 ( .A(A[2]), .B(B[185]), .Z(n17416) );
  NANDN U19212 ( .A(n17435), .B(n17436), .Z(n17413) );
  AND U19213 ( .A(A[0]), .B(B[186]), .Z(n17436) );
  XOR U19214 ( .A(n17418), .B(n17437), .Z(n17415) );
  NAND U19215 ( .A(A[0]), .B(B[187]), .Z(n17437) );
  NAND U19216 ( .A(B[186]), .B(A[1]), .Z(n17418) );
  NAND U19217 ( .A(n17438), .B(n17439), .Z(n1835) );
  NANDN U19218 ( .A(n17440), .B(n17441), .Z(n17439) );
  OR U19219 ( .A(n17442), .B(n17443), .Z(n17441) );
  NAND U19220 ( .A(n17443), .B(n17442), .Z(n17438) );
  XOR U19221 ( .A(n1837), .B(n1836), .Z(\A1[184] ) );
  XOR U19222 ( .A(n17443), .B(n17444), .Z(n1836) );
  XNOR U19223 ( .A(n17442), .B(n17440), .Z(n17444) );
  AND U19224 ( .A(n17445), .B(n17446), .Z(n17440) );
  NANDN U19225 ( .A(n17447), .B(n17448), .Z(n17446) );
  NANDN U19226 ( .A(n17449), .B(n17450), .Z(n17448) );
  AND U19227 ( .A(B[183]), .B(A[3]), .Z(n17442) );
  XNOR U19228 ( .A(n17432), .B(n17451), .Z(n17443) );
  XNOR U19229 ( .A(n17430), .B(n17433), .Z(n17451) );
  NAND U19230 ( .A(A[2]), .B(B[184]), .Z(n17433) );
  NANDN U19231 ( .A(n17452), .B(n17453), .Z(n17430) );
  AND U19232 ( .A(A[0]), .B(B[185]), .Z(n17453) );
  XOR U19233 ( .A(n17435), .B(n17454), .Z(n17432) );
  NAND U19234 ( .A(A[0]), .B(B[186]), .Z(n17454) );
  NAND U19235 ( .A(B[185]), .B(A[1]), .Z(n17435) );
  NAND U19236 ( .A(n17455), .B(n17456), .Z(n1837) );
  NANDN U19237 ( .A(n17457), .B(n17458), .Z(n17456) );
  OR U19238 ( .A(n17459), .B(n17460), .Z(n17458) );
  NAND U19239 ( .A(n17460), .B(n17459), .Z(n17455) );
  XOR U19240 ( .A(n1839), .B(n1838), .Z(\A1[183] ) );
  XOR U19241 ( .A(n17460), .B(n17461), .Z(n1838) );
  XNOR U19242 ( .A(n17459), .B(n17457), .Z(n17461) );
  AND U19243 ( .A(n17462), .B(n17463), .Z(n17457) );
  NANDN U19244 ( .A(n17464), .B(n17465), .Z(n17463) );
  NANDN U19245 ( .A(n17466), .B(n17467), .Z(n17465) );
  AND U19246 ( .A(B[182]), .B(A[3]), .Z(n17459) );
  XNOR U19247 ( .A(n17449), .B(n17468), .Z(n17460) );
  XNOR U19248 ( .A(n17447), .B(n17450), .Z(n17468) );
  NAND U19249 ( .A(A[2]), .B(B[183]), .Z(n17450) );
  NANDN U19250 ( .A(n17469), .B(n17470), .Z(n17447) );
  AND U19251 ( .A(A[0]), .B(B[184]), .Z(n17470) );
  XOR U19252 ( .A(n17452), .B(n17471), .Z(n17449) );
  NAND U19253 ( .A(A[0]), .B(B[185]), .Z(n17471) );
  NAND U19254 ( .A(B[184]), .B(A[1]), .Z(n17452) );
  NAND U19255 ( .A(n17472), .B(n17473), .Z(n1839) );
  NANDN U19256 ( .A(n17474), .B(n17475), .Z(n17473) );
  OR U19257 ( .A(n17476), .B(n17477), .Z(n17475) );
  NAND U19258 ( .A(n17477), .B(n17476), .Z(n17472) );
  XOR U19259 ( .A(n1841), .B(n1840), .Z(\A1[182] ) );
  XOR U19260 ( .A(n17477), .B(n17478), .Z(n1840) );
  XNOR U19261 ( .A(n17476), .B(n17474), .Z(n17478) );
  AND U19262 ( .A(n17479), .B(n17480), .Z(n17474) );
  NANDN U19263 ( .A(n17481), .B(n17482), .Z(n17480) );
  NANDN U19264 ( .A(n17483), .B(n17484), .Z(n17482) );
  AND U19265 ( .A(B[181]), .B(A[3]), .Z(n17476) );
  XNOR U19266 ( .A(n17466), .B(n17485), .Z(n17477) );
  XNOR U19267 ( .A(n17464), .B(n17467), .Z(n17485) );
  NAND U19268 ( .A(A[2]), .B(B[182]), .Z(n17467) );
  NANDN U19269 ( .A(n17486), .B(n17487), .Z(n17464) );
  AND U19270 ( .A(A[0]), .B(B[183]), .Z(n17487) );
  XOR U19271 ( .A(n17469), .B(n17488), .Z(n17466) );
  NAND U19272 ( .A(A[0]), .B(B[184]), .Z(n17488) );
  NAND U19273 ( .A(B[183]), .B(A[1]), .Z(n17469) );
  NAND U19274 ( .A(n17489), .B(n17490), .Z(n1841) );
  NANDN U19275 ( .A(n17491), .B(n17492), .Z(n17490) );
  OR U19276 ( .A(n17493), .B(n17494), .Z(n17492) );
  NAND U19277 ( .A(n17494), .B(n17493), .Z(n17489) );
  XOR U19278 ( .A(n1843), .B(n1842), .Z(\A1[181] ) );
  XOR U19279 ( .A(n17494), .B(n17495), .Z(n1842) );
  XNOR U19280 ( .A(n17493), .B(n17491), .Z(n17495) );
  AND U19281 ( .A(n17496), .B(n17497), .Z(n17491) );
  NANDN U19282 ( .A(n17498), .B(n17499), .Z(n17497) );
  NANDN U19283 ( .A(n17500), .B(n17501), .Z(n17499) );
  AND U19284 ( .A(B[180]), .B(A[3]), .Z(n17493) );
  XNOR U19285 ( .A(n17483), .B(n17502), .Z(n17494) );
  XNOR U19286 ( .A(n17481), .B(n17484), .Z(n17502) );
  NAND U19287 ( .A(A[2]), .B(B[181]), .Z(n17484) );
  NANDN U19288 ( .A(n17503), .B(n17504), .Z(n17481) );
  AND U19289 ( .A(A[0]), .B(B[182]), .Z(n17504) );
  XOR U19290 ( .A(n17486), .B(n17505), .Z(n17483) );
  NAND U19291 ( .A(A[0]), .B(B[183]), .Z(n17505) );
  NAND U19292 ( .A(B[182]), .B(A[1]), .Z(n17486) );
  NAND U19293 ( .A(n17506), .B(n17507), .Z(n1843) );
  NANDN U19294 ( .A(n17508), .B(n17509), .Z(n17507) );
  OR U19295 ( .A(n17510), .B(n17511), .Z(n17509) );
  NAND U19296 ( .A(n17511), .B(n17510), .Z(n17506) );
  XOR U19297 ( .A(n1845), .B(n1844), .Z(\A1[180] ) );
  XOR U19298 ( .A(n17511), .B(n17512), .Z(n1844) );
  XNOR U19299 ( .A(n17510), .B(n17508), .Z(n17512) );
  AND U19300 ( .A(n17513), .B(n17514), .Z(n17508) );
  NANDN U19301 ( .A(n17515), .B(n17516), .Z(n17514) );
  NANDN U19302 ( .A(n17517), .B(n17518), .Z(n17516) );
  AND U19303 ( .A(B[179]), .B(A[3]), .Z(n17510) );
  XNOR U19304 ( .A(n17500), .B(n17519), .Z(n17511) );
  XNOR U19305 ( .A(n17498), .B(n17501), .Z(n17519) );
  NAND U19306 ( .A(A[2]), .B(B[180]), .Z(n17501) );
  NANDN U19307 ( .A(n17520), .B(n17521), .Z(n17498) );
  AND U19308 ( .A(A[0]), .B(B[181]), .Z(n17521) );
  XOR U19309 ( .A(n17503), .B(n17522), .Z(n17500) );
  NAND U19310 ( .A(A[0]), .B(B[182]), .Z(n17522) );
  NAND U19311 ( .A(B[181]), .B(A[1]), .Z(n17503) );
  NAND U19312 ( .A(n17523), .B(n17524), .Z(n1845) );
  NANDN U19313 ( .A(n17525), .B(n17526), .Z(n17524) );
  OR U19314 ( .A(n17527), .B(n17528), .Z(n17526) );
  NAND U19315 ( .A(n17528), .B(n17527), .Z(n17523) );
  XOR U19316 ( .A(n1827), .B(n1826), .Z(\A1[17] ) );
  XOR U19317 ( .A(n17358), .B(n17529), .Z(n1826) );
  XNOR U19318 ( .A(n17357), .B(n17355), .Z(n17529) );
  AND U19319 ( .A(n17530), .B(n17531), .Z(n17355) );
  NANDN U19320 ( .A(n17532), .B(n17533), .Z(n17531) );
  NANDN U19321 ( .A(n17534), .B(n17535), .Z(n17533) );
  AND U19322 ( .A(B[16]), .B(A[3]), .Z(n17357) );
  XNOR U19323 ( .A(n17347), .B(n17536), .Z(n17358) );
  XNOR U19324 ( .A(n17345), .B(n17348), .Z(n17536) );
  NAND U19325 ( .A(A[2]), .B(B[17]), .Z(n17348) );
  NANDN U19326 ( .A(n17537), .B(n17538), .Z(n17345) );
  AND U19327 ( .A(A[0]), .B(B[18]), .Z(n17538) );
  XOR U19328 ( .A(n17350), .B(n17539), .Z(n17347) );
  NAND U19329 ( .A(A[0]), .B(B[19]), .Z(n17539) );
  NAND U19330 ( .A(B[18]), .B(A[1]), .Z(n17350) );
  NAND U19331 ( .A(n17540), .B(n17541), .Z(n1827) );
  NANDN U19332 ( .A(n17542), .B(n17543), .Z(n17541) );
  OR U19333 ( .A(n17544), .B(n17545), .Z(n17543) );
  NAND U19334 ( .A(n17545), .B(n17544), .Z(n17540) );
  XOR U19335 ( .A(n1847), .B(n1846), .Z(\A1[179] ) );
  XOR U19336 ( .A(n17528), .B(n17546), .Z(n1846) );
  XNOR U19337 ( .A(n17527), .B(n17525), .Z(n17546) );
  AND U19338 ( .A(n17547), .B(n17548), .Z(n17525) );
  NANDN U19339 ( .A(n17549), .B(n17550), .Z(n17548) );
  NANDN U19340 ( .A(n17551), .B(n17552), .Z(n17550) );
  AND U19341 ( .A(B[178]), .B(A[3]), .Z(n17527) );
  XNOR U19342 ( .A(n17517), .B(n17553), .Z(n17528) );
  XNOR U19343 ( .A(n17515), .B(n17518), .Z(n17553) );
  NAND U19344 ( .A(A[2]), .B(B[179]), .Z(n17518) );
  NANDN U19345 ( .A(n17554), .B(n17555), .Z(n17515) );
  AND U19346 ( .A(A[0]), .B(B[180]), .Z(n17555) );
  XOR U19347 ( .A(n17520), .B(n17556), .Z(n17517) );
  NAND U19348 ( .A(A[0]), .B(B[181]), .Z(n17556) );
  NAND U19349 ( .A(B[180]), .B(A[1]), .Z(n17520) );
  NAND U19350 ( .A(n17557), .B(n17558), .Z(n1847) );
  NANDN U19351 ( .A(n17559), .B(n17560), .Z(n17558) );
  OR U19352 ( .A(n17561), .B(n17562), .Z(n17560) );
  NAND U19353 ( .A(n17562), .B(n17561), .Z(n17557) );
  XOR U19354 ( .A(n1851), .B(n1850), .Z(\A1[178] ) );
  XOR U19355 ( .A(n17562), .B(n17563), .Z(n1850) );
  XNOR U19356 ( .A(n17561), .B(n17559), .Z(n17563) );
  AND U19357 ( .A(n17564), .B(n17565), .Z(n17559) );
  NANDN U19358 ( .A(n17566), .B(n17567), .Z(n17565) );
  NANDN U19359 ( .A(n17568), .B(n17569), .Z(n17567) );
  AND U19360 ( .A(B[177]), .B(A[3]), .Z(n17561) );
  XNOR U19361 ( .A(n17551), .B(n17570), .Z(n17562) );
  XNOR U19362 ( .A(n17549), .B(n17552), .Z(n17570) );
  NAND U19363 ( .A(A[2]), .B(B[178]), .Z(n17552) );
  NANDN U19364 ( .A(n17571), .B(n17572), .Z(n17549) );
  AND U19365 ( .A(A[0]), .B(B[179]), .Z(n17572) );
  XOR U19366 ( .A(n17554), .B(n17573), .Z(n17551) );
  NAND U19367 ( .A(A[0]), .B(B[180]), .Z(n17573) );
  NAND U19368 ( .A(B[179]), .B(A[1]), .Z(n17554) );
  NAND U19369 ( .A(n17574), .B(n17575), .Z(n1851) );
  NANDN U19370 ( .A(n17576), .B(n17577), .Z(n17575) );
  OR U19371 ( .A(n17578), .B(n17579), .Z(n17577) );
  NAND U19372 ( .A(n17579), .B(n17578), .Z(n17574) );
  XOR U19373 ( .A(n1853), .B(n1852), .Z(\A1[177] ) );
  XOR U19374 ( .A(n17579), .B(n17580), .Z(n1852) );
  XNOR U19375 ( .A(n17578), .B(n17576), .Z(n17580) );
  AND U19376 ( .A(n17581), .B(n17582), .Z(n17576) );
  NANDN U19377 ( .A(n17583), .B(n17584), .Z(n17582) );
  NANDN U19378 ( .A(n17585), .B(n17586), .Z(n17584) );
  AND U19379 ( .A(B[176]), .B(A[3]), .Z(n17578) );
  XNOR U19380 ( .A(n17568), .B(n17587), .Z(n17579) );
  XNOR U19381 ( .A(n17566), .B(n17569), .Z(n17587) );
  NAND U19382 ( .A(A[2]), .B(B[177]), .Z(n17569) );
  NANDN U19383 ( .A(n17588), .B(n17589), .Z(n17566) );
  AND U19384 ( .A(A[0]), .B(B[178]), .Z(n17589) );
  XOR U19385 ( .A(n17571), .B(n17590), .Z(n17568) );
  NAND U19386 ( .A(A[0]), .B(B[179]), .Z(n17590) );
  NAND U19387 ( .A(B[178]), .B(A[1]), .Z(n17571) );
  NAND U19388 ( .A(n17591), .B(n17592), .Z(n1853) );
  NANDN U19389 ( .A(n17593), .B(n17594), .Z(n17592) );
  OR U19390 ( .A(n17595), .B(n17596), .Z(n17594) );
  NAND U19391 ( .A(n17596), .B(n17595), .Z(n17591) );
  XOR U19392 ( .A(n1855), .B(n1854), .Z(\A1[176] ) );
  XOR U19393 ( .A(n17596), .B(n17597), .Z(n1854) );
  XNOR U19394 ( .A(n17595), .B(n17593), .Z(n17597) );
  AND U19395 ( .A(n17598), .B(n17599), .Z(n17593) );
  NANDN U19396 ( .A(n17600), .B(n17601), .Z(n17599) );
  NANDN U19397 ( .A(n17602), .B(n17603), .Z(n17601) );
  AND U19398 ( .A(B[175]), .B(A[3]), .Z(n17595) );
  XNOR U19399 ( .A(n17585), .B(n17604), .Z(n17596) );
  XNOR U19400 ( .A(n17583), .B(n17586), .Z(n17604) );
  NAND U19401 ( .A(A[2]), .B(B[176]), .Z(n17586) );
  NANDN U19402 ( .A(n17605), .B(n17606), .Z(n17583) );
  AND U19403 ( .A(A[0]), .B(B[177]), .Z(n17606) );
  XOR U19404 ( .A(n17588), .B(n17607), .Z(n17585) );
  NAND U19405 ( .A(A[0]), .B(B[178]), .Z(n17607) );
  NAND U19406 ( .A(B[177]), .B(A[1]), .Z(n17588) );
  NAND U19407 ( .A(n17608), .B(n17609), .Z(n1855) );
  NANDN U19408 ( .A(n17610), .B(n17611), .Z(n17609) );
  OR U19409 ( .A(n17612), .B(n17613), .Z(n17611) );
  NAND U19410 ( .A(n17613), .B(n17612), .Z(n17608) );
  XOR U19411 ( .A(n1857), .B(n1856), .Z(\A1[175] ) );
  XOR U19412 ( .A(n17613), .B(n17614), .Z(n1856) );
  XNOR U19413 ( .A(n17612), .B(n17610), .Z(n17614) );
  AND U19414 ( .A(n17615), .B(n17616), .Z(n17610) );
  NANDN U19415 ( .A(n17617), .B(n17618), .Z(n17616) );
  NANDN U19416 ( .A(n17619), .B(n17620), .Z(n17618) );
  AND U19417 ( .A(B[174]), .B(A[3]), .Z(n17612) );
  XNOR U19418 ( .A(n17602), .B(n17621), .Z(n17613) );
  XNOR U19419 ( .A(n17600), .B(n17603), .Z(n17621) );
  NAND U19420 ( .A(A[2]), .B(B[175]), .Z(n17603) );
  NANDN U19421 ( .A(n17622), .B(n17623), .Z(n17600) );
  AND U19422 ( .A(A[0]), .B(B[176]), .Z(n17623) );
  XOR U19423 ( .A(n17605), .B(n17624), .Z(n17602) );
  NAND U19424 ( .A(A[0]), .B(B[177]), .Z(n17624) );
  NAND U19425 ( .A(B[176]), .B(A[1]), .Z(n17605) );
  NAND U19426 ( .A(n17625), .B(n17626), .Z(n1857) );
  NANDN U19427 ( .A(n17627), .B(n17628), .Z(n17626) );
  OR U19428 ( .A(n17629), .B(n17630), .Z(n17628) );
  NAND U19429 ( .A(n17630), .B(n17629), .Z(n17625) );
  XOR U19430 ( .A(n1859), .B(n1858), .Z(\A1[174] ) );
  XOR U19431 ( .A(n17630), .B(n17631), .Z(n1858) );
  XNOR U19432 ( .A(n17629), .B(n17627), .Z(n17631) );
  AND U19433 ( .A(n17632), .B(n17633), .Z(n17627) );
  NANDN U19434 ( .A(n17634), .B(n17635), .Z(n17633) );
  NANDN U19435 ( .A(n17636), .B(n17637), .Z(n17635) );
  AND U19436 ( .A(B[173]), .B(A[3]), .Z(n17629) );
  XNOR U19437 ( .A(n17619), .B(n17638), .Z(n17630) );
  XNOR U19438 ( .A(n17617), .B(n17620), .Z(n17638) );
  NAND U19439 ( .A(A[2]), .B(B[174]), .Z(n17620) );
  NANDN U19440 ( .A(n17639), .B(n17640), .Z(n17617) );
  AND U19441 ( .A(A[0]), .B(B[175]), .Z(n17640) );
  XOR U19442 ( .A(n17622), .B(n17641), .Z(n17619) );
  NAND U19443 ( .A(A[0]), .B(B[176]), .Z(n17641) );
  NAND U19444 ( .A(B[175]), .B(A[1]), .Z(n17622) );
  NAND U19445 ( .A(n17642), .B(n17643), .Z(n1859) );
  NANDN U19446 ( .A(n17644), .B(n17645), .Z(n17643) );
  OR U19447 ( .A(n17646), .B(n17647), .Z(n17645) );
  NAND U19448 ( .A(n17647), .B(n17646), .Z(n17642) );
  XOR U19449 ( .A(n1861), .B(n1860), .Z(\A1[173] ) );
  XOR U19450 ( .A(n17647), .B(n17648), .Z(n1860) );
  XNOR U19451 ( .A(n17646), .B(n17644), .Z(n17648) );
  AND U19452 ( .A(n17649), .B(n17650), .Z(n17644) );
  NANDN U19453 ( .A(n17651), .B(n17652), .Z(n17650) );
  NANDN U19454 ( .A(n17653), .B(n17654), .Z(n17652) );
  AND U19455 ( .A(B[172]), .B(A[3]), .Z(n17646) );
  XNOR U19456 ( .A(n17636), .B(n17655), .Z(n17647) );
  XNOR U19457 ( .A(n17634), .B(n17637), .Z(n17655) );
  NAND U19458 ( .A(A[2]), .B(B[173]), .Z(n17637) );
  NANDN U19459 ( .A(n17656), .B(n17657), .Z(n17634) );
  AND U19460 ( .A(A[0]), .B(B[174]), .Z(n17657) );
  XOR U19461 ( .A(n17639), .B(n17658), .Z(n17636) );
  NAND U19462 ( .A(A[0]), .B(B[175]), .Z(n17658) );
  NAND U19463 ( .A(B[174]), .B(A[1]), .Z(n17639) );
  NAND U19464 ( .A(n17659), .B(n17660), .Z(n1861) );
  NANDN U19465 ( .A(n17661), .B(n17662), .Z(n17660) );
  OR U19466 ( .A(n17663), .B(n17664), .Z(n17662) );
  NAND U19467 ( .A(n17664), .B(n17663), .Z(n17659) );
  XOR U19468 ( .A(n1863), .B(n1862), .Z(\A1[172] ) );
  XOR U19469 ( .A(n17664), .B(n17665), .Z(n1862) );
  XNOR U19470 ( .A(n17663), .B(n17661), .Z(n17665) );
  AND U19471 ( .A(n17666), .B(n17667), .Z(n17661) );
  NANDN U19472 ( .A(n17668), .B(n17669), .Z(n17667) );
  NANDN U19473 ( .A(n17670), .B(n17671), .Z(n17669) );
  AND U19474 ( .A(B[171]), .B(A[3]), .Z(n17663) );
  XNOR U19475 ( .A(n17653), .B(n17672), .Z(n17664) );
  XNOR U19476 ( .A(n17651), .B(n17654), .Z(n17672) );
  NAND U19477 ( .A(A[2]), .B(B[172]), .Z(n17654) );
  NANDN U19478 ( .A(n17673), .B(n17674), .Z(n17651) );
  AND U19479 ( .A(A[0]), .B(B[173]), .Z(n17674) );
  XOR U19480 ( .A(n17656), .B(n17675), .Z(n17653) );
  NAND U19481 ( .A(A[0]), .B(B[174]), .Z(n17675) );
  NAND U19482 ( .A(B[173]), .B(A[1]), .Z(n17656) );
  NAND U19483 ( .A(n17676), .B(n17677), .Z(n1863) );
  NANDN U19484 ( .A(n17678), .B(n17679), .Z(n17677) );
  OR U19485 ( .A(n17680), .B(n17681), .Z(n17679) );
  NAND U19486 ( .A(n17681), .B(n17680), .Z(n17676) );
  XOR U19487 ( .A(n1865), .B(n1864), .Z(\A1[171] ) );
  XOR U19488 ( .A(n17681), .B(n17682), .Z(n1864) );
  XNOR U19489 ( .A(n17680), .B(n17678), .Z(n17682) );
  AND U19490 ( .A(n17683), .B(n17684), .Z(n17678) );
  NANDN U19491 ( .A(n17685), .B(n17686), .Z(n17684) );
  NANDN U19492 ( .A(n17687), .B(n17688), .Z(n17686) );
  AND U19493 ( .A(B[170]), .B(A[3]), .Z(n17680) );
  XNOR U19494 ( .A(n17670), .B(n17689), .Z(n17681) );
  XNOR U19495 ( .A(n17668), .B(n17671), .Z(n17689) );
  NAND U19496 ( .A(A[2]), .B(B[171]), .Z(n17671) );
  NANDN U19497 ( .A(n17690), .B(n17691), .Z(n17668) );
  AND U19498 ( .A(A[0]), .B(B[172]), .Z(n17691) );
  XOR U19499 ( .A(n17673), .B(n17692), .Z(n17670) );
  NAND U19500 ( .A(A[0]), .B(B[173]), .Z(n17692) );
  NAND U19501 ( .A(B[172]), .B(A[1]), .Z(n17673) );
  NAND U19502 ( .A(n17693), .B(n17694), .Z(n1865) );
  NANDN U19503 ( .A(n17695), .B(n17696), .Z(n17694) );
  OR U19504 ( .A(n17697), .B(n17698), .Z(n17696) );
  NAND U19505 ( .A(n17698), .B(n17697), .Z(n17693) );
  XOR U19506 ( .A(n1867), .B(n1866), .Z(\A1[170] ) );
  XOR U19507 ( .A(n17698), .B(n17699), .Z(n1866) );
  XNOR U19508 ( .A(n17697), .B(n17695), .Z(n17699) );
  AND U19509 ( .A(n17700), .B(n17701), .Z(n17695) );
  NANDN U19510 ( .A(n17702), .B(n17703), .Z(n17701) );
  NANDN U19511 ( .A(n17704), .B(n17705), .Z(n17703) );
  AND U19512 ( .A(B[169]), .B(A[3]), .Z(n17697) );
  XNOR U19513 ( .A(n17687), .B(n17706), .Z(n17698) );
  XNOR U19514 ( .A(n17685), .B(n17688), .Z(n17706) );
  NAND U19515 ( .A(A[2]), .B(B[170]), .Z(n17688) );
  NANDN U19516 ( .A(n17707), .B(n17708), .Z(n17685) );
  AND U19517 ( .A(A[0]), .B(B[171]), .Z(n17708) );
  XOR U19518 ( .A(n17690), .B(n17709), .Z(n17687) );
  NAND U19519 ( .A(A[0]), .B(B[172]), .Z(n17709) );
  NAND U19520 ( .A(B[171]), .B(A[1]), .Z(n17690) );
  NAND U19521 ( .A(n17710), .B(n17711), .Z(n1867) );
  NANDN U19522 ( .A(n17712), .B(n17713), .Z(n17711) );
  OR U19523 ( .A(n17714), .B(n17715), .Z(n17713) );
  NAND U19524 ( .A(n17715), .B(n17714), .Z(n17710) );
  XOR U19525 ( .A(n1849), .B(n1848), .Z(\A1[16] ) );
  XOR U19526 ( .A(n17545), .B(n17716), .Z(n1848) );
  XNOR U19527 ( .A(n17544), .B(n17542), .Z(n17716) );
  AND U19528 ( .A(n17717), .B(n17718), .Z(n17542) );
  NANDN U19529 ( .A(n17719), .B(n17720), .Z(n17718) );
  NANDN U19530 ( .A(n17721), .B(n17722), .Z(n17720) );
  AND U19531 ( .A(B[15]), .B(A[3]), .Z(n17544) );
  XNOR U19532 ( .A(n17534), .B(n17723), .Z(n17545) );
  XNOR U19533 ( .A(n17532), .B(n17535), .Z(n17723) );
  NAND U19534 ( .A(A[2]), .B(B[16]), .Z(n17535) );
  NANDN U19535 ( .A(n17724), .B(n17725), .Z(n17532) );
  AND U19536 ( .A(A[0]), .B(B[17]), .Z(n17725) );
  XOR U19537 ( .A(n17537), .B(n17726), .Z(n17534) );
  NAND U19538 ( .A(A[0]), .B(B[18]), .Z(n17726) );
  NAND U19539 ( .A(B[17]), .B(A[1]), .Z(n17537) );
  NAND U19540 ( .A(n17727), .B(n17728), .Z(n1849) );
  NANDN U19541 ( .A(n17729), .B(n17730), .Z(n17728) );
  OR U19542 ( .A(n17731), .B(n17732), .Z(n17730) );
  NAND U19543 ( .A(n17732), .B(n17731), .Z(n17727) );
  XOR U19544 ( .A(n1869), .B(n1868), .Z(\A1[169] ) );
  XOR U19545 ( .A(n17715), .B(n17733), .Z(n1868) );
  XNOR U19546 ( .A(n17714), .B(n17712), .Z(n17733) );
  AND U19547 ( .A(n17734), .B(n17735), .Z(n17712) );
  NANDN U19548 ( .A(n17736), .B(n17737), .Z(n17735) );
  NANDN U19549 ( .A(n17738), .B(n17739), .Z(n17737) );
  AND U19550 ( .A(B[168]), .B(A[3]), .Z(n17714) );
  XNOR U19551 ( .A(n17704), .B(n17740), .Z(n17715) );
  XNOR U19552 ( .A(n17702), .B(n17705), .Z(n17740) );
  NAND U19553 ( .A(A[2]), .B(B[169]), .Z(n17705) );
  NANDN U19554 ( .A(n17741), .B(n17742), .Z(n17702) );
  AND U19555 ( .A(A[0]), .B(B[170]), .Z(n17742) );
  XOR U19556 ( .A(n17707), .B(n17743), .Z(n17704) );
  NAND U19557 ( .A(A[0]), .B(B[171]), .Z(n17743) );
  NAND U19558 ( .A(B[170]), .B(A[1]), .Z(n17707) );
  NAND U19559 ( .A(n17744), .B(n17745), .Z(n1869) );
  NANDN U19560 ( .A(n17746), .B(n17747), .Z(n17745) );
  OR U19561 ( .A(n17748), .B(n17749), .Z(n17747) );
  NAND U19562 ( .A(n17749), .B(n17748), .Z(n17744) );
  XOR U19563 ( .A(n1873), .B(n1872), .Z(\A1[168] ) );
  XOR U19564 ( .A(n17749), .B(n17750), .Z(n1872) );
  XNOR U19565 ( .A(n17748), .B(n17746), .Z(n17750) );
  AND U19566 ( .A(n17751), .B(n17752), .Z(n17746) );
  NANDN U19567 ( .A(n17753), .B(n17754), .Z(n17752) );
  NANDN U19568 ( .A(n17755), .B(n17756), .Z(n17754) );
  AND U19569 ( .A(B[167]), .B(A[3]), .Z(n17748) );
  XNOR U19570 ( .A(n17738), .B(n17757), .Z(n17749) );
  XNOR U19571 ( .A(n17736), .B(n17739), .Z(n17757) );
  NAND U19572 ( .A(A[2]), .B(B[168]), .Z(n17739) );
  NANDN U19573 ( .A(n17758), .B(n17759), .Z(n17736) );
  AND U19574 ( .A(A[0]), .B(B[169]), .Z(n17759) );
  XOR U19575 ( .A(n17741), .B(n17760), .Z(n17738) );
  NAND U19576 ( .A(A[0]), .B(B[170]), .Z(n17760) );
  NAND U19577 ( .A(B[169]), .B(A[1]), .Z(n17741) );
  NAND U19578 ( .A(n17761), .B(n17762), .Z(n1873) );
  NANDN U19579 ( .A(n17763), .B(n17764), .Z(n17762) );
  OR U19580 ( .A(n17765), .B(n17766), .Z(n17764) );
  NAND U19581 ( .A(n17766), .B(n17765), .Z(n17761) );
  XOR U19582 ( .A(n1875), .B(n1874), .Z(\A1[167] ) );
  XOR U19583 ( .A(n17766), .B(n17767), .Z(n1874) );
  XNOR U19584 ( .A(n17765), .B(n17763), .Z(n17767) );
  AND U19585 ( .A(n17768), .B(n17769), .Z(n17763) );
  NANDN U19586 ( .A(n17770), .B(n17771), .Z(n17769) );
  NANDN U19587 ( .A(n17772), .B(n17773), .Z(n17771) );
  AND U19588 ( .A(B[166]), .B(A[3]), .Z(n17765) );
  XNOR U19589 ( .A(n17755), .B(n17774), .Z(n17766) );
  XNOR U19590 ( .A(n17753), .B(n17756), .Z(n17774) );
  NAND U19591 ( .A(A[2]), .B(B[167]), .Z(n17756) );
  NANDN U19592 ( .A(n17775), .B(n17776), .Z(n17753) );
  AND U19593 ( .A(A[0]), .B(B[168]), .Z(n17776) );
  XOR U19594 ( .A(n17758), .B(n17777), .Z(n17755) );
  NAND U19595 ( .A(A[0]), .B(B[169]), .Z(n17777) );
  NAND U19596 ( .A(B[168]), .B(A[1]), .Z(n17758) );
  NAND U19597 ( .A(n17778), .B(n17779), .Z(n1875) );
  NANDN U19598 ( .A(n17780), .B(n17781), .Z(n17779) );
  OR U19599 ( .A(n17782), .B(n17783), .Z(n17781) );
  NAND U19600 ( .A(n17783), .B(n17782), .Z(n17778) );
  XOR U19601 ( .A(n1877), .B(n1876), .Z(\A1[166] ) );
  XOR U19602 ( .A(n17783), .B(n17784), .Z(n1876) );
  XNOR U19603 ( .A(n17782), .B(n17780), .Z(n17784) );
  AND U19604 ( .A(n17785), .B(n17786), .Z(n17780) );
  NANDN U19605 ( .A(n17787), .B(n17788), .Z(n17786) );
  NANDN U19606 ( .A(n17789), .B(n17790), .Z(n17788) );
  AND U19607 ( .A(B[165]), .B(A[3]), .Z(n17782) );
  XNOR U19608 ( .A(n17772), .B(n17791), .Z(n17783) );
  XNOR U19609 ( .A(n17770), .B(n17773), .Z(n17791) );
  NAND U19610 ( .A(A[2]), .B(B[166]), .Z(n17773) );
  NANDN U19611 ( .A(n17792), .B(n17793), .Z(n17770) );
  AND U19612 ( .A(A[0]), .B(B[167]), .Z(n17793) );
  XOR U19613 ( .A(n17775), .B(n17794), .Z(n17772) );
  NAND U19614 ( .A(A[0]), .B(B[168]), .Z(n17794) );
  NAND U19615 ( .A(B[167]), .B(A[1]), .Z(n17775) );
  NAND U19616 ( .A(n17795), .B(n17796), .Z(n1877) );
  NANDN U19617 ( .A(n17797), .B(n17798), .Z(n17796) );
  OR U19618 ( .A(n17799), .B(n17800), .Z(n17798) );
  NAND U19619 ( .A(n17800), .B(n17799), .Z(n17795) );
  XOR U19620 ( .A(n1879), .B(n1878), .Z(\A1[165] ) );
  XOR U19621 ( .A(n17800), .B(n17801), .Z(n1878) );
  XNOR U19622 ( .A(n17799), .B(n17797), .Z(n17801) );
  AND U19623 ( .A(n17802), .B(n17803), .Z(n17797) );
  NANDN U19624 ( .A(n17804), .B(n17805), .Z(n17803) );
  NANDN U19625 ( .A(n17806), .B(n17807), .Z(n17805) );
  AND U19626 ( .A(B[164]), .B(A[3]), .Z(n17799) );
  XNOR U19627 ( .A(n17789), .B(n17808), .Z(n17800) );
  XNOR U19628 ( .A(n17787), .B(n17790), .Z(n17808) );
  NAND U19629 ( .A(A[2]), .B(B[165]), .Z(n17790) );
  NANDN U19630 ( .A(n17809), .B(n17810), .Z(n17787) );
  AND U19631 ( .A(A[0]), .B(B[166]), .Z(n17810) );
  XOR U19632 ( .A(n17792), .B(n17811), .Z(n17789) );
  NAND U19633 ( .A(A[0]), .B(B[167]), .Z(n17811) );
  NAND U19634 ( .A(B[166]), .B(A[1]), .Z(n17792) );
  NAND U19635 ( .A(n17812), .B(n17813), .Z(n1879) );
  NANDN U19636 ( .A(n17814), .B(n17815), .Z(n17813) );
  OR U19637 ( .A(n17816), .B(n17817), .Z(n17815) );
  NAND U19638 ( .A(n17817), .B(n17816), .Z(n17812) );
  XOR U19639 ( .A(n1881), .B(n1880), .Z(\A1[164] ) );
  XOR U19640 ( .A(n17817), .B(n17818), .Z(n1880) );
  XNOR U19641 ( .A(n17816), .B(n17814), .Z(n17818) );
  AND U19642 ( .A(n17819), .B(n17820), .Z(n17814) );
  NANDN U19643 ( .A(n17821), .B(n17822), .Z(n17820) );
  NANDN U19644 ( .A(n17823), .B(n17824), .Z(n17822) );
  AND U19645 ( .A(B[163]), .B(A[3]), .Z(n17816) );
  XNOR U19646 ( .A(n17806), .B(n17825), .Z(n17817) );
  XNOR U19647 ( .A(n17804), .B(n17807), .Z(n17825) );
  NAND U19648 ( .A(A[2]), .B(B[164]), .Z(n17807) );
  NANDN U19649 ( .A(n17826), .B(n17827), .Z(n17804) );
  AND U19650 ( .A(A[0]), .B(B[165]), .Z(n17827) );
  XOR U19651 ( .A(n17809), .B(n17828), .Z(n17806) );
  NAND U19652 ( .A(A[0]), .B(B[166]), .Z(n17828) );
  NAND U19653 ( .A(B[165]), .B(A[1]), .Z(n17809) );
  NAND U19654 ( .A(n17829), .B(n17830), .Z(n1881) );
  NANDN U19655 ( .A(n17831), .B(n17832), .Z(n17830) );
  OR U19656 ( .A(n17833), .B(n17834), .Z(n17832) );
  NAND U19657 ( .A(n17834), .B(n17833), .Z(n17829) );
  XOR U19658 ( .A(n1883), .B(n1882), .Z(\A1[163] ) );
  XOR U19659 ( .A(n17834), .B(n17835), .Z(n1882) );
  XNOR U19660 ( .A(n17833), .B(n17831), .Z(n17835) );
  AND U19661 ( .A(n17836), .B(n17837), .Z(n17831) );
  NANDN U19662 ( .A(n17838), .B(n17839), .Z(n17837) );
  NANDN U19663 ( .A(n17840), .B(n17841), .Z(n17839) );
  AND U19664 ( .A(B[162]), .B(A[3]), .Z(n17833) );
  XNOR U19665 ( .A(n17823), .B(n17842), .Z(n17834) );
  XNOR U19666 ( .A(n17821), .B(n17824), .Z(n17842) );
  NAND U19667 ( .A(A[2]), .B(B[163]), .Z(n17824) );
  NANDN U19668 ( .A(n17843), .B(n17844), .Z(n17821) );
  AND U19669 ( .A(A[0]), .B(B[164]), .Z(n17844) );
  XOR U19670 ( .A(n17826), .B(n17845), .Z(n17823) );
  NAND U19671 ( .A(A[0]), .B(B[165]), .Z(n17845) );
  NAND U19672 ( .A(B[164]), .B(A[1]), .Z(n17826) );
  NAND U19673 ( .A(n17846), .B(n17847), .Z(n1883) );
  NANDN U19674 ( .A(n17848), .B(n17849), .Z(n17847) );
  OR U19675 ( .A(n17850), .B(n17851), .Z(n17849) );
  NAND U19676 ( .A(n17851), .B(n17850), .Z(n17846) );
  XOR U19677 ( .A(n1885), .B(n1884), .Z(\A1[162] ) );
  XOR U19678 ( .A(n17851), .B(n17852), .Z(n1884) );
  XNOR U19679 ( .A(n17850), .B(n17848), .Z(n17852) );
  AND U19680 ( .A(n17853), .B(n17854), .Z(n17848) );
  NANDN U19681 ( .A(n17855), .B(n17856), .Z(n17854) );
  NANDN U19682 ( .A(n17857), .B(n17858), .Z(n17856) );
  AND U19683 ( .A(B[161]), .B(A[3]), .Z(n17850) );
  XNOR U19684 ( .A(n17840), .B(n17859), .Z(n17851) );
  XNOR U19685 ( .A(n17838), .B(n17841), .Z(n17859) );
  NAND U19686 ( .A(A[2]), .B(B[162]), .Z(n17841) );
  NANDN U19687 ( .A(n17860), .B(n17861), .Z(n17838) );
  AND U19688 ( .A(A[0]), .B(B[163]), .Z(n17861) );
  XOR U19689 ( .A(n17843), .B(n17862), .Z(n17840) );
  NAND U19690 ( .A(A[0]), .B(B[164]), .Z(n17862) );
  NAND U19691 ( .A(B[163]), .B(A[1]), .Z(n17843) );
  NAND U19692 ( .A(n17863), .B(n17864), .Z(n1885) );
  NANDN U19693 ( .A(n17865), .B(n17866), .Z(n17864) );
  OR U19694 ( .A(n17867), .B(n17868), .Z(n17866) );
  NAND U19695 ( .A(n17868), .B(n17867), .Z(n17863) );
  XOR U19696 ( .A(n1887), .B(n1886), .Z(\A1[161] ) );
  XOR U19697 ( .A(n17868), .B(n17869), .Z(n1886) );
  XNOR U19698 ( .A(n17867), .B(n17865), .Z(n17869) );
  AND U19699 ( .A(n17870), .B(n17871), .Z(n17865) );
  NANDN U19700 ( .A(n17872), .B(n17873), .Z(n17871) );
  NANDN U19701 ( .A(n17874), .B(n17875), .Z(n17873) );
  AND U19702 ( .A(B[160]), .B(A[3]), .Z(n17867) );
  XNOR U19703 ( .A(n17857), .B(n17876), .Z(n17868) );
  XNOR U19704 ( .A(n17855), .B(n17858), .Z(n17876) );
  NAND U19705 ( .A(A[2]), .B(B[161]), .Z(n17858) );
  NANDN U19706 ( .A(n17877), .B(n17878), .Z(n17855) );
  AND U19707 ( .A(A[0]), .B(B[162]), .Z(n17878) );
  XOR U19708 ( .A(n17860), .B(n17879), .Z(n17857) );
  NAND U19709 ( .A(A[0]), .B(B[163]), .Z(n17879) );
  NAND U19710 ( .A(B[162]), .B(A[1]), .Z(n17860) );
  NAND U19711 ( .A(n17880), .B(n17881), .Z(n1887) );
  NANDN U19712 ( .A(n17882), .B(n17883), .Z(n17881) );
  OR U19713 ( .A(n17884), .B(n17885), .Z(n17883) );
  NAND U19714 ( .A(n17885), .B(n17884), .Z(n17880) );
  XOR U19715 ( .A(n1889), .B(n1888), .Z(\A1[160] ) );
  XOR U19716 ( .A(n17885), .B(n17886), .Z(n1888) );
  XNOR U19717 ( .A(n17884), .B(n17882), .Z(n17886) );
  AND U19718 ( .A(n17887), .B(n17888), .Z(n17882) );
  NANDN U19719 ( .A(n17889), .B(n17890), .Z(n17888) );
  NANDN U19720 ( .A(n17891), .B(n17892), .Z(n17890) );
  AND U19721 ( .A(B[159]), .B(A[3]), .Z(n17884) );
  XNOR U19722 ( .A(n17874), .B(n17893), .Z(n17885) );
  XNOR U19723 ( .A(n17872), .B(n17875), .Z(n17893) );
  NAND U19724 ( .A(A[2]), .B(B[160]), .Z(n17875) );
  NANDN U19725 ( .A(n17894), .B(n17895), .Z(n17872) );
  AND U19726 ( .A(A[0]), .B(B[161]), .Z(n17895) );
  XOR U19727 ( .A(n17877), .B(n17896), .Z(n17874) );
  NAND U19728 ( .A(A[0]), .B(B[162]), .Z(n17896) );
  NAND U19729 ( .A(B[161]), .B(A[1]), .Z(n17877) );
  NAND U19730 ( .A(n17897), .B(n17898), .Z(n1889) );
  NANDN U19731 ( .A(n17899), .B(n17900), .Z(n17898) );
  OR U19732 ( .A(n17901), .B(n17902), .Z(n17900) );
  NAND U19733 ( .A(n17902), .B(n17901), .Z(n17897) );
  XOR U19734 ( .A(n1871), .B(n1870), .Z(\A1[15] ) );
  XOR U19735 ( .A(n17732), .B(n17903), .Z(n1870) );
  XNOR U19736 ( .A(n17731), .B(n17729), .Z(n17903) );
  AND U19737 ( .A(n17904), .B(n17905), .Z(n17729) );
  NANDN U19738 ( .A(n17906), .B(n17907), .Z(n17905) );
  NANDN U19739 ( .A(n17908), .B(n17909), .Z(n17907) );
  AND U19740 ( .A(B[14]), .B(A[3]), .Z(n17731) );
  XNOR U19741 ( .A(n17721), .B(n17910), .Z(n17732) );
  XNOR U19742 ( .A(n17719), .B(n17722), .Z(n17910) );
  NAND U19743 ( .A(A[2]), .B(B[15]), .Z(n17722) );
  NANDN U19744 ( .A(n17911), .B(n17912), .Z(n17719) );
  AND U19745 ( .A(A[0]), .B(B[16]), .Z(n17912) );
  XOR U19746 ( .A(n17724), .B(n17913), .Z(n17721) );
  NAND U19747 ( .A(A[0]), .B(B[17]), .Z(n17913) );
  NAND U19748 ( .A(B[16]), .B(A[1]), .Z(n17724) );
  NAND U19749 ( .A(n17914), .B(n17915), .Z(n1871) );
  NANDN U19750 ( .A(n17916), .B(n17917), .Z(n17915) );
  OR U19751 ( .A(n17918), .B(n17919), .Z(n17917) );
  NAND U19752 ( .A(n17919), .B(n17918), .Z(n17914) );
  XOR U19753 ( .A(n1891), .B(n1890), .Z(\A1[159] ) );
  XOR U19754 ( .A(n17902), .B(n17920), .Z(n1890) );
  XNOR U19755 ( .A(n17901), .B(n17899), .Z(n17920) );
  AND U19756 ( .A(n17921), .B(n17922), .Z(n17899) );
  NANDN U19757 ( .A(n17923), .B(n17924), .Z(n17922) );
  NANDN U19758 ( .A(n17925), .B(n17926), .Z(n17924) );
  AND U19759 ( .A(B[158]), .B(A[3]), .Z(n17901) );
  XNOR U19760 ( .A(n17891), .B(n17927), .Z(n17902) );
  XNOR U19761 ( .A(n17889), .B(n17892), .Z(n17927) );
  NAND U19762 ( .A(A[2]), .B(B[159]), .Z(n17892) );
  NANDN U19763 ( .A(n17928), .B(n17929), .Z(n17889) );
  AND U19764 ( .A(A[0]), .B(B[160]), .Z(n17929) );
  XOR U19765 ( .A(n17894), .B(n17930), .Z(n17891) );
  NAND U19766 ( .A(A[0]), .B(B[161]), .Z(n17930) );
  NAND U19767 ( .A(B[160]), .B(A[1]), .Z(n17894) );
  NAND U19768 ( .A(n17931), .B(n17932), .Z(n1891) );
  NANDN U19769 ( .A(n17933), .B(n17934), .Z(n17932) );
  OR U19770 ( .A(n17935), .B(n17936), .Z(n17934) );
  NAND U19771 ( .A(n17936), .B(n17935), .Z(n17931) );
  XOR U19772 ( .A(n1895), .B(n1894), .Z(\A1[158] ) );
  XOR U19773 ( .A(n17936), .B(n17937), .Z(n1894) );
  XNOR U19774 ( .A(n17935), .B(n17933), .Z(n17937) );
  AND U19775 ( .A(n17938), .B(n17939), .Z(n17933) );
  NANDN U19776 ( .A(n17940), .B(n17941), .Z(n17939) );
  NANDN U19777 ( .A(n17942), .B(n17943), .Z(n17941) );
  AND U19778 ( .A(B[157]), .B(A[3]), .Z(n17935) );
  XNOR U19779 ( .A(n17925), .B(n17944), .Z(n17936) );
  XNOR U19780 ( .A(n17923), .B(n17926), .Z(n17944) );
  NAND U19781 ( .A(A[2]), .B(B[158]), .Z(n17926) );
  NANDN U19782 ( .A(n17945), .B(n17946), .Z(n17923) );
  AND U19783 ( .A(A[0]), .B(B[159]), .Z(n17946) );
  XOR U19784 ( .A(n17928), .B(n17947), .Z(n17925) );
  NAND U19785 ( .A(A[0]), .B(B[160]), .Z(n17947) );
  NAND U19786 ( .A(B[159]), .B(A[1]), .Z(n17928) );
  NAND U19787 ( .A(n17948), .B(n17949), .Z(n1895) );
  NANDN U19788 ( .A(n17950), .B(n17951), .Z(n17949) );
  OR U19789 ( .A(n17952), .B(n17953), .Z(n17951) );
  NAND U19790 ( .A(n17953), .B(n17952), .Z(n17948) );
  XOR U19791 ( .A(n1897), .B(n1896), .Z(\A1[157] ) );
  XOR U19792 ( .A(n17953), .B(n17954), .Z(n1896) );
  XNOR U19793 ( .A(n17952), .B(n17950), .Z(n17954) );
  AND U19794 ( .A(n17955), .B(n17956), .Z(n17950) );
  NANDN U19795 ( .A(n17957), .B(n17958), .Z(n17956) );
  NANDN U19796 ( .A(n17959), .B(n17960), .Z(n17958) );
  AND U19797 ( .A(B[156]), .B(A[3]), .Z(n17952) );
  XNOR U19798 ( .A(n17942), .B(n17961), .Z(n17953) );
  XNOR U19799 ( .A(n17940), .B(n17943), .Z(n17961) );
  NAND U19800 ( .A(A[2]), .B(B[157]), .Z(n17943) );
  NANDN U19801 ( .A(n17962), .B(n17963), .Z(n17940) );
  AND U19802 ( .A(A[0]), .B(B[158]), .Z(n17963) );
  XOR U19803 ( .A(n17945), .B(n17964), .Z(n17942) );
  NAND U19804 ( .A(A[0]), .B(B[159]), .Z(n17964) );
  NAND U19805 ( .A(B[158]), .B(A[1]), .Z(n17945) );
  NAND U19806 ( .A(n17965), .B(n17966), .Z(n1897) );
  NANDN U19807 ( .A(n17967), .B(n17968), .Z(n17966) );
  OR U19808 ( .A(n17969), .B(n17970), .Z(n17968) );
  NAND U19809 ( .A(n17970), .B(n17969), .Z(n17965) );
  XOR U19810 ( .A(n1899), .B(n1898), .Z(\A1[156] ) );
  XOR U19811 ( .A(n17970), .B(n17971), .Z(n1898) );
  XNOR U19812 ( .A(n17969), .B(n17967), .Z(n17971) );
  AND U19813 ( .A(n17972), .B(n17973), .Z(n17967) );
  NANDN U19814 ( .A(n17974), .B(n17975), .Z(n17973) );
  NANDN U19815 ( .A(n17976), .B(n17977), .Z(n17975) );
  AND U19816 ( .A(B[155]), .B(A[3]), .Z(n17969) );
  XNOR U19817 ( .A(n17959), .B(n17978), .Z(n17970) );
  XNOR U19818 ( .A(n17957), .B(n17960), .Z(n17978) );
  NAND U19819 ( .A(A[2]), .B(B[156]), .Z(n17960) );
  NANDN U19820 ( .A(n17979), .B(n17980), .Z(n17957) );
  AND U19821 ( .A(A[0]), .B(B[157]), .Z(n17980) );
  XOR U19822 ( .A(n17962), .B(n17981), .Z(n17959) );
  NAND U19823 ( .A(A[0]), .B(B[158]), .Z(n17981) );
  NAND U19824 ( .A(B[157]), .B(A[1]), .Z(n17962) );
  NAND U19825 ( .A(n17982), .B(n17983), .Z(n1899) );
  NANDN U19826 ( .A(n17984), .B(n17985), .Z(n17983) );
  OR U19827 ( .A(n17986), .B(n17987), .Z(n17985) );
  NAND U19828 ( .A(n17987), .B(n17986), .Z(n17982) );
  XOR U19829 ( .A(n1901), .B(n1900), .Z(\A1[155] ) );
  XOR U19830 ( .A(n17987), .B(n17988), .Z(n1900) );
  XNOR U19831 ( .A(n17986), .B(n17984), .Z(n17988) );
  AND U19832 ( .A(n17989), .B(n17990), .Z(n17984) );
  NANDN U19833 ( .A(n17991), .B(n17992), .Z(n17990) );
  NANDN U19834 ( .A(n17993), .B(n17994), .Z(n17992) );
  AND U19835 ( .A(B[154]), .B(A[3]), .Z(n17986) );
  XNOR U19836 ( .A(n17976), .B(n17995), .Z(n17987) );
  XNOR U19837 ( .A(n17974), .B(n17977), .Z(n17995) );
  NAND U19838 ( .A(A[2]), .B(B[155]), .Z(n17977) );
  NANDN U19839 ( .A(n17996), .B(n17997), .Z(n17974) );
  AND U19840 ( .A(A[0]), .B(B[156]), .Z(n17997) );
  XOR U19841 ( .A(n17979), .B(n17998), .Z(n17976) );
  NAND U19842 ( .A(A[0]), .B(B[157]), .Z(n17998) );
  NAND U19843 ( .A(B[156]), .B(A[1]), .Z(n17979) );
  NAND U19844 ( .A(n17999), .B(n18000), .Z(n1901) );
  NANDN U19845 ( .A(n18001), .B(n18002), .Z(n18000) );
  OR U19846 ( .A(n18003), .B(n18004), .Z(n18002) );
  NAND U19847 ( .A(n18004), .B(n18003), .Z(n17999) );
  XOR U19848 ( .A(n1903), .B(n1902), .Z(\A1[154] ) );
  XOR U19849 ( .A(n18004), .B(n18005), .Z(n1902) );
  XNOR U19850 ( .A(n18003), .B(n18001), .Z(n18005) );
  AND U19851 ( .A(n18006), .B(n18007), .Z(n18001) );
  NANDN U19852 ( .A(n18008), .B(n18009), .Z(n18007) );
  NANDN U19853 ( .A(n18010), .B(n18011), .Z(n18009) );
  AND U19854 ( .A(B[153]), .B(A[3]), .Z(n18003) );
  XNOR U19855 ( .A(n17993), .B(n18012), .Z(n18004) );
  XNOR U19856 ( .A(n17991), .B(n17994), .Z(n18012) );
  NAND U19857 ( .A(A[2]), .B(B[154]), .Z(n17994) );
  NANDN U19858 ( .A(n18013), .B(n18014), .Z(n17991) );
  AND U19859 ( .A(A[0]), .B(B[155]), .Z(n18014) );
  XOR U19860 ( .A(n17996), .B(n18015), .Z(n17993) );
  NAND U19861 ( .A(A[0]), .B(B[156]), .Z(n18015) );
  NAND U19862 ( .A(B[155]), .B(A[1]), .Z(n17996) );
  NAND U19863 ( .A(n18016), .B(n18017), .Z(n1903) );
  NANDN U19864 ( .A(n18018), .B(n18019), .Z(n18017) );
  OR U19865 ( .A(n18020), .B(n18021), .Z(n18019) );
  NAND U19866 ( .A(n18021), .B(n18020), .Z(n18016) );
  XOR U19867 ( .A(n1905), .B(n1904), .Z(\A1[153] ) );
  XOR U19868 ( .A(n18021), .B(n18022), .Z(n1904) );
  XNOR U19869 ( .A(n18020), .B(n18018), .Z(n18022) );
  AND U19870 ( .A(n18023), .B(n18024), .Z(n18018) );
  NANDN U19871 ( .A(n18025), .B(n18026), .Z(n18024) );
  NANDN U19872 ( .A(n18027), .B(n18028), .Z(n18026) );
  AND U19873 ( .A(B[152]), .B(A[3]), .Z(n18020) );
  XNOR U19874 ( .A(n18010), .B(n18029), .Z(n18021) );
  XNOR U19875 ( .A(n18008), .B(n18011), .Z(n18029) );
  NAND U19876 ( .A(A[2]), .B(B[153]), .Z(n18011) );
  NANDN U19877 ( .A(n18030), .B(n18031), .Z(n18008) );
  AND U19878 ( .A(A[0]), .B(B[154]), .Z(n18031) );
  XOR U19879 ( .A(n18013), .B(n18032), .Z(n18010) );
  NAND U19880 ( .A(A[0]), .B(B[155]), .Z(n18032) );
  NAND U19881 ( .A(B[154]), .B(A[1]), .Z(n18013) );
  NAND U19882 ( .A(n18033), .B(n18034), .Z(n1905) );
  NANDN U19883 ( .A(n18035), .B(n18036), .Z(n18034) );
  OR U19884 ( .A(n18037), .B(n18038), .Z(n18036) );
  NAND U19885 ( .A(n18038), .B(n18037), .Z(n18033) );
  XOR U19886 ( .A(n1907), .B(n1906), .Z(\A1[152] ) );
  XOR U19887 ( .A(n18038), .B(n18039), .Z(n1906) );
  XNOR U19888 ( .A(n18037), .B(n18035), .Z(n18039) );
  AND U19889 ( .A(n18040), .B(n18041), .Z(n18035) );
  NANDN U19890 ( .A(n18042), .B(n18043), .Z(n18041) );
  NANDN U19891 ( .A(n18044), .B(n18045), .Z(n18043) );
  AND U19892 ( .A(B[151]), .B(A[3]), .Z(n18037) );
  XNOR U19893 ( .A(n18027), .B(n18046), .Z(n18038) );
  XNOR U19894 ( .A(n18025), .B(n18028), .Z(n18046) );
  NAND U19895 ( .A(A[2]), .B(B[152]), .Z(n18028) );
  NANDN U19896 ( .A(n18047), .B(n18048), .Z(n18025) );
  AND U19897 ( .A(A[0]), .B(B[153]), .Z(n18048) );
  XOR U19898 ( .A(n18030), .B(n18049), .Z(n18027) );
  NAND U19899 ( .A(A[0]), .B(B[154]), .Z(n18049) );
  NAND U19900 ( .A(B[153]), .B(A[1]), .Z(n18030) );
  NAND U19901 ( .A(n18050), .B(n18051), .Z(n1907) );
  NANDN U19902 ( .A(n18052), .B(n18053), .Z(n18051) );
  OR U19903 ( .A(n18054), .B(n18055), .Z(n18053) );
  NAND U19904 ( .A(n18055), .B(n18054), .Z(n18050) );
  XOR U19905 ( .A(n1909), .B(n1908), .Z(\A1[151] ) );
  XOR U19906 ( .A(n18055), .B(n18056), .Z(n1908) );
  XNOR U19907 ( .A(n18054), .B(n18052), .Z(n18056) );
  AND U19908 ( .A(n18057), .B(n18058), .Z(n18052) );
  NANDN U19909 ( .A(n18059), .B(n18060), .Z(n18058) );
  NANDN U19910 ( .A(n18061), .B(n18062), .Z(n18060) );
  AND U19911 ( .A(B[150]), .B(A[3]), .Z(n18054) );
  XNOR U19912 ( .A(n18044), .B(n18063), .Z(n18055) );
  XNOR U19913 ( .A(n18042), .B(n18045), .Z(n18063) );
  NAND U19914 ( .A(A[2]), .B(B[151]), .Z(n18045) );
  NANDN U19915 ( .A(n18064), .B(n18065), .Z(n18042) );
  AND U19916 ( .A(A[0]), .B(B[152]), .Z(n18065) );
  XOR U19917 ( .A(n18047), .B(n18066), .Z(n18044) );
  NAND U19918 ( .A(A[0]), .B(B[153]), .Z(n18066) );
  NAND U19919 ( .A(B[152]), .B(A[1]), .Z(n18047) );
  NAND U19920 ( .A(n18067), .B(n18068), .Z(n1909) );
  NANDN U19921 ( .A(n18069), .B(n18070), .Z(n18068) );
  OR U19922 ( .A(n18071), .B(n18072), .Z(n18070) );
  NAND U19923 ( .A(n18072), .B(n18071), .Z(n18067) );
  XOR U19924 ( .A(n1911), .B(n1910), .Z(\A1[150] ) );
  XOR U19925 ( .A(n18072), .B(n18073), .Z(n1910) );
  XNOR U19926 ( .A(n18071), .B(n18069), .Z(n18073) );
  AND U19927 ( .A(n18074), .B(n18075), .Z(n18069) );
  NANDN U19928 ( .A(n18076), .B(n18077), .Z(n18075) );
  NANDN U19929 ( .A(n18078), .B(n18079), .Z(n18077) );
  AND U19930 ( .A(B[149]), .B(A[3]), .Z(n18071) );
  XNOR U19931 ( .A(n18061), .B(n18080), .Z(n18072) );
  XNOR U19932 ( .A(n18059), .B(n18062), .Z(n18080) );
  NAND U19933 ( .A(A[2]), .B(B[150]), .Z(n18062) );
  NANDN U19934 ( .A(n18081), .B(n18082), .Z(n18059) );
  AND U19935 ( .A(A[0]), .B(B[151]), .Z(n18082) );
  XOR U19936 ( .A(n18064), .B(n18083), .Z(n18061) );
  NAND U19937 ( .A(A[0]), .B(B[152]), .Z(n18083) );
  NAND U19938 ( .A(B[151]), .B(A[1]), .Z(n18064) );
  NAND U19939 ( .A(n18084), .B(n18085), .Z(n1911) );
  NANDN U19940 ( .A(n18086), .B(n18087), .Z(n18085) );
  OR U19941 ( .A(n18088), .B(n18089), .Z(n18087) );
  NAND U19942 ( .A(n18089), .B(n18088), .Z(n18084) );
  XOR U19943 ( .A(n1893), .B(n1892), .Z(\A1[14] ) );
  XOR U19944 ( .A(n17919), .B(n18090), .Z(n1892) );
  XNOR U19945 ( .A(n17918), .B(n17916), .Z(n18090) );
  AND U19946 ( .A(n18091), .B(n18092), .Z(n17916) );
  NANDN U19947 ( .A(n18093), .B(n18094), .Z(n18092) );
  NANDN U19948 ( .A(n18095), .B(n18096), .Z(n18094) );
  AND U19949 ( .A(B[13]), .B(A[3]), .Z(n17918) );
  XNOR U19950 ( .A(n17908), .B(n18097), .Z(n17919) );
  XNOR U19951 ( .A(n17906), .B(n17909), .Z(n18097) );
  NAND U19952 ( .A(A[2]), .B(B[14]), .Z(n17909) );
  NANDN U19953 ( .A(n18098), .B(n18099), .Z(n17906) );
  AND U19954 ( .A(A[0]), .B(B[15]), .Z(n18099) );
  XOR U19955 ( .A(n17911), .B(n18100), .Z(n17908) );
  NAND U19956 ( .A(A[0]), .B(B[16]), .Z(n18100) );
  NAND U19957 ( .A(B[15]), .B(A[1]), .Z(n17911) );
  NAND U19958 ( .A(n18101), .B(n18102), .Z(n1893) );
  NANDN U19959 ( .A(n18103), .B(n18104), .Z(n18102) );
  OR U19960 ( .A(n18105), .B(n18106), .Z(n18104) );
  NAND U19961 ( .A(n18106), .B(n18105), .Z(n18101) );
  XOR U19962 ( .A(n1913), .B(n1912), .Z(\A1[149] ) );
  XOR U19963 ( .A(n18089), .B(n18107), .Z(n1912) );
  XNOR U19964 ( .A(n18088), .B(n18086), .Z(n18107) );
  AND U19965 ( .A(n18108), .B(n18109), .Z(n18086) );
  NANDN U19966 ( .A(n18110), .B(n18111), .Z(n18109) );
  NANDN U19967 ( .A(n18112), .B(n18113), .Z(n18111) );
  AND U19968 ( .A(B[148]), .B(A[3]), .Z(n18088) );
  XNOR U19969 ( .A(n18078), .B(n18114), .Z(n18089) );
  XNOR U19970 ( .A(n18076), .B(n18079), .Z(n18114) );
  NAND U19971 ( .A(A[2]), .B(B[149]), .Z(n18079) );
  NANDN U19972 ( .A(n18115), .B(n18116), .Z(n18076) );
  AND U19973 ( .A(A[0]), .B(B[150]), .Z(n18116) );
  XOR U19974 ( .A(n18081), .B(n18117), .Z(n18078) );
  NAND U19975 ( .A(A[0]), .B(B[151]), .Z(n18117) );
  NAND U19976 ( .A(B[150]), .B(A[1]), .Z(n18081) );
  NAND U19977 ( .A(n18118), .B(n18119), .Z(n1913) );
  NANDN U19978 ( .A(n18120), .B(n18121), .Z(n18119) );
  OR U19979 ( .A(n18122), .B(n18123), .Z(n18121) );
  NAND U19980 ( .A(n18123), .B(n18122), .Z(n18118) );
  XOR U19981 ( .A(n1917), .B(n1916), .Z(\A1[148] ) );
  XOR U19982 ( .A(n18123), .B(n18124), .Z(n1916) );
  XNOR U19983 ( .A(n18122), .B(n18120), .Z(n18124) );
  AND U19984 ( .A(n18125), .B(n18126), .Z(n18120) );
  NANDN U19985 ( .A(n18127), .B(n18128), .Z(n18126) );
  NANDN U19986 ( .A(n18129), .B(n18130), .Z(n18128) );
  AND U19987 ( .A(B[147]), .B(A[3]), .Z(n18122) );
  XNOR U19988 ( .A(n18112), .B(n18131), .Z(n18123) );
  XNOR U19989 ( .A(n18110), .B(n18113), .Z(n18131) );
  NAND U19990 ( .A(A[2]), .B(B[148]), .Z(n18113) );
  NANDN U19991 ( .A(n18132), .B(n18133), .Z(n18110) );
  AND U19992 ( .A(A[0]), .B(B[149]), .Z(n18133) );
  XOR U19993 ( .A(n18115), .B(n18134), .Z(n18112) );
  NAND U19994 ( .A(A[0]), .B(B[150]), .Z(n18134) );
  NAND U19995 ( .A(B[149]), .B(A[1]), .Z(n18115) );
  NAND U19996 ( .A(n18135), .B(n18136), .Z(n1917) );
  NANDN U19997 ( .A(n18137), .B(n18138), .Z(n18136) );
  OR U19998 ( .A(n18139), .B(n18140), .Z(n18138) );
  NAND U19999 ( .A(n18140), .B(n18139), .Z(n18135) );
  XOR U20000 ( .A(n1919), .B(n1918), .Z(\A1[147] ) );
  XOR U20001 ( .A(n18140), .B(n18141), .Z(n1918) );
  XNOR U20002 ( .A(n18139), .B(n18137), .Z(n18141) );
  AND U20003 ( .A(n18142), .B(n18143), .Z(n18137) );
  NANDN U20004 ( .A(n18144), .B(n18145), .Z(n18143) );
  NANDN U20005 ( .A(n18146), .B(n18147), .Z(n18145) );
  AND U20006 ( .A(B[146]), .B(A[3]), .Z(n18139) );
  XNOR U20007 ( .A(n18129), .B(n18148), .Z(n18140) );
  XNOR U20008 ( .A(n18127), .B(n18130), .Z(n18148) );
  NAND U20009 ( .A(A[2]), .B(B[147]), .Z(n18130) );
  NANDN U20010 ( .A(n18149), .B(n18150), .Z(n18127) );
  AND U20011 ( .A(A[0]), .B(B[148]), .Z(n18150) );
  XOR U20012 ( .A(n18132), .B(n18151), .Z(n18129) );
  NAND U20013 ( .A(A[0]), .B(B[149]), .Z(n18151) );
  NAND U20014 ( .A(B[148]), .B(A[1]), .Z(n18132) );
  NAND U20015 ( .A(n18152), .B(n18153), .Z(n1919) );
  NANDN U20016 ( .A(n18154), .B(n18155), .Z(n18153) );
  OR U20017 ( .A(n18156), .B(n18157), .Z(n18155) );
  NAND U20018 ( .A(n18157), .B(n18156), .Z(n18152) );
  XOR U20019 ( .A(n1921), .B(n1920), .Z(\A1[146] ) );
  XOR U20020 ( .A(n18157), .B(n18158), .Z(n1920) );
  XNOR U20021 ( .A(n18156), .B(n18154), .Z(n18158) );
  AND U20022 ( .A(n18159), .B(n18160), .Z(n18154) );
  NANDN U20023 ( .A(n18161), .B(n18162), .Z(n18160) );
  NANDN U20024 ( .A(n18163), .B(n18164), .Z(n18162) );
  AND U20025 ( .A(B[145]), .B(A[3]), .Z(n18156) );
  XNOR U20026 ( .A(n18146), .B(n18165), .Z(n18157) );
  XNOR U20027 ( .A(n18144), .B(n18147), .Z(n18165) );
  NAND U20028 ( .A(A[2]), .B(B[146]), .Z(n18147) );
  NANDN U20029 ( .A(n18166), .B(n18167), .Z(n18144) );
  AND U20030 ( .A(A[0]), .B(B[147]), .Z(n18167) );
  XOR U20031 ( .A(n18149), .B(n18168), .Z(n18146) );
  NAND U20032 ( .A(A[0]), .B(B[148]), .Z(n18168) );
  NAND U20033 ( .A(B[147]), .B(A[1]), .Z(n18149) );
  NAND U20034 ( .A(n18169), .B(n18170), .Z(n1921) );
  NANDN U20035 ( .A(n18171), .B(n18172), .Z(n18170) );
  OR U20036 ( .A(n18173), .B(n18174), .Z(n18172) );
  NAND U20037 ( .A(n18174), .B(n18173), .Z(n18169) );
  XOR U20038 ( .A(n1923), .B(n1922), .Z(\A1[145] ) );
  XOR U20039 ( .A(n18174), .B(n18175), .Z(n1922) );
  XNOR U20040 ( .A(n18173), .B(n18171), .Z(n18175) );
  AND U20041 ( .A(n18176), .B(n18177), .Z(n18171) );
  NANDN U20042 ( .A(n18178), .B(n18179), .Z(n18177) );
  NANDN U20043 ( .A(n18180), .B(n18181), .Z(n18179) );
  AND U20044 ( .A(B[144]), .B(A[3]), .Z(n18173) );
  XNOR U20045 ( .A(n18163), .B(n18182), .Z(n18174) );
  XNOR U20046 ( .A(n18161), .B(n18164), .Z(n18182) );
  NAND U20047 ( .A(A[2]), .B(B[145]), .Z(n18164) );
  NANDN U20048 ( .A(n18183), .B(n18184), .Z(n18161) );
  AND U20049 ( .A(A[0]), .B(B[146]), .Z(n18184) );
  XOR U20050 ( .A(n18166), .B(n18185), .Z(n18163) );
  NAND U20051 ( .A(A[0]), .B(B[147]), .Z(n18185) );
  NAND U20052 ( .A(B[146]), .B(A[1]), .Z(n18166) );
  NAND U20053 ( .A(n18186), .B(n18187), .Z(n1923) );
  NANDN U20054 ( .A(n18188), .B(n18189), .Z(n18187) );
  OR U20055 ( .A(n18190), .B(n18191), .Z(n18189) );
  NAND U20056 ( .A(n18191), .B(n18190), .Z(n18186) );
  XOR U20057 ( .A(n1925), .B(n1924), .Z(\A1[144] ) );
  XOR U20058 ( .A(n18191), .B(n18192), .Z(n1924) );
  XNOR U20059 ( .A(n18190), .B(n18188), .Z(n18192) );
  AND U20060 ( .A(n18193), .B(n18194), .Z(n18188) );
  NANDN U20061 ( .A(n18195), .B(n18196), .Z(n18194) );
  NANDN U20062 ( .A(n18197), .B(n18198), .Z(n18196) );
  AND U20063 ( .A(B[143]), .B(A[3]), .Z(n18190) );
  XNOR U20064 ( .A(n18180), .B(n18199), .Z(n18191) );
  XNOR U20065 ( .A(n18178), .B(n18181), .Z(n18199) );
  NAND U20066 ( .A(A[2]), .B(B[144]), .Z(n18181) );
  NANDN U20067 ( .A(n18200), .B(n18201), .Z(n18178) );
  AND U20068 ( .A(A[0]), .B(B[145]), .Z(n18201) );
  XOR U20069 ( .A(n18183), .B(n18202), .Z(n18180) );
  NAND U20070 ( .A(A[0]), .B(B[146]), .Z(n18202) );
  NAND U20071 ( .A(B[145]), .B(A[1]), .Z(n18183) );
  NAND U20072 ( .A(n18203), .B(n18204), .Z(n1925) );
  NANDN U20073 ( .A(n18205), .B(n18206), .Z(n18204) );
  OR U20074 ( .A(n18207), .B(n18208), .Z(n18206) );
  NAND U20075 ( .A(n18208), .B(n18207), .Z(n18203) );
  XOR U20076 ( .A(n1927), .B(n1926), .Z(\A1[143] ) );
  XOR U20077 ( .A(n18208), .B(n18209), .Z(n1926) );
  XNOR U20078 ( .A(n18207), .B(n18205), .Z(n18209) );
  AND U20079 ( .A(n18210), .B(n18211), .Z(n18205) );
  NANDN U20080 ( .A(n18212), .B(n18213), .Z(n18211) );
  NANDN U20081 ( .A(n18214), .B(n18215), .Z(n18213) );
  AND U20082 ( .A(B[142]), .B(A[3]), .Z(n18207) );
  XNOR U20083 ( .A(n18197), .B(n18216), .Z(n18208) );
  XNOR U20084 ( .A(n18195), .B(n18198), .Z(n18216) );
  NAND U20085 ( .A(A[2]), .B(B[143]), .Z(n18198) );
  NANDN U20086 ( .A(n18217), .B(n18218), .Z(n18195) );
  AND U20087 ( .A(A[0]), .B(B[144]), .Z(n18218) );
  XOR U20088 ( .A(n18200), .B(n18219), .Z(n18197) );
  NAND U20089 ( .A(A[0]), .B(B[145]), .Z(n18219) );
  NAND U20090 ( .A(B[144]), .B(A[1]), .Z(n18200) );
  NAND U20091 ( .A(n18220), .B(n18221), .Z(n1927) );
  NANDN U20092 ( .A(n18222), .B(n18223), .Z(n18221) );
  OR U20093 ( .A(n18224), .B(n18225), .Z(n18223) );
  NAND U20094 ( .A(n18225), .B(n18224), .Z(n18220) );
  XOR U20095 ( .A(n1929), .B(n1928), .Z(\A1[142] ) );
  XOR U20096 ( .A(n18225), .B(n18226), .Z(n1928) );
  XNOR U20097 ( .A(n18224), .B(n18222), .Z(n18226) );
  AND U20098 ( .A(n18227), .B(n18228), .Z(n18222) );
  NANDN U20099 ( .A(n18229), .B(n18230), .Z(n18228) );
  NANDN U20100 ( .A(n18231), .B(n18232), .Z(n18230) );
  AND U20101 ( .A(B[141]), .B(A[3]), .Z(n18224) );
  XNOR U20102 ( .A(n18214), .B(n18233), .Z(n18225) );
  XNOR U20103 ( .A(n18212), .B(n18215), .Z(n18233) );
  NAND U20104 ( .A(A[2]), .B(B[142]), .Z(n18215) );
  NANDN U20105 ( .A(n18234), .B(n18235), .Z(n18212) );
  AND U20106 ( .A(A[0]), .B(B[143]), .Z(n18235) );
  XOR U20107 ( .A(n18217), .B(n18236), .Z(n18214) );
  NAND U20108 ( .A(A[0]), .B(B[144]), .Z(n18236) );
  NAND U20109 ( .A(B[143]), .B(A[1]), .Z(n18217) );
  NAND U20110 ( .A(n18237), .B(n18238), .Z(n1929) );
  NANDN U20111 ( .A(n18239), .B(n18240), .Z(n18238) );
  OR U20112 ( .A(n18241), .B(n18242), .Z(n18240) );
  NAND U20113 ( .A(n18242), .B(n18241), .Z(n18237) );
  XOR U20114 ( .A(n1931), .B(n1930), .Z(\A1[141] ) );
  XOR U20115 ( .A(n18242), .B(n18243), .Z(n1930) );
  XNOR U20116 ( .A(n18241), .B(n18239), .Z(n18243) );
  AND U20117 ( .A(n18244), .B(n18245), .Z(n18239) );
  NANDN U20118 ( .A(n18246), .B(n18247), .Z(n18245) );
  NANDN U20119 ( .A(n18248), .B(n18249), .Z(n18247) );
  AND U20120 ( .A(B[140]), .B(A[3]), .Z(n18241) );
  XNOR U20121 ( .A(n18231), .B(n18250), .Z(n18242) );
  XNOR U20122 ( .A(n18229), .B(n18232), .Z(n18250) );
  NAND U20123 ( .A(A[2]), .B(B[141]), .Z(n18232) );
  NANDN U20124 ( .A(n18251), .B(n18252), .Z(n18229) );
  AND U20125 ( .A(A[0]), .B(B[142]), .Z(n18252) );
  XOR U20126 ( .A(n18234), .B(n18253), .Z(n18231) );
  NAND U20127 ( .A(A[0]), .B(B[143]), .Z(n18253) );
  NAND U20128 ( .A(B[142]), .B(A[1]), .Z(n18234) );
  NAND U20129 ( .A(n18254), .B(n18255), .Z(n1931) );
  NANDN U20130 ( .A(n18256), .B(n18257), .Z(n18255) );
  OR U20131 ( .A(n18258), .B(n18259), .Z(n18257) );
  NAND U20132 ( .A(n18259), .B(n18258), .Z(n18254) );
  XOR U20133 ( .A(n1933), .B(n1932), .Z(\A1[140] ) );
  XOR U20134 ( .A(n18259), .B(n18260), .Z(n1932) );
  XNOR U20135 ( .A(n18258), .B(n18256), .Z(n18260) );
  AND U20136 ( .A(n18261), .B(n18262), .Z(n18256) );
  NANDN U20137 ( .A(n18263), .B(n18264), .Z(n18262) );
  NANDN U20138 ( .A(n18265), .B(n18266), .Z(n18264) );
  AND U20139 ( .A(B[139]), .B(A[3]), .Z(n18258) );
  XNOR U20140 ( .A(n18248), .B(n18267), .Z(n18259) );
  XNOR U20141 ( .A(n18246), .B(n18249), .Z(n18267) );
  NAND U20142 ( .A(A[2]), .B(B[140]), .Z(n18249) );
  NANDN U20143 ( .A(n18268), .B(n18269), .Z(n18246) );
  AND U20144 ( .A(A[0]), .B(B[141]), .Z(n18269) );
  XOR U20145 ( .A(n18251), .B(n18270), .Z(n18248) );
  NAND U20146 ( .A(A[0]), .B(B[142]), .Z(n18270) );
  NAND U20147 ( .A(B[141]), .B(A[1]), .Z(n18251) );
  NAND U20148 ( .A(n18271), .B(n18272), .Z(n1933) );
  NANDN U20149 ( .A(n18273), .B(n18274), .Z(n18272) );
  OR U20150 ( .A(n18275), .B(n18276), .Z(n18274) );
  NAND U20151 ( .A(n18276), .B(n18275), .Z(n18271) );
  XOR U20152 ( .A(n1915), .B(n1914), .Z(\A1[13] ) );
  XOR U20153 ( .A(n18106), .B(n18277), .Z(n1914) );
  XNOR U20154 ( .A(n18105), .B(n18103), .Z(n18277) );
  AND U20155 ( .A(n18278), .B(n18279), .Z(n18103) );
  NANDN U20156 ( .A(n18280), .B(n18281), .Z(n18279) );
  NANDN U20157 ( .A(n18282), .B(n18283), .Z(n18281) );
  AND U20158 ( .A(B[12]), .B(A[3]), .Z(n18105) );
  XNOR U20159 ( .A(n18095), .B(n18284), .Z(n18106) );
  XNOR U20160 ( .A(n18093), .B(n18096), .Z(n18284) );
  NAND U20161 ( .A(A[2]), .B(B[13]), .Z(n18096) );
  NANDN U20162 ( .A(n18285), .B(n18286), .Z(n18093) );
  AND U20163 ( .A(A[0]), .B(B[14]), .Z(n18286) );
  XOR U20164 ( .A(n18098), .B(n18287), .Z(n18095) );
  NAND U20165 ( .A(A[0]), .B(B[15]), .Z(n18287) );
  NAND U20166 ( .A(B[14]), .B(A[1]), .Z(n18098) );
  NAND U20167 ( .A(n18288), .B(n18289), .Z(n1915) );
  NANDN U20168 ( .A(n18290), .B(n18291), .Z(n18289) );
  OR U20169 ( .A(n18292), .B(n18293), .Z(n18291) );
  NAND U20170 ( .A(n18293), .B(n18292), .Z(n18288) );
  XOR U20171 ( .A(n1935), .B(n1934), .Z(\A1[139] ) );
  XOR U20172 ( .A(n18276), .B(n18294), .Z(n1934) );
  XNOR U20173 ( .A(n18275), .B(n18273), .Z(n18294) );
  AND U20174 ( .A(n18295), .B(n18296), .Z(n18273) );
  NANDN U20175 ( .A(n18297), .B(n18298), .Z(n18296) );
  NANDN U20176 ( .A(n18299), .B(n18300), .Z(n18298) );
  AND U20177 ( .A(B[138]), .B(A[3]), .Z(n18275) );
  XNOR U20178 ( .A(n18265), .B(n18301), .Z(n18276) );
  XNOR U20179 ( .A(n18263), .B(n18266), .Z(n18301) );
  NAND U20180 ( .A(A[2]), .B(B[139]), .Z(n18266) );
  NANDN U20181 ( .A(n18302), .B(n18303), .Z(n18263) );
  AND U20182 ( .A(A[0]), .B(B[140]), .Z(n18303) );
  XOR U20183 ( .A(n18268), .B(n18304), .Z(n18265) );
  NAND U20184 ( .A(A[0]), .B(B[141]), .Z(n18304) );
  NAND U20185 ( .A(B[140]), .B(A[1]), .Z(n18268) );
  NAND U20186 ( .A(n18305), .B(n18306), .Z(n1935) );
  NANDN U20187 ( .A(n18307), .B(n18308), .Z(n18306) );
  OR U20188 ( .A(n18309), .B(n18310), .Z(n18308) );
  NAND U20189 ( .A(n18310), .B(n18309), .Z(n18305) );
  XOR U20190 ( .A(n1939), .B(n1938), .Z(\A1[138] ) );
  XOR U20191 ( .A(n18310), .B(n18311), .Z(n1938) );
  XNOR U20192 ( .A(n18309), .B(n18307), .Z(n18311) );
  AND U20193 ( .A(n18312), .B(n18313), .Z(n18307) );
  NANDN U20194 ( .A(n18314), .B(n18315), .Z(n18313) );
  NANDN U20195 ( .A(n18316), .B(n18317), .Z(n18315) );
  AND U20196 ( .A(B[137]), .B(A[3]), .Z(n18309) );
  XNOR U20197 ( .A(n18299), .B(n18318), .Z(n18310) );
  XNOR U20198 ( .A(n18297), .B(n18300), .Z(n18318) );
  NAND U20199 ( .A(A[2]), .B(B[138]), .Z(n18300) );
  NANDN U20200 ( .A(n18319), .B(n18320), .Z(n18297) );
  AND U20201 ( .A(A[0]), .B(B[139]), .Z(n18320) );
  XOR U20202 ( .A(n18302), .B(n18321), .Z(n18299) );
  NAND U20203 ( .A(A[0]), .B(B[140]), .Z(n18321) );
  NAND U20204 ( .A(B[139]), .B(A[1]), .Z(n18302) );
  NAND U20205 ( .A(n18322), .B(n18323), .Z(n1939) );
  NANDN U20206 ( .A(n18324), .B(n18325), .Z(n18323) );
  OR U20207 ( .A(n18326), .B(n18327), .Z(n18325) );
  NAND U20208 ( .A(n18327), .B(n18326), .Z(n18322) );
  XOR U20209 ( .A(n1941), .B(n1940), .Z(\A1[137] ) );
  XOR U20210 ( .A(n18327), .B(n18328), .Z(n1940) );
  XNOR U20211 ( .A(n18326), .B(n18324), .Z(n18328) );
  AND U20212 ( .A(n18329), .B(n18330), .Z(n18324) );
  NANDN U20213 ( .A(n18331), .B(n18332), .Z(n18330) );
  NANDN U20214 ( .A(n18333), .B(n18334), .Z(n18332) );
  AND U20215 ( .A(B[136]), .B(A[3]), .Z(n18326) );
  XNOR U20216 ( .A(n18316), .B(n18335), .Z(n18327) );
  XNOR U20217 ( .A(n18314), .B(n18317), .Z(n18335) );
  NAND U20218 ( .A(A[2]), .B(B[137]), .Z(n18317) );
  NANDN U20219 ( .A(n18336), .B(n18337), .Z(n18314) );
  AND U20220 ( .A(A[0]), .B(B[138]), .Z(n18337) );
  XOR U20221 ( .A(n18319), .B(n18338), .Z(n18316) );
  NAND U20222 ( .A(A[0]), .B(B[139]), .Z(n18338) );
  NAND U20223 ( .A(B[138]), .B(A[1]), .Z(n18319) );
  NAND U20224 ( .A(n18339), .B(n18340), .Z(n1941) );
  NANDN U20225 ( .A(n18341), .B(n18342), .Z(n18340) );
  OR U20226 ( .A(n18343), .B(n18344), .Z(n18342) );
  NAND U20227 ( .A(n18344), .B(n18343), .Z(n18339) );
  XOR U20228 ( .A(n1943), .B(n1942), .Z(\A1[136] ) );
  XOR U20229 ( .A(n18344), .B(n18345), .Z(n1942) );
  XNOR U20230 ( .A(n18343), .B(n18341), .Z(n18345) );
  AND U20231 ( .A(n18346), .B(n18347), .Z(n18341) );
  NANDN U20232 ( .A(n18348), .B(n18349), .Z(n18347) );
  NANDN U20233 ( .A(n18350), .B(n18351), .Z(n18349) );
  AND U20234 ( .A(B[135]), .B(A[3]), .Z(n18343) );
  XNOR U20235 ( .A(n18333), .B(n18352), .Z(n18344) );
  XNOR U20236 ( .A(n18331), .B(n18334), .Z(n18352) );
  NAND U20237 ( .A(A[2]), .B(B[136]), .Z(n18334) );
  NANDN U20238 ( .A(n18353), .B(n18354), .Z(n18331) );
  AND U20239 ( .A(A[0]), .B(B[137]), .Z(n18354) );
  XOR U20240 ( .A(n18336), .B(n18355), .Z(n18333) );
  NAND U20241 ( .A(A[0]), .B(B[138]), .Z(n18355) );
  NAND U20242 ( .A(B[137]), .B(A[1]), .Z(n18336) );
  NAND U20243 ( .A(n18356), .B(n18357), .Z(n1943) );
  NANDN U20244 ( .A(n18358), .B(n18359), .Z(n18357) );
  OR U20245 ( .A(n18360), .B(n18361), .Z(n18359) );
  NAND U20246 ( .A(n18361), .B(n18360), .Z(n18356) );
  XOR U20247 ( .A(n1945), .B(n1944), .Z(\A1[135] ) );
  XOR U20248 ( .A(n18361), .B(n18362), .Z(n1944) );
  XNOR U20249 ( .A(n18360), .B(n18358), .Z(n18362) );
  AND U20250 ( .A(n18363), .B(n18364), .Z(n18358) );
  NANDN U20251 ( .A(n18365), .B(n18366), .Z(n18364) );
  NANDN U20252 ( .A(n18367), .B(n18368), .Z(n18366) );
  AND U20253 ( .A(B[134]), .B(A[3]), .Z(n18360) );
  XNOR U20254 ( .A(n18350), .B(n18369), .Z(n18361) );
  XNOR U20255 ( .A(n18348), .B(n18351), .Z(n18369) );
  NAND U20256 ( .A(A[2]), .B(B[135]), .Z(n18351) );
  NANDN U20257 ( .A(n18370), .B(n18371), .Z(n18348) );
  AND U20258 ( .A(A[0]), .B(B[136]), .Z(n18371) );
  XOR U20259 ( .A(n18353), .B(n18372), .Z(n18350) );
  NAND U20260 ( .A(A[0]), .B(B[137]), .Z(n18372) );
  NAND U20261 ( .A(B[136]), .B(A[1]), .Z(n18353) );
  NAND U20262 ( .A(n18373), .B(n18374), .Z(n1945) );
  NANDN U20263 ( .A(n18375), .B(n18376), .Z(n18374) );
  OR U20264 ( .A(n18377), .B(n18378), .Z(n18376) );
  NAND U20265 ( .A(n18378), .B(n18377), .Z(n18373) );
  XOR U20266 ( .A(n1947), .B(n1946), .Z(\A1[134] ) );
  XOR U20267 ( .A(n18378), .B(n18379), .Z(n1946) );
  XNOR U20268 ( .A(n18377), .B(n18375), .Z(n18379) );
  AND U20269 ( .A(n18380), .B(n18381), .Z(n18375) );
  NANDN U20270 ( .A(n18382), .B(n18383), .Z(n18381) );
  NANDN U20271 ( .A(n18384), .B(n18385), .Z(n18383) );
  AND U20272 ( .A(B[133]), .B(A[3]), .Z(n18377) );
  XNOR U20273 ( .A(n18367), .B(n18386), .Z(n18378) );
  XNOR U20274 ( .A(n18365), .B(n18368), .Z(n18386) );
  NAND U20275 ( .A(A[2]), .B(B[134]), .Z(n18368) );
  NANDN U20276 ( .A(n18387), .B(n18388), .Z(n18365) );
  AND U20277 ( .A(A[0]), .B(B[135]), .Z(n18388) );
  XOR U20278 ( .A(n18370), .B(n18389), .Z(n18367) );
  NAND U20279 ( .A(A[0]), .B(B[136]), .Z(n18389) );
  NAND U20280 ( .A(B[135]), .B(A[1]), .Z(n18370) );
  NAND U20281 ( .A(n18390), .B(n18391), .Z(n1947) );
  NANDN U20282 ( .A(n18392), .B(n18393), .Z(n18391) );
  OR U20283 ( .A(n18394), .B(n18395), .Z(n18393) );
  NAND U20284 ( .A(n18395), .B(n18394), .Z(n18390) );
  XOR U20285 ( .A(n1949), .B(n1948), .Z(\A1[133] ) );
  XOR U20286 ( .A(n18395), .B(n18396), .Z(n1948) );
  XNOR U20287 ( .A(n18394), .B(n18392), .Z(n18396) );
  AND U20288 ( .A(n18397), .B(n18398), .Z(n18392) );
  NANDN U20289 ( .A(n18399), .B(n18400), .Z(n18398) );
  NANDN U20290 ( .A(n18401), .B(n18402), .Z(n18400) );
  AND U20291 ( .A(B[132]), .B(A[3]), .Z(n18394) );
  XNOR U20292 ( .A(n18384), .B(n18403), .Z(n18395) );
  XNOR U20293 ( .A(n18382), .B(n18385), .Z(n18403) );
  NAND U20294 ( .A(A[2]), .B(B[133]), .Z(n18385) );
  NANDN U20295 ( .A(n18404), .B(n18405), .Z(n18382) );
  AND U20296 ( .A(A[0]), .B(B[134]), .Z(n18405) );
  XOR U20297 ( .A(n18387), .B(n18406), .Z(n18384) );
  NAND U20298 ( .A(A[0]), .B(B[135]), .Z(n18406) );
  NAND U20299 ( .A(B[134]), .B(A[1]), .Z(n18387) );
  NAND U20300 ( .A(n18407), .B(n18408), .Z(n1949) );
  NANDN U20301 ( .A(n18409), .B(n18410), .Z(n18408) );
  OR U20302 ( .A(n18411), .B(n18412), .Z(n18410) );
  NAND U20303 ( .A(n18412), .B(n18411), .Z(n18407) );
  XOR U20304 ( .A(n1951), .B(n1950), .Z(\A1[132] ) );
  XOR U20305 ( .A(n18412), .B(n18413), .Z(n1950) );
  XNOR U20306 ( .A(n18411), .B(n18409), .Z(n18413) );
  AND U20307 ( .A(n18414), .B(n18415), .Z(n18409) );
  NANDN U20308 ( .A(n18416), .B(n18417), .Z(n18415) );
  NANDN U20309 ( .A(n18418), .B(n18419), .Z(n18417) );
  AND U20310 ( .A(B[131]), .B(A[3]), .Z(n18411) );
  XNOR U20311 ( .A(n18401), .B(n18420), .Z(n18412) );
  XNOR U20312 ( .A(n18399), .B(n18402), .Z(n18420) );
  NAND U20313 ( .A(A[2]), .B(B[132]), .Z(n18402) );
  NANDN U20314 ( .A(n18421), .B(n18422), .Z(n18399) );
  AND U20315 ( .A(A[0]), .B(B[133]), .Z(n18422) );
  XOR U20316 ( .A(n18404), .B(n18423), .Z(n18401) );
  NAND U20317 ( .A(A[0]), .B(B[134]), .Z(n18423) );
  NAND U20318 ( .A(B[133]), .B(A[1]), .Z(n18404) );
  NAND U20319 ( .A(n18424), .B(n18425), .Z(n1951) );
  NANDN U20320 ( .A(n18426), .B(n18427), .Z(n18425) );
  OR U20321 ( .A(n18428), .B(n18429), .Z(n18427) );
  NAND U20322 ( .A(n18429), .B(n18428), .Z(n18424) );
  XOR U20323 ( .A(n1953), .B(n1952), .Z(\A1[131] ) );
  XOR U20324 ( .A(n18429), .B(n18430), .Z(n1952) );
  XNOR U20325 ( .A(n18428), .B(n18426), .Z(n18430) );
  AND U20326 ( .A(n18431), .B(n18432), .Z(n18426) );
  NANDN U20327 ( .A(n18433), .B(n18434), .Z(n18432) );
  NANDN U20328 ( .A(n18435), .B(n18436), .Z(n18434) );
  AND U20329 ( .A(B[130]), .B(A[3]), .Z(n18428) );
  XNOR U20330 ( .A(n18418), .B(n18437), .Z(n18429) );
  XNOR U20331 ( .A(n18416), .B(n18419), .Z(n18437) );
  NAND U20332 ( .A(A[2]), .B(B[131]), .Z(n18419) );
  NANDN U20333 ( .A(n18438), .B(n18439), .Z(n18416) );
  AND U20334 ( .A(A[0]), .B(B[132]), .Z(n18439) );
  XOR U20335 ( .A(n18421), .B(n18440), .Z(n18418) );
  NAND U20336 ( .A(A[0]), .B(B[133]), .Z(n18440) );
  NAND U20337 ( .A(B[132]), .B(A[1]), .Z(n18421) );
  NAND U20338 ( .A(n18441), .B(n18442), .Z(n1953) );
  NANDN U20339 ( .A(n18443), .B(n18444), .Z(n18442) );
  OR U20340 ( .A(n18445), .B(n18446), .Z(n18444) );
  NAND U20341 ( .A(n18446), .B(n18445), .Z(n18441) );
  XOR U20342 ( .A(n1955), .B(n1954), .Z(\A1[130] ) );
  XOR U20343 ( .A(n18446), .B(n18447), .Z(n1954) );
  XNOR U20344 ( .A(n18445), .B(n18443), .Z(n18447) );
  AND U20345 ( .A(n18448), .B(n18449), .Z(n18443) );
  NANDN U20346 ( .A(n18450), .B(n18451), .Z(n18449) );
  NANDN U20347 ( .A(n18452), .B(n18453), .Z(n18451) );
  AND U20348 ( .A(B[129]), .B(A[3]), .Z(n18445) );
  XNOR U20349 ( .A(n18435), .B(n18454), .Z(n18446) );
  XNOR U20350 ( .A(n18433), .B(n18436), .Z(n18454) );
  NAND U20351 ( .A(A[2]), .B(B[130]), .Z(n18436) );
  NANDN U20352 ( .A(n18455), .B(n18456), .Z(n18433) );
  AND U20353 ( .A(A[0]), .B(B[131]), .Z(n18456) );
  XOR U20354 ( .A(n18438), .B(n18457), .Z(n18435) );
  NAND U20355 ( .A(A[0]), .B(B[132]), .Z(n18457) );
  NAND U20356 ( .A(B[131]), .B(A[1]), .Z(n18438) );
  NAND U20357 ( .A(n18458), .B(n18459), .Z(n1955) );
  NANDN U20358 ( .A(n18460), .B(n18461), .Z(n18459) );
  OR U20359 ( .A(n18462), .B(n18463), .Z(n18461) );
  NAND U20360 ( .A(n18463), .B(n18462), .Z(n18458) );
  XOR U20361 ( .A(n1937), .B(n1936), .Z(\A1[12] ) );
  XOR U20362 ( .A(n18293), .B(n18464), .Z(n1936) );
  XNOR U20363 ( .A(n18292), .B(n18290), .Z(n18464) );
  AND U20364 ( .A(n18465), .B(n18466), .Z(n18290) );
  NANDN U20365 ( .A(n18467), .B(n18468), .Z(n18466) );
  NANDN U20366 ( .A(n18469), .B(n18470), .Z(n18468) );
  AND U20367 ( .A(B[11]), .B(A[3]), .Z(n18292) );
  XNOR U20368 ( .A(n18282), .B(n18471), .Z(n18293) );
  XNOR U20369 ( .A(n18280), .B(n18283), .Z(n18471) );
  NAND U20370 ( .A(A[2]), .B(B[12]), .Z(n18283) );
  NANDN U20371 ( .A(n18472), .B(n18473), .Z(n18280) );
  AND U20372 ( .A(A[0]), .B(B[13]), .Z(n18473) );
  XOR U20373 ( .A(n18285), .B(n18474), .Z(n18282) );
  NAND U20374 ( .A(A[0]), .B(B[14]), .Z(n18474) );
  NAND U20375 ( .A(B[13]), .B(A[1]), .Z(n18285) );
  NAND U20376 ( .A(n18475), .B(n18476), .Z(n1937) );
  NANDN U20377 ( .A(n18477), .B(n18478), .Z(n18476) );
  OR U20378 ( .A(n18479), .B(n18480), .Z(n18478) );
  NAND U20379 ( .A(n18480), .B(n18479), .Z(n18475) );
  XOR U20380 ( .A(n1957), .B(n1956), .Z(\A1[129] ) );
  XOR U20381 ( .A(n18463), .B(n18481), .Z(n1956) );
  XNOR U20382 ( .A(n18462), .B(n18460), .Z(n18481) );
  AND U20383 ( .A(n18482), .B(n18483), .Z(n18460) );
  NANDN U20384 ( .A(n18484), .B(n18485), .Z(n18483) );
  NANDN U20385 ( .A(n18486), .B(n18487), .Z(n18485) );
  AND U20386 ( .A(B[128]), .B(A[3]), .Z(n18462) );
  XNOR U20387 ( .A(n18452), .B(n18488), .Z(n18463) );
  XNOR U20388 ( .A(n18450), .B(n18453), .Z(n18488) );
  NAND U20389 ( .A(A[2]), .B(B[129]), .Z(n18453) );
  NANDN U20390 ( .A(n18489), .B(n18490), .Z(n18450) );
  AND U20391 ( .A(A[0]), .B(B[130]), .Z(n18490) );
  XOR U20392 ( .A(n18455), .B(n18491), .Z(n18452) );
  NAND U20393 ( .A(A[0]), .B(B[131]), .Z(n18491) );
  NAND U20394 ( .A(B[130]), .B(A[1]), .Z(n18455) );
  NAND U20395 ( .A(n18492), .B(n18493), .Z(n1957) );
  NANDN U20396 ( .A(n18494), .B(n18495), .Z(n18493) );
  OR U20397 ( .A(n18496), .B(n18497), .Z(n18495) );
  NAND U20398 ( .A(n18497), .B(n18496), .Z(n18492) );
  XOR U20399 ( .A(n1961), .B(n1960), .Z(\A1[128] ) );
  XOR U20400 ( .A(n18497), .B(n18498), .Z(n1960) );
  XNOR U20401 ( .A(n18496), .B(n18494), .Z(n18498) );
  AND U20402 ( .A(n18499), .B(n18500), .Z(n18494) );
  NANDN U20403 ( .A(n18501), .B(n18502), .Z(n18500) );
  NANDN U20404 ( .A(n18503), .B(n18504), .Z(n18502) );
  AND U20405 ( .A(B[127]), .B(A[3]), .Z(n18496) );
  XNOR U20406 ( .A(n18486), .B(n18505), .Z(n18497) );
  XNOR U20407 ( .A(n18484), .B(n18487), .Z(n18505) );
  NAND U20408 ( .A(A[2]), .B(B[128]), .Z(n18487) );
  NANDN U20409 ( .A(n18506), .B(n18507), .Z(n18484) );
  AND U20410 ( .A(A[0]), .B(B[129]), .Z(n18507) );
  XOR U20411 ( .A(n18489), .B(n18508), .Z(n18486) );
  NAND U20412 ( .A(A[0]), .B(B[130]), .Z(n18508) );
  NAND U20413 ( .A(B[129]), .B(A[1]), .Z(n18489) );
  NAND U20414 ( .A(n18509), .B(n18510), .Z(n1961) );
  NANDN U20415 ( .A(n18511), .B(n18512), .Z(n18510) );
  OR U20416 ( .A(n18513), .B(n18514), .Z(n18512) );
  NAND U20417 ( .A(n18514), .B(n18513), .Z(n18509) );
  XOR U20418 ( .A(n1963), .B(n1962), .Z(\A1[127] ) );
  XOR U20419 ( .A(n18514), .B(n18515), .Z(n1962) );
  XNOR U20420 ( .A(n18513), .B(n18511), .Z(n18515) );
  AND U20421 ( .A(n18516), .B(n18517), .Z(n18511) );
  NANDN U20422 ( .A(n18518), .B(n18519), .Z(n18517) );
  NANDN U20423 ( .A(n18520), .B(n18521), .Z(n18519) );
  AND U20424 ( .A(B[126]), .B(A[3]), .Z(n18513) );
  XNOR U20425 ( .A(n18503), .B(n18522), .Z(n18514) );
  XNOR U20426 ( .A(n18501), .B(n18504), .Z(n18522) );
  NAND U20427 ( .A(A[2]), .B(B[127]), .Z(n18504) );
  NANDN U20428 ( .A(n18523), .B(n18524), .Z(n18501) );
  AND U20429 ( .A(A[0]), .B(B[128]), .Z(n18524) );
  XOR U20430 ( .A(n18506), .B(n18525), .Z(n18503) );
  NAND U20431 ( .A(A[0]), .B(B[129]), .Z(n18525) );
  NAND U20432 ( .A(B[128]), .B(A[1]), .Z(n18506) );
  NAND U20433 ( .A(n18526), .B(n18527), .Z(n1963) );
  NANDN U20434 ( .A(n18528), .B(n18529), .Z(n18527) );
  OR U20435 ( .A(n18530), .B(n18531), .Z(n18529) );
  NAND U20436 ( .A(n18531), .B(n18530), .Z(n18526) );
  XOR U20437 ( .A(n1965), .B(n1964), .Z(\A1[126] ) );
  XOR U20438 ( .A(n18531), .B(n18532), .Z(n1964) );
  XNOR U20439 ( .A(n18530), .B(n18528), .Z(n18532) );
  AND U20440 ( .A(n18533), .B(n18534), .Z(n18528) );
  NANDN U20441 ( .A(n18535), .B(n18536), .Z(n18534) );
  NANDN U20442 ( .A(n18537), .B(n18538), .Z(n18536) );
  AND U20443 ( .A(B[125]), .B(A[3]), .Z(n18530) );
  XNOR U20444 ( .A(n18520), .B(n18539), .Z(n18531) );
  XNOR U20445 ( .A(n18518), .B(n18521), .Z(n18539) );
  NAND U20446 ( .A(A[2]), .B(B[126]), .Z(n18521) );
  NANDN U20447 ( .A(n18540), .B(n18541), .Z(n18518) );
  AND U20448 ( .A(A[0]), .B(B[127]), .Z(n18541) );
  XOR U20449 ( .A(n18523), .B(n18542), .Z(n18520) );
  NAND U20450 ( .A(A[0]), .B(B[128]), .Z(n18542) );
  NAND U20451 ( .A(B[127]), .B(A[1]), .Z(n18523) );
  NAND U20452 ( .A(n18543), .B(n18544), .Z(n1965) );
  NANDN U20453 ( .A(n18545), .B(n18546), .Z(n18544) );
  OR U20454 ( .A(n18547), .B(n18548), .Z(n18546) );
  NAND U20455 ( .A(n18548), .B(n18547), .Z(n18543) );
  XOR U20456 ( .A(n1967), .B(n1966), .Z(\A1[125] ) );
  XOR U20457 ( .A(n18548), .B(n18549), .Z(n1966) );
  XNOR U20458 ( .A(n18547), .B(n18545), .Z(n18549) );
  AND U20459 ( .A(n18550), .B(n18551), .Z(n18545) );
  NANDN U20460 ( .A(n18552), .B(n18553), .Z(n18551) );
  NANDN U20461 ( .A(n18554), .B(n18555), .Z(n18553) );
  AND U20462 ( .A(B[124]), .B(A[3]), .Z(n18547) );
  XNOR U20463 ( .A(n18537), .B(n18556), .Z(n18548) );
  XNOR U20464 ( .A(n18535), .B(n18538), .Z(n18556) );
  NAND U20465 ( .A(A[2]), .B(B[125]), .Z(n18538) );
  NANDN U20466 ( .A(n18557), .B(n18558), .Z(n18535) );
  AND U20467 ( .A(A[0]), .B(B[126]), .Z(n18558) );
  XOR U20468 ( .A(n18540), .B(n18559), .Z(n18537) );
  NAND U20469 ( .A(A[0]), .B(B[127]), .Z(n18559) );
  NAND U20470 ( .A(B[126]), .B(A[1]), .Z(n18540) );
  NAND U20471 ( .A(n18560), .B(n18561), .Z(n1967) );
  NANDN U20472 ( .A(n18562), .B(n18563), .Z(n18561) );
  OR U20473 ( .A(n18564), .B(n18565), .Z(n18563) );
  NAND U20474 ( .A(n18565), .B(n18564), .Z(n18560) );
  XOR U20475 ( .A(n1969), .B(n1968), .Z(\A1[124] ) );
  XOR U20476 ( .A(n18565), .B(n18566), .Z(n1968) );
  XNOR U20477 ( .A(n18564), .B(n18562), .Z(n18566) );
  AND U20478 ( .A(n18567), .B(n18568), .Z(n18562) );
  NANDN U20479 ( .A(n18569), .B(n18570), .Z(n18568) );
  NANDN U20480 ( .A(n18571), .B(n18572), .Z(n18570) );
  AND U20481 ( .A(B[123]), .B(A[3]), .Z(n18564) );
  XNOR U20482 ( .A(n18554), .B(n18573), .Z(n18565) );
  XNOR U20483 ( .A(n18552), .B(n18555), .Z(n18573) );
  NAND U20484 ( .A(A[2]), .B(B[124]), .Z(n18555) );
  NANDN U20485 ( .A(n18574), .B(n18575), .Z(n18552) );
  AND U20486 ( .A(A[0]), .B(B[125]), .Z(n18575) );
  XOR U20487 ( .A(n18557), .B(n18576), .Z(n18554) );
  NAND U20488 ( .A(A[0]), .B(B[126]), .Z(n18576) );
  NAND U20489 ( .A(B[125]), .B(A[1]), .Z(n18557) );
  NAND U20490 ( .A(n18577), .B(n18578), .Z(n1969) );
  NANDN U20491 ( .A(n18579), .B(n18580), .Z(n18578) );
  OR U20492 ( .A(n18581), .B(n18582), .Z(n18580) );
  NAND U20493 ( .A(n18582), .B(n18581), .Z(n18577) );
  XOR U20494 ( .A(n1971), .B(n1970), .Z(\A1[123] ) );
  XOR U20495 ( .A(n18582), .B(n18583), .Z(n1970) );
  XNOR U20496 ( .A(n18581), .B(n18579), .Z(n18583) );
  AND U20497 ( .A(n18584), .B(n18585), .Z(n18579) );
  NANDN U20498 ( .A(n18586), .B(n18587), .Z(n18585) );
  NANDN U20499 ( .A(n18588), .B(n18589), .Z(n18587) );
  AND U20500 ( .A(B[122]), .B(A[3]), .Z(n18581) );
  XNOR U20501 ( .A(n18571), .B(n18590), .Z(n18582) );
  XNOR U20502 ( .A(n18569), .B(n18572), .Z(n18590) );
  NAND U20503 ( .A(A[2]), .B(B[123]), .Z(n18572) );
  NANDN U20504 ( .A(n18591), .B(n18592), .Z(n18569) );
  AND U20505 ( .A(A[0]), .B(B[124]), .Z(n18592) );
  XOR U20506 ( .A(n18574), .B(n18593), .Z(n18571) );
  NAND U20507 ( .A(A[0]), .B(B[125]), .Z(n18593) );
  NAND U20508 ( .A(B[124]), .B(A[1]), .Z(n18574) );
  NAND U20509 ( .A(n18594), .B(n18595), .Z(n1971) );
  NANDN U20510 ( .A(n18596), .B(n18597), .Z(n18595) );
  OR U20511 ( .A(n18598), .B(n18599), .Z(n18597) );
  NAND U20512 ( .A(n18599), .B(n18598), .Z(n18594) );
  XOR U20513 ( .A(n1973), .B(n1972), .Z(\A1[122] ) );
  XOR U20514 ( .A(n18599), .B(n18600), .Z(n1972) );
  XNOR U20515 ( .A(n18598), .B(n18596), .Z(n18600) );
  AND U20516 ( .A(n18601), .B(n18602), .Z(n18596) );
  NANDN U20517 ( .A(n18603), .B(n18604), .Z(n18602) );
  NANDN U20518 ( .A(n18605), .B(n18606), .Z(n18604) );
  AND U20519 ( .A(B[121]), .B(A[3]), .Z(n18598) );
  XNOR U20520 ( .A(n18588), .B(n18607), .Z(n18599) );
  XNOR U20521 ( .A(n18586), .B(n18589), .Z(n18607) );
  NAND U20522 ( .A(A[2]), .B(B[122]), .Z(n18589) );
  NANDN U20523 ( .A(n18608), .B(n18609), .Z(n18586) );
  AND U20524 ( .A(A[0]), .B(B[123]), .Z(n18609) );
  XOR U20525 ( .A(n18591), .B(n18610), .Z(n18588) );
  NAND U20526 ( .A(A[0]), .B(B[124]), .Z(n18610) );
  NAND U20527 ( .A(B[123]), .B(A[1]), .Z(n18591) );
  NAND U20528 ( .A(n18611), .B(n18612), .Z(n1973) );
  NANDN U20529 ( .A(n18613), .B(n18614), .Z(n18612) );
  OR U20530 ( .A(n18615), .B(n18616), .Z(n18614) );
  NAND U20531 ( .A(n18616), .B(n18615), .Z(n18611) );
  XOR U20532 ( .A(n1975), .B(n1974), .Z(\A1[121] ) );
  XOR U20533 ( .A(n18616), .B(n18617), .Z(n1974) );
  XNOR U20534 ( .A(n18615), .B(n18613), .Z(n18617) );
  AND U20535 ( .A(n18618), .B(n18619), .Z(n18613) );
  NANDN U20536 ( .A(n18620), .B(n18621), .Z(n18619) );
  NANDN U20537 ( .A(n18622), .B(n18623), .Z(n18621) );
  AND U20538 ( .A(B[120]), .B(A[3]), .Z(n18615) );
  XNOR U20539 ( .A(n18605), .B(n18624), .Z(n18616) );
  XNOR U20540 ( .A(n18603), .B(n18606), .Z(n18624) );
  NAND U20541 ( .A(A[2]), .B(B[121]), .Z(n18606) );
  NANDN U20542 ( .A(n18625), .B(n18626), .Z(n18603) );
  AND U20543 ( .A(A[0]), .B(B[122]), .Z(n18626) );
  XOR U20544 ( .A(n18608), .B(n18627), .Z(n18605) );
  NAND U20545 ( .A(A[0]), .B(B[123]), .Z(n18627) );
  NAND U20546 ( .A(B[122]), .B(A[1]), .Z(n18608) );
  NAND U20547 ( .A(n18628), .B(n18629), .Z(n1975) );
  NANDN U20548 ( .A(n18630), .B(n18631), .Z(n18629) );
  OR U20549 ( .A(n18632), .B(n18633), .Z(n18631) );
  NAND U20550 ( .A(n18633), .B(n18632), .Z(n18628) );
  XOR U20551 ( .A(n1977), .B(n1976), .Z(\A1[120] ) );
  XOR U20552 ( .A(n18633), .B(n18634), .Z(n1976) );
  XNOR U20553 ( .A(n18632), .B(n18630), .Z(n18634) );
  AND U20554 ( .A(n18635), .B(n18636), .Z(n18630) );
  NANDN U20555 ( .A(n18637), .B(n18638), .Z(n18636) );
  NANDN U20556 ( .A(n18639), .B(n18640), .Z(n18638) );
  AND U20557 ( .A(B[119]), .B(A[3]), .Z(n18632) );
  XNOR U20558 ( .A(n18622), .B(n18641), .Z(n18633) );
  XNOR U20559 ( .A(n18620), .B(n18623), .Z(n18641) );
  NAND U20560 ( .A(A[2]), .B(B[120]), .Z(n18623) );
  NANDN U20561 ( .A(n18642), .B(n18643), .Z(n18620) );
  AND U20562 ( .A(A[0]), .B(B[121]), .Z(n18643) );
  XOR U20563 ( .A(n18625), .B(n18644), .Z(n18622) );
  NAND U20564 ( .A(A[0]), .B(B[122]), .Z(n18644) );
  NAND U20565 ( .A(B[121]), .B(A[1]), .Z(n18625) );
  NAND U20566 ( .A(n18645), .B(n18646), .Z(n1977) );
  NANDN U20567 ( .A(n18647), .B(n18648), .Z(n18646) );
  OR U20568 ( .A(n18649), .B(n18650), .Z(n18648) );
  NAND U20569 ( .A(n18650), .B(n18649), .Z(n18645) );
  XOR U20570 ( .A(n1959), .B(n1958), .Z(\A1[11] ) );
  XOR U20571 ( .A(n18480), .B(n18651), .Z(n1958) );
  XNOR U20572 ( .A(n18479), .B(n18477), .Z(n18651) );
  AND U20573 ( .A(n18652), .B(n18653), .Z(n18477) );
  NANDN U20574 ( .A(n18654), .B(n18655), .Z(n18653) );
  NANDN U20575 ( .A(n18656), .B(n18657), .Z(n18655) );
  AND U20576 ( .A(A[3]), .B(B[10]), .Z(n18479) );
  XNOR U20577 ( .A(n18469), .B(n18658), .Z(n18480) );
  XNOR U20578 ( .A(n18467), .B(n18470), .Z(n18658) );
  NAND U20579 ( .A(A[2]), .B(B[11]), .Z(n18470) );
  NANDN U20580 ( .A(n18659), .B(n18660), .Z(n18467) );
  AND U20581 ( .A(A[0]), .B(B[12]), .Z(n18660) );
  XOR U20582 ( .A(n18472), .B(n18661), .Z(n18469) );
  NAND U20583 ( .A(A[0]), .B(B[13]), .Z(n18661) );
  NAND U20584 ( .A(B[12]), .B(A[1]), .Z(n18472) );
  NAND U20585 ( .A(n18662), .B(n18663), .Z(n1959) );
  NANDN U20586 ( .A(n18664), .B(n18665), .Z(n18663) );
  OR U20587 ( .A(n18666), .B(n18667), .Z(n18665) );
  NAND U20588 ( .A(n18667), .B(n18666), .Z(n18662) );
  XOR U20589 ( .A(n1979), .B(n1978), .Z(\A1[119] ) );
  XOR U20590 ( .A(n18650), .B(n18668), .Z(n1978) );
  XNOR U20591 ( .A(n18649), .B(n18647), .Z(n18668) );
  AND U20592 ( .A(n18669), .B(n18670), .Z(n18647) );
  NANDN U20593 ( .A(n18671), .B(n18672), .Z(n18670) );
  NANDN U20594 ( .A(n18673), .B(n18674), .Z(n18672) );
  AND U20595 ( .A(B[118]), .B(A[3]), .Z(n18649) );
  XNOR U20596 ( .A(n18639), .B(n18675), .Z(n18650) );
  XNOR U20597 ( .A(n18637), .B(n18640), .Z(n18675) );
  NAND U20598 ( .A(A[2]), .B(B[119]), .Z(n18640) );
  NANDN U20599 ( .A(n18676), .B(n18677), .Z(n18637) );
  AND U20600 ( .A(A[0]), .B(B[120]), .Z(n18677) );
  XOR U20601 ( .A(n18642), .B(n18678), .Z(n18639) );
  NAND U20602 ( .A(A[0]), .B(B[121]), .Z(n18678) );
  NAND U20603 ( .A(B[120]), .B(A[1]), .Z(n18642) );
  NAND U20604 ( .A(n18679), .B(n18680), .Z(n1979) );
  NANDN U20605 ( .A(n18681), .B(n18682), .Z(n18680) );
  OR U20606 ( .A(n18683), .B(n18684), .Z(n18682) );
  NAND U20607 ( .A(n18684), .B(n18683), .Z(n18679) );
  XOR U20608 ( .A(n1983), .B(n1982), .Z(\A1[118] ) );
  XOR U20609 ( .A(n18684), .B(n18685), .Z(n1982) );
  XNOR U20610 ( .A(n18683), .B(n18681), .Z(n18685) );
  AND U20611 ( .A(n18686), .B(n18687), .Z(n18681) );
  NANDN U20612 ( .A(n18688), .B(n18689), .Z(n18687) );
  NANDN U20613 ( .A(n18690), .B(n18691), .Z(n18689) );
  AND U20614 ( .A(B[117]), .B(A[3]), .Z(n18683) );
  XNOR U20615 ( .A(n18673), .B(n18692), .Z(n18684) );
  XNOR U20616 ( .A(n18671), .B(n18674), .Z(n18692) );
  NAND U20617 ( .A(A[2]), .B(B[118]), .Z(n18674) );
  NANDN U20618 ( .A(n18693), .B(n18694), .Z(n18671) );
  AND U20619 ( .A(A[0]), .B(B[119]), .Z(n18694) );
  XOR U20620 ( .A(n18676), .B(n18695), .Z(n18673) );
  NAND U20621 ( .A(A[0]), .B(B[120]), .Z(n18695) );
  NAND U20622 ( .A(B[119]), .B(A[1]), .Z(n18676) );
  NAND U20623 ( .A(n18696), .B(n18697), .Z(n1983) );
  NANDN U20624 ( .A(n18698), .B(n18699), .Z(n18697) );
  OR U20625 ( .A(n18700), .B(n18701), .Z(n18699) );
  NAND U20626 ( .A(n18701), .B(n18700), .Z(n18696) );
  XOR U20627 ( .A(n1985), .B(n1984), .Z(\A1[117] ) );
  XOR U20628 ( .A(n18701), .B(n18702), .Z(n1984) );
  XNOR U20629 ( .A(n18700), .B(n18698), .Z(n18702) );
  AND U20630 ( .A(n18703), .B(n18704), .Z(n18698) );
  NANDN U20631 ( .A(n18705), .B(n18706), .Z(n18704) );
  NANDN U20632 ( .A(n18707), .B(n18708), .Z(n18706) );
  AND U20633 ( .A(B[116]), .B(A[3]), .Z(n18700) );
  XNOR U20634 ( .A(n18690), .B(n18709), .Z(n18701) );
  XNOR U20635 ( .A(n18688), .B(n18691), .Z(n18709) );
  NAND U20636 ( .A(A[2]), .B(B[117]), .Z(n18691) );
  NANDN U20637 ( .A(n18710), .B(n18711), .Z(n18688) );
  AND U20638 ( .A(A[0]), .B(B[118]), .Z(n18711) );
  XOR U20639 ( .A(n18693), .B(n18712), .Z(n18690) );
  NAND U20640 ( .A(A[0]), .B(B[119]), .Z(n18712) );
  NAND U20641 ( .A(B[118]), .B(A[1]), .Z(n18693) );
  NAND U20642 ( .A(n18713), .B(n18714), .Z(n1985) );
  NANDN U20643 ( .A(n18715), .B(n18716), .Z(n18714) );
  OR U20644 ( .A(n18717), .B(n18718), .Z(n18716) );
  NAND U20645 ( .A(n18718), .B(n18717), .Z(n18713) );
  XOR U20646 ( .A(n1987), .B(n1986), .Z(\A1[116] ) );
  XOR U20647 ( .A(n18718), .B(n18719), .Z(n1986) );
  XNOR U20648 ( .A(n18717), .B(n18715), .Z(n18719) );
  AND U20649 ( .A(n18720), .B(n18721), .Z(n18715) );
  NANDN U20650 ( .A(n18722), .B(n18723), .Z(n18721) );
  NANDN U20651 ( .A(n18724), .B(n18725), .Z(n18723) );
  AND U20652 ( .A(B[115]), .B(A[3]), .Z(n18717) );
  XNOR U20653 ( .A(n18707), .B(n18726), .Z(n18718) );
  XNOR U20654 ( .A(n18705), .B(n18708), .Z(n18726) );
  NAND U20655 ( .A(A[2]), .B(B[116]), .Z(n18708) );
  NANDN U20656 ( .A(n18727), .B(n18728), .Z(n18705) );
  AND U20657 ( .A(A[0]), .B(B[117]), .Z(n18728) );
  XOR U20658 ( .A(n18710), .B(n18729), .Z(n18707) );
  NAND U20659 ( .A(A[0]), .B(B[118]), .Z(n18729) );
  NAND U20660 ( .A(B[117]), .B(A[1]), .Z(n18710) );
  NAND U20661 ( .A(n18730), .B(n18731), .Z(n1987) );
  NANDN U20662 ( .A(n18732), .B(n18733), .Z(n18731) );
  OR U20663 ( .A(n18734), .B(n18735), .Z(n18733) );
  NAND U20664 ( .A(n18735), .B(n18734), .Z(n18730) );
  XOR U20665 ( .A(n1989), .B(n1988), .Z(\A1[115] ) );
  XOR U20666 ( .A(n18735), .B(n18736), .Z(n1988) );
  XNOR U20667 ( .A(n18734), .B(n18732), .Z(n18736) );
  AND U20668 ( .A(n18737), .B(n18738), .Z(n18732) );
  NANDN U20669 ( .A(n18739), .B(n18740), .Z(n18738) );
  NANDN U20670 ( .A(n18741), .B(n18742), .Z(n18740) );
  AND U20671 ( .A(B[114]), .B(A[3]), .Z(n18734) );
  XNOR U20672 ( .A(n18724), .B(n18743), .Z(n18735) );
  XNOR U20673 ( .A(n18722), .B(n18725), .Z(n18743) );
  NAND U20674 ( .A(A[2]), .B(B[115]), .Z(n18725) );
  NANDN U20675 ( .A(n18744), .B(n18745), .Z(n18722) );
  AND U20676 ( .A(A[0]), .B(B[116]), .Z(n18745) );
  XOR U20677 ( .A(n18727), .B(n18746), .Z(n18724) );
  NAND U20678 ( .A(A[0]), .B(B[117]), .Z(n18746) );
  NAND U20679 ( .A(B[116]), .B(A[1]), .Z(n18727) );
  NAND U20680 ( .A(n18747), .B(n18748), .Z(n1989) );
  NANDN U20681 ( .A(n18749), .B(n18750), .Z(n18748) );
  OR U20682 ( .A(n18751), .B(n18752), .Z(n18750) );
  NAND U20683 ( .A(n18752), .B(n18751), .Z(n18747) );
  XOR U20684 ( .A(n1991), .B(n1990), .Z(\A1[114] ) );
  XOR U20685 ( .A(n18752), .B(n18753), .Z(n1990) );
  XNOR U20686 ( .A(n18751), .B(n18749), .Z(n18753) );
  AND U20687 ( .A(n18754), .B(n18755), .Z(n18749) );
  NANDN U20688 ( .A(n18756), .B(n18757), .Z(n18755) );
  NANDN U20689 ( .A(n18758), .B(n18759), .Z(n18757) );
  AND U20690 ( .A(B[113]), .B(A[3]), .Z(n18751) );
  XNOR U20691 ( .A(n18741), .B(n18760), .Z(n18752) );
  XNOR U20692 ( .A(n18739), .B(n18742), .Z(n18760) );
  NAND U20693 ( .A(A[2]), .B(B[114]), .Z(n18742) );
  NANDN U20694 ( .A(n18761), .B(n18762), .Z(n18739) );
  AND U20695 ( .A(A[0]), .B(B[115]), .Z(n18762) );
  XOR U20696 ( .A(n18744), .B(n18763), .Z(n18741) );
  NAND U20697 ( .A(A[0]), .B(B[116]), .Z(n18763) );
  NAND U20698 ( .A(B[115]), .B(A[1]), .Z(n18744) );
  NAND U20699 ( .A(n18764), .B(n18765), .Z(n1991) );
  NANDN U20700 ( .A(n18766), .B(n18767), .Z(n18765) );
  OR U20701 ( .A(n18768), .B(n18769), .Z(n18767) );
  NAND U20702 ( .A(n18769), .B(n18768), .Z(n18764) );
  XOR U20703 ( .A(n1993), .B(n1992), .Z(\A1[113] ) );
  XOR U20704 ( .A(n18769), .B(n18770), .Z(n1992) );
  XNOR U20705 ( .A(n18768), .B(n18766), .Z(n18770) );
  AND U20706 ( .A(n18771), .B(n18772), .Z(n18766) );
  NANDN U20707 ( .A(n18773), .B(n18774), .Z(n18772) );
  NANDN U20708 ( .A(n18775), .B(n18776), .Z(n18774) );
  AND U20709 ( .A(B[112]), .B(A[3]), .Z(n18768) );
  XNOR U20710 ( .A(n18758), .B(n18777), .Z(n18769) );
  XNOR U20711 ( .A(n18756), .B(n18759), .Z(n18777) );
  NAND U20712 ( .A(A[2]), .B(B[113]), .Z(n18759) );
  NANDN U20713 ( .A(n18778), .B(n18779), .Z(n18756) );
  AND U20714 ( .A(A[0]), .B(B[114]), .Z(n18779) );
  XOR U20715 ( .A(n18761), .B(n18780), .Z(n18758) );
  NAND U20716 ( .A(A[0]), .B(B[115]), .Z(n18780) );
  NAND U20717 ( .A(B[114]), .B(A[1]), .Z(n18761) );
  NAND U20718 ( .A(n18781), .B(n18782), .Z(n1993) );
  NANDN U20719 ( .A(n18783), .B(n18784), .Z(n18782) );
  OR U20720 ( .A(n18785), .B(n18786), .Z(n18784) );
  NAND U20721 ( .A(n18786), .B(n18785), .Z(n18781) );
  XOR U20722 ( .A(n1995), .B(n1994), .Z(\A1[112] ) );
  XOR U20723 ( .A(n18786), .B(n18787), .Z(n1994) );
  XNOR U20724 ( .A(n18785), .B(n18783), .Z(n18787) );
  AND U20725 ( .A(n18788), .B(n18789), .Z(n18783) );
  NANDN U20726 ( .A(n18790), .B(n18791), .Z(n18789) );
  NANDN U20727 ( .A(n18792), .B(n18793), .Z(n18791) );
  AND U20728 ( .A(B[111]), .B(A[3]), .Z(n18785) );
  XNOR U20729 ( .A(n18775), .B(n18794), .Z(n18786) );
  XNOR U20730 ( .A(n18773), .B(n18776), .Z(n18794) );
  NAND U20731 ( .A(A[2]), .B(B[112]), .Z(n18776) );
  NANDN U20732 ( .A(n18795), .B(n18796), .Z(n18773) );
  AND U20733 ( .A(A[0]), .B(B[113]), .Z(n18796) );
  XOR U20734 ( .A(n18778), .B(n18797), .Z(n18775) );
  NAND U20735 ( .A(A[0]), .B(B[114]), .Z(n18797) );
  NAND U20736 ( .A(B[113]), .B(A[1]), .Z(n18778) );
  NAND U20737 ( .A(n18798), .B(n18799), .Z(n1995) );
  NANDN U20738 ( .A(n18800), .B(n18801), .Z(n18799) );
  OR U20739 ( .A(n18802), .B(n18803), .Z(n18801) );
  NAND U20740 ( .A(n18803), .B(n18802), .Z(n18798) );
  XOR U20741 ( .A(n1997), .B(n1996), .Z(\A1[111] ) );
  XOR U20742 ( .A(n18803), .B(n18804), .Z(n1996) );
  XNOR U20743 ( .A(n18802), .B(n18800), .Z(n18804) );
  AND U20744 ( .A(n18805), .B(n18806), .Z(n18800) );
  NANDN U20745 ( .A(n18807), .B(n18808), .Z(n18806) );
  NANDN U20746 ( .A(n18809), .B(n18810), .Z(n18808) );
  AND U20747 ( .A(B[110]), .B(A[3]), .Z(n18802) );
  XNOR U20748 ( .A(n18792), .B(n18811), .Z(n18803) );
  XNOR U20749 ( .A(n18790), .B(n18793), .Z(n18811) );
  NAND U20750 ( .A(A[2]), .B(B[111]), .Z(n18793) );
  NANDN U20751 ( .A(n18812), .B(n18813), .Z(n18790) );
  AND U20752 ( .A(A[0]), .B(B[112]), .Z(n18813) );
  XOR U20753 ( .A(n18795), .B(n18814), .Z(n18792) );
  NAND U20754 ( .A(A[0]), .B(B[113]), .Z(n18814) );
  NAND U20755 ( .A(B[112]), .B(A[1]), .Z(n18795) );
  NAND U20756 ( .A(n18815), .B(n18816), .Z(n1997) );
  NANDN U20757 ( .A(n18817), .B(n18818), .Z(n18816) );
  OR U20758 ( .A(n18819), .B(n18820), .Z(n18818) );
  NAND U20759 ( .A(n18820), .B(n18819), .Z(n18815) );
  XOR U20760 ( .A(n1999), .B(n1998), .Z(\A1[110] ) );
  XOR U20761 ( .A(n18820), .B(n18821), .Z(n1998) );
  XNOR U20762 ( .A(n18819), .B(n18817), .Z(n18821) );
  AND U20763 ( .A(n18822), .B(n18823), .Z(n18817) );
  NANDN U20764 ( .A(n18824), .B(n18825), .Z(n18823) );
  NANDN U20765 ( .A(n18826), .B(n18827), .Z(n18825) );
  AND U20766 ( .A(B[109]), .B(A[3]), .Z(n18819) );
  XNOR U20767 ( .A(n18809), .B(n18828), .Z(n18820) );
  XNOR U20768 ( .A(n18807), .B(n18810), .Z(n18828) );
  NAND U20769 ( .A(A[2]), .B(B[110]), .Z(n18810) );
  NANDN U20770 ( .A(n18829), .B(n18830), .Z(n18807) );
  AND U20771 ( .A(A[0]), .B(B[111]), .Z(n18830) );
  XOR U20772 ( .A(n18812), .B(n18831), .Z(n18809) );
  NAND U20773 ( .A(A[0]), .B(B[112]), .Z(n18831) );
  NAND U20774 ( .A(B[111]), .B(A[1]), .Z(n18812) );
  NAND U20775 ( .A(n18832), .B(n18833), .Z(n1999) );
  NANDN U20776 ( .A(n18834), .B(n18835), .Z(n18833) );
  OR U20777 ( .A(n18836), .B(n18837), .Z(n18835) );
  NAND U20778 ( .A(n18837), .B(n18836), .Z(n18832) );
  XOR U20779 ( .A(n1981), .B(n1980), .Z(\A1[10] ) );
  XOR U20780 ( .A(n18667), .B(n18838), .Z(n1980) );
  XNOR U20781 ( .A(n18666), .B(n18664), .Z(n18838) );
  AND U20782 ( .A(n18839), .B(n18840), .Z(n18664) );
  NANDN U20783 ( .A(n18841), .B(n18842), .Z(n18840) );
  NANDN U20784 ( .A(n18843), .B(n18844), .Z(n18842) );
  OR U20785 ( .A(n18844), .B(n18), .Z(n18839) );
  AND U20786 ( .A(A[3]), .B(B[9]), .Z(n18666) );
  XNOR U20787 ( .A(n18656), .B(n18845), .Z(n18667) );
  XNOR U20788 ( .A(n18654), .B(n18657), .Z(n18845) );
  NANDN U20789 ( .A(n21), .B(A[2]), .Z(n18657) );
  NANDN U20790 ( .A(n18846), .B(n18847), .Z(n18654) );
  AND U20791 ( .A(A[0]), .B(B[11]), .Z(n18847) );
  XOR U20792 ( .A(n18659), .B(n18848), .Z(n18656) );
  NAND U20793 ( .A(A[0]), .B(B[12]), .Z(n18848) );
  NAND U20794 ( .A(B[11]), .B(A[1]), .Z(n18659) );
  NAND U20795 ( .A(n18849), .B(n18850), .Z(n1981) );
  NANDN U20796 ( .A(n2077), .B(n18851), .Z(n18850) );
  NANDN U20797 ( .A(n18852), .B(n2075), .Z(n18851) );
  NANDN U20798 ( .A(n26), .B(B[8]), .Z(n2077) );
  OR U20799 ( .A(n2075), .B(n19), .Z(n18849) );
  NAND U20800 ( .A(n18853), .B(n18854), .Z(n18852) );
  NANDN U20801 ( .A(n3944), .B(n18855), .Z(n18854) );
  NANDN U20802 ( .A(n20), .B(n18856), .Z(n18855) );
  NAND U20803 ( .A(B[8]), .B(A[2]), .Z(n3944) );
  NANDN U20804 ( .A(n18857), .B(n22), .Z(n18853) );
  NANDN U20805 ( .A(n5831), .B(n18858), .Z(n18856) );
  ANDN U20806 ( .B(A[0]), .A(n24), .Z(n18858) );
  NAND U20807 ( .A(B[8]), .B(A[1]), .Z(n5831) );
  XNOR U20808 ( .A(n18859), .B(n18860), .Z(n18857) );
  NANDN U20809 ( .A(n21), .B(A[0]), .Z(n18860) );
  XNOR U20810 ( .A(n18), .B(n18861), .Z(n2075) );
  XNOR U20811 ( .A(n18841), .B(n18844), .Z(n18861) );
  NANDN U20812 ( .A(n24), .B(A[2]), .Z(n18844) );
  NANDN U20813 ( .A(n18859), .B(n18862), .Z(n18841) );
  ANDN U20814 ( .B(A[0]), .A(n21), .Z(n18862) );
  NANDN U20815 ( .A(n24), .B(A[1]), .Z(n18859) );
  XOR U20816 ( .A(n18846), .B(n18863), .Z(n18843) );
  NAND U20817 ( .A(A[0]), .B(B[11]), .Z(n18863) );
  NANDN U20818 ( .A(n21), .B(A[1]), .Z(n18846) );
  XOR U20819 ( .A(n2001), .B(n2000), .Z(\A1[109] ) );
  XOR U20820 ( .A(n18837), .B(n18864), .Z(n2000) );
  XNOR U20821 ( .A(n18836), .B(n18834), .Z(n18864) );
  AND U20822 ( .A(n18865), .B(n18866), .Z(n18834) );
  NANDN U20823 ( .A(n18867), .B(n18868), .Z(n18866) );
  NANDN U20824 ( .A(n18869), .B(n18870), .Z(n18868) );
  AND U20825 ( .A(B[108]), .B(A[3]), .Z(n18836) );
  XNOR U20826 ( .A(n18826), .B(n18871), .Z(n18837) );
  XNOR U20827 ( .A(n18824), .B(n18827), .Z(n18871) );
  NAND U20828 ( .A(A[2]), .B(B[109]), .Z(n18827) );
  NANDN U20829 ( .A(n18872), .B(n18873), .Z(n18824) );
  AND U20830 ( .A(A[0]), .B(B[110]), .Z(n18873) );
  XOR U20831 ( .A(n18829), .B(n18874), .Z(n18826) );
  NAND U20832 ( .A(A[0]), .B(B[111]), .Z(n18874) );
  NAND U20833 ( .A(B[110]), .B(A[1]), .Z(n18829) );
  NAND U20834 ( .A(n18875), .B(n18876), .Z(n2001) );
  NANDN U20835 ( .A(n18877), .B(n18878), .Z(n18876) );
  OR U20836 ( .A(n18879), .B(n18880), .Z(n18878) );
  NAND U20837 ( .A(n18880), .B(n18879), .Z(n18875) );
  XOR U20838 ( .A(n2005), .B(n2004), .Z(\A1[108] ) );
  XOR U20839 ( .A(n18880), .B(n18881), .Z(n2004) );
  XNOR U20840 ( .A(n18879), .B(n18877), .Z(n18881) );
  AND U20841 ( .A(n18882), .B(n18883), .Z(n18877) );
  NANDN U20842 ( .A(n18884), .B(n18885), .Z(n18883) );
  NANDN U20843 ( .A(n18886), .B(n18887), .Z(n18885) );
  AND U20844 ( .A(B[107]), .B(A[3]), .Z(n18879) );
  XNOR U20845 ( .A(n18869), .B(n18888), .Z(n18880) );
  XNOR U20846 ( .A(n18867), .B(n18870), .Z(n18888) );
  NAND U20847 ( .A(A[2]), .B(B[108]), .Z(n18870) );
  NANDN U20848 ( .A(n18889), .B(n18890), .Z(n18867) );
  AND U20849 ( .A(A[0]), .B(B[109]), .Z(n18890) );
  XOR U20850 ( .A(n18872), .B(n18891), .Z(n18869) );
  NAND U20851 ( .A(A[0]), .B(B[110]), .Z(n18891) );
  NAND U20852 ( .A(B[109]), .B(A[1]), .Z(n18872) );
  NAND U20853 ( .A(n18892), .B(n18893), .Z(n2005) );
  NANDN U20854 ( .A(n18894), .B(n18895), .Z(n18893) );
  OR U20855 ( .A(n18896), .B(n18897), .Z(n18895) );
  NAND U20856 ( .A(n18897), .B(n18896), .Z(n18892) );
  XOR U20857 ( .A(n2007), .B(n2006), .Z(\A1[107] ) );
  XOR U20858 ( .A(n18897), .B(n18898), .Z(n2006) );
  XNOR U20859 ( .A(n18896), .B(n18894), .Z(n18898) );
  AND U20860 ( .A(n18899), .B(n18900), .Z(n18894) );
  NANDN U20861 ( .A(n18901), .B(n18902), .Z(n18900) );
  NANDN U20862 ( .A(n18903), .B(n18904), .Z(n18902) );
  AND U20863 ( .A(B[106]), .B(A[3]), .Z(n18896) );
  XNOR U20864 ( .A(n18886), .B(n18905), .Z(n18897) );
  XNOR U20865 ( .A(n18884), .B(n18887), .Z(n18905) );
  NAND U20866 ( .A(A[2]), .B(B[107]), .Z(n18887) );
  NANDN U20867 ( .A(n18906), .B(n18907), .Z(n18884) );
  AND U20868 ( .A(A[0]), .B(B[108]), .Z(n18907) );
  XOR U20869 ( .A(n18889), .B(n18908), .Z(n18886) );
  NAND U20870 ( .A(A[0]), .B(B[109]), .Z(n18908) );
  NAND U20871 ( .A(B[108]), .B(A[1]), .Z(n18889) );
  NAND U20872 ( .A(n18909), .B(n18910), .Z(n2007) );
  NANDN U20873 ( .A(n18911), .B(n18912), .Z(n18910) );
  OR U20874 ( .A(n18913), .B(n18914), .Z(n18912) );
  NAND U20875 ( .A(n18914), .B(n18913), .Z(n18909) );
  XOR U20876 ( .A(n2009), .B(n2008), .Z(\A1[106] ) );
  XOR U20877 ( .A(n18914), .B(n18915), .Z(n2008) );
  XNOR U20878 ( .A(n18913), .B(n18911), .Z(n18915) );
  AND U20879 ( .A(n18916), .B(n18917), .Z(n18911) );
  NANDN U20880 ( .A(n18918), .B(n18919), .Z(n18917) );
  NANDN U20881 ( .A(n18920), .B(n18921), .Z(n18919) );
  AND U20882 ( .A(B[105]), .B(A[3]), .Z(n18913) );
  XNOR U20883 ( .A(n18903), .B(n18922), .Z(n18914) );
  XNOR U20884 ( .A(n18901), .B(n18904), .Z(n18922) );
  NAND U20885 ( .A(A[2]), .B(B[106]), .Z(n18904) );
  NANDN U20886 ( .A(n18923), .B(n18924), .Z(n18901) );
  AND U20887 ( .A(A[0]), .B(B[107]), .Z(n18924) );
  XOR U20888 ( .A(n18906), .B(n18925), .Z(n18903) );
  NAND U20889 ( .A(A[0]), .B(B[108]), .Z(n18925) );
  NAND U20890 ( .A(B[107]), .B(A[1]), .Z(n18906) );
  NAND U20891 ( .A(n18926), .B(n18927), .Z(n2009) );
  NANDN U20892 ( .A(n18928), .B(n18929), .Z(n18927) );
  OR U20893 ( .A(n18930), .B(n18931), .Z(n18929) );
  NAND U20894 ( .A(n18931), .B(n18930), .Z(n18926) );
  XOR U20895 ( .A(n2011), .B(n2010), .Z(\A1[105] ) );
  XOR U20896 ( .A(n18931), .B(n18932), .Z(n2010) );
  XNOR U20897 ( .A(n18930), .B(n18928), .Z(n18932) );
  AND U20898 ( .A(n18933), .B(n18934), .Z(n18928) );
  NANDN U20899 ( .A(n18935), .B(n18936), .Z(n18934) );
  NANDN U20900 ( .A(n18937), .B(n18938), .Z(n18936) );
  AND U20901 ( .A(B[104]), .B(A[3]), .Z(n18930) );
  XNOR U20902 ( .A(n18920), .B(n18939), .Z(n18931) );
  XNOR U20903 ( .A(n18918), .B(n18921), .Z(n18939) );
  NAND U20904 ( .A(A[2]), .B(B[105]), .Z(n18921) );
  NANDN U20905 ( .A(n18940), .B(n18941), .Z(n18918) );
  AND U20906 ( .A(A[0]), .B(B[106]), .Z(n18941) );
  XOR U20907 ( .A(n18923), .B(n18942), .Z(n18920) );
  NAND U20908 ( .A(A[0]), .B(B[107]), .Z(n18942) );
  NAND U20909 ( .A(B[106]), .B(A[1]), .Z(n18923) );
  NAND U20910 ( .A(n18943), .B(n18944), .Z(n2011) );
  NANDN U20911 ( .A(n18945), .B(n18946), .Z(n18944) );
  OR U20912 ( .A(n18947), .B(n18948), .Z(n18946) );
  NAND U20913 ( .A(n18948), .B(n18947), .Z(n18943) );
  XOR U20914 ( .A(n2013), .B(n2012), .Z(\A1[104] ) );
  XOR U20915 ( .A(n18948), .B(n18949), .Z(n2012) );
  XNOR U20916 ( .A(n18947), .B(n18945), .Z(n18949) );
  AND U20917 ( .A(n18950), .B(n18951), .Z(n18945) );
  NANDN U20918 ( .A(n18952), .B(n18953), .Z(n18951) );
  NANDN U20919 ( .A(n18954), .B(n18955), .Z(n18953) );
  AND U20920 ( .A(B[103]), .B(A[3]), .Z(n18947) );
  XNOR U20921 ( .A(n18937), .B(n18956), .Z(n18948) );
  XNOR U20922 ( .A(n18935), .B(n18938), .Z(n18956) );
  NAND U20923 ( .A(A[2]), .B(B[104]), .Z(n18938) );
  NANDN U20924 ( .A(n18957), .B(n18958), .Z(n18935) );
  AND U20925 ( .A(A[0]), .B(B[105]), .Z(n18958) );
  XOR U20926 ( .A(n18940), .B(n18959), .Z(n18937) );
  NAND U20927 ( .A(A[0]), .B(B[106]), .Z(n18959) );
  NAND U20928 ( .A(B[105]), .B(A[1]), .Z(n18940) );
  NAND U20929 ( .A(n18960), .B(n18961), .Z(n2013) );
  NANDN U20930 ( .A(n18962), .B(n18963), .Z(n18961) );
  OR U20931 ( .A(n18964), .B(n18965), .Z(n18963) );
  NAND U20932 ( .A(n18965), .B(n18964), .Z(n18960) );
  XOR U20933 ( .A(n2015), .B(n2014), .Z(\A1[103] ) );
  XOR U20934 ( .A(n18965), .B(n18966), .Z(n2014) );
  XNOR U20935 ( .A(n18964), .B(n18962), .Z(n18966) );
  AND U20936 ( .A(n18967), .B(n18968), .Z(n18962) );
  NANDN U20937 ( .A(n18969), .B(n18970), .Z(n18968) );
  NANDN U20938 ( .A(n18971), .B(n18972), .Z(n18970) );
  AND U20939 ( .A(B[102]), .B(A[3]), .Z(n18964) );
  XNOR U20940 ( .A(n18954), .B(n18973), .Z(n18965) );
  XNOR U20941 ( .A(n18952), .B(n18955), .Z(n18973) );
  NAND U20942 ( .A(A[2]), .B(B[103]), .Z(n18955) );
  NANDN U20943 ( .A(n18974), .B(n18975), .Z(n18952) );
  AND U20944 ( .A(A[0]), .B(B[104]), .Z(n18975) );
  XOR U20945 ( .A(n18957), .B(n18976), .Z(n18954) );
  NAND U20946 ( .A(A[0]), .B(B[105]), .Z(n18976) );
  NAND U20947 ( .A(B[104]), .B(A[1]), .Z(n18957) );
  NAND U20948 ( .A(n18977), .B(n18978), .Z(n2015) );
  NANDN U20949 ( .A(n18979), .B(n18980), .Z(n18978) );
  OR U20950 ( .A(n18981), .B(n18982), .Z(n18980) );
  NAND U20951 ( .A(n18982), .B(n18981), .Z(n18977) );
  XOR U20952 ( .A(n2017), .B(n2016), .Z(\A1[102] ) );
  XOR U20953 ( .A(n18982), .B(n18983), .Z(n2016) );
  XNOR U20954 ( .A(n18981), .B(n18979), .Z(n18983) );
  AND U20955 ( .A(n18984), .B(n18985), .Z(n18979) );
  NANDN U20956 ( .A(n18986), .B(n18987), .Z(n18985) );
  NANDN U20957 ( .A(n18988), .B(n18989), .Z(n18987) );
  AND U20958 ( .A(B[101]), .B(A[3]), .Z(n18981) );
  XNOR U20959 ( .A(n18971), .B(n18990), .Z(n18982) );
  XNOR U20960 ( .A(n18969), .B(n18972), .Z(n18990) );
  NAND U20961 ( .A(A[2]), .B(B[102]), .Z(n18972) );
  NANDN U20962 ( .A(n18991), .B(n18992), .Z(n18969) );
  AND U20963 ( .A(A[0]), .B(B[103]), .Z(n18992) );
  XOR U20964 ( .A(n18974), .B(n18993), .Z(n18971) );
  NAND U20965 ( .A(A[0]), .B(B[104]), .Z(n18993) );
  NAND U20966 ( .A(B[103]), .B(A[1]), .Z(n18974) );
  NAND U20967 ( .A(n18994), .B(n18995), .Z(n2017) );
  NANDN U20968 ( .A(n18996), .B(n18997), .Z(n18995) );
  OR U20969 ( .A(n18998), .B(n18999), .Z(n18997) );
  NAND U20970 ( .A(n18999), .B(n18998), .Z(n18994) );
  XNOR U20972 ( .A(n2020), .B(n19000), .Z(\A1[1024] ) );
  NANDN U20973 ( .A(n26), .B(B[1023]), .Z(n19000) );
  NAND U20974 ( .A(n19001), .B(n19002), .Z(n2020) );
  NANDN U20975 ( .A(n19004), .B(n19005), .Z(n19003) );
  NANDN U20976 ( .A(n19005), .B(n19004), .Z(n19001) );
  XOR U20977 ( .A(n2022), .B(n2021), .Z(\A1[1023] ) );
  XNOR U20978 ( .A(n19006), .B(n19007), .Z(n2021) );
  XOR U20979 ( .A(n19004), .B(n19005), .Z(n19007) );
  NANDN U20980 ( .A(n3), .B(A[2]), .Z(n19005) );
  ANDN U20981 ( .B(B[1022]), .A(n26), .Z(n19004) );
  NAND U20982 ( .A(n19008), .B(n19009), .Z(n19006) );
  OR U20983 ( .A(n19010), .B(n19011), .Z(n19008) );
  NAND U20984 ( .A(n19012), .B(n19013), .Z(n2022) );
  NANDN U20985 ( .A(n19014), .B(n19015), .Z(n19013) );
  OR U20986 ( .A(n19016), .B(n19017), .Z(n19015) );
  NANDN U20987 ( .A(n2), .B(n19016), .Z(n19012) );
  XOR U20988 ( .A(n2024), .B(n2023), .Z(\A1[1022] ) );
  XNOR U20989 ( .A(n2), .B(n19018), .Z(n2023) );
  XNOR U20990 ( .A(n19016), .B(n19014), .Z(n19018) );
  AND U20991 ( .A(n19019), .B(n19020), .Z(n19014) );
  NANDN U20992 ( .A(n19021), .B(n19022), .Z(n19020) );
  NANDN U20993 ( .A(n19023), .B(n19024), .Z(n19022) );
  AND U20994 ( .A(B[1021]), .B(A[3]), .Z(n19016) );
  XOR U20995 ( .A(n19011), .B(n19025), .Z(n19017) );
  XNOR U20996 ( .A(n19009), .B(n19010), .Z(n19025) );
  NAND U20997 ( .A(A[2]), .B(B[1022]), .Z(n19010) );
  NAND U20998 ( .A(B[1023]), .B(n19026), .Z(n19009) );
  ANDN U20999 ( .B(A[0]), .A(n19027), .Z(n19026) );
  NANDN U21000 ( .A(n3), .B(A[1]), .Z(n19011) );
  NAND U21001 ( .A(n19028), .B(n19029), .Z(n2024) );
  NANDN U21002 ( .A(n19030), .B(n19031), .Z(n19029) );
  OR U21003 ( .A(n19032), .B(n19033), .Z(n19031) );
  NAND U21004 ( .A(n19033), .B(n19032), .Z(n19028) );
  XOR U21005 ( .A(n2026), .B(n2025), .Z(\A1[1021] ) );
  XOR U21006 ( .A(n19033), .B(n19034), .Z(n2025) );
  XNOR U21007 ( .A(n19032), .B(n19030), .Z(n19034) );
  AND U21008 ( .A(n19035), .B(n19036), .Z(n19030) );
  NANDN U21009 ( .A(n19037), .B(n19038), .Z(n19036) );
  NANDN U21010 ( .A(n19039), .B(n19040), .Z(n19038) );
  AND U21011 ( .A(B[1020]), .B(A[3]), .Z(n19032) );
  XNOR U21012 ( .A(n19023), .B(n19041), .Z(n19033) );
  XNOR U21013 ( .A(n19021), .B(n19024), .Z(n19041) );
  NAND U21014 ( .A(A[2]), .B(B[1021]), .Z(n19024) );
  NANDN U21015 ( .A(n19042), .B(n19043), .Z(n19021) );
  AND U21016 ( .A(A[0]), .B(B[1022]), .Z(n19043) );
  XOR U21017 ( .A(n19027), .B(n19044), .Z(n19023) );
  NANDN U21018 ( .A(n3), .B(A[0]), .Z(n19044) );
  NAND U21019 ( .A(B[1022]), .B(A[1]), .Z(n19027) );
  NAND U21020 ( .A(n19045), .B(n19046), .Z(n2026) );
  NANDN U21021 ( .A(n19047), .B(n19048), .Z(n19046) );
  OR U21022 ( .A(n19049), .B(n19050), .Z(n19048) );
  NAND U21023 ( .A(n19050), .B(n19049), .Z(n19045) );
  XOR U21024 ( .A(n2028), .B(n2027), .Z(\A1[1020] ) );
  XOR U21025 ( .A(n19050), .B(n19051), .Z(n2027) );
  XNOR U21026 ( .A(n19049), .B(n19047), .Z(n19051) );
  AND U21027 ( .A(n19052), .B(n19053), .Z(n19047) );
  NANDN U21028 ( .A(n19054), .B(n19055), .Z(n19053) );
  NANDN U21029 ( .A(n19056), .B(n19057), .Z(n19055) );
  AND U21030 ( .A(B[1019]), .B(A[3]), .Z(n19049) );
  XNOR U21031 ( .A(n19039), .B(n19058), .Z(n19050) );
  XNOR U21032 ( .A(n19037), .B(n19040), .Z(n19058) );
  NAND U21033 ( .A(A[2]), .B(B[1020]), .Z(n19040) );
  NANDN U21034 ( .A(n19059), .B(n19060), .Z(n19037) );
  AND U21035 ( .A(A[0]), .B(B[1021]), .Z(n19060) );
  XOR U21036 ( .A(n19042), .B(n19061), .Z(n19039) );
  NAND U21037 ( .A(A[0]), .B(B[1022]), .Z(n19061) );
  NAND U21038 ( .A(B[1021]), .B(A[1]), .Z(n19042) );
  NAND U21039 ( .A(n19062), .B(n19063), .Z(n2028) );
  NANDN U21040 ( .A(n19064), .B(n19065), .Z(n19063) );
  OR U21041 ( .A(n19066), .B(n19067), .Z(n19065) );
  NAND U21042 ( .A(n19067), .B(n19066), .Z(n19062) );
  XOR U21043 ( .A(n2019), .B(n2018), .Z(\A1[101] ) );
  XOR U21044 ( .A(n18999), .B(n19068), .Z(n2018) );
  XNOR U21045 ( .A(n18998), .B(n18996), .Z(n19068) );
  AND U21046 ( .A(n19069), .B(n19070), .Z(n18996) );
  NANDN U21047 ( .A(n19071), .B(n19072), .Z(n19070) );
  NANDN U21048 ( .A(n19073), .B(n19074), .Z(n19072) );
  AND U21049 ( .A(A[3]), .B(B[100]), .Z(n18998) );
  XNOR U21050 ( .A(n18988), .B(n19075), .Z(n18999) );
  XNOR U21051 ( .A(n18986), .B(n18989), .Z(n19075) );
  NAND U21052 ( .A(A[2]), .B(B[101]), .Z(n18989) );
  NANDN U21053 ( .A(n19076), .B(n19077), .Z(n18986) );
  AND U21054 ( .A(A[0]), .B(B[102]), .Z(n19077) );
  XOR U21055 ( .A(n18991), .B(n19078), .Z(n18988) );
  NAND U21056 ( .A(A[0]), .B(B[103]), .Z(n19078) );
  NAND U21057 ( .A(B[102]), .B(A[1]), .Z(n18991) );
  NAND U21058 ( .A(n19079), .B(n19080), .Z(n2019) );
  NANDN U21059 ( .A(n19081), .B(n19082), .Z(n19080) );
  OR U21060 ( .A(n19083), .B(n19084), .Z(n19082) );
  NAND U21061 ( .A(n19084), .B(n19083), .Z(n19079) );
  XOR U21062 ( .A(n2030), .B(n2029), .Z(\A1[1019] ) );
  XOR U21063 ( .A(n19067), .B(n19085), .Z(n2029) );
  XNOR U21064 ( .A(n19066), .B(n19064), .Z(n19085) );
  AND U21065 ( .A(n19086), .B(n19087), .Z(n19064) );
  NANDN U21066 ( .A(n19088), .B(n19089), .Z(n19087) );
  NANDN U21067 ( .A(n19090), .B(n19091), .Z(n19089) );
  AND U21068 ( .A(B[1018]), .B(A[3]), .Z(n19066) );
  XNOR U21069 ( .A(n19056), .B(n19092), .Z(n19067) );
  XNOR U21070 ( .A(n19054), .B(n19057), .Z(n19092) );
  NAND U21071 ( .A(A[2]), .B(B[1019]), .Z(n19057) );
  NANDN U21072 ( .A(n19093), .B(n19094), .Z(n19054) );
  AND U21073 ( .A(A[0]), .B(B[1020]), .Z(n19094) );
  XOR U21074 ( .A(n19059), .B(n19095), .Z(n19056) );
  NAND U21075 ( .A(A[0]), .B(B[1021]), .Z(n19095) );
  NAND U21076 ( .A(B[1020]), .B(A[1]), .Z(n19059) );
  NAND U21077 ( .A(n19096), .B(n19097), .Z(n2030) );
  NANDN U21078 ( .A(n19098), .B(n19099), .Z(n19097) );
  OR U21079 ( .A(n19100), .B(n19101), .Z(n19099) );
  NAND U21080 ( .A(n19101), .B(n19100), .Z(n19096) );
  XOR U21081 ( .A(n2034), .B(n2033), .Z(\A1[1018] ) );
  XOR U21082 ( .A(n19101), .B(n19102), .Z(n2033) );
  XNOR U21083 ( .A(n19100), .B(n19098), .Z(n19102) );
  AND U21084 ( .A(n19103), .B(n19104), .Z(n19098) );
  NANDN U21085 ( .A(n19105), .B(n19106), .Z(n19104) );
  NANDN U21086 ( .A(n19107), .B(n19108), .Z(n19106) );
  AND U21087 ( .A(B[1017]), .B(A[3]), .Z(n19100) );
  XNOR U21088 ( .A(n19090), .B(n19109), .Z(n19101) );
  XNOR U21089 ( .A(n19088), .B(n19091), .Z(n19109) );
  NAND U21090 ( .A(A[2]), .B(B[1018]), .Z(n19091) );
  NANDN U21091 ( .A(n19110), .B(n19111), .Z(n19088) );
  AND U21092 ( .A(A[0]), .B(B[1019]), .Z(n19111) );
  XOR U21093 ( .A(n19093), .B(n19112), .Z(n19090) );
  NAND U21094 ( .A(A[0]), .B(B[1020]), .Z(n19112) );
  NAND U21095 ( .A(B[1019]), .B(A[1]), .Z(n19093) );
  NAND U21096 ( .A(n19113), .B(n19114), .Z(n2034) );
  NANDN U21097 ( .A(n19115), .B(n19116), .Z(n19114) );
  OR U21098 ( .A(n19117), .B(n19118), .Z(n19116) );
  NAND U21099 ( .A(n19118), .B(n19117), .Z(n19113) );
  XOR U21100 ( .A(n2036), .B(n2035), .Z(\A1[1017] ) );
  XOR U21101 ( .A(n19118), .B(n19119), .Z(n2035) );
  XNOR U21102 ( .A(n19117), .B(n19115), .Z(n19119) );
  AND U21103 ( .A(n19120), .B(n19121), .Z(n19115) );
  NANDN U21104 ( .A(n19122), .B(n19123), .Z(n19121) );
  NANDN U21105 ( .A(n19124), .B(n19125), .Z(n19123) );
  AND U21106 ( .A(B[1016]), .B(A[3]), .Z(n19117) );
  XNOR U21107 ( .A(n19107), .B(n19126), .Z(n19118) );
  XNOR U21108 ( .A(n19105), .B(n19108), .Z(n19126) );
  NAND U21109 ( .A(A[2]), .B(B[1017]), .Z(n19108) );
  NANDN U21110 ( .A(n19127), .B(n19128), .Z(n19105) );
  AND U21111 ( .A(A[0]), .B(B[1018]), .Z(n19128) );
  XOR U21112 ( .A(n19110), .B(n19129), .Z(n19107) );
  NAND U21113 ( .A(A[0]), .B(B[1019]), .Z(n19129) );
  NAND U21114 ( .A(B[1018]), .B(A[1]), .Z(n19110) );
  NAND U21115 ( .A(n19130), .B(n19131), .Z(n2036) );
  NANDN U21116 ( .A(n19132), .B(n19133), .Z(n19131) );
  OR U21117 ( .A(n19134), .B(n19135), .Z(n19133) );
  NAND U21118 ( .A(n19135), .B(n19134), .Z(n19130) );
  XOR U21119 ( .A(n2038), .B(n2037), .Z(\A1[1016] ) );
  XOR U21120 ( .A(n19135), .B(n19136), .Z(n2037) );
  XNOR U21121 ( .A(n19134), .B(n19132), .Z(n19136) );
  AND U21122 ( .A(n19137), .B(n19138), .Z(n19132) );
  NANDN U21123 ( .A(n19139), .B(n19140), .Z(n19138) );
  NANDN U21124 ( .A(n19141), .B(n19142), .Z(n19140) );
  AND U21125 ( .A(B[1015]), .B(A[3]), .Z(n19134) );
  XNOR U21126 ( .A(n19124), .B(n19143), .Z(n19135) );
  XNOR U21127 ( .A(n19122), .B(n19125), .Z(n19143) );
  NAND U21128 ( .A(A[2]), .B(B[1016]), .Z(n19125) );
  NANDN U21129 ( .A(n19144), .B(n19145), .Z(n19122) );
  AND U21130 ( .A(A[0]), .B(B[1017]), .Z(n19145) );
  XOR U21131 ( .A(n19127), .B(n19146), .Z(n19124) );
  NAND U21132 ( .A(A[0]), .B(B[1018]), .Z(n19146) );
  NAND U21133 ( .A(B[1017]), .B(A[1]), .Z(n19127) );
  NAND U21134 ( .A(n19147), .B(n19148), .Z(n2038) );
  NANDN U21135 ( .A(n19149), .B(n19150), .Z(n19148) );
  OR U21136 ( .A(n19151), .B(n19152), .Z(n19150) );
  NAND U21137 ( .A(n19152), .B(n19151), .Z(n19147) );
  XOR U21138 ( .A(n2040), .B(n2039), .Z(\A1[1015] ) );
  XOR U21139 ( .A(n19152), .B(n19153), .Z(n2039) );
  XNOR U21140 ( .A(n19151), .B(n19149), .Z(n19153) );
  AND U21141 ( .A(n19154), .B(n19155), .Z(n19149) );
  NANDN U21142 ( .A(n19156), .B(n19157), .Z(n19155) );
  NANDN U21143 ( .A(n19158), .B(n19159), .Z(n19157) );
  AND U21144 ( .A(B[1014]), .B(A[3]), .Z(n19151) );
  XNOR U21145 ( .A(n19141), .B(n19160), .Z(n19152) );
  XNOR U21146 ( .A(n19139), .B(n19142), .Z(n19160) );
  NAND U21147 ( .A(A[2]), .B(B[1015]), .Z(n19142) );
  NANDN U21148 ( .A(n19161), .B(n19162), .Z(n19139) );
  AND U21149 ( .A(A[0]), .B(B[1016]), .Z(n19162) );
  XOR U21150 ( .A(n19144), .B(n19163), .Z(n19141) );
  NAND U21151 ( .A(A[0]), .B(B[1017]), .Z(n19163) );
  NAND U21152 ( .A(B[1016]), .B(A[1]), .Z(n19144) );
  NAND U21153 ( .A(n19164), .B(n19165), .Z(n2040) );
  NANDN U21154 ( .A(n19166), .B(n19167), .Z(n19165) );
  OR U21155 ( .A(n19168), .B(n19169), .Z(n19167) );
  NAND U21156 ( .A(n19169), .B(n19168), .Z(n19164) );
  XOR U21157 ( .A(n2042), .B(n2041), .Z(\A1[1014] ) );
  XOR U21158 ( .A(n19169), .B(n19170), .Z(n2041) );
  XNOR U21159 ( .A(n19168), .B(n19166), .Z(n19170) );
  AND U21160 ( .A(n19171), .B(n19172), .Z(n19166) );
  NANDN U21161 ( .A(n19173), .B(n19174), .Z(n19172) );
  NANDN U21162 ( .A(n19175), .B(n19176), .Z(n19174) );
  AND U21163 ( .A(B[1013]), .B(A[3]), .Z(n19168) );
  XNOR U21164 ( .A(n19158), .B(n19177), .Z(n19169) );
  XNOR U21165 ( .A(n19156), .B(n19159), .Z(n19177) );
  NAND U21166 ( .A(A[2]), .B(B[1014]), .Z(n19159) );
  NANDN U21167 ( .A(n19178), .B(n19179), .Z(n19156) );
  AND U21168 ( .A(A[0]), .B(B[1015]), .Z(n19179) );
  XOR U21169 ( .A(n19161), .B(n19180), .Z(n19158) );
  NAND U21170 ( .A(A[0]), .B(B[1016]), .Z(n19180) );
  NAND U21171 ( .A(B[1015]), .B(A[1]), .Z(n19161) );
  NAND U21172 ( .A(n19181), .B(n19182), .Z(n2042) );
  NANDN U21173 ( .A(n19183), .B(n19184), .Z(n19182) );
  OR U21174 ( .A(n19185), .B(n19186), .Z(n19184) );
  NAND U21175 ( .A(n19186), .B(n19185), .Z(n19181) );
  XOR U21176 ( .A(n2044), .B(n2043), .Z(\A1[1013] ) );
  XOR U21177 ( .A(n19186), .B(n19187), .Z(n2043) );
  XNOR U21178 ( .A(n19185), .B(n19183), .Z(n19187) );
  AND U21179 ( .A(n19188), .B(n19189), .Z(n19183) );
  NANDN U21180 ( .A(n19190), .B(n19191), .Z(n19189) );
  NANDN U21181 ( .A(n19192), .B(n19193), .Z(n19191) );
  AND U21182 ( .A(B[1012]), .B(A[3]), .Z(n19185) );
  XNOR U21183 ( .A(n19175), .B(n19194), .Z(n19186) );
  XNOR U21184 ( .A(n19173), .B(n19176), .Z(n19194) );
  NAND U21185 ( .A(A[2]), .B(B[1013]), .Z(n19176) );
  NANDN U21186 ( .A(n19195), .B(n19196), .Z(n19173) );
  AND U21187 ( .A(A[0]), .B(B[1014]), .Z(n19196) );
  XOR U21188 ( .A(n19178), .B(n19197), .Z(n19175) );
  NAND U21189 ( .A(A[0]), .B(B[1015]), .Z(n19197) );
  NAND U21190 ( .A(B[1014]), .B(A[1]), .Z(n19178) );
  NAND U21191 ( .A(n19198), .B(n19199), .Z(n2044) );
  NANDN U21192 ( .A(n19200), .B(n19201), .Z(n19199) );
  OR U21193 ( .A(n19202), .B(n19203), .Z(n19201) );
  NAND U21194 ( .A(n19203), .B(n19202), .Z(n19198) );
  XOR U21195 ( .A(n2046), .B(n2045), .Z(\A1[1012] ) );
  XOR U21196 ( .A(n19203), .B(n19204), .Z(n2045) );
  XNOR U21197 ( .A(n19202), .B(n19200), .Z(n19204) );
  AND U21198 ( .A(n19205), .B(n19206), .Z(n19200) );
  NANDN U21199 ( .A(n19207), .B(n19208), .Z(n19206) );
  NANDN U21200 ( .A(n19209), .B(n19210), .Z(n19208) );
  AND U21201 ( .A(B[1011]), .B(A[3]), .Z(n19202) );
  XNOR U21202 ( .A(n19192), .B(n19211), .Z(n19203) );
  XNOR U21203 ( .A(n19190), .B(n19193), .Z(n19211) );
  NAND U21204 ( .A(A[2]), .B(B[1012]), .Z(n19193) );
  NANDN U21205 ( .A(n19212), .B(n19213), .Z(n19190) );
  AND U21206 ( .A(A[0]), .B(B[1013]), .Z(n19213) );
  XOR U21207 ( .A(n19195), .B(n19214), .Z(n19192) );
  NAND U21208 ( .A(A[0]), .B(B[1014]), .Z(n19214) );
  NAND U21209 ( .A(B[1013]), .B(A[1]), .Z(n19195) );
  NAND U21210 ( .A(n19215), .B(n19216), .Z(n2046) );
  NANDN U21211 ( .A(n19217), .B(n19218), .Z(n19216) );
  OR U21212 ( .A(n19219), .B(n19220), .Z(n19218) );
  NAND U21213 ( .A(n19220), .B(n19219), .Z(n19215) );
  XOR U21214 ( .A(n2048), .B(n2047), .Z(\A1[1011] ) );
  XOR U21215 ( .A(n19220), .B(n19221), .Z(n2047) );
  XNOR U21216 ( .A(n19219), .B(n19217), .Z(n19221) );
  AND U21217 ( .A(n19222), .B(n19223), .Z(n19217) );
  NANDN U21218 ( .A(n19224), .B(n19225), .Z(n19223) );
  NANDN U21219 ( .A(n19226), .B(n19227), .Z(n19225) );
  AND U21220 ( .A(B[1010]), .B(A[3]), .Z(n19219) );
  XNOR U21221 ( .A(n19209), .B(n19228), .Z(n19220) );
  XNOR U21222 ( .A(n19207), .B(n19210), .Z(n19228) );
  NAND U21223 ( .A(A[2]), .B(B[1011]), .Z(n19210) );
  NANDN U21224 ( .A(n19229), .B(n19230), .Z(n19207) );
  AND U21225 ( .A(A[0]), .B(B[1012]), .Z(n19230) );
  XOR U21226 ( .A(n19212), .B(n19231), .Z(n19209) );
  NAND U21227 ( .A(A[0]), .B(B[1013]), .Z(n19231) );
  NAND U21228 ( .A(B[1012]), .B(A[1]), .Z(n19212) );
  NAND U21229 ( .A(n19232), .B(n19233), .Z(n2048) );
  NANDN U21230 ( .A(n19234), .B(n19235), .Z(n19233) );
  OR U21231 ( .A(n19236), .B(n19237), .Z(n19235) );
  NAND U21232 ( .A(n19237), .B(n19236), .Z(n19232) );
  XOR U21233 ( .A(n2050), .B(n2049), .Z(\A1[1010] ) );
  XOR U21234 ( .A(n19237), .B(n19238), .Z(n2049) );
  XNOR U21235 ( .A(n19236), .B(n19234), .Z(n19238) );
  AND U21236 ( .A(n19239), .B(n19240), .Z(n19234) );
  NANDN U21237 ( .A(n19241), .B(n19242), .Z(n19240) );
  NANDN U21238 ( .A(n19243), .B(n19244), .Z(n19242) );
  AND U21239 ( .A(B[1009]), .B(A[3]), .Z(n19236) );
  XNOR U21240 ( .A(n19226), .B(n19245), .Z(n19237) );
  XNOR U21241 ( .A(n19224), .B(n19227), .Z(n19245) );
  NAND U21242 ( .A(A[2]), .B(B[1010]), .Z(n19227) );
  NANDN U21243 ( .A(n19246), .B(n19247), .Z(n19224) );
  AND U21244 ( .A(A[0]), .B(B[1011]), .Z(n19247) );
  XOR U21245 ( .A(n19229), .B(n19248), .Z(n19226) );
  NAND U21246 ( .A(A[0]), .B(B[1012]), .Z(n19248) );
  NAND U21247 ( .A(B[1011]), .B(A[1]), .Z(n19229) );
  NAND U21248 ( .A(n19249), .B(n19250), .Z(n2050) );
  NANDN U21249 ( .A(n19251), .B(n19252), .Z(n19250) );
  OR U21250 ( .A(n19253), .B(n19254), .Z(n19252) );
  NAND U21251 ( .A(n19254), .B(n19253), .Z(n19249) );
  XOR U21252 ( .A(n2032), .B(n2031), .Z(\A1[100] ) );
  XOR U21253 ( .A(n19084), .B(n19255), .Z(n2031) );
  XNOR U21254 ( .A(n19083), .B(n19081), .Z(n19255) );
  AND U21255 ( .A(n19256), .B(n19257), .Z(n19081) );
  NANDN U21256 ( .A(n19258), .B(n19259), .Z(n19257) );
  NANDN U21257 ( .A(n19260), .B(n19261), .Z(n19259) );
  OR U21258 ( .A(n19261), .B(n11), .Z(n19256) );
  AND U21259 ( .A(A[3]), .B(B[99]), .Z(n19083) );
  XNOR U21260 ( .A(n19073), .B(n19262), .Z(n19084) );
  XNOR U21261 ( .A(n19071), .B(n19074), .Z(n19262) );
  NANDN U21262 ( .A(n14), .B(A[2]), .Z(n19074) );
  NANDN U21263 ( .A(n19263), .B(n19264), .Z(n19071) );
  AND U21264 ( .A(A[0]), .B(B[101]), .Z(n19264) );
  XOR U21265 ( .A(n19076), .B(n19265), .Z(n19073) );
  NAND U21266 ( .A(A[0]), .B(B[102]), .Z(n19265) );
  NAND U21267 ( .A(B[101]), .B(A[1]), .Z(n19076) );
  NAND U21268 ( .A(n19266), .B(n19267), .Z(n2032) );
  NANDN U21269 ( .A(n2086), .B(n19268), .Z(n19267) );
  NANDN U21270 ( .A(n19269), .B(n2084), .Z(n19268) );
  NANDN U21271 ( .A(n26), .B(B[98]), .Z(n2086) );
  OR U21272 ( .A(n2084), .B(n12), .Z(n19266) );
  NAND U21273 ( .A(n19270), .B(n19271), .Z(n19269) );
  NANDN U21274 ( .A(n2262), .B(n19272), .Z(n19271) );
  NANDN U21275 ( .A(n13), .B(n19273), .Z(n19272) );
  NAND U21276 ( .A(B[98]), .B(A[2]), .Z(n2262) );
  NANDN U21277 ( .A(n19274), .B(n15), .Z(n19270) );
  NANDN U21278 ( .A(n2449), .B(n19275), .Z(n19273) );
  ANDN U21279 ( .B(A[0]), .A(n17), .Z(n19275) );
  NAND U21280 ( .A(B[98]), .B(A[1]), .Z(n2449) );
  XNOR U21281 ( .A(n19276), .B(n19277), .Z(n19274) );
  NANDN U21282 ( .A(n14), .B(A[0]), .Z(n19277) );
  XNOR U21283 ( .A(n11), .B(n19278), .Z(n2084) );
  XNOR U21284 ( .A(n19258), .B(n19261), .Z(n19278) );
  NANDN U21285 ( .A(n17), .B(A[2]), .Z(n19261) );
  NANDN U21286 ( .A(n19276), .B(n19279), .Z(n19258) );
  ANDN U21287 ( .B(A[0]), .A(n14), .Z(n19279) );
  NANDN U21288 ( .A(n17), .B(A[1]), .Z(n19276) );
  XOR U21289 ( .A(n19263), .B(n19280), .Z(n19260) );
  NAND U21290 ( .A(A[0]), .B(B[101]), .Z(n19280) );
  NANDN U21291 ( .A(n14), .B(A[1]), .Z(n19263) );
  XOR U21292 ( .A(n2052), .B(n2051), .Z(\A1[1009] ) );
  XOR U21293 ( .A(n19254), .B(n19281), .Z(n2051) );
  XNOR U21294 ( .A(n19253), .B(n19251), .Z(n19281) );
  AND U21295 ( .A(n19282), .B(n19283), .Z(n19251) );
  NANDN U21296 ( .A(n19284), .B(n19285), .Z(n19283) );
  NANDN U21297 ( .A(n19286), .B(n19287), .Z(n19285) );
  AND U21298 ( .A(B[1008]), .B(A[3]), .Z(n19253) );
  XNOR U21299 ( .A(n19243), .B(n19288), .Z(n19254) );
  XNOR U21300 ( .A(n19241), .B(n19244), .Z(n19288) );
  NAND U21301 ( .A(A[2]), .B(B[1009]), .Z(n19244) );
  NANDN U21302 ( .A(n19289), .B(n19290), .Z(n19241) );
  AND U21303 ( .A(A[0]), .B(B[1010]), .Z(n19290) );
  XOR U21304 ( .A(n19246), .B(n19291), .Z(n19243) );
  NAND U21305 ( .A(A[0]), .B(B[1011]), .Z(n19291) );
  NAND U21306 ( .A(B[1010]), .B(A[1]), .Z(n19246) );
  NAND U21307 ( .A(n19292), .B(n19293), .Z(n2052) );
  NANDN U21308 ( .A(n19294), .B(n19295), .Z(n19293) );
  OR U21309 ( .A(n19296), .B(n19297), .Z(n19295) );
  NAND U21310 ( .A(n19297), .B(n19296), .Z(n19292) );
  XOR U21311 ( .A(n2056), .B(n2055), .Z(\A1[1008] ) );
  XOR U21312 ( .A(n19297), .B(n19298), .Z(n2055) );
  XNOR U21313 ( .A(n19296), .B(n19294), .Z(n19298) );
  AND U21314 ( .A(n19299), .B(n19300), .Z(n19294) );
  NANDN U21315 ( .A(n19301), .B(n19302), .Z(n19300) );
  NANDN U21316 ( .A(n19303), .B(n19304), .Z(n19302) );
  AND U21317 ( .A(B[1007]), .B(A[3]), .Z(n19296) );
  XNOR U21318 ( .A(n19286), .B(n19305), .Z(n19297) );
  XNOR U21319 ( .A(n19284), .B(n19287), .Z(n19305) );
  NAND U21320 ( .A(A[2]), .B(B[1008]), .Z(n19287) );
  NANDN U21321 ( .A(n19306), .B(n19307), .Z(n19284) );
  AND U21322 ( .A(A[0]), .B(B[1009]), .Z(n19307) );
  XOR U21323 ( .A(n19289), .B(n19308), .Z(n19286) );
  NAND U21324 ( .A(A[0]), .B(B[1010]), .Z(n19308) );
  NAND U21325 ( .A(B[1009]), .B(A[1]), .Z(n19289) );
  NAND U21326 ( .A(n19309), .B(n19310), .Z(n2056) );
  NANDN U21327 ( .A(n19311), .B(n19312), .Z(n19310) );
  OR U21328 ( .A(n19313), .B(n19314), .Z(n19312) );
  NAND U21329 ( .A(n19314), .B(n19313), .Z(n19309) );
  XOR U21330 ( .A(n2058), .B(n2057), .Z(\A1[1007] ) );
  XOR U21331 ( .A(n19314), .B(n19315), .Z(n2057) );
  XNOR U21332 ( .A(n19313), .B(n19311), .Z(n19315) );
  AND U21333 ( .A(n19316), .B(n19317), .Z(n19311) );
  NANDN U21334 ( .A(n19318), .B(n19319), .Z(n19317) );
  NANDN U21335 ( .A(n19320), .B(n19321), .Z(n19319) );
  AND U21336 ( .A(B[1006]), .B(A[3]), .Z(n19313) );
  XNOR U21337 ( .A(n19303), .B(n19322), .Z(n19314) );
  XNOR U21338 ( .A(n19301), .B(n19304), .Z(n19322) );
  NAND U21339 ( .A(A[2]), .B(B[1007]), .Z(n19304) );
  NANDN U21340 ( .A(n19323), .B(n19324), .Z(n19301) );
  AND U21341 ( .A(A[0]), .B(B[1008]), .Z(n19324) );
  XOR U21342 ( .A(n19306), .B(n19325), .Z(n19303) );
  NAND U21343 ( .A(A[0]), .B(B[1009]), .Z(n19325) );
  NAND U21344 ( .A(B[1008]), .B(A[1]), .Z(n19306) );
  NAND U21345 ( .A(n19326), .B(n19327), .Z(n2058) );
  NANDN U21346 ( .A(n19328), .B(n19329), .Z(n19327) );
  OR U21347 ( .A(n19330), .B(n19331), .Z(n19329) );
  NAND U21348 ( .A(n19331), .B(n19330), .Z(n19326) );
  XOR U21349 ( .A(n2060), .B(n2059), .Z(\A1[1006] ) );
  XOR U21350 ( .A(n19331), .B(n19332), .Z(n2059) );
  XNOR U21351 ( .A(n19330), .B(n19328), .Z(n19332) );
  AND U21352 ( .A(n19333), .B(n19334), .Z(n19328) );
  NANDN U21353 ( .A(n19335), .B(n19336), .Z(n19334) );
  NANDN U21354 ( .A(n19337), .B(n19338), .Z(n19336) );
  AND U21355 ( .A(B[1005]), .B(A[3]), .Z(n19330) );
  XNOR U21356 ( .A(n19320), .B(n19339), .Z(n19331) );
  XNOR U21357 ( .A(n19318), .B(n19321), .Z(n19339) );
  NAND U21358 ( .A(A[2]), .B(B[1006]), .Z(n19321) );
  NANDN U21359 ( .A(n19340), .B(n19341), .Z(n19318) );
  AND U21360 ( .A(A[0]), .B(B[1007]), .Z(n19341) );
  XOR U21361 ( .A(n19323), .B(n19342), .Z(n19320) );
  NAND U21362 ( .A(A[0]), .B(B[1008]), .Z(n19342) );
  NAND U21363 ( .A(B[1007]), .B(A[1]), .Z(n19323) );
  NAND U21364 ( .A(n19343), .B(n19344), .Z(n2060) );
  NANDN U21365 ( .A(n19345), .B(n19346), .Z(n19344) );
  OR U21366 ( .A(n19347), .B(n19348), .Z(n19346) );
  NAND U21367 ( .A(n19348), .B(n19347), .Z(n19343) );
  XOR U21368 ( .A(n2062), .B(n2061), .Z(\A1[1005] ) );
  XOR U21369 ( .A(n19348), .B(n19349), .Z(n2061) );
  XNOR U21370 ( .A(n19347), .B(n19345), .Z(n19349) );
  AND U21371 ( .A(n19350), .B(n19351), .Z(n19345) );
  NANDN U21372 ( .A(n19352), .B(n19353), .Z(n19351) );
  NANDN U21373 ( .A(n19354), .B(n19355), .Z(n19353) );
  AND U21374 ( .A(B[1004]), .B(A[3]), .Z(n19347) );
  XNOR U21375 ( .A(n19337), .B(n19356), .Z(n19348) );
  XNOR U21376 ( .A(n19335), .B(n19338), .Z(n19356) );
  NAND U21377 ( .A(A[2]), .B(B[1005]), .Z(n19338) );
  NANDN U21378 ( .A(n19357), .B(n19358), .Z(n19335) );
  AND U21379 ( .A(A[0]), .B(B[1006]), .Z(n19358) );
  XOR U21380 ( .A(n19340), .B(n19359), .Z(n19337) );
  NAND U21381 ( .A(A[0]), .B(B[1007]), .Z(n19359) );
  NAND U21382 ( .A(B[1006]), .B(A[1]), .Z(n19340) );
  NAND U21383 ( .A(n19360), .B(n19361), .Z(n2062) );
  NANDN U21384 ( .A(n19362), .B(n19363), .Z(n19361) );
  OR U21385 ( .A(n19364), .B(n19365), .Z(n19363) );
  NAND U21386 ( .A(n19365), .B(n19364), .Z(n19360) );
  XOR U21387 ( .A(n2064), .B(n2063), .Z(\A1[1004] ) );
  XOR U21388 ( .A(n19365), .B(n19366), .Z(n2063) );
  XNOR U21389 ( .A(n19364), .B(n19362), .Z(n19366) );
  AND U21390 ( .A(n19367), .B(n19368), .Z(n19362) );
  NANDN U21391 ( .A(n19369), .B(n19370), .Z(n19368) );
  NANDN U21392 ( .A(n19371), .B(n19372), .Z(n19370) );
  AND U21393 ( .A(B[1003]), .B(A[3]), .Z(n19364) );
  XNOR U21394 ( .A(n19354), .B(n19373), .Z(n19365) );
  XNOR U21395 ( .A(n19352), .B(n19355), .Z(n19373) );
  NAND U21396 ( .A(A[2]), .B(B[1004]), .Z(n19355) );
  NANDN U21397 ( .A(n19374), .B(n19375), .Z(n19352) );
  AND U21398 ( .A(A[0]), .B(B[1005]), .Z(n19375) );
  XOR U21399 ( .A(n19357), .B(n19376), .Z(n19354) );
  NAND U21400 ( .A(A[0]), .B(B[1006]), .Z(n19376) );
  NAND U21401 ( .A(B[1005]), .B(A[1]), .Z(n19357) );
  NAND U21402 ( .A(n19377), .B(n19378), .Z(n2064) );
  NANDN U21403 ( .A(n19379), .B(n19380), .Z(n19378) );
  OR U21404 ( .A(n19381), .B(n19382), .Z(n19380) );
  NAND U21405 ( .A(n19382), .B(n19381), .Z(n19377) );
  XOR U21406 ( .A(n2066), .B(n2065), .Z(\A1[1003] ) );
  XOR U21407 ( .A(n19382), .B(n19383), .Z(n2065) );
  XNOR U21408 ( .A(n19381), .B(n19379), .Z(n19383) );
  AND U21409 ( .A(n19384), .B(n19385), .Z(n19379) );
  NANDN U21410 ( .A(n19386), .B(n19387), .Z(n19385) );
  NANDN U21411 ( .A(n19388), .B(n19389), .Z(n19387) );
  AND U21412 ( .A(B[1002]), .B(A[3]), .Z(n19381) );
  XNOR U21413 ( .A(n19371), .B(n19390), .Z(n19382) );
  XNOR U21414 ( .A(n19369), .B(n19372), .Z(n19390) );
  NAND U21415 ( .A(A[2]), .B(B[1003]), .Z(n19372) );
  NANDN U21416 ( .A(n19391), .B(n19392), .Z(n19369) );
  AND U21417 ( .A(A[0]), .B(B[1004]), .Z(n19392) );
  XOR U21418 ( .A(n19374), .B(n19393), .Z(n19371) );
  NAND U21419 ( .A(A[0]), .B(B[1005]), .Z(n19393) );
  NAND U21420 ( .A(B[1004]), .B(A[1]), .Z(n19374) );
  NAND U21421 ( .A(n19394), .B(n19395), .Z(n2066) );
  NANDN U21422 ( .A(n19396), .B(n19397), .Z(n19395) );
  OR U21423 ( .A(n19398), .B(n19399), .Z(n19397) );
  NAND U21424 ( .A(n19399), .B(n19398), .Z(n19394) );
  XOR U21425 ( .A(n2068), .B(n2067), .Z(\A1[1002] ) );
  XOR U21426 ( .A(n19399), .B(n19400), .Z(n2067) );
  XNOR U21427 ( .A(n19398), .B(n19396), .Z(n19400) );
  AND U21428 ( .A(n19401), .B(n19402), .Z(n19396) );
  NANDN U21429 ( .A(n19403), .B(n19404), .Z(n19402) );
  NANDN U21430 ( .A(n19405), .B(n19406), .Z(n19404) );
  AND U21431 ( .A(B[1001]), .B(A[3]), .Z(n19398) );
  XNOR U21432 ( .A(n19388), .B(n19407), .Z(n19399) );
  XNOR U21433 ( .A(n19386), .B(n19389), .Z(n19407) );
  NAND U21434 ( .A(A[2]), .B(B[1002]), .Z(n19389) );
  NANDN U21435 ( .A(n19408), .B(n19409), .Z(n19386) );
  AND U21436 ( .A(A[0]), .B(B[1003]), .Z(n19409) );
  XOR U21437 ( .A(n19391), .B(n19410), .Z(n19388) );
  NAND U21438 ( .A(A[0]), .B(B[1004]), .Z(n19410) );
  NAND U21439 ( .A(B[1003]), .B(A[1]), .Z(n19391) );
  NAND U21440 ( .A(n19411), .B(n19412), .Z(n2068) );
  NANDN U21441 ( .A(n19413), .B(n19414), .Z(n19412) );
  OR U21442 ( .A(n19415), .B(n19416), .Z(n19414) );
  NAND U21443 ( .A(n19416), .B(n19415), .Z(n19411) );
  XOR U21444 ( .A(n2070), .B(n2069), .Z(\A1[1001] ) );
  XOR U21445 ( .A(n19416), .B(n19417), .Z(n2069) );
  XNOR U21446 ( .A(n19415), .B(n19413), .Z(n19417) );
  AND U21447 ( .A(n19418), .B(n19419), .Z(n19413) );
  NANDN U21448 ( .A(n19420), .B(n19421), .Z(n19419) );
  NANDN U21449 ( .A(n19422), .B(n19423), .Z(n19421) );
  AND U21450 ( .A(A[3]), .B(B[1000]), .Z(n19415) );
  XNOR U21451 ( .A(n19405), .B(n19424), .Z(n19416) );
  XNOR U21452 ( .A(n19403), .B(n19406), .Z(n19424) );
  NAND U21453 ( .A(A[2]), .B(B[1001]), .Z(n19406) );
  NANDN U21454 ( .A(n19425), .B(n19426), .Z(n19403) );
  AND U21455 ( .A(A[0]), .B(B[1002]), .Z(n19426) );
  XOR U21456 ( .A(n19408), .B(n19427), .Z(n19405) );
  NAND U21457 ( .A(A[0]), .B(B[1003]), .Z(n19427) );
  NAND U21458 ( .A(B[1002]), .B(A[1]), .Z(n19408) );
  NAND U21459 ( .A(n19428), .B(n19429), .Z(n2070) );
  NANDN U21460 ( .A(n19430), .B(n19431), .Z(n19429) );
  OR U21461 ( .A(n19432), .B(n19433), .Z(n19431) );
  NAND U21462 ( .A(n19433), .B(n19432), .Z(n19428) );
  XOR U21463 ( .A(n2072), .B(n2071), .Z(\A1[1000] ) );
  XOR U21464 ( .A(n19433), .B(n19434), .Z(n2071) );
  XNOR U21465 ( .A(n19432), .B(n19430), .Z(n19434) );
  AND U21466 ( .A(n19435), .B(n19436), .Z(n19430) );
  NANDN U21467 ( .A(n19437), .B(n19438), .Z(n19436) );
  NANDN U21468 ( .A(n19439), .B(n19440), .Z(n19438) );
  OR U21469 ( .A(n19440), .B(n4), .Z(n19435) );
  AND U21470 ( .A(A[3]), .B(B[999]), .Z(n19432) );
  XNOR U21471 ( .A(n19422), .B(n19441), .Z(n19433) );
  XNOR U21472 ( .A(n19420), .B(n19423), .Z(n19441) );
  NANDN U21473 ( .A(n7), .B(A[2]), .Z(n19423) );
  NANDN U21474 ( .A(n19442), .B(n19443), .Z(n19420) );
  AND U21475 ( .A(A[0]), .B(B[1001]), .Z(n19443) );
  XOR U21476 ( .A(n19425), .B(n19444), .Z(n19422) );
  NAND U21477 ( .A(A[0]), .B(B[1002]), .Z(n19444) );
  NAND U21478 ( .A(B[1001]), .B(A[1]), .Z(n19425) );
  NAND U21479 ( .A(n19445), .B(n19446), .Z(n2072) );
  NANDN U21480 ( .A(n2095), .B(n19447), .Z(n19446) );
  NANDN U21481 ( .A(n19448), .B(n2093), .Z(n19447) );
  NANDN U21482 ( .A(n26), .B(B[998]), .Z(n2095) );
  OR U21483 ( .A(n2093), .B(n5), .Z(n19445) );
  NAND U21484 ( .A(n19449), .B(n19450), .Z(n19448) );
  NANDN U21485 ( .A(n2110), .B(n19451), .Z(n19450) );
  NANDN U21486 ( .A(n6), .B(n19452), .Z(n19451) );
  NAND U21487 ( .A(B[998]), .B(A[2]), .Z(n2110) );
  NANDN U21488 ( .A(n19453), .B(n8), .Z(n19449) );
  NANDN U21489 ( .A(n2127), .B(n19454), .Z(n19452) );
  ANDN U21490 ( .B(A[0]), .A(n10), .Z(n19454) );
  NAND U21491 ( .A(B[998]), .B(A[1]), .Z(n2127) );
  XNOR U21492 ( .A(n19455), .B(n19456), .Z(n19453) );
  NANDN U21493 ( .A(n7), .B(A[0]), .Z(n19456) );
  XNOR U21494 ( .A(n4), .B(n19457), .Z(n2093) );
  XNOR U21495 ( .A(n19437), .B(n19440), .Z(n19457) );
  NANDN U21496 ( .A(n10), .B(A[2]), .Z(n19440) );
  NANDN U21497 ( .A(n19455), .B(n19458), .Z(n19437) );
  ANDN U21498 ( .B(A[0]), .A(n7), .Z(n19458) );
  NANDN U21499 ( .A(n10), .B(A[1]), .Z(n19455) );
  XOR U21500 ( .A(n19442), .B(n19459), .Z(n19439) );
  NAND U21501 ( .A(A[0]), .B(B[1001]), .Z(n19459) );
  NANDN U21502 ( .A(n7), .B(A[1]), .Z(n19442) );
  XOR U21503 ( .A(n17150), .B(n19460), .Z(\A1[0] ) );
  XNOR U21504 ( .A(n17147), .B(n17149), .Z(n19460) );
  ANDN U21505 ( .B(n29), .A(n28), .Z(n17149) );
  NAND U21506 ( .A(B[0]), .B(A[1]), .Z(n28) );
  AND U21507 ( .A(A[0]), .B(B[1]), .Z(n29) );
  NAND U21508 ( .A(B[0]), .B(A[2]), .Z(n17147) );
  XOR U21509 ( .A(n17152), .B(n19461), .Z(n17150) );
  NAND U21510 ( .A(A[0]), .B(B[2]), .Z(n19461) );
  NAND U21511 ( .A(B[1]), .B(A[1]), .Z(n17152) );
endmodule


module mult_N1024_CC256 ( clk, rst, a, b, c );
  input [1023:0] a;
  input [3:0] b;
  output [1023:0] c;
  input clk, rst;

  wire   [1023:4] swire;
  wire   [1023:0] clocal;
  wire   [2047:1024] sreg;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;

  DFF \sreg_reg[1024]  ( .D(swire[4]), .CLK(clk), .RST(rst), .Q(sreg[1024]) );
  DFF \sreg_reg[1025]  ( .D(swire[5]), .CLK(clk), .RST(rst), .Q(sreg[1025]) );
  DFF \sreg_reg[1026]  ( .D(swire[6]), .CLK(clk), .RST(rst), .Q(sreg[1026]) );
  DFF \sreg_reg[1027]  ( .D(swire[7]), .CLK(clk), .RST(rst), .Q(sreg[1027]) );
  DFF \sreg_reg[1028]  ( .D(swire[8]), .CLK(clk), .RST(rst), .Q(sreg[1028]) );
  DFF \sreg_reg[1029]  ( .D(swire[9]), .CLK(clk), .RST(rst), .Q(sreg[1029]) );
  DFF \sreg_reg[1030]  ( .D(swire[10]), .CLK(clk), .RST(rst), .Q(sreg[1030])
         );
  DFF \sreg_reg[1031]  ( .D(swire[11]), .CLK(clk), .RST(rst), .Q(sreg[1031])
         );
  DFF \sreg_reg[1032]  ( .D(swire[12]), .CLK(clk), .RST(rst), .Q(sreg[1032])
         );
  DFF \sreg_reg[1033]  ( .D(swire[13]), .CLK(clk), .RST(rst), .Q(sreg[1033])
         );
  DFF \sreg_reg[1034]  ( .D(swire[14]), .CLK(clk), .RST(rst), .Q(sreg[1034])
         );
  DFF \sreg_reg[1035]  ( .D(swire[15]), .CLK(clk), .RST(rst), .Q(sreg[1035])
         );
  DFF \sreg_reg[1036]  ( .D(swire[16]), .CLK(clk), .RST(rst), .Q(sreg[1036])
         );
  DFF \sreg_reg[1037]  ( .D(swire[17]), .CLK(clk), .RST(rst), .Q(sreg[1037])
         );
  DFF \sreg_reg[1038]  ( .D(swire[18]), .CLK(clk), .RST(rst), .Q(sreg[1038])
         );
  DFF \sreg_reg[1039]  ( .D(swire[19]), .CLK(clk), .RST(rst), .Q(sreg[1039])
         );
  DFF \sreg_reg[1040]  ( .D(swire[20]), .CLK(clk), .RST(rst), .Q(sreg[1040])
         );
  DFF \sreg_reg[1041]  ( .D(swire[21]), .CLK(clk), .RST(rst), .Q(sreg[1041])
         );
  DFF \sreg_reg[1042]  ( .D(swire[22]), .CLK(clk), .RST(rst), .Q(sreg[1042])
         );
  DFF \sreg_reg[1043]  ( .D(swire[23]), .CLK(clk), .RST(rst), .Q(sreg[1043])
         );
  DFF \sreg_reg[1044]  ( .D(swire[24]), .CLK(clk), .RST(rst), .Q(sreg[1044])
         );
  DFF \sreg_reg[1045]  ( .D(swire[25]), .CLK(clk), .RST(rst), .Q(sreg[1045])
         );
  DFF \sreg_reg[1046]  ( .D(swire[26]), .CLK(clk), .RST(rst), .Q(sreg[1046])
         );
  DFF \sreg_reg[1047]  ( .D(swire[27]), .CLK(clk), .RST(rst), .Q(sreg[1047])
         );
  DFF \sreg_reg[1048]  ( .D(swire[28]), .CLK(clk), .RST(rst), .Q(sreg[1048])
         );
  DFF \sreg_reg[1049]  ( .D(swire[29]), .CLK(clk), .RST(rst), .Q(sreg[1049])
         );
  DFF \sreg_reg[1050]  ( .D(swire[30]), .CLK(clk), .RST(rst), .Q(sreg[1050])
         );
  DFF \sreg_reg[1051]  ( .D(swire[31]), .CLK(clk), .RST(rst), .Q(sreg[1051])
         );
  DFF \sreg_reg[1052]  ( .D(swire[32]), .CLK(clk), .RST(rst), .Q(sreg[1052])
         );
  DFF \sreg_reg[1053]  ( .D(swire[33]), .CLK(clk), .RST(rst), .Q(sreg[1053])
         );
  DFF \sreg_reg[1054]  ( .D(swire[34]), .CLK(clk), .RST(rst), .Q(sreg[1054])
         );
  DFF \sreg_reg[1055]  ( .D(swire[35]), .CLK(clk), .RST(rst), .Q(sreg[1055])
         );
  DFF \sreg_reg[1056]  ( .D(swire[36]), .CLK(clk), .RST(rst), .Q(sreg[1056])
         );
  DFF \sreg_reg[1057]  ( .D(swire[37]), .CLK(clk), .RST(rst), .Q(sreg[1057])
         );
  DFF \sreg_reg[1058]  ( .D(swire[38]), .CLK(clk), .RST(rst), .Q(sreg[1058])
         );
  DFF \sreg_reg[1059]  ( .D(swire[39]), .CLK(clk), .RST(rst), .Q(sreg[1059])
         );
  DFF \sreg_reg[1060]  ( .D(swire[40]), .CLK(clk), .RST(rst), .Q(sreg[1060])
         );
  DFF \sreg_reg[1061]  ( .D(swire[41]), .CLK(clk), .RST(rst), .Q(sreg[1061])
         );
  DFF \sreg_reg[1062]  ( .D(swire[42]), .CLK(clk), .RST(rst), .Q(sreg[1062])
         );
  DFF \sreg_reg[1063]  ( .D(swire[43]), .CLK(clk), .RST(rst), .Q(sreg[1063])
         );
  DFF \sreg_reg[1064]  ( .D(swire[44]), .CLK(clk), .RST(rst), .Q(sreg[1064])
         );
  DFF \sreg_reg[1065]  ( .D(swire[45]), .CLK(clk), .RST(rst), .Q(sreg[1065])
         );
  DFF \sreg_reg[1066]  ( .D(swire[46]), .CLK(clk), .RST(rst), .Q(sreg[1066])
         );
  DFF \sreg_reg[1067]  ( .D(swire[47]), .CLK(clk), .RST(rst), .Q(sreg[1067])
         );
  DFF \sreg_reg[1068]  ( .D(swire[48]), .CLK(clk), .RST(rst), .Q(sreg[1068])
         );
  DFF \sreg_reg[1069]  ( .D(swire[49]), .CLK(clk), .RST(rst), .Q(sreg[1069])
         );
  DFF \sreg_reg[1070]  ( .D(swire[50]), .CLK(clk), .RST(rst), .Q(sreg[1070])
         );
  DFF \sreg_reg[1071]  ( .D(swire[51]), .CLK(clk), .RST(rst), .Q(sreg[1071])
         );
  DFF \sreg_reg[1072]  ( .D(swire[52]), .CLK(clk), .RST(rst), .Q(sreg[1072])
         );
  DFF \sreg_reg[1073]  ( .D(swire[53]), .CLK(clk), .RST(rst), .Q(sreg[1073])
         );
  DFF \sreg_reg[1074]  ( .D(swire[54]), .CLK(clk), .RST(rst), .Q(sreg[1074])
         );
  DFF \sreg_reg[1075]  ( .D(swire[55]), .CLK(clk), .RST(rst), .Q(sreg[1075])
         );
  DFF \sreg_reg[1076]  ( .D(swire[56]), .CLK(clk), .RST(rst), .Q(sreg[1076])
         );
  DFF \sreg_reg[1077]  ( .D(swire[57]), .CLK(clk), .RST(rst), .Q(sreg[1077])
         );
  DFF \sreg_reg[1078]  ( .D(swire[58]), .CLK(clk), .RST(rst), .Q(sreg[1078])
         );
  DFF \sreg_reg[1079]  ( .D(swire[59]), .CLK(clk), .RST(rst), .Q(sreg[1079])
         );
  DFF \sreg_reg[1080]  ( .D(swire[60]), .CLK(clk), .RST(rst), .Q(sreg[1080])
         );
  DFF \sreg_reg[1081]  ( .D(swire[61]), .CLK(clk), .RST(rst), .Q(sreg[1081])
         );
  DFF \sreg_reg[1082]  ( .D(swire[62]), .CLK(clk), .RST(rst), .Q(sreg[1082])
         );
  DFF \sreg_reg[1083]  ( .D(swire[63]), .CLK(clk), .RST(rst), .Q(sreg[1083])
         );
  DFF \sreg_reg[1084]  ( .D(swire[64]), .CLK(clk), .RST(rst), .Q(sreg[1084])
         );
  DFF \sreg_reg[1085]  ( .D(swire[65]), .CLK(clk), .RST(rst), .Q(sreg[1085])
         );
  DFF \sreg_reg[1086]  ( .D(swire[66]), .CLK(clk), .RST(rst), .Q(sreg[1086])
         );
  DFF \sreg_reg[1087]  ( .D(swire[67]), .CLK(clk), .RST(rst), .Q(sreg[1087])
         );
  DFF \sreg_reg[1088]  ( .D(swire[68]), .CLK(clk), .RST(rst), .Q(sreg[1088])
         );
  DFF \sreg_reg[1089]  ( .D(swire[69]), .CLK(clk), .RST(rst), .Q(sreg[1089])
         );
  DFF \sreg_reg[1090]  ( .D(swire[70]), .CLK(clk), .RST(rst), .Q(sreg[1090])
         );
  DFF \sreg_reg[1091]  ( .D(swire[71]), .CLK(clk), .RST(rst), .Q(sreg[1091])
         );
  DFF \sreg_reg[1092]  ( .D(swire[72]), .CLK(clk), .RST(rst), .Q(sreg[1092])
         );
  DFF \sreg_reg[1093]  ( .D(swire[73]), .CLK(clk), .RST(rst), .Q(sreg[1093])
         );
  DFF \sreg_reg[1094]  ( .D(swire[74]), .CLK(clk), .RST(rst), .Q(sreg[1094])
         );
  DFF \sreg_reg[1095]  ( .D(swire[75]), .CLK(clk), .RST(rst), .Q(sreg[1095])
         );
  DFF \sreg_reg[1096]  ( .D(swire[76]), .CLK(clk), .RST(rst), .Q(sreg[1096])
         );
  DFF \sreg_reg[1097]  ( .D(swire[77]), .CLK(clk), .RST(rst), .Q(sreg[1097])
         );
  DFF \sreg_reg[1098]  ( .D(swire[78]), .CLK(clk), .RST(rst), .Q(sreg[1098])
         );
  DFF \sreg_reg[1099]  ( .D(swire[79]), .CLK(clk), .RST(rst), .Q(sreg[1099])
         );
  DFF \sreg_reg[1100]  ( .D(swire[80]), .CLK(clk), .RST(rst), .Q(sreg[1100])
         );
  DFF \sreg_reg[1101]  ( .D(swire[81]), .CLK(clk), .RST(rst), .Q(sreg[1101])
         );
  DFF \sreg_reg[1102]  ( .D(swire[82]), .CLK(clk), .RST(rst), .Q(sreg[1102])
         );
  DFF \sreg_reg[1103]  ( .D(swire[83]), .CLK(clk), .RST(rst), .Q(sreg[1103])
         );
  DFF \sreg_reg[1104]  ( .D(swire[84]), .CLK(clk), .RST(rst), .Q(sreg[1104])
         );
  DFF \sreg_reg[1105]  ( .D(swire[85]), .CLK(clk), .RST(rst), .Q(sreg[1105])
         );
  DFF \sreg_reg[1106]  ( .D(swire[86]), .CLK(clk), .RST(rst), .Q(sreg[1106])
         );
  DFF \sreg_reg[1107]  ( .D(swire[87]), .CLK(clk), .RST(rst), .Q(sreg[1107])
         );
  DFF \sreg_reg[1108]  ( .D(swire[88]), .CLK(clk), .RST(rst), .Q(sreg[1108])
         );
  DFF \sreg_reg[1109]  ( .D(swire[89]), .CLK(clk), .RST(rst), .Q(sreg[1109])
         );
  DFF \sreg_reg[1110]  ( .D(swire[90]), .CLK(clk), .RST(rst), .Q(sreg[1110])
         );
  DFF \sreg_reg[1111]  ( .D(swire[91]), .CLK(clk), .RST(rst), .Q(sreg[1111])
         );
  DFF \sreg_reg[1112]  ( .D(swire[92]), .CLK(clk), .RST(rst), .Q(sreg[1112])
         );
  DFF \sreg_reg[1113]  ( .D(swire[93]), .CLK(clk), .RST(rst), .Q(sreg[1113])
         );
  DFF \sreg_reg[1114]  ( .D(swire[94]), .CLK(clk), .RST(rst), .Q(sreg[1114])
         );
  DFF \sreg_reg[1115]  ( .D(swire[95]), .CLK(clk), .RST(rst), .Q(sreg[1115])
         );
  DFF \sreg_reg[1116]  ( .D(swire[96]), .CLK(clk), .RST(rst), .Q(sreg[1116])
         );
  DFF \sreg_reg[1117]  ( .D(swire[97]), .CLK(clk), .RST(rst), .Q(sreg[1117])
         );
  DFF \sreg_reg[1118]  ( .D(swire[98]), .CLK(clk), .RST(rst), .Q(sreg[1118])
         );
  DFF \sreg_reg[1119]  ( .D(swire[99]), .CLK(clk), .RST(rst), .Q(sreg[1119])
         );
  DFF \sreg_reg[1120]  ( .D(swire[100]), .CLK(clk), .RST(rst), .Q(sreg[1120])
         );
  DFF \sreg_reg[1121]  ( .D(swire[101]), .CLK(clk), .RST(rst), .Q(sreg[1121])
         );
  DFF \sreg_reg[1122]  ( .D(swire[102]), .CLK(clk), .RST(rst), .Q(sreg[1122])
         );
  DFF \sreg_reg[1123]  ( .D(swire[103]), .CLK(clk), .RST(rst), .Q(sreg[1123])
         );
  DFF \sreg_reg[1124]  ( .D(swire[104]), .CLK(clk), .RST(rst), .Q(sreg[1124])
         );
  DFF \sreg_reg[1125]  ( .D(swire[105]), .CLK(clk), .RST(rst), .Q(sreg[1125])
         );
  DFF \sreg_reg[1126]  ( .D(swire[106]), .CLK(clk), .RST(rst), .Q(sreg[1126])
         );
  DFF \sreg_reg[1127]  ( .D(swire[107]), .CLK(clk), .RST(rst), .Q(sreg[1127])
         );
  DFF \sreg_reg[1128]  ( .D(swire[108]), .CLK(clk), .RST(rst), .Q(sreg[1128])
         );
  DFF \sreg_reg[1129]  ( .D(swire[109]), .CLK(clk), .RST(rst), .Q(sreg[1129])
         );
  DFF \sreg_reg[1130]  ( .D(swire[110]), .CLK(clk), .RST(rst), .Q(sreg[1130])
         );
  DFF \sreg_reg[1131]  ( .D(swire[111]), .CLK(clk), .RST(rst), .Q(sreg[1131])
         );
  DFF \sreg_reg[1132]  ( .D(swire[112]), .CLK(clk), .RST(rst), .Q(sreg[1132])
         );
  DFF \sreg_reg[1133]  ( .D(swire[113]), .CLK(clk), .RST(rst), .Q(sreg[1133])
         );
  DFF \sreg_reg[1134]  ( .D(swire[114]), .CLK(clk), .RST(rst), .Q(sreg[1134])
         );
  DFF \sreg_reg[1135]  ( .D(swire[115]), .CLK(clk), .RST(rst), .Q(sreg[1135])
         );
  DFF \sreg_reg[1136]  ( .D(swire[116]), .CLK(clk), .RST(rst), .Q(sreg[1136])
         );
  DFF \sreg_reg[1137]  ( .D(swire[117]), .CLK(clk), .RST(rst), .Q(sreg[1137])
         );
  DFF \sreg_reg[1138]  ( .D(swire[118]), .CLK(clk), .RST(rst), .Q(sreg[1138])
         );
  DFF \sreg_reg[1139]  ( .D(swire[119]), .CLK(clk), .RST(rst), .Q(sreg[1139])
         );
  DFF \sreg_reg[1140]  ( .D(swire[120]), .CLK(clk), .RST(rst), .Q(sreg[1140])
         );
  DFF \sreg_reg[1141]  ( .D(swire[121]), .CLK(clk), .RST(rst), .Q(sreg[1141])
         );
  DFF \sreg_reg[1142]  ( .D(swire[122]), .CLK(clk), .RST(rst), .Q(sreg[1142])
         );
  DFF \sreg_reg[1143]  ( .D(swire[123]), .CLK(clk), .RST(rst), .Q(sreg[1143])
         );
  DFF \sreg_reg[1144]  ( .D(swire[124]), .CLK(clk), .RST(rst), .Q(sreg[1144])
         );
  DFF \sreg_reg[1145]  ( .D(swire[125]), .CLK(clk), .RST(rst), .Q(sreg[1145])
         );
  DFF \sreg_reg[1146]  ( .D(swire[126]), .CLK(clk), .RST(rst), .Q(sreg[1146])
         );
  DFF \sreg_reg[1147]  ( .D(swire[127]), .CLK(clk), .RST(rst), .Q(sreg[1147])
         );
  DFF \sreg_reg[1148]  ( .D(swire[128]), .CLK(clk), .RST(rst), .Q(sreg[1148])
         );
  DFF \sreg_reg[1149]  ( .D(swire[129]), .CLK(clk), .RST(rst), .Q(sreg[1149])
         );
  DFF \sreg_reg[1150]  ( .D(swire[130]), .CLK(clk), .RST(rst), .Q(sreg[1150])
         );
  DFF \sreg_reg[1151]  ( .D(swire[131]), .CLK(clk), .RST(rst), .Q(sreg[1151])
         );
  DFF \sreg_reg[1152]  ( .D(swire[132]), .CLK(clk), .RST(rst), .Q(sreg[1152])
         );
  DFF \sreg_reg[1153]  ( .D(swire[133]), .CLK(clk), .RST(rst), .Q(sreg[1153])
         );
  DFF \sreg_reg[1154]  ( .D(swire[134]), .CLK(clk), .RST(rst), .Q(sreg[1154])
         );
  DFF \sreg_reg[1155]  ( .D(swire[135]), .CLK(clk), .RST(rst), .Q(sreg[1155])
         );
  DFF \sreg_reg[1156]  ( .D(swire[136]), .CLK(clk), .RST(rst), .Q(sreg[1156])
         );
  DFF \sreg_reg[1157]  ( .D(swire[137]), .CLK(clk), .RST(rst), .Q(sreg[1157])
         );
  DFF \sreg_reg[1158]  ( .D(swire[138]), .CLK(clk), .RST(rst), .Q(sreg[1158])
         );
  DFF \sreg_reg[1159]  ( .D(swire[139]), .CLK(clk), .RST(rst), .Q(sreg[1159])
         );
  DFF \sreg_reg[1160]  ( .D(swire[140]), .CLK(clk), .RST(rst), .Q(sreg[1160])
         );
  DFF \sreg_reg[1161]  ( .D(swire[141]), .CLK(clk), .RST(rst), .Q(sreg[1161])
         );
  DFF \sreg_reg[1162]  ( .D(swire[142]), .CLK(clk), .RST(rst), .Q(sreg[1162])
         );
  DFF \sreg_reg[1163]  ( .D(swire[143]), .CLK(clk), .RST(rst), .Q(sreg[1163])
         );
  DFF \sreg_reg[1164]  ( .D(swire[144]), .CLK(clk), .RST(rst), .Q(sreg[1164])
         );
  DFF \sreg_reg[1165]  ( .D(swire[145]), .CLK(clk), .RST(rst), .Q(sreg[1165])
         );
  DFF \sreg_reg[1166]  ( .D(swire[146]), .CLK(clk), .RST(rst), .Q(sreg[1166])
         );
  DFF \sreg_reg[1167]  ( .D(swire[147]), .CLK(clk), .RST(rst), .Q(sreg[1167])
         );
  DFF \sreg_reg[1168]  ( .D(swire[148]), .CLK(clk), .RST(rst), .Q(sreg[1168])
         );
  DFF \sreg_reg[1169]  ( .D(swire[149]), .CLK(clk), .RST(rst), .Q(sreg[1169])
         );
  DFF \sreg_reg[1170]  ( .D(swire[150]), .CLK(clk), .RST(rst), .Q(sreg[1170])
         );
  DFF \sreg_reg[1171]  ( .D(swire[151]), .CLK(clk), .RST(rst), .Q(sreg[1171])
         );
  DFF \sreg_reg[1172]  ( .D(swire[152]), .CLK(clk), .RST(rst), .Q(sreg[1172])
         );
  DFF \sreg_reg[1173]  ( .D(swire[153]), .CLK(clk), .RST(rst), .Q(sreg[1173])
         );
  DFF \sreg_reg[1174]  ( .D(swire[154]), .CLK(clk), .RST(rst), .Q(sreg[1174])
         );
  DFF \sreg_reg[1175]  ( .D(swire[155]), .CLK(clk), .RST(rst), .Q(sreg[1175])
         );
  DFF \sreg_reg[1176]  ( .D(swire[156]), .CLK(clk), .RST(rst), .Q(sreg[1176])
         );
  DFF \sreg_reg[1177]  ( .D(swire[157]), .CLK(clk), .RST(rst), .Q(sreg[1177])
         );
  DFF \sreg_reg[1178]  ( .D(swire[158]), .CLK(clk), .RST(rst), .Q(sreg[1178])
         );
  DFF \sreg_reg[1179]  ( .D(swire[159]), .CLK(clk), .RST(rst), .Q(sreg[1179])
         );
  DFF \sreg_reg[1180]  ( .D(swire[160]), .CLK(clk), .RST(rst), .Q(sreg[1180])
         );
  DFF \sreg_reg[1181]  ( .D(swire[161]), .CLK(clk), .RST(rst), .Q(sreg[1181])
         );
  DFF \sreg_reg[1182]  ( .D(swire[162]), .CLK(clk), .RST(rst), .Q(sreg[1182])
         );
  DFF \sreg_reg[1183]  ( .D(swire[163]), .CLK(clk), .RST(rst), .Q(sreg[1183])
         );
  DFF \sreg_reg[1184]  ( .D(swire[164]), .CLK(clk), .RST(rst), .Q(sreg[1184])
         );
  DFF \sreg_reg[1185]  ( .D(swire[165]), .CLK(clk), .RST(rst), .Q(sreg[1185])
         );
  DFF \sreg_reg[1186]  ( .D(swire[166]), .CLK(clk), .RST(rst), .Q(sreg[1186])
         );
  DFF \sreg_reg[1187]  ( .D(swire[167]), .CLK(clk), .RST(rst), .Q(sreg[1187])
         );
  DFF \sreg_reg[1188]  ( .D(swire[168]), .CLK(clk), .RST(rst), .Q(sreg[1188])
         );
  DFF \sreg_reg[1189]  ( .D(swire[169]), .CLK(clk), .RST(rst), .Q(sreg[1189])
         );
  DFF \sreg_reg[1190]  ( .D(swire[170]), .CLK(clk), .RST(rst), .Q(sreg[1190])
         );
  DFF \sreg_reg[1191]  ( .D(swire[171]), .CLK(clk), .RST(rst), .Q(sreg[1191])
         );
  DFF \sreg_reg[1192]  ( .D(swire[172]), .CLK(clk), .RST(rst), .Q(sreg[1192])
         );
  DFF \sreg_reg[1193]  ( .D(swire[173]), .CLK(clk), .RST(rst), .Q(sreg[1193])
         );
  DFF \sreg_reg[1194]  ( .D(swire[174]), .CLK(clk), .RST(rst), .Q(sreg[1194])
         );
  DFF \sreg_reg[1195]  ( .D(swire[175]), .CLK(clk), .RST(rst), .Q(sreg[1195])
         );
  DFF \sreg_reg[1196]  ( .D(swire[176]), .CLK(clk), .RST(rst), .Q(sreg[1196])
         );
  DFF \sreg_reg[1197]  ( .D(swire[177]), .CLK(clk), .RST(rst), .Q(sreg[1197])
         );
  DFF \sreg_reg[1198]  ( .D(swire[178]), .CLK(clk), .RST(rst), .Q(sreg[1198])
         );
  DFF \sreg_reg[1199]  ( .D(swire[179]), .CLK(clk), .RST(rst), .Q(sreg[1199])
         );
  DFF \sreg_reg[1200]  ( .D(swire[180]), .CLK(clk), .RST(rst), .Q(sreg[1200])
         );
  DFF \sreg_reg[1201]  ( .D(swire[181]), .CLK(clk), .RST(rst), .Q(sreg[1201])
         );
  DFF \sreg_reg[1202]  ( .D(swire[182]), .CLK(clk), .RST(rst), .Q(sreg[1202])
         );
  DFF \sreg_reg[1203]  ( .D(swire[183]), .CLK(clk), .RST(rst), .Q(sreg[1203])
         );
  DFF \sreg_reg[1204]  ( .D(swire[184]), .CLK(clk), .RST(rst), .Q(sreg[1204])
         );
  DFF \sreg_reg[1205]  ( .D(swire[185]), .CLK(clk), .RST(rst), .Q(sreg[1205])
         );
  DFF \sreg_reg[1206]  ( .D(swire[186]), .CLK(clk), .RST(rst), .Q(sreg[1206])
         );
  DFF \sreg_reg[1207]  ( .D(swire[187]), .CLK(clk), .RST(rst), .Q(sreg[1207])
         );
  DFF \sreg_reg[1208]  ( .D(swire[188]), .CLK(clk), .RST(rst), .Q(sreg[1208])
         );
  DFF \sreg_reg[1209]  ( .D(swire[189]), .CLK(clk), .RST(rst), .Q(sreg[1209])
         );
  DFF \sreg_reg[1210]  ( .D(swire[190]), .CLK(clk), .RST(rst), .Q(sreg[1210])
         );
  DFF \sreg_reg[1211]  ( .D(swire[191]), .CLK(clk), .RST(rst), .Q(sreg[1211])
         );
  DFF \sreg_reg[1212]  ( .D(swire[192]), .CLK(clk), .RST(rst), .Q(sreg[1212])
         );
  DFF \sreg_reg[1213]  ( .D(swire[193]), .CLK(clk), .RST(rst), .Q(sreg[1213])
         );
  DFF \sreg_reg[1214]  ( .D(swire[194]), .CLK(clk), .RST(rst), .Q(sreg[1214])
         );
  DFF \sreg_reg[1215]  ( .D(swire[195]), .CLK(clk), .RST(rst), .Q(sreg[1215])
         );
  DFF \sreg_reg[1216]  ( .D(swire[196]), .CLK(clk), .RST(rst), .Q(sreg[1216])
         );
  DFF \sreg_reg[1217]  ( .D(swire[197]), .CLK(clk), .RST(rst), .Q(sreg[1217])
         );
  DFF \sreg_reg[1218]  ( .D(swire[198]), .CLK(clk), .RST(rst), .Q(sreg[1218])
         );
  DFF \sreg_reg[1219]  ( .D(swire[199]), .CLK(clk), .RST(rst), .Q(sreg[1219])
         );
  DFF \sreg_reg[1220]  ( .D(swire[200]), .CLK(clk), .RST(rst), .Q(sreg[1220])
         );
  DFF \sreg_reg[1221]  ( .D(swire[201]), .CLK(clk), .RST(rst), .Q(sreg[1221])
         );
  DFF \sreg_reg[1222]  ( .D(swire[202]), .CLK(clk), .RST(rst), .Q(sreg[1222])
         );
  DFF \sreg_reg[1223]  ( .D(swire[203]), .CLK(clk), .RST(rst), .Q(sreg[1223])
         );
  DFF \sreg_reg[1224]  ( .D(swire[204]), .CLK(clk), .RST(rst), .Q(sreg[1224])
         );
  DFF \sreg_reg[1225]  ( .D(swire[205]), .CLK(clk), .RST(rst), .Q(sreg[1225])
         );
  DFF \sreg_reg[1226]  ( .D(swire[206]), .CLK(clk), .RST(rst), .Q(sreg[1226])
         );
  DFF \sreg_reg[1227]  ( .D(swire[207]), .CLK(clk), .RST(rst), .Q(sreg[1227])
         );
  DFF \sreg_reg[1228]  ( .D(swire[208]), .CLK(clk), .RST(rst), .Q(sreg[1228])
         );
  DFF \sreg_reg[1229]  ( .D(swire[209]), .CLK(clk), .RST(rst), .Q(sreg[1229])
         );
  DFF \sreg_reg[1230]  ( .D(swire[210]), .CLK(clk), .RST(rst), .Q(sreg[1230])
         );
  DFF \sreg_reg[1231]  ( .D(swire[211]), .CLK(clk), .RST(rst), .Q(sreg[1231])
         );
  DFF \sreg_reg[1232]  ( .D(swire[212]), .CLK(clk), .RST(rst), .Q(sreg[1232])
         );
  DFF \sreg_reg[1233]  ( .D(swire[213]), .CLK(clk), .RST(rst), .Q(sreg[1233])
         );
  DFF \sreg_reg[1234]  ( .D(swire[214]), .CLK(clk), .RST(rst), .Q(sreg[1234])
         );
  DFF \sreg_reg[1235]  ( .D(swire[215]), .CLK(clk), .RST(rst), .Q(sreg[1235])
         );
  DFF \sreg_reg[1236]  ( .D(swire[216]), .CLK(clk), .RST(rst), .Q(sreg[1236])
         );
  DFF \sreg_reg[1237]  ( .D(swire[217]), .CLK(clk), .RST(rst), .Q(sreg[1237])
         );
  DFF \sreg_reg[1238]  ( .D(swire[218]), .CLK(clk), .RST(rst), .Q(sreg[1238])
         );
  DFF \sreg_reg[1239]  ( .D(swire[219]), .CLK(clk), .RST(rst), .Q(sreg[1239])
         );
  DFF \sreg_reg[1240]  ( .D(swire[220]), .CLK(clk), .RST(rst), .Q(sreg[1240])
         );
  DFF \sreg_reg[1241]  ( .D(swire[221]), .CLK(clk), .RST(rst), .Q(sreg[1241])
         );
  DFF \sreg_reg[1242]  ( .D(swire[222]), .CLK(clk), .RST(rst), .Q(sreg[1242])
         );
  DFF \sreg_reg[1243]  ( .D(swire[223]), .CLK(clk), .RST(rst), .Q(sreg[1243])
         );
  DFF \sreg_reg[1244]  ( .D(swire[224]), .CLK(clk), .RST(rst), .Q(sreg[1244])
         );
  DFF \sreg_reg[1245]  ( .D(swire[225]), .CLK(clk), .RST(rst), .Q(sreg[1245])
         );
  DFF \sreg_reg[1246]  ( .D(swire[226]), .CLK(clk), .RST(rst), .Q(sreg[1246])
         );
  DFF \sreg_reg[1247]  ( .D(swire[227]), .CLK(clk), .RST(rst), .Q(sreg[1247])
         );
  DFF \sreg_reg[1248]  ( .D(swire[228]), .CLK(clk), .RST(rst), .Q(sreg[1248])
         );
  DFF \sreg_reg[1249]  ( .D(swire[229]), .CLK(clk), .RST(rst), .Q(sreg[1249])
         );
  DFF \sreg_reg[1250]  ( .D(swire[230]), .CLK(clk), .RST(rst), .Q(sreg[1250])
         );
  DFF \sreg_reg[1251]  ( .D(swire[231]), .CLK(clk), .RST(rst), .Q(sreg[1251])
         );
  DFF \sreg_reg[1252]  ( .D(swire[232]), .CLK(clk), .RST(rst), .Q(sreg[1252])
         );
  DFF \sreg_reg[1253]  ( .D(swire[233]), .CLK(clk), .RST(rst), .Q(sreg[1253])
         );
  DFF \sreg_reg[1254]  ( .D(swire[234]), .CLK(clk), .RST(rst), .Q(sreg[1254])
         );
  DFF \sreg_reg[1255]  ( .D(swire[235]), .CLK(clk), .RST(rst), .Q(sreg[1255])
         );
  DFF \sreg_reg[1256]  ( .D(swire[236]), .CLK(clk), .RST(rst), .Q(sreg[1256])
         );
  DFF \sreg_reg[1257]  ( .D(swire[237]), .CLK(clk), .RST(rst), .Q(sreg[1257])
         );
  DFF \sreg_reg[1258]  ( .D(swire[238]), .CLK(clk), .RST(rst), .Q(sreg[1258])
         );
  DFF \sreg_reg[1259]  ( .D(swire[239]), .CLK(clk), .RST(rst), .Q(sreg[1259])
         );
  DFF \sreg_reg[1260]  ( .D(swire[240]), .CLK(clk), .RST(rst), .Q(sreg[1260])
         );
  DFF \sreg_reg[1261]  ( .D(swire[241]), .CLK(clk), .RST(rst), .Q(sreg[1261])
         );
  DFF \sreg_reg[1262]  ( .D(swire[242]), .CLK(clk), .RST(rst), .Q(sreg[1262])
         );
  DFF \sreg_reg[1263]  ( .D(swire[243]), .CLK(clk), .RST(rst), .Q(sreg[1263])
         );
  DFF \sreg_reg[1264]  ( .D(swire[244]), .CLK(clk), .RST(rst), .Q(sreg[1264])
         );
  DFF \sreg_reg[1265]  ( .D(swire[245]), .CLK(clk), .RST(rst), .Q(sreg[1265])
         );
  DFF \sreg_reg[1266]  ( .D(swire[246]), .CLK(clk), .RST(rst), .Q(sreg[1266])
         );
  DFF \sreg_reg[1267]  ( .D(swire[247]), .CLK(clk), .RST(rst), .Q(sreg[1267])
         );
  DFF \sreg_reg[1268]  ( .D(swire[248]), .CLK(clk), .RST(rst), .Q(sreg[1268])
         );
  DFF \sreg_reg[1269]  ( .D(swire[249]), .CLK(clk), .RST(rst), .Q(sreg[1269])
         );
  DFF \sreg_reg[1270]  ( .D(swire[250]), .CLK(clk), .RST(rst), .Q(sreg[1270])
         );
  DFF \sreg_reg[1271]  ( .D(swire[251]), .CLK(clk), .RST(rst), .Q(sreg[1271])
         );
  DFF \sreg_reg[1272]  ( .D(swire[252]), .CLK(clk), .RST(rst), .Q(sreg[1272])
         );
  DFF \sreg_reg[1273]  ( .D(swire[253]), .CLK(clk), .RST(rst), .Q(sreg[1273])
         );
  DFF \sreg_reg[1274]  ( .D(swire[254]), .CLK(clk), .RST(rst), .Q(sreg[1274])
         );
  DFF \sreg_reg[1275]  ( .D(swire[255]), .CLK(clk), .RST(rst), .Q(sreg[1275])
         );
  DFF \sreg_reg[1276]  ( .D(swire[256]), .CLK(clk), .RST(rst), .Q(sreg[1276])
         );
  DFF \sreg_reg[1277]  ( .D(swire[257]), .CLK(clk), .RST(rst), .Q(sreg[1277])
         );
  DFF \sreg_reg[1278]  ( .D(swire[258]), .CLK(clk), .RST(rst), .Q(sreg[1278])
         );
  DFF \sreg_reg[1279]  ( .D(swire[259]), .CLK(clk), .RST(rst), .Q(sreg[1279])
         );
  DFF \sreg_reg[1280]  ( .D(swire[260]), .CLK(clk), .RST(rst), .Q(sreg[1280])
         );
  DFF \sreg_reg[1281]  ( .D(swire[261]), .CLK(clk), .RST(rst), .Q(sreg[1281])
         );
  DFF \sreg_reg[1282]  ( .D(swire[262]), .CLK(clk), .RST(rst), .Q(sreg[1282])
         );
  DFF \sreg_reg[1283]  ( .D(swire[263]), .CLK(clk), .RST(rst), .Q(sreg[1283])
         );
  DFF \sreg_reg[1284]  ( .D(swire[264]), .CLK(clk), .RST(rst), .Q(sreg[1284])
         );
  DFF \sreg_reg[1285]  ( .D(swire[265]), .CLK(clk), .RST(rst), .Q(sreg[1285])
         );
  DFF \sreg_reg[1286]  ( .D(swire[266]), .CLK(clk), .RST(rst), .Q(sreg[1286])
         );
  DFF \sreg_reg[1287]  ( .D(swire[267]), .CLK(clk), .RST(rst), .Q(sreg[1287])
         );
  DFF \sreg_reg[1288]  ( .D(swire[268]), .CLK(clk), .RST(rst), .Q(sreg[1288])
         );
  DFF \sreg_reg[1289]  ( .D(swire[269]), .CLK(clk), .RST(rst), .Q(sreg[1289])
         );
  DFF \sreg_reg[1290]  ( .D(swire[270]), .CLK(clk), .RST(rst), .Q(sreg[1290])
         );
  DFF \sreg_reg[1291]  ( .D(swire[271]), .CLK(clk), .RST(rst), .Q(sreg[1291])
         );
  DFF \sreg_reg[1292]  ( .D(swire[272]), .CLK(clk), .RST(rst), .Q(sreg[1292])
         );
  DFF \sreg_reg[1293]  ( .D(swire[273]), .CLK(clk), .RST(rst), .Q(sreg[1293])
         );
  DFF \sreg_reg[1294]  ( .D(swire[274]), .CLK(clk), .RST(rst), .Q(sreg[1294])
         );
  DFF \sreg_reg[1295]  ( .D(swire[275]), .CLK(clk), .RST(rst), .Q(sreg[1295])
         );
  DFF \sreg_reg[1296]  ( .D(swire[276]), .CLK(clk), .RST(rst), .Q(sreg[1296])
         );
  DFF \sreg_reg[1297]  ( .D(swire[277]), .CLK(clk), .RST(rst), .Q(sreg[1297])
         );
  DFF \sreg_reg[1298]  ( .D(swire[278]), .CLK(clk), .RST(rst), .Q(sreg[1298])
         );
  DFF \sreg_reg[1299]  ( .D(swire[279]), .CLK(clk), .RST(rst), .Q(sreg[1299])
         );
  DFF \sreg_reg[1300]  ( .D(swire[280]), .CLK(clk), .RST(rst), .Q(sreg[1300])
         );
  DFF \sreg_reg[1301]  ( .D(swire[281]), .CLK(clk), .RST(rst), .Q(sreg[1301])
         );
  DFF \sreg_reg[1302]  ( .D(swire[282]), .CLK(clk), .RST(rst), .Q(sreg[1302])
         );
  DFF \sreg_reg[1303]  ( .D(swire[283]), .CLK(clk), .RST(rst), .Q(sreg[1303])
         );
  DFF \sreg_reg[1304]  ( .D(swire[284]), .CLK(clk), .RST(rst), .Q(sreg[1304])
         );
  DFF \sreg_reg[1305]  ( .D(swire[285]), .CLK(clk), .RST(rst), .Q(sreg[1305])
         );
  DFF \sreg_reg[1306]  ( .D(swire[286]), .CLK(clk), .RST(rst), .Q(sreg[1306])
         );
  DFF \sreg_reg[1307]  ( .D(swire[287]), .CLK(clk), .RST(rst), .Q(sreg[1307])
         );
  DFF \sreg_reg[1308]  ( .D(swire[288]), .CLK(clk), .RST(rst), .Q(sreg[1308])
         );
  DFF \sreg_reg[1309]  ( .D(swire[289]), .CLK(clk), .RST(rst), .Q(sreg[1309])
         );
  DFF \sreg_reg[1310]  ( .D(swire[290]), .CLK(clk), .RST(rst), .Q(sreg[1310])
         );
  DFF \sreg_reg[1311]  ( .D(swire[291]), .CLK(clk), .RST(rst), .Q(sreg[1311])
         );
  DFF \sreg_reg[1312]  ( .D(swire[292]), .CLK(clk), .RST(rst), .Q(sreg[1312])
         );
  DFF \sreg_reg[1313]  ( .D(swire[293]), .CLK(clk), .RST(rst), .Q(sreg[1313])
         );
  DFF \sreg_reg[1314]  ( .D(swire[294]), .CLK(clk), .RST(rst), .Q(sreg[1314])
         );
  DFF \sreg_reg[1315]  ( .D(swire[295]), .CLK(clk), .RST(rst), .Q(sreg[1315])
         );
  DFF \sreg_reg[1316]  ( .D(swire[296]), .CLK(clk), .RST(rst), .Q(sreg[1316])
         );
  DFF \sreg_reg[1317]  ( .D(swire[297]), .CLK(clk), .RST(rst), .Q(sreg[1317])
         );
  DFF \sreg_reg[1318]  ( .D(swire[298]), .CLK(clk), .RST(rst), .Q(sreg[1318])
         );
  DFF \sreg_reg[1319]  ( .D(swire[299]), .CLK(clk), .RST(rst), .Q(sreg[1319])
         );
  DFF \sreg_reg[1320]  ( .D(swire[300]), .CLK(clk), .RST(rst), .Q(sreg[1320])
         );
  DFF \sreg_reg[1321]  ( .D(swire[301]), .CLK(clk), .RST(rst), .Q(sreg[1321])
         );
  DFF \sreg_reg[1322]  ( .D(swire[302]), .CLK(clk), .RST(rst), .Q(sreg[1322])
         );
  DFF \sreg_reg[1323]  ( .D(swire[303]), .CLK(clk), .RST(rst), .Q(sreg[1323])
         );
  DFF \sreg_reg[1324]  ( .D(swire[304]), .CLK(clk), .RST(rst), .Q(sreg[1324])
         );
  DFF \sreg_reg[1325]  ( .D(swire[305]), .CLK(clk), .RST(rst), .Q(sreg[1325])
         );
  DFF \sreg_reg[1326]  ( .D(swire[306]), .CLK(clk), .RST(rst), .Q(sreg[1326])
         );
  DFF \sreg_reg[1327]  ( .D(swire[307]), .CLK(clk), .RST(rst), .Q(sreg[1327])
         );
  DFF \sreg_reg[1328]  ( .D(swire[308]), .CLK(clk), .RST(rst), .Q(sreg[1328])
         );
  DFF \sreg_reg[1329]  ( .D(swire[309]), .CLK(clk), .RST(rst), .Q(sreg[1329])
         );
  DFF \sreg_reg[1330]  ( .D(swire[310]), .CLK(clk), .RST(rst), .Q(sreg[1330])
         );
  DFF \sreg_reg[1331]  ( .D(swire[311]), .CLK(clk), .RST(rst), .Q(sreg[1331])
         );
  DFF \sreg_reg[1332]  ( .D(swire[312]), .CLK(clk), .RST(rst), .Q(sreg[1332])
         );
  DFF \sreg_reg[1333]  ( .D(swire[313]), .CLK(clk), .RST(rst), .Q(sreg[1333])
         );
  DFF \sreg_reg[1334]  ( .D(swire[314]), .CLK(clk), .RST(rst), .Q(sreg[1334])
         );
  DFF \sreg_reg[1335]  ( .D(swire[315]), .CLK(clk), .RST(rst), .Q(sreg[1335])
         );
  DFF \sreg_reg[1336]  ( .D(swire[316]), .CLK(clk), .RST(rst), .Q(sreg[1336])
         );
  DFF \sreg_reg[1337]  ( .D(swire[317]), .CLK(clk), .RST(rst), .Q(sreg[1337])
         );
  DFF \sreg_reg[1338]  ( .D(swire[318]), .CLK(clk), .RST(rst), .Q(sreg[1338])
         );
  DFF \sreg_reg[1339]  ( .D(swire[319]), .CLK(clk), .RST(rst), .Q(sreg[1339])
         );
  DFF \sreg_reg[1340]  ( .D(swire[320]), .CLK(clk), .RST(rst), .Q(sreg[1340])
         );
  DFF \sreg_reg[1341]  ( .D(swire[321]), .CLK(clk), .RST(rst), .Q(sreg[1341])
         );
  DFF \sreg_reg[1342]  ( .D(swire[322]), .CLK(clk), .RST(rst), .Q(sreg[1342])
         );
  DFF \sreg_reg[1343]  ( .D(swire[323]), .CLK(clk), .RST(rst), .Q(sreg[1343])
         );
  DFF \sreg_reg[1344]  ( .D(swire[324]), .CLK(clk), .RST(rst), .Q(sreg[1344])
         );
  DFF \sreg_reg[1345]  ( .D(swire[325]), .CLK(clk), .RST(rst), .Q(sreg[1345])
         );
  DFF \sreg_reg[1346]  ( .D(swire[326]), .CLK(clk), .RST(rst), .Q(sreg[1346])
         );
  DFF \sreg_reg[1347]  ( .D(swire[327]), .CLK(clk), .RST(rst), .Q(sreg[1347])
         );
  DFF \sreg_reg[1348]  ( .D(swire[328]), .CLK(clk), .RST(rst), .Q(sreg[1348])
         );
  DFF \sreg_reg[1349]  ( .D(swire[329]), .CLK(clk), .RST(rst), .Q(sreg[1349])
         );
  DFF \sreg_reg[1350]  ( .D(swire[330]), .CLK(clk), .RST(rst), .Q(sreg[1350])
         );
  DFF \sreg_reg[1351]  ( .D(swire[331]), .CLK(clk), .RST(rst), .Q(sreg[1351])
         );
  DFF \sreg_reg[1352]  ( .D(swire[332]), .CLK(clk), .RST(rst), .Q(sreg[1352])
         );
  DFF \sreg_reg[1353]  ( .D(swire[333]), .CLK(clk), .RST(rst), .Q(sreg[1353])
         );
  DFF \sreg_reg[1354]  ( .D(swire[334]), .CLK(clk), .RST(rst), .Q(sreg[1354])
         );
  DFF \sreg_reg[1355]  ( .D(swire[335]), .CLK(clk), .RST(rst), .Q(sreg[1355])
         );
  DFF \sreg_reg[1356]  ( .D(swire[336]), .CLK(clk), .RST(rst), .Q(sreg[1356])
         );
  DFF \sreg_reg[1357]  ( .D(swire[337]), .CLK(clk), .RST(rst), .Q(sreg[1357])
         );
  DFF \sreg_reg[1358]  ( .D(swire[338]), .CLK(clk), .RST(rst), .Q(sreg[1358])
         );
  DFF \sreg_reg[1359]  ( .D(swire[339]), .CLK(clk), .RST(rst), .Q(sreg[1359])
         );
  DFF \sreg_reg[1360]  ( .D(swire[340]), .CLK(clk), .RST(rst), .Q(sreg[1360])
         );
  DFF \sreg_reg[1361]  ( .D(swire[341]), .CLK(clk), .RST(rst), .Q(sreg[1361])
         );
  DFF \sreg_reg[1362]  ( .D(swire[342]), .CLK(clk), .RST(rst), .Q(sreg[1362])
         );
  DFF \sreg_reg[1363]  ( .D(swire[343]), .CLK(clk), .RST(rst), .Q(sreg[1363])
         );
  DFF \sreg_reg[1364]  ( .D(swire[344]), .CLK(clk), .RST(rst), .Q(sreg[1364])
         );
  DFF \sreg_reg[1365]  ( .D(swire[345]), .CLK(clk), .RST(rst), .Q(sreg[1365])
         );
  DFF \sreg_reg[1366]  ( .D(swire[346]), .CLK(clk), .RST(rst), .Q(sreg[1366])
         );
  DFF \sreg_reg[1367]  ( .D(swire[347]), .CLK(clk), .RST(rst), .Q(sreg[1367])
         );
  DFF \sreg_reg[1368]  ( .D(swire[348]), .CLK(clk), .RST(rst), .Q(sreg[1368])
         );
  DFF \sreg_reg[1369]  ( .D(swire[349]), .CLK(clk), .RST(rst), .Q(sreg[1369])
         );
  DFF \sreg_reg[1370]  ( .D(swire[350]), .CLK(clk), .RST(rst), .Q(sreg[1370])
         );
  DFF \sreg_reg[1371]  ( .D(swire[351]), .CLK(clk), .RST(rst), .Q(sreg[1371])
         );
  DFF \sreg_reg[1372]  ( .D(swire[352]), .CLK(clk), .RST(rst), .Q(sreg[1372])
         );
  DFF \sreg_reg[1373]  ( .D(swire[353]), .CLK(clk), .RST(rst), .Q(sreg[1373])
         );
  DFF \sreg_reg[1374]  ( .D(swire[354]), .CLK(clk), .RST(rst), .Q(sreg[1374])
         );
  DFF \sreg_reg[1375]  ( .D(swire[355]), .CLK(clk), .RST(rst), .Q(sreg[1375])
         );
  DFF \sreg_reg[1376]  ( .D(swire[356]), .CLK(clk), .RST(rst), .Q(sreg[1376])
         );
  DFF \sreg_reg[1377]  ( .D(swire[357]), .CLK(clk), .RST(rst), .Q(sreg[1377])
         );
  DFF \sreg_reg[1378]  ( .D(swire[358]), .CLK(clk), .RST(rst), .Q(sreg[1378])
         );
  DFF \sreg_reg[1379]  ( .D(swire[359]), .CLK(clk), .RST(rst), .Q(sreg[1379])
         );
  DFF \sreg_reg[1380]  ( .D(swire[360]), .CLK(clk), .RST(rst), .Q(sreg[1380])
         );
  DFF \sreg_reg[1381]  ( .D(swire[361]), .CLK(clk), .RST(rst), .Q(sreg[1381])
         );
  DFF \sreg_reg[1382]  ( .D(swire[362]), .CLK(clk), .RST(rst), .Q(sreg[1382])
         );
  DFF \sreg_reg[1383]  ( .D(swire[363]), .CLK(clk), .RST(rst), .Q(sreg[1383])
         );
  DFF \sreg_reg[1384]  ( .D(swire[364]), .CLK(clk), .RST(rst), .Q(sreg[1384])
         );
  DFF \sreg_reg[1385]  ( .D(swire[365]), .CLK(clk), .RST(rst), .Q(sreg[1385])
         );
  DFF \sreg_reg[1386]  ( .D(swire[366]), .CLK(clk), .RST(rst), .Q(sreg[1386])
         );
  DFF \sreg_reg[1387]  ( .D(swire[367]), .CLK(clk), .RST(rst), .Q(sreg[1387])
         );
  DFF \sreg_reg[1388]  ( .D(swire[368]), .CLK(clk), .RST(rst), .Q(sreg[1388])
         );
  DFF \sreg_reg[1389]  ( .D(swire[369]), .CLK(clk), .RST(rst), .Q(sreg[1389])
         );
  DFF \sreg_reg[1390]  ( .D(swire[370]), .CLK(clk), .RST(rst), .Q(sreg[1390])
         );
  DFF \sreg_reg[1391]  ( .D(swire[371]), .CLK(clk), .RST(rst), .Q(sreg[1391])
         );
  DFF \sreg_reg[1392]  ( .D(swire[372]), .CLK(clk), .RST(rst), .Q(sreg[1392])
         );
  DFF \sreg_reg[1393]  ( .D(swire[373]), .CLK(clk), .RST(rst), .Q(sreg[1393])
         );
  DFF \sreg_reg[1394]  ( .D(swire[374]), .CLK(clk), .RST(rst), .Q(sreg[1394])
         );
  DFF \sreg_reg[1395]  ( .D(swire[375]), .CLK(clk), .RST(rst), .Q(sreg[1395])
         );
  DFF \sreg_reg[1396]  ( .D(swire[376]), .CLK(clk), .RST(rst), .Q(sreg[1396])
         );
  DFF \sreg_reg[1397]  ( .D(swire[377]), .CLK(clk), .RST(rst), .Q(sreg[1397])
         );
  DFF \sreg_reg[1398]  ( .D(swire[378]), .CLK(clk), .RST(rst), .Q(sreg[1398])
         );
  DFF \sreg_reg[1399]  ( .D(swire[379]), .CLK(clk), .RST(rst), .Q(sreg[1399])
         );
  DFF \sreg_reg[1400]  ( .D(swire[380]), .CLK(clk), .RST(rst), .Q(sreg[1400])
         );
  DFF \sreg_reg[1401]  ( .D(swire[381]), .CLK(clk), .RST(rst), .Q(sreg[1401])
         );
  DFF \sreg_reg[1402]  ( .D(swire[382]), .CLK(clk), .RST(rst), .Q(sreg[1402])
         );
  DFF \sreg_reg[1403]  ( .D(swire[383]), .CLK(clk), .RST(rst), .Q(sreg[1403])
         );
  DFF \sreg_reg[1404]  ( .D(swire[384]), .CLK(clk), .RST(rst), .Q(sreg[1404])
         );
  DFF \sreg_reg[1405]  ( .D(swire[385]), .CLK(clk), .RST(rst), .Q(sreg[1405])
         );
  DFF \sreg_reg[1406]  ( .D(swire[386]), .CLK(clk), .RST(rst), .Q(sreg[1406])
         );
  DFF \sreg_reg[1407]  ( .D(swire[387]), .CLK(clk), .RST(rst), .Q(sreg[1407])
         );
  DFF \sreg_reg[1408]  ( .D(swire[388]), .CLK(clk), .RST(rst), .Q(sreg[1408])
         );
  DFF \sreg_reg[1409]  ( .D(swire[389]), .CLK(clk), .RST(rst), .Q(sreg[1409])
         );
  DFF \sreg_reg[1410]  ( .D(swire[390]), .CLK(clk), .RST(rst), .Q(sreg[1410])
         );
  DFF \sreg_reg[1411]  ( .D(swire[391]), .CLK(clk), .RST(rst), .Q(sreg[1411])
         );
  DFF \sreg_reg[1412]  ( .D(swire[392]), .CLK(clk), .RST(rst), .Q(sreg[1412])
         );
  DFF \sreg_reg[1413]  ( .D(swire[393]), .CLK(clk), .RST(rst), .Q(sreg[1413])
         );
  DFF \sreg_reg[1414]  ( .D(swire[394]), .CLK(clk), .RST(rst), .Q(sreg[1414])
         );
  DFF \sreg_reg[1415]  ( .D(swire[395]), .CLK(clk), .RST(rst), .Q(sreg[1415])
         );
  DFF \sreg_reg[1416]  ( .D(swire[396]), .CLK(clk), .RST(rst), .Q(sreg[1416])
         );
  DFF \sreg_reg[1417]  ( .D(swire[397]), .CLK(clk), .RST(rst), .Q(sreg[1417])
         );
  DFF \sreg_reg[1418]  ( .D(swire[398]), .CLK(clk), .RST(rst), .Q(sreg[1418])
         );
  DFF \sreg_reg[1419]  ( .D(swire[399]), .CLK(clk), .RST(rst), .Q(sreg[1419])
         );
  DFF \sreg_reg[1420]  ( .D(swire[400]), .CLK(clk), .RST(rst), .Q(sreg[1420])
         );
  DFF \sreg_reg[1421]  ( .D(swire[401]), .CLK(clk), .RST(rst), .Q(sreg[1421])
         );
  DFF \sreg_reg[1422]  ( .D(swire[402]), .CLK(clk), .RST(rst), .Q(sreg[1422])
         );
  DFF \sreg_reg[1423]  ( .D(swire[403]), .CLK(clk), .RST(rst), .Q(sreg[1423])
         );
  DFF \sreg_reg[1424]  ( .D(swire[404]), .CLK(clk), .RST(rst), .Q(sreg[1424])
         );
  DFF \sreg_reg[1425]  ( .D(swire[405]), .CLK(clk), .RST(rst), .Q(sreg[1425])
         );
  DFF \sreg_reg[1426]  ( .D(swire[406]), .CLK(clk), .RST(rst), .Q(sreg[1426])
         );
  DFF \sreg_reg[1427]  ( .D(swire[407]), .CLK(clk), .RST(rst), .Q(sreg[1427])
         );
  DFF \sreg_reg[1428]  ( .D(swire[408]), .CLK(clk), .RST(rst), .Q(sreg[1428])
         );
  DFF \sreg_reg[1429]  ( .D(swire[409]), .CLK(clk), .RST(rst), .Q(sreg[1429])
         );
  DFF \sreg_reg[1430]  ( .D(swire[410]), .CLK(clk), .RST(rst), .Q(sreg[1430])
         );
  DFF \sreg_reg[1431]  ( .D(swire[411]), .CLK(clk), .RST(rst), .Q(sreg[1431])
         );
  DFF \sreg_reg[1432]  ( .D(swire[412]), .CLK(clk), .RST(rst), .Q(sreg[1432])
         );
  DFF \sreg_reg[1433]  ( .D(swire[413]), .CLK(clk), .RST(rst), .Q(sreg[1433])
         );
  DFF \sreg_reg[1434]  ( .D(swire[414]), .CLK(clk), .RST(rst), .Q(sreg[1434])
         );
  DFF \sreg_reg[1435]  ( .D(swire[415]), .CLK(clk), .RST(rst), .Q(sreg[1435])
         );
  DFF \sreg_reg[1436]  ( .D(swire[416]), .CLK(clk), .RST(rst), .Q(sreg[1436])
         );
  DFF \sreg_reg[1437]  ( .D(swire[417]), .CLK(clk), .RST(rst), .Q(sreg[1437])
         );
  DFF \sreg_reg[1438]  ( .D(swire[418]), .CLK(clk), .RST(rst), .Q(sreg[1438])
         );
  DFF \sreg_reg[1439]  ( .D(swire[419]), .CLK(clk), .RST(rst), .Q(sreg[1439])
         );
  DFF \sreg_reg[1440]  ( .D(swire[420]), .CLK(clk), .RST(rst), .Q(sreg[1440])
         );
  DFF \sreg_reg[1441]  ( .D(swire[421]), .CLK(clk), .RST(rst), .Q(sreg[1441])
         );
  DFF \sreg_reg[1442]  ( .D(swire[422]), .CLK(clk), .RST(rst), .Q(sreg[1442])
         );
  DFF \sreg_reg[1443]  ( .D(swire[423]), .CLK(clk), .RST(rst), .Q(sreg[1443])
         );
  DFF \sreg_reg[1444]  ( .D(swire[424]), .CLK(clk), .RST(rst), .Q(sreg[1444])
         );
  DFF \sreg_reg[1445]  ( .D(swire[425]), .CLK(clk), .RST(rst), .Q(sreg[1445])
         );
  DFF \sreg_reg[1446]  ( .D(swire[426]), .CLK(clk), .RST(rst), .Q(sreg[1446])
         );
  DFF \sreg_reg[1447]  ( .D(swire[427]), .CLK(clk), .RST(rst), .Q(sreg[1447])
         );
  DFF \sreg_reg[1448]  ( .D(swire[428]), .CLK(clk), .RST(rst), .Q(sreg[1448])
         );
  DFF \sreg_reg[1449]  ( .D(swire[429]), .CLK(clk), .RST(rst), .Q(sreg[1449])
         );
  DFF \sreg_reg[1450]  ( .D(swire[430]), .CLK(clk), .RST(rst), .Q(sreg[1450])
         );
  DFF \sreg_reg[1451]  ( .D(swire[431]), .CLK(clk), .RST(rst), .Q(sreg[1451])
         );
  DFF \sreg_reg[1452]  ( .D(swire[432]), .CLK(clk), .RST(rst), .Q(sreg[1452])
         );
  DFF \sreg_reg[1453]  ( .D(swire[433]), .CLK(clk), .RST(rst), .Q(sreg[1453])
         );
  DFF \sreg_reg[1454]  ( .D(swire[434]), .CLK(clk), .RST(rst), .Q(sreg[1454])
         );
  DFF \sreg_reg[1455]  ( .D(swire[435]), .CLK(clk), .RST(rst), .Q(sreg[1455])
         );
  DFF \sreg_reg[1456]  ( .D(swire[436]), .CLK(clk), .RST(rst), .Q(sreg[1456])
         );
  DFF \sreg_reg[1457]  ( .D(swire[437]), .CLK(clk), .RST(rst), .Q(sreg[1457])
         );
  DFF \sreg_reg[1458]  ( .D(swire[438]), .CLK(clk), .RST(rst), .Q(sreg[1458])
         );
  DFF \sreg_reg[1459]  ( .D(swire[439]), .CLK(clk), .RST(rst), .Q(sreg[1459])
         );
  DFF \sreg_reg[1460]  ( .D(swire[440]), .CLK(clk), .RST(rst), .Q(sreg[1460])
         );
  DFF \sreg_reg[1461]  ( .D(swire[441]), .CLK(clk), .RST(rst), .Q(sreg[1461])
         );
  DFF \sreg_reg[1462]  ( .D(swire[442]), .CLK(clk), .RST(rst), .Q(sreg[1462])
         );
  DFF \sreg_reg[1463]  ( .D(swire[443]), .CLK(clk), .RST(rst), .Q(sreg[1463])
         );
  DFF \sreg_reg[1464]  ( .D(swire[444]), .CLK(clk), .RST(rst), .Q(sreg[1464])
         );
  DFF \sreg_reg[1465]  ( .D(swire[445]), .CLK(clk), .RST(rst), .Q(sreg[1465])
         );
  DFF \sreg_reg[1466]  ( .D(swire[446]), .CLK(clk), .RST(rst), .Q(sreg[1466])
         );
  DFF \sreg_reg[1467]  ( .D(swire[447]), .CLK(clk), .RST(rst), .Q(sreg[1467])
         );
  DFF \sreg_reg[1468]  ( .D(swire[448]), .CLK(clk), .RST(rst), .Q(sreg[1468])
         );
  DFF \sreg_reg[1469]  ( .D(swire[449]), .CLK(clk), .RST(rst), .Q(sreg[1469])
         );
  DFF \sreg_reg[1470]  ( .D(swire[450]), .CLK(clk), .RST(rst), .Q(sreg[1470])
         );
  DFF \sreg_reg[1471]  ( .D(swire[451]), .CLK(clk), .RST(rst), .Q(sreg[1471])
         );
  DFF \sreg_reg[1472]  ( .D(swire[452]), .CLK(clk), .RST(rst), .Q(sreg[1472])
         );
  DFF \sreg_reg[1473]  ( .D(swire[453]), .CLK(clk), .RST(rst), .Q(sreg[1473])
         );
  DFF \sreg_reg[1474]  ( .D(swire[454]), .CLK(clk), .RST(rst), .Q(sreg[1474])
         );
  DFF \sreg_reg[1475]  ( .D(swire[455]), .CLK(clk), .RST(rst), .Q(sreg[1475])
         );
  DFF \sreg_reg[1476]  ( .D(swire[456]), .CLK(clk), .RST(rst), .Q(sreg[1476])
         );
  DFF \sreg_reg[1477]  ( .D(swire[457]), .CLK(clk), .RST(rst), .Q(sreg[1477])
         );
  DFF \sreg_reg[1478]  ( .D(swire[458]), .CLK(clk), .RST(rst), .Q(sreg[1478])
         );
  DFF \sreg_reg[1479]  ( .D(swire[459]), .CLK(clk), .RST(rst), .Q(sreg[1479])
         );
  DFF \sreg_reg[1480]  ( .D(swire[460]), .CLK(clk), .RST(rst), .Q(sreg[1480])
         );
  DFF \sreg_reg[1481]  ( .D(swire[461]), .CLK(clk), .RST(rst), .Q(sreg[1481])
         );
  DFF \sreg_reg[1482]  ( .D(swire[462]), .CLK(clk), .RST(rst), .Q(sreg[1482])
         );
  DFF \sreg_reg[1483]  ( .D(swire[463]), .CLK(clk), .RST(rst), .Q(sreg[1483])
         );
  DFF \sreg_reg[1484]  ( .D(swire[464]), .CLK(clk), .RST(rst), .Q(sreg[1484])
         );
  DFF \sreg_reg[1485]  ( .D(swire[465]), .CLK(clk), .RST(rst), .Q(sreg[1485])
         );
  DFF \sreg_reg[1486]  ( .D(swire[466]), .CLK(clk), .RST(rst), .Q(sreg[1486])
         );
  DFF \sreg_reg[1487]  ( .D(swire[467]), .CLK(clk), .RST(rst), .Q(sreg[1487])
         );
  DFF \sreg_reg[1488]  ( .D(swire[468]), .CLK(clk), .RST(rst), .Q(sreg[1488])
         );
  DFF \sreg_reg[1489]  ( .D(swire[469]), .CLK(clk), .RST(rst), .Q(sreg[1489])
         );
  DFF \sreg_reg[1490]  ( .D(swire[470]), .CLK(clk), .RST(rst), .Q(sreg[1490])
         );
  DFF \sreg_reg[1491]  ( .D(swire[471]), .CLK(clk), .RST(rst), .Q(sreg[1491])
         );
  DFF \sreg_reg[1492]  ( .D(swire[472]), .CLK(clk), .RST(rst), .Q(sreg[1492])
         );
  DFF \sreg_reg[1493]  ( .D(swire[473]), .CLK(clk), .RST(rst), .Q(sreg[1493])
         );
  DFF \sreg_reg[1494]  ( .D(swire[474]), .CLK(clk), .RST(rst), .Q(sreg[1494])
         );
  DFF \sreg_reg[1495]  ( .D(swire[475]), .CLK(clk), .RST(rst), .Q(sreg[1495])
         );
  DFF \sreg_reg[1496]  ( .D(swire[476]), .CLK(clk), .RST(rst), .Q(sreg[1496])
         );
  DFF \sreg_reg[1497]  ( .D(swire[477]), .CLK(clk), .RST(rst), .Q(sreg[1497])
         );
  DFF \sreg_reg[1498]  ( .D(swire[478]), .CLK(clk), .RST(rst), .Q(sreg[1498])
         );
  DFF \sreg_reg[1499]  ( .D(swire[479]), .CLK(clk), .RST(rst), .Q(sreg[1499])
         );
  DFF \sreg_reg[1500]  ( .D(swire[480]), .CLK(clk), .RST(rst), .Q(sreg[1500])
         );
  DFF \sreg_reg[1501]  ( .D(swire[481]), .CLK(clk), .RST(rst), .Q(sreg[1501])
         );
  DFF \sreg_reg[1502]  ( .D(swire[482]), .CLK(clk), .RST(rst), .Q(sreg[1502])
         );
  DFF \sreg_reg[1503]  ( .D(swire[483]), .CLK(clk), .RST(rst), .Q(sreg[1503])
         );
  DFF \sreg_reg[1504]  ( .D(swire[484]), .CLK(clk), .RST(rst), .Q(sreg[1504])
         );
  DFF \sreg_reg[1505]  ( .D(swire[485]), .CLK(clk), .RST(rst), .Q(sreg[1505])
         );
  DFF \sreg_reg[1506]  ( .D(swire[486]), .CLK(clk), .RST(rst), .Q(sreg[1506])
         );
  DFF \sreg_reg[1507]  ( .D(swire[487]), .CLK(clk), .RST(rst), .Q(sreg[1507])
         );
  DFF \sreg_reg[1508]  ( .D(swire[488]), .CLK(clk), .RST(rst), .Q(sreg[1508])
         );
  DFF \sreg_reg[1509]  ( .D(swire[489]), .CLK(clk), .RST(rst), .Q(sreg[1509])
         );
  DFF \sreg_reg[1510]  ( .D(swire[490]), .CLK(clk), .RST(rst), .Q(sreg[1510])
         );
  DFF \sreg_reg[1511]  ( .D(swire[491]), .CLK(clk), .RST(rst), .Q(sreg[1511])
         );
  DFF \sreg_reg[1512]  ( .D(swire[492]), .CLK(clk), .RST(rst), .Q(sreg[1512])
         );
  DFF \sreg_reg[1513]  ( .D(swire[493]), .CLK(clk), .RST(rst), .Q(sreg[1513])
         );
  DFF \sreg_reg[1514]  ( .D(swire[494]), .CLK(clk), .RST(rst), .Q(sreg[1514])
         );
  DFF \sreg_reg[1515]  ( .D(swire[495]), .CLK(clk), .RST(rst), .Q(sreg[1515])
         );
  DFF \sreg_reg[1516]  ( .D(swire[496]), .CLK(clk), .RST(rst), .Q(sreg[1516])
         );
  DFF \sreg_reg[1517]  ( .D(swire[497]), .CLK(clk), .RST(rst), .Q(sreg[1517])
         );
  DFF \sreg_reg[1518]  ( .D(swire[498]), .CLK(clk), .RST(rst), .Q(sreg[1518])
         );
  DFF \sreg_reg[1519]  ( .D(swire[499]), .CLK(clk), .RST(rst), .Q(sreg[1519])
         );
  DFF \sreg_reg[1520]  ( .D(swire[500]), .CLK(clk), .RST(rst), .Q(sreg[1520])
         );
  DFF \sreg_reg[1521]  ( .D(swire[501]), .CLK(clk), .RST(rst), .Q(sreg[1521])
         );
  DFF \sreg_reg[1522]  ( .D(swire[502]), .CLK(clk), .RST(rst), .Q(sreg[1522])
         );
  DFF \sreg_reg[1523]  ( .D(swire[503]), .CLK(clk), .RST(rst), .Q(sreg[1523])
         );
  DFF \sreg_reg[1524]  ( .D(swire[504]), .CLK(clk), .RST(rst), .Q(sreg[1524])
         );
  DFF \sreg_reg[1525]  ( .D(swire[505]), .CLK(clk), .RST(rst), .Q(sreg[1525])
         );
  DFF \sreg_reg[1526]  ( .D(swire[506]), .CLK(clk), .RST(rst), .Q(sreg[1526])
         );
  DFF \sreg_reg[1527]  ( .D(swire[507]), .CLK(clk), .RST(rst), .Q(sreg[1527])
         );
  DFF \sreg_reg[1528]  ( .D(swire[508]), .CLK(clk), .RST(rst), .Q(sreg[1528])
         );
  DFF \sreg_reg[1529]  ( .D(swire[509]), .CLK(clk), .RST(rst), .Q(sreg[1529])
         );
  DFF \sreg_reg[1530]  ( .D(swire[510]), .CLK(clk), .RST(rst), .Q(sreg[1530])
         );
  DFF \sreg_reg[1531]  ( .D(swire[511]), .CLK(clk), .RST(rst), .Q(sreg[1531])
         );
  DFF \sreg_reg[1532]  ( .D(swire[512]), .CLK(clk), .RST(rst), .Q(sreg[1532])
         );
  DFF \sreg_reg[1533]  ( .D(swire[513]), .CLK(clk), .RST(rst), .Q(sreg[1533])
         );
  DFF \sreg_reg[1534]  ( .D(swire[514]), .CLK(clk), .RST(rst), .Q(sreg[1534])
         );
  DFF \sreg_reg[1535]  ( .D(swire[515]), .CLK(clk), .RST(rst), .Q(sreg[1535])
         );
  DFF \sreg_reg[1536]  ( .D(swire[516]), .CLK(clk), .RST(rst), .Q(sreg[1536])
         );
  DFF \sreg_reg[1537]  ( .D(swire[517]), .CLK(clk), .RST(rst), .Q(sreg[1537])
         );
  DFF \sreg_reg[1538]  ( .D(swire[518]), .CLK(clk), .RST(rst), .Q(sreg[1538])
         );
  DFF \sreg_reg[1539]  ( .D(swire[519]), .CLK(clk), .RST(rst), .Q(sreg[1539])
         );
  DFF \sreg_reg[1540]  ( .D(swire[520]), .CLK(clk), .RST(rst), .Q(sreg[1540])
         );
  DFF \sreg_reg[1541]  ( .D(swire[521]), .CLK(clk), .RST(rst), .Q(sreg[1541])
         );
  DFF \sreg_reg[1542]  ( .D(swire[522]), .CLK(clk), .RST(rst), .Q(sreg[1542])
         );
  DFF \sreg_reg[1543]  ( .D(swire[523]), .CLK(clk), .RST(rst), .Q(sreg[1543])
         );
  DFF \sreg_reg[1544]  ( .D(swire[524]), .CLK(clk), .RST(rst), .Q(sreg[1544])
         );
  DFF \sreg_reg[1545]  ( .D(swire[525]), .CLK(clk), .RST(rst), .Q(sreg[1545])
         );
  DFF \sreg_reg[1546]  ( .D(swire[526]), .CLK(clk), .RST(rst), .Q(sreg[1546])
         );
  DFF \sreg_reg[1547]  ( .D(swire[527]), .CLK(clk), .RST(rst), .Q(sreg[1547])
         );
  DFF \sreg_reg[1548]  ( .D(swire[528]), .CLK(clk), .RST(rst), .Q(sreg[1548])
         );
  DFF \sreg_reg[1549]  ( .D(swire[529]), .CLK(clk), .RST(rst), .Q(sreg[1549])
         );
  DFF \sreg_reg[1550]  ( .D(swire[530]), .CLK(clk), .RST(rst), .Q(sreg[1550])
         );
  DFF \sreg_reg[1551]  ( .D(swire[531]), .CLK(clk), .RST(rst), .Q(sreg[1551])
         );
  DFF \sreg_reg[1552]  ( .D(swire[532]), .CLK(clk), .RST(rst), .Q(sreg[1552])
         );
  DFF \sreg_reg[1553]  ( .D(swire[533]), .CLK(clk), .RST(rst), .Q(sreg[1553])
         );
  DFF \sreg_reg[1554]  ( .D(swire[534]), .CLK(clk), .RST(rst), .Q(sreg[1554])
         );
  DFF \sreg_reg[1555]  ( .D(swire[535]), .CLK(clk), .RST(rst), .Q(sreg[1555])
         );
  DFF \sreg_reg[1556]  ( .D(swire[536]), .CLK(clk), .RST(rst), .Q(sreg[1556])
         );
  DFF \sreg_reg[1557]  ( .D(swire[537]), .CLK(clk), .RST(rst), .Q(sreg[1557])
         );
  DFF \sreg_reg[1558]  ( .D(swire[538]), .CLK(clk), .RST(rst), .Q(sreg[1558])
         );
  DFF \sreg_reg[1559]  ( .D(swire[539]), .CLK(clk), .RST(rst), .Q(sreg[1559])
         );
  DFF \sreg_reg[1560]  ( .D(swire[540]), .CLK(clk), .RST(rst), .Q(sreg[1560])
         );
  DFF \sreg_reg[1561]  ( .D(swire[541]), .CLK(clk), .RST(rst), .Q(sreg[1561])
         );
  DFF \sreg_reg[1562]  ( .D(swire[542]), .CLK(clk), .RST(rst), .Q(sreg[1562])
         );
  DFF \sreg_reg[1563]  ( .D(swire[543]), .CLK(clk), .RST(rst), .Q(sreg[1563])
         );
  DFF \sreg_reg[1564]  ( .D(swire[544]), .CLK(clk), .RST(rst), .Q(sreg[1564])
         );
  DFF \sreg_reg[1565]  ( .D(swire[545]), .CLK(clk), .RST(rst), .Q(sreg[1565])
         );
  DFF \sreg_reg[1566]  ( .D(swire[546]), .CLK(clk), .RST(rst), .Q(sreg[1566])
         );
  DFF \sreg_reg[1567]  ( .D(swire[547]), .CLK(clk), .RST(rst), .Q(sreg[1567])
         );
  DFF \sreg_reg[1568]  ( .D(swire[548]), .CLK(clk), .RST(rst), .Q(sreg[1568])
         );
  DFF \sreg_reg[1569]  ( .D(swire[549]), .CLK(clk), .RST(rst), .Q(sreg[1569])
         );
  DFF \sreg_reg[1570]  ( .D(swire[550]), .CLK(clk), .RST(rst), .Q(sreg[1570])
         );
  DFF \sreg_reg[1571]  ( .D(swire[551]), .CLK(clk), .RST(rst), .Q(sreg[1571])
         );
  DFF \sreg_reg[1572]  ( .D(swire[552]), .CLK(clk), .RST(rst), .Q(sreg[1572])
         );
  DFF \sreg_reg[1573]  ( .D(swire[553]), .CLK(clk), .RST(rst), .Q(sreg[1573])
         );
  DFF \sreg_reg[1574]  ( .D(swire[554]), .CLK(clk), .RST(rst), .Q(sreg[1574])
         );
  DFF \sreg_reg[1575]  ( .D(swire[555]), .CLK(clk), .RST(rst), .Q(sreg[1575])
         );
  DFF \sreg_reg[1576]  ( .D(swire[556]), .CLK(clk), .RST(rst), .Q(sreg[1576])
         );
  DFF \sreg_reg[1577]  ( .D(swire[557]), .CLK(clk), .RST(rst), .Q(sreg[1577])
         );
  DFF \sreg_reg[1578]  ( .D(swire[558]), .CLK(clk), .RST(rst), .Q(sreg[1578])
         );
  DFF \sreg_reg[1579]  ( .D(swire[559]), .CLK(clk), .RST(rst), .Q(sreg[1579])
         );
  DFF \sreg_reg[1580]  ( .D(swire[560]), .CLK(clk), .RST(rst), .Q(sreg[1580])
         );
  DFF \sreg_reg[1581]  ( .D(swire[561]), .CLK(clk), .RST(rst), .Q(sreg[1581])
         );
  DFF \sreg_reg[1582]  ( .D(swire[562]), .CLK(clk), .RST(rst), .Q(sreg[1582])
         );
  DFF \sreg_reg[1583]  ( .D(swire[563]), .CLK(clk), .RST(rst), .Q(sreg[1583])
         );
  DFF \sreg_reg[1584]  ( .D(swire[564]), .CLK(clk), .RST(rst), .Q(sreg[1584])
         );
  DFF \sreg_reg[1585]  ( .D(swire[565]), .CLK(clk), .RST(rst), .Q(sreg[1585])
         );
  DFF \sreg_reg[1586]  ( .D(swire[566]), .CLK(clk), .RST(rst), .Q(sreg[1586])
         );
  DFF \sreg_reg[1587]  ( .D(swire[567]), .CLK(clk), .RST(rst), .Q(sreg[1587])
         );
  DFF \sreg_reg[1588]  ( .D(swire[568]), .CLK(clk), .RST(rst), .Q(sreg[1588])
         );
  DFF \sreg_reg[1589]  ( .D(swire[569]), .CLK(clk), .RST(rst), .Q(sreg[1589])
         );
  DFF \sreg_reg[1590]  ( .D(swire[570]), .CLK(clk), .RST(rst), .Q(sreg[1590])
         );
  DFF \sreg_reg[1591]  ( .D(swire[571]), .CLK(clk), .RST(rst), .Q(sreg[1591])
         );
  DFF \sreg_reg[1592]  ( .D(swire[572]), .CLK(clk), .RST(rst), .Q(sreg[1592])
         );
  DFF \sreg_reg[1593]  ( .D(swire[573]), .CLK(clk), .RST(rst), .Q(sreg[1593])
         );
  DFF \sreg_reg[1594]  ( .D(swire[574]), .CLK(clk), .RST(rst), .Q(sreg[1594])
         );
  DFF \sreg_reg[1595]  ( .D(swire[575]), .CLK(clk), .RST(rst), .Q(sreg[1595])
         );
  DFF \sreg_reg[1596]  ( .D(swire[576]), .CLK(clk), .RST(rst), .Q(sreg[1596])
         );
  DFF \sreg_reg[1597]  ( .D(swire[577]), .CLK(clk), .RST(rst), .Q(sreg[1597])
         );
  DFF \sreg_reg[1598]  ( .D(swire[578]), .CLK(clk), .RST(rst), .Q(sreg[1598])
         );
  DFF \sreg_reg[1599]  ( .D(swire[579]), .CLK(clk), .RST(rst), .Q(sreg[1599])
         );
  DFF \sreg_reg[1600]  ( .D(swire[580]), .CLK(clk), .RST(rst), .Q(sreg[1600])
         );
  DFF \sreg_reg[1601]  ( .D(swire[581]), .CLK(clk), .RST(rst), .Q(sreg[1601])
         );
  DFF \sreg_reg[1602]  ( .D(swire[582]), .CLK(clk), .RST(rst), .Q(sreg[1602])
         );
  DFF \sreg_reg[1603]  ( .D(swire[583]), .CLK(clk), .RST(rst), .Q(sreg[1603])
         );
  DFF \sreg_reg[1604]  ( .D(swire[584]), .CLK(clk), .RST(rst), .Q(sreg[1604])
         );
  DFF \sreg_reg[1605]  ( .D(swire[585]), .CLK(clk), .RST(rst), .Q(sreg[1605])
         );
  DFF \sreg_reg[1606]  ( .D(swire[586]), .CLK(clk), .RST(rst), .Q(sreg[1606])
         );
  DFF \sreg_reg[1607]  ( .D(swire[587]), .CLK(clk), .RST(rst), .Q(sreg[1607])
         );
  DFF \sreg_reg[1608]  ( .D(swire[588]), .CLK(clk), .RST(rst), .Q(sreg[1608])
         );
  DFF \sreg_reg[1609]  ( .D(swire[589]), .CLK(clk), .RST(rst), .Q(sreg[1609])
         );
  DFF \sreg_reg[1610]  ( .D(swire[590]), .CLK(clk), .RST(rst), .Q(sreg[1610])
         );
  DFF \sreg_reg[1611]  ( .D(swire[591]), .CLK(clk), .RST(rst), .Q(sreg[1611])
         );
  DFF \sreg_reg[1612]  ( .D(swire[592]), .CLK(clk), .RST(rst), .Q(sreg[1612])
         );
  DFF \sreg_reg[1613]  ( .D(swire[593]), .CLK(clk), .RST(rst), .Q(sreg[1613])
         );
  DFF \sreg_reg[1614]  ( .D(swire[594]), .CLK(clk), .RST(rst), .Q(sreg[1614])
         );
  DFF \sreg_reg[1615]  ( .D(swire[595]), .CLK(clk), .RST(rst), .Q(sreg[1615])
         );
  DFF \sreg_reg[1616]  ( .D(swire[596]), .CLK(clk), .RST(rst), .Q(sreg[1616])
         );
  DFF \sreg_reg[1617]  ( .D(swire[597]), .CLK(clk), .RST(rst), .Q(sreg[1617])
         );
  DFF \sreg_reg[1618]  ( .D(swire[598]), .CLK(clk), .RST(rst), .Q(sreg[1618])
         );
  DFF \sreg_reg[1619]  ( .D(swire[599]), .CLK(clk), .RST(rst), .Q(sreg[1619])
         );
  DFF \sreg_reg[1620]  ( .D(swire[600]), .CLK(clk), .RST(rst), .Q(sreg[1620])
         );
  DFF \sreg_reg[1621]  ( .D(swire[601]), .CLK(clk), .RST(rst), .Q(sreg[1621])
         );
  DFF \sreg_reg[1622]  ( .D(swire[602]), .CLK(clk), .RST(rst), .Q(sreg[1622])
         );
  DFF \sreg_reg[1623]  ( .D(swire[603]), .CLK(clk), .RST(rst), .Q(sreg[1623])
         );
  DFF \sreg_reg[1624]  ( .D(swire[604]), .CLK(clk), .RST(rst), .Q(sreg[1624])
         );
  DFF \sreg_reg[1625]  ( .D(swire[605]), .CLK(clk), .RST(rst), .Q(sreg[1625])
         );
  DFF \sreg_reg[1626]  ( .D(swire[606]), .CLK(clk), .RST(rst), .Q(sreg[1626])
         );
  DFF \sreg_reg[1627]  ( .D(swire[607]), .CLK(clk), .RST(rst), .Q(sreg[1627])
         );
  DFF \sreg_reg[1628]  ( .D(swire[608]), .CLK(clk), .RST(rst), .Q(sreg[1628])
         );
  DFF \sreg_reg[1629]  ( .D(swire[609]), .CLK(clk), .RST(rst), .Q(sreg[1629])
         );
  DFF \sreg_reg[1630]  ( .D(swire[610]), .CLK(clk), .RST(rst), .Q(sreg[1630])
         );
  DFF \sreg_reg[1631]  ( .D(swire[611]), .CLK(clk), .RST(rst), .Q(sreg[1631])
         );
  DFF \sreg_reg[1632]  ( .D(swire[612]), .CLK(clk), .RST(rst), .Q(sreg[1632])
         );
  DFF \sreg_reg[1633]  ( .D(swire[613]), .CLK(clk), .RST(rst), .Q(sreg[1633])
         );
  DFF \sreg_reg[1634]  ( .D(swire[614]), .CLK(clk), .RST(rst), .Q(sreg[1634])
         );
  DFF \sreg_reg[1635]  ( .D(swire[615]), .CLK(clk), .RST(rst), .Q(sreg[1635])
         );
  DFF \sreg_reg[1636]  ( .D(swire[616]), .CLK(clk), .RST(rst), .Q(sreg[1636])
         );
  DFF \sreg_reg[1637]  ( .D(swire[617]), .CLK(clk), .RST(rst), .Q(sreg[1637])
         );
  DFF \sreg_reg[1638]  ( .D(swire[618]), .CLK(clk), .RST(rst), .Q(sreg[1638])
         );
  DFF \sreg_reg[1639]  ( .D(swire[619]), .CLK(clk), .RST(rst), .Q(sreg[1639])
         );
  DFF \sreg_reg[1640]  ( .D(swire[620]), .CLK(clk), .RST(rst), .Q(sreg[1640])
         );
  DFF \sreg_reg[1641]  ( .D(swire[621]), .CLK(clk), .RST(rst), .Q(sreg[1641])
         );
  DFF \sreg_reg[1642]  ( .D(swire[622]), .CLK(clk), .RST(rst), .Q(sreg[1642])
         );
  DFF \sreg_reg[1643]  ( .D(swire[623]), .CLK(clk), .RST(rst), .Q(sreg[1643])
         );
  DFF \sreg_reg[1644]  ( .D(swire[624]), .CLK(clk), .RST(rst), .Q(sreg[1644])
         );
  DFF \sreg_reg[1645]  ( .D(swire[625]), .CLK(clk), .RST(rst), .Q(sreg[1645])
         );
  DFF \sreg_reg[1646]  ( .D(swire[626]), .CLK(clk), .RST(rst), .Q(sreg[1646])
         );
  DFF \sreg_reg[1647]  ( .D(swire[627]), .CLK(clk), .RST(rst), .Q(sreg[1647])
         );
  DFF \sreg_reg[1648]  ( .D(swire[628]), .CLK(clk), .RST(rst), .Q(sreg[1648])
         );
  DFF \sreg_reg[1649]  ( .D(swire[629]), .CLK(clk), .RST(rst), .Q(sreg[1649])
         );
  DFF \sreg_reg[1650]  ( .D(swire[630]), .CLK(clk), .RST(rst), .Q(sreg[1650])
         );
  DFF \sreg_reg[1651]  ( .D(swire[631]), .CLK(clk), .RST(rst), .Q(sreg[1651])
         );
  DFF \sreg_reg[1652]  ( .D(swire[632]), .CLK(clk), .RST(rst), .Q(sreg[1652])
         );
  DFF \sreg_reg[1653]  ( .D(swire[633]), .CLK(clk), .RST(rst), .Q(sreg[1653])
         );
  DFF \sreg_reg[1654]  ( .D(swire[634]), .CLK(clk), .RST(rst), .Q(sreg[1654])
         );
  DFF \sreg_reg[1655]  ( .D(swire[635]), .CLK(clk), .RST(rst), .Q(sreg[1655])
         );
  DFF \sreg_reg[1656]  ( .D(swire[636]), .CLK(clk), .RST(rst), .Q(sreg[1656])
         );
  DFF \sreg_reg[1657]  ( .D(swire[637]), .CLK(clk), .RST(rst), .Q(sreg[1657])
         );
  DFF \sreg_reg[1658]  ( .D(swire[638]), .CLK(clk), .RST(rst), .Q(sreg[1658])
         );
  DFF \sreg_reg[1659]  ( .D(swire[639]), .CLK(clk), .RST(rst), .Q(sreg[1659])
         );
  DFF \sreg_reg[1660]  ( .D(swire[640]), .CLK(clk), .RST(rst), .Q(sreg[1660])
         );
  DFF \sreg_reg[1661]  ( .D(swire[641]), .CLK(clk), .RST(rst), .Q(sreg[1661])
         );
  DFF \sreg_reg[1662]  ( .D(swire[642]), .CLK(clk), .RST(rst), .Q(sreg[1662])
         );
  DFF \sreg_reg[1663]  ( .D(swire[643]), .CLK(clk), .RST(rst), .Q(sreg[1663])
         );
  DFF \sreg_reg[1664]  ( .D(swire[644]), .CLK(clk), .RST(rst), .Q(sreg[1664])
         );
  DFF \sreg_reg[1665]  ( .D(swire[645]), .CLK(clk), .RST(rst), .Q(sreg[1665])
         );
  DFF \sreg_reg[1666]  ( .D(swire[646]), .CLK(clk), .RST(rst), .Q(sreg[1666])
         );
  DFF \sreg_reg[1667]  ( .D(swire[647]), .CLK(clk), .RST(rst), .Q(sreg[1667])
         );
  DFF \sreg_reg[1668]  ( .D(swire[648]), .CLK(clk), .RST(rst), .Q(sreg[1668])
         );
  DFF \sreg_reg[1669]  ( .D(swire[649]), .CLK(clk), .RST(rst), .Q(sreg[1669])
         );
  DFF \sreg_reg[1670]  ( .D(swire[650]), .CLK(clk), .RST(rst), .Q(sreg[1670])
         );
  DFF \sreg_reg[1671]  ( .D(swire[651]), .CLK(clk), .RST(rst), .Q(sreg[1671])
         );
  DFF \sreg_reg[1672]  ( .D(swire[652]), .CLK(clk), .RST(rst), .Q(sreg[1672])
         );
  DFF \sreg_reg[1673]  ( .D(swire[653]), .CLK(clk), .RST(rst), .Q(sreg[1673])
         );
  DFF \sreg_reg[1674]  ( .D(swire[654]), .CLK(clk), .RST(rst), .Q(sreg[1674])
         );
  DFF \sreg_reg[1675]  ( .D(swire[655]), .CLK(clk), .RST(rst), .Q(sreg[1675])
         );
  DFF \sreg_reg[1676]  ( .D(swire[656]), .CLK(clk), .RST(rst), .Q(sreg[1676])
         );
  DFF \sreg_reg[1677]  ( .D(swire[657]), .CLK(clk), .RST(rst), .Q(sreg[1677])
         );
  DFF \sreg_reg[1678]  ( .D(swire[658]), .CLK(clk), .RST(rst), .Q(sreg[1678])
         );
  DFF \sreg_reg[1679]  ( .D(swire[659]), .CLK(clk), .RST(rst), .Q(sreg[1679])
         );
  DFF \sreg_reg[1680]  ( .D(swire[660]), .CLK(clk), .RST(rst), .Q(sreg[1680])
         );
  DFF \sreg_reg[1681]  ( .D(swire[661]), .CLK(clk), .RST(rst), .Q(sreg[1681])
         );
  DFF \sreg_reg[1682]  ( .D(swire[662]), .CLK(clk), .RST(rst), .Q(sreg[1682])
         );
  DFF \sreg_reg[1683]  ( .D(swire[663]), .CLK(clk), .RST(rst), .Q(sreg[1683])
         );
  DFF \sreg_reg[1684]  ( .D(swire[664]), .CLK(clk), .RST(rst), .Q(sreg[1684])
         );
  DFF \sreg_reg[1685]  ( .D(swire[665]), .CLK(clk), .RST(rst), .Q(sreg[1685])
         );
  DFF \sreg_reg[1686]  ( .D(swire[666]), .CLK(clk), .RST(rst), .Q(sreg[1686])
         );
  DFF \sreg_reg[1687]  ( .D(swire[667]), .CLK(clk), .RST(rst), .Q(sreg[1687])
         );
  DFF \sreg_reg[1688]  ( .D(swire[668]), .CLK(clk), .RST(rst), .Q(sreg[1688])
         );
  DFF \sreg_reg[1689]  ( .D(swire[669]), .CLK(clk), .RST(rst), .Q(sreg[1689])
         );
  DFF \sreg_reg[1690]  ( .D(swire[670]), .CLK(clk), .RST(rst), .Q(sreg[1690])
         );
  DFF \sreg_reg[1691]  ( .D(swire[671]), .CLK(clk), .RST(rst), .Q(sreg[1691])
         );
  DFF \sreg_reg[1692]  ( .D(swire[672]), .CLK(clk), .RST(rst), .Q(sreg[1692])
         );
  DFF \sreg_reg[1693]  ( .D(swire[673]), .CLK(clk), .RST(rst), .Q(sreg[1693])
         );
  DFF \sreg_reg[1694]  ( .D(swire[674]), .CLK(clk), .RST(rst), .Q(sreg[1694])
         );
  DFF \sreg_reg[1695]  ( .D(swire[675]), .CLK(clk), .RST(rst), .Q(sreg[1695])
         );
  DFF \sreg_reg[1696]  ( .D(swire[676]), .CLK(clk), .RST(rst), .Q(sreg[1696])
         );
  DFF \sreg_reg[1697]  ( .D(swire[677]), .CLK(clk), .RST(rst), .Q(sreg[1697])
         );
  DFF \sreg_reg[1698]  ( .D(swire[678]), .CLK(clk), .RST(rst), .Q(sreg[1698])
         );
  DFF \sreg_reg[1699]  ( .D(swire[679]), .CLK(clk), .RST(rst), .Q(sreg[1699])
         );
  DFF \sreg_reg[1700]  ( .D(swire[680]), .CLK(clk), .RST(rst), .Q(sreg[1700])
         );
  DFF \sreg_reg[1701]  ( .D(swire[681]), .CLK(clk), .RST(rst), .Q(sreg[1701])
         );
  DFF \sreg_reg[1702]  ( .D(swire[682]), .CLK(clk), .RST(rst), .Q(sreg[1702])
         );
  DFF \sreg_reg[1703]  ( .D(swire[683]), .CLK(clk), .RST(rst), .Q(sreg[1703])
         );
  DFF \sreg_reg[1704]  ( .D(swire[684]), .CLK(clk), .RST(rst), .Q(sreg[1704])
         );
  DFF \sreg_reg[1705]  ( .D(swire[685]), .CLK(clk), .RST(rst), .Q(sreg[1705])
         );
  DFF \sreg_reg[1706]  ( .D(swire[686]), .CLK(clk), .RST(rst), .Q(sreg[1706])
         );
  DFF \sreg_reg[1707]  ( .D(swire[687]), .CLK(clk), .RST(rst), .Q(sreg[1707])
         );
  DFF \sreg_reg[1708]  ( .D(swire[688]), .CLK(clk), .RST(rst), .Q(sreg[1708])
         );
  DFF \sreg_reg[1709]  ( .D(swire[689]), .CLK(clk), .RST(rst), .Q(sreg[1709])
         );
  DFF \sreg_reg[1710]  ( .D(swire[690]), .CLK(clk), .RST(rst), .Q(sreg[1710])
         );
  DFF \sreg_reg[1711]  ( .D(swire[691]), .CLK(clk), .RST(rst), .Q(sreg[1711])
         );
  DFF \sreg_reg[1712]  ( .D(swire[692]), .CLK(clk), .RST(rst), .Q(sreg[1712])
         );
  DFF \sreg_reg[1713]  ( .D(swire[693]), .CLK(clk), .RST(rst), .Q(sreg[1713])
         );
  DFF \sreg_reg[1714]  ( .D(swire[694]), .CLK(clk), .RST(rst), .Q(sreg[1714])
         );
  DFF \sreg_reg[1715]  ( .D(swire[695]), .CLK(clk), .RST(rst), .Q(sreg[1715])
         );
  DFF \sreg_reg[1716]  ( .D(swire[696]), .CLK(clk), .RST(rst), .Q(sreg[1716])
         );
  DFF \sreg_reg[1717]  ( .D(swire[697]), .CLK(clk), .RST(rst), .Q(sreg[1717])
         );
  DFF \sreg_reg[1718]  ( .D(swire[698]), .CLK(clk), .RST(rst), .Q(sreg[1718])
         );
  DFF \sreg_reg[1719]  ( .D(swire[699]), .CLK(clk), .RST(rst), .Q(sreg[1719])
         );
  DFF \sreg_reg[1720]  ( .D(swire[700]), .CLK(clk), .RST(rst), .Q(sreg[1720])
         );
  DFF \sreg_reg[1721]  ( .D(swire[701]), .CLK(clk), .RST(rst), .Q(sreg[1721])
         );
  DFF \sreg_reg[1722]  ( .D(swire[702]), .CLK(clk), .RST(rst), .Q(sreg[1722])
         );
  DFF \sreg_reg[1723]  ( .D(swire[703]), .CLK(clk), .RST(rst), .Q(sreg[1723])
         );
  DFF \sreg_reg[1724]  ( .D(swire[704]), .CLK(clk), .RST(rst), .Q(sreg[1724])
         );
  DFF \sreg_reg[1725]  ( .D(swire[705]), .CLK(clk), .RST(rst), .Q(sreg[1725])
         );
  DFF \sreg_reg[1726]  ( .D(swire[706]), .CLK(clk), .RST(rst), .Q(sreg[1726])
         );
  DFF \sreg_reg[1727]  ( .D(swire[707]), .CLK(clk), .RST(rst), .Q(sreg[1727])
         );
  DFF \sreg_reg[1728]  ( .D(swire[708]), .CLK(clk), .RST(rst), .Q(sreg[1728])
         );
  DFF \sreg_reg[1729]  ( .D(swire[709]), .CLK(clk), .RST(rst), .Q(sreg[1729])
         );
  DFF \sreg_reg[1730]  ( .D(swire[710]), .CLK(clk), .RST(rst), .Q(sreg[1730])
         );
  DFF \sreg_reg[1731]  ( .D(swire[711]), .CLK(clk), .RST(rst), .Q(sreg[1731])
         );
  DFF \sreg_reg[1732]  ( .D(swire[712]), .CLK(clk), .RST(rst), .Q(sreg[1732])
         );
  DFF \sreg_reg[1733]  ( .D(swire[713]), .CLK(clk), .RST(rst), .Q(sreg[1733])
         );
  DFF \sreg_reg[1734]  ( .D(swire[714]), .CLK(clk), .RST(rst), .Q(sreg[1734])
         );
  DFF \sreg_reg[1735]  ( .D(swire[715]), .CLK(clk), .RST(rst), .Q(sreg[1735])
         );
  DFF \sreg_reg[1736]  ( .D(swire[716]), .CLK(clk), .RST(rst), .Q(sreg[1736])
         );
  DFF \sreg_reg[1737]  ( .D(swire[717]), .CLK(clk), .RST(rst), .Q(sreg[1737])
         );
  DFF \sreg_reg[1738]  ( .D(swire[718]), .CLK(clk), .RST(rst), .Q(sreg[1738])
         );
  DFF \sreg_reg[1739]  ( .D(swire[719]), .CLK(clk), .RST(rst), .Q(sreg[1739])
         );
  DFF \sreg_reg[1740]  ( .D(swire[720]), .CLK(clk), .RST(rst), .Q(sreg[1740])
         );
  DFF \sreg_reg[1741]  ( .D(swire[721]), .CLK(clk), .RST(rst), .Q(sreg[1741])
         );
  DFF \sreg_reg[1742]  ( .D(swire[722]), .CLK(clk), .RST(rst), .Q(sreg[1742])
         );
  DFF \sreg_reg[1743]  ( .D(swire[723]), .CLK(clk), .RST(rst), .Q(sreg[1743])
         );
  DFF \sreg_reg[1744]  ( .D(swire[724]), .CLK(clk), .RST(rst), .Q(sreg[1744])
         );
  DFF \sreg_reg[1745]  ( .D(swire[725]), .CLK(clk), .RST(rst), .Q(sreg[1745])
         );
  DFF \sreg_reg[1746]  ( .D(swire[726]), .CLK(clk), .RST(rst), .Q(sreg[1746])
         );
  DFF \sreg_reg[1747]  ( .D(swire[727]), .CLK(clk), .RST(rst), .Q(sreg[1747])
         );
  DFF \sreg_reg[1748]  ( .D(swire[728]), .CLK(clk), .RST(rst), .Q(sreg[1748])
         );
  DFF \sreg_reg[1749]  ( .D(swire[729]), .CLK(clk), .RST(rst), .Q(sreg[1749])
         );
  DFF \sreg_reg[1750]  ( .D(swire[730]), .CLK(clk), .RST(rst), .Q(sreg[1750])
         );
  DFF \sreg_reg[1751]  ( .D(swire[731]), .CLK(clk), .RST(rst), .Q(sreg[1751])
         );
  DFF \sreg_reg[1752]  ( .D(swire[732]), .CLK(clk), .RST(rst), .Q(sreg[1752])
         );
  DFF \sreg_reg[1753]  ( .D(swire[733]), .CLK(clk), .RST(rst), .Q(sreg[1753])
         );
  DFF \sreg_reg[1754]  ( .D(swire[734]), .CLK(clk), .RST(rst), .Q(sreg[1754])
         );
  DFF \sreg_reg[1755]  ( .D(swire[735]), .CLK(clk), .RST(rst), .Q(sreg[1755])
         );
  DFF \sreg_reg[1756]  ( .D(swire[736]), .CLK(clk), .RST(rst), .Q(sreg[1756])
         );
  DFF \sreg_reg[1757]  ( .D(swire[737]), .CLK(clk), .RST(rst), .Q(sreg[1757])
         );
  DFF \sreg_reg[1758]  ( .D(swire[738]), .CLK(clk), .RST(rst), .Q(sreg[1758])
         );
  DFF \sreg_reg[1759]  ( .D(swire[739]), .CLK(clk), .RST(rst), .Q(sreg[1759])
         );
  DFF \sreg_reg[1760]  ( .D(swire[740]), .CLK(clk), .RST(rst), .Q(sreg[1760])
         );
  DFF \sreg_reg[1761]  ( .D(swire[741]), .CLK(clk), .RST(rst), .Q(sreg[1761])
         );
  DFF \sreg_reg[1762]  ( .D(swire[742]), .CLK(clk), .RST(rst), .Q(sreg[1762])
         );
  DFF \sreg_reg[1763]  ( .D(swire[743]), .CLK(clk), .RST(rst), .Q(sreg[1763])
         );
  DFF \sreg_reg[1764]  ( .D(swire[744]), .CLK(clk), .RST(rst), .Q(sreg[1764])
         );
  DFF \sreg_reg[1765]  ( .D(swire[745]), .CLK(clk), .RST(rst), .Q(sreg[1765])
         );
  DFF \sreg_reg[1766]  ( .D(swire[746]), .CLK(clk), .RST(rst), .Q(sreg[1766])
         );
  DFF \sreg_reg[1767]  ( .D(swire[747]), .CLK(clk), .RST(rst), .Q(sreg[1767])
         );
  DFF \sreg_reg[1768]  ( .D(swire[748]), .CLK(clk), .RST(rst), .Q(sreg[1768])
         );
  DFF \sreg_reg[1769]  ( .D(swire[749]), .CLK(clk), .RST(rst), .Q(sreg[1769])
         );
  DFF \sreg_reg[1770]  ( .D(swire[750]), .CLK(clk), .RST(rst), .Q(sreg[1770])
         );
  DFF \sreg_reg[1771]  ( .D(swire[751]), .CLK(clk), .RST(rst), .Q(sreg[1771])
         );
  DFF \sreg_reg[1772]  ( .D(swire[752]), .CLK(clk), .RST(rst), .Q(sreg[1772])
         );
  DFF \sreg_reg[1773]  ( .D(swire[753]), .CLK(clk), .RST(rst), .Q(sreg[1773])
         );
  DFF \sreg_reg[1774]  ( .D(swire[754]), .CLK(clk), .RST(rst), .Q(sreg[1774])
         );
  DFF \sreg_reg[1775]  ( .D(swire[755]), .CLK(clk), .RST(rst), .Q(sreg[1775])
         );
  DFF \sreg_reg[1776]  ( .D(swire[756]), .CLK(clk), .RST(rst), .Q(sreg[1776])
         );
  DFF \sreg_reg[1777]  ( .D(swire[757]), .CLK(clk), .RST(rst), .Q(sreg[1777])
         );
  DFF \sreg_reg[1778]  ( .D(swire[758]), .CLK(clk), .RST(rst), .Q(sreg[1778])
         );
  DFF \sreg_reg[1779]  ( .D(swire[759]), .CLK(clk), .RST(rst), .Q(sreg[1779])
         );
  DFF \sreg_reg[1780]  ( .D(swire[760]), .CLK(clk), .RST(rst), .Q(sreg[1780])
         );
  DFF \sreg_reg[1781]  ( .D(swire[761]), .CLK(clk), .RST(rst), .Q(sreg[1781])
         );
  DFF \sreg_reg[1782]  ( .D(swire[762]), .CLK(clk), .RST(rst), .Q(sreg[1782])
         );
  DFF \sreg_reg[1783]  ( .D(swire[763]), .CLK(clk), .RST(rst), .Q(sreg[1783])
         );
  DFF \sreg_reg[1784]  ( .D(swire[764]), .CLK(clk), .RST(rst), .Q(sreg[1784])
         );
  DFF \sreg_reg[1785]  ( .D(swire[765]), .CLK(clk), .RST(rst), .Q(sreg[1785])
         );
  DFF \sreg_reg[1786]  ( .D(swire[766]), .CLK(clk), .RST(rst), .Q(sreg[1786])
         );
  DFF \sreg_reg[1787]  ( .D(swire[767]), .CLK(clk), .RST(rst), .Q(sreg[1787])
         );
  DFF \sreg_reg[1788]  ( .D(swire[768]), .CLK(clk), .RST(rst), .Q(sreg[1788])
         );
  DFF \sreg_reg[1789]  ( .D(swire[769]), .CLK(clk), .RST(rst), .Q(sreg[1789])
         );
  DFF \sreg_reg[1790]  ( .D(swire[770]), .CLK(clk), .RST(rst), .Q(sreg[1790])
         );
  DFF \sreg_reg[1791]  ( .D(swire[771]), .CLK(clk), .RST(rst), .Q(sreg[1791])
         );
  DFF \sreg_reg[1792]  ( .D(swire[772]), .CLK(clk), .RST(rst), .Q(sreg[1792])
         );
  DFF \sreg_reg[1793]  ( .D(swire[773]), .CLK(clk), .RST(rst), .Q(sreg[1793])
         );
  DFF \sreg_reg[1794]  ( .D(swire[774]), .CLK(clk), .RST(rst), .Q(sreg[1794])
         );
  DFF \sreg_reg[1795]  ( .D(swire[775]), .CLK(clk), .RST(rst), .Q(sreg[1795])
         );
  DFF \sreg_reg[1796]  ( .D(swire[776]), .CLK(clk), .RST(rst), .Q(sreg[1796])
         );
  DFF \sreg_reg[1797]  ( .D(swire[777]), .CLK(clk), .RST(rst), .Q(sreg[1797])
         );
  DFF \sreg_reg[1798]  ( .D(swire[778]), .CLK(clk), .RST(rst), .Q(sreg[1798])
         );
  DFF \sreg_reg[1799]  ( .D(swire[779]), .CLK(clk), .RST(rst), .Q(sreg[1799])
         );
  DFF \sreg_reg[1800]  ( .D(swire[780]), .CLK(clk), .RST(rst), .Q(sreg[1800])
         );
  DFF \sreg_reg[1801]  ( .D(swire[781]), .CLK(clk), .RST(rst), .Q(sreg[1801])
         );
  DFF \sreg_reg[1802]  ( .D(swire[782]), .CLK(clk), .RST(rst), .Q(sreg[1802])
         );
  DFF \sreg_reg[1803]  ( .D(swire[783]), .CLK(clk), .RST(rst), .Q(sreg[1803])
         );
  DFF \sreg_reg[1804]  ( .D(swire[784]), .CLK(clk), .RST(rst), .Q(sreg[1804])
         );
  DFF \sreg_reg[1805]  ( .D(swire[785]), .CLK(clk), .RST(rst), .Q(sreg[1805])
         );
  DFF \sreg_reg[1806]  ( .D(swire[786]), .CLK(clk), .RST(rst), .Q(sreg[1806])
         );
  DFF \sreg_reg[1807]  ( .D(swire[787]), .CLK(clk), .RST(rst), .Q(sreg[1807])
         );
  DFF \sreg_reg[1808]  ( .D(swire[788]), .CLK(clk), .RST(rst), .Q(sreg[1808])
         );
  DFF \sreg_reg[1809]  ( .D(swire[789]), .CLK(clk), .RST(rst), .Q(sreg[1809])
         );
  DFF \sreg_reg[1810]  ( .D(swire[790]), .CLK(clk), .RST(rst), .Q(sreg[1810])
         );
  DFF \sreg_reg[1811]  ( .D(swire[791]), .CLK(clk), .RST(rst), .Q(sreg[1811])
         );
  DFF \sreg_reg[1812]  ( .D(swire[792]), .CLK(clk), .RST(rst), .Q(sreg[1812])
         );
  DFF \sreg_reg[1813]  ( .D(swire[793]), .CLK(clk), .RST(rst), .Q(sreg[1813])
         );
  DFF \sreg_reg[1814]  ( .D(swire[794]), .CLK(clk), .RST(rst), .Q(sreg[1814])
         );
  DFF \sreg_reg[1815]  ( .D(swire[795]), .CLK(clk), .RST(rst), .Q(sreg[1815])
         );
  DFF \sreg_reg[1816]  ( .D(swire[796]), .CLK(clk), .RST(rst), .Q(sreg[1816])
         );
  DFF \sreg_reg[1817]  ( .D(swire[797]), .CLK(clk), .RST(rst), .Q(sreg[1817])
         );
  DFF \sreg_reg[1818]  ( .D(swire[798]), .CLK(clk), .RST(rst), .Q(sreg[1818])
         );
  DFF \sreg_reg[1819]  ( .D(swire[799]), .CLK(clk), .RST(rst), .Q(sreg[1819])
         );
  DFF \sreg_reg[1820]  ( .D(swire[800]), .CLK(clk), .RST(rst), .Q(sreg[1820])
         );
  DFF \sreg_reg[1821]  ( .D(swire[801]), .CLK(clk), .RST(rst), .Q(sreg[1821])
         );
  DFF \sreg_reg[1822]  ( .D(swire[802]), .CLK(clk), .RST(rst), .Q(sreg[1822])
         );
  DFF \sreg_reg[1823]  ( .D(swire[803]), .CLK(clk), .RST(rst), .Q(sreg[1823])
         );
  DFF \sreg_reg[1824]  ( .D(swire[804]), .CLK(clk), .RST(rst), .Q(sreg[1824])
         );
  DFF \sreg_reg[1825]  ( .D(swire[805]), .CLK(clk), .RST(rst), .Q(sreg[1825])
         );
  DFF \sreg_reg[1826]  ( .D(swire[806]), .CLK(clk), .RST(rst), .Q(sreg[1826])
         );
  DFF \sreg_reg[1827]  ( .D(swire[807]), .CLK(clk), .RST(rst), .Q(sreg[1827])
         );
  DFF \sreg_reg[1828]  ( .D(swire[808]), .CLK(clk), .RST(rst), .Q(sreg[1828])
         );
  DFF \sreg_reg[1829]  ( .D(swire[809]), .CLK(clk), .RST(rst), .Q(sreg[1829])
         );
  DFF \sreg_reg[1830]  ( .D(swire[810]), .CLK(clk), .RST(rst), .Q(sreg[1830])
         );
  DFF \sreg_reg[1831]  ( .D(swire[811]), .CLK(clk), .RST(rst), .Q(sreg[1831])
         );
  DFF \sreg_reg[1832]  ( .D(swire[812]), .CLK(clk), .RST(rst), .Q(sreg[1832])
         );
  DFF \sreg_reg[1833]  ( .D(swire[813]), .CLK(clk), .RST(rst), .Q(sreg[1833])
         );
  DFF \sreg_reg[1834]  ( .D(swire[814]), .CLK(clk), .RST(rst), .Q(sreg[1834])
         );
  DFF \sreg_reg[1835]  ( .D(swire[815]), .CLK(clk), .RST(rst), .Q(sreg[1835])
         );
  DFF \sreg_reg[1836]  ( .D(swire[816]), .CLK(clk), .RST(rst), .Q(sreg[1836])
         );
  DFF \sreg_reg[1837]  ( .D(swire[817]), .CLK(clk), .RST(rst), .Q(sreg[1837])
         );
  DFF \sreg_reg[1838]  ( .D(swire[818]), .CLK(clk), .RST(rst), .Q(sreg[1838])
         );
  DFF \sreg_reg[1839]  ( .D(swire[819]), .CLK(clk), .RST(rst), .Q(sreg[1839])
         );
  DFF \sreg_reg[1840]  ( .D(swire[820]), .CLK(clk), .RST(rst), .Q(sreg[1840])
         );
  DFF \sreg_reg[1841]  ( .D(swire[821]), .CLK(clk), .RST(rst), .Q(sreg[1841])
         );
  DFF \sreg_reg[1842]  ( .D(swire[822]), .CLK(clk), .RST(rst), .Q(sreg[1842])
         );
  DFF \sreg_reg[1843]  ( .D(swire[823]), .CLK(clk), .RST(rst), .Q(sreg[1843])
         );
  DFF \sreg_reg[1844]  ( .D(swire[824]), .CLK(clk), .RST(rst), .Q(sreg[1844])
         );
  DFF \sreg_reg[1845]  ( .D(swire[825]), .CLK(clk), .RST(rst), .Q(sreg[1845])
         );
  DFF \sreg_reg[1846]  ( .D(swire[826]), .CLK(clk), .RST(rst), .Q(sreg[1846])
         );
  DFF \sreg_reg[1847]  ( .D(swire[827]), .CLK(clk), .RST(rst), .Q(sreg[1847])
         );
  DFF \sreg_reg[1848]  ( .D(swire[828]), .CLK(clk), .RST(rst), .Q(sreg[1848])
         );
  DFF \sreg_reg[1849]  ( .D(swire[829]), .CLK(clk), .RST(rst), .Q(sreg[1849])
         );
  DFF \sreg_reg[1850]  ( .D(swire[830]), .CLK(clk), .RST(rst), .Q(sreg[1850])
         );
  DFF \sreg_reg[1851]  ( .D(swire[831]), .CLK(clk), .RST(rst), .Q(sreg[1851])
         );
  DFF \sreg_reg[1852]  ( .D(swire[832]), .CLK(clk), .RST(rst), .Q(sreg[1852])
         );
  DFF \sreg_reg[1853]  ( .D(swire[833]), .CLK(clk), .RST(rst), .Q(sreg[1853])
         );
  DFF \sreg_reg[1854]  ( .D(swire[834]), .CLK(clk), .RST(rst), .Q(sreg[1854])
         );
  DFF \sreg_reg[1855]  ( .D(swire[835]), .CLK(clk), .RST(rst), .Q(sreg[1855])
         );
  DFF \sreg_reg[1856]  ( .D(swire[836]), .CLK(clk), .RST(rst), .Q(sreg[1856])
         );
  DFF \sreg_reg[1857]  ( .D(swire[837]), .CLK(clk), .RST(rst), .Q(sreg[1857])
         );
  DFF \sreg_reg[1858]  ( .D(swire[838]), .CLK(clk), .RST(rst), .Q(sreg[1858])
         );
  DFF \sreg_reg[1859]  ( .D(swire[839]), .CLK(clk), .RST(rst), .Q(sreg[1859])
         );
  DFF \sreg_reg[1860]  ( .D(swire[840]), .CLK(clk), .RST(rst), .Q(sreg[1860])
         );
  DFF \sreg_reg[1861]  ( .D(swire[841]), .CLK(clk), .RST(rst), .Q(sreg[1861])
         );
  DFF \sreg_reg[1862]  ( .D(swire[842]), .CLK(clk), .RST(rst), .Q(sreg[1862])
         );
  DFF \sreg_reg[1863]  ( .D(swire[843]), .CLK(clk), .RST(rst), .Q(sreg[1863])
         );
  DFF \sreg_reg[1864]  ( .D(swire[844]), .CLK(clk), .RST(rst), .Q(sreg[1864])
         );
  DFF \sreg_reg[1865]  ( .D(swire[845]), .CLK(clk), .RST(rst), .Q(sreg[1865])
         );
  DFF \sreg_reg[1866]  ( .D(swire[846]), .CLK(clk), .RST(rst), .Q(sreg[1866])
         );
  DFF \sreg_reg[1867]  ( .D(swire[847]), .CLK(clk), .RST(rst), .Q(sreg[1867])
         );
  DFF \sreg_reg[1868]  ( .D(swire[848]), .CLK(clk), .RST(rst), .Q(sreg[1868])
         );
  DFF \sreg_reg[1869]  ( .D(swire[849]), .CLK(clk), .RST(rst), .Q(sreg[1869])
         );
  DFF \sreg_reg[1870]  ( .D(swire[850]), .CLK(clk), .RST(rst), .Q(sreg[1870])
         );
  DFF \sreg_reg[1871]  ( .D(swire[851]), .CLK(clk), .RST(rst), .Q(sreg[1871])
         );
  DFF \sreg_reg[1872]  ( .D(swire[852]), .CLK(clk), .RST(rst), .Q(sreg[1872])
         );
  DFF \sreg_reg[1873]  ( .D(swire[853]), .CLK(clk), .RST(rst), .Q(sreg[1873])
         );
  DFF \sreg_reg[1874]  ( .D(swire[854]), .CLK(clk), .RST(rst), .Q(sreg[1874])
         );
  DFF \sreg_reg[1875]  ( .D(swire[855]), .CLK(clk), .RST(rst), .Q(sreg[1875])
         );
  DFF \sreg_reg[1876]  ( .D(swire[856]), .CLK(clk), .RST(rst), .Q(sreg[1876])
         );
  DFF \sreg_reg[1877]  ( .D(swire[857]), .CLK(clk), .RST(rst), .Q(sreg[1877])
         );
  DFF \sreg_reg[1878]  ( .D(swire[858]), .CLK(clk), .RST(rst), .Q(sreg[1878])
         );
  DFF \sreg_reg[1879]  ( .D(swire[859]), .CLK(clk), .RST(rst), .Q(sreg[1879])
         );
  DFF \sreg_reg[1880]  ( .D(swire[860]), .CLK(clk), .RST(rst), .Q(sreg[1880])
         );
  DFF \sreg_reg[1881]  ( .D(swire[861]), .CLK(clk), .RST(rst), .Q(sreg[1881])
         );
  DFF \sreg_reg[1882]  ( .D(swire[862]), .CLK(clk), .RST(rst), .Q(sreg[1882])
         );
  DFF \sreg_reg[1883]  ( .D(swire[863]), .CLK(clk), .RST(rst), .Q(sreg[1883])
         );
  DFF \sreg_reg[1884]  ( .D(swire[864]), .CLK(clk), .RST(rst), .Q(sreg[1884])
         );
  DFF \sreg_reg[1885]  ( .D(swire[865]), .CLK(clk), .RST(rst), .Q(sreg[1885])
         );
  DFF \sreg_reg[1886]  ( .D(swire[866]), .CLK(clk), .RST(rst), .Q(sreg[1886])
         );
  DFF \sreg_reg[1887]  ( .D(swire[867]), .CLK(clk), .RST(rst), .Q(sreg[1887])
         );
  DFF \sreg_reg[1888]  ( .D(swire[868]), .CLK(clk), .RST(rst), .Q(sreg[1888])
         );
  DFF \sreg_reg[1889]  ( .D(swire[869]), .CLK(clk), .RST(rst), .Q(sreg[1889])
         );
  DFF \sreg_reg[1890]  ( .D(swire[870]), .CLK(clk), .RST(rst), .Q(sreg[1890])
         );
  DFF \sreg_reg[1891]  ( .D(swire[871]), .CLK(clk), .RST(rst), .Q(sreg[1891])
         );
  DFF \sreg_reg[1892]  ( .D(swire[872]), .CLK(clk), .RST(rst), .Q(sreg[1892])
         );
  DFF \sreg_reg[1893]  ( .D(swire[873]), .CLK(clk), .RST(rst), .Q(sreg[1893])
         );
  DFF \sreg_reg[1894]  ( .D(swire[874]), .CLK(clk), .RST(rst), .Q(sreg[1894])
         );
  DFF \sreg_reg[1895]  ( .D(swire[875]), .CLK(clk), .RST(rst), .Q(sreg[1895])
         );
  DFF \sreg_reg[1896]  ( .D(swire[876]), .CLK(clk), .RST(rst), .Q(sreg[1896])
         );
  DFF \sreg_reg[1897]  ( .D(swire[877]), .CLK(clk), .RST(rst), .Q(sreg[1897])
         );
  DFF \sreg_reg[1898]  ( .D(swire[878]), .CLK(clk), .RST(rst), .Q(sreg[1898])
         );
  DFF \sreg_reg[1899]  ( .D(swire[879]), .CLK(clk), .RST(rst), .Q(sreg[1899])
         );
  DFF \sreg_reg[1900]  ( .D(swire[880]), .CLK(clk), .RST(rst), .Q(sreg[1900])
         );
  DFF \sreg_reg[1901]  ( .D(swire[881]), .CLK(clk), .RST(rst), .Q(sreg[1901])
         );
  DFF \sreg_reg[1902]  ( .D(swire[882]), .CLK(clk), .RST(rst), .Q(sreg[1902])
         );
  DFF \sreg_reg[1903]  ( .D(swire[883]), .CLK(clk), .RST(rst), .Q(sreg[1903])
         );
  DFF \sreg_reg[1904]  ( .D(swire[884]), .CLK(clk), .RST(rst), .Q(sreg[1904])
         );
  DFF \sreg_reg[1905]  ( .D(swire[885]), .CLK(clk), .RST(rst), .Q(sreg[1905])
         );
  DFF \sreg_reg[1906]  ( .D(swire[886]), .CLK(clk), .RST(rst), .Q(sreg[1906])
         );
  DFF \sreg_reg[1907]  ( .D(swire[887]), .CLK(clk), .RST(rst), .Q(sreg[1907])
         );
  DFF \sreg_reg[1908]  ( .D(swire[888]), .CLK(clk), .RST(rst), .Q(sreg[1908])
         );
  DFF \sreg_reg[1909]  ( .D(swire[889]), .CLK(clk), .RST(rst), .Q(sreg[1909])
         );
  DFF \sreg_reg[1910]  ( .D(swire[890]), .CLK(clk), .RST(rst), .Q(sreg[1910])
         );
  DFF \sreg_reg[1911]  ( .D(swire[891]), .CLK(clk), .RST(rst), .Q(sreg[1911])
         );
  DFF \sreg_reg[1912]  ( .D(swire[892]), .CLK(clk), .RST(rst), .Q(sreg[1912])
         );
  DFF \sreg_reg[1913]  ( .D(swire[893]), .CLK(clk), .RST(rst), .Q(sreg[1913])
         );
  DFF \sreg_reg[1914]  ( .D(swire[894]), .CLK(clk), .RST(rst), .Q(sreg[1914])
         );
  DFF \sreg_reg[1915]  ( .D(swire[895]), .CLK(clk), .RST(rst), .Q(sreg[1915])
         );
  DFF \sreg_reg[1916]  ( .D(swire[896]), .CLK(clk), .RST(rst), .Q(sreg[1916])
         );
  DFF \sreg_reg[1917]  ( .D(swire[897]), .CLK(clk), .RST(rst), .Q(sreg[1917])
         );
  DFF \sreg_reg[1918]  ( .D(swire[898]), .CLK(clk), .RST(rst), .Q(sreg[1918])
         );
  DFF \sreg_reg[1919]  ( .D(swire[899]), .CLK(clk), .RST(rst), .Q(sreg[1919])
         );
  DFF \sreg_reg[1920]  ( .D(swire[900]), .CLK(clk), .RST(rst), .Q(sreg[1920])
         );
  DFF \sreg_reg[1921]  ( .D(swire[901]), .CLK(clk), .RST(rst), .Q(sreg[1921])
         );
  DFF \sreg_reg[1922]  ( .D(swire[902]), .CLK(clk), .RST(rst), .Q(sreg[1922])
         );
  DFF \sreg_reg[1923]  ( .D(swire[903]), .CLK(clk), .RST(rst), .Q(sreg[1923])
         );
  DFF \sreg_reg[1924]  ( .D(swire[904]), .CLK(clk), .RST(rst), .Q(sreg[1924])
         );
  DFF \sreg_reg[1925]  ( .D(swire[905]), .CLK(clk), .RST(rst), .Q(sreg[1925])
         );
  DFF \sreg_reg[1926]  ( .D(swire[906]), .CLK(clk), .RST(rst), .Q(sreg[1926])
         );
  DFF \sreg_reg[1927]  ( .D(swire[907]), .CLK(clk), .RST(rst), .Q(sreg[1927])
         );
  DFF \sreg_reg[1928]  ( .D(swire[908]), .CLK(clk), .RST(rst), .Q(sreg[1928])
         );
  DFF \sreg_reg[1929]  ( .D(swire[909]), .CLK(clk), .RST(rst), .Q(sreg[1929])
         );
  DFF \sreg_reg[1930]  ( .D(swire[910]), .CLK(clk), .RST(rst), .Q(sreg[1930])
         );
  DFF \sreg_reg[1931]  ( .D(swire[911]), .CLK(clk), .RST(rst), .Q(sreg[1931])
         );
  DFF \sreg_reg[1932]  ( .D(swire[912]), .CLK(clk), .RST(rst), .Q(sreg[1932])
         );
  DFF \sreg_reg[1933]  ( .D(swire[913]), .CLK(clk), .RST(rst), .Q(sreg[1933])
         );
  DFF \sreg_reg[1934]  ( .D(swire[914]), .CLK(clk), .RST(rst), .Q(sreg[1934])
         );
  DFF \sreg_reg[1935]  ( .D(swire[915]), .CLK(clk), .RST(rst), .Q(sreg[1935])
         );
  DFF \sreg_reg[1936]  ( .D(swire[916]), .CLK(clk), .RST(rst), .Q(sreg[1936])
         );
  DFF \sreg_reg[1937]  ( .D(swire[917]), .CLK(clk), .RST(rst), .Q(sreg[1937])
         );
  DFF \sreg_reg[1938]  ( .D(swire[918]), .CLK(clk), .RST(rst), .Q(sreg[1938])
         );
  DFF \sreg_reg[1939]  ( .D(swire[919]), .CLK(clk), .RST(rst), .Q(sreg[1939])
         );
  DFF \sreg_reg[1940]  ( .D(swire[920]), .CLK(clk), .RST(rst), .Q(sreg[1940])
         );
  DFF \sreg_reg[1941]  ( .D(swire[921]), .CLK(clk), .RST(rst), .Q(sreg[1941])
         );
  DFF \sreg_reg[1942]  ( .D(swire[922]), .CLK(clk), .RST(rst), .Q(sreg[1942])
         );
  DFF \sreg_reg[1943]  ( .D(swire[923]), .CLK(clk), .RST(rst), .Q(sreg[1943])
         );
  DFF \sreg_reg[1944]  ( .D(swire[924]), .CLK(clk), .RST(rst), .Q(sreg[1944])
         );
  DFF \sreg_reg[1945]  ( .D(swire[925]), .CLK(clk), .RST(rst), .Q(sreg[1945])
         );
  DFF \sreg_reg[1946]  ( .D(swire[926]), .CLK(clk), .RST(rst), .Q(sreg[1946])
         );
  DFF \sreg_reg[1947]  ( .D(swire[927]), .CLK(clk), .RST(rst), .Q(sreg[1947])
         );
  DFF \sreg_reg[1948]  ( .D(swire[928]), .CLK(clk), .RST(rst), .Q(sreg[1948])
         );
  DFF \sreg_reg[1949]  ( .D(swire[929]), .CLK(clk), .RST(rst), .Q(sreg[1949])
         );
  DFF \sreg_reg[1950]  ( .D(swire[930]), .CLK(clk), .RST(rst), .Q(sreg[1950])
         );
  DFF \sreg_reg[1951]  ( .D(swire[931]), .CLK(clk), .RST(rst), .Q(sreg[1951])
         );
  DFF \sreg_reg[1952]  ( .D(swire[932]), .CLK(clk), .RST(rst), .Q(sreg[1952])
         );
  DFF \sreg_reg[1953]  ( .D(swire[933]), .CLK(clk), .RST(rst), .Q(sreg[1953])
         );
  DFF \sreg_reg[1954]  ( .D(swire[934]), .CLK(clk), .RST(rst), .Q(sreg[1954])
         );
  DFF \sreg_reg[1955]  ( .D(swire[935]), .CLK(clk), .RST(rst), .Q(sreg[1955])
         );
  DFF \sreg_reg[1956]  ( .D(swire[936]), .CLK(clk), .RST(rst), .Q(sreg[1956])
         );
  DFF \sreg_reg[1957]  ( .D(swire[937]), .CLK(clk), .RST(rst), .Q(sreg[1957])
         );
  DFF \sreg_reg[1958]  ( .D(swire[938]), .CLK(clk), .RST(rst), .Q(sreg[1958])
         );
  DFF \sreg_reg[1959]  ( .D(swire[939]), .CLK(clk), .RST(rst), .Q(sreg[1959])
         );
  DFF \sreg_reg[1960]  ( .D(swire[940]), .CLK(clk), .RST(rst), .Q(sreg[1960])
         );
  DFF \sreg_reg[1961]  ( .D(swire[941]), .CLK(clk), .RST(rst), .Q(sreg[1961])
         );
  DFF \sreg_reg[1962]  ( .D(swire[942]), .CLK(clk), .RST(rst), .Q(sreg[1962])
         );
  DFF \sreg_reg[1963]  ( .D(swire[943]), .CLK(clk), .RST(rst), .Q(sreg[1963])
         );
  DFF \sreg_reg[1964]  ( .D(swire[944]), .CLK(clk), .RST(rst), .Q(sreg[1964])
         );
  DFF \sreg_reg[1965]  ( .D(swire[945]), .CLK(clk), .RST(rst), .Q(sreg[1965])
         );
  DFF \sreg_reg[1966]  ( .D(swire[946]), .CLK(clk), .RST(rst), .Q(sreg[1966])
         );
  DFF \sreg_reg[1967]  ( .D(swire[947]), .CLK(clk), .RST(rst), .Q(sreg[1967])
         );
  DFF \sreg_reg[1968]  ( .D(swire[948]), .CLK(clk), .RST(rst), .Q(sreg[1968])
         );
  DFF \sreg_reg[1969]  ( .D(swire[949]), .CLK(clk), .RST(rst), .Q(sreg[1969])
         );
  DFF \sreg_reg[1970]  ( .D(swire[950]), .CLK(clk), .RST(rst), .Q(sreg[1970])
         );
  DFF \sreg_reg[1971]  ( .D(swire[951]), .CLK(clk), .RST(rst), .Q(sreg[1971])
         );
  DFF \sreg_reg[1972]  ( .D(swire[952]), .CLK(clk), .RST(rst), .Q(sreg[1972])
         );
  DFF \sreg_reg[1973]  ( .D(swire[953]), .CLK(clk), .RST(rst), .Q(sreg[1973])
         );
  DFF \sreg_reg[1974]  ( .D(swire[954]), .CLK(clk), .RST(rst), .Q(sreg[1974])
         );
  DFF \sreg_reg[1975]  ( .D(swire[955]), .CLK(clk), .RST(rst), .Q(sreg[1975])
         );
  DFF \sreg_reg[1976]  ( .D(swire[956]), .CLK(clk), .RST(rst), .Q(sreg[1976])
         );
  DFF \sreg_reg[1977]  ( .D(swire[957]), .CLK(clk), .RST(rst), .Q(sreg[1977])
         );
  DFF \sreg_reg[1978]  ( .D(swire[958]), .CLK(clk), .RST(rst), .Q(sreg[1978])
         );
  DFF \sreg_reg[1979]  ( .D(swire[959]), .CLK(clk), .RST(rst), .Q(sreg[1979])
         );
  DFF \sreg_reg[1980]  ( .D(swire[960]), .CLK(clk), .RST(rst), .Q(sreg[1980])
         );
  DFF \sreg_reg[1981]  ( .D(swire[961]), .CLK(clk), .RST(rst), .Q(sreg[1981])
         );
  DFF \sreg_reg[1982]  ( .D(swire[962]), .CLK(clk), .RST(rst), .Q(sreg[1982])
         );
  DFF \sreg_reg[1983]  ( .D(swire[963]), .CLK(clk), .RST(rst), .Q(sreg[1983])
         );
  DFF \sreg_reg[1984]  ( .D(swire[964]), .CLK(clk), .RST(rst), .Q(sreg[1984])
         );
  DFF \sreg_reg[1985]  ( .D(swire[965]), .CLK(clk), .RST(rst), .Q(sreg[1985])
         );
  DFF \sreg_reg[1986]  ( .D(swire[966]), .CLK(clk), .RST(rst), .Q(sreg[1986])
         );
  DFF \sreg_reg[1987]  ( .D(swire[967]), .CLK(clk), .RST(rst), .Q(sreg[1987])
         );
  DFF \sreg_reg[1988]  ( .D(swire[968]), .CLK(clk), .RST(rst), .Q(sreg[1988])
         );
  DFF \sreg_reg[1989]  ( .D(swire[969]), .CLK(clk), .RST(rst), .Q(sreg[1989])
         );
  DFF \sreg_reg[1990]  ( .D(swire[970]), .CLK(clk), .RST(rst), .Q(sreg[1990])
         );
  DFF \sreg_reg[1991]  ( .D(swire[971]), .CLK(clk), .RST(rst), .Q(sreg[1991])
         );
  DFF \sreg_reg[1992]  ( .D(swire[972]), .CLK(clk), .RST(rst), .Q(sreg[1992])
         );
  DFF \sreg_reg[1993]  ( .D(swire[973]), .CLK(clk), .RST(rst), .Q(sreg[1993])
         );
  DFF \sreg_reg[1994]  ( .D(swire[974]), .CLK(clk), .RST(rst), .Q(sreg[1994])
         );
  DFF \sreg_reg[1995]  ( .D(swire[975]), .CLK(clk), .RST(rst), .Q(sreg[1995])
         );
  DFF \sreg_reg[1996]  ( .D(swire[976]), .CLK(clk), .RST(rst), .Q(sreg[1996])
         );
  DFF \sreg_reg[1997]  ( .D(swire[977]), .CLK(clk), .RST(rst), .Q(sreg[1997])
         );
  DFF \sreg_reg[1998]  ( .D(swire[978]), .CLK(clk), .RST(rst), .Q(sreg[1998])
         );
  DFF \sreg_reg[1999]  ( .D(swire[979]), .CLK(clk), .RST(rst), .Q(sreg[1999])
         );
  DFF \sreg_reg[2000]  ( .D(swire[980]), .CLK(clk), .RST(rst), .Q(sreg[2000])
         );
  DFF \sreg_reg[2001]  ( .D(swire[981]), .CLK(clk), .RST(rst), .Q(sreg[2001])
         );
  DFF \sreg_reg[2002]  ( .D(swire[982]), .CLK(clk), .RST(rst), .Q(sreg[2002])
         );
  DFF \sreg_reg[2003]  ( .D(swire[983]), .CLK(clk), .RST(rst), .Q(sreg[2003])
         );
  DFF \sreg_reg[2004]  ( .D(swire[984]), .CLK(clk), .RST(rst), .Q(sreg[2004])
         );
  DFF \sreg_reg[2005]  ( .D(swire[985]), .CLK(clk), .RST(rst), .Q(sreg[2005])
         );
  DFF \sreg_reg[2006]  ( .D(swire[986]), .CLK(clk), .RST(rst), .Q(sreg[2006])
         );
  DFF \sreg_reg[2007]  ( .D(swire[987]), .CLK(clk), .RST(rst), .Q(sreg[2007])
         );
  DFF \sreg_reg[2008]  ( .D(swire[988]), .CLK(clk), .RST(rst), .Q(sreg[2008])
         );
  DFF \sreg_reg[2009]  ( .D(swire[989]), .CLK(clk), .RST(rst), .Q(sreg[2009])
         );
  DFF \sreg_reg[2010]  ( .D(swire[990]), .CLK(clk), .RST(rst), .Q(sreg[2010])
         );
  DFF \sreg_reg[2011]  ( .D(swire[991]), .CLK(clk), .RST(rst), .Q(sreg[2011])
         );
  DFF \sreg_reg[2012]  ( .D(swire[992]), .CLK(clk), .RST(rst), .Q(sreg[2012])
         );
  DFF \sreg_reg[2013]  ( .D(swire[993]), .CLK(clk), .RST(rst), .Q(sreg[2013])
         );
  DFF \sreg_reg[2014]  ( .D(swire[994]), .CLK(clk), .RST(rst), .Q(sreg[2014])
         );
  DFF \sreg_reg[2015]  ( .D(swire[995]), .CLK(clk), .RST(rst), .Q(sreg[2015])
         );
  DFF \sreg_reg[2016]  ( .D(swire[996]), .CLK(clk), .RST(rst), .Q(sreg[2016])
         );
  DFF \sreg_reg[2017]  ( .D(swire[997]), .CLK(clk), .RST(rst), .Q(sreg[2017])
         );
  DFF \sreg_reg[2018]  ( .D(swire[998]), .CLK(clk), .RST(rst), .Q(sreg[2018])
         );
  DFF \sreg_reg[2019]  ( .D(swire[999]), .CLK(clk), .RST(rst), .Q(sreg[2019])
         );
  DFF \sreg_reg[2020]  ( .D(swire[1000]), .CLK(clk), .RST(rst), .Q(sreg[2020])
         );
  DFF \sreg_reg[2021]  ( .D(swire[1001]), .CLK(clk), .RST(rst), .Q(sreg[2021])
         );
  DFF \sreg_reg[2022]  ( .D(swire[1002]), .CLK(clk), .RST(rst), .Q(sreg[2022])
         );
  DFF \sreg_reg[2023]  ( .D(swire[1003]), .CLK(clk), .RST(rst), .Q(sreg[2023])
         );
  DFF \sreg_reg[2024]  ( .D(swire[1004]), .CLK(clk), .RST(rst), .Q(sreg[2024])
         );
  DFF \sreg_reg[2025]  ( .D(swire[1005]), .CLK(clk), .RST(rst), .Q(sreg[2025])
         );
  DFF \sreg_reg[2026]  ( .D(swire[1006]), .CLK(clk), .RST(rst), .Q(sreg[2026])
         );
  DFF \sreg_reg[2027]  ( .D(swire[1007]), .CLK(clk), .RST(rst), .Q(sreg[2027])
         );
  DFF \sreg_reg[2028]  ( .D(swire[1008]), .CLK(clk), .RST(rst), .Q(sreg[2028])
         );
  DFF \sreg_reg[2029]  ( .D(swire[1009]), .CLK(clk), .RST(rst), .Q(sreg[2029])
         );
  DFF \sreg_reg[2030]  ( .D(swire[1010]), .CLK(clk), .RST(rst), .Q(sreg[2030])
         );
  DFF \sreg_reg[2031]  ( .D(swire[1011]), .CLK(clk), .RST(rst), .Q(sreg[2031])
         );
  DFF \sreg_reg[2032]  ( .D(swire[1012]), .CLK(clk), .RST(rst), .Q(sreg[2032])
         );
  DFF \sreg_reg[2033]  ( .D(swire[1013]), .CLK(clk), .RST(rst), .Q(sreg[2033])
         );
  DFF \sreg_reg[2034]  ( .D(swire[1014]), .CLK(clk), .RST(rst), .Q(sreg[2034])
         );
  DFF \sreg_reg[2035]  ( .D(swire[1015]), .CLK(clk), .RST(rst), .Q(sreg[2035])
         );
  DFF \sreg_reg[2036]  ( .D(swire[1016]), .CLK(clk), .RST(rst), .Q(sreg[2036])
         );
  DFF \sreg_reg[2037]  ( .D(swire[1017]), .CLK(clk), .RST(rst), .Q(sreg[2037])
         );
  DFF \sreg_reg[2038]  ( .D(swire[1018]), .CLK(clk), .RST(rst), .Q(sreg[2038])
         );
  DFF \sreg_reg[2039]  ( .D(swire[1019]), .CLK(clk), .RST(rst), .Q(sreg[2039])
         );
  DFF \sreg_reg[2040]  ( .D(swire[1020]), .CLK(clk), .RST(rst), .Q(sreg[2040])
         );
  DFF \sreg_reg[2041]  ( .D(swire[1021]), .CLK(clk), .RST(rst), .Q(sreg[2041])
         );
  DFF \sreg_reg[2042]  ( .D(swire[1022]), .CLK(clk), .RST(rst), .Q(sreg[2042])
         );
  DFF \sreg_reg[2043]  ( .D(swire[1023]), .CLK(clk), .RST(rst), .Q(sreg[2043])
         );
  DFF \sreg_reg[1023]  ( .D(c[1023]), .CLK(clk), .RST(rst), .Q(c[1019]) );
  DFF \sreg_reg[1022]  ( .D(c[1022]), .CLK(clk), .RST(rst), .Q(c[1018]) );
  DFF \sreg_reg[1021]  ( .D(c[1021]), .CLK(clk), .RST(rst), .Q(c[1017]) );
  DFF \sreg_reg[1020]  ( .D(c[1020]), .CLK(clk), .RST(rst), .Q(c[1016]) );
  DFF \sreg_reg[1019]  ( .D(c[1019]), .CLK(clk), .RST(rst), .Q(c[1015]) );
  DFF \sreg_reg[1018]  ( .D(c[1018]), .CLK(clk), .RST(rst), .Q(c[1014]) );
  DFF \sreg_reg[1017]  ( .D(c[1017]), .CLK(clk), .RST(rst), .Q(c[1013]) );
  DFF \sreg_reg[1016]  ( .D(c[1016]), .CLK(clk), .RST(rst), .Q(c[1012]) );
  DFF \sreg_reg[1015]  ( .D(c[1015]), .CLK(clk), .RST(rst), .Q(c[1011]) );
  DFF \sreg_reg[1014]  ( .D(c[1014]), .CLK(clk), .RST(rst), .Q(c[1010]) );
  DFF \sreg_reg[1013]  ( .D(c[1013]), .CLK(clk), .RST(rst), .Q(c[1009]) );
  DFF \sreg_reg[1012]  ( .D(c[1012]), .CLK(clk), .RST(rst), .Q(c[1008]) );
  DFF \sreg_reg[1011]  ( .D(c[1011]), .CLK(clk), .RST(rst), .Q(c[1007]) );
  DFF \sreg_reg[1010]  ( .D(c[1010]), .CLK(clk), .RST(rst), .Q(c[1006]) );
  DFF \sreg_reg[1009]  ( .D(c[1009]), .CLK(clk), .RST(rst), .Q(c[1005]) );
  DFF \sreg_reg[1008]  ( .D(c[1008]), .CLK(clk), .RST(rst), .Q(c[1004]) );
  DFF \sreg_reg[1007]  ( .D(c[1007]), .CLK(clk), .RST(rst), .Q(c[1003]) );
  DFF \sreg_reg[1006]  ( .D(c[1006]), .CLK(clk), .RST(rst), .Q(c[1002]) );
  DFF \sreg_reg[1005]  ( .D(c[1005]), .CLK(clk), .RST(rst), .Q(c[1001]) );
  DFF \sreg_reg[1004]  ( .D(c[1004]), .CLK(clk), .RST(rst), .Q(c[1000]) );
  DFF \sreg_reg[1003]  ( .D(c[1003]), .CLK(clk), .RST(rst), .Q(c[999]) );
  DFF \sreg_reg[1002]  ( .D(c[1002]), .CLK(clk), .RST(rst), .Q(c[998]) );
  DFF \sreg_reg[1001]  ( .D(c[1001]), .CLK(clk), .RST(rst), .Q(c[997]) );
  DFF \sreg_reg[1000]  ( .D(c[1000]), .CLK(clk), .RST(rst), .Q(c[996]) );
  DFF \sreg_reg[999]  ( .D(c[999]), .CLK(clk), .RST(rst), .Q(c[995]) );
  DFF \sreg_reg[998]  ( .D(c[998]), .CLK(clk), .RST(rst), .Q(c[994]) );
  DFF \sreg_reg[997]  ( .D(c[997]), .CLK(clk), .RST(rst), .Q(c[993]) );
  DFF \sreg_reg[996]  ( .D(c[996]), .CLK(clk), .RST(rst), .Q(c[992]) );
  DFF \sreg_reg[995]  ( .D(c[995]), .CLK(clk), .RST(rst), .Q(c[991]) );
  DFF \sreg_reg[994]  ( .D(c[994]), .CLK(clk), .RST(rst), .Q(c[990]) );
  DFF \sreg_reg[993]  ( .D(c[993]), .CLK(clk), .RST(rst), .Q(c[989]) );
  DFF \sreg_reg[992]  ( .D(c[992]), .CLK(clk), .RST(rst), .Q(c[988]) );
  DFF \sreg_reg[991]  ( .D(c[991]), .CLK(clk), .RST(rst), .Q(c[987]) );
  DFF \sreg_reg[990]  ( .D(c[990]), .CLK(clk), .RST(rst), .Q(c[986]) );
  DFF \sreg_reg[989]  ( .D(c[989]), .CLK(clk), .RST(rst), .Q(c[985]) );
  DFF \sreg_reg[988]  ( .D(c[988]), .CLK(clk), .RST(rst), .Q(c[984]) );
  DFF \sreg_reg[987]  ( .D(c[987]), .CLK(clk), .RST(rst), .Q(c[983]) );
  DFF \sreg_reg[986]  ( .D(c[986]), .CLK(clk), .RST(rst), .Q(c[982]) );
  DFF \sreg_reg[985]  ( .D(c[985]), .CLK(clk), .RST(rst), .Q(c[981]) );
  DFF \sreg_reg[984]  ( .D(c[984]), .CLK(clk), .RST(rst), .Q(c[980]) );
  DFF \sreg_reg[983]  ( .D(c[983]), .CLK(clk), .RST(rst), .Q(c[979]) );
  DFF \sreg_reg[982]  ( .D(c[982]), .CLK(clk), .RST(rst), .Q(c[978]) );
  DFF \sreg_reg[981]  ( .D(c[981]), .CLK(clk), .RST(rst), .Q(c[977]) );
  DFF \sreg_reg[980]  ( .D(c[980]), .CLK(clk), .RST(rst), .Q(c[976]) );
  DFF \sreg_reg[979]  ( .D(c[979]), .CLK(clk), .RST(rst), .Q(c[975]) );
  DFF \sreg_reg[978]  ( .D(c[978]), .CLK(clk), .RST(rst), .Q(c[974]) );
  DFF \sreg_reg[977]  ( .D(c[977]), .CLK(clk), .RST(rst), .Q(c[973]) );
  DFF \sreg_reg[976]  ( .D(c[976]), .CLK(clk), .RST(rst), .Q(c[972]) );
  DFF \sreg_reg[975]  ( .D(c[975]), .CLK(clk), .RST(rst), .Q(c[971]) );
  DFF \sreg_reg[974]  ( .D(c[974]), .CLK(clk), .RST(rst), .Q(c[970]) );
  DFF \sreg_reg[973]  ( .D(c[973]), .CLK(clk), .RST(rst), .Q(c[969]) );
  DFF \sreg_reg[972]  ( .D(c[972]), .CLK(clk), .RST(rst), .Q(c[968]) );
  DFF \sreg_reg[971]  ( .D(c[971]), .CLK(clk), .RST(rst), .Q(c[967]) );
  DFF \sreg_reg[970]  ( .D(c[970]), .CLK(clk), .RST(rst), .Q(c[966]) );
  DFF \sreg_reg[969]  ( .D(c[969]), .CLK(clk), .RST(rst), .Q(c[965]) );
  DFF \sreg_reg[968]  ( .D(c[968]), .CLK(clk), .RST(rst), .Q(c[964]) );
  DFF \sreg_reg[967]  ( .D(c[967]), .CLK(clk), .RST(rst), .Q(c[963]) );
  DFF \sreg_reg[966]  ( .D(c[966]), .CLK(clk), .RST(rst), .Q(c[962]) );
  DFF \sreg_reg[965]  ( .D(c[965]), .CLK(clk), .RST(rst), .Q(c[961]) );
  DFF \sreg_reg[964]  ( .D(c[964]), .CLK(clk), .RST(rst), .Q(c[960]) );
  DFF \sreg_reg[963]  ( .D(c[963]), .CLK(clk), .RST(rst), .Q(c[959]) );
  DFF \sreg_reg[962]  ( .D(c[962]), .CLK(clk), .RST(rst), .Q(c[958]) );
  DFF \sreg_reg[961]  ( .D(c[961]), .CLK(clk), .RST(rst), .Q(c[957]) );
  DFF \sreg_reg[960]  ( .D(c[960]), .CLK(clk), .RST(rst), .Q(c[956]) );
  DFF \sreg_reg[959]  ( .D(c[959]), .CLK(clk), .RST(rst), .Q(c[955]) );
  DFF \sreg_reg[958]  ( .D(c[958]), .CLK(clk), .RST(rst), .Q(c[954]) );
  DFF \sreg_reg[957]  ( .D(c[957]), .CLK(clk), .RST(rst), .Q(c[953]) );
  DFF \sreg_reg[956]  ( .D(c[956]), .CLK(clk), .RST(rst), .Q(c[952]) );
  DFF \sreg_reg[955]  ( .D(c[955]), .CLK(clk), .RST(rst), .Q(c[951]) );
  DFF \sreg_reg[954]  ( .D(c[954]), .CLK(clk), .RST(rst), .Q(c[950]) );
  DFF \sreg_reg[953]  ( .D(c[953]), .CLK(clk), .RST(rst), .Q(c[949]) );
  DFF \sreg_reg[952]  ( .D(c[952]), .CLK(clk), .RST(rst), .Q(c[948]) );
  DFF \sreg_reg[951]  ( .D(c[951]), .CLK(clk), .RST(rst), .Q(c[947]) );
  DFF \sreg_reg[950]  ( .D(c[950]), .CLK(clk), .RST(rst), .Q(c[946]) );
  DFF \sreg_reg[949]  ( .D(c[949]), .CLK(clk), .RST(rst), .Q(c[945]) );
  DFF \sreg_reg[948]  ( .D(c[948]), .CLK(clk), .RST(rst), .Q(c[944]) );
  DFF \sreg_reg[947]  ( .D(c[947]), .CLK(clk), .RST(rst), .Q(c[943]) );
  DFF \sreg_reg[946]  ( .D(c[946]), .CLK(clk), .RST(rst), .Q(c[942]) );
  DFF \sreg_reg[945]  ( .D(c[945]), .CLK(clk), .RST(rst), .Q(c[941]) );
  DFF \sreg_reg[944]  ( .D(c[944]), .CLK(clk), .RST(rst), .Q(c[940]) );
  DFF \sreg_reg[943]  ( .D(c[943]), .CLK(clk), .RST(rst), .Q(c[939]) );
  DFF \sreg_reg[942]  ( .D(c[942]), .CLK(clk), .RST(rst), .Q(c[938]) );
  DFF \sreg_reg[941]  ( .D(c[941]), .CLK(clk), .RST(rst), .Q(c[937]) );
  DFF \sreg_reg[940]  ( .D(c[940]), .CLK(clk), .RST(rst), .Q(c[936]) );
  DFF \sreg_reg[939]  ( .D(c[939]), .CLK(clk), .RST(rst), .Q(c[935]) );
  DFF \sreg_reg[938]  ( .D(c[938]), .CLK(clk), .RST(rst), .Q(c[934]) );
  DFF \sreg_reg[937]  ( .D(c[937]), .CLK(clk), .RST(rst), .Q(c[933]) );
  DFF \sreg_reg[936]  ( .D(c[936]), .CLK(clk), .RST(rst), .Q(c[932]) );
  DFF \sreg_reg[935]  ( .D(c[935]), .CLK(clk), .RST(rst), .Q(c[931]) );
  DFF \sreg_reg[934]  ( .D(c[934]), .CLK(clk), .RST(rst), .Q(c[930]) );
  DFF \sreg_reg[933]  ( .D(c[933]), .CLK(clk), .RST(rst), .Q(c[929]) );
  DFF \sreg_reg[932]  ( .D(c[932]), .CLK(clk), .RST(rst), .Q(c[928]) );
  DFF \sreg_reg[931]  ( .D(c[931]), .CLK(clk), .RST(rst), .Q(c[927]) );
  DFF \sreg_reg[930]  ( .D(c[930]), .CLK(clk), .RST(rst), .Q(c[926]) );
  DFF \sreg_reg[929]  ( .D(c[929]), .CLK(clk), .RST(rst), .Q(c[925]) );
  DFF \sreg_reg[928]  ( .D(c[928]), .CLK(clk), .RST(rst), .Q(c[924]) );
  DFF \sreg_reg[927]  ( .D(c[927]), .CLK(clk), .RST(rst), .Q(c[923]) );
  DFF \sreg_reg[926]  ( .D(c[926]), .CLK(clk), .RST(rst), .Q(c[922]) );
  DFF \sreg_reg[925]  ( .D(c[925]), .CLK(clk), .RST(rst), .Q(c[921]) );
  DFF \sreg_reg[924]  ( .D(c[924]), .CLK(clk), .RST(rst), .Q(c[920]) );
  DFF \sreg_reg[923]  ( .D(c[923]), .CLK(clk), .RST(rst), .Q(c[919]) );
  DFF \sreg_reg[922]  ( .D(c[922]), .CLK(clk), .RST(rst), .Q(c[918]) );
  DFF \sreg_reg[921]  ( .D(c[921]), .CLK(clk), .RST(rst), .Q(c[917]) );
  DFF \sreg_reg[920]  ( .D(c[920]), .CLK(clk), .RST(rst), .Q(c[916]) );
  DFF \sreg_reg[919]  ( .D(c[919]), .CLK(clk), .RST(rst), .Q(c[915]) );
  DFF \sreg_reg[918]  ( .D(c[918]), .CLK(clk), .RST(rst), .Q(c[914]) );
  DFF \sreg_reg[917]  ( .D(c[917]), .CLK(clk), .RST(rst), .Q(c[913]) );
  DFF \sreg_reg[916]  ( .D(c[916]), .CLK(clk), .RST(rst), .Q(c[912]) );
  DFF \sreg_reg[915]  ( .D(c[915]), .CLK(clk), .RST(rst), .Q(c[911]) );
  DFF \sreg_reg[914]  ( .D(c[914]), .CLK(clk), .RST(rst), .Q(c[910]) );
  DFF \sreg_reg[913]  ( .D(c[913]), .CLK(clk), .RST(rst), .Q(c[909]) );
  DFF \sreg_reg[912]  ( .D(c[912]), .CLK(clk), .RST(rst), .Q(c[908]) );
  DFF \sreg_reg[911]  ( .D(c[911]), .CLK(clk), .RST(rst), .Q(c[907]) );
  DFF \sreg_reg[910]  ( .D(c[910]), .CLK(clk), .RST(rst), .Q(c[906]) );
  DFF \sreg_reg[909]  ( .D(c[909]), .CLK(clk), .RST(rst), .Q(c[905]) );
  DFF \sreg_reg[908]  ( .D(c[908]), .CLK(clk), .RST(rst), .Q(c[904]) );
  DFF \sreg_reg[907]  ( .D(c[907]), .CLK(clk), .RST(rst), .Q(c[903]) );
  DFF \sreg_reg[906]  ( .D(c[906]), .CLK(clk), .RST(rst), .Q(c[902]) );
  DFF \sreg_reg[905]  ( .D(c[905]), .CLK(clk), .RST(rst), .Q(c[901]) );
  DFF \sreg_reg[904]  ( .D(c[904]), .CLK(clk), .RST(rst), .Q(c[900]) );
  DFF \sreg_reg[903]  ( .D(c[903]), .CLK(clk), .RST(rst), .Q(c[899]) );
  DFF \sreg_reg[902]  ( .D(c[902]), .CLK(clk), .RST(rst), .Q(c[898]) );
  DFF \sreg_reg[901]  ( .D(c[901]), .CLK(clk), .RST(rst), .Q(c[897]) );
  DFF \sreg_reg[900]  ( .D(c[900]), .CLK(clk), .RST(rst), .Q(c[896]) );
  DFF \sreg_reg[899]  ( .D(c[899]), .CLK(clk), .RST(rst), .Q(c[895]) );
  DFF \sreg_reg[898]  ( .D(c[898]), .CLK(clk), .RST(rst), .Q(c[894]) );
  DFF \sreg_reg[897]  ( .D(c[897]), .CLK(clk), .RST(rst), .Q(c[893]) );
  DFF \sreg_reg[896]  ( .D(c[896]), .CLK(clk), .RST(rst), .Q(c[892]) );
  DFF \sreg_reg[895]  ( .D(c[895]), .CLK(clk), .RST(rst), .Q(c[891]) );
  DFF \sreg_reg[894]  ( .D(c[894]), .CLK(clk), .RST(rst), .Q(c[890]) );
  DFF \sreg_reg[893]  ( .D(c[893]), .CLK(clk), .RST(rst), .Q(c[889]) );
  DFF \sreg_reg[892]  ( .D(c[892]), .CLK(clk), .RST(rst), .Q(c[888]) );
  DFF \sreg_reg[891]  ( .D(c[891]), .CLK(clk), .RST(rst), .Q(c[887]) );
  DFF \sreg_reg[890]  ( .D(c[890]), .CLK(clk), .RST(rst), .Q(c[886]) );
  DFF \sreg_reg[889]  ( .D(c[889]), .CLK(clk), .RST(rst), .Q(c[885]) );
  DFF \sreg_reg[888]  ( .D(c[888]), .CLK(clk), .RST(rst), .Q(c[884]) );
  DFF \sreg_reg[887]  ( .D(c[887]), .CLK(clk), .RST(rst), .Q(c[883]) );
  DFF \sreg_reg[886]  ( .D(c[886]), .CLK(clk), .RST(rst), .Q(c[882]) );
  DFF \sreg_reg[885]  ( .D(c[885]), .CLK(clk), .RST(rst), .Q(c[881]) );
  DFF \sreg_reg[884]  ( .D(c[884]), .CLK(clk), .RST(rst), .Q(c[880]) );
  DFF \sreg_reg[883]  ( .D(c[883]), .CLK(clk), .RST(rst), .Q(c[879]) );
  DFF \sreg_reg[882]  ( .D(c[882]), .CLK(clk), .RST(rst), .Q(c[878]) );
  DFF \sreg_reg[881]  ( .D(c[881]), .CLK(clk), .RST(rst), .Q(c[877]) );
  DFF \sreg_reg[880]  ( .D(c[880]), .CLK(clk), .RST(rst), .Q(c[876]) );
  DFF \sreg_reg[879]  ( .D(c[879]), .CLK(clk), .RST(rst), .Q(c[875]) );
  DFF \sreg_reg[878]  ( .D(c[878]), .CLK(clk), .RST(rst), .Q(c[874]) );
  DFF \sreg_reg[877]  ( .D(c[877]), .CLK(clk), .RST(rst), .Q(c[873]) );
  DFF \sreg_reg[876]  ( .D(c[876]), .CLK(clk), .RST(rst), .Q(c[872]) );
  DFF \sreg_reg[875]  ( .D(c[875]), .CLK(clk), .RST(rst), .Q(c[871]) );
  DFF \sreg_reg[874]  ( .D(c[874]), .CLK(clk), .RST(rst), .Q(c[870]) );
  DFF \sreg_reg[873]  ( .D(c[873]), .CLK(clk), .RST(rst), .Q(c[869]) );
  DFF \sreg_reg[872]  ( .D(c[872]), .CLK(clk), .RST(rst), .Q(c[868]) );
  DFF \sreg_reg[871]  ( .D(c[871]), .CLK(clk), .RST(rst), .Q(c[867]) );
  DFF \sreg_reg[870]  ( .D(c[870]), .CLK(clk), .RST(rst), .Q(c[866]) );
  DFF \sreg_reg[869]  ( .D(c[869]), .CLK(clk), .RST(rst), .Q(c[865]) );
  DFF \sreg_reg[868]  ( .D(c[868]), .CLK(clk), .RST(rst), .Q(c[864]) );
  DFF \sreg_reg[867]  ( .D(c[867]), .CLK(clk), .RST(rst), .Q(c[863]) );
  DFF \sreg_reg[866]  ( .D(c[866]), .CLK(clk), .RST(rst), .Q(c[862]) );
  DFF \sreg_reg[865]  ( .D(c[865]), .CLK(clk), .RST(rst), .Q(c[861]) );
  DFF \sreg_reg[864]  ( .D(c[864]), .CLK(clk), .RST(rst), .Q(c[860]) );
  DFF \sreg_reg[863]  ( .D(c[863]), .CLK(clk), .RST(rst), .Q(c[859]) );
  DFF \sreg_reg[862]  ( .D(c[862]), .CLK(clk), .RST(rst), .Q(c[858]) );
  DFF \sreg_reg[861]  ( .D(c[861]), .CLK(clk), .RST(rst), .Q(c[857]) );
  DFF \sreg_reg[860]  ( .D(c[860]), .CLK(clk), .RST(rst), .Q(c[856]) );
  DFF \sreg_reg[859]  ( .D(c[859]), .CLK(clk), .RST(rst), .Q(c[855]) );
  DFF \sreg_reg[858]  ( .D(c[858]), .CLK(clk), .RST(rst), .Q(c[854]) );
  DFF \sreg_reg[857]  ( .D(c[857]), .CLK(clk), .RST(rst), .Q(c[853]) );
  DFF \sreg_reg[856]  ( .D(c[856]), .CLK(clk), .RST(rst), .Q(c[852]) );
  DFF \sreg_reg[855]  ( .D(c[855]), .CLK(clk), .RST(rst), .Q(c[851]) );
  DFF \sreg_reg[854]  ( .D(c[854]), .CLK(clk), .RST(rst), .Q(c[850]) );
  DFF \sreg_reg[853]  ( .D(c[853]), .CLK(clk), .RST(rst), .Q(c[849]) );
  DFF \sreg_reg[852]  ( .D(c[852]), .CLK(clk), .RST(rst), .Q(c[848]) );
  DFF \sreg_reg[851]  ( .D(c[851]), .CLK(clk), .RST(rst), .Q(c[847]) );
  DFF \sreg_reg[850]  ( .D(c[850]), .CLK(clk), .RST(rst), .Q(c[846]) );
  DFF \sreg_reg[849]  ( .D(c[849]), .CLK(clk), .RST(rst), .Q(c[845]) );
  DFF \sreg_reg[848]  ( .D(c[848]), .CLK(clk), .RST(rst), .Q(c[844]) );
  DFF \sreg_reg[847]  ( .D(c[847]), .CLK(clk), .RST(rst), .Q(c[843]) );
  DFF \sreg_reg[846]  ( .D(c[846]), .CLK(clk), .RST(rst), .Q(c[842]) );
  DFF \sreg_reg[845]  ( .D(c[845]), .CLK(clk), .RST(rst), .Q(c[841]) );
  DFF \sreg_reg[844]  ( .D(c[844]), .CLK(clk), .RST(rst), .Q(c[840]) );
  DFF \sreg_reg[843]  ( .D(c[843]), .CLK(clk), .RST(rst), .Q(c[839]) );
  DFF \sreg_reg[842]  ( .D(c[842]), .CLK(clk), .RST(rst), .Q(c[838]) );
  DFF \sreg_reg[841]  ( .D(c[841]), .CLK(clk), .RST(rst), .Q(c[837]) );
  DFF \sreg_reg[840]  ( .D(c[840]), .CLK(clk), .RST(rst), .Q(c[836]) );
  DFF \sreg_reg[839]  ( .D(c[839]), .CLK(clk), .RST(rst), .Q(c[835]) );
  DFF \sreg_reg[838]  ( .D(c[838]), .CLK(clk), .RST(rst), .Q(c[834]) );
  DFF \sreg_reg[837]  ( .D(c[837]), .CLK(clk), .RST(rst), .Q(c[833]) );
  DFF \sreg_reg[836]  ( .D(c[836]), .CLK(clk), .RST(rst), .Q(c[832]) );
  DFF \sreg_reg[835]  ( .D(c[835]), .CLK(clk), .RST(rst), .Q(c[831]) );
  DFF \sreg_reg[834]  ( .D(c[834]), .CLK(clk), .RST(rst), .Q(c[830]) );
  DFF \sreg_reg[833]  ( .D(c[833]), .CLK(clk), .RST(rst), .Q(c[829]) );
  DFF \sreg_reg[832]  ( .D(c[832]), .CLK(clk), .RST(rst), .Q(c[828]) );
  DFF \sreg_reg[831]  ( .D(c[831]), .CLK(clk), .RST(rst), .Q(c[827]) );
  DFF \sreg_reg[830]  ( .D(c[830]), .CLK(clk), .RST(rst), .Q(c[826]) );
  DFF \sreg_reg[829]  ( .D(c[829]), .CLK(clk), .RST(rst), .Q(c[825]) );
  DFF \sreg_reg[828]  ( .D(c[828]), .CLK(clk), .RST(rst), .Q(c[824]) );
  DFF \sreg_reg[827]  ( .D(c[827]), .CLK(clk), .RST(rst), .Q(c[823]) );
  DFF \sreg_reg[826]  ( .D(c[826]), .CLK(clk), .RST(rst), .Q(c[822]) );
  DFF \sreg_reg[825]  ( .D(c[825]), .CLK(clk), .RST(rst), .Q(c[821]) );
  DFF \sreg_reg[824]  ( .D(c[824]), .CLK(clk), .RST(rst), .Q(c[820]) );
  DFF \sreg_reg[823]  ( .D(c[823]), .CLK(clk), .RST(rst), .Q(c[819]) );
  DFF \sreg_reg[822]  ( .D(c[822]), .CLK(clk), .RST(rst), .Q(c[818]) );
  DFF \sreg_reg[821]  ( .D(c[821]), .CLK(clk), .RST(rst), .Q(c[817]) );
  DFF \sreg_reg[820]  ( .D(c[820]), .CLK(clk), .RST(rst), .Q(c[816]) );
  DFF \sreg_reg[819]  ( .D(c[819]), .CLK(clk), .RST(rst), .Q(c[815]) );
  DFF \sreg_reg[818]  ( .D(c[818]), .CLK(clk), .RST(rst), .Q(c[814]) );
  DFF \sreg_reg[817]  ( .D(c[817]), .CLK(clk), .RST(rst), .Q(c[813]) );
  DFF \sreg_reg[816]  ( .D(c[816]), .CLK(clk), .RST(rst), .Q(c[812]) );
  DFF \sreg_reg[815]  ( .D(c[815]), .CLK(clk), .RST(rst), .Q(c[811]) );
  DFF \sreg_reg[814]  ( .D(c[814]), .CLK(clk), .RST(rst), .Q(c[810]) );
  DFF \sreg_reg[813]  ( .D(c[813]), .CLK(clk), .RST(rst), .Q(c[809]) );
  DFF \sreg_reg[812]  ( .D(c[812]), .CLK(clk), .RST(rst), .Q(c[808]) );
  DFF \sreg_reg[811]  ( .D(c[811]), .CLK(clk), .RST(rst), .Q(c[807]) );
  DFF \sreg_reg[810]  ( .D(c[810]), .CLK(clk), .RST(rst), .Q(c[806]) );
  DFF \sreg_reg[809]  ( .D(c[809]), .CLK(clk), .RST(rst), .Q(c[805]) );
  DFF \sreg_reg[808]  ( .D(c[808]), .CLK(clk), .RST(rst), .Q(c[804]) );
  DFF \sreg_reg[807]  ( .D(c[807]), .CLK(clk), .RST(rst), .Q(c[803]) );
  DFF \sreg_reg[806]  ( .D(c[806]), .CLK(clk), .RST(rst), .Q(c[802]) );
  DFF \sreg_reg[805]  ( .D(c[805]), .CLK(clk), .RST(rst), .Q(c[801]) );
  DFF \sreg_reg[804]  ( .D(c[804]), .CLK(clk), .RST(rst), .Q(c[800]) );
  DFF \sreg_reg[803]  ( .D(c[803]), .CLK(clk), .RST(rst), .Q(c[799]) );
  DFF \sreg_reg[802]  ( .D(c[802]), .CLK(clk), .RST(rst), .Q(c[798]) );
  DFF \sreg_reg[801]  ( .D(c[801]), .CLK(clk), .RST(rst), .Q(c[797]) );
  DFF \sreg_reg[800]  ( .D(c[800]), .CLK(clk), .RST(rst), .Q(c[796]) );
  DFF \sreg_reg[799]  ( .D(c[799]), .CLK(clk), .RST(rst), .Q(c[795]) );
  DFF \sreg_reg[798]  ( .D(c[798]), .CLK(clk), .RST(rst), .Q(c[794]) );
  DFF \sreg_reg[797]  ( .D(c[797]), .CLK(clk), .RST(rst), .Q(c[793]) );
  DFF \sreg_reg[796]  ( .D(c[796]), .CLK(clk), .RST(rst), .Q(c[792]) );
  DFF \sreg_reg[795]  ( .D(c[795]), .CLK(clk), .RST(rst), .Q(c[791]) );
  DFF \sreg_reg[794]  ( .D(c[794]), .CLK(clk), .RST(rst), .Q(c[790]) );
  DFF \sreg_reg[793]  ( .D(c[793]), .CLK(clk), .RST(rst), .Q(c[789]) );
  DFF \sreg_reg[792]  ( .D(c[792]), .CLK(clk), .RST(rst), .Q(c[788]) );
  DFF \sreg_reg[791]  ( .D(c[791]), .CLK(clk), .RST(rst), .Q(c[787]) );
  DFF \sreg_reg[790]  ( .D(c[790]), .CLK(clk), .RST(rst), .Q(c[786]) );
  DFF \sreg_reg[789]  ( .D(c[789]), .CLK(clk), .RST(rst), .Q(c[785]) );
  DFF \sreg_reg[788]  ( .D(c[788]), .CLK(clk), .RST(rst), .Q(c[784]) );
  DFF \sreg_reg[787]  ( .D(c[787]), .CLK(clk), .RST(rst), .Q(c[783]) );
  DFF \sreg_reg[786]  ( .D(c[786]), .CLK(clk), .RST(rst), .Q(c[782]) );
  DFF \sreg_reg[785]  ( .D(c[785]), .CLK(clk), .RST(rst), .Q(c[781]) );
  DFF \sreg_reg[784]  ( .D(c[784]), .CLK(clk), .RST(rst), .Q(c[780]) );
  DFF \sreg_reg[783]  ( .D(c[783]), .CLK(clk), .RST(rst), .Q(c[779]) );
  DFF \sreg_reg[782]  ( .D(c[782]), .CLK(clk), .RST(rst), .Q(c[778]) );
  DFF \sreg_reg[781]  ( .D(c[781]), .CLK(clk), .RST(rst), .Q(c[777]) );
  DFF \sreg_reg[780]  ( .D(c[780]), .CLK(clk), .RST(rst), .Q(c[776]) );
  DFF \sreg_reg[779]  ( .D(c[779]), .CLK(clk), .RST(rst), .Q(c[775]) );
  DFF \sreg_reg[778]  ( .D(c[778]), .CLK(clk), .RST(rst), .Q(c[774]) );
  DFF \sreg_reg[777]  ( .D(c[777]), .CLK(clk), .RST(rst), .Q(c[773]) );
  DFF \sreg_reg[776]  ( .D(c[776]), .CLK(clk), .RST(rst), .Q(c[772]) );
  DFF \sreg_reg[775]  ( .D(c[775]), .CLK(clk), .RST(rst), .Q(c[771]) );
  DFF \sreg_reg[774]  ( .D(c[774]), .CLK(clk), .RST(rst), .Q(c[770]) );
  DFF \sreg_reg[773]  ( .D(c[773]), .CLK(clk), .RST(rst), .Q(c[769]) );
  DFF \sreg_reg[772]  ( .D(c[772]), .CLK(clk), .RST(rst), .Q(c[768]) );
  DFF \sreg_reg[771]  ( .D(c[771]), .CLK(clk), .RST(rst), .Q(c[767]) );
  DFF \sreg_reg[770]  ( .D(c[770]), .CLK(clk), .RST(rst), .Q(c[766]) );
  DFF \sreg_reg[769]  ( .D(c[769]), .CLK(clk), .RST(rst), .Q(c[765]) );
  DFF \sreg_reg[768]  ( .D(c[768]), .CLK(clk), .RST(rst), .Q(c[764]) );
  DFF \sreg_reg[767]  ( .D(c[767]), .CLK(clk), .RST(rst), .Q(c[763]) );
  DFF \sreg_reg[766]  ( .D(c[766]), .CLK(clk), .RST(rst), .Q(c[762]) );
  DFF \sreg_reg[765]  ( .D(c[765]), .CLK(clk), .RST(rst), .Q(c[761]) );
  DFF \sreg_reg[764]  ( .D(c[764]), .CLK(clk), .RST(rst), .Q(c[760]) );
  DFF \sreg_reg[763]  ( .D(c[763]), .CLK(clk), .RST(rst), .Q(c[759]) );
  DFF \sreg_reg[762]  ( .D(c[762]), .CLK(clk), .RST(rst), .Q(c[758]) );
  DFF \sreg_reg[761]  ( .D(c[761]), .CLK(clk), .RST(rst), .Q(c[757]) );
  DFF \sreg_reg[760]  ( .D(c[760]), .CLK(clk), .RST(rst), .Q(c[756]) );
  DFF \sreg_reg[759]  ( .D(c[759]), .CLK(clk), .RST(rst), .Q(c[755]) );
  DFF \sreg_reg[758]  ( .D(c[758]), .CLK(clk), .RST(rst), .Q(c[754]) );
  DFF \sreg_reg[757]  ( .D(c[757]), .CLK(clk), .RST(rst), .Q(c[753]) );
  DFF \sreg_reg[756]  ( .D(c[756]), .CLK(clk), .RST(rst), .Q(c[752]) );
  DFF \sreg_reg[755]  ( .D(c[755]), .CLK(clk), .RST(rst), .Q(c[751]) );
  DFF \sreg_reg[754]  ( .D(c[754]), .CLK(clk), .RST(rst), .Q(c[750]) );
  DFF \sreg_reg[753]  ( .D(c[753]), .CLK(clk), .RST(rst), .Q(c[749]) );
  DFF \sreg_reg[752]  ( .D(c[752]), .CLK(clk), .RST(rst), .Q(c[748]) );
  DFF \sreg_reg[751]  ( .D(c[751]), .CLK(clk), .RST(rst), .Q(c[747]) );
  DFF \sreg_reg[750]  ( .D(c[750]), .CLK(clk), .RST(rst), .Q(c[746]) );
  DFF \sreg_reg[749]  ( .D(c[749]), .CLK(clk), .RST(rst), .Q(c[745]) );
  DFF \sreg_reg[748]  ( .D(c[748]), .CLK(clk), .RST(rst), .Q(c[744]) );
  DFF \sreg_reg[747]  ( .D(c[747]), .CLK(clk), .RST(rst), .Q(c[743]) );
  DFF \sreg_reg[746]  ( .D(c[746]), .CLK(clk), .RST(rst), .Q(c[742]) );
  DFF \sreg_reg[745]  ( .D(c[745]), .CLK(clk), .RST(rst), .Q(c[741]) );
  DFF \sreg_reg[744]  ( .D(c[744]), .CLK(clk), .RST(rst), .Q(c[740]) );
  DFF \sreg_reg[743]  ( .D(c[743]), .CLK(clk), .RST(rst), .Q(c[739]) );
  DFF \sreg_reg[742]  ( .D(c[742]), .CLK(clk), .RST(rst), .Q(c[738]) );
  DFF \sreg_reg[741]  ( .D(c[741]), .CLK(clk), .RST(rst), .Q(c[737]) );
  DFF \sreg_reg[740]  ( .D(c[740]), .CLK(clk), .RST(rst), .Q(c[736]) );
  DFF \sreg_reg[739]  ( .D(c[739]), .CLK(clk), .RST(rst), .Q(c[735]) );
  DFF \sreg_reg[738]  ( .D(c[738]), .CLK(clk), .RST(rst), .Q(c[734]) );
  DFF \sreg_reg[737]  ( .D(c[737]), .CLK(clk), .RST(rst), .Q(c[733]) );
  DFF \sreg_reg[736]  ( .D(c[736]), .CLK(clk), .RST(rst), .Q(c[732]) );
  DFF \sreg_reg[735]  ( .D(c[735]), .CLK(clk), .RST(rst), .Q(c[731]) );
  DFF \sreg_reg[734]  ( .D(c[734]), .CLK(clk), .RST(rst), .Q(c[730]) );
  DFF \sreg_reg[733]  ( .D(c[733]), .CLK(clk), .RST(rst), .Q(c[729]) );
  DFF \sreg_reg[732]  ( .D(c[732]), .CLK(clk), .RST(rst), .Q(c[728]) );
  DFF \sreg_reg[731]  ( .D(c[731]), .CLK(clk), .RST(rst), .Q(c[727]) );
  DFF \sreg_reg[730]  ( .D(c[730]), .CLK(clk), .RST(rst), .Q(c[726]) );
  DFF \sreg_reg[729]  ( .D(c[729]), .CLK(clk), .RST(rst), .Q(c[725]) );
  DFF \sreg_reg[728]  ( .D(c[728]), .CLK(clk), .RST(rst), .Q(c[724]) );
  DFF \sreg_reg[727]  ( .D(c[727]), .CLK(clk), .RST(rst), .Q(c[723]) );
  DFF \sreg_reg[726]  ( .D(c[726]), .CLK(clk), .RST(rst), .Q(c[722]) );
  DFF \sreg_reg[725]  ( .D(c[725]), .CLK(clk), .RST(rst), .Q(c[721]) );
  DFF \sreg_reg[724]  ( .D(c[724]), .CLK(clk), .RST(rst), .Q(c[720]) );
  DFF \sreg_reg[723]  ( .D(c[723]), .CLK(clk), .RST(rst), .Q(c[719]) );
  DFF \sreg_reg[722]  ( .D(c[722]), .CLK(clk), .RST(rst), .Q(c[718]) );
  DFF \sreg_reg[721]  ( .D(c[721]), .CLK(clk), .RST(rst), .Q(c[717]) );
  DFF \sreg_reg[720]  ( .D(c[720]), .CLK(clk), .RST(rst), .Q(c[716]) );
  DFF \sreg_reg[719]  ( .D(c[719]), .CLK(clk), .RST(rst), .Q(c[715]) );
  DFF \sreg_reg[718]  ( .D(c[718]), .CLK(clk), .RST(rst), .Q(c[714]) );
  DFF \sreg_reg[717]  ( .D(c[717]), .CLK(clk), .RST(rst), .Q(c[713]) );
  DFF \sreg_reg[716]  ( .D(c[716]), .CLK(clk), .RST(rst), .Q(c[712]) );
  DFF \sreg_reg[715]  ( .D(c[715]), .CLK(clk), .RST(rst), .Q(c[711]) );
  DFF \sreg_reg[714]  ( .D(c[714]), .CLK(clk), .RST(rst), .Q(c[710]) );
  DFF \sreg_reg[713]  ( .D(c[713]), .CLK(clk), .RST(rst), .Q(c[709]) );
  DFF \sreg_reg[712]  ( .D(c[712]), .CLK(clk), .RST(rst), .Q(c[708]) );
  DFF \sreg_reg[711]  ( .D(c[711]), .CLK(clk), .RST(rst), .Q(c[707]) );
  DFF \sreg_reg[710]  ( .D(c[710]), .CLK(clk), .RST(rst), .Q(c[706]) );
  DFF \sreg_reg[709]  ( .D(c[709]), .CLK(clk), .RST(rst), .Q(c[705]) );
  DFF \sreg_reg[708]  ( .D(c[708]), .CLK(clk), .RST(rst), .Q(c[704]) );
  DFF \sreg_reg[707]  ( .D(c[707]), .CLK(clk), .RST(rst), .Q(c[703]) );
  DFF \sreg_reg[706]  ( .D(c[706]), .CLK(clk), .RST(rst), .Q(c[702]) );
  DFF \sreg_reg[705]  ( .D(c[705]), .CLK(clk), .RST(rst), .Q(c[701]) );
  DFF \sreg_reg[704]  ( .D(c[704]), .CLK(clk), .RST(rst), .Q(c[700]) );
  DFF \sreg_reg[703]  ( .D(c[703]), .CLK(clk), .RST(rst), .Q(c[699]) );
  DFF \sreg_reg[702]  ( .D(c[702]), .CLK(clk), .RST(rst), .Q(c[698]) );
  DFF \sreg_reg[701]  ( .D(c[701]), .CLK(clk), .RST(rst), .Q(c[697]) );
  DFF \sreg_reg[700]  ( .D(c[700]), .CLK(clk), .RST(rst), .Q(c[696]) );
  DFF \sreg_reg[699]  ( .D(c[699]), .CLK(clk), .RST(rst), .Q(c[695]) );
  DFF \sreg_reg[698]  ( .D(c[698]), .CLK(clk), .RST(rst), .Q(c[694]) );
  DFF \sreg_reg[697]  ( .D(c[697]), .CLK(clk), .RST(rst), .Q(c[693]) );
  DFF \sreg_reg[696]  ( .D(c[696]), .CLK(clk), .RST(rst), .Q(c[692]) );
  DFF \sreg_reg[695]  ( .D(c[695]), .CLK(clk), .RST(rst), .Q(c[691]) );
  DFF \sreg_reg[694]  ( .D(c[694]), .CLK(clk), .RST(rst), .Q(c[690]) );
  DFF \sreg_reg[693]  ( .D(c[693]), .CLK(clk), .RST(rst), .Q(c[689]) );
  DFF \sreg_reg[692]  ( .D(c[692]), .CLK(clk), .RST(rst), .Q(c[688]) );
  DFF \sreg_reg[691]  ( .D(c[691]), .CLK(clk), .RST(rst), .Q(c[687]) );
  DFF \sreg_reg[690]  ( .D(c[690]), .CLK(clk), .RST(rst), .Q(c[686]) );
  DFF \sreg_reg[689]  ( .D(c[689]), .CLK(clk), .RST(rst), .Q(c[685]) );
  DFF \sreg_reg[688]  ( .D(c[688]), .CLK(clk), .RST(rst), .Q(c[684]) );
  DFF \sreg_reg[687]  ( .D(c[687]), .CLK(clk), .RST(rst), .Q(c[683]) );
  DFF \sreg_reg[686]  ( .D(c[686]), .CLK(clk), .RST(rst), .Q(c[682]) );
  DFF \sreg_reg[685]  ( .D(c[685]), .CLK(clk), .RST(rst), .Q(c[681]) );
  DFF \sreg_reg[684]  ( .D(c[684]), .CLK(clk), .RST(rst), .Q(c[680]) );
  DFF \sreg_reg[683]  ( .D(c[683]), .CLK(clk), .RST(rst), .Q(c[679]) );
  DFF \sreg_reg[682]  ( .D(c[682]), .CLK(clk), .RST(rst), .Q(c[678]) );
  DFF \sreg_reg[681]  ( .D(c[681]), .CLK(clk), .RST(rst), .Q(c[677]) );
  DFF \sreg_reg[680]  ( .D(c[680]), .CLK(clk), .RST(rst), .Q(c[676]) );
  DFF \sreg_reg[679]  ( .D(c[679]), .CLK(clk), .RST(rst), .Q(c[675]) );
  DFF \sreg_reg[678]  ( .D(c[678]), .CLK(clk), .RST(rst), .Q(c[674]) );
  DFF \sreg_reg[677]  ( .D(c[677]), .CLK(clk), .RST(rst), .Q(c[673]) );
  DFF \sreg_reg[676]  ( .D(c[676]), .CLK(clk), .RST(rst), .Q(c[672]) );
  DFF \sreg_reg[675]  ( .D(c[675]), .CLK(clk), .RST(rst), .Q(c[671]) );
  DFF \sreg_reg[674]  ( .D(c[674]), .CLK(clk), .RST(rst), .Q(c[670]) );
  DFF \sreg_reg[673]  ( .D(c[673]), .CLK(clk), .RST(rst), .Q(c[669]) );
  DFF \sreg_reg[672]  ( .D(c[672]), .CLK(clk), .RST(rst), .Q(c[668]) );
  DFF \sreg_reg[671]  ( .D(c[671]), .CLK(clk), .RST(rst), .Q(c[667]) );
  DFF \sreg_reg[670]  ( .D(c[670]), .CLK(clk), .RST(rst), .Q(c[666]) );
  DFF \sreg_reg[669]  ( .D(c[669]), .CLK(clk), .RST(rst), .Q(c[665]) );
  DFF \sreg_reg[668]  ( .D(c[668]), .CLK(clk), .RST(rst), .Q(c[664]) );
  DFF \sreg_reg[667]  ( .D(c[667]), .CLK(clk), .RST(rst), .Q(c[663]) );
  DFF \sreg_reg[666]  ( .D(c[666]), .CLK(clk), .RST(rst), .Q(c[662]) );
  DFF \sreg_reg[665]  ( .D(c[665]), .CLK(clk), .RST(rst), .Q(c[661]) );
  DFF \sreg_reg[664]  ( .D(c[664]), .CLK(clk), .RST(rst), .Q(c[660]) );
  DFF \sreg_reg[663]  ( .D(c[663]), .CLK(clk), .RST(rst), .Q(c[659]) );
  DFF \sreg_reg[662]  ( .D(c[662]), .CLK(clk), .RST(rst), .Q(c[658]) );
  DFF \sreg_reg[661]  ( .D(c[661]), .CLK(clk), .RST(rst), .Q(c[657]) );
  DFF \sreg_reg[660]  ( .D(c[660]), .CLK(clk), .RST(rst), .Q(c[656]) );
  DFF \sreg_reg[659]  ( .D(c[659]), .CLK(clk), .RST(rst), .Q(c[655]) );
  DFF \sreg_reg[658]  ( .D(c[658]), .CLK(clk), .RST(rst), .Q(c[654]) );
  DFF \sreg_reg[657]  ( .D(c[657]), .CLK(clk), .RST(rst), .Q(c[653]) );
  DFF \sreg_reg[656]  ( .D(c[656]), .CLK(clk), .RST(rst), .Q(c[652]) );
  DFF \sreg_reg[655]  ( .D(c[655]), .CLK(clk), .RST(rst), .Q(c[651]) );
  DFF \sreg_reg[654]  ( .D(c[654]), .CLK(clk), .RST(rst), .Q(c[650]) );
  DFF \sreg_reg[653]  ( .D(c[653]), .CLK(clk), .RST(rst), .Q(c[649]) );
  DFF \sreg_reg[652]  ( .D(c[652]), .CLK(clk), .RST(rst), .Q(c[648]) );
  DFF \sreg_reg[651]  ( .D(c[651]), .CLK(clk), .RST(rst), .Q(c[647]) );
  DFF \sreg_reg[650]  ( .D(c[650]), .CLK(clk), .RST(rst), .Q(c[646]) );
  DFF \sreg_reg[649]  ( .D(c[649]), .CLK(clk), .RST(rst), .Q(c[645]) );
  DFF \sreg_reg[648]  ( .D(c[648]), .CLK(clk), .RST(rst), .Q(c[644]) );
  DFF \sreg_reg[647]  ( .D(c[647]), .CLK(clk), .RST(rst), .Q(c[643]) );
  DFF \sreg_reg[646]  ( .D(c[646]), .CLK(clk), .RST(rst), .Q(c[642]) );
  DFF \sreg_reg[645]  ( .D(c[645]), .CLK(clk), .RST(rst), .Q(c[641]) );
  DFF \sreg_reg[644]  ( .D(c[644]), .CLK(clk), .RST(rst), .Q(c[640]) );
  DFF \sreg_reg[643]  ( .D(c[643]), .CLK(clk), .RST(rst), .Q(c[639]) );
  DFF \sreg_reg[642]  ( .D(c[642]), .CLK(clk), .RST(rst), .Q(c[638]) );
  DFF \sreg_reg[641]  ( .D(c[641]), .CLK(clk), .RST(rst), .Q(c[637]) );
  DFF \sreg_reg[640]  ( .D(c[640]), .CLK(clk), .RST(rst), .Q(c[636]) );
  DFF \sreg_reg[639]  ( .D(c[639]), .CLK(clk), .RST(rst), .Q(c[635]) );
  DFF \sreg_reg[638]  ( .D(c[638]), .CLK(clk), .RST(rst), .Q(c[634]) );
  DFF \sreg_reg[637]  ( .D(c[637]), .CLK(clk), .RST(rst), .Q(c[633]) );
  DFF \sreg_reg[636]  ( .D(c[636]), .CLK(clk), .RST(rst), .Q(c[632]) );
  DFF \sreg_reg[635]  ( .D(c[635]), .CLK(clk), .RST(rst), .Q(c[631]) );
  DFF \sreg_reg[634]  ( .D(c[634]), .CLK(clk), .RST(rst), .Q(c[630]) );
  DFF \sreg_reg[633]  ( .D(c[633]), .CLK(clk), .RST(rst), .Q(c[629]) );
  DFF \sreg_reg[632]  ( .D(c[632]), .CLK(clk), .RST(rst), .Q(c[628]) );
  DFF \sreg_reg[631]  ( .D(c[631]), .CLK(clk), .RST(rst), .Q(c[627]) );
  DFF \sreg_reg[630]  ( .D(c[630]), .CLK(clk), .RST(rst), .Q(c[626]) );
  DFF \sreg_reg[629]  ( .D(c[629]), .CLK(clk), .RST(rst), .Q(c[625]) );
  DFF \sreg_reg[628]  ( .D(c[628]), .CLK(clk), .RST(rst), .Q(c[624]) );
  DFF \sreg_reg[627]  ( .D(c[627]), .CLK(clk), .RST(rst), .Q(c[623]) );
  DFF \sreg_reg[626]  ( .D(c[626]), .CLK(clk), .RST(rst), .Q(c[622]) );
  DFF \sreg_reg[625]  ( .D(c[625]), .CLK(clk), .RST(rst), .Q(c[621]) );
  DFF \sreg_reg[624]  ( .D(c[624]), .CLK(clk), .RST(rst), .Q(c[620]) );
  DFF \sreg_reg[623]  ( .D(c[623]), .CLK(clk), .RST(rst), .Q(c[619]) );
  DFF \sreg_reg[622]  ( .D(c[622]), .CLK(clk), .RST(rst), .Q(c[618]) );
  DFF \sreg_reg[621]  ( .D(c[621]), .CLK(clk), .RST(rst), .Q(c[617]) );
  DFF \sreg_reg[620]  ( .D(c[620]), .CLK(clk), .RST(rst), .Q(c[616]) );
  DFF \sreg_reg[619]  ( .D(c[619]), .CLK(clk), .RST(rst), .Q(c[615]) );
  DFF \sreg_reg[618]  ( .D(c[618]), .CLK(clk), .RST(rst), .Q(c[614]) );
  DFF \sreg_reg[617]  ( .D(c[617]), .CLK(clk), .RST(rst), .Q(c[613]) );
  DFF \sreg_reg[616]  ( .D(c[616]), .CLK(clk), .RST(rst), .Q(c[612]) );
  DFF \sreg_reg[615]  ( .D(c[615]), .CLK(clk), .RST(rst), .Q(c[611]) );
  DFF \sreg_reg[614]  ( .D(c[614]), .CLK(clk), .RST(rst), .Q(c[610]) );
  DFF \sreg_reg[613]  ( .D(c[613]), .CLK(clk), .RST(rst), .Q(c[609]) );
  DFF \sreg_reg[612]  ( .D(c[612]), .CLK(clk), .RST(rst), .Q(c[608]) );
  DFF \sreg_reg[611]  ( .D(c[611]), .CLK(clk), .RST(rst), .Q(c[607]) );
  DFF \sreg_reg[610]  ( .D(c[610]), .CLK(clk), .RST(rst), .Q(c[606]) );
  DFF \sreg_reg[609]  ( .D(c[609]), .CLK(clk), .RST(rst), .Q(c[605]) );
  DFF \sreg_reg[608]  ( .D(c[608]), .CLK(clk), .RST(rst), .Q(c[604]) );
  DFF \sreg_reg[607]  ( .D(c[607]), .CLK(clk), .RST(rst), .Q(c[603]) );
  DFF \sreg_reg[606]  ( .D(c[606]), .CLK(clk), .RST(rst), .Q(c[602]) );
  DFF \sreg_reg[605]  ( .D(c[605]), .CLK(clk), .RST(rst), .Q(c[601]) );
  DFF \sreg_reg[604]  ( .D(c[604]), .CLK(clk), .RST(rst), .Q(c[600]) );
  DFF \sreg_reg[603]  ( .D(c[603]), .CLK(clk), .RST(rst), .Q(c[599]) );
  DFF \sreg_reg[602]  ( .D(c[602]), .CLK(clk), .RST(rst), .Q(c[598]) );
  DFF \sreg_reg[601]  ( .D(c[601]), .CLK(clk), .RST(rst), .Q(c[597]) );
  DFF \sreg_reg[600]  ( .D(c[600]), .CLK(clk), .RST(rst), .Q(c[596]) );
  DFF \sreg_reg[599]  ( .D(c[599]), .CLK(clk), .RST(rst), .Q(c[595]) );
  DFF \sreg_reg[598]  ( .D(c[598]), .CLK(clk), .RST(rst), .Q(c[594]) );
  DFF \sreg_reg[597]  ( .D(c[597]), .CLK(clk), .RST(rst), .Q(c[593]) );
  DFF \sreg_reg[596]  ( .D(c[596]), .CLK(clk), .RST(rst), .Q(c[592]) );
  DFF \sreg_reg[595]  ( .D(c[595]), .CLK(clk), .RST(rst), .Q(c[591]) );
  DFF \sreg_reg[594]  ( .D(c[594]), .CLK(clk), .RST(rst), .Q(c[590]) );
  DFF \sreg_reg[593]  ( .D(c[593]), .CLK(clk), .RST(rst), .Q(c[589]) );
  DFF \sreg_reg[592]  ( .D(c[592]), .CLK(clk), .RST(rst), .Q(c[588]) );
  DFF \sreg_reg[591]  ( .D(c[591]), .CLK(clk), .RST(rst), .Q(c[587]) );
  DFF \sreg_reg[590]  ( .D(c[590]), .CLK(clk), .RST(rst), .Q(c[586]) );
  DFF \sreg_reg[589]  ( .D(c[589]), .CLK(clk), .RST(rst), .Q(c[585]) );
  DFF \sreg_reg[588]  ( .D(c[588]), .CLK(clk), .RST(rst), .Q(c[584]) );
  DFF \sreg_reg[587]  ( .D(c[587]), .CLK(clk), .RST(rst), .Q(c[583]) );
  DFF \sreg_reg[586]  ( .D(c[586]), .CLK(clk), .RST(rst), .Q(c[582]) );
  DFF \sreg_reg[585]  ( .D(c[585]), .CLK(clk), .RST(rst), .Q(c[581]) );
  DFF \sreg_reg[584]  ( .D(c[584]), .CLK(clk), .RST(rst), .Q(c[580]) );
  DFF \sreg_reg[583]  ( .D(c[583]), .CLK(clk), .RST(rst), .Q(c[579]) );
  DFF \sreg_reg[582]  ( .D(c[582]), .CLK(clk), .RST(rst), .Q(c[578]) );
  DFF \sreg_reg[581]  ( .D(c[581]), .CLK(clk), .RST(rst), .Q(c[577]) );
  DFF \sreg_reg[580]  ( .D(c[580]), .CLK(clk), .RST(rst), .Q(c[576]) );
  DFF \sreg_reg[579]  ( .D(c[579]), .CLK(clk), .RST(rst), .Q(c[575]) );
  DFF \sreg_reg[578]  ( .D(c[578]), .CLK(clk), .RST(rst), .Q(c[574]) );
  DFF \sreg_reg[577]  ( .D(c[577]), .CLK(clk), .RST(rst), .Q(c[573]) );
  DFF \sreg_reg[576]  ( .D(c[576]), .CLK(clk), .RST(rst), .Q(c[572]) );
  DFF \sreg_reg[575]  ( .D(c[575]), .CLK(clk), .RST(rst), .Q(c[571]) );
  DFF \sreg_reg[574]  ( .D(c[574]), .CLK(clk), .RST(rst), .Q(c[570]) );
  DFF \sreg_reg[573]  ( .D(c[573]), .CLK(clk), .RST(rst), .Q(c[569]) );
  DFF \sreg_reg[572]  ( .D(c[572]), .CLK(clk), .RST(rst), .Q(c[568]) );
  DFF \sreg_reg[571]  ( .D(c[571]), .CLK(clk), .RST(rst), .Q(c[567]) );
  DFF \sreg_reg[570]  ( .D(c[570]), .CLK(clk), .RST(rst), .Q(c[566]) );
  DFF \sreg_reg[569]  ( .D(c[569]), .CLK(clk), .RST(rst), .Q(c[565]) );
  DFF \sreg_reg[568]  ( .D(c[568]), .CLK(clk), .RST(rst), .Q(c[564]) );
  DFF \sreg_reg[567]  ( .D(c[567]), .CLK(clk), .RST(rst), .Q(c[563]) );
  DFF \sreg_reg[566]  ( .D(c[566]), .CLK(clk), .RST(rst), .Q(c[562]) );
  DFF \sreg_reg[565]  ( .D(c[565]), .CLK(clk), .RST(rst), .Q(c[561]) );
  DFF \sreg_reg[564]  ( .D(c[564]), .CLK(clk), .RST(rst), .Q(c[560]) );
  DFF \sreg_reg[563]  ( .D(c[563]), .CLK(clk), .RST(rst), .Q(c[559]) );
  DFF \sreg_reg[562]  ( .D(c[562]), .CLK(clk), .RST(rst), .Q(c[558]) );
  DFF \sreg_reg[561]  ( .D(c[561]), .CLK(clk), .RST(rst), .Q(c[557]) );
  DFF \sreg_reg[560]  ( .D(c[560]), .CLK(clk), .RST(rst), .Q(c[556]) );
  DFF \sreg_reg[559]  ( .D(c[559]), .CLK(clk), .RST(rst), .Q(c[555]) );
  DFF \sreg_reg[558]  ( .D(c[558]), .CLK(clk), .RST(rst), .Q(c[554]) );
  DFF \sreg_reg[557]  ( .D(c[557]), .CLK(clk), .RST(rst), .Q(c[553]) );
  DFF \sreg_reg[556]  ( .D(c[556]), .CLK(clk), .RST(rst), .Q(c[552]) );
  DFF \sreg_reg[555]  ( .D(c[555]), .CLK(clk), .RST(rst), .Q(c[551]) );
  DFF \sreg_reg[554]  ( .D(c[554]), .CLK(clk), .RST(rst), .Q(c[550]) );
  DFF \sreg_reg[553]  ( .D(c[553]), .CLK(clk), .RST(rst), .Q(c[549]) );
  DFF \sreg_reg[552]  ( .D(c[552]), .CLK(clk), .RST(rst), .Q(c[548]) );
  DFF \sreg_reg[551]  ( .D(c[551]), .CLK(clk), .RST(rst), .Q(c[547]) );
  DFF \sreg_reg[550]  ( .D(c[550]), .CLK(clk), .RST(rst), .Q(c[546]) );
  DFF \sreg_reg[549]  ( .D(c[549]), .CLK(clk), .RST(rst), .Q(c[545]) );
  DFF \sreg_reg[548]  ( .D(c[548]), .CLK(clk), .RST(rst), .Q(c[544]) );
  DFF \sreg_reg[547]  ( .D(c[547]), .CLK(clk), .RST(rst), .Q(c[543]) );
  DFF \sreg_reg[546]  ( .D(c[546]), .CLK(clk), .RST(rst), .Q(c[542]) );
  DFF \sreg_reg[545]  ( .D(c[545]), .CLK(clk), .RST(rst), .Q(c[541]) );
  DFF \sreg_reg[544]  ( .D(c[544]), .CLK(clk), .RST(rst), .Q(c[540]) );
  DFF \sreg_reg[543]  ( .D(c[543]), .CLK(clk), .RST(rst), .Q(c[539]) );
  DFF \sreg_reg[542]  ( .D(c[542]), .CLK(clk), .RST(rst), .Q(c[538]) );
  DFF \sreg_reg[541]  ( .D(c[541]), .CLK(clk), .RST(rst), .Q(c[537]) );
  DFF \sreg_reg[540]  ( .D(c[540]), .CLK(clk), .RST(rst), .Q(c[536]) );
  DFF \sreg_reg[539]  ( .D(c[539]), .CLK(clk), .RST(rst), .Q(c[535]) );
  DFF \sreg_reg[538]  ( .D(c[538]), .CLK(clk), .RST(rst), .Q(c[534]) );
  DFF \sreg_reg[537]  ( .D(c[537]), .CLK(clk), .RST(rst), .Q(c[533]) );
  DFF \sreg_reg[536]  ( .D(c[536]), .CLK(clk), .RST(rst), .Q(c[532]) );
  DFF \sreg_reg[535]  ( .D(c[535]), .CLK(clk), .RST(rst), .Q(c[531]) );
  DFF \sreg_reg[534]  ( .D(c[534]), .CLK(clk), .RST(rst), .Q(c[530]) );
  DFF \sreg_reg[533]  ( .D(c[533]), .CLK(clk), .RST(rst), .Q(c[529]) );
  DFF \sreg_reg[532]  ( .D(c[532]), .CLK(clk), .RST(rst), .Q(c[528]) );
  DFF \sreg_reg[531]  ( .D(c[531]), .CLK(clk), .RST(rst), .Q(c[527]) );
  DFF \sreg_reg[530]  ( .D(c[530]), .CLK(clk), .RST(rst), .Q(c[526]) );
  DFF \sreg_reg[529]  ( .D(c[529]), .CLK(clk), .RST(rst), .Q(c[525]) );
  DFF \sreg_reg[528]  ( .D(c[528]), .CLK(clk), .RST(rst), .Q(c[524]) );
  DFF \sreg_reg[527]  ( .D(c[527]), .CLK(clk), .RST(rst), .Q(c[523]) );
  DFF \sreg_reg[526]  ( .D(c[526]), .CLK(clk), .RST(rst), .Q(c[522]) );
  DFF \sreg_reg[525]  ( .D(c[525]), .CLK(clk), .RST(rst), .Q(c[521]) );
  DFF \sreg_reg[524]  ( .D(c[524]), .CLK(clk), .RST(rst), .Q(c[520]) );
  DFF \sreg_reg[523]  ( .D(c[523]), .CLK(clk), .RST(rst), .Q(c[519]) );
  DFF \sreg_reg[522]  ( .D(c[522]), .CLK(clk), .RST(rst), .Q(c[518]) );
  DFF \sreg_reg[521]  ( .D(c[521]), .CLK(clk), .RST(rst), .Q(c[517]) );
  DFF \sreg_reg[520]  ( .D(c[520]), .CLK(clk), .RST(rst), .Q(c[516]) );
  DFF \sreg_reg[519]  ( .D(c[519]), .CLK(clk), .RST(rst), .Q(c[515]) );
  DFF \sreg_reg[518]  ( .D(c[518]), .CLK(clk), .RST(rst), .Q(c[514]) );
  DFF \sreg_reg[517]  ( .D(c[517]), .CLK(clk), .RST(rst), .Q(c[513]) );
  DFF \sreg_reg[516]  ( .D(c[516]), .CLK(clk), .RST(rst), .Q(c[512]) );
  DFF \sreg_reg[515]  ( .D(c[515]), .CLK(clk), .RST(rst), .Q(c[511]) );
  DFF \sreg_reg[514]  ( .D(c[514]), .CLK(clk), .RST(rst), .Q(c[510]) );
  DFF \sreg_reg[513]  ( .D(c[513]), .CLK(clk), .RST(rst), .Q(c[509]) );
  DFF \sreg_reg[512]  ( .D(c[512]), .CLK(clk), .RST(rst), .Q(c[508]) );
  DFF \sreg_reg[511]  ( .D(c[511]), .CLK(clk), .RST(rst), .Q(c[507]) );
  DFF \sreg_reg[510]  ( .D(c[510]), .CLK(clk), .RST(rst), .Q(c[506]) );
  DFF \sreg_reg[509]  ( .D(c[509]), .CLK(clk), .RST(rst), .Q(c[505]) );
  DFF \sreg_reg[508]  ( .D(c[508]), .CLK(clk), .RST(rst), .Q(c[504]) );
  DFF \sreg_reg[507]  ( .D(c[507]), .CLK(clk), .RST(rst), .Q(c[503]) );
  DFF \sreg_reg[506]  ( .D(c[506]), .CLK(clk), .RST(rst), .Q(c[502]) );
  DFF \sreg_reg[505]  ( .D(c[505]), .CLK(clk), .RST(rst), .Q(c[501]) );
  DFF \sreg_reg[504]  ( .D(c[504]), .CLK(clk), .RST(rst), .Q(c[500]) );
  DFF \sreg_reg[503]  ( .D(c[503]), .CLK(clk), .RST(rst), .Q(c[499]) );
  DFF \sreg_reg[502]  ( .D(c[502]), .CLK(clk), .RST(rst), .Q(c[498]) );
  DFF \sreg_reg[501]  ( .D(c[501]), .CLK(clk), .RST(rst), .Q(c[497]) );
  DFF \sreg_reg[500]  ( .D(c[500]), .CLK(clk), .RST(rst), .Q(c[496]) );
  DFF \sreg_reg[499]  ( .D(c[499]), .CLK(clk), .RST(rst), .Q(c[495]) );
  DFF \sreg_reg[498]  ( .D(c[498]), .CLK(clk), .RST(rst), .Q(c[494]) );
  DFF \sreg_reg[497]  ( .D(c[497]), .CLK(clk), .RST(rst), .Q(c[493]) );
  DFF \sreg_reg[496]  ( .D(c[496]), .CLK(clk), .RST(rst), .Q(c[492]) );
  DFF \sreg_reg[495]  ( .D(c[495]), .CLK(clk), .RST(rst), .Q(c[491]) );
  DFF \sreg_reg[494]  ( .D(c[494]), .CLK(clk), .RST(rst), .Q(c[490]) );
  DFF \sreg_reg[493]  ( .D(c[493]), .CLK(clk), .RST(rst), .Q(c[489]) );
  DFF \sreg_reg[492]  ( .D(c[492]), .CLK(clk), .RST(rst), .Q(c[488]) );
  DFF \sreg_reg[491]  ( .D(c[491]), .CLK(clk), .RST(rst), .Q(c[487]) );
  DFF \sreg_reg[490]  ( .D(c[490]), .CLK(clk), .RST(rst), .Q(c[486]) );
  DFF \sreg_reg[489]  ( .D(c[489]), .CLK(clk), .RST(rst), .Q(c[485]) );
  DFF \sreg_reg[488]  ( .D(c[488]), .CLK(clk), .RST(rst), .Q(c[484]) );
  DFF \sreg_reg[487]  ( .D(c[487]), .CLK(clk), .RST(rst), .Q(c[483]) );
  DFF \sreg_reg[486]  ( .D(c[486]), .CLK(clk), .RST(rst), .Q(c[482]) );
  DFF \sreg_reg[485]  ( .D(c[485]), .CLK(clk), .RST(rst), .Q(c[481]) );
  DFF \sreg_reg[484]  ( .D(c[484]), .CLK(clk), .RST(rst), .Q(c[480]) );
  DFF \sreg_reg[483]  ( .D(c[483]), .CLK(clk), .RST(rst), .Q(c[479]) );
  DFF \sreg_reg[482]  ( .D(c[482]), .CLK(clk), .RST(rst), .Q(c[478]) );
  DFF \sreg_reg[481]  ( .D(c[481]), .CLK(clk), .RST(rst), .Q(c[477]) );
  DFF \sreg_reg[480]  ( .D(c[480]), .CLK(clk), .RST(rst), .Q(c[476]) );
  DFF \sreg_reg[479]  ( .D(c[479]), .CLK(clk), .RST(rst), .Q(c[475]) );
  DFF \sreg_reg[478]  ( .D(c[478]), .CLK(clk), .RST(rst), .Q(c[474]) );
  DFF \sreg_reg[477]  ( .D(c[477]), .CLK(clk), .RST(rst), .Q(c[473]) );
  DFF \sreg_reg[476]  ( .D(c[476]), .CLK(clk), .RST(rst), .Q(c[472]) );
  DFF \sreg_reg[475]  ( .D(c[475]), .CLK(clk), .RST(rst), .Q(c[471]) );
  DFF \sreg_reg[474]  ( .D(c[474]), .CLK(clk), .RST(rst), .Q(c[470]) );
  DFF \sreg_reg[473]  ( .D(c[473]), .CLK(clk), .RST(rst), .Q(c[469]) );
  DFF \sreg_reg[472]  ( .D(c[472]), .CLK(clk), .RST(rst), .Q(c[468]) );
  DFF \sreg_reg[471]  ( .D(c[471]), .CLK(clk), .RST(rst), .Q(c[467]) );
  DFF \sreg_reg[470]  ( .D(c[470]), .CLK(clk), .RST(rst), .Q(c[466]) );
  DFF \sreg_reg[469]  ( .D(c[469]), .CLK(clk), .RST(rst), .Q(c[465]) );
  DFF \sreg_reg[468]  ( .D(c[468]), .CLK(clk), .RST(rst), .Q(c[464]) );
  DFF \sreg_reg[467]  ( .D(c[467]), .CLK(clk), .RST(rst), .Q(c[463]) );
  DFF \sreg_reg[466]  ( .D(c[466]), .CLK(clk), .RST(rst), .Q(c[462]) );
  DFF \sreg_reg[465]  ( .D(c[465]), .CLK(clk), .RST(rst), .Q(c[461]) );
  DFF \sreg_reg[464]  ( .D(c[464]), .CLK(clk), .RST(rst), .Q(c[460]) );
  DFF \sreg_reg[463]  ( .D(c[463]), .CLK(clk), .RST(rst), .Q(c[459]) );
  DFF \sreg_reg[462]  ( .D(c[462]), .CLK(clk), .RST(rst), .Q(c[458]) );
  DFF \sreg_reg[461]  ( .D(c[461]), .CLK(clk), .RST(rst), .Q(c[457]) );
  DFF \sreg_reg[460]  ( .D(c[460]), .CLK(clk), .RST(rst), .Q(c[456]) );
  DFF \sreg_reg[459]  ( .D(c[459]), .CLK(clk), .RST(rst), .Q(c[455]) );
  DFF \sreg_reg[458]  ( .D(c[458]), .CLK(clk), .RST(rst), .Q(c[454]) );
  DFF \sreg_reg[457]  ( .D(c[457]), .CLK(clk), .RST(rst), .Q(c[453]) );
  DFF \sreg_reg[456]  ( .D(c[456]), .CLK(clk), .RST(rst), .Q(c[452]) );
  DFF \sreg_reg[455]  ( .D(c[455]), .CLK(clk), .RST(rst), .Q(c[451]) );
  DFF \sreg_reg[454]  ( .D(c[454]), .CLK(clk), .RST(rst), .Q(c[450]) );
  DFF \sreg_reg[453]  ( .D(c[453]), .CLK(clk), .RST(rst), .Q(c[449]) );
  DFF \sreg_reg[452]  ( .D(c[452]), .CLK(clk), .RST(rst), .Q(c[448]) );
  DFF \sreg_reg[451]  ( .D(c[451]), .CLK(clk), .RST(rst), .Q(c[447]) );
  DFF \sreg_reg[450]  ( .D(c[450]), .CLK(clk), .RST(rst), .Q(c[446]) );
  DFF \sreg_reg[449]  ( .D(c[449]), .CLK(clk), .RST(rst), .Q(c[445]) );
  DFF \sreg_reg[448]  ( .D(c[448]), .CLK(clk), .RST(rst), .Q(c[444]) );
  DFF \sreg_reg[447]  ( .D(c[447]), .CLK(clk), .RST(rst), .Q(c[443]) );
  DFF \sreg_reg[446]  ( .D(c[446]), .CLK(clk), .RST(rst), .Q(c[442]) );
  DFF \sreg_reg[445]  ( .D(c[445]), .CLK(clk), .RST(rst), .Q(c[441]) );
  DFF \sreg_reg[444]  ( .D(c[444]), .CLK(clk), .RST(rst), .Q(c[440]) );
  DFF \sreg_reg[443]  ( .D(c[443]), .CLK(clk), .RST(rst), .Q(c[439]) );
  DFF \sreg_reg[442]  ( .D(c[442]), .CLK(clk), .RST(rst), .Q(c[438]) );
  DFF \sreg_reg[441]  ( .D(c[441]), .CLK(clk), .RST(rst), .Q(c[437]) );
  DFF \sreg_reg[440]  ( .D(c[440]), .CLK(clk), .RST(rst), .Q(c[436]) );
  DFF \sreg_reg[439]  ( .D(c[439]), .CLK(clk), .RST(rst), .Q(c[435]) );
  DFF \sreg_reg[438]  ( .D(c[438]), .CLK(clk), .RST(rst), .Q(c[434]) );
  DFF \sreg_reg[437]  ( .D(c[437]), .CLK(clk), .RST(rst), .Q(c[433]) );
  DFF \sreg_reg[436]  ( .D(c[436]), .CLK(clk), .RST(rst), .Q(c[432]) );
  DFF \sreg_reg[435]  ( .D(c[435]), .CLK(clk), .RST(rst), .Q(c[431]) );
  DFF \sreg_reg[434]  ( .D(c[434]), .CLK(clk), .RST(rst), .Q(c[430]) );
  DFF \sreg_reg[433]  ( .D(c[433]), .CLK(clk), .RST(rst), .Q(c[429]) );
  DFF \sreg_reg[432]  ( .D(c[432]), .CLK(clk), .RST(rst), .Q(c[428]) );
  DFF \sreg_reg[431]  ( .D(c[431]), .CLK(clk), .RST(rst), .Q(c[427]) );
  DFF \sreg_reg[430]  ( .D(c[430]), .CLK(clk), .RST(rst), .Q(c[426]) );
  DFF \sreg_reg[429]  ( .D(c[429]), .CLK(clk), .RST(rst), .Q(c[425]) );
  DFF \sreg_reg[428]  ( .D(c[428]), .CLK(clk), .RST(rst), .Q(c[424]) );
  DFF \sreg_reg[427]  ( .D(c[427]), .CLK(clk), .RST(rst), .Q(c[423]) );
  DFF \sreg_reg[426]  ( .D(c[426]), .CLK(clk), .RST(rst), .Q(c[422]) );
  DFF \sreg_reg[425]  ( .D(c[425]), .CLK(clk), .RST(rst), .Q(c[421]) );
  DFF \sreg_reg[424]  ( .D(c[424]), .CLK(clk), .RST(rst), .Q(c[420]) );
  DFF \sreg_reg[423]  ( .D(c[423]), .CLK(clk), .RST(rst), .Q(c[419]) );
  DFF \sreg_reg[422]  ( .D(c[422]), .CLK(clk), .RST(rst), .Q(c[418]) );
  DFF \sreg_reg[421]  ( .D(c[421]), .CLK(clk), .RST(rst), .Q(c[417]) );
  DFF \sreg_reg[420]  ( .D(c[420]), .CLK(clk), .RST(rst), .Q(c[416]) );
  DFF \sreg_reg[419]  ( .D(c[419]), .CLK(clk), .RST(rst), .Q(c[415]) );
  DFF \sreg_reg[418]  ( .D(c[418]), .CLK(clk), .RST(rst), .Q(c[414]) );
  DFF \sreg_reg[417]  ( .D(c[417]), .CLK(clk), .RST(rst), .Q(c[413]) );
  DFF \sreg_reg[416]  ( .D(c[416]), .CLK(clk), .RST(rst), .Q(c[412]) );
  DFF \sreg_reg[415]  ( .D(c[415]), .CLK(clk), .RST(rst), .Q(c[411]) );
  DFF \sreg_reg[414]  ( .D(c[414]), .CLK(clk), .RST(rst), .Q(c[410]) );
  DFF \sreg_reg[413]  ( .D(c[413]), .CLK(clk), .RST(rst), .Q(c[409]) );
  DFF \sreg_reg[412]  ( .D(c[412]), .CLK(clk), .RST(rst), .Q(c[408]) );
  DFF \sreg_reg[411]  ( .D(c[411]), .CLK(clk), .RST(rst), .Q(c[407]) );
  DFF \sreg_reg[410]  ( .D(c[410]), .CLK(clk), .RST(rst), .Q(c[406]) );
  DFF \sreg_reg[409]  ( .D(c[409]), .CLK(clk), .RST(rst), .Q(c[405]) );
  DFF \sreg_reg[408]  ( .D(c[408]), .CLK(clk), .RST(rst), .Q(c[404]) );
  DFF \sreg_reg[407]  ( .D(c[407]), .CLK(clk), .RST(rst), .Q(c[403]) );
  DFF \sreg_reg[406]  ( .D(c[406]), .CLK(clk), .RST(rst), .Q(c[402]) );
  DFF \sreg_reg[405]  ( .D(c[405]), .CLK(clk), .RST(rst), .Q(c[401]) );
  DFF \sreg_reg[404]  ( .D(c[404]), .CLK(clk), .RST(rst), .Q(c[400]) );
  DFF \sreg_reg[403]  ( .D(c[403]), .CLK(clk), .RST(rst), .Q(c[399]) );
  DFF \sreg_reg[402]  ( .D(c[402]), .CLK(clk), .RST(rst), .Q(c[398]) );
  DFF \sreg_reg[401]  ( .D(c[401]), .CLK(clk), .RST(rst), .Q(c[397]) );
  DFF \sreg_reg[400]  ( .D(c[400]), .CLK(clk), .RST(rst), .Q(c[396]) );
  DFF \sreg_reg[399]  ( .D(c[399]), .CLK(clk), .RST(rst), .Q(c[395]) );
  DFF \sreg_reg[398]  ( .D(c[398]), .CLK(clk), .RST(rst), .Q(c[394]) );
  DFF \sreg_reg[397]  ( .D(c[397]), .CLK(clk), .RST(rst), .Q(c[393]) );
  DFF \sreg_reg[396]  ( .D(c[396]), .CLK(clk), .RST(rst), .Q(c[392]) );
  DFF \sreg_reg[395]  ( .D(c[395]), .CLK(clk), .RST(rst), .Q(c[391]) );
  DFF \sreg_reg[394]  ( .D(c[394]), .CLK(clk), .RST(rst), .Q(c[390]) );
  DFF \sreg_reg[393]  ( .D(c[393]), .CLK(clk), .RST(rst), .Q(c[389]) );
  DFF \sreg_reg[392]  ( .D(c[392]), .CLK(clk), .RST(rst), .Q(c[388]) );
  DFF \sreg_reg[391]  ( .D(c[391]), .CLK(clk), .RST(rst), .Q(c[387]) );
  DFF \sreg_reg[390]  ( .D(c[390]), .CLK(clk), .RST(rst), .Q(c[386]) );
  DFF \sreg_reg[389]  ( .D(c[389]), .CLK(clk), .RST(rst), .Q(c[385]) );
  DFF \sreg_reg[388]  ( .D(c[388]), .CLK(clk), .RST(rst), .Q(c[384]) );
  DFF \sreg_reg[387]  ( .D(c[387]), .CLK(clk), .RST(rst), .Q(c[383]) );
  DFF \sreg_reg[386]  ( .D(c[386]), .CLK(clk), .RST(rst), .Q(c[382]) );
  DFF \sreg_reg[385]  ( .D(c[385]), .CLK(clk), .RST(rst), .Q(c[381]) );
  DFF \sreg_reg[384]  ( .D(c[384]), .CLK(clk), .RST(rst), .Q(c[380]) );
  DFF \sreg_reg[383]  ( .D(c[383]), .CLK(clk), .RST(rst), .Q(c[379]) );
  DFF \sreg_reg[382]  ( .D(c[382]), .CLK(clk), .RST(rst), .Q(c[378]) );
  DFF \sreg_reg[381]  ( .D(c[381]), .CLK(clk), .RST(rst), .Q(c[377]) );
  DFF \sreg_reg[380]  ( .D(c[380]), .CLK(clk), .RST(rst), .Q(c[376]) );
  DFF \sreg_reg[379]  ( .D(c[379]), .CLK(clk), .RST(rst), .Q(c[375]) );
  DFF \sreg_reg[378]  ( .D(c[378]), .CLK(clk), .RST(rst), .Q(c[374]) );
  DFF \sreg_reg[377]  ( .D(c[377]), .CLK(clk), .RST(rst), .Q(c[373]) );
  DFF \sreg_reg[376]  ( .D(c[376]), .CLK(clk), .RST(rst), .Q(c[372]) );
  DFF \sreg_reg[375]  ( .D(c[375]), .CLK(clk), .RST(rst), .Q(c[371]) );
  DFF \sreg_reg[374]  ( .D(c[374]), .CLK(clk), .RST(rst), .Q(c[370]) );
  DFF \sreg_reg[373]  ( .D(c[373]), .CLK(clk), .RST(rst), .Q(c[369]) );
  DFF \sreg_reg[372]  ( .D(c[372]), .CLK(clk), .RST(rst), .Q(c[368]) );
  DFF \sreg_reg[371]  ( .D(c[371]), .CLK(clk), .RST(rst), .Q(c[367]) );
  DFF \sreg_reg[370]  ( .D(c[370]), .CLK(clk), .RST(rst), .Q(c[366]) );
  DFF \sreg_reg[369]  ( .D(c[369]), .CLK(clk), .RST(rst), .Q(c[365]) );
  DFF \sreg_reg[368]  ( .D(c[368]), .CLK(clk), .RST(rst), .Q(c[364]) );
  DFF \sreg_reg[367]  ( .D(c[367]), .CLK(clk), .RST(rst), .Q(c[363]) );
  DFF \sreg_reg[366]  ( .D(c[366]), .CLK(clk), .RST(rst), .Q(c[362]) );
  DFF \sreg_reg[365]  ( .D(c[365]), .CLK(clk), .RST(rst), .Q(c[361]) );
  DFF \sreg_reg[364]  ( .D(c[364]), .CLK(clk), .RST(rst), .Q(c[360]) );
  DFF \sreg_reg[363]  ( .D(c[363]), .CLK(clk), .RST(rst), .Q(c[359]) );
  DFF \sreg_reg[362]  ( .D(c[362]), .CLK(clk), .RST(rst), .Q(c[358]) );
  DFF \sreg_reg[361]  ( .D(c[361]), .CLK(clk), .RST(rst), .Q(c[357]) );
  DFF \sreg_reg[360]  ( .D(c[360]), .CLK(clk), .RST(rst), .Q(c[356]) );
  DFF \sreg_reg[359]  ( .D(c[359]), .CLK(clk), .RST(rst), .Q(c[355]) );
  DFF \sreg_reg[358]  ( .D(c[358]), .CLK(clk), .RST(rst), .Q(c[354]) );
  DFF \sreg_reg[357]  ( .D(c[357]), .CLK(clk), .RST(rst), .Q(c[353]) );
  DFF \sreg_reg[356]  ( .D(c[356]), .CLK(clk), .RST(rst), .Q(c[352]) );
  DFF \sreg_reg[355]  ( .D(c[355]), .CLK(clk), .RST(rst), .Q(c[351]) );
  DFF \sreg_reg[354]  ( .D(c[354]), .CLK(clk), .RST(rst), .Q(c[350]) );
  DFF \sreg_reg[353]  ( .D(c[353]), .CLK(clk), .RST(rst), .Q(c[349]) );
  DFF \sreg_reg[352]  ( .D(c[352]), .CLK(clk), .RST(rst), .Q(c[348]) );
  DFF \sreg_reg[351]  ( .D(c[351]), .CLK(clk), .RST(rst), .Q(c[347]) );
  DFF \sreg_reg[350]  ( .D(c[350]), .CLK(clk), .RST(rst), .Q(c[346]) );
  DFF \sreg_reg[349]  ( .D(c[349]), .CLK(clk), .RST(rst), .Q(c[345]) );
  DFF \sreg_reg[348]  ( .D(c[348]), .CLK(clk), .RST(rst), .Q(c[344]) );
  DFF \sreg_reg[347]  ( .D(c[347]), .CLK(clk), .RST(rst), .Q(c[343]) );
  DFF \sreg_reg[346]  ( .D(c[346]), .CLK(clk), .RST(rst), .Q(c[342]) );
  DFF \sreg_reg[345]  ( .D(c[345]), .CLK(clk), .RST(rst), .Q(c[341]) );
  DFF \sreg_reg[344]  ( .D(c[344]), .CLK(clk), .RST(rst), .Q(c[340]) );
  DFF \sreg_reg[343]  ( .D(c[343]), .CLK(clk), .RST(rst), .Q(c[339]) );
  DFF \sreg_reg[342]  ( .D(c[342]), .CLK(clk), .RST(rst), .Q(c[338]) );
  DFF \sreg_reg[341]  ( .D(c[341]), .CLK(clk), .RST(rst), .Q(c[337]) );
  DFF \sreg_reg[340]  ( .D(c[340]), .CLK(clk), .RST(rst), .Q(c[336]) );
  DFF \sreg_reg[339]  ( .D(c[339]), .CLK(clk), .RST(rst), .Q(c[335]) );
  DFF \sreg_reg[338]  ( .D(c[338]), .CLK(clk), .RST(rst), .Q(c[334]) );
  DFF \sreg_reg[337]  ( .D(c[337]), .CLK(clk), .RST(rst), .Q(c[333]) );
  DFF \sreg_reg[336]  ( .D(c[336]), .CLK(clk), .RST(rst), .Q(c[332]) );
  DFF \sreg_reg[335]  ( .D(c[335]), .CLK(clk), .RST(rst), .Q(c[331]) );
  DFF \sreg_reg[334]  ( .D(c[334]), .CLK(clk), .RST(rst), .Q(c[330]) );
  DFF \sreg_reg[333]  ( .D(c[333]), .CLK(clk), .RST(rst), .Q(c[329]) );
  DFF \sreg_reg[332]  ( .D(c[332]), .CLK(clk), .RST(rst), .Q(c[328]) );
  DFF \sreg_reg[331]  ( .D(c[331]), .CLK(clk), .RST(rst), .Q(c[327]) );
  DFF \sreg_reg[330]  ( .D(c[330]), .CLK(clk), .RST(rst), .Q(c[326]) );
  DFF \sreg_reg[329]  ( .D(c[329]), .CLK(clk), .RST(rst), .Q(c[325]) );
  DFF \sreg_reg[328]  ( .D(c[328]), .CLK(clk), .RST(rst), .Q(c[324]) );
  DFF \sreg_reg[327]  ( .D(c[327]), .CLK(clk), .RST(rst), .Q(c[323]) );
  DFF \sreg_reg[326]  ( .D(c[326]), .CLK(clk), .RST(rst), .Q(c[322]) );
  DFF \sreg_reg[325]  ( .D(c[325]), .CLK(clk), .RST(rst), .Q(c[321]) );
  DFF \sreg_reg[324]  ( .D(c[324]), .CLK(clk), .RST(rst), .Q(c[320]) );
  DFF \sreg_reg[323]  ( .D(c[323]), .CLK(clk), .RST(rst), .Q(c[319]) );
  DFF \sreg_reg[322]  ( .D(c[322]), .CLK(clk), .RST(rst), .Q(c[318]) );
  DFF \sreg_reg[321]  ( .D(c[321]), .CLK(clk), .RST(rst), .Q(c[317]) );
  DFF \sreg_reg[320]  ( .D(c[320]), .CLK(clk), .RST(rst), .Q(c[316]) );
  DFF \sreg_reg[319]  ( .D(c[319]), .CLK(clk), .RST(rst), .Q(c[315]) );
  DFF \sreg_reg[318]  ( .D(c[318]), .CLK(clk), .RST(rst), .Q(c[314]) );
  DFF \sreg_reg[317]  ( .D(c[317]), .CLK(clk), .RST(rst), .Q(c[313]) );
  DFF \sreg_reg[316]  ( .D(c[316]), .CLK(clk), .RST(rst), .Q(c[312]) );
  DFF \sreg_reg[315]  ( .D(c[315]), .CLK(clk), .RST(rst), .Q(c[311]) );
  DFF \sreg_reg[314]  ( .D(c[314]), .CLK(clk), .RST(rst), .Q(c[310]) );
  DFF \sreg_reg[313]  ( .D(c[313]), .CLK(clk), .RST(rst), .Q(c[309]) );
  DFF \sreg_reg[312]  ( .D(c[312]), .CLK(clk), .RST(rst), .Q(c[308]) );
  DFF \sreg_reg[311]  ( .D(c[311]), .CLK(clk), .RST(rst), .Q(c[307]) );
  DFF \sreg_reg[310]  ( .D(c[310]), .CLK(clk), .RST(rst), .Q(c[306]) );
  DFF \sreg_reg[309]  ( .D(c[309]), .CLK(clk), .RST(rst), .Q(c[305]) );
  DFF \sreg_reg[308]  ( .D(c[308]), .CLK(clk), .RST(rst), .Q(c[304]) );
  DFF \sreg_reg[307]  ( .D(c[307]), .CLK(clk), .RST(rst), .Q(c[303]) );
  DFF \sreg_reg[306]  ( .D(c[306]), .CLK(clk), .RST(rst), .Q(c[302]) );
  DFF \sreg_reg[305]  ( .D(c[305]), .CLK(clk), .RST(rst), .Q(c[301]) );
  DFF \sreg_reg[304]  ( .D(c[304]), .CLK(clk), .RST(rst), .Q(c[300]) );
  DFF \sreg_reg[303]  ( .D(c[303]), .CLK(clk), .RST(rst), .Q(c[299]) );
  DFF \sreg_reg[302]  ( .D(c[302]), .CLK(clk), .RST(rst), .Q(c[298]) );
  DFF \sreg_reg[301]  ( .D(c[301]), .CLK(clk), .RST(rst), .Q(c[297]) );
  DFF \sreg_reg[300]  ( .D(c[300]), .CLK(clk), .RST(rst), .Q(c[296]) );
  DFF \sreg_reg[299]  ( .D(c[299]), .CLK(clk), .RST(rst), .Q(c[295]) );
  DFF \sreg_reg[298]  ( .D(c[298]), .CLK(clk), .RST(rst), .Q(c[294]) );
  DFF \sreg_reg[297]  ( .D(c[297]), .CLK(clk), .RST(rst), .Q(c[293]) );
  DFF \sreg_reg[296]  ( .D(c[296]), .CLK(clk), .RST(rst), .Q(c[292]) );
  DFF \sreg_reg[295]  ( .D(c[295]), .CLK(clk), .RST(rst), .Q(c[291]) );
  DFF \sreg_reg[294]  ( .D(c[294]), .CLK(clk), .RST(rst), .Q(c[290]) );
  DFF \sreg_reg[293]  ( .D(c[293]), .CLK(clk), .RST(rst), .Q(c[289]) );
  DFF \sreg_reg[292]  ( .D(c[292]), .CLK(clk), .RST(rst), .Q(c[288]) );
  DFF \sreg_reg[291]  ( .D(c[291]), .CLK(clk), .RST(rst), .Q(c[287]) );
  DFF \sreg_reg[290]  ( .D(c[290]), .CLK(clk), .RST(rst), .Q(c[286]) );
  DFF \sreg_reg[289]  ( .D(c[289]), .CLK(clk), .RST(rst), .Q(c[285]) );
  DFF \sreg_reg[288]  ( .D(c[288]), .CLK(clk), .RST(rst), .Q(c[284]) );
  DFF \sreg_reg[287]  ( .D(c[287]), .CLK(clk), .RST(rst), .Q(c[283]) );
  DFF \sreg_reg[286]  ( .D(c[286]), .CLK(clk), .RST(rst), .Q(c[282]) );
  DFF \sreg_reg[285]  ( .D(c[285]), .CLK(clk), .RST(rst), .Q(c[281]) );
  DFF \sreg_reg[284]  ( .D(c[284]), .CLK(clk), .RST(rst), .Q(c[280]) );
  DFF \sreg_reg[283]  ( .D(c[283]), .CLK(clk), .RST(rst), .Q(c[279]) );
  DFF \sreg_reg[282]  ( .D(c[282]), .CLK(clk), .RST(rst), .Q(c[278]) );
  DFF \sreg_reg[281]  ( .D(c[281]), .CLK(clk), .RST(rst), .Q(c[277]) );
  DFF \sreg_reg[280]  ( .D(c[280]), .CLK(clk), .RST(rst), .Q(c[276]) );
  DFF \sreg_reg[279]  ( .D(c[279]), .CLK(clk), .RST(rst), .Q(c[275]) );
  DFF \sreg_reg[278]  ( .D(c[278]), .CLK(clk), .RST(rst), .Q(c[274]) );
  DFF \sreg_reg[277]  ( .D(c[277]), .CLK(clk), .RST(rst), .Q(c[273]) );
  DFF \sreg_reg[276]  ( .D(c[276]), .CLK(clk), .RST(rst), .Q(c[272]) );
  DFF \sreg_reg[275]  ( .D(c[275]), .CLK(clk), .RST(rst), .Q(c[271]) );
  DFF \sreg_reg[274]  ( .D(c[274]), .CLK(clk), .RST(rst), .Q(c[270]) );
  DFF \sreg_reg[273]  ( .D(c[273]), .CLK(clk), .RST(rst), .Q(c[269]) );
  DFF \sreg_reg[272]  ( .D(c[272]), .CLK(clk), .RST(rst), .Q(c[268]) );
  DFF \sreg_reg[271]  ( .D(c[271]), .CLK(clk), .RST(rst), .Q(c[267]) );
  DFF \sreg_reg[270]  ( .D(c[270]), .CLK(clk), .RST(rst), .Q(c[266]) );
  DFF \sreg_reg[269]  ( .D(c[269]), .CLK(clk), .RST(rst), .Q(c[265]) );
  DFF \sreg_reg[268]  ( .D(c[268]), .CLK(clk), .RST(rst), .Q(c[264]) );
  DFF \sreg_reg[267]  ( .D(c[267]), .CLK(clk), .RST(rst), .Q(c[263]) );
  DFF \sreg_reg[266]  ( .D(c[266]), .CLK(clk), .RST(rst), .Q(c[262]) );
  DFF \sreg_reg[265]  ( .D(c[265]), .CLK(clk), .RST(rst), .Q(c[261]) );
  DFF \sreg_reg[264]  ( .D(c[264]), .CLK(clk), .RST(rst), .Q(c[260]) );
  DFF \sreg_reg[263]  ( .D(c[263]), .CLK(clk), .RST(rst), .Q(c[259]) );
  DFF \sreg_reg[262]  ( .D(c[262]), .CLK(clk), .RST(rst), .Q(c[258]) );
  DFF \sreg_reg[261]  ( .D(c[261]), .CLK(clk), .RST(rst), .Q(c[257]) );
  DFF \sreg_reg[260]  ( .D(c[260]), .CLK(clk), .RST(rst), .Q(c[256]) );
  DFF \sreg_reg[259]  ( .D(c[259]), .CLK(clk), .RST(rst), .Q(c[255]) );
  DFF \sreg_reg[258]  ( .D(c[258]), .CLK(clk), .RST(rst), .Q(c[254]) );
  DFF \sreg_reg[257]  ( .D(c[257]), .CLK(clk), .RST(rst), .Q(c[253]) );
  DFF \sreg_reg[256]  ( .D(c[256]), .CLK(clk), .RST(rst), .Q(c[252]) );
  DFF \sreg_reg[255]  ( .D(c[255]), .CLK(clk), .RST(rst), .Q(c[251]) );
  DFF \sreg_reg[254]  ( .D(c[254]), .CLK(clk), .RST(rst), .Q(c[250]) );
  DFF \sreg_reg[253]  ( .D(c[253]), .CLK(clk), .RST(rst), .Q(c[249]) );
  DFF \sreg_reg[252]  ( .D(c[252]), .CLK(clk), .RST(rst), .Q(c[248]) );
  DFF \sreg_reg[251]  ( .D(c[251]), .CLK(clk), .RST(rst), .Q(c[247]) );
  DFF \sreg_reg[250]  ( .D(c[250]), .CLK(clk), .RST(rst), .Q(c[246]) );
  DFF \sreg_reg[249]  ( .D(c[249]), .CLK(clk), .RST(rst), .Q(c[245]) );
  DFF \sreg_reg[248]  ( .D(c[248]), .CLK(clk), .RST(rst), .Q(c[244]) );
  DFF \sreg_reg[247]  ( .D(c[247]), .CLK(clk), .RST(rst), .Q(c[243]) );
  DFF \sreg_reg[246]  ( .D(c[246]), .CLK(clk), .RST(rst), .Q(c[242]) );
  DFF \sreg_reg[245]  ( .D(c[245]), .CLK(clk), .RST(rst), .Q(c[241]) );
  DFF \sreg_reg[244]  ( .D(c[244]), .CLK(clk), .RST(rst), .Q(c[240]) );
  DFF \sreg_reg[243]  ( .D(c[243]), .CLK(clk), .RST(rst), .Q(c[239]) );
  DFF \sreg_reg[242]  ( .D(c[242]), .CLK(clk), .RST(rst), .Q(c[238]) );
  DFF \sreg_reg[241]  ( .D(c[241]), .CLK(clk), .RST(rst), .Q(c[237]) );
  DFF \sreg_reg[240]  ( .D(c[240]), .CLK(clk), .RST(rst), .Q(c[236]) );
  DFF \sreg_reg[239]  ( .D(c[239]), .CLK(clk), .RST(rst), .Q(c[235]) );
  DFF \sreg_reg[238]  ( .D(c[238]), .CLK(clk), .RST(rst), .Q(c[234]) );
  DFF \sreg_reg[237]  ( .D(c[237]), .CLK(clk), .RST(rst), .Q(c[233]) );
  DFF \sreg_reg[236]  ( .D(c[236]), .CLK(clk), .RST(rst), .Q(c[232]) );
  DFF \sreg_reg[235]  ( .D(c[235]), .CLK(clk), .RST(rst), .Q(c[231]) );
  DFF \sreg_reg[234]  ( .D(c[234]), .CLK(clk), .RST(rst), .Q(c[230]) );
  DFF \sreg_reg[233]  ( .D(c[233]), .CLK(clk), .RST(rst), .Q(c[229]) );
  DFF \sreg_reg[232]  ( .D(c[232]), .CLK(clk), .RST(rst), .Q(c[228]) );
  DFF \sreg_reg[231]  ( .D(c[231]), .CLK(clk), .RST(rst), .Q(c[227]) );
  DFF \sreg_reg[230]  ( .D(c[230]), .CLK(clk), .RST(rst), .Q(c[226]) );
  DFF \sreg_reg[229]  ( .D(c[229]), .CLK(clk), .RST(rst), .Q(c[225]) );
  DFF \sreg_reg[228]  ( .D(c[228]), .CLK(clk), .RST(rst), .Q(c[224]) );
  DFF \sreg_reg[227]  ( .D(c[227]), .CLK(clk), .RST(rst), .Q(c[223]) );
  DFF \sreg_reg[226]  ( .D(c[226]), .CLK(clk), .RST(rst), .Q(c[222]) );
  DFF \sreg_reg[225]  ( .D(c[225]), .CLK(clk), .RST(rst), .Q(c[221]) );
  DFF \sreg_reg[224]  ( .D(c[224]), .CLK(clk), .RST(rst), .Q(c[220]) );
  DFF \sreg_reg[223]  ( .D(c[223]), .CLK(clk), .RST(rst), .Q(c[219]) );
  DFF \sreg_reg[222]  ( .D(c[222]), .CLK(clk), .RST(rst), .Q(c[218]) );
  DFF \sreg_reg[221]  ( .D(c[221]), .CLK(clk), .RST(rst), .Q(c[217]) );
  DFF \sreg_reg[220]  ( .D(c[220]), .CLK(clk), .RST(rst), .Q(c[216]) );
  DFF \sreg_reg[219]  ( .D(c[219]), .CLK(clk), .RST(rst), .Q(c[215]) );
  DFF \sreg_reg[218]  ( .D(c[218]), .CLK(clk), .RST(rst), .Q(c[214]) );
  DFF \sreg_reg[217]  ( .D(c[217]), .CLK(clk), .RST(rst), .Q(c[213]) );
  DFF \sreg_reg[216]  ( .D(c[216]), .CLK(clk), .RST(rst), .Q(c[212]) );
  DFF \sreg_reg[215]  ( .D(c[215]), .CLK(clk), .RST(rst), .Q(c[211]) );
  DFF \sreg_reg[214]  ( .D(c[214]), .CLK(clk), .RST(rst), .Q(c[210]) );
  DFF \sreg_reg[213]  ( .D(c[213]), .CLK(clk), .RST(rst), .Q(c[209]) );
  DFF \sreg_reg[212]  ( .D(c[212]), .CLK(clk), .RST(rst), .Q(c[208]) );
  DFF \sreg_reg[211]  ( .D(c[211]), .CLK(clk), .RST(rst), .Q(c[207]) );
  DFF \sreg_reg[210]  ( .D(c[210]), .CLK(clk), .RST(rst), .Q(c[206]) );
  DFF \sreg_reg[209]  ( .D(c[209]), .CLK(clk), .RST(rst), .Q(c[205]) );
  DFF \sreg_reg[208]  ( .D(c[208]), .CLK(clk), .RST(rst), .Q(c[204]) );
  DFF \sreg_reg[207]  ( .D(c[207]), .CLK(clk), .RST(rst), .Q(c[203]) );
  DFF \sreg_reg[206]  ( .D(c[206]), .CLK(clk), .RST(rst), .Q(c[202]) );
  DFF \sreg_reg[205]  ( .D(c[205]), .CLK(clk), .RST(rst), .Q(c[201]) );
  DFF \sreg_reg[204]  ( .D(c[204]), .CLK(clk), .RST(rst), .Q(c[200]) );
  DFF \sreg_reg[203]  ( .D(c[203]), .CLK(clk), .RST(rst), .Q(c[199]) );
  DFF \sreg_reg[202]  ( .D(c[202]), .CLK(clk), .RST(rst), .Q(c[198]) );
  DFF \sreg_reg[201]  ( .D(c[201]), .CLK(clk), .RST(rst), .Q(c[197]) );
  DFF \sreg_reg[200]  ( .D(c[200]), .CLK(clk), .RST(rst), .Q(c[196]) );
  DFF \sreg_reg[199]  ( .D(c[199]), .CLK(clk), .RST(rst), .Q(c[195]) );
  DFF \sreg_reg[198]  ( .D(c[198]), .CLK(clk), .RST(rst), .Q(c[194]) );
  DFF \sreg_reg[197]  ( .D(c[197]), .CLK(clk), .RST(rst), .Q(c[193]) );
  DFF \sreg_reg[196]  ( .D(c[196]), .CLK(clk), .RST(rst), .Q(c[192]) );
  DFF \sreg_reg[195]  ( .D(c[195]), .CLK(clk), .RST(rst), .Q(c[191]) );
  DFF \sreg_reg[194]  ( .D(c[194]), .CLK(clk), .RST(rst), .Q(c[190]) );
  DFF \sreg_reg[193]  ( .D(c[193]), .CLK(clk), .RST(rst), .Q(c[189]) );
  DFF \sreg_reg[192]  ( .D(c[192]), .CLK(clk), .RST(rst), .Q(c[188]) );
  DFF \sreg_reg[191]  ( .D(c[191]), .CLK(clk), .RST(rst), .Q(c[187]) );
  DFF \sreg_reg[190]  ( .D(c[190]), .CLK(clk), .RST(rst), .Q(c[186]) );
  DFF \sreg_reg[189]  ( .D(c[189]), .CLK(clk), .RST(rst), .Q(c[185]) );
  DFF \sreg_reg[188]  ( .D(c[188]), .CLK(clk), .RST(rst), .Q(c[184]) );
  DFF \sreg_reg[187]  ( .D(c[187]), .CLK(clk), .RST(rst), .Q(c[183]) );
  DFF \sreg_reg[186]  ( .D(c[186]), .CLK(clk), .RST(rst), .Q(c[182]) );
  DFF \sreg_reg[185]  ( .D(c[185]), .CLK(clk), .RST(rst), .Q(c[181]) );
  DFF \sreg_reg[184]  ( .D(c[184]), .CLK(clk), .RST(rst), .Q(c[180]) );
  DFF \sreg_reg[183]  ( .D(c[183]), .CLK(clk), .RST(rst), .Q(c[179]) );
  DFF \sreg_reg[182]  ( .D(c[182]), .CLK(clk), .RST(rst), .Q(c[178]) );
  DFF \sreg_reg[181]  ( .D(c[181]), .CLK(clk), .RST(rst), .Q(c[177]) );
  DFF \sreg_reg[180]  ( .D(c[180]), .CLK(clk), .RST(rst), .Q(c[176]) );
  DFF \sreg_reg[179]  ( .D(c[179]), .CLK(clk), .RST(rst), .Q(c[175]) );
  DFF \sreg_reg[178]  ( .D(c[178]), .CLK(clk), .RST(rst), .Q(c[174]) );
  DFF \sreg_reg[177]  ( .D(c[177]), .CLK(clk), .RST(rst), .Q(c[173]) );
  DFF \sreg_reg[176]  ( .D(c[176]), .CLK(clk), .RST(rst), .Q(c[172]) );
  DFF \sreg_reg[175]  ( .D(c[175]), .CLK(clk), .RST(rst), .Q(c[171]) );
  DFF \sreg_reg[174]  ( .D(c[174]), .CLK(clk), .RST(rst), .Q(c[170]) );
  DFF \sreg_reg[173]  ( .D(c[173]), .CLK(clk), .RST(rst), .Q(c[169]) );
  DFF \sreg_reg[172]  ( .D(c[172]), .CLK(clk), .RST(rst), .Q(c[168]) );
  DFF \sreg_reg[171]  ( .D(c[171]), .CLK(clk), .RST(rst), .Q(c[167]) );
  DFF \sreg_reg[170]  ( .D(c[170]), .CLK(clk), .RST(rst), .Q(c[166]) );
  DFF \sreg_reg[169]  ( .D(c[169]), .CLK(clk), .RST(rst), .Q(c[165]) );
  DFF \sreg_reg[168]  ( .D(c[168]), .CLK(clk), .RST(rst), .Q(c[164]) );
  DFF \sreg_reg[167]  ( .D(c[167]), .CLK(clk), .RST(rst), .Q(c[163]) );
  DFF \sreg_reg[166]  ( .D(c[166]), .CLK(clk), .RST(rst), .Q(c[162]) );
  DFF \sreg_reg[165]  ( .D(c[165]), .CLK(clk), .RST(rst), .Q(c[161]) );
  DFF \sreg_reg[164]  ( .D(c[164]), .CLK(clk), .RST(rst), .Q(c[160]) );
  DFF \sreg_reg[163]  ( .D(c[163]), .CLK(clk), .RST(rst), .Q(c[159]) );
  DFF \sreg_reg[162]  ( .D(c[162]), .CLK(clk), .RST(rst), .Q(c[158]) );
  DFF \sreg_reg[161]  ( .D(c[161]), .CLK(clk), .RST(rst), .Q(c[157]) );
  DFF \sreg_reg[160]  ( .D(c[160]), .CLK(clk), .RST(rst), .Q(c[156]) );
  DFF \sreg_reg[159]  ( .D(c[159]), .CLK(clk), .RST(rst), .Q(c[155]) );
  DFF \sreg_reg[158]  ( .D(c[158]), .CLK(clk), .RST(rst), .Q(c[154]) );
  DFF \sreg_reg[157]  ( .D(c[157]), .CLK(clk), .RST(rst), .Q(c[153]) );
  DFF \sreg_reg[156]  ( .D(c[156]), .CLK(clk), .RST(rst), .Q(c[152]) );
  DFF \sreg_reg[155]  ( .D(c[155]), .CLK(clk), .RST(rst), .Q(c[151]) );
  DFF \sreg_reg[154]  ( .D(c[154]), .CLK(clk), .RST(rst), .Q(c[150]) );
  DFF \sreg_reg[153]  ( .D(c[153]), .CLK(clk), .RST(rst), .Q(c[149]) );
  DFF \sreg_reg[152]  ( .D(c[152]), .CLK(clk), .RST(rst), .Q(c[148]) );
  DFF \sreg_reg[151]  ( .D(c[151]), .CLK(clk), .RST(rst), .Q(c[147]) );
  DFF \sreg_reg[150]  ( .D(c[150]), .CLK(clk), .RST(rst), .Q(c[146]) );
  DFF \sreg_reg[149]  ( .D(c[149]), .CLK(clk), .RST(rst), .Q(c[145]) );
  DFF \sreg_reg[148]  ( .D(c[148]), .CLK(clk), .RST(rst), .Q(c[144]) );
  DFF \sreg_reg[147]  ( .D(c[147]), .CLK(clk), .RST(rst), .Q(c[143]) );
  DFF \sreg_reg[146]  ( .D(c[146]), .CLK(clk), .RST(rst), .Q(c[142]) );
  DFF \sreg_reg[145]  ( .D(c[145]), .CLK(clk), .RST(rst), .Q(c[141]) );
  DFF \sreg_reg[144]  ( .D(c[144]), .CLK(clk), .RST(rst), .Q(c[140]) );
  DFF \sreg_reg[143]  ( .D(c[143]), .CLK(clk), .RST(rst), .Q(c[139]) );
  DFF \sreg_reg[142]  ( .D(c[142]), .CLK(clk), .RST(rst), .Q(c[138]) );
  DFF \sreg_reg[141]  ( .D(c[141]), .CLK(clk), .RST(rst), .Q(c[137]) );
  DFF \sreg_reg[140]  ( .D(c[140]), .CLK(clk), .RST(rst), .Q(c[136]) );
  DFF \sreg_reg[139]  ( .D(c[139]), .CLK(clk), .RST(rst), .Q(c[135]) );
  DFF \sreg_reg[138]  ( .D(c[138]), .CLK(clk), .RST(rst), .Q(c[134]) );
  DFF \sreg_reg[137]  ( .D(c[137]), .CLK(clk), .RST(rst), .Q(c[133]) );
  DFF \sreg_reg[136]  ( .D(c[136]), .CLK(clk), .RST(rst), .Q(c[132]) );
  DFF \sreg_reg[135]  ( .D(c[135]), .CLK(clk), .RST(rst), .Q(c[131]) );
  DFF \sreg_reg[134]  ( .D(c[134]), .CLK(clk), .RST(rst), .Q(c[130]) );
  DFF \sreg_reg[133]  ( .D(c[133]), .CLK(clk), .RST(rst), .Q(c[129]) );
  DFF \sreg_reg[132]  ( .D(c[132]), .CLK(clk), .RST(rst), .Q(c[128]) );
  DFF \sreg_reg[131]  ( .D(c[131]), .CLK(clk), .RST(rst), .Q(c[127]) );
  DFF \sreg_reg[130]  ( .D(c[130]), .CLK(clk), .RST(rst), .Q(c[126]) );
  DFF \sreg_reg[129]  ( .D(c[129]), .CLK(clk), .RST(rst), .Q(c[125]) );
  DFF \sreg_reg[128]  ( .D(c[128]), .CLK(clk), .RST(rst), .Q(c[124]) );
  DFF \sreg_reg[127]  ( .D(c[127]), .CLK(clk), .RST(rst), .Q(c[123]) );
  DFF \sreg_reg[126]  ( .D(c[126]), .CLK(clk), .RST(rst), .Q(c[122]) );
  DFF \sreg_reg[125]  ( .D(c[125]), .CLK(clk), .RST(rst), .Q(c[121]) );
  DFF \sreg_reg[124]  ( .D(c[124]), .CLK(clk), .RST(rst), .Q(c[120]) );
  DFF \sreg_reg[123]  ( .D(c[123]), .CLK(clk), .RST(rst), .Q(c[119]) );
  DFF \sreg_reg[122]  ( .D(c[122]), .CLK(clk), .RST(rst), .Q(c[118]) );
  DFF \sreg_reg[121]  ( .D(c[121]), .CLK(clk), .RST(rst), .Q(c[117]) );
  DFF \sreg_reg[120]  ( .D(c[120]), .CLK(clk), .RST(rst), .Q(c[116]) );
  DFF \sreg_reg[119]  ( .D(c[119]), .CLK(clk), .RST(rst), .Q(c[115]) );
  DFF \sreg_reg[118]  ( .D(c[118]), .CLK(clk), .RST(rst), .Q(c[114]) );
  DFF \sreg_reg[117]  ( .D(c[117]), .CLK(clk), .RST(rst), .Q(c[113]) );
  DFF \sreg_reg[116]  ( .D(c[116]), .CLK(clk), .RST(rst), .Q(c[112]) );
  DFF \sreg_reg[115]  ( .D(c[115]), .CLK(clk), .RST(rst), .Q(c[111]) );
  DFF \sreg_reg[114]  ( .D(c[114]), .CLK(clk), .RST(rst), .Q(c[110]) );
  DFF \sreg_reg[113]  ( .D(c[113]), .CLK(clk), .RST(rst), .Q(c[109]) );
  DFF \sreg_reg[112]  ( .D(c[112]), .CLK(clk), .RST(rst), .Q(c[108]) );
  DFF \sreg_reg[111]  ( .D(c[111]), .CLK(clk), .RST(rst), .Q(c[107]) );
  DFF \sreg_reg[110]  ( .D(c[110]), .CLK(clk), .RST(rst), .Q(c[106]) );
  DFF \sreg_reg[109]  ( .D(c[109]), .CLK(clk), .RST(rst), .Q(c[105]) );
  DFF \sreg_reg[108]  ( .D(c[108]), .CLK(clk), .RST(rst), .Q(c[104]) );
  DFF \sreg_reg[107]  ( .D(c[107]), .CLK(clk), .RST(rst), .Q(c[103]) );
  DFF \sreg_reg[106]  ( .D(c[106]), .CLK(clk), .RST(rst), .Q(c[102]) );
  DFF \sreg_reg[105]  ( .D(c[105]), .CLK(clk), .RST(rst), .Q(c[101]) );
  DFF \sreg_reg[104]  ( .D(c[104]), .CLK(clk), .RST(rst), .Q(c[100]) );
  DFF \sreg_reg[103]  ( .D(c[103]), .CLK(clk), .RST(rst), .Q(c[99]) );
  DFF \sreg_reg[102]  ( .D(c[102]), .CLK(clk), .RST(rst), .Q(c[98]) );
  DFF \sreg_reg[101]  ( .D(c[101]), .CLK(clk), .RST(rst), .Q(c[97]) );
  DFF \sreg_reg[100]  ( .D(c[100]), .CLK(clk), .RST(rst), .Q(c[96]) );
  DFF \sreg_reg[99]  ( .D(c[99]), .CLK(clk), .RST(rst), .Q(c[95]) );
  DFF \sreg_reg[98]  ( .D(c[98]), .CLK(clk), .RST(rst), .Q(c[94]) );
  DFF \sreg_reg[97]  ( .D(c[97]), .CLK(clk), .RST(rst), .Q(c[93]) );
  DFF \sreg_reg[96]  ( .D(c[96]), .CLK(clk), .RST(rst), .Q(c[92]) );
  DFF \sreg_reg[95]  ( .D(c[95]), .CLK(clk), .RST(rst), .Q(c[91]) );
  DFF \sreg_reg[94]  ( .D(c[94]), .CLK(clk), .RST(rst), .Q(c[90]) );
  DFF \sreg_reg[93]  ( .D(c[93]), .CLK(clk), .RST(rst), .Q(c[89]) );
  DFF \sreg_reg[92]  ( .D(c[92]), .CLK(clk), .RST(rst), .Q(c[88]) );
  DFF \sreg_reg[91]  ( .D(c[91]), .CLK(clk), .RST(rst), .Q(c[87]) );
  DFF \sreg_reg[90]  ( .D(c[90]), .CLK(clk), .RST(rst), .Q(c[86]) );
  DFF \sreg_reg[89]  ( .D(c[89]), .CLK(clk), .RST(rst), .Q(c[85]) );
  DFF \sreg_reg[88]  ( .D(c[88]), .CLK(clk), .RST(rst), .Q(c[84]) );
  DFF \sreg_reg[87]  ( .D(c[87]), .CLK(clk), .RST(rst), .Q(c[83]) );
  DFF \sreg_reg[86]  ( .D(c[86]), .CLK(clk), .RST(rst), .Q(c[82]) );
  DFF \sreg_reg[85]  ( .D(c[85]), .CLK(clk), .RST(rst), .Q(c[81]) );
  DFF \sreg_reg[84]  ( .D(c[84]), .CLK(clk), .RST(rst), .Q(c[80]) );
  DFF \sreg_reg[83]  ( .D(c[83]), .CLK(clk), .RST(rst), .Q(c[79]) );
  DFF \sreg_reg[82]  ( .D(c[82]), .CLK(clk), .RST(rst), .Q(c[78]) );
  DFF \sreg_reg[81]  ( .D(c[81]), .CLK(clk), .RST(rst), .Q(c[77]) );
  DFF \sreg_reg[80]  ( .D(c[80]), .CLK(clk), .RST(rst), .Q(c[76]) );
  DFF \sreg_reg[79]  ( .D(c[79]), .CLK(clk), .RST(rst), .Q(c[75]) );
  DFF \sreg_reg[78]  ( .D(c[78]), .CLK(clk), .RST(rst), .Q(c[74]) );
  DFF \sreg_reg[77]  ( .D(c[77]), .CLK(clk), .RST(rst), .Q(c[73]) );
  DFF \sreg_reg[76]  ( .D(c[76]), .CLK(clk), .RST(rst), .Q(c[72]) );
  DFF \sreg_reg[75]  ( .D(c[75]), .CLK(clk), .RST(rst), .Q(c[71]) );
  DFF \sreg_reg[74]  ( .D(c[74]), .CLK(clk), .RST(rst), .Q(c[70]) );
  DFF \sreg_reg[73]  ( .D(c[73]), .CLK(clk), .RST(rst), .Q(c[69]) );
  DFF \sreg_reg[72]  ( .D(c[72]), .CLK(clk), .RST(rst), .Q(c[68]) );
  DFF \sreg_reg[71]  ( .D(c[71]), .CLK(clk), .RST(rst), .Q(c[67]) );
  DFF \sreg_reg[70]  ( .D(c[70]), .CLK(clk), .RST(rst), .Q(c[66]) );
  DFF \sreg_reg[69]  ( .D(c[69]), .CLK(clk), .RST(rst), .Q(c[65]) );
  DFF \sreg_reg[68]  ( .D(c[68]), .CLK(clk), .RST(rst), .Q(c[64]) );
  DFF \sreg_reg[67]  ( .D(c[67]), .CLK(clk), .RST(rst), .Q(c[63]) );
  DFF \sreg_reg[66]  ( .D(c[66]), .CLK(clk), .RST(rst), .Q(c[62]) );
  DFF \sreg_reg[65]  ( .D(c[65]), .CLK(clk), .RST(rst), .Q(c[61]) );
  DFF \sreg_reg[64]  ( .D(c[64]), .CLK(clk), .RST(rst), .Q(c[60]) );
  DFF \sreg_reg[63]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[59]) );
  DFF \sreg_reg[62]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[58]) );
  DFF \sreg_reg[61]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[57]) );
  DFF \sreg_reg[60]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[56]) );
  DFF \sreg_reg[59]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[55]) );
  DFF \sreg_reg[58]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[54]) );
  DFF \sreg_reg[57]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[53]) );
  DFF \sreg_reg[56]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[52]) );
  DFF \sreg_reg[55]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[51]) );
  DFF \sreg_reg[54]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[50]) );
  DFF \sreg_reg[53]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[49]) );
  DFF \sreg_reg[52]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[48]) );
  DFF \sreg_reg[51]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[50]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[49]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[48]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[47]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[46]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[45]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[44]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[43]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[42]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[41]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[40]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[39]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[38]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[37]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[36]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[35]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[34]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[33]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[32]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[31]  ( .D(c[31]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[30]  ( .D(c[30]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[29]  ( .D(c[29]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[28]  ( .D(c[28]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[27]  ( .D(c[27]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[26]  ( .D(c[26]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[25]  ( .D(c[25]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[24]  ( .D(c[24]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[23]  ( .D(c[23]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[22]  ( .D(c[22]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[21]  ( .D(c[21]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[20]  ( .D(c[20]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[19]  ( .D(c[19]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[18]  ( .D(c[18]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[17]  ( .D(c[17]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[16]  ( .D(c[16]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[15]  ( .D(c[15]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[14]  ( .D(c[14]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[13]  ( .D(c[13]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[12]  ( .D(c[12]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[11]  ( .D(c[11]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[10]  ( .D(c[10]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[9]  ( .D(c[9]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[8]  ( .D(c[8]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[7]  ( .D(c[7]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[6]  ( .D(c[6]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[5]  ( .D(c[5]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[4]  ( .D(c[4]), .CLK(clk), .RST(rst), .Q(c[0]) );
  ADD_N1024_2 ADD_ ( .A({1'b0, 1'b0, 1'b0, 1'b0, sreg[2043:1024]}), .B(clocal), 
        .CI(1'b0), .S({swire, c[1023:1020]}) );
  mult_N1024_CC256_DW02_mult_0 mult_44 ( .A(b), .B(a), .TC(1'b0), .PRODUCT({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, clocal}) );
endmodule

