
module matrixMult_N_M_3_N8_M32 ( clk, rst, x, y, o );
  input [31:0] x;
  input [31:0] y;
  output [31:0] o;
  input clk, rst;
  wire   N33, N34, N35, N38, N40, N41, N42, N44, N45, N46, N47, N48, N49, N50,
         N51, N52, N53, N55, N57, N58, N59, N61, N62, N63, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
         n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
         n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
         n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
         n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
         n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
         n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
         n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
         n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
         n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
         n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
         n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
         n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
         n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
         n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
         n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
         n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
         n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
         n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
         n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
         n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
         n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
         n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
         n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
         n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
         n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
         n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
         n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
         n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
         n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
         n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
         n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224;

  DFF \o_reg[31]  ( .D(n6252), .CLK(clk), .RST(rst), .Q(o[31]) );
  DFF \o_reg[30]  ( .D(N63), .CLK(clk), .RST(rst), .Q(o[30]) );
  DFF \o_reg[29]  ( .D(N62), .CLK(clk), .RST(rst), .Q(o[29]) );
  DFF \o_reg[28]  ( .D(N61), .CLK(clk), .RST(rst), .Q(o[28]) );
  DFF \o_reg[27]  ( .D(n6253), .CLK(clk), .RST(rst), .Q(o[27]) );
  DFF \o_reg[26]  ( .D(N59), .CLK(clk), .RST(rst), .Q(o[26]) );
  DFF \o_reg[25]  ( .D(N58), .CLK(clk), .RST(rst), .Q(o[25]) );
  DFF \o_reg[24]  ( .D(N57), .CLK(clk), .RST(rst), .Q(o[24]) );
  DFF \o_reg[23]  ( .D(n6254), .CLK(clk), .RST(rst), .Q(o[23]) );
  DFF \o_reg[22]  ( .D(N55), .CLK(clk), .RST(rst), .Q(o[22]) );
  DFF \o_reg[21]  ( .D(n6255), .CLK(clk), .RST(rst), .Q(o[21]) );
  DFF \o_reg[20]  ( .D(N53), .CLK(clk), .RST(rst), .Q(o[20]) );
  DFF \o_reg[19]  ( .D(N52), .CLK(clk), .RST(rst), .Q(o[19]) );
  DFF \o_reg[18]  ( .D(N51), .CLK(clk), .RST(rst), .Q(o[18]) );
  DFF \o_reg[17]  ( .D(N50), .CLK(clk), .RST(rst), .Q(o[17]) );
  DFF \o_reg[16]  ( .D(N49), .CLK(clk), .RST(rst), .Q(o[16]) );
  DFF \o_reg[15]  ( .D(N48), .CLK(clk), .RST(rst), .Q(o[15]) );
  DFF \o_reg[14]  ( .D(N47), .CLK(clk), .RST(rst), .Q(o[14]) );
  DFF \o_reg[13]  ( .D(N46), .CLK(clk), .RST(rst), .Q(o[13]) );
  DFF \o_reg[12]  ( .D(N45), .CLK(clk), .RST(rst), .Q(o[12]) );
  DFF \o_reg[11]  ( .D(N44), .CLK(clk), .RST(rst), .Q(o[11]) );
  DFF \o_reg[10]  ( .D(n6256), .CLK(clk), .RST(rst), .Q(o[10]) );
  DFF \o_reg[9]  ( .D(N42), .CLK(clk), .RST(rst), .Q(o[9]) );
  DFF \o_reg[8]  ( .D(N41), .CLK(clk), .RST(rst), .Q(o[8]) );
  DFF \o_reg[7]  ( .D(N40), .CLK(clk), .RST(rst), .Q(o[7]) );
  DFF \o_reg[6]  ( .D(n6257), .CLK(clk), .RST(rst), .Q(o[6]) );
  DFF \o_reg[5]  ( .D(N38), .CLK(clk), .RST(rst), .Q(o[5]) );
  DFF \o_reg[4]  ( .D(n6258), .CLK(clk), .RST(rst), .Q(o[4]) );
  DFF \o_reg[3]  ( .D(n6259), .CLK(clk), .RST(rst), .Q(o[3]) );
  DFF \o_reg[2]  ( .D(N35), .CLK(clk), .RST(rst), .Q(o[2]) );
  DFF \o_reg[1]  ( .D(N34), .CLK(clk), .RST(rst), .Q(o[1]) );
  DFF \o_reg[0]  ( .D(N33), .CLK(clk), .RST(rst), .Q(o[0]) );
  NAND U3272 ( .A(n7487), .B(n7486), .Z(n6260) );
  NANDN U3273 ( .A(n7485), .B(n7484), .Z(n6261) );
  NAND U3274 ( .A(n6260), .B(n6261), .Z(n7595) );
  XNOR U3275 ( .A(n8895), .B(n8894), .Z(n8818) );
  XNOR U3276 ( .A(n7044), .B(n7043), .Z(n6998) );
  XNOR U3277 ( .A(n6827), .B(n6826), .Z(n6828) );
  XNOR U3278 ( .A(n6933), .B(n6932), .Z(n6936) );
  XOR U3279 ( .A(n7602), .B(n7601), .Z(n7598) );
  XNOR U3280 ( .A(n6644), .B(n6643), .Z(n6646) );
  XNOR U3281 ( .A(n8818), .B(n8817), .Z(n8899) );
  NAND U3282 ( .A(n8566), .B(n8565), .Z(n6262) );
  NANDN U3283 ( .A(n8564), .B(n8563), .Z(n6263) );
  AND U3284 ( .A(n6262), .B(n6263), .Z(n8734) );
  XNOR U3285 ( .A(n7086), .B(n7085), .Z(n7088) );
  XNOR U3286 ( .A(n7051), .B(n7050), .Z(n7001) );
  NAND U3287 ( .A(n7309), .B(n7308), .Z(n6264) );
  NAND U3288 ( .A(n7306), .B(n7307), .Z(n6265) );
  AND U3289 ( .A(n6264), .B(n6265), .Z(n7387) );
  XNOR U3290 ( .A(n7771), .B(n7770), .Z(n7773) );
  XNOR U3291 ( .A(n7755), .B(n7754), .Z(n7717) );
  XNOR U3292 ( .A(n6833), .B(n6832), .Z(n6843) );
  XNOR U3293 ( .A(n6838), .B(n6837), .Z(n6839) );
  XNOR U3294 ( .A(n7005), .B(n7004), .Z(n7006) );
  XNOR U3295 ( .A(n6894), .B(n6893), .Z(n6896) );
  NAND U3296 ( .A(n7444), .B(n7445), .Z(n6266) );
  NANDN U3297 ( .A(n7447), .B(n7446), .Z(n6267) );
  NAND U3298 ( .A(n6266), .B(n6267), .Z(n7534) );
  XNOR U3299 ( .A(n7070), .B(n7069), .Z(n7109) );
  XNOR U3300 ( .A(n8594), .B(n8593), .Z(n8579) );
  XOR U3301 ( .A(n8647), .B(n8646), .Z(n8588) );
  XNOR U3302 ( .A(n6939), .B(n6938), .Z(n6955) );
  XNOR U3303 ( .A(n7250), .B(n7249), .Z(n7251) );
  XNOR U3304 ( .A(n8901), .B(n8900), .Z(n8761) );
  NAND U3305 ( .A(n6410), .B(n6398), .Z(n6268) );
  NAND U3306 ( .A(n6382), .B(n6383), .Z(n6269) );
  AND U3307 ( .A(n6268), .B(n6269), .Z(n6385) );
  XNOR U3308 ( .A(n6404), .B(n6403), .Z(n6406) );
  NAND U3309 ( .A(n6642), .B(n6641), .Z(n6270) );
  NAND U3310 ( .A(n6639), .B(n6640), .Z(n6271) );
  AND U3311 ( .A(n6270), .B(n6271), .Z(n6649) );
  XOR U3312 ( .A(n6877), .B(n6876), .Z(n6881) );
  XNOR U3313 ( .A(n7057), .B(n7056), .Z(n6972) );
  XOR U3314 ( .A(n7945), .B(n7944), .Z(n6272) );
  NANDN U3315 ( .A(n7946), .B(n6272), .Z(n6273) );
  NAND U3316 ( .A(n7945), .B(n7944), .Z(n6274) );
  AND U3317 ( .A(n6273), .B(n6274), .Z(n7954) );
  XNOR U3318 ( .A(n8093), .B(n8092), .Z(n8095) );
  XNOR U3319 ( .A(n8953), .B(n8952), .Z(n8955) );
  XNOR U3320 ( .A(n8740), .B(n8739), .Z(n8733) );
  XOR U3321 ( .A(n9218), .B(n9217), .Z(n9216) );
  XNOR U3322 ( .A(n6855), .B(n6854), .Z(n6856) );
  XNOR U3323 ( .A(n7042), .B(n7041), .Z(n7043) );
  NAND U3324 ( .A(n7088), .B(n7087), .Z(n6275) );
  NANDN U3325 ( .A(n7086), .B(n7085), .Z(n6276) );
  AND U3326 ( .A(n6275), .B(n6276), .Z(n7204) );
  XNOR U3327 ( .A(n7495), .B(n7494), .Z(n7496) );
  XNOR U3328 ( .A(n6773), .B(n6772), .Z(n6774) );
  XNOR U3329 ( .A(n6756), .B(n6755), .Z(n6758) );
  XNOR U3330 ( .A(n6821), .B(n6820), .Z(n6822) );
  XNOR U3331 ( .A(n7019), .B(n7018), .Z(n7021) );
  XNOR U3332 ( .A(n6908), .B(n6907), .Z(n6900) );
  XNOR U3333 ( .A(n7436), .B(n7435), .Z(n7415) );
  NAND U3334 ( .A(n7313), .B(n7312), .Z(n6277) );
  NAND U3335 ( .A(n7310), .B(n7311), .Z(n6278) );
  AND U3336 ( .A(n6277), .B(n6278), .Z(n7389) );
  XOR U3337 ( .A(n7330), .B(n7329), .Z(n7332) );
  NAND U3338 ( .A(n7443), .B(n7442), .Z(n6279) );
  NAND U3339 ( .A(n7440), .B(n7441), .Z(n6280) );
  NAND U3340 ( .A(n6279), .B(n6280), .Z(n7535) );
  NAND U3341 ( .A(n7717), .B(n7718), .Z(n6281) );
  NANDN U3342 ( .A(n7720), .B(n7719), .Z(n6282) );
  AND U3343 ( .A(n6281), .B(n6282), .Z(n7883) );
  NAND U3344 ( .A(n7614), .B(n7613), .Z(n6283) );
  NANDN U3345 ( .A(n7612), .B(n7611), .Z(n6284) );
  AND U3346 ( .A(n6283), .B(n6284), .Z(n7712) );
  NAND U3347 ( .A(n7919), .B(n7918), .Z(n6285) );
  NANDN U3348 ( .A(n7917), .B(n7916), .Z(n6286) );
  AND U3349 ( .A(n6285), .B(n6286), .Z(n8074) );
  NAND U3350 ( .A(n7095), .B(n6628), .Z(n6287) );
  NANDN U3351 ( .A(n6528), .B(n6527), .Z(n6288) );
  AND U3352 ( .A(n6287), .B(n6288), .Z(n6575) );
  XNOR U3353 ( .A(n6937), .B(n6936), .Z(n6938) );
  XNOR U3354 ( .A(n6809), .B(n6808), .Z(n6811) );
  XOR U3355 ( .A(n7142), .B(n7141), .Z(n7111) );
  NAND U3356 ( .A(n7774), .B(n7775), .Z(n6289) );
  NANDN U3357 ( .A(n7777), .B(n7776), .Z(n6290) );
  NAND U3358 ( .A(n6289), .B(n6290), .Z(n7877) );
  NAND U3359 ( .A(n8143), .B(n8142), .Z(n6291) );
  NANDN U3360 ( .A(n8141), .B(n8140), .Z(n6292) );
  AND U3361 ( .A(n6291), .B(n6292), .Z(n8301) );
  XNOR U3362 ( .A(n8586), .B(n8585), .Z(n8587) );
  XNOR U3363 ( .A(n8639), .B(n8638), .Z(n8641) );
  XOR U3364 ( .A(n6951), .B(n6950), .Z(n6888) );
  XNOR U3365 ( .A(n7256), .B(n7255), .Z(n7257) );
  XNOR U3366 ( .A(n8816), .B(n8815), .Z(n8817) );
  XNOR U3367 ( .A(n8800), .B(n8799), .Z(n8804) );
  XNOR U3368 ( .A(n8582), .B(n8581), .Z(n8568) );
  XOR U3369 ( .A(n6456), .B(n6457), .Z(n6293) );
  NANDN U3370 ( .A(n6458), .B(n6293), .Z(n6294) );
  NAND U3371 ( .A(n6456), .B(n6457), .Z(n6295) );
  AND U3372 ( .A(n6294), .B(n6295), .Z(n6459) );
  NAND U3373 ( .A(n8913), .B(n8910), .Z(n6296) );
  NANDN U3374 ( .A(n8913), .B(n6649), .Z(n6297) );
  NANDN U3375 ( .A(n8911), .B(n6297), .Z(n6298) );
  NAND U3376 ( .A(n6296), .B(n6298), .Z(n6726) );
  XOR U3377 ( .A(n6972), .B(n6971), .Z(n6974) );
  XNOR U3378 ( .A(n7252), .B(n7251), .Z(n7160) );
  NAND U3379 ( .A(n7466), .B(n7467), .Z(n6299) );
  NANDN U3380 ( .A(n7469), .B(n7468), .Z(n6300) );
  NAND U3381 ( .A(n6299), .B(n6300), .Z(n7590) );
  NAND U3382 ( .A(n7962), .B(n7961), .Z(n6301) );
  NAND U3383 ( .A(n7959), .B(n7960), .Z(n6302) );
  AND U3384 ( .A(n6301), .B(n6302), .Z(n8236) );
  XNOR U3385 ( .A(n8770), .B(n8769), .Z(n8895) );
  XNOR U3386 ( .A(n8963), .B(n8962), .Z(n8961) );
  NAND U3387 ( .A(n6963), .B(n6960), .Z(n6303) );
  NANDN U3388 ( .A(n6963), .B(n6962), .Z(n6304) );
  NANDN U3389 ( .A(n6961), .B(n6304), .Z(n6305) );
  NAND U3390 ( .A(n6303), .B(n6305), .Z(n6977) );
  XNOR U3391 ( .A(n7950), .B(n7949), .Z(n7945) );
  NAND U3392 ( .A(n8736), .B(n8735), .Z(n6306) );
  NAND U3393 ( .A(n8733), .B(n8734), .Z(n6307) );
  AND U3394 ( .A(n6306), .B(n6307), .Z(n8922) );
  XNOR U3395 ( .A(n6906), .B(n6905), .Z(n6907) );
  XNOR U3396 ( .A(n6912), .B(n6911), .Z(n6913) );
  XNOR U3397 ( .A(n6999), .B(n6998), .Z(n7000) );
  NAND U3398 ( .A(n7773), .B(n7772), .Z(n6308) );
  NANDN U3399 ( .A(n7771), .B(n7770), .Z(n6309) );
  NAND U3400 ( .A(n6308), .B(n6309), .Z(n7846) );
  NAND U3401 ( .A(n7985), .B(n7986), .Z(n6310) );
  NANDN U3402 ( .A(n7988), .B(n7987), .Z(n6311) );
  NAND U3403 ( .A(n6310), .B(n6311), .Z(n8134) );
  XNOR U3404 ( .A(n6630), .B(n6629), .Z(n6605) );
  XNOR U3405 ( .A(n6683), .B(n6682), .Z(n6684) );
  XNOR U3406 ( .A(n6763), .B(o[12]), .Z(n6775) );
  XNOR U3407 ( .A(n6688), .B(o[11]), .Z(n6697) );
  XNOR U3408 ( .A(n6836), .B(o[13]), .Z(n6829) );
  XNOR U3409 ( .A(n7049), .B(n7048), .Z(n7050) );
  XNOR U3410 ( .A(n6931), .B(n6930), .Z(n6932) );
  XNOR U3411 ( .A(n7140), .B(n7139), .Z(n7141) );
  NAND U3412 ( .A(n7321), .B(n7320), .Z(n6312) );
  NAND U3413 ( .A(n7319), .B(n7318), .Z(n6313) );
  NAND U3414 ( .A(n6312), .B(n6313), .Z(n7446) );
  NAND U3415 ( .A(n7317), .B(n7316), .Z(n6314) );
  NAND U3416 ( .A(n7314), .B(n7315), .Z(n6315) );
  AND U3417 ( .A(n6314), .B(n6315), .Z(n7417) );
  NAND U3418 ( .A(n7293), .B(n7292), .Z(n6316) );
  NANDN U3419 ( .A(n7291), .B(n7290), .Z(n6317) );
  NAND U3420 ( .A(n6316), .B(n6317), .Z(n7442) );
  NAND U3421 ( .A(n7224), .B(n7223), .Z(n6318) );
  NANDN U3422 ( .A(n7222), .B(n7221), .Z(n6319) );
  AND U3423 ( .A(n6318), .B(n6319), .Z(n7335) );
  NAND U3424 ( .A(n7389), .B(n7388), .Z(n6320) );
  NAND U3425 ( .A(n7387), .B(n7386), .Z(n6321) );
  NAND U3426 ( .A(n6320), .B(n6321), .Z(n7573) );
  NAND U3427 ( .A(n7975), .B(n7976), .Z(n6322) );
  NANDN U3428 ( .A(n7978), .B(n7977), .Z(n6323) );
  AND U3429 ( .A(n6322), .B(n6323), .Z(n8141) );
  XNOR U3430 ( .A(n8341), .B(n8340), .Z(n8343) );
  XOR U3431 ( .A(n8467), .B(n8466), .Z(n8469) );
  NAND U3432 ( .A(n6618), .B(n6617), .Z(n6324) );
  NANDN U3433 ( .A(n7495), .B(n7024), .Z(n6325) );
  NAND U3434 ( .A(n6324), .B(n6325), .Z(n6715) );
  XNOR U3435 ( .A(n6752), .B(n6751), .Z(n6745) );
  XNOR U3436 ( .A(n6823), .B(n6822), .Z(n6814) );
  XNOR U3437 ( .A(n6949), .B(n6948), .Z(n6950) );
  XNOR U3438 ( .A(n6840), .B(n6839), .Z(n6808) );
  XOR U3439 ( .A(n7076), .B(n7075), .Z(n7067) );
  XNOR U3440 ( .A(n7007), .B(n7006), .Z(n6993) );
  XOR U3441 ( .A(n6989), .B(n6988), .Z(n7055) );
  NAND U3442 ( .A(n7524), .B(n7525), .Z(n6326) );
  NANDN U3443 ( .A(n7527), .B(n7526), .Z(n6327) );
  AND U3444 ( .A(n6326), .B(n6327), .Z(n7693) );
  NAND U3445 ( .A(n7630), .B(n7629), .Z(n6328) );
  NANDN U3446 ( .A(n7628), .B(n7627), .Z(n6329) );
  AND U3447 ( .A(n6328), .B(n6329), .Z(n7809) );
  NAND U3448 ( .A(n7885), .B(n7884), .Z(n6330) );
  NANDN U3449 ( .A(n7883), .B(n7882), .Z(n6331) );
  AND U3450 ( .A(n6330), .B(n6331), .Z(n8077) );
  NAND U3451 ( .A(n7799), .B(n7798), .Z(n6332) );
  NAND U3452 ( .A(n7797), .B(n7796), .Z(n6333) );
  NAND U3453 ( .A(n6332), .B(n6333), .Z(n7932) );
  XNOR U3454 ( .A(n8580), .B(n8579), .Z(n8581) );
  XOR U3455 ( .A(n6846), .B(n6845), .Z(n6871) );
  XOR U3456 ( .A(n6955), .B(n6954), .Z(n6957) );
  XNOR U3457 ( .A(n7355), .B(n7354), .Z(n7357) );
  NAND U3458 ( .A(n7271), .B(n7270), .Z(n6334) );
  NAND U3459 ( .A(n7268), .B(n7269), .Z(n6335) );
  AND U3460 ( .A(n6334), .B(n6335), .Z(n7467) );
  XNOR U3461 ( .A(n8812), .B(n8811), .Z(n8750) );
  XNOR U3462 ( .A(n8995), .B(n8994), .Z(n8993) );
  XNOR U3463 ( .A(n9176), .B(n9175), .Z(n9178) );
  XNOR U3464 ( .A(n8804), .B(n8803), .Z(n8806) );
  XNOR U3465 ( .A(n8786), .B(n8785), .Z(n8788) );
  XNOR U3466 ( .A(n8618), .B(n8617), .Z(n8570) );
  NAND U3467 ( .A(n8554), .B(n8553), .Z(n6336) );
  NAND U3468 ( .A(n8296), .B(n8297), .Z(n6337) );
  AND U3469 ( .A(n6336), .B(n6337), .Z(n8564) );
  XOR U3470 ( .A(n6653), .B(n6652), .Z(n6645) );
  XNOR U3471 ( .A(n6875), .B(n6874), .Z(n6876) );
  XOR U3472 ( .A(n7160), .B(n7159), .Z(n7162) );
  NAND U3473 ( .A(n7595), .B(n7596), .Z(n6338) );
  NANDN U3474 ( .A(n7598), .B(n7597), .Z(n6339) );
  NAND U3475 ( .A(n6338), .B(n6339), .Z(n7949) );
  NAND U3476 ( .A(n8238), .B(n8237), .Z(n6340) );
  NAND U3477 ( .A(n8235), .B(n8236), .Z(n6341) );
  AND U3478 ( .A(n6340), .B(n6341), .Z(n8527) );
  XNOR U3479 ( .A(n8893), .B(n8892), .Z(n8894) );
  XNOR U3480 ( .A(n9200), .B(n9199), .Z(n9198) );
  XNOR U3481 ( .A(n8946), .B(n8947), .Z(n8949) );
  XOR U3482 ( .A(n8744), .B(n8743), .Z(n8746) );
  NAND U3483 ( .A(n8907), .B(n8906), .Z(n6342) );
  NAND U3484 ( .A(n6384), .B(n6385), .Z(n6343) );
  AND U3485 ( .A(n6342), .B(n6343), .Z(n6456) );
  XOR U3486 ( .A(n6516), .B(n6515), .Z(n6344) );
  NANDN U3487 ( .A(n6517), .B(n6344), .Z(n6345) );
  NAND U3488 ( .A(n6516), .B(n6515), .Z(n6346) );
  AND U3489 ( .A(n6345), .B(n6346), .Z(n6642) );
  XOR U3490 ( .A(n6977), .B(n6978), .Z(n6347) );
  NANDN U3491 ( .A(n6979), .B(n6347), .Z(n6348) );
  NAND U3492 ( .A(n6977), .B(n6978), .Z(n6349) );
  AND U3493 ( .A(n6348), .B(n6349), .Z(n7147) );
  NAND U3494 ( .A(n8915), .B(n8914), .Z(n6350) );
  NAND U3495 ( .A(n7587), .B(n7588), .Z(n6351) );
  NAND U3496 ( .A(n6350), .B(n6351), .Z(n7944) );
  XNOR U3497 ( .A(n8923), .B(n8922), .Z(n8921) );
  AND U3498 ( .A(x[0]), .B(y[0]), .Z(n7024) );
  XOR U3499 ( .A(n7024), .B(o[0]), .Z(N33) );
  NAND U3500 ( .A(x[1]), .B(y[0]), .Z(n6387) );
  AND U3501 ( .A(x[0]), .B(y[1]), .Z(n6354) );
  XNOR U3502 ( .A(n6354), .B(o[1]), .Z(n6357) );
  XOR U3503 ( .A(n6387), .B(n6357), .Z(n6356) );
  NAND U3504 ( .A(n7024), .B(o[0]), .Z(n6355) );
  XNOR U3505 ( .A(n6356), .B(n6355), .Z(N34) );
  AND U3506 ( .A(y[2]), .B(x[0]), .Z(n6377) );
  XOR U3507 ( .A(n6377), .B(o[2]), .Z(n6393) );
  AND U3508 ( .A(y[0]), .B(x[2]), .Z(n6353) );
  NAND U3509 ( .A(y[1]), .B(x[1]), .Z(n6352) );
  XNOR U3510 ( .A(n6353), .B(n6352), .Z(n6389) );
  AND U3511 ( .A(n6354), .B(o[1]), .Z(n6388) );
  XNOR U3512 ( .A(n6389), .B(n6388), .Z(n6392) );
  XNOR U3513 ( .A(n6393), .B(n6392), .Z(n6395) );
  AND U3514 ( .A(n6356), .B(n6355), .Z(n6359) );
  NAND U3515 ( .A(n6387), .B(n6357), .Z(n6358) );
  NANDN U3516 ( .A(n6359), .B(n6358), .Z(n6394) );
  XNOR U3517 ( .A(n6395), .B(n6394), .Z(N35) );
  NAND U3518 ( .A(x[3]), .B(y[1]), .Z(n6364) );
  ANDN U3519 ( .B(o[4]), .A(n6364), .Z(n6422) );
  AND U3520 ( .A(y[0]), .B(x[5]), .Z(n6361) );
  NAND U3521 ( .A(x[0]), .B(y[5]), .Z(n6360) );
  XNOR U3522 ( .A(n6361), .B(n6360), .Z(n6421) );
  XOR U3523 ( .A(n6422), .B(n6421), .Z(n6418) );
  AND U3524 ( .A(y[3]), .B(x[2]), .Z(n6416) );
  NAND U3525 ( .A(x[4]), .B(y[1]), .Z(n6425) );
  XNOR U3526 ( .A(o[5]), .B(n6425), .Z(n6412) );
  AND U3527 ( .A(y[4]), .B(x[1]), .Z(n6363) );
  NAND U3528 ( .A(y[2]), .B(x[3]), .Z(n6362) );
  XNOR U3529 ( .A(n6363), .B(n6362), .Z(n6411) );
  XNOR U3530 ( .A(n6412), .B(n6411), .Z(n6415) );
  XNOR U3531 ( .A(n6416), .B(n6415), .Z(n6417) );
  XOR U3532 ( .A(n6418), .B(n6417), .Z(n6463) );
  AND U3533 ( .A(x[1]), .B(y[3]), .Z(n6586) );
  AND U3534 ( .A(y[2]), .B(x[2]), .Z(n6531) );
  NAND U3535 ( .A(n6586), .B(n6531), .Z(n6366) );
  XNOR U3536 ( .A(o[4]), .B(n6364), .Z(n6372) );
  XOR U3537 ( .A(n6586), .B(n6531), .Z(n6371) );
  NAND U3538 ( .A(n6372), .B(n6371), .Z(n6365) );
  NAND U3539 ( .A(n6366), .B(n6365), .Z(n6462) );
  AND U3540 ( .A(x[4]), .B(y[0]), .Z(n6368) );
  AND U3541 ( .A(y[4]), .B(x[0]), .Z(n6367) );
  NAND U3542 ( .A(n6368), .B(n6367), .Z(n6370) );
  AND U3543 ( .A(x[2]), .B(y[1]), .Z(n6386) );
  AND U3544 ( .A(n6386), .B(o[3]), .Z(n6374) );
  XOR U3545 ( .A(n6368), .B(n6367), .Z(n6373) );
  NAND U3546 ( .A(n6374), .B(n6373), .Z(n6369) );
  NAND U3547 ( .A(n6370), .B(n6369), .Z(n6461) );
  XNOR U3548 ( .A(n6462), .B(n6461), .Z(n6464) );
  XOR U3549 ( .A(n6463), .B(n6464), .Z(n6458) );
  XOR U3550 ( .A(n6372), .B(n6371), .Z(n6404) );
  XNOR U3551 ( .A(n6374), .B(n6373), .Z(n6403) );
  AND U3552 ( .A(y[3]), .B(x[0]), .Z(n6376) );
  AND U3553 ( .A(x[3]), .B(y[0]), .Z(n6375) );
  NAND U3554 ( .A(n6376), .B(n6375), .Z(n6379) );
  XOR U3555 ( .A(n6376), .B(n6375), .Z(n6381) );
  AND U3556 ( .A(n6377), .B(o[2]), .Z(n6380) );
  NAND U3557 ( .A(n6381), .B(n6380), .Z(n6378) );
  AND U3558 ( .A(n6379), .B(n6378), .Z(n6405) );
  XOR U3559 ( .A(n6406), .B(n6405), .Z(n6384) );
  XOR U3560 ( .A(n6381), .B(n6380), .Z(n6382) );
  XOR U3561 ( .A(o[3]), .B(n6386), .Z(n6383) );
  XOR U3562 ( .A(n6383), .B(n6382), .Z(n6398) );
  AND U3563 ( .A(y[2]), .B(x[1]), .Z(n6410) );
  XOR U3564 ( .A(n6385), .B(n6384), .Z(n8907) );
  NANDN U3565 ( .A(n6387), .B(n6386), .Z(n6391) );
  NAND U3566 ( .A(n6389), .B(n6388), .Z(n6390) );
  AND U3567 ( .A(n6391), .B(n6390), .Z(n6400) );
  NANDN U3568 ( .A(n6393), .B(n6392), .Z(n6397) );
  NAND U3569 ( .A(n6395), .B(n6394), .Z(n6396) );
  AND U3570 ( .A(n6397), .B(n6396), .Z(n6399) );
  NANDN U3571 ( .A(n6400), .B(n6399), .Z(n6402) );
  XOR U3572 ( .A(n6410), .B(n6398), .Z(n8905) );
  XNOR U3573 ( .A(n6400), .B(n6399), .Z(n8904) );
  NAND U3574 ( .A(n8905), .B(n8904), .Z(n6401) );
  AND U3575 ( .A(n6402), .B(n6401), .Z(n8906) );
  NANDN U3576 ( .A(n6404), .B(n6403), .Z(n6408) );
  NAND U3577 ( .A(n6406), .B(n6405), .Z(n6407) );
  AND U3578 ( .A(n6408), .B(n6407), .Z(n6457) );
  XOR U3579 ( .A(n6456), .B(n6457), .Z(n6409) );
  XNOR U3580 ( .A(n6458), .B(n6409), .Z(N38) );
  AND U3581 ( .A(x[3]), .B(y[4]), .Z(n6490) );
  NAND U3582 ( .A(n6490), .B(n6410), .Z(n6414) );
  NAND U3583 ( .A(n6412), .B(n6411), .Z(n6413) );
  AND U3584 ( .A(n6414), .B(n6413), .Z(n6427) );
  NANDN U3585 ( .A(n6416), .B(n6415), .Z(n6420) );
  NANDN U3586 ( .A(n6418), .B(n6417), .Z(n6419) );
  AND U3587 ( .A(n6420), .B(n6419), .Z(n6426) );
  NANDN U3588 ( .A(n6427), .B(n6426), .Z(n6429) );
  AND U3589 ( .A(y[5]), .B(x[5]), .Z(n6635) );
  NAND U3590 ( .A(n7024), .B(n6635), .Z(n6424) );
  NAND U3591 ( .A(n6422), .B(n6421), .Z(n6423) );
  AND U3592 ( .A(n6424), .B(n6423), .Z(n6449) );
  ANDN U3593 ( .B(o[5]), .A(n6425), .Z(n6437) );
  AND U3594 ( .A(x[0]), .B(y[6]), .Z(n6435) );
  NAND U3595 ( .A(x[6]), .B(y[0]), .Z(n6436) );
  XOR U3596 ( .A(n6435), .B(n6436), .Z(n6438) );
  XNOR U3597 ( .A(n6437), .B(n6438), .Z(n6448) );
  XNOR U3598 ( .A(n6449), .B(n6448), .Z(n6450) );
  NAND U3599 ( .A(x[5]), .B(y[1]), .Z(n6447) );
  XNOR U3600 ( .A(o[6]), .B(n6447), .Z(n6444) );
  AND U3601 ( .A(y[5]), .B(x[1]), .Z(n6441) );
  NAND U3602 ( .A(y[2]), .B(x[4]), .Z(n6442) );
  XNOR U3603 ( .A(n6441), .B(n6442), .Z(n6443) );
  XOR U3604 ( .A(n6444), .B(n6443), .Z(n6431) );
  AND U3605 ( .A(x[2]), .B(y[4]), .Z(n6925) );
  NAND U3606 ( .A(x[3]), .B(y[3]), .Z(n6430) );
  XOR U3607 ( .A(n6925), .B(n6430), .Z(n6432) );
  XOR U3608 ( .A(n6431), .B(n6432), .Z(n6451) );
  XNOR U3609 ( .A(n6450), .B(n6451), .Z(n6455) );
  XNOR U3610 ( .A(n6427), .B(n6426), .Z(n6454) );
  NAND U3611 ( .A(n6455), .B(n6454), .Z(n6428) );
  AND U3612 ( .A(n6429), .B(n6428), .Z(n6508) );
  NAND U3613 ( .A(x[6]), .B(y[1]), .Z(n6475) );
  XNOR U3614 ( .A(o[7]), .B(n6475), .Z(n6470) );
  AND U3615 ( .A(x[1]), .B(y[6]), .Z(n6849) );
  AND U3616 ( .A(x[5]), .B(y[2]), .Z(n6596) );
  XOR U3617 ( .A(n6849), .B(n6596), .Z(n6469) );
  XOR U3618 ( .A(n6470), .B(n6469), .Z(n6483) );
  NANDN U3619 ( .A(n6430), .B(n6925), .Z(n6434) );
  NANDN U3620 ( .A(n6432), .B(n6431), .Z(n6433) );
  AND U3621 ( .A(n6434), .B(n6433), .Z(n6482) );
  XNOR U3622 ( .A(n6483), .B(n6482), .Z(n6484) );
  NANDN U3623 ( .A(n6436), .B(n6435), .Z(n6440) );
  NANDN U3624 ( .A(n6438), .B(n6437), .Z(n6439) );
  NAND U3625 ( .A(n6440), .B(n6439), .Z(n6485) );
  XNOR U3626 ( .A(n6484), .B(n6485), .Z(n6502) );
  NANDN U3627 ( .A(n6442), .B(n6441), .Z(n6446) );
  NAND U3628 ( .A(n6444), .B(n6443), .Z(n6445) );
  AND U3629 ( .A(n6446), .B(n6445), .Z(n6478) );
  AND U3630 ( .A(y[7]), .B(x[0]), .Z(n6494) );
  AND U3631 ( .A(x[7]), .B(y[0]), .Z(n6495) );
  XOR U3632 ( .A(n6494), .B(n6495), .Z(n6497) );
  ANDN U3633 ( .B(o[6]), .A(n6447), .Z(n6496) );
  XOR U3634 ( .A(n6497), .B(n6496), .Z(n6477) );
  AND U3635 ( .A(y[5]), .B(x[2]), .Z(n6488) );
  AND U3636 ( .A(y[3]), .B(x[4]), .Z(n6489) );
  XOR U3637 ( .A(n6488), .B(n6489), .Z(n6491) );
  XNOR U3638 ( .A(n6491), .B(n6490), .Z(n6476) );
  XOR U3639 ( .A(n6477), .B(n6476), .Z(n6479) );
  XOR U3640 ( .A(n6478), .B(n6479), .Z(n6503) );
  XNOR U3641 ( .A(n6502), .B(n6503), .Z(n6504) );
  NANDN U3642 ( .A(n6449), .B(n6448), .Z(n6453) );
  NANDN U3643 ( .A(n6451), .B(n6450), .Z(n6452) );
  NAND U3644 ( .A(n6453), .B(n6452), .Z(n6505) );
  XOR U3645 ( .A(n6504), .B(n6505), .Z(n6509) );
  XNOR U3646 ( .A(n6508), .B(n6509), .Z(n6511) );
  XOR U3647 ( .A(n6455), .B(n6454), .Z(n6460) );
  NANDN U3648 ( .A(n6460), .B(n6459), .Z(n6468) );
  XNOR U3649 ( .A(n6460), .B(n6459), .Z(n8909) );
  NAND U3650 ( .A(n6462), .B(n6461), .Z(n6466) );
  NANDN U3651 ( .A(n6464), .B(n6463), .Z(n6465) );
  AND U3652 ( .A(n6466), .B(n6465), .Z(n8908) );
  NAND U3653 ( .A(n8909), .B(n8908), .Z(n6467) );
  NAND U3654 ( .A(n6468), .B(n6467), .Z(n6510) );
  XNOR U3655 ( .A(n6511), .B(n6510), .Z(N40) );
  NAND U3656 ( .A(n6596), .B(n6849), .Z(n6472) );
  NAND U3657 ( .A(n6470), .B(n6469), .Z(n6471) );
  AND U3658 ( .A(n6472), .B(n6471), .Z(n6543) );
  NAND U3659 ( .A(x[3]), .B(y[5]), .Z(n6537) );
  AND U3660 ( .A(y[6]), .B(x[2]), .Z(n6474) );
  NAND U3661 ( .A(x[6]), .B(y[2]), .Z(n6473) );
  XNOR U3662 ( .A(n6474), .B(n6473), .Z(n6533) );
  AND U3663 ( .A(y[4]), .B(x[4]), .Z(n6532) );
  XNOR U3664 ( .A(n6533), .B(n6532), .Z(n6536) );
  XOR U3665 ( .A(n6537), .B(n6536), .Z(n6539) );
  ANDN U3666 ( .B(o[7]), .A(n6475), .Z(n6528) );
  NAND U3667 ( .A(x[5]), .B(y[3]), .Z(n7095) );
  NAND U3668 ( .A(y[7]), .B(x[1]), .Z(n6628) );
  XOR U3669 ( .A(n7095), .B(n6628), .Z(n6527) );
  XNOR U3670 ( .A(n6528), .B(n6527), .Z(n6538) );
  XNOR U3671 ( .A(n6539), .B(n6538), .Z(n6542) );
  XNOR U3672 ( .A(n6543), .B(n6542), .Z(n6545) );
  NANDN U3673 ( .A(n6477), .B(n6476), .Z(n6481) );
  NANDN U3674 ( .A(n6479), .B(n6478), .Z(n6480) );
  AND U3675 ( .A(n6481), .B(n6480), .Z(n6544) );
  XOR U3676 ( .A(n6545), .B(n6544), .Z(n6556) );
  NANDN U3677 ( .A(n6483), .B(n6482), .Z(n6487) );
  NANDN U3678 ( .A(n6485), .B(n6484), .Z(n6486) );
  AND U3679 ( .A(n6487), .B(n6486), .Z(n6555) );
  NAND U3680 ( .A(n6489), .B(n6488), .Z(n6493) );
  NAND U3681 ( .A(n6491), .B(n6490), .Z(n6492) );
  AND U3682 ( .A(n6493), .B(n6492), .Z(n6551) );
  NAND U3683 ( .A(n6495), .B(n6494), .Z(n6499) );
  NAND U3684 ( .A(n6497), .B(n6496), .Z(n6498) );
  AND U3685 ( .A(n6499), .B(n6498), .Z(n6549) );
  NAND U3686 ( .A(x[7]), .B(y[1]), .Z(n6526) );
  XNOR U3687 ( .A(o[8]), .B(n6526), .Z(n6518) );
  AND U3688 ( .A(x[8]), .B(y[0]), .Z(n6501) );
  NAND U3689 ( .A(x[0]), .B(y[8]), .Z(n6500) );
  XOR U3690 ( .A(n6501), .B(n6500), .Z(n6519) );
  XNOR U3691 ( .A(n6518), .B(n6519), .Z(n6548) );
  XNOR U3692 ( .A(n6549), .B(n6548), .Z(n6550) );
  XOR U3693 ( .A(n6551), .B(n6550), .Z(n6554) );
  XOR U3694 ( .A(n6555), .B(n6554), .Z(n6557) );
  XOR U3695 ( .A(n6556), .B(n6557), .Z(n6516) );
  NANDN U3696 ( .A(n6503), .B(n6502), .Z(n6507) );
  NANDN U3697 ( .A(n6505), .B(n6504), .Z(n6506) );
  NAND U3698 ( .A(n6507), .B(n6506), .Z(n6515) );
  NANDN U3699 ( .A(n6509), .B(n6508), .Z(n6513) );
  NAND U3700 ( .A(n6511), .B(n6510), .Z(n6512) );
  AND U3701 ( .A(n6513), .B(n6512), .Z(n6517) );
  XOR U3702 ( .A(n6515), .B(n6517), .Z(n6514) );
  XOR U3703 ( .A(n6516), .B(n6514), .Z(N41) );
  NAND U3704 ( .A(y[8]), .B(x[8]), .Z(n7086) );
  NANDN U3705 ( .A(n7086), .B(n7024), .Z(n6521) );
  NANDN U3706 ( .A(n6519), .B(n6518), .Z(n6520) );
  AND U3707 ( .A(n6521), .B(n6520), .Z(n6568) );
  NAND U3708 ( .A(y[1]), .B(x[8]), .Z(n6595) );
  XNOR U3709 ( .A(o[9]), .B(n6595), .Z(n6583) );
  AND U3710 ( .A(x[9]), .B(y[0]), .Z(n6523) );
  NAND U3711 ( .A(y[9]), .B(x[0]), .Z(n6522) );
  XNOR U3712 ( .A(n6523), .B(n6522), .Z(n6582) );
  XOR U3713 ( .A(n6583), .B(n6582), .Z(n6567) );
  AND U3714 ( .A(x[7]), .B(y[2]), .Z(n6525) );
  NAND U3715 ( .A(y[4]), .B(x[5]), .Z(n6524) );
  XNOR U3716 ( .A(n6525), .B(n6524), .Z(n6598) );
  ANDN U3717 ( .B(o[8]), .A(n6526), .Z(n6597) );
  XNOR U3718 ( .A(n6598), .B(n6597), .Z(n6566) );
  XOR U3719 ( .A(n6567), .B(n6566), .Z(n6569) );
  XNOR U3720 ( .A(n6568), .B(n6569), .Z(n6576) );
  AND U3721 ( .A(y[3]), .B(x[6]), .Z(n6530) );
  NAND U3722 ( .A(x[1]), .B(y[8]), .Z(n6529) );
  XNOR U3723 ( .A(n6530), .B(n6529), .Z(n6588) );
  AND U3724 ( .A(y[5]), .B(x[4]), .Z(n6587) );
  XOR U3725 ( .A(n6588), .B(n6587), .Z(n6563) );
  AND U3726 ( .A(y[7]), .B(x[2]), .Z(n6561) );
  NAND U3727 ( .A(x[3]), .B(y[6]), .Z(n6560) );
  XNOR U3728 ( .A(n6561), .B(n6560), .Z(n6562) );
  XNOR U3729 ( .A(n6563), .B(n6562), .Z(n6574) );
  XOR U3730 ( .A(n6575), .B(n6574), .Z(n6577) );
  XOR U3731 ( .A(n6576), .B(n6577), .Z(n6652) );
  AND U3732 ( .A(x[6]), .B(y[6]), .Z(n6779) );
  NAND U3733 ( .A(n6779), .B(n6531), .Z(n6535) );
  NAND U3734 ( .A(n6533), .B(n6532), .Z(n6534) );
  NAND U3735 ( .A(n6535), .B(n6534), .Z(n6650) );
  NAND U3736 ( .A(n6537), .B(n6536), .Z(n6541) );
  NAND U3737 ( .A(n6539), .B(n6538), .Z(n6540) );
  AND U3738 ( .A(n6541), .B(n6540), .Z(n6651) );
  XNOR U3739 ( .A(n6650), .B(n6651), .Z(n6653) );
  NANDN U3740 ( .A(n6543), .B(n6542), .Z(n6547) );
  NAND U3741 ( .A(n6545), .B(n6544), .Z(n6546) );
  AND U3742 ( .A(n6547), .B(n6546), .Z(n6643) );
  NANDN U3743 ( .A(n6549), .B(n6548), .Z(n6553) );
  NANDN U3744 ( .A(n6551), .B(n6550), .Z(n6552) );
  NAND U3745 ( .A(n6553), .B(n6552), .Z(n6644) );
  XNOR U3746 ( .A(n6645), .B(n6646), .Z(n6639) );
  NANDN U3747 ( .A(n6555), .B(n6554), .Z(n6559) );
  OR U3748 ( .A(n6557), .B(n6556), .Z(n6558) );
  AND U3749 ( .A(n6559), .B(n6558), .Z(n6640) );
  XOR U3750 ( .A(n6639), .B(n6640), .Z(n6641) );
  XOR U3751 ( .A(n6642), .B(n6641), .Z(N42) );
  NANDN U3752 ( .A(n6561), .B(n6560), .Z(n6565) );
  NANDN U3753 ( .A(n6563), .B(n6562), .Z(n6564) );
  AND U3754 ( .A(n6565), .B(n6564), .Z(n6573) );
  NANDN U3755 ( .A(n6567), .B(n6566), .Z(n6571) );
  NANDN U3756 ( .A(n6569), .B(n6568), .Z(n6570) );
  NAND U3757 ( .A(n6571), .B(n6570), .Z(n6572) );
  NANDN U3758 ( .A(n6573), .B(n6572), .Z(n6581) );
  XOR U3759 ( .A(n6573), .B(n6572), .Z(n6658) );
  NANDN U3760 ( .A(n6575), .B(n6574), .Z(n6579) );
  NANDN U3761 ( .A(n6577), .B(n6576), .Z(n6578) );
  AND U3762 ( .A(n6579), .B(n6578), .Z(n6659) );
  OR U3763 ( .A(n6658), .B(n6659), .Z(n6580) );
  AND U3764 ( .A(n6581), .B(n6580), .Z(n6722) );
  AND U3765 ( .A(x[9]), .B(y[9]), .Z(n7178) );
  IV U3766 ( .A(n7178), .Z(n7291) );
  NANDN U3767 ( .A(n7291), .B(n7024), .Z(n6585) );
  NAND U3768 ( .A(n6583), .B(n6582), .Z(n6584) );
  AND U3769 ( .A(n6585), .B(n6584), .Z(n6602) );
  NAND U3770 ( .A(y[8]), .B(x[6]), .Z(n6931) );
  NANDN U3771 ( .A(n6931), .B(n6586), .Z(n6590) );
  NAND U3772 ( .A(n6588), .B(n6587), .Z(n6589) );
  AND U3773 ( .A(n6590), .B(n6589), .Z(n6606) );
  AND U3774 ( .A(y[9]), .B(x[1]), .Z(n6592) );
  NAND U3775 ( .A(y[7]), .B(x[3]), .Z(n6591) );
  XNOR U3776 ( .A(n6592), .B(n6591), .Z(n6629) );
  NAND U3777 ( .A(y[8]), .B(x[2]), .Z(n6630) );
  XNOR U3778 ( .A(n6606), .B(n6605), .Z(n6608) );
  AND U3779 ( .A(x[10]), .B(y[0]), .Z(n6594) );
  NAND U3780 ( .A(x[0]), .B(y[10]), .Z(n6593) );
  XNOR U3781 ( .A(n6594), .B(n6593), .Z(n6618) );
  ANDN U3782 ( .B(o[9]), .A(n6595), .Z(n6617) );
  XOR U3783 ( .A(n6618), .B(n6617), .Z(n6607) );
  XNOR U3784 ( .A(n6608), .B(n6607), .Z(n6601) );
  NAND U3785 ( .A(n6602), .B(n6601), .Z(n6604) );
  NAND U3786 ( .A(y[1]), .B(x[9]), .Z(n6619) );
  XNOR U3787 ( .A(o[10]), .B(n6619), .Z(n6633) );
  NAND U3788 ( .A(y[2]), .B(x[8]), .Z(n6634) );
  XNOR U3789 ( .A(n6633), .B(n6634), .Z(n6636) );
  XOR U3790 ( .A(n6636), .B(n6635), .Z(n6623) );
  AND U3791 ( .A(y[3]), .B(x[7]), .Z(n6611) );
  NAND U3792 ( .A(x[4]), .B(y[6]), .Z(n6612) );
  XNOR U3793 ( .A(n6611), .B(n6612), .Z(n6614) );
  AND U3794 ( .A(x[6]), .B(y[4]), .Z(n6613) );
  XNOR U3795 ( .A(n6614), .B(n6613), .Z(n6622) );
  XNOR U3796 ( .A(n6623), .B(n6622), .Z(n6624) );
  NAND U3797 ( .A(y[4]), .B(x[7]), .Z(n6683) );
  NANDN U3798 ( .A(n6683), .B(n6596), .Z(n6600) );
  NAND U3799 ( .A(n6598), .B(n6597), .Z(n6599) );
  NAND U3800 ( .A(n6600), .B(n6599), .Z(n6625) );
  XOR U3801 ( .A(n6624), .B(n6625), .Z(n6656) );
  XOR U3802 ( .A(n6602), .B(n6601), .Z(n6657) );
  NANDN U3803 ( .A(n6656), .B(n6657), .Z(n6603) );
  AND U3804 ( .A(n6604), .B(n6603), .Z(n6720) );
  NANDN U3805 ( .A(n6606), .B(n6605), .Z(n6610) );
  NAND U3806 ( .A(n6608), .B(n6607), .Z(n6609) );
  AND U3807 ( .A(n6610), .B(n6609), .Z(n6710) );
  NANDN U3808 ( .A(n6612), .B(n6611), .Z(n6616) );
  NAND U3809 ( .A(n6614), .B(n6613), .Z(n6615) );
  AND U3810 ( .A(n6616), .B(n6615), .Z(n6708) );
  NAND U3811 ( .A(y[10]), .B(x[10]), .Z(n7495) );
  ANDN U3812 ( .B(o[10]), .A(n6619), .Z(n6678) );
  AND U3813 ( .A(x[11]), .B(y[0]), .Z(n6621) );
  NAND U3814 ( .A(y[11]), .B(x[0]), .Z(n6620) );
  XOR U3815 ( .A(n6621), .B(n6620), .Z(n6679) );
  XNOR U3816 ( .A(n6678), .B(n6679), .Z(n6714) );
  AND U3817 ( .A(x[1]), .B(y[10]), .Z(n6695) );
  NAND U3818 ( .A(y[5]), .B(x[6]), .Z(n6696) );
  XNOR U3819 ( .A(n6695), .B(n6696), .Z(n6698) );
  NAND U3820 ( .A(y[1]), .B(x[10]), .Z(n6688) );
  XOR U3821 ( .A(n6698), .B(n6697), .Z(n6713) );
  XOR U3822 ( .A(n6714), .B(n6713), .Z(n6716) );
  XOR U3823 ( .A(n6715), .B(n6716), .Z(n6707) );
  XNOR U3824 ( .A(n6708), .B(n6707), .Z(n6709) );
  XOR U3825 ( .A(n6710), .B(n6709), .Z(n6668) );
  NANDN U3826 ( .A(n6623), .B(n6622), .Z(n6627) );
  NANDN U3827 ( .A(n6625), .B(n6624), .Z(n6626) );
  NAND U3828 ( .A(n6627), .B(n6626), .Z(n6667) );
  AND U3829 ( .A(y[2]), .B(x[9]), .Z(n6682) );
  NAND U3830 ( .A(y[3]), .B(x[8]), .Z(n6685) );
  XNOR U3831 ( .A(n6684), .B(n6685), .Z(n6703) );
  NAND U3832 ( .A(x[3]), .B(y[8]), .Z(n6701) );
  AND U3833 ( .A(x[2]), .B(y[9]), .Z(n6689) );
  NAND U3834 ( .A(x[5]), .B(y[6]), .Z(n6690) );
  XNOR U3835 ( .A(n6689), .B(n6690), .Z(n6691) );
  NAND U3836 ( .A(y[7]), .B(x[4]), .Z(n6692) );
  XNOR U3837 ( .A(n6691), .B(n6692), .Z(n6702) );
  XOR U3838 ( .A(n6701), .B(n6702), .Z(n6704) );
  XOR U3839 ( .A(n6703), .B(n6704), .Z(n6674) );
  AND U3840 ( .A(x[3]), .B(y[9]), .Z(n6757) );
  NANDN U3841 ( .A(n6628), .B(n6757), .Z(n6632) );
  NANDN U3842 ( .A(n6630), .B(n6629), .Z(n6631) );
  AND U3843 ( .A(n6632), .B(n6631), .Z(n6673) );
  NANDN U3844 ( .A(n6634), .B(n6633), .Z(n6638) );
  NAND U3845 ( .A(n6636), .B(n6635), .Z(n6637) );
  NAND U3846 ( .A(n6638), .B(n6637), .Z(n6672) );
  XOR U3847 ( .A(n6673), .B(n6672), .Z(n6675) );
  XNOR U3848 ( .A(n6674), .B(n6675), .Z(n6666) );
  XOR U3849 ( .A(n6667), .B(n6666), .Z(n6669) );
  XOR U3850 ( .A(n6668), .B(n6669), .Z(n6719) );
  XNOR U3851 ( .A(n6720), .B(n6719), .Z(n6721) );
  XNOR U3852 ( .A(n6722), .B(n6721), .Z(n6728) );
  IV U3853 ( .A(n6649), .Z(n8910) );
  NANDN U3854 ( .A(n6644), .B(n6643), .Z(n6648) );
  NAND U3855 ( .A(n6646), .B(n6645), .Z(n6647) );
  NAND U3856 ( .A(n6648), .B(n6647), .Z(n8911) );
  NAND U3857 ( .A(n6651), .B(n6650), .Z(n6655) );
  NANDN U3858 ( .A(n6653), .B(n6652), .Z(n6654) );
  AND U3859 ( .A(n6655), .B(n6654), .Z(n6663) );
  XNOR U3860 ( .A(n6657), .B(n6656), .Z(n6661) );
  XOR U3861 ( .A(n6659), .B(n6658), .Z(n6660) );
  XOR U3862 ( .A(n6661), .B(n6660), .Z(n6662) );
  XNOR U3863 ( .A(n6663), .B(n6662), .Z(n8913) );
  NAND U3864 ( .A(n6661), .B(n6660), .Z(n6665) );
  NAND U3865 ( .A(n6663), .B(n6662), .Z(n6664) );
  NAND U3866 ( .A(n6665), .B(n6664), .Z(n6725) );
  XNOR U3867 ( .A(n6726), .B(n6725), .Z(n6727) );
  XNOR U3868 ( .A(n6728), .B(n6727), .Z(N44) );
  NAND U3869 ( .A(n6667), .B(n6666), .Z(n6671) );
  NAND U3870 ( .A(n6669), .B(n6668), .Z(n6670) );
  NAND U3871 ( .A(n6671), .B(n6670), .Z(n6803) );
  NANDN U3872 ( .A(n6673), .B(n6672), .Z(n6677) );
  OR U3873 ( .A(n6675), .B(n6674), .Z(n6676) );
  AND U3874 ( .A(n6677), .B(n6676), .Z(n6792) );
  NAND U3875 ( .A(x[11]), .B(y[11]), .Z(n7771) );
  NANDN U3876 ( .A(n7771), .B(n7024), .Z(n6681) );
  NANDN U3877 ( .A(n6679), .B(n6678), .Z(n6680) );
  AND U3878 ( .A(n6681), .B(n6680), .Z(n6769) );
  NANDN U3879 ( .A(n6683), .B(n6682), .Z(n6687) );
  NANDN U3880 ( .A(n6685), .B(n6684), .Z(n6686) );
  AND U3881 ( .A(n6687), .B(n6686), .Z(n6767) );
  ANDN U3882 ( .B(o[11]), .A(n6688), .Z(n6781) );
  NAND U3883 ( .A(x[1]), .B(y[11]), .Z(n6778) );
  XNOR U3884 ( .A(n6778), .B(n6779), .Z(n6780) );
  XOR U3885 ( .A(n6781), .B(n6780), .Z(n6766) );
  XNOR U3886 ( .A(n6767), .B(n6766), .Z(n6768) );
  XNOR U3887 ( .A(n6769), .B(n6768), .Z(n6790) );
  AND U3888 ( .A(x[2]), .B(y[10]), .Z(n6755) );
  NAND U3889 ( .A(y[4]), .B(x[8]), .Z(n6756) );
  XOR U3890 ( .A(n6758), .B(n6757), .Z(n6744) );
  NAND U3891 ( .A(y[1]), .B(x[11]), .Z(n6763) );
  AND U3892 ( .A(y[12]), .B(x[0]), .Z(n6772) );
  NAND U3893 ( .A(y[0]), .B(x[12]), .Z(n6773) );
  XNOR U3894 ( .A(n6775), .B(n6774), .Z(n6743) );
  XNOR U3895 ( .A(n6744), .B(n6743), .Z(n6746) );
  AND U3896 ( .A(y[8]), .B(x[4]), .Z(n6785) );
  AND U3897 ( .A(y[2]), .B(x[10]), .Z(n6784) );
  XOR U3898 ( .A(n6785), .B(n6784), .Z(n6787) );
  AND U3899 ( .A(y[3]), .B(x[9]), .Z(n6786) );
  XOR U3900 ( .A(n6787), .B(n6786), .Z(n6752) );
  NAND U3901 ( .A(y[5]), .B(x[7]), .Z(n6750) );
  NAND U3902 ( .A(x[5]), .B(y[7]), .Z(n6749) );
  XOR U3903 ( .A(n6750), .B(n6749), .Z(n6751) );
  XOR U3904 ( .A(n6746), .B(n6745), .Z(n6740) );
  NANDN U3905 ( .A(n6690), .B(n6689), .Z(n6694) );
  NANDN U3906 ( .A(n6692), .B(n6691), .Z(n6693) );
  AND U3907 ( .A(n6694), .B(n6693), .Z(n6738) );
  NANDN U3908 ( .A(n6696), .B(n6695), .Z(n6700) );
  NAND U3909 ( .A(n6698), .B(n6697), .Z(n6699) );
  NAND U3910 ( .A(n6700), .B(n6699), .Z(n6737) );
  XNOR U3911 ( .A(n6738), .B(n6737), .Z(n6739) );
  XOR U3912 ( .A(n6740), .B(n6739), .Z(n6791) );
  XOR U3913 ( .A(n6790), .B(n6791), .Z(n6793) );
  XNOR U3914 ( .A(n6792), .B(n6793), .Z(n6802) );
  XOR U3915 ( .A(n6803), .B(n6802), .Z(n6805) );
  NANDN U3916 ( .A(n6702), .B(n6701), .Z(n6706) );
  OR U3917 ( .A(n6704), .B(n6703), .Z(n6705) );
  AND U3918 ( .A(n6706), .B(n6705), .Z(n6732) );
  NANDN U3919 ( .A(n6708), .B(n6707), .Z(n6712) );
  NANDN U3920 ( .A(n6710), .B(n6709), .Z(n6711) );
  AND U3921 ( .A(n6712), .B(n6711), .Z(n6731) );
  XNOR U3922 ( .A(n6732), .B(n6731), .Z(n6733) );
  NAND U3923 ( .A(n6714), .B(n6713), .Z(n6718) );
  NAND U3924 ( .A(n6716), .B(n6715), .Z(n6717) );
  NAND U3925 ( .A(n6718), .B(n6717), .Z(n6734) );
  XNOR U3926 ( .A(n6733), .B(n6734), .Z(n6804) );
  XOR U3927 ( .A(n6805), .B(n6804), .Z(n6797) );
  NANDN U3928 ( .A(n6720), .B(n6719), .Z(n6724) );
  NANDN U3929 ( .A(n6722), .B(n6721), .Z(n6723) );
  AND U3930 ( .A(n6724), .B(n6723), .Z(n6796) );
  XNOR U3931 ( .A(n6797), .B(n6796), .Z(n6799) );
  NANDN U3932 ( .A(n6726), .B(n6725), .Z(n6730) );
  NAND U3933 ( .A(n6728), .B(n6727), .Z(n6729) );
  AND U3934 ( .A(n6730), .B(n6729), .Z(n6798) );
  XOR U3935 ( .A(n6799), .B(n6798), .Z(N45) );
  NANDN U3936 ( .A(n6732), .B(n6731), .Z(n6736) );
  NANDN U3937 ( .A(n6734), .B(n6733), .Z(n6735) );
  AND U3938 ( .A(n6736), .B(n6735), .Z(n6877) );
  NANDN U3939 ( .A(n6738), .B(n6737), .Z(n6742) );
  NANDN U3940 ( .A(n6740), .B(n6739), .Z(n6741) );
  AND U3941 ( .A(n6742), .B(n6741), .Z(n6863) );
  NANDN U3942 ( .A(n6744), .B(n6743), .Z(n6748) );
  NAND U3943 ( .A(n6746), .B(n6745), .Z(n6747) );
  AND U3944 ( .A(n6748), .B(n6747), .Z(n6869) );
  NAND U3945 ( .A(n6750), .B(n6749), .Z(n6754) );
  NANDN U3946 ( .A(n6752), .B(n6751), .Z(n6753) );
  AND U3947 ( .A(n6754), .B(n6753), .Z(n6868) );
  XOR U3948 ( .A(n6869), .B(n6868), .Z(n6870) );
  NANDN U3949 ( .A(n6756), .B(n6755), .Z(n6760) );
  NAND U3950 ( .A(n6758), .B(n6757), .Z(n6759) );
  AND U3951 ( .A(n6760), .B(n6759), .Z(n6846) );
  AND U3952 ( .A(y[6]), .B(x[7]), .Z(n6762) );
  NAND U3953 ( .A(y[12]), .B(x[1]), .Z(n6761) );
  XNOR U3954 ( .A(n6762), .B(n6761), .Z(n6851) );
  ANDN U3955 ( .B(o[12]), .A(n6763), .Z(n6850) );
  XOR U3956 ( .A(n6851), .B(n6850), .Z(n6844) );
  AND U3957 ( .A(x[9]), .B(y[4]), .Z(n6765) );
  NAND U3958 ( .A(y[11]), .B(x[2]), .Z(n6764) );
  XNOR U3959 ( .A(n6765), .B(n6764), .Z(n6832) );
  NAND U3960 ( .A(y[7]), .B(x[6]), .Z(n6833) );
  XOR U3961 ( .A(n6844), .B(n6843), .Z(n6845) );
  XNOR U3962 ( .A(n6870), .B(n6871), .Z(n6862) );
  XNOR U3963 ( .A(n6863), .B(n6862), .Z(n6865) );
  NANDN U3964 ( .A(n6767), .B(n6766), .Z(n6771) );
  NANDN U3965 ( .A(n6769), .B(n6768), .Z(n6770) );
  NAND U3966 ( .A(n6771), .B(n6770), .Z(n6810) );
  NANDN U3967 ( .A(n6773), .B(n6772), .Z(n6777) );
  NAND U3968 ( .A(n6775), .B(n6774), .Z(n6776) );
  AND U3969 ( .A(n6777), .B(n6776), .Z(n6838) );
  AND U3970 ( .A(y[3]), .B(x[10]), .Z(n6857) );
  AND U3971 ( .A(y[2]), .B(x[11]), .Z(n6855) );
  NAND U3972 ( .A(y[5]), .B(x[8]), .Z(n6854) );
  XOR U3973 ( .A(n6857), .B(n6856), .Z(n6837) );
  NANDN U3974 ( .A(n6779), .B(n6778), .Z(n6783) );
  NANDN U3975 ( .A(n6781), .B(n6780), .Z(n6782) );
  NAND U3976 ( .A(n6783), .B(n6782), .Z(n6840) );
  NAND U3977 ( .A(n6785), .B(n6784), .Z(n6789) );
  NAND U3978 ( .A(n6787), .B(n6786), .Z(n6788) );
  NAND U3979 ( .A(n6789), .B(n6788), .Z(n6816) );
  NAND U3980 ( .A(y[1]), .B(x[12]), .Z(n6836) );
  AND U3981 ( .A(x[0]), .B(y[13]), .Z(n6826) );
  NAND U3982 ( .A(x[13]), .B(y[0]), .Z(n6827) );
  XOR U3983 ( .A(n6829), .B(n6828), .Z(n6815) );
  AND U3984 ( .A(x[5]), .B(y[8]), .Z(n6820) );
  NAND U3985 ( .A(x[3]), .B(y[10]), .Z(n6821) );
  NAND U3986 ( .A(x[4]), .B(y[9]), .Z(n6823) );
  XOR U3987 ( .A(n6815), .B(n6814), .Z(n6817) );
  XNOR U3988 ( .A(n6816), .B(n6817), .Z(n6809) );
  XOR U3989 ( .A(n6810), .B(n6811), .Z(n6864) );
  XOR U3990 ( .A(n6865), .B(n6864), .Z(n6875) );
  NANDN U3991 ( .A(n6791), .B(n6790), .Z(n6795) );
  OR U3992 ( .A(n6793), .B(n6792), .Z(n6794) );
  AND U3993 ( .A(n6795), .B(n6794), .Z(n6874) );
  NANDN U3994 ( .A(n6797), .B(n6796), .Z(n6801) );
  NAND U3995 ( .A(n6799), .B(n6798), .Z(n6800) );
  NAND U3996 ( .A(n6801), .B(n6800), .Z(n6880) );
  XOR U3997 ( .A(n6881), .B(n6880), .Z(n6883) );
  NAND U3998 ( .A(n6803), .B(n6802), .Z(n6807) );
  NAND U3999 ( .A(n6805), .B(n6804), .Z(n6806) );
  AND U4000 ( .A(n6807), .B(n6806), .Z(n6882) );
  XOR U4001 ( .A(n6883), .B(n6882), .Z(N46) );
  NANDN U4002 ( .A(n6809), .B(n6808), .Z(n6813) );
  NAND U4003 ( .A(n6811), .B(n6810), .Z(n6812) );
  NAND U4004 ( .A(n6813), .B(n6812), .Z(n6889) );
  NAND U4005 ( .A(n6815), .B(n6814), .Z(n6819) );
  NAND U4006 ( .A(n6817), .B(n6816), .Z(n6818) );
  AND U4007 ( .A(n6819), .B(n6818), .Z(n6956) );
  NANDN U4008 ( .A(n6821), .B(n6820), .Z(n6825) );
  NANDN U4009 ( .A(n6823), .B(n6822), .Z(n6824) );
  AND U4010 ( .A(n6825), .B(n6824), .Z(n6939) );
  NANDN U4011 ( .A(n6827), .B(n6826), .Z(n6831) );
  NAND U4012 ( .A(n6829), .B(n6828), .Z(n6830) );
  AND U4013 ( .A(n6831), .B(n6830), .Z(n6937) );
  AND U4014 ( .A(y[3]), .B(x[11]), .Z(n6930) );
  NAND U4015 ( .A(x[1]), .B(y[13]), .Z(n6933) );
  AND U4016 ( .A(x[9]), .B(y[11]), .Z(n7542) );
  NAND U4017 ( .A(n7542), .B(n6925), .Z(n6835) );
  NANDN U4018 ( .A(n6833), .B(n6832), .Z(n6834) );
  NAND U4019 ( .A(n6835), .B(n6834), .Z(n6945) );
  ANDN U4020 ( .B(o[13]), .A(n6836), .Z(n6914) );
  AND U4021 ( .A(y[14]), .B(x[0]), .Z(n6911) );
  NAND U4022 ( .A(x[14]), .B(y[0]), .Z(n6912) );
  XOR U4023 ( .A(n6914), .B(n6913), .Z(n6943) );
  NAND U4024 ( .A(x[13]), .B(y[1]), .Z(n6922) );
  XNOR U4025 ( .A(o[14]), .B(n6922), .Z(n6919) );
  AND U4026 ( .A(y[2]), .B(x[12]), .Z(n7186) );
  AND U4027 ( .A(y[7]), .B(x[7]), .Z(n6917) );
  XOR U4028 ( .A(n7186), .B(n6917), .Z(n6918) );
  XOR U4029 ( .A(n6919), .B(n6918), .Z(n6942) );
  XOR U4030 ( .A(n6943), .B(n6942), .Z(n6944) );
  XNOR U4031 ( .A(n6945), .B(n6944), .Z(n6954) );
  XOR U4032 ( .A(n6956), .B(n6957), .Z(n6887) );
  NANDN U4033 ( .A(n6838), .B(n6837), .Z(n6842) );
  NANDN U4034 ( .A(n6840), .B(n6839), .Z(n6841) );
  AND U4035 ( .A(n6842), .B(n6841), .Z(n6951) );
  NAND U4036 ( .A(n6844), .B(n6843), .Z(n6848) );
  NANDN U4037 ( .A(n6846), .B(n6845), .Z(n6847) );
  AND U4038 ( .A(n6848), .B(n6847), .Z(n6949) );
  NAND U4039 ( .A(y[12]), .B(x[7]), .Z(n7436) );
  NANDN U4040 ( .A(n7436), .B(n6849), .Z(n6853) );
  NAND U4041 ( .A(n6851), .B(n6850), .Z(n6852) );
  AND U4042 ( .A(n6853), .B(n6852), .Z(n6894) );
  NANDN U4043 ( .A(n6855), .B(n6854), .Z(n6859) );
  NANDN U4044 ( .A(n6857), .B(n6856), .Z(n6858) );
  AND U4045 ( .A(n6859), .B(n6858), .Z(n6893) );
  AND U4046 ( .A(x[10]), .B(y[4]), .Z(n6861) );
  NAND U4047 ( .A(y[12]), .B(x[2]), .Z(n6860) );
  XNOR U4048 ( .A(n6861), .B(n6860), .Z(n6927) );
  AND U4049 ( .A(y[5]), .B(x[9]), .Z(n6926) );
  XOR U4050 ( .A(n6927), .B(n6926), .Z(n6902) );
  AND U4051 ( .A(x[3]), .B(y[11]), .Z(n6905) );
  NAND U4052 ( .A(y[6]), .B(x[8]), .Z(n6906) );
  NAND U4053 ( .A(x[5]), .B(y[9]), .Z(n6908) );
  AND U4054 ( .A(y[10]), .B(x[4]), .Z(n6899) );
  XOR U4055 ( .A(n6900), .B(n6899), .Z(n6901) );
  XOR U4056 ( .A(n6902), .B(n6901), .Z(n6895) );
  XOR U4057 ( .A(n6896), .B(n6895), .Z(n6948) );
  XOR U4058 ( .A(n6887), .B(n6888), .Z(n6890) );
  XOR U4059 ( .A(n6889), .B(n6890), .Z(n6966) );
  NANDN U4060 ( .A(n6863), .B(n6862), .Z(n6867) );
  NAND U4061 ( .A(n6865), .B(n6864), .Z(n6866) );
  AND U4062 ( .A(n6867), .B(n6866), .Z(n6964) );
  NAND U4063 ( .A(n6869), .B(n6868), .Z(n6873) );
  NANDN U4064 ( .A(n6871), .B(n6870), .Z(n6872) );
  NAND U4065 ( .A(n6873), .B(n6872), .Z(n6965) );
  XNOR U4066 ( .A(n6964), .B(n6965), .Z(n6967) );
  XNOR U4067 ( .A(n6966), .B(n6967), .Z(n6963) );
  NANDN U4068 ( .A(n6875), .B(n6874), .Z(n6879) );
  NANDN U4069 ( .A(n6877), .B(n6876), .Z(n6878) );
  NAND U4070 ( .A(n6879), .B(n6878), .Z(n6961) );
  NAND U4071 ( .A(n6881), .B(n6880), .Z(n6885) );
  NAND U4072 ( .A(n6883), .B(n6882), .Z(n6884) );
  AND U4073 ( .A(n6885), .B(n6884), .Z(n6962) );
  IV U4074 ( .A(n6962), .Z(n6960) );
  XOR U4075 ( .A(n6961), .B(n6960), .Z(n6886) );
  XNOR U4076 ( .A(n6963), .B(n6886), .Z(N47) );
  NANDN U4077 ( .A(n6888), .B(n6887), .Z(n6892) );
  NANDN U4078 ( .A(n6890), .B(n6889), .Z(n6891) );
  NAND U4079 ( .A(n6892), .B(n6891), .Z(n6973) );
  NANDN U4080 ( .A(n6894), .B(n6893), .Z(n6898) );
  NAND U4081 ( .A(n6896), .B(n6895), .Z(n6897) );
  NAND U4082 ( .A(n6898), .B(n6897), .Z(n6988) );
  NAND U4083 ( .A(n6900), .B(n6899), .Z(n6904) );
  NAND U4084 ( .A(n6902), .B(n6901), .Z(n6903) );
  NAND U4085 ( .A(n6904), .B(n6903), .Z(n6986) );
  NANDN U4086 ( .A(n6906), .B(n6905), .Z(n6910) );
  NANDN U4087 ( .A(n6908), .B(n6907), .Z(n6909) );
  AND U4088 ( .A(n6910), .B(n6909), .Z(n7019) );
  NANDN U4089 ( .A(n6912), .B(n6911), .Z(n6916) );
  NAND U4090 ( .A(n6914), .B(n6913), .Z(n6915) );
  NAND U4091 ( .A(n6916), .B(n6915), .Z(n7018) );
  AND U4092 ( .A(x[4]), .B(y[11]), .Z(n7035) );
  NAND U4093 ( .A(y[5]), .B(x[10]), .Z(n7036) );
  XNOR U4094 ( .A(n7035), .B(n7036), .Z(n7037) );
  NAND U4095 ( .A(y[8]), .B(x[7]), .Z(n7038) );
  XNOR U4096 ( .A(n7037), .B(n7038), .Z(n7048) );
  NAND U4097 ( .A(x[6]), .B(y[9]), .Z(n7049) );
  NAND U4098 ( .A(x[5]), .B(y[10]), .Z(n7051) );
  AND U4099 ( .A(x[2]), .B(y[13]), .Z(n7041) );
  NAND U4100 ( .A(x[9]), .B(y[6]), .Z(n7042) );
  NAND U4101 ( .A(x[3]), .B(y[12]), .Z(n7044) );
  AND U4102 ( .A(x[1]), .B(y[14]), .Z(n7029) );
  NAND U4103 ( .A(y[7]), .B(x[8]), .Z(n7030) );
  XNOR U4104 ( .A(n7029), .B(n7030), .Z(n7031) );
  NAND U4105 ( .A(x[14]), .B(y[1]), .Z(n7047) );
  XOR U4106 ( .A(o[15]), .B(n7047), .Z(n7032) );
  XOR U4107 ( .A(n7031), .B(n7032), .Z(n6999) );
  XOR U4108 ( .A(n7001), .B(n7000), .Z(n7020) );
  XOR U4109 ( .A(n7021), .B(n7020), .Z(n6987) );
  XNOR U4110 ( .A(n6986), .B(n6987), .Z(n6989) );
  NAND U4111 ( .A(n7186), .B(n6917), .Z(n6921) );
  AND U4112 ( .A(n6919), .B(n6918), .Z(n6920) );
  ANDN U4113 ( .B(n6921), .A(n6920), .Z(n7007) );
  ANDN U4114 ( .B(o[14]), .A(n6922), .Z(n7025) );
  AND U4115 ( .A(x[15]), .B(y[0]), .Z(n6924) );
  NAND U4116 ( .A(x[0]), .B(y[15]), .Z(n6923) );
  XOR U4117 ( .A(n6924), .B(n6923), .Z(n7026) );
  XNOR U4118 ( .A(n7025), .B(n7026), .Z(n7004) );
  AND U4119 ( .A(y[4]), .B(x[11]), .Z(n7010) );
  NAND U4120 ( .A(x[13]), .B(y[2]), .Z(n7011) );
  XNOR U4121 ( .A(n7010), .B(n7011), .Z(n7012) );
  NAND U4122 ( .A(y[3]), .B(x[12]), .Z(n7013) );
  XOR U4123 ( .A(n7012), .B(n7013), .Z(n7005) );
  NAND U4124 ( .A(y[12]), .B(x[10]), .Z(n7755) );
  NANDN U4125 ( .A(n7755), .B(n6925), .Z(n6929) );
  NAND U4126 ( .A(n6927), .B(n6926), .Z(n6928) );
  NAND U4127 ( .A(n6929), .B(n6928), .Z(n6992) );
  XOR U4128 ( .A(n6993), .B(n6992), .Z(n6995) );
  NANDN U4129 ( .A(n6931), .B(n6930), .Z(n6935) );
  NANDN U4130 ( .A(n6933), .B(n6932), .Z(n6934) );
  NAND U4131 ( .A(n6935), .B(n6934), .Z(n6994) );
  XOR U4132 ( .A(n6995), .B(n6994), .Z(n6983) );
  NANDN U4133 ( .A(n6937), .B(n6936), .Z(n6941) );
  NANDN U4134 ( .A(n6939), .B(n6938), .Z(n6940) );
  NAND U4135 ( .A(n6941), .B(n6940), .Z(n6981) );
  NAND U4136 ( .A(n6943), .B(n6942), .Z(n6947) );
  NAND U4137 ( .A(n6945), .B(n6944), .Z(n6946) );
  NAND U4138 ( .A(n6947), .B(n6946), .Z(n6980) );
  XOR U4139 ( .A(n6981), .B(n6980), .Z(n6982) );
  XNOR U4140 ( .A(n6983), .B(n6982), .Z(n7054) );
  XOR U4141 ( .A(n7055), .B(n7054), .Z(n7056) );
  NANDN U4142 ( .A(n6949), .B(n6948), .Z(n6953) );
  NANDN U4143 ( .A(n6951), .B(n6950), .Z(n6952) );
  NAND U4144 ( .A(n6953), .B(n6952), .Z(n7057) );
  NANDN U4145 ( .A(n6955), .B(n6954), .Z(n6959) );
  NANDN U4146 ( .A(n6957), .B(n6956), .Z(n6958) );
  AND U4147 ( .A(n6959), .B(n6958), .Z(n6971) );
  XOR U4148 ( .A(n6973), .B(n6974), .Z(n6979) );
  NANDN U4149 ( .A(n6965), .B(n6964), .Z(n6969) );
  NAND U4150 ( .A(n6967), .B(n6966), .Z(n6968) );
  AND U4151 ( .A(n6969), .B(n6968), .Z(n6978) );
  XOR U4152 ( .A(n6977), .B(n6978), .Z(n6970) );
  XNOR U4153 ( .A(n6979), .B(n6970), .Z(N48) );
  NANDN U4154 ( .A(n6972), .B(n6971), .Z(n6976) );
  NANDN U4155 ( .A(n6974), .B(n6973), .Z(n6975) );
  AND U4156 ( .A(n6976), .B(n6975), .Z(n7148) );
  NAND U4157 ( .A(n6981), .B(n6980), .Z(n6985) );
  NAND U4158 ( .A(n6983), .B(n6982), .Z(n6984) );
  NAND U4159 ( .A(n6985), .B(n6984), .Z(n7063) );
  NAND U4160 ( .A(n6987), .B(n6986), .Z(n6991) );
  NANDN U4161 ( .A(n6989), .B(n6988), .Z(n6990) );
  NAND U4162 ( .A(n6991), .B(n6990), .Z(n7062) );
  NAND U4163 ( .A(n6993), .B(n6992), .Z(n6997) );
  NAND U4164 ( .A(n6995), .B(n6994), .Z(n6996) );
  NAND U4165 ( .A(n6997), .B(n6996), .Z(n7061) );
  XOR U4166 ( .A(n7062), .B(n7061), .Z(n7064) );
  XOR U4167 ( .A(n7063), .B(n7064), .Z(n7155) );
  NANDN U4168 ( .A(n6999), .B(n6998), .Z(n7003) );
  NAND U4169 ( .A(n7001), .B(n7000), .Z(n7002) );
  AND U4170 ( .A(n7003), .B(n7002), .Z(n7142) );
  NANDN U4171 ( .A(n7005), .B(n7004), .Z(n7009) );
  NANDN U4172 ( .A(n7007), .B(n7006), .Z(n7008) );
  AND U4173 ( .A(n7009), .B(n7008), .Z(n7140) );
  NANDN U4174 ( .A(n7011), .B(n7010), .Z(n7015) );
  NANDN U4175 ( .A(n7013), .B(n7012), .Z(n7014) );
  AND U4176 ( .A(n7015), .B(n7014), .Z(n7124) );
  AND U4177 ( .A(y[11]), .B(x[5]), .Z(n7017) );
  NAND U4178 ( .A(y[3]), .B(x[13]), .Z(n7016) );
  XNOR U4179 ( .A(n7017), .B(n7016), .Z(n7096) );
  NAND U4180 ( .A(y[4]), .B(x[12]), .Z(n7097) );
  XNOR U4181 ( .A(n7096), .B(n7097), .Z(n7121) );
  AND U4182 ( .A(y[7]), .B(x[9]), .Z(n7127) );
  NAND U4183 ( .A(y[14]), .B(x[2]), .Z(n7128) );
  XNOR U4184 ( .A(n7127), .B(n7128), .Z(n7129) );
  NAND U4185 ( .A(x[3]), .B(y[13]), .Z(n7130) );
  XOR U4186 ( .A(n7129), .B(n7130), .Z(n7122) );
  XNOR U4187 ( .A(n7121), .B(n7122), .Z(n7123) );
  XNOR U4188 ( .A(n7124), .B(n7123), .Z(n7139) );
  NANDN U4189 ( .A(n7019), .B(n7018), .Z(n7023) );
  NAND U4190 ( .A(n7021), .B(n7020), .Z(n7022) );
  AND U4191 ( .A(n7023), .B(n7022), .Z(n7110) );
  AND U4192 ( .A(y[15]), .B(x[15]), .Z(n9052) );
  NAND U4193 ( .A(n9052), .B(n7024), .Z(n7028) );
  NANDN U4194 ( .A(n7026), .B(n7025), .Z(n7027) );
  AND U4195 ( .A(n7028), .B(n7027), .Z(n7116) );
  NANDN U4196 ( .A(n7030), .B(n7029), .Z(n7034) );
  NANDN U4197 ( .A(n7032), .B(n7031), .Z(n7033) );
  NAND U4198 ( .A(n7034), .B(n7033), .Z(n7115) );
  XNOR U4199 ( .A(n7116), .B(n7115), .Z(n7118) );
  NANDN U4200 ( .A(n7036), .B(n7035), .Z(n7040) );
  NANDN U4201 ( .A(n7038), .B(n7037), .Z(n7039) );
  AND U4202 ( .A(n7040), .B(n7039), .Z(n7106) );
  AND U4203 ( .A(x[16]), .B(y[0]), .Z(n7079) );
  NAND U4204 ( .A(x[0]), .B(y[16]), .Z(n7080) );
  XNOR U4205 ( .A(n7079), .B(n7080), .Z(n7081) );
  NAND U4206 ( .A(y[1]), .B(x[15]), .Z(n7100) );
  XOR U4207 ( .A(o[16]), .B(n7100), .Z(n7082) );
  XNOR U4208 ( .A(n7081), .B(n7082), .Z(n7103) );
  AND U4209 ( .A(x[7]), .B(y[9]), .Z(n7089) );
  NAND U4210 ( .A(x[6]), .B(y[10]), .Z(n7090) );
  XNOR U4211 ( .A(n7089), .B(n7090), .Z(n7091) );
  NAND U4212 ( .A(y[6]), .B(x[10]), .Z(n7092) );
  XOR U4213 ( .A(n7091), .B(n7092), .Z(n7104) );
  XNOR U4214 ( .A(n7103), .B(n7104), .Z(n7105) );
  XNOR U4215 ( .A(n7106), .B(n7105), .Z(n7117) );
  XOR U4216 ( .A(n7118), .B(n7117), .Z(n7070) );
  NANDN U4217 ( .A(n7042), .B(n7041), .Z(n7046) );
  NANDN U4218 ( .A(n7044), .B(n7043), .Z(n7045) );
  AND U4219 ( .A(n7046), .B(n7045), .Z(n7076) );
  AND U4220 ( .A(y[2]), .B(x[14]), .Z(n7133) );
  NAND U4221 ( .A(y[5]), .B(x[11]), .Z(n7134) );
  XNOR U4222 ( .A(n7133), .B(n7134), .Z(n7135) );
  NAND U4223 ( .A(y[12]), .B(x[4]), .Z(n7136) );
  XNOR U4224 ( .A(n7135), .B(n7136), .Z(n7074) );
  AND U4225 ( .A(y[15]), .B(x[1]), .Z(n7085) );
  ANDN U4226 ( .B(o[15]), .A(n7047), .Z(n7087) );
  XOR U4227 ( .A(n7088), .B(n7087), .Z(n7073) );
  XOR U4228 ( .A(n7074), .B(n7073), .Z(n7075) );
  NANDN U4229 ( .A(n7049), .B(n7048), .Z(n7053) );
  NANDN U4230 ( .A(n7051), .B(n7050), .Z(n7052) );
  AND U4231 ( .A(n7053), .B(n7052), .Z(n7068) );
  XOR U4232 ( .A(n7067), .B(n7068), .Z(n7069) );
  XOR U4233 ( .A(n7110), .B(n7109), .Z(n7112) );
  XNOR U4234 ( .A(n7111), .B(n7112), .Z(n7152) );
  NAND U4235 ( .A(n7055), .B(n7054), .Z(n7059) );
  NANDN U4236 ( .A(n7057), .B(n7056), .Z(n7058) );
  AND U4237 ( .A(n7059), .B(n7058), .Z(n7153) );
  XOR U4238 ( .A(n7152), .B(n7153), .Z(n7154) );
  XOR U4239 ( .A(n7155), .B(n7154), .Z(n7146) );
  IV U4240 ( .A(n7146), .Z(n7145) );
  XOR U4241 ( .A(n7147), .B(n7145), .Z(n7060) );
  XNOR U4242 ( .A(n7148), .B(n7060), .Z(N49) );
  NAND U4243 ( .A(n7062), .B(n7061), .Z(n7066) );
  NAND U4244 ( .A(n7064), .B(n7063), .Z(n7065) );
  NAND U4245 ( .A(n7066), .B(n7065), .Z(n7161) );
  NAND U4246 ( .A(n7068), .B(n7067), .Z(n7072) );
  NANDN U4247 ( .A(n7070), .B(n7069), .Z(n7071) );
  AND U4248 ( .A(n7072), .B(n7071), .Z(n7252) );
  NAND U4249 ( .A(n7074), .B(n7073), .Z(n7078) );
  NANDN U4250 ( .A(n7076), .B(n7075), .Z(n7077) );
  AND U4251 ( .A(n7078), .B(n7077), .Z(n7249) );
  NANDN U4252 ( .A(n7080), .B(n7079), .Z(n7084) );
  NANDN U4253 ( .A(n7082), .B(n7081), .Z(n7083) );
  AND U4254 ( .A(n7084), .B(n7083), .Z(n7200) );
  AND U4255 ( .A(y[7]), .B(x[10]), .Z(n7215) );
  NAND U4256 ( .A(y[15]), .B(x[2]), .Z(n7216) );
  XNOR U4257 ( .A(n7215), .B(n7216), .Z(n7217) );
  NAND U4258 ( .A(x[3]), .B(y[14]), .Z(n7218) );
  XNOR U4259 ( .A(n7217), .B(n7218), .Z(n7197) );
  AND U4260 ( .A(x[0]), .B(y[17]), .Z(n7172) );
  NAND U4261 ( .A(x[17]), .B(y[0]), .Z(n7173) );
  XNOR U4262 ( .A(n7172), .B(n7173), .Z(n7174) );
  NAND U4263 ( .A(x[16]), .B(y[1]), .Z(n7179) );
  XOR U4264 ( .A(o[17]), .B(n7179), .Z(n7175) );
  XOR U4265 ( .A(n7174), .B(n7175), .Z(n7198) );
  XNOR U4266 ( .A(n7197), .B(n7198), .Z(n7199) );
  XNOR U4267 ( .A(n7200), .B(n7199), .Z(n7206) );
  NANDN U4268 ( .A(n7090), .B(n7089), .Z(n7094) );
  NANDN U4269 ( .A(n7092), .B(n7091), .Z(n7093) );
  NAND U4270 ( .A(n7094), .B(n7093), .Z(n7203) );
  XNOR U4271 ( .A(n7204), .B(n7203), .Z(n7205) );
  XOR U4272 ( .A(n7206), .B(n7205), .Z(n7244) );
  AND U4273 ( .A(x[13]), .B(y[11]), .Z(n8028) );
  NANDN U4274 ( .A(n7095), .B(n8028), .Z(n7099) );
  NANDN U4275 ( .A(n7097), .B(n7096), .Z(n7098) );
  AND U4276 ( .A(n7099), .B(n7098), .Z(n7193) );
  AND U4277 ( .A(y[8]), .B(x[9]), .Z(n7221) );
  NAND U4278 ( .A(x[1]), .B(y[16]), .Z(n7222) );
  XNOR U4279 ( .A(n7221), .B(n7222), .Z(n7224) );
  ANDN U4280 ( .B(o[16]), .A(n7100), .Z(n7223) );
  XOR U4281 ( .A(n7224), .B(n7223), .Z(n7191) );
  AND U4282 ( .A(x[15]), .B(y[2]), .Z(n7102) );
  NAND U4283 ( .A(x[12]), .B(y[5]), .Z(n7101) );
  XNOR U4284 ( .A(n7102), .B(n7101), .Z(n7187) );
  NAND U4285 ( .A(x[14]), .B(y[3]), .Z(n7188) );
  XOR U4286 ( .A(n7187), .B(n7188), .Z(n7192) );
  XOR U4287 ( .A(n7191), .B(n7192), .Z(n7194) );
  XNOR U4288 ( .A(n7193), .B(n7194), .Z(n7243) );
  XNOR U4289 ( .A(n7244), .B(n7243), .Z(n7245) );
  NANDN U4290 ( .A(n7104), .B(n7103), .Z(n7108) );
  NANDN U4291 ( .A(n7106), .B(n7105), .Z(n7107) );
  NAND U4292 ( .A(n7108), .B(n7107), .Z(n7246) );
  XOR U4293 ( .A(n7245), .B(n7246), .Z(n7250) );
  NAND U4294 ( .A(n7110), .B(n7109), .Z(n7114) );
  NAND U4295 ( .A(n7112), .B(n7111), .Z(n7113) );
  NAND U4296 ( .A(n7114), .B(n7113), .Z(n7258) );
  NANDN U4297 ( .A(n7116), .B(n7115), .Z(n7120) );
  NAND U4298 ( .A(n7118), .B(n7117), .Z(n7119) );
  AND U4299 ( .A(n7120), .B(n7119), .Z(n7239) );
  NANDN U4300 ( .A(n7122), .B(n7121), .Z(n7126) );
  NANDN U4301 ( .A(n7124), .B(n7123), .Z(n7125) );
  AND U4302 ( .A(n7126), .B(n7125), .Z(n7238) );
  NANDN U4303 ( .A(n7128), .B(n7127), .Z(n7132) );
  NANDN U4304 ( .A(n7130), .B(n7129), .Z(n7131) );
  AND U4305 ( .A(n7132), .B(n7131), .Z(n7210) );
  NANDN U4306 ( .A(n7134), .B(n7133), .Z(n7138) );
  NANDN U4307 ( .A(n7136), .B(n7135), .Z(n7137) );
  NAND U4308 ( .A(n7138), .B(n7137), .Z(n7209) );
  XNOR U4309 ( .A(n7210), .B(n7209), .Z(n7211) );
  AND U4310 ( .A(y[9]), .B(x[8]), .Z(n7225) );
  NAND U4311 ( .A(x[5]), .B(y[12]), .Z(n7226) );
  XNOR U4312 ( .A(n7225), .B(n7226), .Z(n7227) );
  NAND U4313 ( .A(x[6]), .B(y[11]), .Z(n7228) );
  XNOR U4314 ( .A(n7227), .B(n7228), .Z(n7231) );
  NAND U4315 ( .A(x[7]), .B(y[10]), .Z(n7232) );
  XNOR U4316 ( .A(n7231), .B(n7232), .Z(n7233) );
  AND U4317 ( .A(x[4]), .B(y[13]), .Z(n7180) );
  NAND U4318 ( .A(x[13]), .B(y[4]), .Z(n7181) );
  XNOR U4319 ( .A(n7180), .B(n7181), .Z(n7182) );
  NAND U4320 ( .A(y[6]), .B(x[11]), .Z(n7183) );
  XOR U4321 ( .A(n7182), .B(n7183), .Z(n7234) );
  XOR U4322 ( .A(n7233), .B(n7234), .Z(n7212) );
  XNOR U4323 ( .A(n7211), .B(n7212), .Z(n7237) );
  XOR U4324 ( .A(n7238), .B(n7237), .Z(n7240) );
  XOR U4325 ( .A(n7239), .B(n7240), .Z(n7256) );
  NANDN U4326 ( .A(n7140), .B(n7139), .Z(n7144) );
  NANDN U4327 ( .A(n7142), .B(n7141), .Z(n7143) );
  AND U4328 ( .A(n7144), .B(n7143), .Z(n7255) );
  XNOR U4329 ( .A(n7258), .B(n7257), .Z(n7159) );
  XOR U4330 ( .A(n7161), .B(n7162), .Z(n7168) );
  OR U4331 ( .A(n7147), .B(n7145), .Z(n7151) );
  ANDN U4332 ( .B(n7147), .A(n7146), .Z(n7149) );
  OR U4333 ( .A(n7149), .B(n7148), .Z(n7150) );
  AND U4334 ( .A(n7151), .B(n7150), .Z(n7167) );
  NAND U4335 ( .A(n7153), .B(n7152), .Z(n7157) );
  NAND U4336 ( .A(n7155), .B(n7154), .Z(n7156) );
  NAND U4337 ( .A(n7157), .B(n7156), .Z(n7166) );
  IV U4338 ( .A(n7166), .Z(n7165) );
  XOR U4339 ( .A(n7167), .B(n7165), .Z(n7158) );
  XNOR U4340 ( .A(n7168), .B(n7158), .Z(N50) );
  NANDN U4341 ( .A(n7160), .B(n7159), .Z(n7164) );
  NANDN U4342 ( .A(n7162), .B(n7161), .Z(n7163) );
  AND U4343 ( .A(n7164), .B(n7163), .Z(n7350) );
  OR U4344 ( .A(n7167), .B(n7165), .Z(n7171) );
  ANDN U4345 ( .B(n7167), .A(n7166), .Z(n7169) );
  OR U4346 ( .A(n7169), .B(n7168), .Z(n7170) );
  AND U4347 ( .A(n7171), .B(n7170), .Z(n7349) );
  AND U4348 ( .A(x[6]), .B(y[12]), .Z(n7279) );
  AND U4349 ( .A(x[5]), .B(y[13]), .Z(n7278) );
  XOR U4350 ( .A(n7279), .B(n7278), .Z(n7281) );
  AND U4351 ( .A(y[14]), .B(x[4]), .Z(n7319) );
  AND U4352 ( .A(y[10]), .B(x[8]), .Z(n7318) );
  XOR U4353 ( .A(n7319), .B(n7318), .Z(n7321) );
  AND U4354 ( .A(x[7]), .B(y[11]), .Z(n7320) );
  XOR U4355 ( .A(n7321), .B(n7320), .Z(n7280) );
  XNOR U4356 ( .A(n7281), .B(n7280), .Z(n7331) );
  AND U4357 ( .A(y[2]), .B(x[16]), .Z(n7285) );
  AND U4358 ( .A(y[7]), .B(x[11]), .Z(n7284) );
  XOR U4359 ( .A(n7285), .B(n7284), .Z(n7287) );
  AND U4360 ( .A(x[2]), .B(y[16]), .Z(n7286) );
  XOR U4361 ( .A(n7287), .B(n7286), .Z(n7330) );
  NANDN U4362 ( .A(n7173), .B(n7172), .Z(n7177) );
  NANDN U4363 ( .A(n7175), .B(n7174), .Z(n7176) );
  AND U4364 ( .A(n7177), .B(n7176), .Z(n7329) );
  XOR U4365 ( .A(n7331), .B(n7332), .Z(n7325) );
  AND U4366 ( .A(y[3]), .B(x[15]), .Z(n7290) );
  XOR U4367 ( .A(n7290), .B(n7178), .Z(n7293) );
  AND U4368 ( .A(x[14]), .B(y[4]), .Z(n7292) );
  XOR U4369 ( .A(n7293), .B(n7292), .Z(n7301) );
  AND U4370 ( .A(x[1]), .B(y[17]), .Z(n7311) );
  AND U4371 ( .A(y[8]), .B(x[10]), .Z(n7310) );
  XOR U4372 ( .A(n7311), .B(n7310), .Z(n7313) );
  ANDN U4373 ( .B(o[17]), .A(n7179), .Z(n7312) );
  XNOR U4374 ( .A(n7313), .B(n7312), .Z(n7300) );
  XNOR U4375 ( .A(n7301), .B(n7300), .Z(n7303) );
  NANDN U4376 ( .A(n7181), .B(n7180), .Z(n7185) );
  NANDN U4377 ( .A(n7183), .B(n7182), .Z(n7184) );
  AND U4378 ( .A(n7185), .B(n7184), .Z(n7302) );
  XOR U4379 ( .A(n7303), .B(n7302), .Z(n7324) );
  AND U4380 ( .A(y[5]), .B(x[15]), .Z(n7432) );
  IV U4381 ( .A(n7432), .Z(n7541) );
  NANDN U4382 ( .A(n7541), .B(n7186), .Z(n7190) );
  NANDN U4383 ( .A(n7188), .B(n7187), .Z(n7189) );
  NAND U4384 ( .A(n7190), .B(n7189), .Z(n7323) );
  XOR U4385 ( .A(n7324), .B(n7323), .Z(n7326) );
  XOR U4386 ( .A(n7325), .B(n7326), .Z(n7268) );
  NANDN U4387 ( .A(n7192), .B(n7191), .Z(n7196) );
  OR U4388 ( .A(n7194), .B(n7193), .Z(n7195) );
  AND U4389 ( .A(n7196), .B(n7195), .Z(n7341) );
  NANDN U4390 ( .A(n7198), .B(n7197), .Z(n7202) );
  NANDN U4391 ( .A(n7200), .B(n7199), .Z(n7201) );
  NAND U4392 ( .A(n7202), .B(n7201), .Z(n7342) );
  XNOR U4393 ( .A(n7341), .B(n7342), .Z(n7343) );
  NANDN U4394 ( .A(n7204), .B(n7203), .Z(n7208) );
  NAND U4395 ( .A(n7206), .B(n7205), .Z(n7207) );
  NAND U4396 ( .A(n7208), .B(n7207), .Z(n7344) );
  XNOR U4397 ( .A(n7343), .B(n7344), .Z(n7269) );
  XOR U4398 ( .A(n7268), .B(n7269), .Z(n7271) );
  NANDN U4399 ( .A(n7210), .B(n7209), .Z(n7214) );
  NANDN U4400 ( .A(n7212), .B(n7211), .Z(n7213) );
  AND U4401 ( .A(n7214), .B(n7213), .Z(n7274) );
  NANDN U4402 ( .A(n7216), .B(n7215), .Z(n7220) );
  NANDN U4403 ( .A(n7218), .B(n7217), .Z(n7219) );
  NAND U4404 ( .A(n7220), .B(n7219), .Z(n7296) );
  AND U4405 ( .A(y[15]), .B(x[3]), .Z(n7315) );
  AND U4406 ( .A(x[13]), .B(y[5]), .Z(n7314) );
  XOR U4407 ( .A(n7315), .B(n7314), .Z(n7317) );
  AND U4408 ( .A(y[6]), .B(x[12]), .Z(n7316) );
  XOR U4409 ( .A(n7317), .B(n7316), .Z(n7295) );
  NAND U4410 ( .A(x[17]), .B(y[1]), .Z(n7322) );
  XNOR U4411 ( .A(o[18]), .B(n7322), .Z(n7309) );
  AND U4412 ( .A(x[0]), .B(y[18]), .Z(n7307) );
  AND U4413 ( .A(y[0]), .B(x[18]), .Z(n7306) );
  XOR U4414 ( .A(n7307), .B(n7306), .Z(n7308) );
  XOR U4415 ( .A(n7309), .B(n7308), .Z(n7294) );
  XOR U4416 ( .A(n7295), .B(n7294), .Z(n7297) );
  XNOR U4417 ( .A(n7296), .B(n7297), .Z(n7338) );
  NANDN U4418 ( .A(n7226), .B(n7225), .Z(n7230) );
  NANDN U4419 ( .A(n7228), .B(n7227), .Z(n7229) );
  NAND U4420 ( .A(n7230), .B(n7229), .Z(n7336) );
  XNOR U4421 ( .A(n7335), .B(n7336), .Z(n7337) );
  XOR U4422 ( .A(n7338), .B(n7337), .Z(n7272) );
  NANDN U4423 ( .A(n7232), .B(n7231), .Z(n7236) );
  NANDN U4424 ( .A(n7234), .B(n7233), .Z(n7235) );
  NAND U4425 ( .A(n7236), .B(n7235), .Z(n7273) );
  XOR U4426 ( .A(n7272), .B(n7273), .Z(n7275) );
  XNOR U4427 ( .A(n7274), .B(n7275), .Z(n7270) );
  XOR U4428 ( .A(n7271), .B(n7270), .Z(n7265) );
  NANDN U4429 ( .A(n7238), .B(n7237), .Z(n7242) );
  OR U4430 ( .A(n7240), .B(n7239), .Z(n7241) );
  AND U4431 ( .A(n7242), .B(n7241), .Z(n7263) );
  NANDN U4432 ( .A(n7244), .B(n7243), .Z(n7248) );
  NANDN U4433 ( .A(n7246), .B(n7245), .Z(n7247) );
  AND U4434 ( .A(n7248), .B(n7247), .Z(n7262) );
  XNOR U4435 ( .A(n7263), .B(n7262), .Z(n7264) );
  XNOR U4436 ( .A(n7265), .B(n7264), .Z(n7354) );
  NANDN U4437 ( .A(n7250), .B(n7249), .Z(n7254) );
  NANDN U4438 ( .A(n7252), .B(n7251), .Z(n7253) );
  NAND U4439 ( .A(n7254), .B(n7253), .Z(n7355) );
  NANDN U4440 ( .A(n7256), .B(n7255), .Z(n7260) );
  NAND U4441 ( .A(n7258), .B(n7257), .Z(n7259) );
  AND U4442 ( .A(n7260), .B(n7259), .Z(n7356) );
  XOR U4443 ( .A(n7357), .B(n7356), .Z(n7348) );
  IV U4444 ( .A(n7348), .Z(n7347) );
  XOR U4445 ( .A(n7349), .B(n7347), .Z(n7261) );
  XNOR U4446 ( .A(n7350), .B(n7261), .Z(N51) );
  NANDN U4447 ( .A(n7263), .B(n7262), .Z(n7267) );
  NANDN U4448 ( .A(n7265), .B(n7264), .Z(n7266) );
  AND U4449 ( .A(n7267), .B(n7266), .Z(n7469) );
  NANDN U4450 ( .A(n7273), .B(n7272), .Z(n7277) );
  NANDN U4451 ( .A(n7275), .B(n7274), .Z(n7276) );
  NAND U4452 ( .A(n7277), .B(n7276), .Z(n7450) );
  NAND U4453 ( .A(n7279), .B(n7278), .Z(n7283) );
  NAND U4454 ( .A(n7281), .B(n7280), .Z(n7282) );
  NAND U4455 ( .A(n7283), .B(n7282), .Z(n7382) );
  NAND U4456 ( .A(n7285), .B(n7284), .Z(n7289) );
  NAND U4457 ( .A(n7287), .B(n7286), .Z(n7288) );
  NAND U4458 ( .A(n7289), .B(n7288), .Z(n7380) );
  AND U4459 ( .A(x[1]), .B(y[18]), .Z(n7390) );
  NAND U4460 ( .A(x[8]), .B(y[11]), .Z(n7391) );
  XNOR U4461 ( .A(n7390), .B(n7391), .Z(n7392) );
  NAND U4462 ( .A(y[5]), .B(x[14]), .Z(n7393) );
  XNOR U4463 ( .A(n7392), .B(n7393), .Z(n7441) );
  AND U4464 ( .A(x[2]), .B(y[17]), .Z(n7426) );
  NAND U4465 ( .A(x[13]), .B(y[6]), .Z(n7427) );
  XNOR U4466 ( .A(n7426), .B(n7427), .Z(n7429) );
  AND U4467 ( .A(y[7]), .B(x[12]), .Z(n7428) );
  XOR U4468 ( .A(n7429), .B(n7428), .Z(n7440) );
  XOR U4469 ( .A(n7441), .B(n7440), .Z(n7443) );
  XOR U4470 ( .A(n7442), .B(n7443), .Z(n7381) );
  XOR U4471 ( .A(n7380), .B(n7381), .Z(n7383) );
  XOR U4472 ( .A(n7382), .B(n7383), .Z(n7449) );
  NAND U4473 ( .A(n7295), .B(n7294), .Z(n7299) );
  NAND U4474 ( .A(n7297), .B(n7296), .Z(n7298) );
  NAND U4475 ( .A(n7299), .B(n7298), .Z(n7374) );
  NANDN U4476 ( .A(n7301), .B(n7300), .Z(n7305) );
  NAND U4477 ( .A(n7303), .B(n7302), .Z(n7304) );
  AND U4478 ( .A(n7305), .B(n7304), .Z(n7375) );
  XOR U4479 ( .A(n7374), .B(n7375), .Z(n7376) );
  AND U4480 ( .A(y[10]), .B(x[9]), .Z(n7420) );
  NAND U4481 ( .A(y[3]), .B(x[16]), .Z(n7421) );
  XNOR U4482 ( .A(n7420), .B(n7421), .Z(n7422) );
  NAND U4483 ( .A(y[4]), .B(x[15]), .Z(n7423) );
  XOR U4484 ( .A(n7422), .B(n7423), .Z(n7386) );
  XOR U4485 ( .A(n7386), .B(n7387), .Z(n7388) );
  XNOR U4486 ( .A(n7388), .B(n7389), .Z(n7370) );
  AND U4487 ( .A(x[3]), .B(y[16]), .Z(n7433) );
  NAND U4488 ( .A(y[8]), .B(x[11]), .Z(n7434) );
  XNOR U4489 ( .A(n7433), .B(n7434), .Z(n7435) );
  NAND U4490 ( .A(y[1]), .B(x[18]), .Z(n7439) );
  XNOR U4491 ( .A(o[19]), .B(n7439), .Z(n7399) );
  AND U4492 ( .A(y[2]), .B(x[17]), .Z(n7396) );
  NAND U4493 ( .A(y[9]), .B(x[10]), .Z(n7397) );
  XNOR U4494 ( .A(n7396), .B(n7397), .Z(n7398) );
  XNOR U4495 ( .A(n7399), .B(n7398), .Z(n7414) );
  XNOR U4496 ( .A(n7415), .B(n7414), .Z(n7416) );
  XNOR U4497 ( .A(n7416), .B(n7417), .Z(n7368) );
  ANDN U4498 ( .B(o[18]), .A(n7322), .Z(n7411) );
  AND U4499 ( .A(x[0]), .B(y[19]), .Z(n7409) );
  NAND U4500 ( .A(x[19]), .B(y[0]), .Z(n7408) );
  XNOR U4501 ( .A(n7409), .B(n7408), .Z(n7410) );
  XOR U4502 ( .A(n7411), .B(n7410), .Z(n7445) );
  AND U4503 ( .A(x[5]), .B(y[14]), .Z(n7402) );
  NAND U4504 ( .A(x[6]), .B(y[13]), .Z(n7403) );
  XNOR U4505 ( .A(n7402), .B(n7403), .Z(n7405) );
  AND U4506 ( .A(y[15]), .B(x[4]), .Z(n7404) );
  XOR U4507 ( .A(n7405), .B(n7404), .Z(n7444) );
  XNOR U4508 ( .A(n7445), .B(n7444), .Z(n7447) );
  XOR U4509 ( .A(n7446), .B(n7447), .Z(n7369) );
  XOR U4510 ( .A(n7368), .B(n7369), .Z(n7371) );
  XOR U4511 ( .A(n7370), .B(n7371), .Z(n7377) );
  XOR U4512 ( .A(n7376), .B(n7377), .Z(n7448) );
  XOR U4513 ( .A(n7449), .B(n7448), .Z(n7451) );
  XOR U4514 ( .A(n7450), .B(n7451), .Z(n7457) );
  NANDN U4515 ( .A(n7324), .B(n7323), .Z(n7328) );
  NANDN U4516 ( .A(n7326), .B(n7325), .Z(n7327) );
  NAND U4517 ( .A(n7328), .B(n7327), .Z(n7462) );
  NANDN U4518 ( .A(n7330), .B(n7329), .Z(n7334) );
  NANDN U4519 ( .A(n7332), .B(n7331), .Z(n7333) );
  AND U4520 ( .A(n7334), .B(n7333), .Z(n7461) );
  NANDN U4521 ( .A(n7336), .B(n7335), .Z(n7340) );
  NAND U4522 ( .A(n7338), .B(n7337), .Z(n7339) );
  AND U4523 ( .A(n7340), .B(n7339), .Z(n7460) );
  XOR U4524 ( .A(n7461), .B(n7460), .Z(n7463) );
  XOR U4525 ( .A(n7462), .B(n7463), .Z(n7454) );
  NANDN U4526 ( .A(n7342), .B(n7341), .Z(n7346) );
  NANDN U4527 ( .A(n7344), .B(n7343), .Z(n7345) );
  NAND U4528 ( .A(n7346), .B(n7345), .Z(n7455) );
  XNOR U4529 ( .A(n7454), .B(n7455), .Z(n7456) );
  XOR U4530 ( .A(n7457), .B(n7456), .Z(n7466) );
  XOR U4531 ( .A(n7467), .B(n7466), .Z(n7468) );
  XOR U4532 ( .A(n7469), .B(n7468), .Z(n7364) );
  OR U4533 ( .A(n7349), .B(n7347), .Z(n7353) );
  ANDN U4534 ( .B(n7349), .A(n7348), .Z(n7351) );
  OR U4535 ( .A(n7351), .B(n7350), .Z(n7352) );
  AND U4536 ( .A(n7353), .B(n7352), .Z(n7363) );
  NANDN U4537 ( .A(n7355), .B(n7354), .Z(n7359) );
  NAND U4538 ( .A(n7357), .B(n7356), .Z(n7358) );
  NAND U4539 ( .A(n7359), .B(n7358), .Z(n7362) );
  IV U4540 ( .A(n7362), .Z(n7361) );
  XOR U4541 ( .A(n7363), .B(n7361), .Z(n7360) );
  XNOR U4542 ( .A(n7364), .B(n7360), .Z(N52) );
  OR U4543 ( .A(n7363), .B(n7361), .Z(n7367) );
  ANDN U4544 ( .B(n7363), .A(n7362), .Z(n7365) );
  OR U4545 ( .A(n7365), .B(n7364), .Z(n7366) );
  AND U4546 ( .A(n7367), .B(n7366), .Z(n7592) );
  NANDN U4547 ( .A(n7369), .B(n7368), .Z(n7373) );
  NANDN U4548 ( .A(n7371), .B(n7370), .Z(n7372) );
  AND U4549 ( .A(n7373), .B(n7372), .Z(n7477) );
  NAND U4550 ( .A(n7375), .B(n7374), .Z(n7379) );
  NANDN U4551 ( .A(n7377), .B(n7376), .Z(n7378) );
  AND U4552 ( .A(n7379), .B(n7378), .Z(n7476) );
  XOR U4553 ( .A(n7477), .B(n7476), .Z(n7479) );
  NAND U4554 ( .A(n7381), .B(n7380), .Z(n7385) );
  NAND U4555 ( .A(n7383), .B(n7382), .Z(n7384) );
  AND U4556 ( .A(n7385), .B(n7384), .Z(n7478) );
  XOR U4557 ( .A(n7479), .B(n7478), .Z(n7471) );
  NANDN U4558 ( .A(n7391), .B(n7390), .Z(n7395) );
  NANDN U4559 ( .A(n7393), .B(n7392), .Z(n7394) );
  AND U4560 ( .A(n7395), .B(n7394), .Z(n7519) );
  NANDN U4561 ( .A(n7397), .B(n7396), .Z(n7401) );
  NAND U4562 ( .A(n7399), .B(n7398), .Z(n7400) );
  NAND U4563 ( .A(n7401), .B(n7400), .Z(n7518) );
  XNOR U4564 ( .A(n7519), .B(n7518), .Z(n7520) );
  AND U4565 ( .A(x[13]), .B(y[7]), .Z(n7500) );
  NAND U4566 ( .A(x[3]), .B(y[17]), .Z(n7501) );
  XNOR U4567 ( .A(n7500), .B(n7501), .Z(n7502) );
  NAND U4568 ( .A(y[12]), .B(x[8]), .Z(n7503) );
  XNOR U4569 ( .A(n7502), .B(n7503), .Z(n7561) );
  AND U4570 ( .A(y[15]), .B(x[5]), .Z(n7506) );
  NAND U4571 ( .A(x[4]), .B(y[16]), .Z(n7507) );
  XNOR U4572 ( .A(n7506), .B(n7507), .Z(n7508) );
  NAND U4573 ( .A(x[7]), .B(y[13]), .Z(n7509) );
  XNOR U4574 ( .A(n7508), .B(n7509), .Z(n7559) );
  NAND U4575 ( .A(x[6]), .B(y[14]), .Z(n7560) );
  XOR U4576 ( .A(n7559), .B(n7560), .Z(n7562) );
  XOR U4577 ( .A(n7561), .B(n7562), .Z(n7521) );
  XOR U4578 ( .A(n7520), .B(n7521), .Z(n7572) );
  NANDN U4579 ( .A(n7403), .B(n7402), .Z(n7407) );
  NAND U4580 ( .A(n7405), .B(n7404), .Z(n7406) );
  AND U4581 ( .A(n7407), .B(n7406), .Z(n7567) );
  AND U4582 ( .A(y[8]), .B(x[12]), .Z(n7553) );
  NAND U4583 ( .A(y[2]), .B(x[18]), .Z(n7554) );
  XNOR U4584 ( .A(n7553), .B(n7554), .Z(n7555) );
  NAND U4585 ( .A(y[3]), .B(x[17]), .Z(n7556) );
  XNOR U4586 ( .A(n7555), .B(n7556), .Z(n7565) );
  NANDN U4587 ( .A(n7409), .B(n7408), .Z(n7413) );
  NANDN U4588 ( .A(n7411), .B(n7410), .Z(n7412) );
  NAND U4589 ( .A(n7413), .B(n7412), .Z(n7566) );
  XOR U4590 ( .A(n7565), .B(n7566), .Z(n7568) );
  XNOR U4591 ( .A(n7567), .B(n7568), .Z(n7571) );
  XOR U4592 ( .A(n7572), .B(n7571), .Z(n7574) );
  XOR U4593 ( .A(n7573), .B(n7574), .Z(n7485) );
  NANDN U4594 ( .A(n7415), .B(n7414), .Z(n7419) );
  NAND U4595 ( .A(n7417), .B(n7416), .Z(n7418) );
  AND U4596 ( .A(n7419), .B(n7418), .Z(n7484) );
  XNOR U4597 ( .A(n7485), .B(n7484), .Z(n7487) );
  NANDN U4598 ( .A(n7421), .B(n7420), .Z(n7425) );
  NANDN U4599 ( .A(n7423), .B(n7422), .Z(n7424) );
  AND U4600 ( .A(n7425), .B(n7424), .Z(n7489) );
  NANDN U4601 ( .A(n7427), .B(n7426), .Z(n7431) );
  NAND U4602 ( .A(n7429), .B(n7428), .Z(n7430) );
  AND U4603 ( .A(n7431), .B(n7430), .Z(n7527) );
  AND U4604 ( .A(x[14]), .B(y[6]), .Z(n7544) );
  XOR U4605 ( .A(n7542), .B(n7432), .Z(n7543) );
  XOR U4606 ( .A(n7544), .B(n7543), .Z(n7524) );
  AND U4607 ( .A(x[16]), .B(y[4]), .Z(n7494) );
  NAND U4608 ( .A(x[2]), .B(y[18]), .Z(n7497) );
  XNOR U4609 ( .A(n7496), .B(n7497), .Z(n7525) );
  XOR U4610 ( .A(n7524), .B(n7525), .Z(n7526) );
  XNOR U4611 ( .A(n7527), .B(n7526), .Z(n7488) );
  XNOR U4612 ( .A(n7489), .B(n7488), .Z(n7490) );
  NANDN U4613 ( .A(n7434), .B(n7433), .Z(n7438) );
  NANDN U4614 ( .A(n7436), .B(n7435), .Z(n7437) );
  AND U4615 ( .A(n7438), .B(n7437), .Z(n7531) );
  ANDN U4616 ( .B(o[19]), .A(n7439), .Z(n7514) );
  AND U4617 ( .A(y[20]), .B(x[0]), .Z(n7513) );
  NAND U4618 ( .A(x[20]), .B(y[0]), .Z(n7512) );
  XOR U4619 ( .A(n7513), .B(n7512), .Z(n7515) );
  XOR U4620 ( .A(n7514), .B(n7515), .Z(n7529) );
  AND U4621 ( .A(x[19]), .B(y[1]), .Z(n7540) );
  XOR U4622 ( .A(o[20]), .B(n7540), .Z(n7549) );
  AND U4623 ( .A(y[9]), .B(x[11]), .Z(n7547) );
  NAND U4624 ( .A(x[1]), .B(y[19]), .Z(n7548) );
  XOR U4625 ( .A(n7547), .B(n7548), .Z(n7550) );
  XNOR U4626 ( .A(n7549), .B(n7550), .Z(n7528) );
  XNOR U4627 ( .A(n7529), .B(n7528), .Z(n7530) );
  XOR U4628 ( .A(n7531), .B(n7530), .Z(n7491) );
  XNOR U4629 ( .A(n7490), .B(n7491), .Z(n7537) );
  XOR U4630 ( .A(n7535), .B(n7534), .Z(n7536) );
  XOR U4631 ( .A(n7537), .B(n7536), .Z(n7486) );
  XOR U4632 ( .A(n7487), .B(n7486), .Z(n7470) );
  XNOR U4633 ( .A(n7471), .B(n7470), .Z(n7473) );
  NANDN U4634 ( .A(n7449), .B(n7448), .Z(n7453) );
  NANDN U4635 ( .A(n7451), .B(n7450), .Z(n7452) );
  AND U4636 ( .A(n7453), .B(n7452), .Z(n7472) );
  XOR U4637 ( .A(n7473), .B(n7472), .Z(n7582) );
  NANDN U4638 ( .A(n7455), .B(n7454), .Z(n7459) );
  NAND U4639 ( .A(n7457), .B(n7456), .Z(n7458) );
  AND U4640 ( .A(n7459), .B(n7458), .Z(n7581) );
  XNOR U4641 ( .A(n7582), .B(n7581), .Z(n7583) );
  NAND U4642 ( .A(n7461), .B(n7460), .Z(n7465) );
  NAND U4643 ( .A(n7463), .B(n7462), .Z(n7464) );
  NAND U4644 ( .A(n7465), .B(n7464), .Z(n7584) );
  XNOR U4645 ( .A(n7583), .B(n7584), .Z(n7589) );
  XNOR U4646 ( .A(n7589), .B(n7590), .Z(n7591) );
  XNOR U4647 ( .A(n7592), .B(n7591), .Z(N53) );
  NANDN U4648 ( .A(n7471), .B(n7470), .Z(n7475) );
  NAND U4649 ( .A(n7473), .B(n7472), .Z(n7474) );
  AND U4650 ( .A(n7475), .B(n7474), .Z(n7483) );
  NAND U4651 ( .A(n7477), .B(n7476), .Z(n7481) );
  NAND U4652 ( .A(n7479), .B(n7478), .Z(n7480) );
  NAND U4653 ( .A(n7481), .B(n7480), .Z(n7482) );
  NAND U4654 ( .A(n7483), .B(n7482), .Z(n7578) );
  XOR U4655 ( .A(n7483), .B(n7482), .Z(n7579) );
  NANDN U4656 ( .A(n7489), .B(n7488), .Z(n7493) );
  NANDN U4657 ( .A(n7491), .B(n7490), .Z(n7492) );
  AND U4658 ( .A(n7493), .B(n7492), .Z(n7701) );
  NANDN U4659 ( .A(n7495), .B(n7494), .Z(n7499) );
  NANDN U4660 ( .A(n7497), .B(n7496), .Z(n7498) );
  AND U4661 ( .A(n7499), .B(n7498), .Z(n7628) );
  NANDN U4662 ( .A(n7501), .B(n7500), .Z(n7505) );
  NANDN U4663 ( .A(n7503), .B(n7502), .Z(n7504) );
  AND U4664 ( .A(n7505), .B(n7504), .Z(n7618) );
  NAND U4665 ( .A(x[1]), .B(y[20]), .Z(n7676) );
  NAND U4666 ( .A(x[10]), .B(y[11]), .Z(n7675) );
  NAND U4667 ( .A(y[3]), .B(x[18]), .Z(n7674) );
  XNOR U4668 ( .A(n7675), .B(n7674), .Z(n7677) );
  XOR U4669 ( .A(n7676), .B(n7677), .Z(n7616) );
  NAND U4670 ( .A(x[20]), .B(y[1]), .Z(n7661) );
  XNOR U4671 ( .A(o[21]), .B(n7661), .Z(n7646) );
  AND U4672 ( .A(x[19]), .B(y[2]), .Z(n7644) );
  AND U4673 ( .A(y[10]), .B(x[11]), .Z(n7643) );
  XOR U4674 ( .A(n7644), .B(n7643), .Z(n7645) );
  XOR U4675 ( .A(n7646), .B(n7645), .Z(n7615) );
  XOR U4676 ( .A(n7616), .B(n7615), .Z(n7617) );
  XNOR U4677 ( .A(n7618), .B(n7617), .Z(n7627) );
  XNOR U4678 ( .A(n7628), .B(n7627), .Z(n7630) );
  NANDN U4679 ( .A(n7507), .B(n7506), .Z(n7511) );
  NANDN U4680 ( .A(n7509), .B(n7508), .Z(n7510) );
  AND U4681 ( .A(n7511), .B(n7510), .Z(n7612) );
  NANDN U4682 ( .A(n7513), .B(n7512), .Z(n7517) );
  OR U4683 ( .A(n7515), .B(n7514), .Z(n7516) );
  AND U4684 ( .A(n7517), .B(n7516), .Z(n7611) );
  XNOR U4685 ( .A(n7612), .B(n7611), .Z(n7614) );
  AND U4686 ( .A(y[7]), .B(x[14]), .Z(n7669) );
  AND U4687 ( .A(y[15]), .B(x[6]), .Z(n7668) );
  XOR U4688 ( .A(n7669), .B(n7668), .Z(n7671) );
  AND U4689 ( .A(y[14]), .B(x[7]), .Z(n7670) );
  XOR U4690 ( .A(n7671), .B(n7670), .Z(n7634) );
  NAND U4691 ( .A(x[8]), .B(y[13]), .Z(n7632) );
  NAND U4692 ( .A(y[12]), .B(x[9]), .Z(n7631) );
  XOR U4693 ( .A(n7632), .B(n7631), .Z(n7633) );
  XNOR U4694 ( .A(n7634), .B(n7633), .Z(n7652) );
  AND U4695 ( .A(x[3]), .B(y[18]), .Z(n7656) );
  AND U4696 ( .A(x[13]), .B(y[8]), .Z(n7655) );
  XOR U4697 ( .A(n7656), .B(n7655), .Z(n7658) );
  AND U4698 ( .A(x[4]), .B(y[17]), .Z(n7657) );
  XOR U4699 ( .A(n7658), .B(n7657), .Z(n7650) );
  AND U4700 ( .A(y[9]), .B(x[12]), .Z(n7638) );
  AND U4701 ( .A(y[4]), .B(x[17]), .Z(n7637) );
  XOR U4702 ( .A(n7638), .B(n7637), .Z(n7640) );
  AND U4703 ( .A(x[2]), .B(y[19]), .Z(n7639) );
  XOR U4704 ( .A(n7640), .B(n7639), .Z(n7649) );
  XOR U4705 ( .A(n7650), .B(n7649), .Z(n7651) );
  XNOR U4706 ( .A(n7652), .B(n7651), .Z(n7613) );
  XOR U4707 ( .A(n7614), .B(n7613), .Z(n7629) );
  XOR U4708 ( .A(n7630), .B(n7629), .Z(n7698) );
  NANDN U4709 ( .A(n7519), .B(n7518), .Z(n7523) );
  NANDN U4710 ( .A(n7521), .B(n7520), .Z(n7522) );
  AND U4711 ( .A(n7523), .B(n7522), .Z(n7695) );
  NANDN U4712 ( .A(n7529), .B(n7528), .Z(n7533) );
  NANDN U4713 ( .A(n7531), .B(n7530), .Z(n7532) );
  NAND U4714 ( .A(n7533), .B(n7532), .Z(n7692) );
  XNOR U4715 ( .A(n7693), .B(n7692), .Z(n7694) );
  XOR U4716 ( .A(n7695), .B(n7694), .Z(n7699) );
  XNOR U4717 ( .A(n7698), .B(n7699), .Z(n7700) );
  XNOR U4718 ( .A(n7701), .B(n7700), .Z(n7596) );
  XOR U4719 ( .A(n7595), .B(n7596), .Z(n7597) );
  NAND U4720 ( .A(n7535), .B(n7534), .Z(n7539) );
  NAND U4721 ( .A(n7537), .B(n7536), .Z(n7538) );
  NAND U4722 ( .A(n7539), .B(n7538), .Z(n7601) );
  AND U4723 ( .A(n7540), .B(o[20]), .Z(n7683) );
  AND U4724 ( .A(x[21]), .B(y[0]), .Z(n7681) );
  AND U4725 ( .A(y[21]), .B(x[0]), .Z(n7680) );
  XOR U4726 ( .A(n7681), .B(n7680), .Z(n7682) );
  XOR U4727 ( .A(n7683), .B(n7682), .Z(n7687) );
  AND U4728 ( .A(y[5]), .B(x[16]), .Z(n7662) );
  NAND U4729 ( .A(x[5]), .B(y[16]), .Z(n7663) );
  XNOR U4730 ( .A(n7662), .B(n7663), .Z(n7665) );
  AND U4731 ( .A(y[6]), .B(x[15]), .Z(n7664) );
  XOR U4732 ( .A(n7665), .B(n7664), .Z(n7686) );
  XOR U4733 ( .A(n7687), .B(n7686), .Z(n7689) );
  NANDN U4734 ( .A(n7542), .B(n7541), .Z(n7546) );
  NANDN U4735 ( .A(n7544), .B(n7543), .Z(n7545) );
  AND U4736 ( .A(n7546), .B(n7545), .Z(n7688) );
  XOR U4737 ( .A(n7689), .B(n7688), .Z(n7608) );
  NANDN U4738 ( .A(n7548), .B(n7547), .Z(n7552) );
  NANDN U4739 ( .A(n7550), .B(n7549), .Z(n7551) );
  AND U4740 ( .A(n7552), .B(n7551), .Z(n7606) );
  NANDN U4741 ( .A(n7554), .B(n7553), .Z(n7558) );
  NANDN U4742 ( .A(n7556), .B(n7555), .Z(n7557) );
  NAND U4743 ( .A(n7558), .B(n7557), .Z(n7605) );
  XNOR U4744 ( .A(n7606), .B(n7605), .Z(n7607) );
  XOR U4745 ( .A(n7608), .B(n7607), .Z(n7622) );
  NANDN U4746 ( .A(n7560), .B(n7559), .Z(n7564) );
  NANDN U4747 ( .A(n7562), .B(n7561), .Z(n7563) );
  AND U4748 ( .A(n7564), .B(n7563), .Z(n7621) );
  XNOR U4749 ( .A(n7622), .B(n7621), .Z(n7623) );
  NANDN U4750 ( .A(n7566), .B(n7565), .Z(n7570) );
  OR U4751 ( .A(n7568), .B(n7567), .Z(n7569) );
  NAND U4752 ( .A(n7570), .B(n7569), .Z(n7624) );
  XOR U4753 ( .A(n7623), .B(n7624), .Z(n7599) );
  NAND U4754 ( .A(n7572), .B(n7571), .Z(n7576) );
  NAND U4755 ( .A(n7574), .B(n7573), .Z(n7575) );
  AND U4756 ( .A(n7576), .B(n7575), .Z(n7600) );
  XNOR U4757 ( .A(n7599), .B(n7600), .Z(n7602) );
  XOR U4758 ( .A(n7597), .B(n7598), .Z(n7580) );
  NAND U4759 ( .A(n7579), .B(n7580), .Z(n7577) );
  NAND U4760 ( .A(n7578), .B(n7577), .Z(n7946) );
  XNOR U4761 ( .A(n7580), .B(n7579), .Z(n7588) );
  NANDN U4762 ( .A(n7582), .B(n7581), .Z(n7586) );
  NANDN U4763 ( .A(n7584), .B(n7583), .Z(n7585) );
  AND U4764 ( .A(n7586), .B(n7585), .Z(n7587) );
  XOR U4765 ( .A(n7588), .B(n7587), .Z(n8915) );
  NANDN U4766 ( .A(n7590), .B(n7589), .Z(n7594) );
  NAND U4767 ( .A(n7592), .B(n7591), .Z(n7593) );
  AND U4768 ( .A(n7594), .B(n7593), .Z(n8914) );
  NAND U4769 ( .A(n7600), .B(n7599), .Z(n7604) );
  NANDN U4770 ( .A(n7602), .B(n7601), .Z(n7603) );
  NAND U4771 ( .A(n7604), .B(n7603), .Z(n7947) );
  NANDN U4772 ( .A(n7606), .B(n7605), .Z(n7610) );
  NAND U4773 ( .A(n7608), .B(n7607), .Z(n7609) );
  AND U4774 ( .A(n7610), .B(n7609), .Z(n7714) );
  NAND U4775 ( .A(n7616), .B(n7615), .Z(n7620) );
  NANDN U4776 ( .A(n7618), .B(n7617), .Z(n7619) );
  NAND U4777 ( .A(n7620), .B(n7619), .Z(n7711) );
  XNOR U4778 ( .A(n7712), .B(n7711), .Z(n7713) );
  XNOR U4779 ( .A(n7714), .B(n7713), .Z(n7705) );
  NANDN U4780 ( .A(n7622), .B(n7621), .Z(n7626) );
  NANDN U4781 ( .A(n7624), .B(n7623), .Z(n7625) );
  NAND U4782 ( .A(n7626), .B(n7625), .Z(n7706) );
  XNOR U4783 ( .A(n7705), .B(n7706), .Z(n7707) );
  NAND U4784 ( .A(n7632), .B(n7631), .Z(n7636) );
  NANDN U4785 ( .A(n7634), .B(n7633), .Z(n7635) );
  AND U4786 ( .A(n7636), .B(n7635), .Z(n7792) );
  NAND U4787 ( .A(n7638), .B(n7637), .Z(n7642) );
  NAND U4788 ( .A(n7640), .B(n7639), .Z(n7641) );
  AND U4789 ( .A(n7642), .B(n7641), .Z(n7760) );
  AND U4790 ( .A(x[5]), .B(y[17]), .Z(n7745) );
  NAND U4791 ( .A(y[5]), .B(x[17]), .Z(n7746) );
  XNOR U4792 ( .A(n7745), .B(n7746), .Z(n7747) );
  NAND U4793 ( .A(x[16]), .B(y[6]), .Z(n7748) );
  XNOR U4794 ( .A(n7747), .B(n7748), .Z(n7758) );
  AND U4795 ( .A(y[10]), .B(x[12]), .Z(n7727) );
  NAND U4796 ( .A(y[4]), .B(x[18]), .Z(n7728) );
  XNOR U4797 ( .A(n7727), .B(n7728), .Z(n7729) );
  NAND U4798 ( .A(x[4]), .B(y[18]), .Z(n7730) );
  XOR U4799 ( .A(n7729), .B(n7730), .Z(n7759) );
  XOR U4800 ( .A(n7758), .B(n7759), .Z(n7761) );
  XOR U4801 ( .A(n7760), .B(n7761), .Z(n7791) );
  NAND U4802 ( .A(n7644), .B(n7643), .Z(n7648) );
  NAND U4803 ( .A(n7646), .B(n7645), .Z(n7647) );
  AND U4804 ( .A(n7648), .B(n7647), .Z(n7790) );
  XOR U4805 ( .A(n7791), .B(n7790), .Z(n7793) );
  XOR U4806 ( .A(n7792), .B(n7793), .Z(n7807) );
  NAND U4807 ( .A(n7650), .B(n7649), .Z(n7654) );
  NANDN U4808 ( .A(n7652), .B(n7651), .Z(n7653) );
  AND U4809 ( .A(n7654), .B(n7653), .Z(n7803) );
  NAND U4810 ( .A(n7656), .B(n7655), .Z(n7660) );
  NAND U4811 ( .A(n7658), .B(n7657), .Z(n7659) );
  AND U4812 ( .A(n7660), .B(n7659), .Z(n7777) );
  AND U4813 ( .A(x[3]), .B(y[19]), .Z(n7764) );
  NAND U4814 ( .A(y[8]), .B(x[14]), .Z(n7765) );
  XNOR U4815 ( .A(n7764), .B(n7765), .Z(n7766) );
  NAND U4816 ( .A(x[19]), .B(y[3]), .Z(n7767) );
  XNOR U4817 ( .A(n7766), .B(n7767), .Z(n7775) );
  AND U4818 ( .A(y[21]), .B(x[1]), .Z(n7770) );
  ANDN U4819 ( .B(o[21]), .A(n7661), .Z(n7772) );
  XOR U4820 ( .A(n7773), .B(n7772), .Z(n7774) );
  XOR U4821 ( .A(n7775), .B(n7774), .Z(n7776) );
  XOR U4822 ( .A(n7777), .B(n7776), .Z(n7796) );
  NANDN U4823 ( .A(n7663), .B(n7662), .Z(n7667) );
  NAND U4824 ( .A(n7665), .B(n7664), .Z(n7666) );
  AND U4825 ( .A(n7667), .B(n7666), .Z(n7720) );
  AND U4826 ( .A(x[20]), .B(y[2]), .Z(n7739) );
  NAND U4827 ( .A(x[13]), .B(y[9]), .Z(n7740) );
  XNOR U4828 ( .A(n7739), .B(n7740), .Z(n7741) );
  NAND U4829 ( .A(x[2]), .B(y[20]), .Z(n7742) );
  XNOR U4830 ( .A(n7741), .B(n7742), .Z(n7718) );
  AND U4831 ( .A(y[7]), .B(x[15]), .Z(n7752) );
  NAND U4832 ( .A(x[6]), .B(y[16]), .Z(n7753) );
  XNOR U4833 ( .A(n7752), .B(n7753), .Z(n7754) );
  XOR U4834 ( .A(n7718), .B(n7717), .Z(n7719) );
  XOR U4835 ( .A(n7720), .B(n7719), .Z(n7797) );
  XOR U4836 ( .A(n7796), .B(n7797), .Z(n7799) );
  NAND U4837 ( .A(n7669), .B(n7668), .Z(n7673) );
  NAND U4838 ( .A(n7671), .B(n7670), .Z(n7672) );
  AND U4839 ( .A(n7673), .B(n7672), .Z(n7780) );
  AND U4840 ( .A(x[21]), .B(y[1]), .Z(n7751) );
  XOR U4841 ( .A(n7751), .B(o[22]), .Z(n7735) );
  AND U4842 ( .A(y[22]), .B(x[0]), .Z(n7734) );
  NAND U4843 ( .A(y[0]), .B(x[22]), .Z(n7733) );
  XOR U4844 ( .A(n7734), .B(n7733), .Z(n7736) );
  XOR U4845 ( .A(n7735), .B(n7736), .Z(n7779) );
  AND U4846 ( .A(y[15]), .B(x[7]), .Z(n7721) );
  NAND U4847 ( .A(y[14]), .B(x[8]), .Z(n7722) );
  XNOR U4848 ( .A(n7721), .B(n7722), .Z(n7723) );
  NAND U4849 ( .A(x[9]), .B(y[13]), .Z(n7724) );
  XNOR U4850 ( .A(n7723), .B(n7724), .Z(n7778) );
  XOR U4851 ( .A(n7779), .B(n7778), .Z(n7781) );
  XOR U4852 ( .A(n7780), .B(n7781), .Z(n7787) );
  NAND U4853 ( .A(n7675), .B(n7674), .Z(n7679) );
  NANDN U4854 ( .A(n7677), .B(n7676), .Z(n7678) );
  AND U4855 ( .A(n7679), .B(n7678), .Z(n7785) );
  NAND U4856 ( .A(n7681), .B(n7680), .Z(n7685) );
  NAND U4857 ( .A(n7683), .B(n7682), .Z(n7684) );
  AND U4858 ( .A(n7685), .B(n7684), .Z(n7784) );
  XNOR U4859 ( .A(n7785), .B(n7784), .Z(n7786) );
  XNOR U4860 ( .A(n7787), .B(n7786), .Z(n7798) );
  XOR U4861 ( .A(n7799), .B(n7798), .Z(n7801) );
  NAND U4862 ( .A(n7687), .B(n7686), .Z(n7691) );
  NAND U4863 ( .A(n7689), .B(n7688), .Z(n7690) );
  NAND U4864 ( .A(n7691), .B(n7690), .Z(n7800) );
  XNOR U4865 ( .A(n7801), .B(n7800), .Z(n7802) );
  XNOR U4866 ( .A(n7803), .B(n7802), .Z(n7806) );
  XNOR U4867 ( .A(n7807), .B(n7806), .Z(n7808) );
  XOR U4868 ( .A(n7809), .B(n7808), .Z(n7708) );
  XNOR U4869 ( .A(n7707), .B(n7708), .Z(n7817) );
  NANDN U4870 ( .A(n7693), .B(n7692), .Z(n7697) );
  NANDN U4871 ( .A(n7695), .B(n7694), .Z(n7696) );
  AND U4872 ( .A(n7697), .B(n7696), .Z(n7815) );
  NANDN U4873 ( .A(n7699), .B(n7698), .Z(n7703) );
  NANDN U4874 ( .A(n7701), .B(n7700), .Z(n7702) );
  NAND U4875 ( .A(n7703), .B(n7702), .Z(n7814) );
  XNOR U4876 ( .A(n7815), .B(n7814), .Z(n7816) );
  XOR U4877 ( .A(n7817), .B(n7816), .Z(n7948) );
  XNOR U4878 ( .A(n7947), .B(n7948), .Z(n7950) );
  XOR U4879 ( .A(n7944), .B(n7945), .Z(n7704) );
  XNOR U4880 ( .A(n7946), .B(n7704), .Z(N55) );
  NANDN U4881 ( .A(n7706), .B(n7705), .Z(n7710) );
  NANDN U4882 ( .A(n7708), .B(n7707), .Z(n7709) );
  NAND U4883 ( .A(n7710), .B(n7709), .Z(n7812) );
  NANDN U4884 ( .A(n7712), .B(n7711), .Z(n7716) );
  NANDN U4885 ( .A(n7714), .B(n7713), .Z(n7715) );
  NAND U4886 ( .A(n7716), .B(n7715), .Z(n7922) );
  AND U4887 ( .A(y[1]), .B(x[22]), .Z(n7897) );
  XOR U4888 ( .A(n7897), .B(o[23]), .Z(n7889) );
  AND U4889 ( .A(x[23]), .B(y[0]), .Z(n7887) );
  NAND U4890 ( .A(y[23]), .B(x[0]), .Z(n7886) );
  XNOR U4891 ( .A(n7887), .B(n7886), .Z(n7888) );
  XOR U4892 ( .A(n7889), .B(n7888), .Z(n7829) );
  NANDN U4893 ( .A(n7722), .B(n7721), .Z(n7726) );
  NANDN U4894 ( .A(n7724), .B(n7723), .Z(n7725) );
  NAND U4895 ( .A(n7726), .B(n7725), .Z(n7828) );
  XOR U4896 ( .A(n7829), .B(n7828), .Z(n7831) );
  AND U4897 ( .A(x[20]), .B(y[3]), .Z(n8496) );
  AND U4898 ( .A(y[7]), .B(x[16]), .Z(n7892) );
  XOR U4899 ( .A(n8496), .B(n7892), .Z(n7894) );
  AND U4900 ( .A(x[19]), .B(y[4]), .Z(n7893) );
  XOR U4901 ( .A(n7894), .B(n7893), .Z(n7830) );
  XOR U4902 ( .A(n7831), .B(n7830), .Z(n7824) );
  NANDN U4903 ( .A(n7728), .B(n7727), .Z(n7732) );
  NANDN U4904 ( .A(n7730), .B(n7729), .Z(n7731) );
  NAND U4905 ( .A(n7732), .B(n7731), .Z(n7822) );
  NANDN U4906 ( .A(n7734), .B(n7733), .Z(n7738) );
  OR U4907 ( .A(n7736), .B(n7735), .Z(n7737) );
  AND U4908 ( .A(n7738), .B(n7737), .Z(n7823) );
  XNOR U4909 ( .A(n7822), .B(n7823), .Z(n7825) );
  XNOR U4910 ( .A(n7824), .B(n7825), .Z(n7882) );
  XNOR U4911 ( .A(n7883), .B(n7882), .Z(n7885) );
  NANDN U4912 ( .A(n7740), .B(n7739), .Z(n7744) );
  NANDN U4913 ( .A(n7742), .B(n7741), .Z(n7743) );
  AND U4914 ( .A(n7744), .B(n7743), .Z(n7917) );
  NANDN U4915 ( .A(n7746), .B(n7745), .Z(n7750) );
  NANDN U4916 ( .A(n7748), .B(n7747), .Z(n7749) );
  NAND U4917 ( .A(n7750), .B(n7749), .Z(n7842) );
  NAND U4918 ( .A(n7751), .B(o[22]), .Z(n7912) );
  NAND U4919 ( .A(x[1]), .B(y[22]), .Z(n7911) );
  NAND U4920 ( .A(x[12]), .B(y[11]), .Z(n7910) );
  XOR U4921 ( .A(n7911), .B(n7910), .Z(n7913) );
  XOR U4922 ( .A(n7912), .B(n7913), .Z(n7841) );
  NAND U4923 ( .A(x[21]), .B(y[2]), .Z(n7860) );
  NAND U4924 ( .A(y[21]), .B(x[2]), .Z(n7859) );
  NAND U4925 ( .A(x[13]), .B(y[10]), .Z(n7858) );
  XNOR U4926 ( .A(n7859), .B(n7858), .Z(n7861) );
  XOR U4927 ( .A(n7860), .B(n7861), .Z(n7840) );
  XNOR U4928 ( .A(n7841), .B(n7840), .Z(n7843) );
  XOR U4929 ( .A(n7842), .B(n7843), .Z(n7916) );
  XNOR U4930 ( .A(n7917), .B(n7916), .Z(n7919) );
  NANDN U4931 ( .A(n7753), .B(n7752), .Z(n7757) );
  NANDN U4932 ( .A(n7755), .B(n7754), .Z(n7756) );
  NAND U4933 ( .A(n7757), .B(n7756), .Z(n7836) );
  AND U4934 ( .A(x[17]), .B(y[6]), .Z(n7855) );
  AND U4935 ( .A(x[5]), .B(y[18]), .Z(n7853) );
  NAND U4936 ( .A(y[5]), .B(x[18]), .Z(n7852) );
  XNOR U4937 ( .A(n7853), .B(n7852), .Z(n7854) );
  XOR U4938 ( .A(n7855), .B(n7854), .Z(n7834) );
  AND U4939 ( .A(x[3]), .B(y[20]), .Z(n7865) );
  AND U4940 ( .A(x[14]), .B(y[9]), .Z(n7864) );
  XOR U4941 ( .A(n7865), .B(n7864), .Z(n7867) );
  AND U4942 ( .A(x[4]), .B(y[19]), .Z(n7866) );
  XOR U4943 ( .A(n7867), .B(n7866), .Z(n7835) );
  XOR U4944 ( .A(n7834), .B(n7835), .Z(n7837) );
  XOR U4945 ( .A(n7836), .B(n7837), .Z(n7918) );
  XOR U4946 ( .A(n7919), .B(n7918), .Z(n7884) );
  XOR U4947 ( .A(n7885), .B(n7884), .Z(n7921) );
  NANDN U4948 ( .A(n7759), .B(n7758), .Z(n7763) );
  OR U4949 ( .A(n7761), .B(n7760), .Z(n7762) );
  NAND U4950 ( .A(n7763), .B(n7762), .Z(n7926) );
  AND U4951 ( .A(y[8]), .B(x[15]), .Z(n7898) );
  NAND U4952 ( .A(x[6]), .B(y[17]), .Z(n7899) );
  XNOR U4953 ( .A(n7898), .B(n7899), .Z(n7901) );
  AND U4954 ( .A(y[12]), .B(x[11]), .Z(n7900) );
  XOR U4955 ( .A(n7901), .B(n7900), .Z(n7872) );
  AND U4956 ( .A(x[10]), .B(y[13]), .Z(n7871) );
  AND U4957 ( .A(x[7]), .B(y[16]), .Z(n7904) );
  NAND U4958 ( .A(y[14]), .B(x[9]), .Z(n7905) );
  XNOR U4959 ( .A(n7904), .B(n7905), .Z(n7907) );
  AND U4960 ( .A(y[15]), .B(x[8]), .Z(n7906) );
  XNOR U4961 ( .A(n7907), .B(n7906), .Z(n7870) );
  XOR U4962 ( .A(n7871), .B(n7870), .Z(n7873) );
  XOR U4963 ( .A(n7872), .B(n7873), .Z(n7849) );
  NANDN U4964 ( .A(n7765), .B(n7764), .Z(n7769) );
  NANDN U4965 ( .A(n7767), .B(n7766), .Z(n7768) );
  AND U4966 ( .A(n7769), .B(n7768), .Z(n7847) );
  XNOR U4967 ( .A(n7847), .B(n7846), .Z(n7848) );
  XNOR U4968 ( .A(n7849), .B(n7848), .Z(n7927) );
  XOR U4969 ( .A(n7926), .B(n7927), .Z(n7929) );
  NANDN U4970 ( .A(n7779), .B(n7778), .Z(n7783) );
  OR U4971 ( .A(n7781), .B(n7780), .Z(n7782) );
  NAND U4972 ( .A(n7783), .B(n7782), .Z(n7876) );
  XOR U4973 ( .A(n7877), .B(n7876), .Z(n7879) );
  NANDN U4974 ( .A(n7785), .B(n7784), .Z(n7789) );
  NANDN U4975 ( .A(n7787), .B(n7786), .Z(n7788) );
  AND U4976 ( .A(n7789), .B(n7788), .Z(n7878) );
  XOR U4977 ( .A(n7879), .B(n7878), .Z(n7928) );
  XOR U4978 ( .A(n7929), .B(n7928), .Z(n7920) );
  XOR U4979 ( .A(n7921), .B(n7920), .Z(n7923) );
  XOR U4980 ( .A(n7922), .B(n7923), .Z(n7941) );
  NANDN U4981 ( .A(n7791), .B(n7790), .Z(n7795) );
  OR U4982 ( .A(n7793), .B(n7792), .Z(n7794) );
  NAND U4983 ( .A(n7795), .B(n7794), .Z(n7933) );
  XOR U4984 ( .A(n7933), .B(n7932), .Z(n7935) );
  NANDN U4985 ( .A(n7801), .B(n7800), .Z(n7805) );
  NANDN U4986 ( .A(n7803), .B(n7802), .Z(n7804) );
  AND U4987 ( .A(n7805), .B(n7804), .Z(n7934) );
  XOR U4988 ( .A(n7935), .B(n7934), .Z(n7939) );
  NANDN U4989 ( .A(n7807), .B(n7806), .Z(n7811) );
  NANDN U4990 ( .A(n7809), .B(n7808), .Z(n7810) );
  AND U4991 ( .A(n7811), .B(n7810), .Z(n7938) );
  XOR U4992 ( .A(n7939), .B(n7938), .Z(n7940) );
  XNOR U4993 ( .A(n7941), .B(n7940), .Z(n7813) );
  NANDN U4994 ( .A(n7812), .B(n7813), .Z(n7821) );
  XNOR U4995 ( .A(n7813), .B(n7812), .Z(n7956) );
  NANDN U4996 ( .A(n7815), .B(n7814), .Z(n7819) );
  NAND U4997 ( .A(n7817), .B(n7816), .Z(n7818) );
  AND U4998 ( .A(n7819), .B(n7818), .Z(n7955) );
  NAND U4999 ( .A(n7956), .B(n7955), .Z(n7820) );
  AND U5000 ( .A(n7821), .B(n7820), .Z(n7960) );
  NAND U5001 ( .A(n7823), .B(n7822), .Z(n7827) );
  NANDN U5002 ( .A(n7825), .B(n7824), .Z(n7826) );
  AND U5003 ( .A(n7827), .B(n7826), .Z(n7972) );
  NAND U5004 ( .A(n7829), .B(n7828), .Z(n7833) );
  NAND U5005 ( .A(n7831), .B(n7830), .Z(n7832) );
  AND U5006 ( .A(n7833), .B(n7832), .Z(n7970) );
  NAND U5007 ( .A(n7835), .B(n7834), .Z(n7839) );
  NAND U5008 ( .A(n7837), .B(n7836), .Z(n7838) );
  AND U5009 ( .A(n7839), .B(n7838), .Z(n7969) );
  XOR U5010 ( .A(n7970), .B(n7969), .Z(n7971) );
  XOR U5011 ( .A(n7972), .B(n7971), .Z(n7964) );
  NANDN U5012 ( .A(n7841), .B(n7840), .Z(n7845) );
  NAND U5013 ( .A(n7843), .B(n7842), .Z(n7844) );
  NAND U5014 ( .A(n7845), .B(n7844), .Z(n7963) );
  XNOR U5015 ( .A(n7964), .B(n7963), .Z(n7965) );
  NANDN U5016 ( .A(n7847), .B(n7846), .Z(n7851) );
  NANDN U5017 ( .A(n7849), .B(n7848), .Z(n7850) );
  AND U5018 ( .A(n7851), .B(n7850), .Z(n8071) );
  AND U5019 ( .A(x[24]), .B(y[0]), .Z(n8056) );
  NAND U5020 ( .A(x[0]), .B(y[24]), .Z(n8057) );
  XNOR U5021 ( .A(n8056), .B(n8057), .Z(n8058) );
  NAND U5022 ( .A(x[23]), .B(y[1]), .Z(n8037) );
  XOR U5023 ( .A(o[24]), .B(n8037), .Z(n8059) );
  XNOR U5024 ( .A(n8058), .B(n8059), .Z(n7986) );
  AND U5025 ( .A(x[7]), .B(y[17]), .Z(n8032) );
  AND U5026 ( .A(y[6]), .B(x[18]), .Z(n8031) );
  XOR U5027 ( .A(n8032), .B(n8031), .Z(n8034) );
  AND U5028 ( .A(y[7]), .B(x[17]), .Z(n8033) );
  XOR U5029 ( .A(n8034), .B(n8033), .Z(n7985) );
  XOR U5030 ( .A(n7986), .B(n7985), .Z(n7987) );
  NANDN U5031 ( .A(n7853), .B(n7852), .Z(n7857) );
  NANDN U5032 ( .A(n7855), .B(n7854), .Z(n7856) );
  NAND U5033 ( .A(n7857), .B(n7856), .Z(n7988) );
  XOR U5034 ( .A(n7987), .B(n7988), .Z(n8003) );
  NAND U5035 ( .A(n7859), .B(n7858), .Z(n7863) );
  NANDN U5036 ( .A(n7861), .B(n7860), .Z(n7862) );
  NAND U5037 ( .A(n7863), .B(n7862), .Z(n8001) );
  NAND U5038 ( .A(n7865), .B(n7864), .Z(n7869) );
  NAND U5039 ( .A(n7867), .B(n7866), .Z(n7868) );
  AND U5040 ( .A(n7869), .B(n7868), .Z(n8002) );
  XNOR U5041 ( .A(n8001), .B(n8002), .Z(n8004) );
  XOR U5042 ( .A(n8003), .B(n8004), .Z(n8069) );
  NANDN U5043 ( .A(n7871), .B(n7870), .Z(n7875) );
  OR U5044 ( .A(n7873), .B(n7872), .Z(n7874) );
  AND U5045 ( .A(n7875), .B(n7874), .Z(n8068) );
  XOR U5046 ( .A(n8069), .B(n8068), .Z(n8070) );
  XOR U5047 ( .A(n8071), .B(n8070), .Z(n7966) );
  XOR U5048 ( .A(n7965), .B(n7966), .Z(n8080) );
  NAND U5049 ( .A(n7877), .B(n7876), .Z(n7881) );
  NAND U5050 ( .A(n7879), .B(n7878), .Z(n7880) );
  AND U5051 ( .A(n7881), .B(n7880), .Z(n8081) );
  XOR U5052 ( .A(n8080), .B(n8081), .Z(n8083) );
  AND U5053 ( .A(y[13]), .B(x[11]), .Z(n8046) );
  AND U5054 ( .A(x[14]), .B(y[10]), .Z(n8045) );
  NAND U5055 ( .A(x[8]), .B(y[16]), .Z(n8044) );
  XOR U5056 ( .A(n8045), .B(n8044), .Z(n8047) );
  XOR U5057 ( .A(n8046), .B(n8047), .Z(n8041) );
  AND U5058 ( .A(y[15]), .B(x[9]), .Z(n8038) );
  NAND U5059 ( .A(y[14]), .B(x[10]), .Z(n8039) );
  XNOR U5060 ( .A(n8038), .B(n8039), .Z(n8040) );
  XOR U5061 ( .A(n8041), .B(n8040), .Z(n8064) );
  NANDN U5062 ( .A(n7887), .B(n7886), .Z(n7891) );
  NANDN U5063 ( .A(n7889), .B(n7888), .Z(n7890) );
  NAND U5064 ( .A(n7891), .B(n7890), .Z(n8063) );
  AND U5065 ( .A(x[3]), .B(y[21]), .Z(n8050) );
  NAND U5066 ( .A(y[9]), .B(x[15]), .Z(n8051) );
  XNOR U5067 ( .A(n8050), .B(n8051), .Z(n8053) );
  AND U5068 ( .A(y[20]), .B(x[4]), .Z(n8052) );
  XNOR U5069 ( .A(n8053), .B(n8052), .Z(n8062) );
  XOR U5070 ( .A(n8063), .B(n8062), .Z(n8065) );
  XOR U5071 ( .A(n8064), .B(n8065), .Z(n8016) );
  NAND U5072 ( .A(n8496), .B(n7892), .Z(n7896) );
  AND U5073 ( .A(n7894), .B(n7893), .Z(n7895) );
  ANDN U5074 ( .B(n7896), .A(n7895), .Z(n7978) );
  AND U5075 ( .A(y[23]), .B(x[1]), .Z(n8027) );
  XOR U5076 ( .A(n8028), .B(n8027), .Z(n8026) );
  AND U5077 ( .A(n7897), .B(o[23]), .Z(n8025) );
  XOR U5078 ( .A(n8026), .B(n8025), .Z(n7976) );
  AND U5079 ( .A(y[2]), .B(x[22]), .Z(n8020) );
  AND U5080 ( .A(y[12]), .B(x[12]), .Z(n8019) );
  XOR U5081 ( .A(n8020), .B(n8019), .Z(n8022) );
  AND U5082 ( .A(x[2]), .B(y[22]), .Z(n8021) );
  XOR U5083 ( .A(n8022), .B(n8021), .Z(n7975) );
  XOR U5084 ( .A(n7976), .B(n7975), .Z(n7977) );
  XNOR U5085 ( .A(n7978), .B(n7977), .Z(n8014) );
  NANDN U5086 ( .A(n7899), .B(n7898), .Z(n7903) );
  NAND U5087 ( .A(n7901), .B(n7900), .Z(n7902) );
  AND U5088 ( .A(n7903), .B(n7902), .Z(n7982) );
  AND U5089 ( .A(x[21]), .B(y[3]), .Z(n7989) );
  NAND U5090 ( .A(y[8]), .B(x[16]), .Z(n7990) );
  XNOR U5091 ( .A(n7989), .B(n7990), .Z(n7991) );
  NAND U5092 ( .A(x[5]), .B(y[19]), .Z(n7992) );
  XNOR U5093 ( .A(n7991), .B(n7992), .Z(n7979) );
  AND U5094 ( .A(x[20]), .B(y[4]), .Z(n7995) );
  NAND U5095 ( .A(x[6]), .B(y[18]), .Z(n7996) );
  XNOR U5096 ( .A(n7995), .B(n7996), .Z(n7997) );
  NAND U5097 ( .A(y[5]), .B(x[19]), .Z(n7998) );
  XOR U5098 ( .A(n7997), .B(n7998), .Z(n7980) );
  XNOR U5099 ( .A(n7979), .B(n7980), .Z(n7981) );
  XNOR U5100 ( .A(n7982), .B(n7981), .Z(n8009) );
  NANDN U5101 ( .A(n7905), .B(n7904), .Z(n7909) );
  NAND U5102 ( .A(n7907), .B(n7906), .Z(n7908) );
  NAND U5103 ( .A(n7909), .B(n7908), .Z(n8007) );
  NAND U5104 ( .A(n7911), .B(n7910), .Z(n7915) );
  NAND U5105 ( .A(n7913), .B(n7912), .Z(n7914) );
  AND U5106 ( .A(n7915), .B(n7914), .Z(n8008) );
  XNOR U5107 ( .A(n8007), .B(n8008), .Z(n8010) );
  XNOR U5108 ( .A(n8009), .B(n8010), .Z(n8013) );
  XOR U5109 ( .A(n8014), .B(n8013), .Z(n8015) );
  XOR U5110 ( .A(n8016), .B(n8015), .Z(n8075) );
  XOR U5111 ( .A(n8075), .B(n8074), .Z(n8076) );
  XOR U5112 ( .A(n8077), .B(n8076), .Z(n8082) );
  XOR U5113 ( .A(n8083), .B(n8082), .Z(n8093) );
  NAND U5114 ( .A(n7921), .B(n7920), .Z(n7925) );
  NAND U5115 ( .A(n7923), .B(n7922), .Z(n7924) );
  NAND U5116 ( .A(n7925), .B(n7924), .Z(n8088) );
  NAND U5117 ( .A(n7927), .B(n7926), .Z(n7931) );
  NAND U5118 ( .A(n7929), .B(n7928), .Z(n7930) );
  NAND U5119 ( .A(n7931), .B(n7930), .Z(n8086) );
  NAND U5120 ( .A(n7933), .B(n7932), .Z(n7937) );
  NAND U5121 ( .A(n7935), .B(n7934), .Z(n7936) );
  AND U5122 ( .A(n7937), .B(n7936), .Z(n8087) );
  XOR U5123 ( .A(n8086), .B(n8087), .Z(n8089) );
  XOR U5124 ( .A(n8088), .B(n8089), .Z(n8092) );
  NAND U5125 ( .A(n7939), .B(n7938), .Z(n7943) );
  NANDN U5126 ( .A(n7941), .B(n7940), .Z(n7942) );
  AND U5127 ( .A(n7943), .B(n7942), .Z(n8094) );
  XOR U5128 ( .A(n8095), .B(n8094), .Z(n7959) );
  XOR U5129 ( .A(n7960), .B(n7959), .Z(n7962) );
  NAND U5130 ( .A(n7948), .B(n7947), .Z(n7952) );
  NANDN U5131 ( .A(n7950), .B(n7949), .Z(n7951) );
  NAND U5132 ( .A(n7952), .B(n7951), .Z(n7953) );
  NANDN U5133 ( .A(n7954), .B(n7953), .Z(n7958) );
  XNOR U5134 ( .A(n7954), .B(n7953), .Z(n8917) );
  XNOR U5135 ( .A(n7956), .B(n7955), .Z(n8916) );
  NAND U5136 ( .A(n8917), .B(n8916), .Z(n7957) );
  NAND U5137 ( .A(n7958), .B(n7957), .Z(n7961) );
  XOR U5138 ( .A(n7962), .B(n7961), .Z(N57) );
  NANDN U5139 ( .A(n7964), .B(n7963), .Z(n7968) );
  NANDN U5140 ( .A(n7966), .B(n7965), .Z(n7967) );
  AND U5141 ( .A(n7968), .B(n7967), .Z(n8226) );
  NAND U5142 ( .A(n7970), .B(n7969), .Z(n7974) );
  NAND U5143 ( .A(n7972), .B(n7971), .Z(n7973) );
  NAND U5144 ( .A(n7974), .B(n7973), .Z(n8223) );
  NANDN U5145 ( .A(n7980), .B(n7979), .Z(n7984) );
  NANDN U5146 ( .A(n7982), .B(n7981), .Z(n7983) );
  NAND U5147 ( .A(n7984), .B(n7983), .Z(n8140) );
  XNOR U5148 ( .A(n8141), .B(n8140), .Z(n8143) );
  NANDN U5149 ( .A(n7990), .B(n7989), .Z(n7994) );
  NANDN U5150 ( .A(n7992), .B(n7991), .Z(n7993) );
  AND U5151 ( .A(n7994), .B(n7993), .Z(n8202) );
  AND U5152 ( .A(y[3]), .B(x[22]), .Z(n8164) );
  AND U5153 ( .A(y[8]), .B(x[17]), .Z(n8163) );
  NAND U5154 ( .A(x[5]), .B(y[20]), .Z(n8162) );
  XOR U5155 ( .A(n8163), .B(n8162), .Z(n8165) );
  XOR U5156 ( .A(n8164), .B(n8165), .Z(n8200) );
  AND U5157 ( .A(x[21]), .B(y[4]), .Z(n8181) );
  NAND U5158 ( .A(y[5]), .B(x[20]), .Z(n8182) );
  XNOR U5159 ( .A(n8181), .B(n8182), .Z(n8183) );
  NAND U5160 ( .A(x[19]), .B(y[6]), .Z(n8184) );
  XNOR U5161 ( .A(n8183), .B(n8184), .Z(n8199) );
  XNOR U5162 ( .A(n8200), .B(n8199), .Z(n8201) );
  XNOR U5163 ( .A(n8202), .B(n8201), .Z(n8135) );
  XOR U5164 ( .A(n8134), .B(n8135), .Z(n8137) );
  NANDN U5165 ( .A(n7996), .B(n7995), .Z(n8000) );
  NANDN U5166 ( .A(n7998), .B(n7997), .Z(n7999) );
  AND U5167 ( .A(n8000), .B(n7999), .Z(n8207) );
  AND U5168 ( .A(y[10]), .B(x[15]), .Z(n8189) );
  AND U5169 ( .A(x[6]), .B(y[19]), .Z(n8188) );
  NAND U5170 ( .A(y[7]), .B(x[18]), .Z(n8187) );
  XOR U5171 ( .A(n8188), .B(n8187), .Z(n8190) );
  XOR U5172 ( .A(n8189), .B(n8190), .Z(n8206) );
  AND U5173 ( .A(x[23]), .B(y[2]), .Z(n8170) );
  AND U5174 ( .A(x[16]), .B(y[9]), .Z(n8169) );
  NAND U5175 ( .A(y[21]), .B(x[4]), .Z(n8168) );
  XOR U5176 ( .A(n8169), .B(n8168), .Z(n8171) );
  XNOR U5177 ( .A(n8170), .B(n8171), .Z(n8205) );
  XOR U5178 ( .A(n8206), .B(n8205), .Z(n8208) );
  XOR U5179 ( .A(n8207), .B(n8208), .Z(n8136) );
  XOR U5180 ( .A(n8137), .B(n8136), .Z(n8142) );
  XOR U5181 ( .A(n8143), .B(n8142), .Z(n8101) );
  NAND U5182 ( .A(n8002), .B(n8001), .Z(n8006) );
  NANDN U5183 ( .A(n8004), .B(n8003), .Z(n8005) );
  NAND U5184 ( .A(n8006), .B(n8005), .Z(n8098) );
  NAND U5185 ( .A(n8008), .B(n8007), .Z(n8012) );
  NANDN U5186 ( .A(n8010), .B(n8009), .Z(n8011) );
  AND U5187 ( .A(n8012), .B(n8011), .Z(n8099) );
  XOR U5188 ( .A(n8098), .B(n8099), .Z(n8100) );
  XNOR U5189 ( .A(n8101), .B(n8100), .Z(n8224) );
  XOR U5190 ( .A(n8223), .B(n8224), .Z(n8225) );
  XOR U5191 ( .A(n8226), .B(n8225), .Z(n8232) );
  NAND U5192 ( .A(n8014), .B(n8013), .Z(n8018) );
  NANDN U5193 ( .A(n8016), .B(n8015), .Z(n8017) );
  AND U5194 ( .A(n8018), .B(n8017), .Z(n8217) );
  NAND U5195 ( .A(n8020), .B(n8019), .Z(n8024) );
  NAND U5196 ( .A(n8022), .B(n8021), .Z(n8023) );
  NAND U5197 ( .A(n8024), .B(n8023), .Z(n8105) );
  AND U5198 ( .A(n8026), .B(n8025), .Z(n8030) );
  NAND U5199 ( .A(n8028), .B(n8027), .Z(n8029) );
  NANDN U5200 ( .A(n8030), .B(n8029), .Z(n8104) );
  XOR U5201 ( .A(n8105), .B(n8104), .Z(n8106) );
  NAND U5202 ( .A(n8032), .B(n8031), .Z(n8036) );
  NAND U5203 ( .A(n8034), .B(n8033), .Z(n8035) );
  NAND U5204 ( .A(n8036), .B(n8035), .Z(n8124) );
  ANDN U5205 ( .B(o[24]), .A(n8037), .Z(n8119) );
  AND U5206 ( .A(x[25]), .B(y[0]), .Z(n8117) );
  NAND U5207 ( .A(y[25]), .B(x[0]), .Z(n8116) );
  XNOR U5208 ( .A(n8117), .B(n8116), .Z(n8118) );
  XOR U5209 ( .A(n8119), .B(n8118), .Z(n8123) );
  AND U5210 ( .A(x[8]), .B(y[17]), .Z(n8113) );
  AND U5211 ( .A(x[9]), .B(y[16]), .Z(n8111) );
  NAND U5212 ( .A(y[15]), .B(x[10]), .Z(n8110) );
  XNOR U5213 ( .A(n8111), .B(n8110), .Z(n8112) );
  XOR U5214 ( .A(n8113), .B(n8112), .Z(n8122) );
  XNOR U5215 ( .A(n8123), .B(n8122), .Z(n8125) );
  XOR U5216 ( .A(n8124), .B(n8125), .Z(n8107) );
  XNOR U5217 ( .A(n8106), .B(n8107), .Z(n8130) );
  NANDN U5218 ( .A(n8039), .B(n8038), .Z(n8043) );
  NANDN U5219 ( .A(n8041), .B(n8040), .Z(n8042) );
  AND U5220 ( .A(n8043), .B(n8042), .Z(n8129) );
  NAND U5221 ( .A(y[14]), .B(x[11]), .Z(n8177) );
  NAND U5222 ( .A(y[13]), .B(x[12]), .Z(n8176) );
  NAND U5223 ( .A(x[7]), .B(y[18]), .Z(n8175) );
  XNOR U5224 ( .A(n8176), .B(n8175), .Z(n8178) );
  XOR U5225 ( .A(n8177), .B(n8178), .Z(n8157) );
  NAND U5226 ( .A(x[13]), .B(y[12]), .Z(n8152) );
  AND U5227 ( .A(x[24]), .B(y[1]), .Z(n8174) );
  XOR U5228 ( .A(o[25]), .B(n8174), .Z(n8151) );
  NAND U5229 ( .A(x[1]), .B(y[24]), .Z(n8150) );
  XOR U5230 ( .A(n8151), .B(n8150), .Z(n8153) );
  XOR U5231 ( .A(n8152), .B(n8153), .Z(n8156) );
  XOR U5232 ( .A(n8157), .B(n8156), .Z(n8158) );
  NANDN U5233 ( .A(n8045), .B(n8044), .Z(n8049) );
  OR U5234 ( .A(n8047), .B(n8046), .Z(n8048) );
  NAND U5235 ( .A(n8049), .B(n8048), .Z(n8159) );
  XNOR U5236 ( .A(n8158), .B(n8159), .Z(n8128) );
  XOR U5237 ( .A(n8129), .B(n8128), .Z(n8131) );
  XOR U5238 ( .A(n8130), .B(n8131), .Z(n8213) );
  NANDN U5239 ( .A(n8051), .B(n8050), .Z(n8055) );
  NAND U5240 ( .A(n8053), .B(n8052), .Z(n8054) );
  AND U5241 ( .A(n8055), .B(n8054), .Z(n8196) );
  NANDN U5242 ( .A(n8057), .B(n8056), .Z(n8061) );
  NANDN U5243 ( .A(n8059), .B(n8058), .Z(n8060) );
  AND U5244 ( .A(n8061), .B(n8060), .Z(n8194) );
  AND U5245 ( .A(x[14]), .B(y[11]), .Z(n8144) );
  NAND U5246 ( .A(y[23]), .B(x[2]), .Z(n8145) );
  XNOR U5247 ( .A(n8144), .B(n8145), .Z(n8146) );
  NAND U5248 ( .A(x[3]), .B(y[22]), .Z(n8147) );
  XNOR U5249 ( .A(n8146), .B(n8147), .Z(n8193) );
  XNOR U5250 ( .A(n8194), .B(n8193), .Z(n8195) );
  XOR U5251 ( .A(n8196), .B(n8195), .Z(n8212) );
  NAND U5252 ( .A(n8063), .B(n8062), .Z(n8067) );
  NAND U5253 ( .A(n8065), .B(n8064), .Z(n8066) );
  NAND U5254 ( .A(n8067), .B(n8066), .Z(n8211) );
  XNOR U5255 ( .A(n8212), .B(n8211), .Z(n8214) );
  XOR U5256 ( .A(n8213), .B(n8214), .Z(n8218) );
  XNOR U5257 ( .A(n8217), .B(n8218), .Z(n8220) );
  NAND U5258 ( .A(n8069), .B(n8068), .Z(n8073) );
  NANDN U5259 ( .A(n8071), .B(n8070), .Z(n8072) );
  AND U5260 ( .A(n8073), .B(n8072), .Z(n8219) );
  XOR U5261 ( .A(n8220), .B(n8219), .Z(n8230) );
  NAND U5262 ( .A(n8075), .B(n8074), .Z(n8079) );
  NAND U5263 ( .A(n8077), .B(n8076), .Z(n8078) );
  AND U5264 ( .A(n8079), .B(n8078), .Z(n8229) );
  XNOR U5265 ( .A(n8230), .B(n8229), .Z(n8231) );
  XOR U5266 ( .A(n8232), .B(n8231), .Z(n8240) );
  NAND U5267 ( .A(n8081), .B(n8080), .Z(n8085) );
  NAND U5268 ( .A(n8083), .B(n8082), .Z(n8084) );
  NAND U5269 ( .A(n8085), .B(n8084), .Z(n8239) );
  XOR U5270 ( .A(n8240), .B(n8239), .Z(n8242) );
  NAND U5271 ( .A(n8087), .B(n8086), .Z(n8091) );
  NAND U5272 ( .A(n8089), .B(n8088), .Z(n8090) );
  AND U5273 ( .A(n8091), .B(n8090), .Z(n8241) );
  XOR U5274 ( .A(n8242), .B(n8241), .Z(n8235) );
  XOR U5275 ( .A(n8236), .B(n8235), .Z(n8238) );
  NANDN U5276 ( .A(n8093), .B(n8092), .Z(n8097) );
  NAND U5277 ( .A(n8095), .B(n8094), .Z(n8096) );
  AND U5278 ( .A(n8097), .B(n8096), .Z(n8237) );
  XNOR U5279 ( .A(n8238), .B(n8237), .Z(N58) );
  NAND U5280 ( .A(n8099), .B(n8098), .Z(n8103) );
  NANDN U5281 ( .A(n8101), .B(n8100), .Z(n8102) );
  AND U5282 ( .A(n8103), .B(n8102), .Z(n8544) );
  NAND U5283 ( .A(n8105), .B(n8104), .Z(n8109) );
  NANDN U5284 ( .A(n8107), .B(n8106), .Z(n8108) );
  AND U5285 ( .A(n8109), .B(n8108), .Z(n8248) );
  NAND U5286 ( .A(y[2]), .B(x[24]), .Z(n8330) );
  NAND U5287 ( .A(x[2]), .B(y[24]), .Z(n8329) );
  NAND U5288 ( .A(x[15]), .B(y[11]), .Z(n8328) );
  XNOR U5289 ( .A(n8329), .B(n8328), .Z(n8331) );
  XOR U5290 ( .A(n8330), .B(n8331), .Z(n8353) );
  NANDN U5291 ( .A(n8111), .B(n8110), .Z(n8115) );
  NANDN U5292 ( .A(n8113), .B(n8112), .Z(n8114) );
  AND U5293 ( .A(n8115), .B(n8114), .Z(n8352) );
  XOR U5294 ( .A(n8353), .B(n8352), .Z(n8354) );
  NANDN U5295 ( .A(n8117), .B(n8116), .Z(n8121) );
  NANDN U5296 ( .A(n8119), .B(n8118), .Z(n8120) );
  NAND U5297 ( .A(n8121), .B(n8120), .Z(n8355) );
  XOR U5298 ( .A(n8354), .B(n8355), .Z(n8245) );
  NAND U5299 ( .A(n8123), .B(n8122), .Z(n8127) );
  NANDN U5300 ( .A(n8125), .B(n8124), .Z(n8126) );
  AND U5301 ( .A(n8127), .B(n8126), .Z(n8246) );
  XOR U5302 ( .A(n8245), .B(n8246), .Z(n8247) );
  XOR U5303 ( .A(n8248), .B(n8247), .Z(n8293) );
  NANDN U5304 ( .A(n8129), .B(n8128), .Z(n8133) );
  NANDN U5305 ( .A(n8131), .B(n8130), .Z(n8132) );
  AND U5306 ( .A(n8133), .B(n8132), .Z(n8291) );
  NAND U5307 ( .A(n8135), .B(n8134), .Z(n8139) );
  NAND U5308 ( .A(n8137), .B(n8136), .Z(n8138) );
  NAND U5309 ( .A(n8139), .B(n8138), .Z(n8290) );
  XNOR U5310 ( .A(n8291), .B(n8290), .Z(n8292) );
  XNOR U5311 ( .A(n8293), .B(n8292), .Z(n8542) );
  AND U5312 ( .A(x[7]), .B(y[19]), .Z(n8252) );
  AND U5313 ( .A(x[6]), .B(y[20]), .Z(n8266) );
  AND U5314 ( .A(y[18]), .B(x[8]), .Z(n8265) );
  XOR U5315 ( .A(n8266), .B(n8265), .Z(n8268) );
  AND U5316 ( .A(x[9]), .B(y[17]), .Z(n8267) );
  XOR U5317 ( .A(n8268), .B(n8267), .Z(n8251) );
  XOR U5318 ( .A(n8252), .B(n8251), .Z(n8254) );
  AND U5319 ( .A(x[5]), .B(y[21]), .Z(n8365) );
  AND U5320 ( .A(y[14]), .B(x[12]), .Z(n8364) );
  XOR U5321 ( .A(n8365), .B(n8364), .Z(n8367) );
  AND U5322 ( .A(x[10]), .B(y[16]), .Z(n8366) );
  XOR U5323 ( .A(n8367), .B(n8366), .Z(n8253) );
  XOR U5324 ( .A(n8254), .B(n8253), .Z(n8337) );
  NANDN U5325 ( .A(n8145), .B(n8144), .Z(n8149) );
  NANDN U5326 ( .A(n8147), .B(n8146), .Z(n8148) );
  NAND U5327 ( .A(n8149), .B(n8148), .Z(n8334) );
  NANDN U5328 ( .A(n8151), .B(n8150), .Z(n8155) );
  NANDN U5329 ( .A(n8153), .B(n8152), .Z(n8154) );
  AND U5330 ( .A(n8155), .B(n8154), .Z(n8335) );
  XOR U5331 ( .A(n8334), .B(n8335), .Z(n8336) );
  XOR U5332 ( .A(n8337), .B(n8336), .Z(n8347) );
  NAND U5333 ( .A(n8157), .B(n8156), .Z(n8161) );
  NANDN U5334 ( .A(n8159), .B(n8158), .Z(n8160) );
  AND U5335 ( .A(n8161), .B(n8160), .Z(n8346) );
  XNOR U5336 ( .A(n8347), .B(n8346), .Z(n8349) );
  NANDN U5337 ( .A(n8163), .B(n8162), .Z(n8167) );
  OR U5338 ( .A(n8165), .B(n8164), .Z(n8166) );
  AND U5339 ( .A(n8167), .B(n8166), .Z(n8305) );
  NANDN U5340 ( .A(n8169), .B(n8168), .Z(n8173) );
  OR U5341 ( .A(n8171), .B(n8170), .Z(n8172) );
  AND U5342 ( .A(n8173), .B(n8172), .Z(n8304) );
  XOR U5343 ( .A(n8305), .B(n8304), .Z(n8307) );
  AND U5344 ( .A(x[14]), .B(y[12]), .Z(n8279) );
  AND U5345 ( .A(n8174), .B(o[25]), .Z(n8278) );
  XOR U5346 ( .A(n8279), .B(n8278), .Z(n8281) );
  AND U5347 ( .A(y[25]), .B(x[1]), .Z(n8280) );
  XOR U5348 ( .A(n8281), .B(n8280), .Z(n8359) );
  AND U5349 ( .A(x[25]), .B(y[1]), .Z(n8271) );
  XOR U5350 ( .A(o[26]), .B(n8271), .Z(n8371) );
  AND U5351 ( .A(y[0]), .B(x[26]), .Z(n8370) );
  XOR U5352 ( .A(n8371), .B(n8370), .Z(n8373) );
  AND U5353 ( .A(y[26]), .B(x[0]), .Z(n8372) );
  XOR U5354 ( .A(n8373), .B(n8372), .Z(n8358) );
  XOR U5355 ( .A(n8359), .B(n8358), .Z(n8361) );
  NAND U5356 ( .A(n8176), .B(n8175), .Z(n8180) );
  NANDN U5357 ( .A(n8178), .B(n8177), .Z(n8179) );
  AND U5358 ( .A(n8180), .B(n8179), .Z(n8360) );
  XOR U5359 ( .A(n8361), .B(n8360), .Z(n8306) );
  XOR U5360 ( .A(n8307), .B(n8306), .Z(n8379) );
  NANDN U5361 ( .A(n8182), .B(n8181), .Z(n8186) );
  NANDN U5362 ( .A(n8184), .B(n8183), .Z(n8185) );
  NAND U5363 ( .A(n8186), .B(n8185), .Z(n8342) );
  NAND U5364 ( .A(x[20]), .B(y[6]), .Z(n8274) );
  NAND U5365 ( .A(x[13]), .B(y[13]), .Z(n8273) );
  NAND U5366 ( .A(y[5]), .B(x[21]), .Z(n8272) );
  XOR U5367 ( .A(n8273), .B(n8272), .Z(n8275) );
  XOR U5368 ( .A(n8274), .B(n8275), .Z(n8341) );
  AND U5369 ( .A(x[23]), .B(y[3]), .Z(n8323) );
  AND U5370 ( .A(x[16]), .B(y[10]), .Z(n8322) );
  XOR U5371 ( .A(n8323), .B(n8322), .Z(n8325) );
  AND U5372 ( .A(y[4]), .B(x[22]), .Z(n8324) );
  XOR U5373 ( .A(n8325), .B(n8324), .Z(n8340) );
  XOR U5374 ( .A(n8342), .B(n8343), .Z(n8377) );
  AND U5375 ( .A(y[15]), .B(x[11]), .Z(n8258) );
  AND U5376 ( .A(x[3]), .B(y[23]), .Z(n8257) );
  XOR U5377 ( .A(n8258), .B(n8257), .Z(n8260) );
  AND U5378 ( .A(y[7]), .B(x[19]), .Z(n8259) );
  XOR U5379 ( .A(n8260), .B(n8259), .Z(n8311) );
  AND U5380 ( .A(x[4]), .B(y[22]), .Z(n8317) );
  AND U5381 ( .A(x[17]), .B(y[9]), .Z(n8316) );
  XOR U5382 ( .A(n8317), .B(n8316), .Z(n8319) );
  AND U5383 ( .A(y[8]), .B(x[18]), .Z(n8318) );
  XOR U5384 ( .A(n8319), .B(n8318), .Z(n8310) );
  XOR U5385 ( .A(n8311), .B(n8310), .Z(n8313) );
  NANDN U5386 ( .A(n8188), .B(n8187), .Z(n8192) );
  OR U5387 ( .A(n8190), .B(n8189), .Z(n8191) );
  AND U5388 ( .A(n8192), .B(n8191), .Z(n8312) );
  XNOR U5389 ( .A(n8313), .B(n8312), .Z(n8376) );
  XNOR U5390 ( .A(n8377), .B(n8376), .Z(n8378) );
  XNOR U5391 ( .A(n8379), .B(n8378), .Z(n8348) );
  XOR U5392 ( .A(n8349), .B(n8348), .Z(n8299) );
  NANDN U5393 ( .A(n8194), .B(n8193), .Z(n8198) );
  NANDN U5394 ( .A(n8196), .B(n8195), .Z(n8197) );
  NAND U5395 ( .A(n8198), .B(n8197), .Z(n8286) );
  NANDN U5396 ( .A(n8200), .B(n8199), .Z(n8204) );
  NANDN U5397 ( .A(n8202), .B(n8201), .Z(n8203) );
  NAND U5398 ( .A(n8204), .B(n8203), .Z(n8285) );
  NANDN U5399 ( .A(n8206), .B(n8205), .Z(n8210) );
  OR U5400 ( .A(n8208), .B(n8207), .Z(n8209) );
  NAND U5401 ( .A(n8210), .B(n8209), .Z(n8284) );
  XOR U5402 ( .A(n8285), .B(n8284), .Z(n8287) );
  XOR U5403 ( .A(n8286), .B(n8287), .Z(n8298) );
  XNOR U5404 ( .A(n8299), .B(n8298), .Z(n8300) );
  XNOR U5405 ( .A(n8301), .B(n8300), .Z(n8541) );
  XOR U5406 ( .A(n8542), .B(n8541), .Z(n8543) );
  XOR U5407 ( .A(n8544), .B(n8543), .Z(n8550) );
  NAND U5408 ( .A(n8212), .B(n8211), .Z(n8216) );
  NANDN U5409 ( .A(n8214), .B(n8213), .Z(n8215) );
  AND U5410 ( .A(n8216), .B(n8215), .Z(n8548) );
  NANDN U5411 ( .A(n8218), .B(n8217), .Z(n8222) );
  NAND U5412 ( .A(n8220), .B(n8219), .Z(n8221) );
  AND U5413 ( .A(n8222), .B(n8221), .Z(n8547) );
  XOR U5414 ( .A(n8548), .B(n8547), .Z(n8549) );
  XOR U5415 ( .A(n8550), .B(n8549), .Z(n8535) );
  NAND U5416 ( .A(n8224), .B(n8223), .Z(n8228) );
  NAND U5417 ( .A(n8226), .B(n8225), .Z(n8227) );
  AND U5418 ( .A(n8228), .B(n8227), .Z(n8534) );
  NANDN U5419 ( .A(n8230), .B(n8229), .Z(n8234) );
  NANDN U5420 ( .A(n8232), .B(n8231), .Z(n8233) );
  AND U5421 ( .A(n8234), .B(n8233), .Z(n8533) );
  XOR U5422 ( .A(n8534), .B(n8533), .Z(n8536) );
  XOR U5423 ( .A(n8535), .B(n8536), .Z(n8528) );
  XNOR U5424 ( .A(n8528), .B(n8527), .Z(n8530) );
  NAND U5425 ( .A(n8240), .B(n8239), .Z(n8244) );
  NAND U5426 ( .A(n8242), .B(n8241), .Z(n8243) );
  AND U5427 ( .A(n8244), .B(n8243), .Z(n8529) );
  XOR U5428 ( .A(n8530), .B(n8529), .Z(N59) );
  NAND U5429 ( .A(n8246), .B(n8245), .Z(n8250) );
  NAND U5430 ( .A(n8248), .B(n8247), .Z(n8249) );
  NAND U5431 ( .A(n8250), .B(n8249), .Z(n8406) );
  NAND U5432 ( .A(n8252), .B(n8251), .Z(n8256) );
  NAND U5433 ( .A(n8254), .B(n8253), .Z(n8255) );
  AND U5434 ( .A(n8256), .B(n8255), .Z(n8402) );
  NAND U5435 ( .A(n8258), .B(n8257), .Z(n8262) );
  NAND U5436 ( .A(n8260), .B(n8259), .Z(n8261) );
  NAND U5437 ( .A(n8262), .B(n8261), .Z(n8480) );
  NAND U5438 ( .A(y[5]), .B(x[22]), .Z(n8426) );
  NAND U5439 ( .A(x[23]), .B(y[4]), .Z(n8425) );
  NAND U5440 ( .A(x[8]), .B(y[19]), .Z(n8424) );
  XOR U5441 ( .A(n8425), .B(n8424), .Z(n8427) );
  XOR U5442 ( .A(n8426), .B(n8427), .Z(n8479) );
  AND U5443 ( .A(x[24]), .B(y[3]), .Z(n8264) );
  NAND U5444 ( .A(x[20]), .B(y[7]), .Z(n8263) );
  XNOR U5445 ( .A(n8264), .B(n8263), .Z(n8498) );
  AND U5446 ( .A(y[20]), .B(x[7]), .Z(n8497) );
  XOR U5447 ( .A(n8498), .B(n8497), .Z(n8478) );
  XNOR U5448 ( .A(n8479), .B(n8478), .Z(n8481) );
  XNOR U5449 ( .A(n8480), .B(n8481), .Z(n8400) );
  NAND U5450 ( .A(n8266), .B(n8265), .Z(n8270) );
  NAND U5451 ( .A(n8268), .B(n8267), .Z(n8269) );
  NAND U5452 ( .A(n8270), .B(n8269), .Z(n8474) );
  AND U5453 ( .A(x[14]), .B(y[13]), .Z(n8443) );
  AND U5454 ( .A(x[1]), .B(y[26]), .Z(n8442) );
  XOR U5455 ( .A(n8443), .B(n8442), .Z(n8445) );
  AND U5456 ( .A(n8271), .B(o[26]), .Z(n8444) );
  XOR U5457 ( .A(n8445), .B(n8444), .Z(n8473) );
  AND U5458 ( .A(y[10]), .B(x[17]), .Z(n8516) );
  AND U5459 ( .A(y[23]), .B(x[4]), .Z(n8515) );
  XOR U5460 ( .A(n8516), .B(n8515), .Z(n8518) );
  AND U5461 ( .A(x[5]), .B(y[22]), .Z(n8517) );
  XOR U5462 ( .A(n8518), .B(n8517), .Z(n8472) );
  XOR U5463 ( .A(n8473), .B(n8472), .Z(n8475) );
  XNOR U5464 ( .A(n8474), .B(n8475), .Z(n8492) );
  NAND U5465 ( .A(n8273), .B(n8272), .Z(n8277) );
  NAND U5466 ( .A(n8275), .B(n8274), .Z(n8276) );
  NAND U5467 ( .A(n8277), .B(n8276), .Z(n8490) );
  NAND U5468 ( .A(n8279), .B(n8278), .Z(n8283) );
  NAND U5469 ( .A(n8281), .B(n8280), .Z(n8282) );
  AND U5470 ( .A(n8283), .B(n8282), .Z(n8491) );
  XNOR U5471 ( .A(n8490), .B(n8491), .Z(n8493) );
  XOR U5472 ( .A(n8492), .B(n8493), .Z(n8401) );
  XOR U5473 ( .A(n8400), .B(n8401), .Z(n8403) );
  XNOR U5474 ( .A(n8402), .B(n8403), .Z(n8407) );
  XOR U5475 ( .A(n8406), .B(n8407), .Z(n8409) );
  NAND U5476 ( .A(n8285), .B(n8284), .Z(n8289) );
  NAND U5477 ( .A(n8287), .B(n8286), .Z(n8288) );
  AND U5478 ( .A(n8289), .B(n8288), .Z(n8408) );
  XOR U5479 ( .A(n8409), .B(n8408), .Z(n8296) );
  NANDN U5480 ( .A(n8291), .B(n8290), .Z(n8295) );
  NANDN U5481 ( .A(n8293), .B(n8292), .Z(n8294) );
  AND U5482 ( .A(n8295), .B(n8294), .Z(n8297) );
  XOR U5483 ( .A(n8297), .B(n8296), .Z(n8553) );
  NANDN U5484 ( .A(n8299), .B(n8298), .Z(n8303) );
  NANDN U5485 ( .A(n8301), .B(n8300), .Z(n8302) );
  AND U5486 ( .A(n8303), .B(n8302), .Z(n8385) );
  NAND U5487 ( .A(n8305), .B(n8304), .Z(n8309) );
  NAND U5488 ( .A(n8307), .B(n8306), .Z(n8308) );
  NAND U5489 ( .A(n8309), .B(n8308), .Z(n8414) );
  NAND U5490 ( .A(n8311), .B(n8310), .Z(n8315) );
  NAND U5491 ( .A(n8313), .B(n8312), .Z(n8314) );
  NAND U5492 ( .A(n8315), .B(n8314), .Z(n8412) );
  NAND U5493 ( .A(n8317), .B(n8316), .Z(n8321) );
  NAND U5494 ( .A(n8319), .B(n8318), .Z(n8320) );
  AND U5495 ( .A(n8321), .B(n8320), .Z(n8468) );
  AND U5496 ( .A(y[18]), .B(x[9]), .Z(n8633) );
  AND U5497 ( .A(x[21]), .B(y[6]), .Z(n8507) );
  XOR U5498 ( .A(n8633), .B(n8507), .Z(n8509) );
  AND U5499 ( .A(x[18]), .B(y[9]), .Z(n8508) );
  XOR U5500 ( .A(n8509), .B(n8508), .Z(n8467) );
  AND U5501 ( .A(y[1]), .B(x[26]), .Z(n8512) );
  XOR U5502 ( .A(o[27]), .B(n8512), .Z(n8524) );
  AND U5503 ( .A(y[27]), .B(x[0]), .Z(n8522) );
  AND U5504 ( .A(y[0]), .B(x[27]), .Z(n8521) );
  XOR U5505 ( .A(n8522), .B(n8521), .Z(n8523) );
  XNOR U5506 ( .A(n8524), .B(n8523), .Z(n8466) );
  XNOR U5507 ( .A(n8468), .B(n8469), .Z(n8463) );
  NAND U5508 ( .A(n8323), .B(n8322), .Z(n8327) );
  NAND U5509 ( .A(n8325), .B(n8324), .Z(n8326) );
  NAND U5510 ( .A(n8327), .B(n8326), .Z(n8460) );
  NAND U5511 ( .A(n8329), .B(n8328), .Z(n8333) );
  NANDN U5512 ( .A(n8331), .B(n8330), .Z(n8332) );
  AND U5513 ( .A(n8333), .B(n8332), .Z(n8461) );
  XOR U5514 ( .A(n8460), .B(n8461), .Z(n8462) );
  XNOR U5515 ( .A(n8463), .B(n8462), .Z(n8413) );
  XOR U5516 ( .A(n8412), .B(n8413), .Z(n8415) );
  XOR U5517 ( .A(n8414), .B(n8415), .Z(n8391) );
  NAND U5518 ( .A(n8335), .B(n8334), .Z(n8339) );
  NAND U5519 ( .A(n8337), .B(n8336), .Z(n8338) );
  AND U5520 ( .A(n8339), .B(n8338), .Z(n8389) );
  NANDN U5521 ( .A(n8341), .B(n8340), .Z(n8345) );
  NAND U5522 ( .A(n8343), .B(n8342), .Z(n8344) );
  AND U5523 ( .A(n8345), .B(n8344), .Z(n8388) );
  XOR U5524 ( .A(n8389), .B(n8388), .Z(n8390) );
  XOR U5525 ( .A(n8391), .B(n8390), .Z(n8383) );
  NANDN U5526 ( .A(n8347), .B(n8346), .Z(n8351) );
  NAND U5527 ( .A(n8349), .B(n8348), .Z(n8350) );
  AND U5528 ( .A(n8351), .B(n8350), .Z(n8397) );
  NAND U5529 ( .A(n8353), .B(n8352), .Z(n8357) );
  NANDN U5530 ( .A(n8355), .B(n8354), .Z(n8356) );
  NAND U5531 ( .A(n8357), .B(n8356), .Z(n8420) );
  NAND U5532 ( .A(n8359), .B(n8358), .Z(n8363) );
  NAND U5533 ( .A(n8361), .B(n8360), .Z(n8362) );
  NAND U5534 ( .A(n8363), .B(n8362), .Z(n8418) );
  AND U5535 ( .A(y[8]), .B(x[19]), .Z(n8502) );
  AND U5536 ( .A(x[25]), .B(y[2]), .Z(n8501) );
  XOR U5537 ( .A(n8502), .B(n8501), .Z(n8504) );
  AND U5538 ( .A(x[6]), .B(y[21]), .Z(n8503) );
  XOR U5539 ( .A(n8504), .B(n8503), .Z(n8485) );
  AND U5540 ( .A(y[12]), .B(x[15]), .Z(n8449) );
  AND U5541 ( .A(y[25]), .B(x[2]), .Z(n8448) );
  XOR U5542 ( .A(n8449), .B(n8448), .Z(n8451) );
  AND U5543 ( .A(x[3]), .B(y[24]), .Z(n8450) );
  XOR U5544 ( .A(n8451), .B(n8450), .Z(n8484) );
  XOR U5545 ( .A(n8485), .B(n8484), .Z(n8487) );
  AND U5546 ( .A(x[16]), .B(y[11]), .Z(n8431) );
  AND U5547 ( .A(x[10]), .B(y[17]), .Z(n8430) );
  XOR U5548 ( .A(n8431), .B(n8430), .Z(n8433) );
  AND U5549 ( .A(x[11]), .B(y[16]), .Z(n8432) );
  XOR U5550 ( .A(n8433), .B(n8432), .Z(n8439) );
  AND U5551 ( .A(x[13]), .B(y[14]), .Z(n8437) );
  AND U5552 ( .A(y[15]), .B(x[12]), .Z(n8436) );
  XOR U5553 ( .A(n8437), .B(n8436), .Z(n8438) );
  XOR U5554 ( .A(n8439), .B(n8438), .Z(n8486) );
  XOR U5555 ( .A(n8487), .B(n8486), .Z(n8456) );
  NAND U5556 ( .A(n8365), .B(n8364), .Z(n8369) );
  NAND U5557 ( .A(n8367), .B(n8366), .Z(n8368) );
  NAND U5558 ( .A(n8369), .B(n8368), .Z(n8455) );
  NAND U5559 ( .A(n8371), .B(n8370), .Z(n8375) );
  NAND U5560 ( .A(n8373), .B(n8372), .Z(n8374) );
  NAND U5561 ( .A(n8375), .B(n8374), .Z(n8454) );
  XNOR U5562 ( .A(n8455), .B(n8454), .Z(n8457) );
  XNOR U5563 ( .A(n8456), .B(n8457), .Z(n8419) );
  XOR U5564 ( .A(n8418), .B(n8419), .Z(n8421) );
  XOR U5565 ( .A(n8420), .B(n8421), .Z(n8395) );
  NANDN U5566 ( .A(n8377), .B(n8376), .Z(n8381) );
  NANDN U5567 ( .A(n8379), .B(n8378), .Z(n8380) );
  AND U5568 ( .A(n8381), .B(n8380), .Z(n8394) );
  XOR U5569 ( .A(n8395), .B(n8394), .Z(n8396) );
  XOR U5570 ( .A(n8397), .B(n8396), .Z(n8382) );
  XOR U5571 ( .A(n8383), .B(n8382), .Z(n8384) );
  XOR U5572 ( .A(n8385), .B(n8384), .Z(n8554) );
  NAND U5573 ( .A(n8383), .B(n8382), .Z(n8387) );
  NANDN U5574 ( .A(n8385), .B(n8384), .Z(n8386) );
  AND U5575 ( .A(n8387), .B(n8386), .Z(n8563) );
  XNOR U5576 ( .A(n8564), .B(n8563), .Z(n8566) );
  NAND U5577 ( .A(n8389), .B(n8388), .Z(n8393) );
  NANDN U5578 ( .A(n8391), .B(n8390), .Z(n8392) );
  AND U5579 ( .A(n8393), .B(n8392), .Z(n8717) );
  NAND U5580 ( .A(n8395), .B(n8394), .Z(n8399) );
  NAND U5581 ( .A(n8397), .B(n8396), .Z(n8398) );
  NAND U5582 ( .A(n8399), .B(n8398), .Z(n8715) );
  NANDN U5583 ( .A(n8401), .B(n8400), .Z(n8405) );
  NANDN U5584 ( .A(n8403), .B(n8402), .Z(n8404) );
  AND U5585 ( .A(n8405), .B(n8404), .Z(n8716) );
  XNOR U5586 ( .A(n8715), .B(n8716), .Z(n8718) );
  XNOR U5587 ( .A(n8717), .B(n8718), .Z(n8724) );
  NAND U5588 ( .A(n8407), .B(n8406), .Z(n8411) );
  NAND U5589 ( .A(n8409), .B(n8408), .Z(n8410) );
  NAND U5590 ( .A(n8411), .B(n8410), .Z(n8722) );
  NAND U5591 ( .A(n8413), .B(n8412), .Z(n8417) );
  NAND U5592 ( .A(n8415), .B(n8414), .Z(n8416) );
  NAND U5593 ( .A(n8417), .B(n8416), .Z(n8710) );
  NAND U5594 ( .A(n8419), .B(n8418), .Z(n8423) );
  NAND U5595 ( .A(n8421), .B(n8420), .Z(n8422) );
  NAND U5596 ( .A(n8423), .B(n8422), .Z(n8709) );
  XOR U5597 ( .A(n8710), .B(n8709), .Z(n8712) );
  AND U5598 ( .A(x[17]), .B(y[11]), .Z(n8622) );
  AND U5599 ( .A(y[6]), .B(x[22]), .Z(n8621) );
  XOR U5600 ( .A(n8622), .B(n8621), .Z(n8624) );
  AND U5601 ( .A(x[4]), .B(y[24]), .Z(n8623) );
  XOR U5602 ( .A(n8624), .B(n8623), .Z(n8651) );
  AND U5603 ( .A(y[10]), .B(x[18]), .Z(n8887) );
  AND U5604 ( .A(x[6]), .B(y[22]), .Z(n8841) );
  AND U5605 ( .A(x[19]), .B(y[9]), .Z(n8683) );
  XOR U5606 ( .A(n8841), .B(n8683), .Z(n8684) );
  XOR U5607 ( .A(n8887), .B(n8684), .Z(n8650) );
  XOR U5608 ( .A(n8651), .B(n8650), .Z(n8653) );
  NAND U5609 ( .A(n8425), .B(n8424), .Z(n8429) );
  NAND U5610 ( .A(n8427), .B(n8426), .Z(n8428) );
  AND U5611 ( .A(n8429), .B(n8428), .Z(n8652) );
  XOR U5612 ( .A(n8653), .B(n8652), .Z(n8585) );
  NAND U5613 ( .A(n8431), .B(n8430), .Z(n8435) );
  NAND U5614 ( .A(n8433), .B(n8432), .Z(n8434) );
  NAND U5615 ( .A(n8435), .B(n8434), .Z(n8705) );
  AND U5616 ( .A(y[17]), .B(x[11]), .Z(n8670) );
  AND U5617 ( .A(y[21]), .B(x[7]), .Z(n8668) );
  AND U5618 ( .A(y[16]), .B(x[12]), .Z(n8667) );
  XOR U5619 ( .A(n8668), .B(n8667), .Z(n8669) );
  XOR U5620 ( .A(n8670), .B(n8669), .Z(n8704) );
  AND U5621 ( .A(x[27]), .B(y[1]), .Z(n8875) );
  XOR U5622 ( .A(o[28]), .B(n8875), .Z(n8698) );
  AND U5623 ( .A(y[2]), .B(x[26]), .Z(n8697) );
  XOR U5624 ( .A(n8698), .B(n8697), .Z(n8700) );
  AND U5625 ( .A(y[13]), .B(x[15]), .Z(n8699) );
  XOR U5626 ( .A(n8700), .B(n8699), .Z(n8703) );
  XOR U5627 ( .A(n8704), .B(n8703), .Z(n8706) );
  XNOR U5628 ( .A(n8705), .B(n8706), .Z(n8586) );
  NAND U5629 ( .A(n8437), .B(n8436), .Z(n8441) );
  NAND U5630 ( .A(n8439), .B(n8438), .Z(n8440) );
  NAND U5631 ( .A(n8441), .B(n8440), .Z(n8646) );
  NAND U5632 ( .A(n8443), .B(n8442), .Z(n8447) );
  NAND U5633 ( .A(n8445), .B(n8444), .Z(n8446) );
  NAND U5634 ( .A(n8447), .B(n8446), .Z(n8645) );
  NAND U5635 ( .A(n8449), .B(n8448), .Z(n8453) );
  NAND U5636 ( .A(n8451), .B(n8450), .Z(n8452) );
  NAND U5637 ( .A(n8453), .B(n8452), .Z(n8644) );
  XNOR U5638 ( .A(n8645), .B(n8644), .Z(n8647) );
  XNOR U5639 ( .A(n8587), .B(n8588), .Z(n8618) );
  NAND U5640 ( .A(n8455), .B(n8454), .Z(n8459) );
  NANDN U5641 ( .A(n8457), .B(n8456), .Z(n8458) );
  AND U5642 ( .A(n8459), .B(n8458), .Z(n8616) );
  NAND U5643 ( .A(n8461), .B(n8460), .Z(n8465) );
  NANDN U5644 ( .A(n8463), .B(n8462), .Z(n8464) );
  AND U5645 ( .A(n8465), .B(n8464), .Z(n8612) );
  NANDN U5646 ( .A(n8467), .B(n8466), .Z(n8471) );
  NANDN U5647 ( .A(n8469), .B(n8468), .Z(n8470) );
  NAND U5648 ( .A(n8471), .B(n8470), .Z(n8609) );
  NAND U5649 ( .A(n8473), .B(n8472), .Z(n8477) );
  NAND U5650 ( .A(n8475), .B(n8474), .Z(n8476) );
  AND U5651 ( .A(n8477), .B(n8476), .Z(n8610) );
  XOR U5652 ( .A(n8609), .B(n8610), .Z(n8611) );
  XOR U5653 ( .A(n8612), .B(n8611), .Z(n8615) );
  XOR U5654 ( .A(n8616), .B(n8615), .Z(n8617) );
  NANDN U5655 ( .A(n8479), .B(n8478), .Z(n8483) );
  NAND U5656 ( .A(n8481), .B(n8480), .Z(n8482) );
  NAND U5657 ( .A(n8483), .B(n8482), .Z(n8574) );
  NAND U5658 ( .A(n8485), .B(n8484), .Z(n8489) );
  NAND U5659 ( .A(n8487), .B(n8486), .Z(n8488) );
  NAND U5660 ( .A(n8489), .B(n8488), .Z(n8573) );
  XOR U5661 ( .A(n8574), .B(n8573), .Z(n8576) );
  NAND U5662 ( .A(n8491), .B(n8490), .Z(n8495) );
  NANDN U5663 ( .A(n8493), .B(n8492), .Z(n8494) );
  AND U5664 ( .A(n8495), .B(n8494), .Z(n8575) );
  XOR U5665 ( .A(n8576), .B(n8575), .Z(n8567) );
  AND U5666 ( .A(y[7]), .B(x[24]), .Z(n9128) );
  NAND U5667 ( .A(n9128), .B(n8496), .Z(n8500) );
  NAND U5668 ( .A(n8498), .B(n8497), .Z(n8499) );
  NAND U5669 ( .A(n8500), .B(n8499), .Z(n8605) );
  AND U5670 ( .A(x[1]), .B(y[27]), .Z(n8664) );
  AND U5671 ( .A(x[14]), .B(y[14]), .Z(n8662) );
  AND U5672 ( .A(x[25]), .B(y[3]), .Z(n8836) );
  XOR U5673 ( .A(n8662), .B(n8836), .Z(n8663) );
  XOR U5674 ( .A(n8664), .B(n8663), .Z(n8604) );
  AND U5675 ( .A(y[26]), .B(x[2]), .Z(n8659) );
  AND U5676 ( .A(y[12]), .B(x[16]), .Z(n8657) );
  AND U5677 ( .A(x[24]), .B(y[4]), .Z(n8656) );
  XOR U5678 ( .A(n8657), .B(n8656), .Z(n8658) );
  XOR U5679 ( .A(n8659), .B(n8658), .Z(n8603) );
  XOR U5680 ( .A(n8604), .B(n8603), .Z(n8606) );
  XOR U5681 ( .A(n8605), .B(n8606), .Z(n8582) );
  NAND U5682 ( .A(n8502), .B(n8501), .Z(n8506) );
  NAND U5683 ( .A(n8504), .B(n8503), .Z(n8505) );
  NAND U5684 ( .A(n8506), .B(n8505), .Z(n8599) );
  AND U5685 ( .A(x[13]), .B(y[15]), .Z(n8694) );
  AND U5686 ( .A(y[25]), .B(x[3]), .Z(n8692) );
  AND U5687 ( .A(y[5]), .B(x[23]), .Z(n8691) );
  XOR U5688 ( .A(n8692), .B(n8691), .Z(n8693) );
  XOR U5689 ( .A(n8694), .B(n8693), .Z(n8598) );
  AND U5690 ( .A(x[5]), .B(y[23]), .Z(n8678) );
  AND U5691 ( .A(y[7]), .B(x[21]), .Z(n8677) );
  XOR U5692 ( .A(n8678), .B(n8677), .Z(n8680) );
  AND U5693 ( .A(x[20]), .B(y[8]), .Z(n8679) );
  XOR U5694 ( .A(n8680), .B(n8679), .Z(n8597) );
  XOR U5695 ( .A(n8598), .B(n8597), .Z(n8600) );
  XOR U5696 ( .A(n8599), .B(n8600), .Z(n8580) );
  AND U5697 ( .A(n8633), .B(n8507), .Z(n8511) );
  NAND U5698 ( .A(n8509), .B(n8508), .Z(n8510) );
  NANDN U5699 ( .A(n8511), .B(n8510), .Z(n8640) );
  NAND U5700 ( .A(n8512), .B(o[27]), .Z(n8628) );
  NAND U5701 ( .A(y[0]), .B(x[28]), .Z(n8627) );
  XOR U5702 ( .A(n8628), .B(n8627), .Z(n8630) );
  NAND U5703 ( .A(x[0]), .B(y[28]), .Z(n8629) );
  XOR U5704 ( .A(n8630), .B(n8629), .Z(n8639) );
  AND U5705 ( .A(y[20]), .B(x[8]), .Z(n8635) );
  AND U5706 ( .A(x[9]), .B(y[19]), .Z(n8514) );
  AND U5707 ( .A(x[10]), .B(y[18]), .Z(n8513) );
  XOR U5708 ( .A(n8514), .B(n8513), .Z(n8634) );
  XOR U5709 ( .A(n8635), .B(n8634), .Z(n8638) );
  XOR U5710 ( .A(n8640), .B(n8641), .Z(n8594) );
  NAND U5711 ( .A(n8516), .B(n8515), .Z(n8520) );
  NAND U5712 ( .A(n8518), .B(n8517), .Z(n8519) );
  AND U5713 ( .A(n8520), .B(n8519), .Z(n8592) );
  NAND U5714 ( .A(n8522), .B(n8521), .Z(n8526) );
  NAND U5715 ( .A(n8524), .B(n8523), .Z(n8525) );
  AND U5716 ( .A(n8526), .B(n8525), .Z(n8591) );
  XOR U5717 ( .A(n8592), .B(n8591), .Z(n8593) );
  XNOR U5718 ( .A(n8567), .B(n8568), .Z(n8569) );
  XNOR U5719 ( .A(n8570), .B(n8569), .Z(n8711) );
  XNOR U5720 ( .A(n8712), .B(n8711), .Z(n8721) );
  XOR U5721 ( .A(n8722), .B(n8721), .Z(n8723) );
  XNOR U5722 ( .A(n8724), .B(n8723), .Z(n8565) );
  XOR U5723 ( .A(n8566), .B(n8565), .Z(n8727) );
  NANDN U5724 ( .A(n8528), .B(n8527), .Z(n8532) );
  NAND U5725 ( .A(n8530), .B(n8529), .Z(n8531) );
  AND U5726 ( .A(n8532), .B(n8531), .Z(n8540) );
  NANDN U5727 ( .A(n8534), .B(n8533), .Z(n8538) );
  OR U5728 ( .A(n8536), .B(n8535), .Z(n8537) );
  AND U5729 ( .A(n8538), .B(n8537), .Z(n8539) );
  NANDN U5730 ( .A(n8540), .B(n8539), .Z(n8556) );
  XNOR U5731 ( .A(n8540), .B(n8539), .Z(n8919) );
  NAND U5732 ( .A(n8542), .B(n8541), .Z(n8546) );
  NAND U5733 ( .A(n8544), .B(n8543), .Z(n8545) );
  AND U5734 ( .A(n8546), .B(n8545), .Z(n8560) );
  NAND U5735 ( .A(n8548), .B(n8547), .Z(n8552) );
  NAND U5736 ( .A(n8550), .B(n8549), .Z(n8551) );
  AND U5737 ( .A(n8552), .B(n8551), .Z(n8557) );
  XNOR U5738 ( .A(n8554), .B(n8553), .Z(n8558) );
  XNOR U5739 ( .A(n8557), .B(n8558), .Z(n8559) );
  XNOR U5740 ( .A(n8560), .B(n8559), .Z(n8918) );
  NAND U5741 ( .A(n8919), .B(n8918), .Z(n8555) );
  NAND U5742 ( .A(n8556), .B(n8555), .Z(n8728) );
  XNOR U5743 ( .A(n8727), .B(n8728), .Z(n8730) );
  NANDN U5744 ( .A(n8558), .B(n8557), .Z(n8562) );
  NAND U5745 ( .A(n8560), .B(n8559), .Z(n8561) );
  NAND U5746 ( .A(n8562), .B(n8561), .Z(n8729) );
  XNOR U5747 ( .A(n8730), .B(n8729), .Z(N61) );
  NANDN U5748 ( .A(n8568), .B(n8567), .Z(n8572) );
  NANDN U5749 ( .A(n8570), .B(n8569), .Z(n8571) );
  AND U5750 ( .A(n8572), .B(n8571), .Z(n8745) );
  NAND U5751 ( .A(n8574), .B(n8573), .Z(n8578) );
  NAND U5752 ( .A(n8576), .B(n8575), .Z(n8577) );
  NAND U5753 ( .A(n8578), .B(n8577), .Z(n8755) );
  NANDN U5754 ( .A(n8580), .B(n8579), .Z(n8584) );
  NANDN U5755 ( .A(n8582), .B(n8581), .Z(n8583) );
  AND U5756 ( .A(n8584), .B(n8583), .Z(n8756) );
  XOR U5757 ( .A(n8755), .B(n8756), .Z(n8758) );
  NANDN U5758 ( .A(n8586), .B(n8585), .Z(n8590) );
  NANDN U5759 ( .A(n8588), .B(n8587), .Z(n8589) );
  NAND U5760 ( .A(n8590), .B(n8589), .Z(n8749) );
  NAND U5761 ( .A(n8592), .B(n8591), .Z(n8596) );
  NANDN U5762 ( .A(n8594), .B(n8593), .Z(n8595) );
  AND U5763 ( .A(n8596), .B(n8595), .Z(n8811) );
  NAND U5764 ( .A(n8598), .B(n8597), .Z(n8602) );
  NAND U5765 ( .A(n8600), .B(n8599), .Z(n8601) );
  NAND U5766 ( .A(n8602), .B(n8601), .Z(n8810) );
  NAND U5767 ( .A(n8604), .B(n8603), .Z(n8608) );
  NAND U5768 ( .A(n8606), .B(n8605), .Z(n8607) );
  NAND U5769 ( .A(n8608), .B(n8607), .Z(n8809) );
  XNOR U5770 ( .A(n8810), .B(n8809), .Z(n8812) );
  XOR U5771 ( .A(n8749), .B(n8750), .Z(n8752) );
  NAND U5772 ( .A(n8610), .B(n8609), .Z(n8614) );
  NAND U5773 ( .A(n8612), .B(n8611), .Z(n8613) );
  AND U5774 ( .A(n8614), .B(n8613), .Z(n8751) );
  XOR U5775 ( .A(n8752), .B(n8751), .Z(n8757) );
  XOR U5776 ( .A(n8758), .B(n8757), .Z(n8764) );
  NAND U5777 ( .A(n8616), .B(n8615), .Z(n8620) );
  NANDN U5778 ( .A(n8618), .B(n8617), .Z(n8619) );
  AND U5779 ( .A(n8620), .B(n8619), .Z(n8762) );
  NAND U5780 ( .A(n8622), .B(n8621), .Z(n8626) );
  NAND U5781 ( .A(n8624), .B(n8623), .Z(n8625) );
  NAND U5782 ( .A(n8626), .B(n8625), .Z(n8797) );
  NAND U5783 ( .A(n8628), .B(n8627), .Z(n8632) );
  NAND U5784 ( .A(n8630), .B(n8629), .Z(n8631) );
  AND U5785 ( .A(n8632), .B(n8631), .Z(n8798) );
  XOR U5786 ( .A(n8797), .B(n8798), .Z(n8799) );
  AND U5787 ( .A(y[19]), .B(x[10]), .Z(n8882) );
  NAND U5788 ( .A(n8633), .B(n8882), .Z(n8637) );
  NAND U5789 ( .A(n8635), .B(n8634), .Z(n8636) );
  NAND U5790 ( .A(n8637), .B(n8636), .Z(n8775) );
  AND U5791 ( .A(y[14]), .B(x[15]), .Z(n8831) );
  AND U5792 ( .A(x[21]), .B(y[8]), .Z(n8830) );
  XOR U5793 ( .A(n8831), .B(n8830), .Z(n8833) );
  AND U5794 ( .A(x[20]), .B(y[9]), .Z(n8832) );
  XOR U5795 ( .A(n8833), .B(n8832), .Z(n8774) );
  AND U5796 ( .A(y[17]), .B(x[12]), .Z(n8822) );
  AND U5797 ( .A(x[1]), .B(y[28]), .Z(n8821) );
  XOR U5798 ( .A(n8822), .B(n8821), .Z(n8824) );
  AND U5799 ( .A(y[7]), .B(x[22]), .Z(n8823) );
  XOR U5800 ( .A(n8824), .B(n8823), .Z(n8773) );
  XOR U5801 ( .A(n8774), .B(n8773), .Z(n8776) );
  XNOR U5802 ( .A(n8775), .B(n8776), .Z(n8800) );
  NANDN U5803 ( .A(n8639), .B(n8638), .Z(n8643) );
  NAND U5804 ( .A(n8641), .B(n8640), .Z(n8642) );
  AND U5805 ( .A(n8643), .B(n8642), .Z(n8803) );
  NAND U5806 ( .A(n8645), .B(n8644), .Z(n8649) );
  NANDN U5807 ( .A(n8647), .B(n8646), .Z(n8648) );
  AND U5808 ( .A(n8649), .B(n8648), .Z(n8805) );
  XOR U5809 ( .A(n8806), .B(n8805), .Z(n8901) );
  NAND U5810 ( .A(n8651), .B(n8650), .Z(n8655) );
  NAND U5811 ( .A(n8653), .B(n8652), .Z(n8654) );
  NAND U5812 ( .A(n8655), .B(n8654), .Z(n8898) );
  NAND U5813 ( .A(n8657), .B(n8656), .Z(n8661) );
  NAND U5814 ( .A(n8659), .B(n8658), .Z(n8660) );
  NAND U5815 ( .A(n8661), .B(n8660), .Z(n8768) );
  NAND U5816 ( .A(n8662), .B(n8836), .Z(n8666) );
  NAND U5817 ( .A(n8664), .B(n8663), .Z(n8665) );
  NAND U5818 ( .A(n8666), .B(n8665), .Z(n8767) );
  XOR U5819 ( .A(n8768), .B(n8767), .Z(n8769) );
  NAND U5820 ( .A(n8668), .B(n8667), .Z(n8672) );
  NAND U5821 ( .A(n8670), .B(n8669), .Z(n8671) );
  NAND U5822 ( .A(n8672), .B(n8671), .Z(n8865) );
  AND U5823 ( .A(x[3]), .B(y[26]), .Z(n8852) );
  AND U5824 ( .A(y[12]), .B(x[17]), .Z(n8851) );
  XOR U5825 ( .A(n8852), .B(n8851), .Z(n8854) );
  AND U5826 ( .A(y[18]), .B(x[11]), .Z(n8853) );
  XOR U5827 ( .A(n8854), .B(n8853), .Z(n8864) );
  AND U5828 ( .A(x[13]), .B(y[16]), .Z(n8847) );
  AND U5829 ( .A(y[5]), .B(x[24]), .Z(n8846) );
  XOR U5830 ( .A(n8847), .B(n8846), .Z(n8848) );
  AND U5831 ( .A(x[23]), .B(y[6]), .Z(n9036) );
  XOR U5832 ( .A(n8848), .B(n9036), .Z(n8863) );
  XOR U5833 ( .A(n8864), .B(n8863), .Z(n8866) );
  XNOR U5834 ( .A(n8865), .B(n8866), .Z(n8770) );
  AND U5835 ( .A(y[11]), .B(x[18]), .Z(n8674) );
  NAND U5836 ( .A(y[10]), .B(x[19]), .Z(n8673) );
  XNOR U5837 ( .A(n8674), .B(n8673), .Z(n8889) );
  AND U5838 ( .A(y[27]), .B(x[2]), .Z(n8888) );
  XOR U5839 ( .A(n8889), .B(n8888), .Z(n8858) );
  NAND U5840 ( .A(o[28]), .B(y[1]), .Z(n8675) );
  XNOR U5841 ( .A(y[2]), .B(n8675), .Z(n8676) );
  AND U5842 ( .A(x[27]), .B(n8676), .Z(n8878) );
  AND U5843 ( .A(x[16]), .B(y[13]), .Z(n8877) );
  XOR U5844 ( .A(n8878), .B(n8877), .Z(n8857) );
  XOR U5845 ( .A(n8858), .B(n8857), .Z(n8860) );
  NAND U5846 ( .A(n8678), .B(n8677), .Z(n8682) );
  NAND U5847 ( .A(n8680), .B(n8679), .Z(n8681) );
  NAND U5848 ( .A(n8682), .B(n8681), .Z(n8859) );
  XOR U5849 ( .A(n8860), .B(n8859), .Z(n8893) );
  NAND U5850 ( .A(n8841), .B(n8683), .Z(n8686) );
  NAND U5851 ( .A(n8887), .B(n8684), .Z(n8685) );
  NAND U5852 ( .A(n8686), .B(n8685), .Z(n8781) );
  AND U5853 ( .A(y[1]), .B(x[28]), .Z(n8829) );
  XOR U5854 ( .A(o[29]), .B(n8829), .Z(n8794) );
  AND U5855 ( .A(x[0]), .B(y[29]), .Z(n8792) );
  AND U5856 ( .A(y[0]), .B(x[29]), .Z(n8791) );
  XOR U5857 ( .A(n8792), .B(n8791), .Z(n8793) );
  XOR U5858 ( .A(n8794), .B(n8793), .Z(n8780) );
  AND U5859 ( .A(y[15]), .B(x[14]), .Z(n8838) );
  AND U5860 ( .A(x[26]), .B(y[3]), .Z(n8688) );
  AND U5861 ( .A(y[4]), .B(x[25]), .Z(n8687) );
  XOR U5862 ( .A(n8688), .B(n8687), .Z(n8837) );
  XOR U5863 ( .A(n8838), .B(n8837), .Z(n8779) );
  XOR U5864 ( .A(n8780), .B(n8779), .Z(n8782) );
  XNOR U5865 ( .A(n8781), .B(n8782), .Z(n8892) );
  NAND U5866 ( .A(y[20]), .B(x[9]), .Z(n8787) );
  AND U5867 ( .A(y[22]), .B(x[7]), .Z(n8690) );
  NAND U5868 ( .A(x[6]), .B(y[23]), .Z(n8689) );
  XNOR U5869 ( .A(n8690), .B(n8689), .Z(n8843) );
  AND U5870 ( .A(y[21]), .B(x[8]), .Z(n8842) );
  XOR U5871 ( .A(n8843), .B(n8842), .Z(n8786) );
  AND U5872 ( .A(x[5]), .B(y[24]), .Z(n8884) );
  AND U5873 ( .A(y[25]), .B(x[4]), .Z(n8881) );
  XOR U5874 ( .A(n8882), .B(n8881), .Z(n8883) );
  XNOR U5875 ( .A(n8884), .B(n8883), .Z(n8785) );
  XOR U5876 ( .A(n8787), .B(n8788), .Z(n8872) );
  NAND U5877 ( .A(n8692), .B(n8691), .Z(n8696) );
  NAND U5878 ( .A(n8694), .B(n8693), .Z(n8695) );
  AND U5879 ( .A(n8696), .B(n8695), .Z(n8870) );
  NAND U5880 ( .A(n8698), .B(n8697), .Z(n8702) );
  NAND U5881 ( .A(n8700), .B(n8699), .Z(n8701) );
  AND U5882 ( .A(n8702), .B(n8701), .Z(n8869) );
  XOR U5883 ( .A(n8870), .B(n8869), .Z(n8871) );
  XOR U5884 ( .A(n8872), .B(n8871), .Z(n8816) );
  NAND U5885 ( .A(n8704), .B(n8703), .Z(n8708) );
  NAND U5886 ( .A(n8706), .B(n8705), .Z(n8707) );
  NAND U5887 ( .A(n8708), .B(n8707), .Z(n8815) );
  XOR U5888 ( .A(n8898), .B(n8899), .Z(n8900) );
  XOR U5889 ( .A(n8762), .B(n8761), .Z(n8763) );
  XOR U5890 ( .A(n8764), .B(n8763), .Z(n8744) );
  NAND U5891 ( .A(n8710), .B(n8709), .Z(n8714) );
  NAND U5892 ( .A(n8712), .B(n8711), .Z(n8713) );
  AND U5893 ( .A(n8714), .B(n8713), .Z(n8743) );
  XNOR U5894 ( .A(n8745), .B(n8746), .Z(n8740) );
  NAND U5895 ( .A(n8716), .B(n8715), .Z(n8720) );
  NANDN U5896 ( .A(n8718), .B(n8717), .Z(n8719) );
  NAND U5897 ( .A(n8720), .B(n8719), .Z(n8737) );
  NAND U5898 ( .A(n8722), .B(n8721), .Z(n8726) );
  NANDN U5899 ( .A(n8724), .B(n8723), .Z(n8725) );
  AND U5900 ( .A(n8726), .B(n8725), .Z(n8738) );
  XOR U5901 ( .A(n8737), .B(n8738), .Z(n8739) );
  XOR U5902 ( .A(n8734), .B(n8733), .Z(n8736) );
  NANDN U5903 ( .A(n8728), .B(n8727), .Z(n8732) );
  NAND U5904 ( .A(n8730), .B(n8729), .Z(n8731) );
  AND U5905 ( .A(n8732), .B(n8731), .Z(n8735) );
  XOR U5906 ( .A(n8736), .B(n8735), .Z(N62) );
  NAND U5907 ( .A(n8738), .B(n8737), .Z(n8742) );
  NANDN U5908 ( .A(n8740), .B(n8739), .Z(n8741) );
  NAND U5909 ( .A(n8742), .B(n8741), .Z(n8923) );
  NANDN U5910 ( .A(n8744), .B(n8743), .Z(n8748) );
  NANDN U5911 ( .A(n8746), .B(n8745), .Z(n8747) );
  NAND U5912 ( .A(n8748), .B(n8747), .Z(n9209) );
  NAND U5913 ( .A(n8750), .B(n8749), .Z(n8754) );
  NAND U5914 ( .A(n8752), .B(n8751), .Z(n8753) );
  AND U5915 ( .A(n8754), .B(n8753), .Z(n9192) );
  NAND U5916 ( .A(n8756), .B(n8755), .Z(n8760) );
  NAND U5917 ( .A(n8758), .B(n8757), .Z(n8759) );
  AND U5918 ( .A(n8760), .B(n8759), .Z(n9194) );
  NAND U5919 ( .A(n8762), .B(n8761), .Z(n8766) );
  NAND U5920 ( .A(n8764), .B(n8763), .Z(n8765) );
  AND U5921 ( .A(n8766), .B(n8765), .Z(n9193) );
  XOR U5922 ( .A(n9194), .B(n9193), .Z(n9191) );
  XOR U5923 ( .A(n9192), .B(n9191), .Z(n9211) );
  NAND U5924 ( .A(n8768), .B(n8767), .Z(n8772) );
  NANDN U5925 ( .A(n8770), .B(n8769), .Z(n8771) );
  AND U5926 ( .A(n8772), .B(n8771), .Z(n9170) );
  NAND U5927 ( .A(n8774), .B(n8773), .Z(n8778) );
  NAND U5928 ( .A(n8776), .B(n8775), .Z(n8777) );
  AND U5929 ( .A(n8778), .B(n8777), .Z(n9169) );
  XOR U5930 ( .A(n9170), .B(n9169), .Z(n9172) );
  NAND U5931 ( .A(n8780), .B(n8779), .Z(n8784) );
  NAND U5932 ( .A(n8782), .B(n8781), .Z(n8783) );
  AND U5933 ( .A(n8784), .B(n8783), .Z(n9171) );
  XOR U5934 ( .A(n9172), .B(n9171), .Z(n8946) );
  NANDN U5935 ( .A(n8786), .B(n8785), .Z(n8790) );
  NAND U5936 ( .A(n8788), .B(n8787), .Z(n8789) );
  NAND U5937 ( .A(n8790), .B(n8789), .Z(n8935) );
  AND U5938 ( .A(y[3]), .B(x[27]), .Z(n9054) );
  AND U5939 ( .A(x[1]), .B(y[29]), .Z(n9053) );
  XOR U5940 ( .A(n9054), .B(n9053), .Z(n9051) );
  XOR U5941 ( .A(n9052), .B(n9051), .Z(n8983) );
  AND U5942 ( .A(y[18]), .B(x[12]), .Z(n9021) );
  AND U5943 ( .A(y[19]), .B(x[11]), .Z(n9023) );
  AND U5944 ( .A(x[13]), .B(y[17]), .Z(n9022) );
  XOR U5945 ( .A(n9023), .B(n9022), .Z(n9020) );
  XOR U5946 ( .A(n9021), .B(n9020), .Z(n9007) );
  AND U5947 ( .A(y[21]), .B(x[9]), .Z(n9009) );
  AND U5948 ( .A(y[20]), .B(x[10]), .Z(n9008) );
  XOR U5949 ( .A(n9009), .B(n9008), .Z(n9006) );
  XOR U5950 ( .A(n9007), .B(n9006), .Z(n8982) );
  XOR U5951 ( .A(n8983), .B(n8982), .Z(n8981) );
  NAND U5952 ( .A(n8792), .B(n8791), .Z(n8796) );
  NAND U5953 ( .A(n8794), .B(n8793), .Z(n8795) );
  NAND U5954 ( .A(n8796), .B(n8795), .Z(n8980) );
  XNOR U5955 ( .A(n8981), .B(n8980), .Z(n8934) );
  XOR U5956 ( .A(n8935), .B(n8934), .Z(n8933) );
  NAND U5957 ( .A(n8798), .B(n8797), .Z(n8802) );
  NANDN U5958 ( .A(n8800), .B(n8799), .Z(n8801) );
  AND U5959 ( .A(n8802), .B(n8801), .Z(n8932) );
  XNOR U5960 ( .A(n8933), .B(n8932), .Z(n8947) );
  NANDN U5961 ( .A(n8804), .B(n8803), .Z(n8808) );
  NAND U5962 ( .A(n8806), .B(n8805), .Z(n8807) );
  AND U5963 ( .A(n8808), .B(n8807), .Z(n8948) );
  XNOR U5964 ( .A(n8949), .B(n8948), .Z(n9215) );
  NAND U5965 ( .A(n8810), .B(n8809), .Z(n8814) );
  NANDN U5966 ( .A(n8812), .B(n8811), .Z(n8813) );
  NAND U5967 ( .A(n8814), .B(n8813), .Z(n8929) );
  NANDN U5968 ( .A(n8816), .B(n8815), .Z(n8820) );
  NANDN U5969 ( .A(n8818), .B(n8817), .Z(n8819) );
  AND U5970 ( .A(n8820), .B(n8819), .Z(n9199) );
  NAND U5971 ( .A(n8822), .B(n8821), .Z(n8826) );
  NAND U5972 ( .A(n8824), .B(n8823), .Z(n8825) );
  AND U5973 ( .A(n8826), .B(n8825), .Z(n8975) );
  AND U5974 ( .A(y[5]), .B(x[25]), .Z(n9035) );
  AND U5975 ( .A(y[6]), .B(x[24]), .Z(n8828) );
  AND U5976 ( .A(y[7]), .B(x[23]), .Z(n8827) );
  XOR U5977 ( .A(n8828), .B(n8827), .Z(n9034) );
  XOR U5978 ( .A(n9035), .B(n9034), .Z(n8995) );
  AND U5979 ( .A(n8829), .B(o[29]), .Z(n9027) );
  AND U5980 ( .A(y[2]), .B(x[28]), .Z(n9029) );
  AND U5981 ( .A(y[14]), .B(x[16]), .Z(n9028) );
  XOR U5982 ( .A(n9029), .B(n9028), .Z(n9026) );
  XNOR U5983 ( .A(n9027), .B(n9026), .Z(n8994) );
  NAND U5984 ( .A(n8831), .B(n8830), .Z(n8835) );
  NAND U5985 ( .A(n8833), .B(n8832), .Z(n8834) );
  AND U5986 ( .A(n8835), .B(n8834), .Z(n8992) );
  XOR U5987 ( .A(n8993), .B(n8992), .Z(n8974) );
  XOR U5988 ( .A(n8975), .B(n8974), .Z(n8973) );
  AND U5989 ( .A(y[4]), .B(x[26]), .Z(n9048) );
  NAND U5990 ( .A(n8836), .B(n9048), .Z(n8840) );
  NAND U5991 ( .A(n8838), .B(n8837), .Z(n8839) );
  AND U5992 ( .A(n8840), .B(n8839), .Z(n8972) );
  XOR U5993 ( .A(n8973), .B(n8972), .Z(n8953) );
  AND U5994 ( .A(y[23]), .B(x[7]), .Z(n9146) );
  AND U5995 ( .A(y[8]), .B(x[22]), .Z(n9148) );
  AND U5996 ( .A(x[21]), .B(y[9]), .Z(n9147) );
  XOR U5997 ( .A(n9148), .B(n9147), .Z(n9145) );
  XOR U5998 ( .A(n9146), .B(n9145), .Z(n9001) );
  AND U5999 ( .A(x[2]), .B(y[28]), .Z(n9047) );
  XOR U6000 ( .A(n9048), .B(n9047), .Z(n9046) );
  AND U6001 ( .A(x[17]), .B(y[13]), .Z(n9045) );
  XOR U6002 ( .A(n9046), .B(n9045), .Z(n9003) );
  NAND U6003 ( .A(n8841), .B(n9146), .Z(n8845) );
  NAND U6004 ( .A(n8843), .B(n8842), .Z(n8844) );
  NAND U6005 ( .A(n8845), .B(n8844), .Z(n9002) );
  XOR U6006 ( .A(n9003), .B(n9002), .Z(n9000) );
  XOR U6007 ( .A(n9001), .B(n9000), .Z(n9176) );
  NAND U6008 ( .A(n8847), .B(n8846), .Z(n8850) );
  NAND U6009 ( .A(n8848), .B(n9036), .Z(n8849) );
  AND U6010 ( .A(n8850), .B(n8849), .Z(n9175) );
  AND U6011 ( .A(x[0]), .B(y[30]), .Z(n9013) );
  AND U6012 ( .A(y[1]), .B(x[29]), .Z(n9121) );
  XOR U6013 ( .A(o[30]), .B(n9121), .Z(n9015) );
  AND U6014 ( .A(y[0]), .B(x[30]), .Z(n9014) );
  XOR U6015 ( .A(n9015), .B(n9014), .Z(n9012) );
  XOR U6016 ( .A(n9013), .B(n9012), .Z(n8963) );
  AND U6017 ( .A(x[14]), .B(y[16]), .Z(n9142) );
  AND U6018 ( .A(x[20]), .B(y[10]), .Z(n9141) );
  XOR U6019 ( .A(n9142), .B(n9141), .Z(n9140) );
  AND U6020 ( .A(y[22]), .B(x[8]), .Z(n9139) );
  XNOR U6021 ( .A(n9140), .B(n9139), .Z(n8962) );
  NAND U6022 ( .A(n8852), .B(n8851), .Z(n8856) );
  NAND U6023 ( .A(n8854), .B(n8853), .Z(n8855) );
  AND U6024 ( .A(n8856), .B(n8855), .Z(n8960) );
  XOR U6025 ( .A(n8961), .B(n8960), .Z(n9177) );
  XNOR U6026 ( .A(n9178), .B(n9177), .Z(n8952) );
  NAND U6027 ( .A(n8858), .B(n8857), .Z(n8862) );
  NAND U6028 ( .A(n8860), .B(n8859), .Z(n8861) );
  NAND U6029 ( .A(n8862), .B(n8861), .Z(n8954) );
  XOR U6030 ( .A(n8955), .B(n8954), .Z(n9200) );
  NAND U6031 ( .A(n8864), .B(n8863), .Z(n8868) );
  NAND U6032 ( .A(n8866), .B(n8865), .Z(n8867) );
  NAND U6033 ( .A(n8868), .B(n8867), .Z(n8940) );
  NAND U6034 ( .A(n8870), .B(n8869), .Z(n8874) );
  NAND U6035 ( .A(n8872), .B(n8871), .Z(n8873) );
  AND U6036 ( .A(n8874), .B(n8873), .Z(n8941) );
  XOR U6037 ( .A(n8940), .B(n8941), .Z(n8939) );
  AND U6038 ( .A(n8875), .B(o[28]), .Z(n8876) );
  NAND U6039 ( .A(y[2]), .B(n8876), .Z(n8880) );
  NAND U6040 ( .A(n8878), .B(n8877), .Z(n8879) );
  NAND U6041 ( .A(n8880), .B(n8879), .Z(n8966) );
  AND U6042 ( .A(n8882), .B(n8881), .Z(n8886) );
  NAND U6043 ( .A(n8884), .B(n8883), .Z(n8885) );
  NANDN U6044 ( .A(n8886), .B(n8885), .Z(n8968) );
  AND U6045 ( .A(x[19]), .B(y[11]), .Z(n9042) );
  NAND U6046 ( .A(n8887), .B(n9042), .Z(n8891) );
  NAND U6047 ( .A(n8889), .B(n8888), .Z(n8890) );
  NAND U6048 ( .A(n8891), .B(n8890), .Z(n8986) );
  AND U6049 ( .A(y[26]), .B(x[4]), .Z(n9058) );
  AND U6050 ( .A(x[3]), .B(y[27]), .Z(n9060) );
  AND U6051 ( .A(y[12]), .B(x[18]), .Z(n9059) );
  XOR U6052 ( .A(n9060), .B(n9059), .Z(n9057) );
  XOR U6053 ( .A(n9058), .B(n9057), .Z(n8989) );
  AND U6054 ( .A(y[25]), .B(x[5]), .Z(n9041) );
  XOR U6055 ( .A(n9042), .B(n9041), .Z(n9040) );
  AND U6056 ( .A(x[6]), .B(y[24]), .Z(n9039) );
  XOR U6057 ( .A(n9040), .B(n9039), .Z(n8988) );
  XOR U6058 ( .A(n8989), .B(n8988), .Z(n8987) );
  XOR U6059 ( .A(n8986), .B(n8987), .Z(n8969) );
  XOR U6060 ( .A(n8968), .B(n8969), .Z(n8967) );
  XOR U6061 ( .A(n8966), .B(n8967), .Z(n8938) );
  XNOR U6062 ( .A(n8939), .B(n8938), .Z(n9197) );
  XNOR U6063 ( .A(n9198), .B(n9197), .Z(n8928) );
  XOR U6064 ( .A(n8929), .B(n8928), .Z(n8927) );
  NANDN U6065 ( .A(n8893), .B(n8892), .Z(n8897) );
  NANDN U6066 ( .A(n8895), .B(n8894), .Z(n8896) );
  AND U6067 ( .A(n8897), .B(n8896), .Z(n8926) );
  XOR U6068 ( .A(n8927), .B(n8926), .Z(n9218) );
  NAND U6069 ( .A(n8899), .B(n8898), .Z(n8903) );
  NANDN U6070 ( .A(n8901), .B(n8900), .Z(n8902) );
  AND U6071 ( .A(n8903), .B(n8902), .Z(n9217) );
  XOR U6072 ( .A(n9215), .B(n9216), .Z(n9212) );
  XNOR U6073 ( .A(n9211), .B(n9212), .Z(n9210) );
  XOR U6074 ( .A(n9209), .B(n9210), .Z(n8920) );
  XNOR U6075 ( .A(n8921), .B(n8920), .Z(N63) );
  XOR U6076 ( .A(n8905), .B(n8904), .Z(n6259) );
  XNOR U6077 ( .A(n8907), .B(n8906), .Z(n6258) );
  XNOR U6078 ( .A(n8909), .B(n8908), .Z(n6257) );
  XOR U6079 ( .A(n8911), .B(n8910), .Z(n8912) );
  XNOR U6080 ( .A(n8913), .B(n8912), .Z(n6256) );
  XOR U6081 ( .A(n8915), .B(n8914), .Z(n6255) );
  XOR U6082 ( .A(n8917), .B(n8916), .Z(n6254) );
  XOR U6083 ( .A(n8919), .B(n8918), .Z(n6253) );
  NAND U6084 ( .A(n8921), .B(n8920), .Z(n8925) );
  NANDN U6085 ( .A(n8923), .B(n8922), .Z(n8924) );
  AND U6086 ( .A(n8925), .B(n8924), .Z(n9208) );
  NAND U6087 ( .A(n8927), .B(n8926), .Z(n8931) );
  NAND U6088 ( .A(n8929), .B(n8928), .Z(n8930) );
  AND U6089 ( .A(n8931), .B(n8930), .Z(n9190) );
  NAND U6090 ( .A(n8933), .B(n8932), .Z(n8937) );
  NAND U6091 ( .A(n8935), .B(n8934), .Z(n8936) );
  AND U6092 ( .A(n8937), .B(n8936), .Z(n8945) );
  NAND U6093 ( .A(n8939), .B(n8938), .Z(n8943) );
  NAND U6094 ( .A(n8941), .B(n8940), .Z(n8942) );
  NAND U6095 ( .A(n8943), .B(n8942), .Z(n8944) );
  XNOR U6096 ( .A(n8945), .B(n8944), .Z(n9188) );
  ANDN U6097 ( .B(n8947), .A(n8946), .Z(n8951) );
  AND U6098 ( .A(n8949), .B(n8948), .Z(n8950) );
  NOR U6099 ( .A(n8951), .B(n8950), .Z(n8959) );
  NANDN U6100 ( .A(n8953), .B(n8952), .Z(n8957) );
  NAND U6101 ( .A(n8955), .B(n8954), .Z(n8956) );
  AND U6102 ( .A(n8957), .B(n8956), .Z(n8958) );
  XNOR U6103 ( .A(n8959), .B(n8958), .Z(n9186) );
  NAND U6104 ( .A(n8961), .B(n8960), .Z(n8965) );
  NANDN U6105 ( .A(n8963), .B(n8962), .Z(n8964) );
  AND U6106 ( .A(n8965), .B(n8964), .Z(n9168) );
  NAND U6107 ( .A(n8967), .B(n8966), .Z(n8971) );
  NAND U6108 ( .A(n8969), .B(n8968), .Z(n8970) );
  AND U6109 ( .A(n8971), .B(n8970), .Z(n8979) );
  NAND U6110 ( .A(n8973), .B(n8972), .Z(n8977) );
  NAND U6111 ( .A(n8975), .B(n8974), .Z(n8976) );
  NAND U6112 ( .A(n8977), .B(n8976), .Z(n8978) );
  XNOR U6113 ( .A(n8979), .B(n8978), .Z(n9166) );
  NAND U6114 ( .A(n8981), .B(n8980), .Z(n8985) );
  NAND U6115 ( .A(n8983), .B(n8982), .Z(n8984) );
  AND U6116 ( .A(n8985), .B(n8984), .Z(n9164) );
  NAND U6117 ( .A(n8987), .B(n8986), .Z(n8991) );
  NAND U6118 ( .A(n8989), .B(n8988), .Z(n8990) );
  AND U6119 ( .A(n8991), .B(n8990), .Z(n8999) );
  NAND U6120 ( .A(n8993), .B(n8992), .Z(n8997) );
  NANDN U6121 ( .A(n8995), .B(n8994), .Z(n8996) );
  NAND U6122 ( .A(n8997), .B(n8996), .Z(n8998) );
  XNOR U6123 ( .A(n8999), .B(n8998), .Z(n9162) );
  NAND U6124 ( .A(n9001), .B(n9000), .Z(n9005) );
  NAND U6125 ( .A(n9003), .B(n9002), .Z(n9004) );
  AND U6126 ( .A(n9005), .B(n9004), .Z(n9160) );
  NAND U6127 ( .A(n9007), .B(n9006), .Z(n9011) );
  NAND U6128 ( .A(n9009), .B(n9008), .Z(n9010) );
  AND U6129 ( .A(n9011), .B(n9010), .Z(n9019) );
  NAND U6130 ( .A(n9013), .B(n9012), .Z(n9017) );
  NAND U6131 ( .A(n9015), .B(n9014), .Z(n9016) );
  NAND U6132 ( .A(n9017), .B(n9016), .Z(n9018) );
  XNOR U6133 ( .A(n9019), .B(n9018), .Z(n9158) );
  NAND U6134 ( .A(n9021), .B(n9020), .Z(n9025) );
  NAND U6135 ( .A(n9023), .B(n9022), .Z(n9024) );
  AND U6136 ( .A(n9025), .B(n9024), .Z(n9033) );
  NAND U6137 ( .A(n9027), .B(n9026), .Z(n9031) );
  NAND U6138 ( .A(n9029), .B(n9028), .Z(n9030) );
  NAND U6139 ( .A(n9031), .B(n9030), .Z(n9032) );
  XNOR U6140 ( .A(n9033), .B(n9032), .Z(n9088) );
  NAND U6141 ( .A(n9035), .B(n9034), .Z(n9038) );
  NAND U6142 ( .A(n9128), .B(n9036), .Z(n9037) );
  AND U6143 ( .A(n9038), .B(n9037), .Z(n9086) );
  NAND U6144 ( .A(n9040), .B(n9039), .Z(n9044) );
  AND U6145 ( .A(n9042), .B(n9041), .Z(n9043) );
  ANDN U6146 ( .B(n9044), .A(n9043), .Z(n9084) );
  NAND U6147 ( .A(n9046), .B(n9045), .Z(n9050) );
  NAND U6148 ( .A(n9048), .B(n9047), .Z(n9049) );
  AND U6149 ( .A(n9050), .B(n9049), .Z(n9082) );
  NAND U6150 ( .A(n9052), .B(n9051), .Z(n9056) );
  NAND U6151 ( .A(n9054), .B(n9053), .Z(n9055) );
  AND U6152 ( .A(n9056), .B(n9055), .Z(n9064) );
  NAND U6153 ( .A(n9058), .B(n9057), .Z(n9062) );
  NAND U6154 ( .A(n9060), .B(n9059), .Z(n9061) );
  NAND U6155 ( .A(n9062), .B(n9061), .Z(n9063) );
  XNOR U6156 ( .A(n9064), .B(n9063), .Z(n9080) );
  AND U6157 ( .A(y[31]), .B(x[0]), .Z(n9066) );
  NAND U6158 ( .A(x[8]), .B(y[23]), .Z(n9065) );
  XNOR U6159 ( .A(n9066), .B(n9065), .Z(n9070) );
  AND U6160 ( .A(y[11]), .B(x[20]), .Z(n9068) );
  NAND U6161 ( .A(y[26]), .B(x[5]), .Z(n9067) );
  XNOR U6162 ( .A(n9068), .B(n9067), .Z(n9069) );
  XOR U6163 ( .A(n9070), .B(n9069), .Z(n9078) );
  AND U6164 ( .A(x[31]), .B(y[0]), .Z(n9072) );
  NAND U6165 ( .A(x[6]), .B(y[25]), .Z(n9071) );
  XNOR U6166 ( .A(n9072), .B(n9071), .Z(n9076) );
  AND U6167 ( .A(x[27]), .B(y[4]), .Z(n9074) );
  NAND U6168 ( .A(y[28]), .B(x[3]), .Z(n9073) );
  XNOR U6169 ( .A(n9074), .B(n9073), .Z(n9075) );
  XNOR U6170 ( .A(n9076), .B(n9075), .Z(n9077) );
  XNOR U6171 ( .A(n9078), .B(n9077), .Z(n9079) );
  XNOR U6172 ( .A(n9080), .B(n9079), .Z(n9081) );
  XNOR U6173 ( .A(n9082), .B(n9081), .Z(n9083) );
  XNOR U6174 ( .A(n9084), .B(n9083), .Z(n9085) );
  XNOR U6175 ( .A(n9086), .B(n9085), .Z(n9087) );
  XOR U6176 ( .A(n9088), .B(n9087), .Z(n9156) );
  AND U6177 ( .A(x[28]), .B(y[3]), .Z(n9090) );
  NAND U6178 ( .A(x[17]), .B(y[14]), .Z(n9089) );
  XNOR U6179 ( .A(n9090), .B(n9089), .Z(n9094) );
  AND U6180 ( .A(x[12]), .B(y[19]), .Z(n9092) );
  NAND U6181 ( .A(x[29]), .B(y[2]), .Z(n9091) );
  XNOR U6182 ( .A(n9092), .B(n9091), .Z(n9093) );
  XOR U6183 ( .A(n9094), .B(n9093), .Z(n9102) );
  AND U6184 ( .A(y[29]), .B(x[2]), .Z(n9096) );
  NAND U6185 ( .A(x[16]), .B(y[15]), .Z(n9095) );
  XNOR U6186 ( .A(n9096), .B(n9095), .Z(n9100) );
  AND U6187 ( .A(y[24]), .B(x[7]), .Z(n9098) );
  NAND U6188 ( .A(x[10]), .B(y[21]), .Z(n9097) );
  XNOR U6189 ( .A(n9098), .B(n9097), .Z(n9099) );
  XNOR U6190 ( .A(n9100), .B(n9099), .Z(n9101) );
  XNOR U6191 ( .A(n9102), .B(n9101), .Z(n9118) );
  AND U6192 ( .A(y[16]), .B(x[15]), .Z(n9104) );
  NAND U6193 ( .A(y[17]), .B(x[14]), .Z(n9103) );
  XNOR U6194 ( .A(n9104), .B(n9103), .Z(n9108) );
  AND U6195 ( .A(x[30]), .B(y[1]), .Z(n9106) );
  NAND U6196 ( .A(x[26]), .B(y[5]), .Z(n9105) );
  XNOR U6197 ( .A(n9106), .B(n9105), .Z(n9107) );
  XOR U6198 ( .A(n9108), .B(n9107), .Z(n9116) );
  AND U6199 ( .A(x[11]), .B(y[20]), .Z(n9110) );
  NAND U6200 ( .A(y[18]), .B(x[13]), .Z(n9109) );
  XNOR U6201 ( .A(n9110), .B(n9109), .Z(n9114) );
  AND U6202 ( .A(x[9]), .B(y[22]), .Z(n9112) );
  NAND U6203 ( .A(x[4]), .B(y[27]), .Z(n9111) );
  XNOR U6204 ( .A(n9112), .B(n9111), .Z(n9113) );
  XNOR U6205 ( .A(n9114), .B(n9113), .Z(n9115) );
  XNOR U6206 ( .A(n9116), .B(n9115), .Z(n9117) );
  XOR U6207 ( .A(n9118), .B(n9117), .Z(n9138) );
  AND U6208 ( .A(y[6]), .B(x[25]), .Z(n9120) );
  NAND U6209 ( .A(y[12]), .B(x[19]), .Z(n9119) );
  XNOR U6210 ( .A(n9120), .B(n9119), .Z(n9136) );
  AND U6211 ( .A(y[13]), .B(x[18]), .Z(n9134) );
  AND U6212 ( .A(n9121), .B(o[30]), .Z(n9132) );
  AND U6213 ( .A(x[22]), .B(y[9]), .Z(n9123) );
  NAND U6214 ( .A(y[10]), .B(x[21]), .Z(n9122) );
  XNOR U6215 ( .A(n9123), .B(n9122), .Z(n9124) );
  XOR U6216 ( .A(o[31]), .B(n9124), .Z(n9130) );
  AND U6217 ( .A(y[30]), .B(x[1]), .Z(n9126) );
  NAND U6218 ( .A(y[8]), .B(x[23]), .Z(n9125) );
  XNOR U6219 ( .A(n9126), .B(n9125), .Z(n9127) );
  XNOR U6220 ( .A(n9128), .B(n9127), .Z(n9129) );
  XNOR U6221 ( .A(n9130), .B(n9129), .Z(n9131) );
  XNOR U6222 ( .A(n9132), .B(n9131), .Z(n9133) );
  XNOR U6223 ( .A(n9134), .B(n9133), .Z(n9135) );
  XNOR U6224 ( .A(n9136), .B(n9135), .Z(n9137) );
  XNOR U6225 ( .A(n9138), .B(n9137), .Z(n9154) );
  NAND U6226 ( .A(n9140), .B(n9139), .Z(n9144) );
  NAND U6227 ( .A(n9142), .B(n9141), .Z(n9143) );
  AND U6228 ( .A(n9144), .B(n9143), .Z(n9152) );
  NAND U6229 ( .A(n9146), .B(n9145), .Z(n9150) );
  NAND U6230 ( .A(n9148), .B(n9147), .Z(n9149) );
  NAND U6231 ( .A(n9150), .B(n9149), .Z(n9151) );
  XNOR U6232 ( .A(n9152), .B(n9151), .Z(n9153) );
  XNOR U6233 ( .A(n9154), .B(n9153), .Z(n9155) );
  XNOR U6234 ( .A(n9156), .B(n9155), .Z(n9157) );
  XNOR U6235 ( .A(n9158), .B(n9157), .Z(n9159) );
  XNOR U6236 ( .A(n9160), .B(n9159), .Z(n9161) );
  XNOR U6237 ( .A(n9162), .B(n9161), .Z(n9163) );
  XNOR U6238 ( .A(n9164), .B(n9163), .Z(n9165) );
  XNOR U6239 ( .A(n9166), .B(n9165), .Z(n9167) );
  XNOR U6240 ( .A(n9168), .B(n9167), .Z(n9184) );
  AND U6241 ( .A(n9170), .B(n9169), .Z(n9174) );
  AND U6242 ( .A(n9172), .B(n9171), .Z(n9173) );
  NOR U6243 ( .A(n9174), .B(n9173), .Z(n9182) );
  NANDN U6244 ( .A(n9176), .B(n9175), .Z(n9180) );
  NAND U6245 ( .A(n9178), .B(n9177), .Z(n9179) );
  AND U6246 ( .A(n9180), .B(n9179), .Z(n9181) );
  XNOR U6247 ( .A(n9182), .B(n9181), .Z(n9183) );
  XNOR U6248 ( .A(n9184), .B(n9183), .Z(n9185) );
  XNOR U6249 ( .A(n9186), .B(n9185), .Z(n9187) );
  XNOR U6250 ( .A(n9188), .B(n9187), .Z(n9189) );
  XNOR U6251 ( .A(n9190), .B(n9189), .Z(n9206) );
  NAND U6252 ( .A(n9192), .B(n9191), .Z(n9196) );
  NAND U6253 ( .A(n9194), .B(n9193), .Z(n9195) );
  AND U6254 ( .A(n9196), .B(n9195), .Z(n9204) );
  NAND U6255 ( .A(n9198), .B(n9197), .Z(n9202) );
  NANDN U6256 ( .A(n9200), .B(n9199), .Z(n9201) );
  NAND U6257 ( .A(n9202), .B(n9201), .Z(n9203) );
  XNOR U6258 ( .A(n9204), .B(n9203), .Z(n9205) );
  XNOR U6259 ( .A(n9206), .B(n9205), .Z(n9207) );
  XNOR U6260 ( .A(n9208), .B(n9207), .Z(n9224) );
  NAND U6261 ( .A(n9210), .B(n9209), .Z(n9214) );
  NANDN U6262 ( .A(n9212), .B(n9211), .Z(n9213) );
  AND U6263 ( .A(n9214), .B(n9213), .Z(n9222) );
  NANDN U6264 ( .A(n9216), .B(n9215), .Z(n9220) );
  NANDN U6265 ( .A(n9218), .B(n9217), .Z(n9219) );
  NAND U6266 ( .A(n9220), .B(n9219), .Z(n9221) );
  XNOR U6267 ( .A(n9222), .B(n9221), .Z(n9223) );
  XNOR U6268 ( .A(n9224), .B(n9223), .Z(n6252) );
endmodule

