
module modmult_step_N512_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [513:0] A;
  input [513:0] B;
  output [513:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560;

  IV U1 ( .A(n2559), .Z(n1) );
  IV U2 ( .A(A[1]), .Z(n2) );
  XNOR U3 ( .A(n3), .B(n4), .Z(DIFF[9]) );
  XOR U4 ( .A(B[9]), .B(A[9]), .Z(n4) );
  XNOR U5 ( .A(n5), .B(n6), .Z(DIFF[99]) );
  XOR U6 ( .A(B[99]), .B(A[99]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(DIFF[98]) );
  XOR U8 ( .A(B[98]), .B(A[98]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(DIFF[97]) );
  XOR U10 ( .A(B[97]), .B(A[97]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(DIFF[96]) );
  XOR U12 ( .A(B[96]), .B(A[96]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(DIFF[95]) );
  XOR U14 ( .A(B[95]), .B(A[95]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(DIFF[94]) );
  XOR U16 ( .A(B[94]), .B(A[94]), .Z(n16) );
  XOR U17 ( .A(n17), .B(n18), .Z(DIFF[93]) );
  XOR U18 ( .A(B[93]), .B(A[93]), .Z(n18) );
  XOR U19 ( .A(n19), .B(n20), .Z(DIFF[92]) );
  XOR U20 ( .A(B[92]), .B(A[92]), .Z(n20) );
  XOR U21 ( .A(n21), .B(n22), .Z(DIFF[91]) );
  XOR U22 ( .A(B[91]), .B(A[91]), .Z(n22) );
  XOR U23 ( .A(n23), .B(n24), .Z(DIFF[90]) );
  XOR U24 ( .A(B[90]), .B(A[90]), .Z(n24) );
  XOR U25 ( .A(n25), .B(n26), .Z(DIFF[8]) );
  XOR U26 ( .A(B[8]), .B(A[8]), .Z(n26) );
  XOR U27 ( .A(n27), .B(n28), .Z(DIFF[89]) );
  XOR U28 ( .A(B[89]), .B(A[89]), .Z(n28) );
  XOR U29 ( .A(n29), .B(n30), .Z(DIFF[88]) );
  XOR U30 ( .A(B[88]), .B(A[88]), .Z(n30) );
  XOR U31 ( .A(n31), .B(n32), .Z(DIFF[87]) );
  XOR U32 ( .A(B[87]), .B(A[87]), .Z(n32) );
  XOR U33 ( .A(n33), .B(n34), .Z(DIFF[86]) );
  XOR U34 ( .A(B[86]), .B(A[86]), .Z(n34) );
  XOR U35 ( .A(n35), .B(n36), .Z(DIFF[85]) );
  XOR U36 ( .A(B[85]), .B(A[85]), .Z(n36) );
  XOR U37 ( .A(n37), .B(n38), .Z(DIFF[84]) );
  XOR U38 ( .A(B[84]), .B(A[84]), .Z(n38) );
  XOR U39 ( .A(n39), .B(n40), .Z(DIFF[83]) );
  XOR U40 ( .A(B[83]), .B(A[83]), .Z(n40) );
  XOR U41 ( .A(n41), .B(n42), .Z(DIFF[82]) );
  XOR U42 ( .A(B[82]), .B(A[82]), .Z(n42) );
  XOR U43 ( .A(n43), .B(n44), .Z(DIFF[81]) );
  XOR U44 ( .A(B[81]), .B(A[81]), .Z(n44) );
  XOR U45 ( .A(n45), .B(n46), .Z(DIFF[80]) );
  XOR U46 ( .A(B[80]), .B(A[80]), .Z(n46) );
  XOR U47 ( .A(n47), .B(n48), .Z(DIFF[7]) );
  XOR U48 ( .A(B[7]), .B(A[7]), .Z(n48) );
  XOR U49 ( .A(n49), .B(n50), .Z(DIFF[79]) );
  XOR U50 ( .A(B[79]), .B(A[79]), .Z(n50) );
  XOR U51 ( .A(n51), .B(n52), .Z(DIFF[78]) );
  XOR U52 ( .A(B[78]), .B(A[78]), .Z(n52) );
  XOR U53 ( .A(n53), .B(n54), .Z(DIFF[77]) );
  XOR U54 ( .A(B[77]), .B(A[77]), .Z(n54) );
  XOR U55 ( .A(n55), .B(n56), .Z(DIFF[76]) );
  XOR U56 ( .A(B[76]), .B(A[76]), .Z(n56) );
  XOR U57 ( .A(n57), .B(n58), .Z(DIFF[75]) );
  XOR U58 ( .A(B[75]), .B(A[75]), .Z(n58) );
  XOR U59 ( .A(n59), .B(n60), .Z(DIFF[74]) );
  XOR U60 ( .A(B[74]), .B(A[74]), .Z(n60) );
  XOR U61 ( .A(n61), .B(n62), .Z(DIFF[73]) );
  XOR U62 ( .A(B[73]), .B(A[73]), .Z(n62) );
  XOR U63 ( .A(n63), .B(n64), .Z(DIFF[72]) );
  XOR U64 ( .A(B[72]), .B(A[72]), .Z(n64) );
  XOR U65 ( .A(n65), .B(n66), .Z(DIFF[71]) );
  XOR U66 ( .A(B[71]), .B(A[71]), .Z(n66) );
  XOR U67 ( .A(n67), .B(n68), .Z(DIFF[70]) );
  XOR U68 ( .A(B[70]), .B(A[70]), .Z(n68) );
  XOR U69 ( .A(n69), .B(n70), .Z(DIFF[6]) );
  XOR U70 ( .A(B[6]), .B(A[6]), .Z(n70) );
  XOR U71 ( .A(n71), .B(n72), .Z(DIFF[69]) );
  XOR U72 ( .A(B[69]), .B(A[69]), .Z(n72) );
  XOR U73 ( .A(n73), .B(n74), .Z(DIFF[68]) );
  XOR U74 ( .A(B[68]), .B(A[68]), .Z(n74) );
  XOR U75 ( .A(n75), .B(n76), .Z(DIFF[67]) );
  XOR U76 ( .A(B[67]), .B(A[67]), .Z(n76) );
  XOR U77 ( .A(n77), .B(n78), .Z(DIFF[66]) );
  XOR U78 ( .A(B[66]), .B(A[66]), .Z(n78) );
  XOR U79 ( .A(n79), .B(n80), .Z(DIFF[65]) );
  XOR U80 ( .A(B[65]), .B(A[65]), .Z(n80) );
  XOR U81 ( .A(n81), .B(n82), .Z(DIFF[64]) );
  XOR U82 ( .A(B[64]), .B(A[64]), .Z(n82) );
  XOR U83 ( .A(n83), .B(n84), .Z(DIFF[63]) );
  XOR U84 ( .A(B[63]), .B(A[63]), .Z(n84) );
  XOR U85 ( .A(n85), .B(n86), .Z(DIFF[62]) );
  XOR U86 ( .A(B[62]), .B(A[62]), .Z(n86) );
  XOR U87 ( .A(n87), .B(n88), .Z(DIFF[61]) );
  XOR U88 ( .A(B[61]), .B(A[61]), .Z(n88) );
  XOR U89 ( .A(n89), .B(n90), .Z(DIFF[60]) );
  XOR U90 ( .A(B[60]), .B(A[60]), .Z(n90) );
  XOR U91 ( .A(n91), .B(n92), .Z(DIFF[5]) );
  XOR U92 ( .A(B[5]), .B(A[5]), .Z(n92) );
  XOR U93 ( .A(n93), .B(n94), .Z(DIFF[59]) );
  XOR U94 ( .A(B[59]), .B(A[59]), .Z(n94) );
  XOR U95 ( .A(n95), .B(n96), .Z(DIFF[58]) );
  XOR U96 ( .A(B[58]), .B(A[58]), .Z(n96) );
  XOR U97 ( .A(n97), .B(n98), .Z(DIFF[57]) );
  XOR U98 ( .A(B[57]), .B(A[57]), .Z(n98) );
  XOR U99 ( .A(n99), .B(n100), .Z(DIFF[56]) );
  XOR U100 ( .A(B[56]), .B(A[56]), .Z(n100) );
  XOR U101 ( .A(n101), .B(n102), .Z(DIFF[55]) );
  XOR U102 ( .A(B[55]), .B(A[55]), .Z(n102) );
  XOR U103 ( .A(n103), .B(n104), .Z(DIFF[54]) );
  XOR U104 ( .A(B[54]), .B(A[54]), .Z(n104) );
  XOR U105 ( .A(n105), .B(n106), .Z(DIFF[53]) );
  XOR U106 ( .A(B[53]), .B(A[53]), .Z(n106) );
  XOR U107 ( .A(n107), .B(n108), .Z(DIFF[52]) );
  XOR U108 ( .A(B[52]), .B(A[52]), .Z(n108) );
  XOR U109 ( .A(n109), .B(n110), .Z(DIFF[51]) );
  XOR U110 ( .A(B[51]), .B(A[51]), .Z(n110) );
  XOR U111 ( .A(A[513]), .B(n111), .Z(DIFF[513]) );
  ANDN U112 ( .B(n112), .A(A[512]), .Z(n111) );
  XOR U113 ( .A(A[512]), .B(n112), .Z(DIFF[512]) );
  AND U114 ( .A(n113), .B(n114), .Z(n112) );
  NANDN U115 ( .A(B[511]), .B(n115), .Z(n114) );
  NANDN U116 ( .A(A[511]), .B(n116), .Z(n115) );
  NANDN U117 ( .A(n116), .B(A[511]), .Z(n113) );
  XOR U118 ( .A(n116), .B(n117), .Z(DIFF[511]) );
  XOR U119 ( .A(B[511]), .B(A[511]), .Z(n117) );
  AND U120 ( .A(n118), .B(n119), .Z(n116) );
  NANDN U121 ( .A(B[510]), .B(n120), .Z(n119) );
  NANDN U122 ( .A(A[510]), .B(n121), .Z(n120) );
  NANDN U123 ( .A(n121), .B(A[510]), .Z(n118) );
  XOR U124 ( .A(n121), .B(n122), .Z(DIFF[510]) );
  XOR U125 ( .A(B[510]), .B(A[510]), .Z(n122) );
  AND U126 ( .A(n123), .B(n124), .Z(n121) );
  NANDN U127 ( .A(B[509]), .B(n125), .Z(n124) );
  NANDN U128 ( .A(A[509]), .B(n126), .Z(n125) );
  NANDN U129 ( .A(n126), .B(A[509]), .Z(n123) );
  XOR U130 ( .A(n127), .B(n128), .Z(DIFF[50]) );
  XOR U131 ( .A(B[50]), .B(A[50]), .Z(n128) );
  XOR U132 ( .A(n126), .B(n129), .Z(DIFF[509]) );
  XOR U133 ( .A(B[509]), .B(A[509]), .Z(n129) );
  AND U134 ( .A(n130), .B(n131), .Z(n126) );
  NANDN U135 ( .A(B[508]), .B(n132), .Z(n131) );
  NANDN U136 ( .A(A[508]), .B(n133), .Z(n132) );
  NANDN U137 ( .A(n133), .B(A[508]), .Z(n130) );
  XOR U138 ( .A(n133), .B(n134), .Z(DIFF[508]) );
  XOR U139 ( .A(B[508]), .B(A[508]), .Z(n134) );
  AND U140 ( .A(n135), .B(n136), .Z(n133) );
  NANDN U141 ( .A(B[507]), .B(n137), .Z(n136) );
  NANDN U142 ( .A(A[507]), .B(n138), .Z(n137) );
  NANDN U143 ( .A(n138), .B(A[507]), .Z(n135) );
  XOR U144 ( .A(n138), .B(n139), .Z(DIFF[507]) );
  XOR U145 ( .A(B[507]), .B(A[507]), .Z(n139) );
  AND U146 ( .A(n140), .B(n141), .Z(n138) );
  NANDN U147 ( .A(B[506]), .B(n142), .Z(n141) );
  NANDN U148 ( .A(A[506]), .B(n143), .Z(n142) );
  NANDN U149 ( .A(n143), .B(A[506]), .Z(n140) );
  XOR U150 ( .A(n143), .B(n144), .Z(DIFF[506]) );
  XOR U151 ( .A(B[506]), .B(A[506]), .Z(n144) );
  AND U152 ( .A(n145), .B(n146), .Z(n143) );
  NANDN U153 ( .A(B[505]), .B(n147), .Z(n146) );
  NANDN U154 ( .A(A[505]), .B(n148), .Z(n147) );
  NANDN U155 ( .A(n148), .B(A[505]), .Z(n145) );
  XOR U156 ( .A(n148), .B(n149), .Z(DIFF[505]) );
  XOR U157 ( .A(B[505]), .B(A[505]), .Z(n149) );
  AND U158 ( .A(n150), .B(n151), .Z(n148) );
  NANDN U159 ( .A(B[504]), .B(n152), .Z(n151) );
  NANDN U160 ( .A(A[504]), .B(n153), .Z(n152) );
  NANDN U161 ( .A(n153), .B(A[504]), .Z(n150) );
  XOR U162 ( .A(n153), .B(n154), .Z(DIFF[504]) );
  XOR U163 ( .A(B[504]), .B(A[504]), .Z(n154) );
  AND U164 ( .A(n155), .B(n156), .Z(n153) );
  NANDN U165 ( .A(B[503]), .B(n157), .Z(n156) );
  NANDN U166 ( .A(A[503]), .B(n158), .Z(n157) );
  NANDN U167 ( .A(n158), .B(A[503]), .Z(n155) );
  XOR U168 ( .A(n158), .B(n159), .Z(DIFF[503]) );
  XOR U169 ( .A(B[503]), .B(A[503]), .Z(n159) );
  AND U170 ( .A(n160), .B(n161), .Z(n158) );
  NANDN U171 ( .A(B[502]), .B(n162), .Z(n161) );
  NANDN U172 ( .A(A[502]), .B(n163), .Z(n162) );
  NANDN U173 ( .A(n163), .B(A[502]), .Z(n160) );
  XOR U174 ( .A(n163), .B(n164), .Z(DIFF[502]) );
  XOR U175 ( .A(B[502]), .B(A[502]), .Z(n164) );
  AND U176 ( .A(n165), .B(n166), .Z(n163) );
  NANDN U177 ( .A(B[501]), .B(n167), .Z(n166) );
  NANDN U178 ( .A(A[501]), .B(n168), .Z(n167) );
  NANDN U179 ( .A(n168), .B(A[501]), .Z(n165) );
  XOR U180 ( .A(n168), .B(n169), .Z(DIFF[501]) );
  XOR U181 ( .A(B[501]), .B(A[501]), .Z(n169) );
  AND U182 ( .A(n170), .B(n171), .Z(n168) );
  NANDN U183 ( .A(B[500]), .B(n172), .Z(n171) );
  NANDN U184 ( .A(A[500]), .B(n173), .Z(n172) );
  NANDN U185 ( .A(n173), .B(A[500]), .Z(n170) );
  XOR U186 ( .A(n173), .B(n174), .Z(DIFF[500]) );
  XOR U187 ( .A(B[500]), .B(A[500]), .Z(n174) );
  AND U188 ( .A(n175), .B(n176), .Z(n173) );
  NANDN U189 ( .A(B[499]), .B(n177), .Z(n176) );
  NANDN U190 ( .A(A[499]), .B(n178), .Z(n177) );
  NANDN U191 ( .A(n178), .B(A[499]), .Z(n175) );
  XOR U192 ( .A(n179), .B(n180), .Z(DIFF[4]) );
  XOR U193 ( .A(B[4]), .B(A[4]), .Z(n180) );
  XOR U194 ( .A(n181), .B(n182), .Z(DIFF[49]) );
  XOR U195 ( .A(B[49]), .B(A[49]), .Z(n182) );
  XOR U196 ( .A(n178), .B(n183), .Z(DIFF[499]) );
  XOR U197 ( .A(B[499]), .B(A[499]), .Z(n183) );
  AND U198 ( .A(n184), .B(n185), .Z(n178) );
  NANDN U199 ( .A(B[498]), .B(n186), .Z(n185) );
  NANDN U200 ( .A(A[498]), .B(n187), .Z(n186) );
  NANDN U201 ( .A(n187), .B(A[498]), .Z(n184) );
  XOR U202 ( .A(n187), .B(n188), .Z(DIFF[498]) );
  XOR U203 ( .A(B[498]), .B(A[498]), .Z(n188) );
  AND U204 ( .A(n189), .B(n190), .Z(n187) );
  NANDN U205 ( .A(B[497]), .B(n191), .Z(n190) );
  NANDN U206 ( .A(A[497]), .B(n192), .Z(n191) );
  NANDN U207 ( .A(n192), .B(A[497]), .Z(n189) );
  XOR U208 ( .A(n192), .B(n193), .Z(DIFF[497]) );
  XOR U209 ( .A(B[497]), .B(A[497]), .Z(n193) );
  AND U210 ( .A(n194), .B(n195), .Z(n192) );
  NANDN U211 ( .A(B[496]), .B(n196), .Z(n195) );
  NANDN U212 ( .A(A[496]), .B(n197), .Z(n196) );
  NANDN U213 ( .A(n197), .B(A[496]), .Z(n194) );
  XOR U214 ( .A(n197), .B(n198), .Z(DIFF[496]) );
  XOR U215 ( .A(B[496]), .B(A[496]), .Z(n198) );
  AND U216 ( .A(n199), .B(n200), .Z(n197) );
  NANDN U217 ( .A(B[495]), .B(n201), .Z(n200) );
  NANDN U218 ( .A(A[495]), .B(n202), .Z(n201) );
  NANDN U219 ( .A(n202), .B(A[495]), .Z(n199) );
  XOR U220 ( .A(n202), .B(n203), .Z(DIFF[495]) );
  XOR U221 ( .A(B[495]), .B(A[495]), .Z(n203) );
  AND U222 ( .A(n204), .B(n205), .Z(n202) );
  NANDN U223 ( .A(B[494]), .B(n206), .Z(n205) );
  NANDN U224 ( .A(A[494]), .B(n207), .Z(n206) );
  NANDN U225 ( .A(n207), .B(A[494]), .Z(n204) );
  XOR U226 ( .A(n207), .B(n208), .Z(DIFF[494]) );
  XOR U227 ( .A(B[494]), .B(A[494]), .Z(n208) );
  AND U228 ( .A(n209), .B(n210), .Z(n207) );
  NANDN U229 ( .A(B[493]), .B(n211), .Z(n210) );
  NANDN U230 ( .A(A[493]), .B(n212), .Z(n211) );
  NANDN U231 ( .A(n212), .B(A[493]), .Z(n209) );
  XOR U232 ( .A(n212), .B(n213), .Z(DIFF[493]) );
  XOR U233 ( .A(B[493]), .B(A[493]), .Z(n213) );
  AND U234 ( .A(n214), .B(n215), .Z(n212) );
  NANDN U235 ( .A(B[492]), .B(n216), .Z(n215) );
  NANDN U236 ( .A(A[492]), .B(n217), .Z(n216) );
  NANDN U237 ( .A(n217), .B(A[492]), .Z(n214) );
  XOR U238 ( .A(n217), .B(n218), .Z(DIFF[492]) );
  XOR U239 ( .A(B[492]), .B(A[492]), .Z(n218) );
  AND U240 ( .A(n219), .B(n220), .Z(n217) );
  NANDN U241 ( .A(B[491]), .B(n221), .Z(n220) );
  NANDN U242 ( .A(A[491]), .B(n222), .Z(n221) );
  NANDN U243 ( .A(n222), .B(A[491]), .Z(n219) );
  XOR U244 ( .A(n222), .B(n223), .Z(DIFF[491]) );
  XOR U245 ( .A(B[491]), .B(A[491]), .Z(n223) );
  AND U246 ( .A(n224), .B(n225), .Z(n222) );
  NANDN U247 ( .A(B[490]), .B(n226), .Z(n225) );
  NANDN U248 ( .A(A[490]), .B(n227), .Z(n226) );
  NANDN U249 ( .A(n227), .B(A[490]), .Z(n224) );
  XOR U250 ( .A(n227), .B(n228), .Z(DIFF[490]) );
  XOR U251 ( .A(B[490]), .B(A[490]), .Z(n228) );
  AND U252 ( .A(n229), .B(n230), .Z(n227) );
  NANDN U253 ( .A(B[489]), .B(n231), .Z(n230) );
  NANDN U254 ( .A(A[489]), .B(n232), .Z(n231) );
  NANDN U255 ( .A(n232), .B(A[489]), .Z(n229) );
  XOR U256 ( .A(n233), .B(n234), .Z(DIFF[48]) );
  XOR U257 ( .A(B[48]), .B(A[48]), .Z(n234) );
  XOR U258 ( .A(n232), .B(n235), .Z(DIFF[489]) );
  XOR U259 ( .A(B[489]), .B(A[489]), .Z(n235) );
  AND U260 ( .A(n236), .B(n237), .Z(n232) );
  NANDN U261 ( .A(B[488]), .B(n238), .Z(n237) );
  NANDN U262 ( .A(A[488]), .B(n239), .Z(n238) );
  NANDN U263 ( .A(n239), .B(A[488]), .Z(n236) );
  XOR U264 ( .A(n239), .B(n240), .Z(DIFF[488]) );
  XOR U265 ( .A(B[488]), .B(A[488]), .Z(n240) );
  AND U266 ( .A(n241), .B(n242), .Z(n239) );
  NANDN U267 ( .A(B[487]), .B(n243), .Z(n242) );
  NANDN U268 ( .A(A[487]), .B(n244), .Z(n243) );
  NANDN U269 ( .A(n244), .B(A[487]), .Z(n241) );
  XOR U270 ( .A(n244), .B(n245), .Z(DIFF[487]) );
  XOR U271 ( .A(B[487]), .B(A[487]), .Z(n245) );
  AND U272 ( .A(n246), .B(n247), .Z(n244) );
  NANDN U273 ( .A(B[486]), .B(n248), .Z(n247) );
  NANDN U274 ( .A(A[486]), .B(n249), .Z(n248) );
  NANDN U275 ( .A(n249), .B(A[486]), .Z(n246) );
  XOR U276 ( .A(n249), .B(n250), .Z(DIFF[486]) );
  XOR U277 ( .A(B[486]), .B(A[486]), .Z(n250) );
  AND U278 ( .A(n251), .B(n252), .Z(n249) );
  NANDN U279 ( .A(B[485]), .B(n253), .Z(n252) );
  NANDN U280 ( .A(A[485]), .B(n254), .Z(n253) );
  NANDN U281 ( .A(n254), .B(A[485]), .Z(n251) );
  XOR U282 ( .A(n254), .B(n255), .Z(DIFF[485]) );
  XOR U283 ( .A(B[485]), .B(A[485]), .Z(n255) );
  AND U284 ( .A(n256), .B(n257), .Z(n254) );
  NANDN U285 ( .A(B[484]), .B(n258), .Z(n257) );
  NANDN U286 ( .A(A[484]), .B(n259), .Z(n258) );
  NANDN U287 ( .A(n259), .B(A[484]), .Z(n256) );
  XOR U288 ( .A(n259), .B(n260), .Z(DIFF[484]) );
  XOR U289 ( .A(B[484]), .B(A[484]), .Z(n260) );
  AND U290 ( .A(n261), .B(n262), .Z(n259) );
  NANDN U291 ( .A(B[483]), .B(n263), .Z(n262) );
  NANDN U292 ( .A(A[483]), .B(n264), .Z(n263) );
  NANDN U293 ( .A(n264), .B(A[483]), .Z(n261) );
  XOR U294 ( .A(n264), .B(n265), .Z(DIFF[483]) );
  XOR U295 ( .A(B[483]), .B(A[483]), .Z(n265) );
  AND U296 ( .A(n266), .B(n267), .Z(n264) );
  NANDN U297 ( .A(B[482]), .B(n268), .Z(n267) );
  NANDN U298 ( .A(A[482]), .B(n269), .Z(n268) );
  NANDN U299 ( .A(n269), .B(A[482]), .Z(n266) );
  XOR U300 ( .A(n269), .B(n270), .Z(DIFF[482]) );
  XOR U301 ( .A(B[482]), .B(A[482]), .Z(n270) );
  AND U302 ( .A(n271), .B(n272), .Z(n269) );
  NANDN U303 ( .A(B[481]), .B(n273), .Z(n272) );
  NANDN U304 ( .A(A[481]), .B(n274), .Z(n273) );
  NANDN U305 ( .A(n274), .B(A[481]), .Z(n271) );
  XOR U306 ( .A(n274), .B(n275), .Z(DIFF[481]) );
  XOR U307 ( .A(B[481]), .B(A[481]), .Z(n275) );
  AND U308 ( .A(n276), .B(n277), .Z(n274) );
  NANDN U309 ( .A(B[480]), .B(n278), .Z(n277) );
  NANDN U310 ( .A(A[480]), .B(n279), .Z(n278) );
  NANDN U311 ( .A(n279), .B(A[480]), .Z(n276) );
  XOR U312 ( .A(n279), .B(n280), .Z(DIFF[480]) );
  XOR U313 ( .A(B[480]), .B(A[480]), .Z(n280) );
  AND U314 ( .A(n281), .B(n282), .Z(n279) );
  NANDN U315 ( .A(B[479]), .B(n283), .Z(n282) );
  NANDN U316 ( .A(A[479]), .B(n284), .Z(n283) );
  NANDN U317 ( .A(n284), .B(A[479]), .Z(n281) );
  XOR U318 ( .A(n285), .B(n286), .Z(DIFF[47]) );
  XOR U319 ( .A(B[47]), .B(A[47]), .Z(n286) );
  XOR U320 ( .A(n284), .B(n287), .Z(DIFF[479]) );
  XOR U321 ( .A(B[479]), .B(A[479]), .Z(n287) );
  AND U322 ( .A(n288), .B(n289), .Z(n284) );
  NANDN U323 ( .A(B[478]), .B(n290), .Z(n289) );
  NANDN U324 ( .A(A[478]), .B(n291), .Z(n290) );
  NANDN U325 ( .A(n291), .B(A[478]), .Z(n288) );
  XOR U326 ( .A(n291), .B(n292), .Z(DIFF[478]) );
  XOR U327 ( .A(B[478]), .B(A[478]), .Z(n292) );
  AND U328 ( .A(n293), .B(n294), .Z(n291) );
  NANDN U329 ( .A(B[477]), .B(n295), .Z(n294) );
  NANDN U330 ( .A(A[477]), .B(n296), .Z(n295) );
  NANDN U331 ( .A(n296), .B(A[477]), .Z(n293) );
  XOR U332 ( .A(n296), .B(n297), .Z(DIFF[477]) );
  XOR U333 ( .A(B[477]), .B(A[477]), .Z(n297) );
  AND U334 ( .A(n298), .B(n299), .Z(n296) );
  NANDN U335 ( .A(B[476]), .B(n300), .Z(n299) );
  NANDN U336 ( .A(A[476]), .B(n301), .Z(n300) );
  NANDN U337 ( .A(n301), .B(A[476]), .Z(n298) );
  XOR U338 ( .A(n301), .B(n302), .Z(DIFF[476]) );
  XOR U339 ( .A(B[476]), .B(A[476]), .Z(n302) );
  AND U340 ( .A(n303), .B(n304), .Z(n301) );
  NANDN U341 ( .A(B[475]), .B(n305), .Z(n304) );
  NANDN U342 ( .A(A[475]), .B(n306), .Z(n305) );
  NANDN U343 ( .A(n306), .B(A[475]), .Z(n303) );
  XOR U344 ( .A(n306), .B(n307), .Z(DIFF[475]) );
  XOR U345 ( .A(B[475]), .B(A[475]), .Z(n307) );
  AND U346 ( .A(n308), .B(n309), .Z(n306) );
  NANDN U347 ( .A(B[474]), .B(n310), .Z(n309) );
  NANDN U348 ( .A(A[474]), .B(n311), .Z(n310) );
  NANDN U349 ( .A(n311), .B(A[474]), .Z(n308) );
  XOR U350 ( .A(n311), .B(n312), .Z(DIFF[474]) );
  XOR U351 ( .A(B[474]), .B(A[474]), .Z(n312) );
  AND U352 ( .A(n313), .B(n314), .Z(n311) );
  NANDN U353 ( .A(B[473]), .B(n315), .Z(n314) );
  NANDN U354 ( .A(A[473]), .B(n316), .Z(n315) );
  NANDN U355 ( .A(n316), .B(A[473]), .Z(n313) );
  XOR U356 ( .A(n316), .B(n317), .Z(DIFF[473]) );
  XOR U357 ( .A(B[473]), .B(A[473]), .Z(n317) );
  AND U358 ( .A(n318), .B(n319), .Z(n316) );
  NANDN U359 ( .A(B[472]), .B(n320), .Z(n319) );
  NANDN U360 ( .A(A[472]), .B(n321), .Z(n320) );
  NANDN U361 ( .A(n321), .B(A[472]), .Z(n318) );
  XOR U362 ( .A(n321), .B(n322), .Z(DIFF[472]) );
  XOR U363 ( .A(B[472]), .B(A[472]), .Z(n322) );
  AND U364 ( .A(n323), .B(n324), .Z(n321) );
  NANDN U365 ( .A(B[471]), .B(n325), .Z(n324) );
  NANDN U366 ( .A(A[471]), .B(n326), .Z(n325) );
  NANDN U367 ( .A(n326), .B(A[471]), .Z(n323) );
  XOR U368 ( .A(n326), .B(n327), .Z(DIFF[471]) );
  XOR U369 ( .A(B[471]), .B(A[471]), .Z(n327) );
  AND U370 ( .A(n328), .B(n329), .Z(n326) );
  NANDN U371 ( .A(B[470]), .B(n330), .Z(n329) );
  NANDN U372 ( .A(A[470]), .B(n331), .Z(n330) );
  NANDN U373 ( .A(n331), .B(A[470]), .Z(n328) );
  XOR U374 ( .A(n331), .B(n332), .Z(DIFF[470]) );
  XOR U375 ( .A(B[470]), .B(A[470]), .Z(n332) );
  AND U376 ( .A(n333), .B(n334), .Z(n331) );
  NANDN U377 ( .A(B[469]), .B(n335), .Z(n334) );
  NANDN U378 ( .A(A[469]), .B(n336), .Z(n335) );
  NANDN U379 ( .A(n336), .B(A[469]), .Z(n333) );
  XOR U380 ( .A(n337), .B(n338), .Z(DIFF[46]) );
  XOR U381 ( .A(B[46]), .B(A[46]), .Z(n338) );
  XOR U382 ( .A(n336), .B(n339), .Z(DIFF[469]) );
  XOR U383 ( .A(B[469]), .B(A[469]), .Z(n339) );
  AND U384 ( .A(n340), .B(n341), .Z(n336) );
  NANDN U385 ( .A(B[468]), .B(n342), .Z(n341) );
  NANDN U386 ( .A(A[468]), .B(n343), .Z(n342) );
  NANDN U387 ( .A(n343), .B(A[468]), .Z(n340) );
  XOR U388 ( .A(n343), .B(n344), .Z(DIFF[468]) );
  XOR U389 ( .A(B[468]), .B(A[468]), .Z(n344) );
  AND U390 ( .A(n345), .B(n346), .Z(n343) );
  NANDN U391 ( .A(B[467]), .B(n347), .Z(n346) );
  NANDN U392 ( .A(A[467]), .B(n348), .Z(n347) );
  NANDN U393 ( .A(n348), .B(A[467]), .Z(n345) );
  XOR U394 ( .A(n348), .B(n349), .Z(DIFF[467]) );
  XOR U395 ( .A(B[467]), .B(A[467]), .Z(n349) );
  AND U396 ( .A(n350), .B(n351), .Z(n348) );
  NANDN U397 ( .A(B[466]), .B(n352), .Z(n351) );
  NANDN U398 ( .A(A[466]), .B(n353), .Z(n352) );
  NANDN U399 ( .A(n353), .B(A[466]), .Z(n350) );
  XOR U400 ( .A(n353), .B(n354), .Z(DIFF[466]) );
  XOR U401 ( .A(B[466]), .B(A[466]), .Z(n354) );
  AND U402 ( .A(n355), .B(n356), .Z(n353) );
  NANDN U403 ( .A(B[465]), .B(n357), .Z(n356) );
  NANDN U404 ( .A(A[465]), .B(n358), .Z(n357) );
  NANDN U405 ( .A(n358), .B(A[465]), .Z(n355) );
  XOR U406 ( .A(n358), .B(n359), .Z(DIFF[465]) );
  XOR U407 ( .A(B[465]), .B(A[465]), .Z(n359) );
  AND U408 ( .A(n360), .B(n361), .Z(n358) );
  NANDN U409 ( .A(B[464]), .B(n362), .Z(n361) );
  NANDN U410 ( .A(A[464]), .B(n363), .Z(n362) );
  NANDN U411 ( .A(n363), .B(A[464]), .Z(n360) );
  XOR U412 ( .A(n363), .B(n364), .Z(DIFF[464]) );
  XOR U413 ( .A(B[464]), .B(A[464]), .Z(n364) );
  AND U414 ( .A(n365), .B(n366), .Z(n363) );
  NANDN U415 ( .A(B[463]), .B(n367), .Z(n366) );
  NANDN U416 ( .A(A[463]), .B(n368), .Z(n367) );
  NANDN U417 ( .A(n368), .B(A[463]), .Z(n365) );
  XOR U418 ( .A(n368), .B(n369), .Z(DIFF[463]) );
  XOR U419 ( .A(B[463]), .B(A[463]), .Z(n369) );
  AND U420 ( .A(n370), .B(n371), .Z(n368) );
  NANDN U421 ( .A(B[462]), .B(n372), .Z(n371) );
  NANDN U422 ( .A(A[462]), .B(n373), .Z(n372) );
  NANDN U423 ( .A(n373), .B(A[462]), .Z(n370) );
  XOR U424 ( .A(n373), .B(n374), .Z(DIFF[462]) );
  XOR U425 ( .A(B[462]), .B(A[462]), .Z(n374) );
  AND U426 ( .A(n375), .B(n376), .Z(n373) );
  NANDN U427 ( .A(B[461]), .B(n377), .Z(n376) );
  NANDN U428 ( .A(A[461]), .B(n378), .Z(n377) );
  NANDN U429 ( .A(n378), .B(A[461]), .Z(n375) );
  XOR U430 ( .A(n378), .B(n379), .Z(DIFF[461]) );
  XOR U431 ( .A(B[461]), .B(A[461]), .Z(n379) );
  AND U432 ( .A(n380), .B(n381), .Z(n378) );
  NANDN U433 ( .A(B[460]), .B(n382), .Z(n381) );
  NANDN U434 ( .A(A[460]), .B(n383), .Z(n382) );
  NANDN U435 ( .A(n383), .B(A[460]), .Z(n380) );
  XOR U436 ( .A(n383), .B(n384), .Z(DIFF[460]) );
  XOR U437 ( .A(B[460]), .B(A[460]), .Z(n384) );
  AND U438 ( .A(n385), .B(n386), .Z(n383) );
  NANDN U439 ( .A(B[459]), .B(n387), .Z(n386) );
  NANDN U440 ( .A(A[459]), .B(n388), .Z(n387) );
  NANDN U441 ( .A(n388), .B(A[459]), .Z(n385) );
  XOR U442 ( .A(n389), .B(n390), .Z(DIFF[45]) );
  XOR U443 ( .A(B[45]), .B(A[45]), .Z(n390) );
  XOR U444 ( .A(n388), .B(n391), .Z(DIFF[459]) );
  XOR U445 ( .A(B[459]), .B(A[459]), .Z(n391) );
  AND U446 ( .A(n392), .B(n393), .Z(n388) );
  NANDN U447 ( .A(B[458]), .B(n394), .Z(n393) );
  NANDN U448 ( .A(A[458]), .B(n395), .Z(n394) );
  NANDN U449 ( .A(n395), .B(A[458]), .Z(n392) );
  XOR U450 ( .A(n395), .B(n396), .Z(DIFF[458]) );
  XOR U451 ( .A(B[458]), .B(A[458]), .Z(n396) );
  AND U452 ( .A(n397), .B(n398), .Z(n395) );
  NANDN U453 ( .A(B[457]), .B(n399), .Z(n398) );
  NANDN U454 ( .A(A[457]), .B(n400), .Z(n399) );
  NANDN U455 ( .A(n400), .B(A[457]), .Z(n397) );
  XOR U456 ( .A(n400), .B(n401), .Z(DIFF[457]) );
  XOR U457 ( .A(B[457]), .B(A[457]), .Z(n401) );
  AND U458 ( .A(n402), .B(n403), .Z(n400) );
  NANDN U459 ( .A(B[456]), .B(n404), .Z(n403) );
  NANDN U460 ( .A(A[456]), .B(n405), .Z(n404) );
  NANDN U461 ( .A(n405), .B(A[456]), .Z(n402) );
  XOR U462 ( .A(n405), .B(n406), .Z(DIFF[456]) );
  XOR U463 ( .A(B[456]), .B(A[456]), .Z(n406) );
  AND U464 ( .A(n407), .B(n408), .Z(n405) );
  NANDN U465 ( .A(B[455]), .B(n409), .Z(n408) );
  NANDN U466 ( .A(A[455]), .B(n410), .Z(n409) );
  NANDN U467 ( .A(n410), .B(A[455]), .Z(n407) );
  XOR U468 ( .A(n410), .B(n411), .Z(DIFF[455]) );
  XOR U469 ( .A(B[455]), .B(A[455]), .Z(n411) );
  AND U470 ( .A(n412), .B(n413), .Z(n410) );
  NANDN U471 ( .A(B[454]), .B(n414), .Z(n413) );
  NANDN U472 ( .A(A[454]), .B(n415), .Z(n414) );
  NANDN U473 ( .A(n415), .B(A[454]), .Z(n412) );
  XOR U474 ( .A(n415), .B(n416), .Z(DIFF[454]) );
  XOR U475 ( .A(B[454]), .B(A[454]), .Z(n416) );
  AND U476 ( .A(n417), .B(n418), .Z(n415) );
  NANDN U477 ( .A(B[453]), .B(n419), .Z(n418) );
  NANDN U478 ( .A(A[453]), .B(n420), .Z(n419) );
  NANDN U479 ( .A(n420), .B(A[453]), .Z(n417) );
  XOR U480 ( .A(n420), .B(n421), .Z(DIFF[453]) );
  XOR U481 ( .A(B[453]), .B(A[453]), .Z(n421) );
  AND U482 ( .A(n422), .B(n423), .Z(n420) );
  NANDN U483 ( .A(B[452]), .B(n424), .Z(n423) );
  NANDN U484 ( .A(A[452]), .B(n425), .Z(n424) );
  NANDN U485 ( .A(n425), .B(A[452]), .Z(n422) );
  XOR U486 ( .A(n425), .B(n426), .Z(DIFF[452]) );
  XOR U487 ( .A(B[452]), .B(A[452]), .Z(n426) );
  AND U488 ( .A(n427), .B(n428), .Z(n425) );
  NANDN U489 ( .A(B[451]), .B(n429), .Z(n428) );
  NANDN U490 ( .A(A[451]), .B(n430), .Z(n429) );
  NANDN U491 ( .A(n430), .B(A[451]), .Z(n427) );
  XOR U492 ( .A(n430), .B(n431), .Z(DIFF[451]) );
  XOR U493 ( .A(B[451]), .B(A[451]), .Z(n431) );
  AND U494 ( .A(n432), .B(n433), .Z(n430) );
  NANDN U495 ( .A(B[450]), .B(n434), .Z(n433) );
  NANDN U496 ( .A(A[450]), .B(n435), .Z(n434) );
  NANDN U497 ( .A(n435), .B(A[450]), .Z(n432) );
  XOR U498 ( .A(n435), .B(n436), .Z(DIFF[450]) );
  XOR U499 ( .A(B[450]), .B(A[450]), .Z(n436) );
  AND U500 ( .A(n437), .B(n438), .Z(n435) );
  NANDN U501 ( .A(B[449]), .B(n439), .Z(n438) );
  NANDN U502 ( .A(A[449]), .B(n440), .Z(n439) );
  NANDN U503 ( .A(n440), .B(A[449]), .Z(n437) );
  XOR U504 ( .A(n441), .B(n442), .Z(DIFF[44]) );
  XOR U505 ( .A(B[44]), .B(A[44]), .Z(n442) );
  XOR U506 ( .A(n440), .B(n443), .Z(DIFF[449]) );
  XOR U507 ( .A(B[449]), .B(A[449]), .Z(n443) );
  AND U508 ( .A(n444), .B(n445), .Z(n440) );
  NANDN U509 ( .A(B[448]), .B(n446), .Z(n445) );
  NANDN U510 ( .A(A[448]), .B(n447), .Z(n446) );
  NANDN U511 ( .A(n447), .B(A[448]), .Z(n444) );
  XOR U512 ( .A(n447), .B(n448), .Z(DIFF[448]) );
  XOR U513 ( .A(B[448]), .B(A[448]), .Z(n448) );
  AND U514 ( .A(n449), .B(n450), .Z(n447) );
  NANDN U515 ( .A(B[447]), .B(n451), .Z(n450) );
  NANDN U516 ( .A(A[447]), .B(n452), .Z(n451) );
  NANDN U517 ( .A(n452), .B(A[447]), .Z(n449) );
  XOR U518 ( .A(n452), .B(n453), .Z(DIFF[447]) );
  XOR U519 ( .A(B[447]), .B(A[447]), .Z(n453) );
  AND U520 ( .A(n454), .B(n455), .Z(n452) );
  NANDN U521 ( .A(B[446]), .B(n456), .Z(n455) );
  NANDN U522 ( .A(A[446]), .B(n457), .Z(n456) );
  NANDN U523 ( .A(n457), .B(A[446]), .Z(n454) );
  XOR U524 ( .A(n457), .B(n458), .Z(DIFF[446]) );
  XOR U525 ( .A(B[446]), .B(A[446]), .Z(n458) );
  AND U526 ( .A(n459), .B(n460), .Z(n457) );
  NANDN U527 ( .A(B[445]), .B(n461), .Z(n460) );
  NANDN U528 ( .A(A[445]), .B(n462), .Z(n461) );
  NANDN U529 ( .A(n462), .B(A[445]), .Z(n459) );
  XOR U530 ( .A(n462), .B(n463), .Z(DIFF[445]) );
  XOR U531 ( .A(B[445]), .B(A[445]), .Z(n463) );
  AND U532 ( .A(n464), .B(n465), .Z(n462) );
  NANDN U533 ( .A(B[444]), .B(n466), .Z(n465) );
  NANDN U534 ( .A(A[444]), .B(n467), .Z(n466) );
  NANDN U535 ( .A(n467), .B(A[444]), .Z(n464) );
  XOR U536 ( .A(n467), .B(n468), .Z(DIFF[444]) );
  XOR U537 ( .A(B[444]), .B(A[444]), .Z(n468) );
  AND U538 ( .A(n469), .B(n470), .Z(n467) );
  NANDN U539 ( .A(B[443]), .B(n471), .Z(n470) );
  NANDN U540 ( .A(A[443]), .B(n472), .Z(n471) );
  NANDN U541 ( .A(n472), .B(A[443]), .Z(n469) );
  XOR U542 ( .A(n472), .B(n473), .Z(DIFF[443]) );
  XOR U543 ( .A(B[443]), .B(A[443]), .Z(n473) );
  AND U544 ( .A(n474), .B(n475), .Z(n472) );
  NANDN U545 ( .A(B[442]), .B(n476), .Z(n475) );
  NANDN U546 ( .A(A[442]), .B(n477), .Z(n476) );
  NANDN U547 ( .A(n477), .B(A[442]), .Z(n474) );
  XOR U548 ( .A(n477), .B(n478), .Z(DIFF[442]) );
  XOR U549 ( .A(B[442]), .B(A[442]), .Z(n478) );
  AND U550 ( .A(n479), .B(n480), .Z(n477) );
  NANDN U551 ( .A(B[441]), .B(n481), .Z(n480) );
  NANDN U552 ( .A(A[441]), .B(n482), .Z(n481) );
  NANDN U553 ( .A(n482), .B(A[441]), .Z(n479) );
  XOR U554 ( .A(n482), .B(n483), .Z(DIFF[441]) );
  XOR U555 ( .A(B[441]), .B(A[441]), .Z(n483) );
  AND U556 ( .A(n484), .B(n485), .Z(n482) );
  NANDN U557 ( .A(B[440]), .B(n486), .Z(n485) );
  NANDN U558 ( .A(A[440]), .B(n487), .Z(n486) );
  NANDN U559 ( .A(n487), .B(A[440]), .Z(n484) );
  XOR U560 ( .A(n487), .B(n488), .Z(DIFF[440]) );
  XOR U561 ( .A(B[440]), .B(A[440]), .Z(n488) );
  AND U562 ( .A(n489), .B(n490), .Z(n487) );
  NANDN U563 ( .A(B[439]), .B(n491), .Z(n490) );
  NANDN U564 ( .A(A[439]), .B(n492), .Z(n491) );
  NANDN U565 ( .A(n492), .B(A[439]), .Z(n489) );
  XOR U566 ( .A(n493), .B(n494), .Z(DIFF[43]) );
  XOR U567 ( .A(B[43]), .B(A[43]), .Z(n494) );
  XOR U568 ( .A(n492), .B(n495), .Z(DIFF[439]) );
  XOR U569 ( .A(B[439]), .B(A[439]), .Z(n495) );
  AND U570 ( .A(n496), .B(n497), .Z(n492) );
  NANDN U571 ( .A(B[438]), .B(n498), .Z(n497) );
  NANDN U572 ( .A(A[438]), .B(n499), .Z(n498) );
  NANDN U573 ( .A(n499), .B(A[438]), .Z(n496) );
  XOR U574 ( .A(n499), .B(n500), .Z(DIFF[438]) );
  XOR U575 ( .A(B[438]), .B(A[438]), .Z(n500) );
  AND U576 ( .A(n501), .B(n502), .Z(n499) );
  NANDN U577 ( .A(B[437]), .B(n503), .Z(n502) );
  NANDN U578 ( .A(A[437]), .B(n504), .Z(n503) );
  NANDN U579 ( .A(n504), .B(A[437]), .Z(n501) );
  XOR U580 ( .A(n504), .B(n505), .Z(DIFF[437]) );
  XOR U581 ( .A(B[437]), .B(A[437]), .Z(n505) );
  AND U582 ( .A(n506), .B(n507), .Z(n504) );
  NANDN U583 ( .A(B[436]), .B(n508), .Z(n507) );
  NANDN U584 ( .A(A[436]), .B(n509), .Z(n508) );
  NANDN U585 ( .A(n509), .B(A[436]), .Z(n506) );
  XOR U586 ( .A(n509), .B(n510), .Z(DIFF[436]) );
  XOR U587 ( .A(B[436]), .B(A[436]), .Z(n510) );
  AND U588 ( .A(n511), .B(n512), .Z(n509) );
  NANDN U589 ( .A(B[435]), .B(n513), .Z(n512) );
  NANDN U590 ( .A(A[435]), .B(n514), .Z(n513) );
  NANDN U591 ( .A(n514), .B(A[435]), .Z(n511) );
  XOR U592 ( .A(n514), .B(n515), .Z(DIFF[435]) );
  XOR U593 ( .A(B[435]), .B(A[435]), .Z(n515) );
  AND U594 ( .A(n516), .B(n517), .Z(n514) );
  NANDN U595 ( .A(B[434]), .B(n518), .Z(n517) );
  NANDN U596 ( .A(A[434]), .B(n519), .Z(n518) );
  NANDN U597 ( .A(n519), .B(A[434]), .Z(n516) );
  XOR U598 ( .A(n519), .B(n520), .Z(DIFF[434]) );
  XOR U599 ( .A(B[434]), .B(A[434]), .Z(n520) );
  AND U600 ( .A(n521), .B(n522), .Z(n519) );
  NANDN U601 ( .A(B[433]), .B(n523), .Z(n522) );
  NANDN U602 ( .A(A[433]), .B(n524), .Z(n523) );
  NANDN U603 ( .A(n524), .B(A[433]), .Z(n521) );
  XOR U604 ( .A(n524), .B(n525), .Z(DIFF[433]) );
  XOR U605 ( .A(B[433]), .B(A[433]), .Z(n525) );
  AND U606 ( .A(n526), .B(n527), .Z(n524) );
  NANDN U607 ( .A(B[432]), .B(n528), .Z(n527) );
  NANDN U608 ( .A(A[432]), .B(n529), .Z(n528) );
  NANDN U609 ( .A(n529), .B(A[432]), .Z(n526) );
  XOR U610 ( .A(n529), .B(n530), .Z(DIFF[432]) );
  XOR U611 ( .A(B[432]), .B(A[432]), .Z(n530) );
  AND U612 ( .A(n531), .B(n532), .Z(n529) );
  NANDN U613 ( .A(B[431]), .B(n533), .Z(n532) );
  NANDN U614 ( .A(A[431]), .B(n534), .Z(n533) );
  NANDN U615 ( .A(n534), .B(A[431]), .Z(n531) );
  XOR U616 ( .A(n534), .B(n535), .Z(DIFF[431]) );
  XOR U617 ( .A(B[431]), .B(A[431]), .Z(n535) );
  AND U618 ( .A(n536), .B(n537), .Z(n534) );
  NANDN U619 ( .A(B[430]), .B(n538), .Z(n537) );
  NANDN U620 ( .A(A[430]), .B(n539), .Z(n538) );
  NANDN U621 ( .A(n539), .B(A[430]), .Z(n536) );
  XOR U622 ( .A(n539), .B(n540), .Z(DIFF[430]) );
  XOR U623 ( .A(B[430]), .B(A[430]), .Z(n540) );
  AND U624 ( .A(n541), .B(n542), .Z(n539) );
  NANDN U625 ( .A(B[429]), .B(n543), .Z(n542) );
  NANDN U626 ( .A(A[429]), .B(n544), .Z(n543) );
  NANDN U627 ( .A(n544), .B(A[429]), .Z(n541) );
  XOR U628 ( .A(n545), .B(n546), .Z(DIFF[42]) );
  XOR U629 ( .A(B[42]), .B(A[42]), .Z(n546) );
  XOR U630 ( .A(n544), .B(n547), .Z(DIFF[429]) );
  XOR U631 ( .A(B[429]), .B(A[429]), .Z(n547) );
  AND U632 ( .A(n548), .B(n549), .Z(n544) );
  NANDN U633 ( .A(B[428]), .B(n550), .Z(n549) );
  NANDN U634 ( .A(A[428]), .B(n551), .Z(n550) );
  NANDN U635 ( .A(n551), .B(A[428]), .Z(n548) );
  XOR U636 ( .A(n551), .B(n552), .Z(DIFF[428]) );
  XOR U637 ( .A(B[428]), .B(A[428]), .Z(n552) );
  AND U638 ( .A(n553), .B(n554), .Z(n551) );
  NANDN U639 ( .A(B[427]), .B(n555), .Z(n554) );
  NANDN U640 ( .A(A[427]), .B(n556), .Z(n555) );
  NANDN U641 ( .A(n556), .B(A[427]), .Z(n553) );
  XOR U642 ( .A(n556), .B(n557), .Z(DIFF[427]) );
  XOR U643 ( .A(B[427]), .B(A[427]), .Z(n557) );
  AND U644 ( .A(n558), .B(n559), .Z(n556) );
  NANDN U645 ( .A(B[426]), .B(n560), .Z(n559) );
  NANDN U646 ( .A(A[426]), .B(n561), .Z(n560) );
  NANDN U647 ( .A(n561), .B(A[426]), .Z(n558) );
  XOR U648 ( .A(n561), .B(n562), .Z(DIFF[426]) );
  XOR U649 ( .A(B[426]), .B(A[426]), .Z(n562) );
  AND U650 ( .A(n563), .B(n564), .Z(n561) );
  NANDN U651 ( .A(B[425]), .B(n565), .Z(n564) );
  NANDN U652 ( .A(A[425]), .B(n566), .Z(n565) );
  NANDN U653 ( .A(n566), .B(A[425]), .Z(n563) );
  XOR U654 ( .A(n566), .B(n567), .Z(DIFF[425]) );
  XOR U655 ( .A(B[425]), .B(A[425]), .Z(n567) );
  AND U656 ( .A(n568), .B(n569), .Z(n566) );
  NANDN U657 ( .A(B[424]), .B(n570), .Z(n569) );
  NANDN U658 ( .A(A[424]), .B(n571), .Z(n570) );
  NANDN U659 ( .A(n571), .B(A[424]), .Z(n568) );
  XOR U660 ( .A(n571), .B(n572), .Z(DIFF[424]) );
  XOR U661 ( .A(B[424]), .B(A[424]), .Z(n572) );
  AND U662 ( .A(n573), .B(n574), .Z(n571) );
  NANDN U663 ( .A(B[423]), .B(n575), .Z(n574) );
  NANDN U664 ( .A(A[423]), .B(n576), .Z(n575) );
  NANDN U665 ( .A(n576), .B(A[423]), .Z(n573) );
  XOR U666 ( .A(n576), .B(n577), .Z(DIFF[423]) );
  XOR U667 ( .A(B[423]), .B(A[423]), .Z(n577) );
  AND U668 ( .A(n578), .B(n579), .Z(n576) );
  NANDN U669 ( .A(B[422]), .B(n580), .Z(n579) );
  NANDN U670 ( .A(A[422]), .B(n581), .Z(n580) );
  NANDN U671 ( .A(n581), .B(A[422]), .Z(n578) );
  XOR U672 ( .A(n581), .B(n582), .Z(DIFF[422]) );
  XOR U673 ( .A(B[422]), .B(A[422]), .Z(n582) );
  AND U674 ( .A(n583), .B(n584), .Z(n581) );
  NANDN U675 ( .A(B[421]), .B(n585), .Z(n584) );
  NANDN U676 ( .A(A[421]), .B(n586), .Z(n585) );
  NANDN U677 ( .A(n586), .B(A[421]), .Z(n583) );
  XOR U678 ( .A(n586), .B(n587), .Z(DIFF[421]) );
  XOR U679 ( .A(B[421]), .B(A[421]), .Z(n587) );
  AND U680 ( .A(n588), .B(n589), .Z(n586) );
  NANDN U681 ( .A(B[420]), .B(n590), .Z(n589) );
  NANDN U682 ( .A(A[420]), .B(n591), .Z(n590) );
  NANDN U683 ( .A(n591), .B(A[420]), .Z(n588) );
  XOR U684 ( .A(n591), .B(n592), .Z(DIFF[420]) );
  XOR U685 ( .A(B[420]), .B(A[420]), .Z(n592) );
  AND U686 ( .A(n593), .B(n594), .Z(n591) );
  NANDN U687 ( .A(B[419]), .B(n595), .Z(n594) );
  NANDN U688 ( .A(A[419]), .B(n596), .Z(n595) );
  NANDN U689 ( .A(n596), .B(A[419]), .Z(n593) );
  XOR U690 ( .A(n597), .B(n598), .Z(DIFF[41]) );
  XOR U691 ( .A(B[41]), .B(A[41]), .Z(n598) );
  XOR U692 ( .A(n596), .B(n599), .Z(DIFF[419]) );
  XOR U693 ( .A(B[419]), .B(A[419]), .Z(n599) );
  AND U694 ( .A(n600), .B(n601), .Z(n596) );
  NANDN U695 ( .A(B[418]), .B(n602), .Z(n601) );
  NANDN U696 ( .A(A[418]), .B(n603), .Z(n602) );
  NANDN U697 ( .A(n603), .B(A[418]), .Z(n600) );
  XOR U698 ( .A(n603), .B(n604), .Z(DIFF[418]) );
  XOR U699 ( .A(B[418]), .B(A[418]), .Z(n604) );
  AND U700 ( .A(n605), .B(n606), .Z(n603) );
  NANDN U701 ( .A(B[417]), .B(n607), .Z(n606) );
  NANDN U702 ( .A(A[417]), .B(n608), .Z(n607) );
  NANDN U703 ( .A(n608), .B(A[417]), .Z(n605) );
  XOR U704 ( .A(n608), .B(n609), .Z(DIFF[417]) );
  XOR U705 ( .A(B[417]), .B(A[417]), .Z(n609) );
  AND U706 ( .A(n610), .B(n611), .Z(n608) );
  NANDN U707 ( .A(B[416]), .B(n612), .Z(n611) );
  NANDN U708 ( .A(A[416]), .B(n613), .Z(n612) );
  NANDN U709 ( .A(n613), .B(A[416]), .Z(n610) );
  XOR U710 ( .A(n613), .B(n614), .Z(DIFF[416]) );
  XOR U711 ( .A(B[416]), .B(A[416]), .Z(n614) );
  AND U712 ( .A(n615), .B(n616), .Z(n613) );
  NANDN U713 ( .A(B[415]), .B(n617), .Z(n616) );
  NANDN U714 ( .A(A[415]), .B(n618), .Z(n617) );
  NANDN U715 ( .A(n618), .B(A[415]), .Z(n615) );
  XOR U716 ( .A(n618), .B(n619), .Z(DIFF[415]) );
  XOR U717 ( .A(B[415]), .B(A[415]), .Z(n619) );
  AND U718 ( .A(n620), .B(n621), .Z(n618) );
  NANDN U719 ( .A(B[414]), .B(n622), .Z(n621) );
  NANDN U720 ( .A(A[414]), .B(n623), .Z(n622) );
  NANDN U721 ( .A(n623), .B(A[414]), .Z(n620) );
  XOR U722 ( .A(n623), .B(n624), .Z(DIFF[414]) );
  XOR U723 ( .A(B[414]), .B(A[414]), .Z(n624) );
  AND U724 ( .A(n625), .B(n626), .Z(n623) );
  NANDN U725 ( .A(B[413]), .B(n627), .Z(n626) );
  NANDN U726 ( .A(A[413]), .B(n628), .Z(n627) );
  NANDN U727 ( .A(n628), .B(A[413]), .Z(n625) );
  XOR U728 ( .A(n628), .B(n629), .Z(DIFF[413]) );
  XOR U729 ( .A(B[413]), .B(A[413]), .Z(n629) );
  AND U730 ( .A(n630), .B(n631), .Z(n628) );
  NANDN U731 ( .A(B[412]), .B(n632), .Z(n631) );
  NANDN U732 ( .A(A[412]), .B(n633), .Z(n632) );
  NANDN U733 ( .A(n633), .B(A[412]), .Z(n630) );
  XOR U734 ( .A(n633), .B(n634), .Z(DIFF[412]) );
  XOR U735 ( .A(B[412]), .B(A[412]), .Z(n634) );
  AND U736 ( .A(n635), .B(n636), .Z(n633) );
  NANDN U737 ( .A(B[411]), .B(n637), .Z(n636) );
  NANDN U738 ( .A(A[411]), .B(n638), .Z(n637) );
  NANDN U739 ( .A(n638), .B(A[411]), .Z(n635) );
  XOR U740 ( .A(n638), .B(n639), .Z(DIFF[411]) );
  XOR U741 ( .A(B[411]), .B(A[411]), .Z(n639) );
  AND U742 ( .A(n640), .B(n641), .Z(n638) );
  NANDN U743 ( .A(B[410]), .B(n642), .Z(n641) );
  NANDN U744 ( .A(A[410]), .B(n643), .Z(n642) );
  NANDN U745 ( .A(n643), .B(A[410]), .Z(n640) );
  XOR U746 ( .A(n643), .B(n644), .Z(DIFF[410]) );
  XOR U747 ( .A(B[410]), .B(A[410]), .Z(n644) );
  AND U748 ( .A(n645), .B(n646), .Z(n643) );
  NANDN U749 ( .A(B[409]), .B(n647), .Z(n646) );
  NANDN U750 ( .A(A[409]), .B(n648), .Z(n647) );
  NANDN U751 ( .A(n648), .B(A[409]), .Z(n645) );
  XOR U752 ( .A(n649), .B(n650), .Z(DIFF[40]) );
  XOR U753 ( .A(B[40]), .B(A[40]), .Z(n650) );
  XOR U754 ( .A(n648), .B(n651), .Z(DIFF[409]) );
  XOR U755 ( .A(B[409]), .B(A[409]), .Z(n651) );
  AND U756 ( .A(n652), .B(n653), .Z(n648) );
  NANDN U757 ( .A(B[408]), .B(n654), .Z(n653) );
  NANDN U758 ( .A(A[408]), .B(n655), .Z(n654) );
  NANDN U759 ( .A(n655), .B(A[408]), .Z(n652) );
  XOR U760 ( .A(n655), .B(n656), .Z(DIFF[408]) );
  XOR U761 ( .A(B[408]), .B(A[408]), .Z(n656) );
  AND U762 ( .A(n657), .B(n658), .Z(n655) );
  NANDN U763 ( .A(B[407]), .B(n659), .Z(n658) );
  NANDN U764 ( .A(A[407]), .B(n660), .Z(n659) );
  NANDN U765 ( .A(n660), .B(A[407]), .Z(n657) );
  XOR U766 ( .A(n660), .B(n661), .Z(DIFF[407]) );
  XOR U767 ( .A(B[407]), .B(A[407]), .Z(n661) );
  AND U768 ( .A(n662), .B(n663), .Z(n660) );
  NANDN U769 ( .A(B[406]), .B(n664), .Z(n663) );
  NANDN U770 ( .A(A[406]), .B(n665), .Z(n664) );
  NANDN U771 ( .A(n665), .B(A[406]), .Z(n662) );
  XOR U772 ( .A(n665), .B(n666), .Z(DIFF[406]) );
  XOR U773 ( .A(B[406]), .B(A[406]), .Z(n666) );
  AND U774 ( .A(n667), .B(n668), .Z(n665) );
  NANDN U775 ( .A(B[405]), .B(n669), .Z(n668) );
  NANDN U776 ( .A(A[405]), .B(n670), .Z(n669) );
  NANDN U777 ( .A(n670), .B(A[405]), .Z(n667) );
  XOR U778 ( .A(n670), .B(n671), .Z(DIFF[405]) );
  XOR U779 ( .A(B[405]), .B(A[405]), .Z(n671) );
  AND U780 ( .A(n672), .B(n673), .Z(n670) );
  NANDN U781 ( .A(B[404]), .B(n674), .Z(n673) );
  NANDN U782 ( .A(A[404]), .B(n675), .Z(n674) );
  NANDN U783 ( .A(n675), .B(A[404]), .Z(n672) );
  XOR U784 ( .A(n675), .B(n676), .Z(DIFF[404]) );
  XOR U785 ( .A(B[404]), .B(A[404]), .Z(n676) );
  AND U786 ( .A(n677), .B(n678), .Z(n675) );
  NANDN U787 ( .A(B[403]), .B(n679), .Z(n678) );
  NANDN U788 ( .A(A[403]), .B(n680), .Z(n679) );
  NANDN U789 ( .A(n680), .B(A[403]), .Z(n677) );
  XOR U790 ( .A(n680), .B(n681), .Z(DIFF[403]) );
  XOR U791 ( .A(B[403]), .B(A[403]), .Z(n681) );
  AND U792 ( .A(n682), .B(n683), .Z(n680) );
  NANDN U793 ( .A(B[402]), .B(n684), .Z(n683) );
  NANDN U794 ( .A(A[402]), .B(n685), .Z(n684) );
  NANDN U795 ( .A(n685), .B(A[402]), .Z(n682) );
  XOR U796 ( .A(n685), .B(n686), .Z(DIFF[402]) );
  XOR U797 ( .A(B[402]), .B(A[402]), .Z(n686) );
  AND U798 ( .A(n687), .B(n688), .Z(n685) );
  NANDN U799 ( .A(B[401]), .B(n689), .Z(n688) );
  NANDN U800 ( .A(A[401]), .B(n690), .Z(n689) );
  NANDN U801 ( .A(n690), .B(A[401]), .Z(n687) );
  XOR U802 ( .A(n690), .B(n691), .Z(DIFF[401]) );
  XOR U803 ( .A(B[401]), .B(A[401]), .Z(n691) );
  AND U804 ( .A(n692), .B(n693), .Z(n690) );
  NANDN U805 ( .A(B[400]), .B(n694), .Z(n693) );
  NANDN U806 ( .A(A[400]), .B(n695), .Z(n694) );
  NANDN U807 ( .A(n695), .B(A[400]), .Z(n692) );
  XOR U808 ( .A(n695), .B(n696), .Z(DIFF[400]) );
  XOR U809 ( .A(B[400]), .B(A[400]), .Z(n696) );
  AND U810 ( .A(n697), .B(n698), .Z(n695) );
  NANDN U811 ( .A(B[399]), .B(n699), .Z(n698) );
  NANDN U812 ( .A(A[399]), .B(n700), .Z(n699) );
  NANDN U813 ( .A(n700), .B(A[399]), .Z(n697) );
  XOR U814 ( .A(n701), .B(n702), .Z(DIFF[3]) );
  XOR U815 ( .A(B[3]), .B(A[3]), .Z(n702) );
  XOR U816 ( .A(n703), .B(n704), .Z(DIFF[39]) );
  XOR U817 ( .A(B[39]), .B(A[39]), .Z(n704) );
  XOR U818 ( .A(n700), .B(n705), .Z(DIFF[399]) );
  XOR U819 ( .A(B[399]), .B(A[399]), .Z(n705) );
  AND U820 ( .A(n706), .B(n707), .Z(n700) );
  NANDN U821 ( .A(B[398]), .B(n708), .Z(n707) );
  NANDN U822 ( .A(A[398]), .B(n709), .Z(n708) );
  NANDN U823 ( .A(n709), .B(A[398]), .Z(n706) );
  XOR U824 ( .A(n709), .B(n710), .Z(DIFF[398]) );
  XOR U825 ( .A(B[398]), .B(A[398]), .Z(n710) );
  AND U826 ( .A(n711), .B(n712), .Z(n709) );
  NANDN U827 ( .A(B[397]), .B(n713), .Z(n712) );
  NANDN U828 ( .A(A[397]), .B(n714), .Z(n713) );
  NANDN U829 ( .A(n714), .B(A[397]), .Z(n711) );
  XOR U830 ( .A(n714), .B(n715), .Z(DIFF[397]) );
  XOR U831 ( .A(B[397]), .B(A[397]), .Z(n715) );
  AND U832 ( .A(n716), .B(n717), .Z(n714) );
  NANDN U833 ( .A(B[396]), .B(n718), .Z(n717) );
  NANDN U834 ( .A(A[396]), .B(n719), .Z(n718) );
  NANDN U835 ( .A(n719), .B(A[396]), .Z(n716) );
  XOR U836 ( .A(n719), .B(n720), .Z(DIFF[396]) );
  XOR U837 ( .A(B[396]), .B(A[396]), .Z(n720) );
  AND U838 ( .A(n721), .B(n722), .Z(n719) );
  NANDN U839 ( .A(B[395]), .B(n723), .Z(n722) );
  NANDN U840 ( .A(A[395]), .B(n724), .Z(n723) );
  NANDN U841 ( .A(n724), .B(A[395]), .Z(n721) );
  XOR U842 ( .A(n724), .B(n725), .Z(DIFF[395]) );
  XOR U843 ( .A(B[395]), .B(A[395]), .Z(n725) );
  AND U844 ( .A(n726), .B(n727), .Z(n724) );
  NANDN U845 ( .A(B[394]), .B(n728), .Z(n727) );
  NANDN U846 ( .A(A[394]), .B(n729), .Z(n728) );
  NANDN U847 ( .A(n729), .B(A[394]), .Z(n726) );
  XOR U848 ( .A(n729), .B(n730), .Z(DIFF[394]) );
  XOR U849 ( .A(B[394]), .B(A[394]), .Z(n730) );
  AND U850 ( .A(n731), .B(n732), .Z(n729) );
  NANDN U851 ( .A(B[393]), .B(n733), .Z(n732) );
  NANDN U852 ( .A(A[393]), .B(n734), .Z(n733) );
  NANDN U853 ( .A(n734), .B(A[393]), .Z(n731) );
  XOR U854 ( .A(n734), .B(n735), .Z(DIFF[393]) );
  XOR U855 ( .A(B[393]), .B(A[393]), .Z(n735) );
  AND U856 ( .A(n736), .B(n737), .Z(n734) );
  NANDN U857 ( .A(B[392]), .B(n738), .Z(n737) );
  NANDN U858 ( .A(A[392]), .B(n739), .Z(n738) );
  NANDN U859 ( .A(n739), .B(A[392]), .Z(n736) );
  XOR U860 ( .A(n739), .B(n740), .Z(DIFF[392]) );
  XOR U861 ( .A(B[392]), .B(A[392]), .Z(n740) );
  AND U862 ( .A(n741), .B(n742), .Z(n739) );
  NANDN U863 ( .A(B[391]), .B(n743), .Z(n742) );
  NANDN U864 ( .A(A[391]), .B(n744), .Z(n743) );
  NANDN U865 ( .A(n744), .B(A[391]), .Z(n741) );
  XOR U866 ( .A(n744), .B(n745), .Z(DIFF[391]) );
  XOR U867 ( .A(B[391]), .B(A[391]), .Z(n745) );
  AND U868 ( .A(n746), .B(n747), .Z(n744) );
  NANDN U869 ( .A(B[390]), .B(n748), .Z(n747) );
  NANDN U870 ( .A(A[390]), .B(n749), .Z(n748) );
  NANDN U871 ( .A(n749), .B(A[390]), .Z(n746) );
  XOR U872 ( .A(n749), .B(n750), .Z(DIFF[390]) );
  XOR U873 ( .A(B[390]), .B(A[390]), .Z(n750) );
  AND U874 ( .A(n751), .B(n752), .Z(n749) );
  NANDN U875 ( .A(B[389]), .B(n753), .Z(n752) );
  NANDN U876 ( .A(A[389]), .B(n754), .Z(n753) );
  NANDN U877 ( .A(n754), .B(A[389]), .Z(n751) );
  XOR U878 ( .A(n755), .B(n756), .Z(DIFF[38]) );
  XOR U879 ( .A(B[38]), .B(A[38]), .Z(n756) );
  XOR U880 ( .A(n754), .B(n757), .Z(DIFF[389]) );
  XOR U881 ( .A(B[389]), .B(A[389]), .Z(n757) );
  AND U882 ( .A(n758), .B(n759), .Z(n754) );
  NANDN U883 ( .A(B[388]), .B(n760), .Z(n759) );
  NANDN U884 ( .A(A[388]), .B(n761), .Z(n760) );
  NANDN U885 ( .A(n761), .B(A[388]), .Z(n758) );
  XOR U886 ( .A(n761), .B(n762), .Z(DIFF[388]) );
  XOR U887 ( .A(B[388]), .B(A[388]), .Z(n762) );
  AND U888 ( .A(n763), .B(n764), .Z(n761) );
  NANDN U889 ( .A(B[387]), .B(n765), .Z(n764) );
  NANDN U890 ( .A(A[387]), .B(n766), .Z(n765) );
  NANDN U891 ( .A(n766), .B(A[387]), .Z(n763) );
  XOR U892 ( .A(n766), .B(n767), .Z(DIFF[387]) );
  XOR U893 ( .A(B[387]), .B(A[387]), .Z(n767) );
  AND U894 ( .A(n768), .B(n769), .Z(n766) );
  NANDN U895 ( .A(B[386]), .B(n770), .Z(n769) );
  NANDN U896 ( .A(A[386]), .B(n771), .Z(n770) );
  NANDN U897 ( .A(n771), .B(A[386]), .Z(n768) );
  XOR U898 ( .A(n771), .B(n772), .Z(DIFF[386]) );
  XOR U899 ( .A(B[386]), .B(A[386]), .Z(n772) );
  AND U900 ( .A(n773), .B(n774), .Z(n771) );
  NANDN U901 ( .A(B[385]), .B(n775), .Z(n774) );
  NANDN U902 ( .A(A[385]), .B(n776), .Z(n775) );
  NANDN U903 ( .A(n776), .B(A[385]), .Z(n773) );
  XOR U904 ( .A(n776), .B(n777), .Z(DIFF[385]) );
  XOR U905 ( .A(B[385]), .B(A[385]), .Z(n777) );
  AND U906 ( .A(n778), .B(n779), .Z(n776) );
  NANDN U907 ( .A(B[384]), .B(n780), .Z(n779) );
  NANDN U908 ( .A(A[384]), .B(n781), .Z(n780) );
  NANDN U909 ( .A(n781), .B(A[384]), .Z(n778) );
  XOR U910 ( .A(n781), .B(n782), .Z(DIFF[384]) );
  XOR U911 ( .A(B[384]), .B(A[384]), .Z(n782) );
  AND U912 ( .A(n783), .B(n784), .Z(n781) );
  NANDN U913 ( .A(B[383]), .B(n785), .Z(n784) );
  NANDN U914 ( .A(A[383]), .B(n786), .Z(n785) );
  NANDN U915 ( .A(n786), .B(A[383]), .Z(n783) );
  XOR U916 ( .A(n786), .B(n787), .Z(DIFF[383]) );
  XOR U917 ( .A(B[383]), .B(A[383]), .Z(n787) );
  AND U918 ( .A(n788), .B(n789), .Z(n786) );
  NANDN U919 ( .A(B[382]), .B(n790), .Z(n789) );
  NANDN U920 ( .A(A[382]), .B(n791), .Z(n790) );
  NANDN U921 ( .A(n791), .B(A[382]), .Z(n788) );
  XOR U922 ( .A(n791), .B(n792), .Z(DIFF[382]) );
  XOR U923 ( .A(B[382]), .B(A[382]), .Z(n792) );
  AND U924 ( .A(n793), .B(n794), .Z(n791) );
  NANDN U925 ( .A(B[381]), .B(n795), .Z(n794) );
  NANDN U926 ( .A(A[381]), .B(n796), .Z(n795) );
  NANDN U927 ( .A(n796), .B(A[381]), .Z(n793) );
  XOR U928 ( .A(n796), .B(n797), .Z(DIFF[381]) );
  XOR U929 ( .A(B[381]), .B(A[381]), .Z(n797) );
  AND U930 ( .A(n798), .B(n799), .Z(n796) );
  NANDN U931 ( .A(B[380]), .B(n800), .Z(n799) );
  NANDN U932 ( .A(A[380]), .B(n801), .Z(n800) );
  NANDN U933 ( .A(n801), .B(A[380]), .Z(n798) );
  XOR U934 ( .A(n801), .B(n802), .Z(DIFF[380]) );
  XOR U935 ( .A(B[380]), .B(A[380]), .Z(n802) );
  AND U936 ( .A(n803), .B(n804), .Z(n801) );
  NANDN U937 ( .A(B[379]), .B(n805), .Z(n804) );
  NANDN U938 ( .A(A[379]), .B(n806), .Z(n805) );
  NANDN U939 ( .A(n806), .B(A[379]), .Z(n803) );
  XOR U940 ( .A(n807), .B(n808), .Z(DIFF[37]) );
  XOR U941 ( .A(B[37]), .B(A[37]), .Z(n808) );
  XOR U942 ( .A(n806), .B(n809), .Z(DIFF[379]) );
  XOR U943 ( .A(B[379]), .B(A[379]), .Z(n809) );
  AND U944 ( .A(n810), .B(n811), .Z(n806) );
  NANDN U945 ( .A(B[378]), .B(n812), .Z(n811) );
  NANDN U946 ( .A(A[378]), .B(n813), .Z(n812) );
  NANDN U947 ( .A(n813), .B(A[378]), .Z(n810) );
  XOR U948 ( .A(n813), .B(n814), .Z(DIFF[378]) );
  XOR U949 ( .A(B[378]), .B(A[378]), .Z(n814) );
  AND U950 ( .A(n815), .B(n816), .Z(n813) );
  NANDN U951 ( .A(B[377]), .B(n817), .Z(n816) );
  NANDN U952 ( .A(A[377]), .B(n818), .Z(n817) );
  NANDN U953 ( .A(n818), .B(A[377]), .Z(n815) );
  XOR U954 ( .A(n818), .B(n819), .Z(DIFF[377]) );
  XOR U955 ( .A(B[377]), .B(A[377]), .Z(n819) );
  AND U956 ( .A(n820), .B(n821), .Z(n818) );
  NANDN U957 ( .A(B[376]), .B(n822), .Z(n821) );
  NANDN U958 ( .A(A[376]), .B(n823), .Z(n822) );
  NANDN U959 ( .A(n823), .B(A[376]), .Z(n820) );
  XOR U960 ( .A(n823), .B(n824), .Z(DIFF[376]) );
  XOR U961 ( .A(B[376]), .B(A[376]), .Z(n824) );
  AND U962 ( .A(n825), .B(n826), .Z(n823) );
  NANDN U963 ( .A(B[375]), .B(n827), .Z(n826) );
  NANDN U964 ( .A(A[375]), .B(n828), .Z(n827) );
  NANDN U965 ( .A(n828), .B(A[375]), .Z(n825) );
  XOR U966 ( .A(n828), .B(n829), .Z(DIFF[375]) );
  XOR U967 ( .A(B[375]), .B(A[375]), .Z(n829) );
  AND U968 ( .A(n830), .B(n831), .Z(n828) );
  NANDN U969 ( .A(B[374]), .B(n832), .Z(n831) );
  NANDN U970 ( .A(A[374]), .B(n833), .Z(n832) );
  NANDN U971 ( .A(n833), .B(A[374]), .Z(n830) );
  XOR U972 ( .A(n833), .B(n834), .Z(DIFF[374]) );
  XOR U973 ( .A(B[374]), .B(A[374]), .Z(n834) );
  AND U974 ( .A(n835), .B(n836), .Z(n833) );
  NANDN U975 ( .A(B[373]), .B(n837), .Z(n836) );
  NANDN U976 ( .A(A[373]), .B(n838), .Z(n837) );
  NANDN U977 ( .A(n838), .B(A[373]), .Z(n835) );
  XOR U978 ( .A(n838), .B(n839), .Z(DIFF[373]) );
  XOR U979 ( .A(B[373]), .B(A[373]), .Z(n839) );
  AND U980 ( .A(n840), .B(n841), .Z(n838) );
  NANDN U981 ( .A(B[372]), .B(n842), .Z(n841) );
  NANDN U982 ( .A(A[372]), .B(n843), .Z(n842) );
  NANDN U983 ( .A(n843), .B(A[372]), .Z(n840) );
  XOR U984 ( .A(n843), .B(n844), .Z(DIFF[372]) );
  XOR U985 ( .A(B[372]), .B(A[372]), .Z(n844) );
  AND U986 ( .A(n845), .B(n846), .Z(n843) );
  NANDN U987 ( .A(B[371]), .B(n847), .Z(n846) );
  NANDN U988 ( .A(A[371]), .B(n848), .Z(n847) );
  NANDN U989 ( .A(n848), .B(A[371]), .Z(n845) );
  XOR U990 ( .A(n848), .B(n849), .Z(DIFF[371]) );
  XOR U991 ( .A(B[371]), .B(A[371]), .Z(n849) );
  AND U992 ( .A(n850), .B(n851), .Z(n848) );
  NANDN U993 ( .A(B[370]), .B(n852), .Z(n851) );
  NANDN U994 ( .A(A[370]), .B(n853), .Z(n852) );
  NANDN U995 ( .A(n853), .B(A[370]), .Z(n850) );
  XOR U996 ( .A(n853), .B(n854), .Z(DIFF[370]) );
  XOR U997 ( .A(B[370]), .B(A[370]), .Z(n854) );
  AND U998 ( .A(n855), .B(n856), .Z(n853) );
  NANDN U999 ( .A(B[369]), .B(n857), .Z(n856) );
  NANDN U1000 ( .A(A[369]), .B(n858), .Z(n857) );
  NANDN U1001 ( .A(n858), .B(A[369]), .Z(n855) );
  XOR U1002 ( .A(n859), .B(n860), .Z(DIFF[36]) );
  XOR U1003 ( .A(B[36]), .B(A[36]), .Z(n860) );
  XOR U1004 ( .A(n858), .B(n861), .Z(DIFF[369]) );
  XOR U1005 ( .A(B[369]), .B(A[369]), .Z(n861) );
  AND U1006 ( .A(n862), .B(n863), .Z(n858) );
  NANDN U1007 ( .A(B[368]), .B(n864), .Z(n863) );
  NANDN U1008 ( .A(A[368]), .B(n865), .Z(n864) );
  NANDN U1009 ( .A(n865), .B(A[368]), .Z(n862) );
  XOR U1010 ( .A(n865), .B(n866), .Z(DIFF[368]) );
  XOR U1011 ( .A(B[368]), .B(A[368]), .Z(n866) );
  AND U1012 ( .A(n867), .B(n868), .Z(n865) );
  NANDN U1013 ( .A(B[367]), .B(n869), .Z(n868) );
  NANDN U1014 ( .A(A[367]), .B(n870), .Z(n869) );
  NANDN U1015 ( .A(n870), .B(A[367]), .Z(n867) );
  XOR U1016 ( .A(n870), .B(n871), .Z(DIFF[367]) );
  XOR U1017 ( .A(B[367]), .B(A[367]), .Z(n871) );
  AND U1018 ( .A(n872), .B(n873), .Z(n870) );
  NANDN U1019 ( .A(B[366]), .B(n874), .Z(n873) );
  NANDN U1020 ( .A(A[366]), .B(n875), .Z(n874) );
  NANDN U1021 ( .A(n875), .B(A[366]), .Z(n872) );
  XOR U1022 ( .A(n875), .B(n876), .Z(DIFF[366]) );
  XOR U1023 ( .A(B[366]), .B(A[366]), .Z(n876) );
  AND U1024 ( .A(n877), .B(n878), .Z(n875) );
  NANDN U1025 ( .A(B[365]), .B(n879), .Z(n878) );
  NANDN U1026 ( .A(A[365]), .B(n880), .Z(n879) );
  NANDN U1027 ( .A(n880), .B(A[365]), .Z(n877) );
  XOR U1028 ( .A(n880), .B(n881), .Z(DIFF[365]) );
  XOR U1029 ( .A(B[365]), .B(A[365]), .Z(n881) );
  AND U1030 ( .A(n882), .B(n883), .Z(n880) );
  NANDN U1031 ( .A(B[364]), .B(n884), .Z(n883) );
  NANDN U1032 ( .A(A[364]), .B(n885), .Z(n884) );
  NANDN U1033 ( .A(n885), .B(A[364]), .Z(n882) );
  XOR U1034 ( .A(n885), .B(n886), .Z(DIFF[364]) );
  XOR U1035 ( .A(B[364]), .B(A[364]), .Z(n886) );
  AND U1036 ( .A(n887), .B(n888), .Z(n885) );
  NANDN U1037 ( .A(B[363]), .B(n889), .Z(n888) );
  NANDN U1038 ( .A(A[363]), .B(n890), .Z(n889) );
  NANDN U1039 ( .A(n890), .B(A[363]), .Z(n887) );
  XOR U1040 ( .A(n890), .B(n891), .Z(DIFF[363]) );
  XOR U1041 ( .A(B[363]), .B(A[363]), .Z(n891) );
  AND U1042 ( .A(n892), .B(n893), .Z(n890) );
  NANDN U1043 ( .A(B[362]), .B(n894), .Z(n893) );
  NANDN U1044 ( .A(A[362]), .B(n895), .Z(n894) );
  NANDN U1045 ( .A(n895), .B(A[362]), .Z(n892) );
  XOR U1046 ( .A(n895), .B(n896), .Z(DIFF[362]) );
  XOR U1047 ( .A(B[362]), .B(A[362]), .Z(n896) );
  AND U1048 ( .A(n897), .B(n898), .Z(n895) );
  NANDN U1049 ( .A(B[361]), .B(n899), .Z(n898) );
  NANDN U1050 ( .A(A[361]), .B(n900), .Z(n899) );
  NANDN U1051 ( .A(n900), .B(A[361]), .Z(n897) );
  XOR U1052 ( .A(n900), .B(n901), .Z(DIFF[361]) );
  XOR U1053 ( .A(B[361]), .B(A[361]), .Z(n901) );
  AND U1054 ( .A(n902), .B(n903), .Z(n900) );
  NANDN U1055 ( .A(B[360]), .B(n904), .Z(n903) );
  NANDN U1056 ( .A(A[360]), .B(n905), .Z(n904) );
  NANDN U1057 ( .A(n905), .B(A[360]), .Z(n902) );
  XOR U1058 ( .A(n905), .B(n906), .Z(DIFF[360]) );
  XOR U1059 ( .A(B[360]), .B(A[360]), .Z(n906) );
  AND U1060 ( .A(n907), .B(n908), .Z(n905) );
  NANDN U1061 ( .A(B[359]), .B(n909), .Z(n908) );
  NANDN U1062 ( .A(A[359]), .B(n910), .Z(n909) );
  NANDN U1063 ( .A(n910), .B(A[359]), .Z(n907) );
  XOR U1064 ( .A(n911), .B(n912), .Z(DIFF[35]) );
  XOR U1065 ( .A(B[35]), .B(A[35]), .Z(n912) );
  XOR U1066 ( .A(n910), .B(n913), .Z(DIFF[359]) );
  XOR U1067 ( .A(B[359]), .B(A[359]), .Z(n913) );
  AND U1068 ( .A(n914), .B(n915), .Z(n910) );
  NANDN U1069 ( .A(B[358]), .B(n916), .Z(n915) );
  NANDN U1070 ( .A(A[358]), .B(n917), .Z(n916) );
  NANDN U1071 ( .A(n917), .B(A[358]), .Z(n914) );
  XOR U1072 ( .A(n917), .B(n918), .Z(DIFF[358]) );
  XOR U1073 ( .A(B[358]), .B(A[358]), .Z(n918) );
  AND U1074 ( .A(n919), .B(n920), .Z(n917) );
  NANDN U1075 ( .A(B[357]), .B(n921), .Z(n920) );
  NANDN U1076 ( .A(A[357]), .B(n922), .Z(n921) );
  NANDN U1077 ( .A(n922), .B(A[357]), .Z(n919) );
  XOR U1078 ( .A(n922), .B(n923), .Z(DIFF[357]) );
  XOR U1079 ( .A(B[357]), .B(A[357]), .Z(n923) );
  AND U1080 ( .A(n924), .B(n925), .Z(n922) );
  NANDN U1081 ( .A(B[356]), .B(n926), .Z(n925) );
  NANDN U1082 ( .A(A[356]), .B(n927), .Z(n926) );
  NANDN U1083 ( .A(n927), .B(A[356]), .Z(n924) );
  XOR U1084 ( .A(n927), .B(n928), .Z(DIFF[356]) );
  XOR U1085 ( .A(B[356]), .B(A[356]), .Z(n928) );
  AND U1086 ( .A(n929), .B(n930), .Z(n927) );
  NANDN U1087 ( .A(B[355]), .B(n931), .Z(n930) );
  NANDN U1088 ( .A(A[355]), .B(n932), .Z(n931) );
  NANDN U1089 ( .A(n932), .B(A[355]), .Z(n929) );
  XOR U1090 ( .A(n932), .B(n933), .Z(DIFF[355]) );
  XOR U1091 ( .A(B[355]), .B(A[355]), .Z(n933) );
  AND U1092 ( .A(n934), .B(n935), .Z(n932) );
  NANDN U1093 ( .A(B[354]), .B(n936), .Z(n935) );
  NANDN U1094 ( .A(A[354]), .B(n937), .Z(n936) );
  NANDN U1095 ( .A(n937), .B(A[354]), .Z(n934) );
  XOR U1096 ( .A(n937), .B(n938), .Z(DIFF[354]) );
  XOR U1097 ( .A(B[354]), .B(A[354]), .Z(n938) );
  AND U1098 ( .A(n939), .B(n940), .Z(n937) );
  NANDN U1099 ( .A(B[353]), .B(n941), .Z(n940) );
  NANDN U1100 ( .A(A[353]), .B(n942), .Z(n941) );
  NANDN U1101 ( .A(n942), .B(A[353]), .Z(n939) );
  XOR U1102 ( .A(n942), .B(n943), .Z(DIFF[353]) );
  XOR U1103 ( .A(B[353]), .B(A[353]), .Z(n943) );
  AND U1104 ( .A(n944), .B(n945), .Z(n942) );
  NANDN U1105 ( .A(B[352]), .B(n946), .Z(n945) );
  NANDN U1106 ( .A(A[352]), .B(n947), .Z(n946) );
  NANDN U1107 ( .A(n947), .B(A[352]), .Z(n944) );
  XOR U1108 ( .A(n947), .B(n948), .Z(DIFF[352]) );
  XOR U1109 ( .A(B[352]), .B(A[352]), .Z(n948) );
  AND U1110 ( .A(n949), .B(n950), .Z(n947) );
  NANDN U1111 ( .A(B[351]), .B(n951), .Z(n950) );
  NANDN U1112 ( .A(A[351]), .B(n952), .Z(n951) );
  NANDN U1113 ( .A(n952), .B(A[351]), .Z(n949) );
  XOR U1114 ( .A(n952), .B(n953), .Z(DIFF[351]) );
  XOR U1115 ( .A(B[351]), .B(A[351]), .Z(n953) );
  AND U1116 ( .A(n954), .B(n955), .Z(n952) );
  NANDN U1117 ( .A(B[350]), .B(n956), .Z(n955) );
  NANDN U1118 ( .A(A[350]), .B(n957), .Z(n956) );
  NANDN U1119 ( .A(n957), .B(A[350]), .Z(n954) );
  XOR U1120 ( .A(n957), .B(n958), .Z(DIFF[350]) );
  XOR U1121 ( .A(B[350]), .B(A[350]), .Z(n958) );
  AND U1122 ( .A(n959), .B(n960), .Z(n957) );
  NANDN U1123 ( .A(B[349]), .B(n961), .Z(n960) );
  NANDN U1124 ( .A(A[349]), .B(n962), .Z(n961) );
  NANDN U1125 ( .A(n962), .B(A[349]), .Z(n959) );
  XOR U1126 ( .A(n963), .B(n964), .Z(DIFF[34]) );
  XOR U1127 ( .A(B[34]), .B(A[34]), .Z(n964) );
  XOR U1128 ( .A(n962), .B(n965), .Z(DIFF[349]) );
  XOR U1129 ( .A(B[349]), .B(A[349]), .Z(n965) );
  AND U1130 ( .A(n966), .B(n967), .Z(n962) );
  NANDN U1131 ( .A(B[348]), .B(n968), .Z(n967) );
  NANDN U1132 ( .A(A[348]), .B(n969), .Z(n968) );
  NANDN U1133 ( .A(n969), .B(A[348]), .Z(n966) );
  XOR U1134 ( .A(n969), .B(n970), .Z(DIFF[348]) );
  XOR U1135 ( .A(B[348]), .B(A[348]), .Z(n970) );
  AND U1136 ( .A(n971), .B(n972), .Z(n969) );
  NANDN U1137 ( .A(B[347]), .B(n973), .Z(n972) );
  NANDN U1138 ( .A(A[347]), .B(n974), .Z(n973) );
  NANDN U1139 ( .A(n974), .B(A[347]), .Z(n971) );
  XOR U1140 ( .A(n974), .B(n975), .Z(DIFF[347]) );
  XOR U1141 ( .A(B[347]), .B(A[347]), .Z(n975) );
  AND U1142 ( .A(n976), .B(n977), .Z(n974) );
  NANDN U1143 ( .A(B[346]), .B(n978), .Z(n977) );
  NANDN U1144 ( .A(A[346]), .B(n979), .Z(n978) );
  NANDN U1145 ( .A(n979), .B(A[346]), .Z(n976) );
  XOR U1146 ( .A(n979), .B(n980), .Z(DIFF[346]) );
  XOR U1147 ( .A(B[346]), .B(A[346]), .Z(n980) );
  AND U1148 ( .A(n981), .B(n982), .Z(n979) );
  NANDN U1149 ( .A(B[345]), .B(n983), .Z(n982) );
  NANDN U1150 ( .A(A[345]), .B(n984), .Z(n983) );
  NANDN U1151 ( .A(n984), .B(A[345]), .Z(n981) );
  XOR U1152 ( .A(n984), .B(n985), .Z(DIFF[345]) );
  XOR U1153 ( .A(B[345]), .B(A[345]), .Z(n985) );
  AND U1154 ( .A(n986), .B(n987), .Z(n984) );
  NANDN U1155 ( .A(B[344]), .B(n988), .Z(n987) );
  NANDN U1156 ( .A(A[344]), .B(n989), .Z(n988) );
  NANDN U1157 ( .A(n989), .B(A[344]), .Z(n986) );
  XOR U1158 ( .A(n989), .B(n990), .Z(DIFF[344]) );
  XOR U1159 ( .A(B[344]), .B(A[344]), .Z(n990) );
  AND U1160 ( .A(n991), .B(n992), .Z(n989) );
  NANDN U1161 ( .A(B[343]), .B(n993), .Z(n992) );
  NANDN U1162 ( .A(A[343]), .B(n994), .Z(n993) );
  NANDN U1163 ( .A(n994), .B(A[343]), .Z(n991) );
  XOR U1164 ( .A(n994), .B(n995), .Z(DIFF[343]) );
  XOR U1165 ( .A(B[343]), .B(A[343]), .Z(n995) );
  AND U1166 ( .A(n996), .B(n997), .Z(n994) );
  NANDN U1167 ( .A(B[342]), .B(n998), .Z(n997) );
  NANDN U1168 ( .A(A[342]), .B(n999), .Z(n998) );
  NANDN U1169 ( .A(n999), .B(A[342]), .Z(n996) );
  XOR U1170 ( .A(n999), .B(n1000), .Z(DIFF[342]) );
  XOR U1171 ( .A(B[342]), .B(A[342]), .Z(n1000) );
  AND U1172 ( .A(n1001), .B(n1002), .Z(n999) );
  NANDN U1173 ( .A(B[341]), .B(n1003), .Z(n1002) );
  NANDN U1174 ( .A(A[341]), .B(n1004), .Z(n1003) );
  NANDN U1175 ( .A(n1004), .B(A[341]), .Z(n1001) );
  XOR U1176 ( .A(n1004), .B(n1005), .Z(DIFF[341]) );
  XOR U1177 ( .A(B[341]), .B(A[341]), .Z(n1005) );
  AND U1178 ( .A(n1006), .B(n1007), .Z(n1004) );
  NANDN U1179 ( .A(B[340]), .B(n1008), .Z(n1007) );
  NANDN U1180 ( .A(A[340]), .B(n1009), .Z(n1008) );
  NANDN U1181 ( .A(n1009), .B(A[340]), .Z(n1006) );
  XOR U1182 ( .A(n1009), .B(n1010), .Z(DIFF[340]) );
  XOR U1183 ( .A(B[340]), .B(A[340]), .Z(n1010) );
  AND U1184 ( .A(n1011), .B(n1012), .Z(n1009) );
  NANDN U1185 ( .A(B[339]), .B(n1013), .Z(n1012) );
  NANDN U1186 ( .A(A[339]), .B(n1014), .Z(n1013) );
  NANDN U1187 ( .A(n1014), .B(A[339]), .Z(n1011) );
  XOR U1188 ( .A(n1015), .B(n1016), .Z(DIFF[33]) );
  XOR U1189 ( .A(B[33]), .B(A[33]), .Z(n1016) );
  XOR U1190 ( .A(n1014), .B(n1017), .Z(DIFF[339]) );
  XOR U1191 ( .A(B[339]), .B(A[339]), .Z(n1017) );
  AND U1192 ( .A(n1018), .B(n1019), .Z(n1014) );
  NANDN U1193 ( .A(B[338]), .B(n1020), .Z(n1019) );
  NANDN U1194 ( .A(A[338]), .B(n1021), .Z(n1020) );
  NANDN U1195 ( .A(n1021), .B(A[338]), .Z(n1018) );
  XOR U1196 ( .A(n1021), .B(n1022), .Z(DIFF[338]) );
  XOR U1197 ( .A(B[338]), .B(A[338]), .Z(n1022) );
  AND U1198 ( .A(n1023), .B(n1024), .Z(n1021) );
  NANDN U1199 ( .A(B[337]), .B(n1025), .Z(n1024) );
  NANDN U1200 ( .A(A[337]), .B(n1026), .Z(n1025) );
  NANDN U1201 ( .A(n1026), .B(A[337]), .Z(n1023) );
  XOR U1202 ( .A(n1026), .B(n1027), .Z(DIFF[337]) );
  XOR U1203 ( .A(B[337]), .B(A[337]), .Z(n1027) );
  AND U1204 ( .A(n1028), .B(n1029), .Z(n1026) );
  NANDN U1205 ( .A(B[336]), .B(n1030), .Z(n1029) );
  NANDN U1206 ( .A(A[336]), .B(n1031), .Z(n1030) );
  NANDN U1207 ( .A(n1031), .B(A[336]), .Z(n1028) );
  XOR U1208 ( .A(n1031), .B(n1032), .Z(DIFF[336]) );
  XOR U1209 ( .A(B[336]), .B(A[336]), .Z(n1032) );
  AND U1210 ( .A(n1033), .B(n1034), .Z(n1031) );
  NANDN U1211 ( .A(B[335]), .B(n1035), .Z(n1034) );
  NANDN U1212 ( .A(A[335]), .B(n1036), .Z(n1035) );
  NANDN U1213 ( .A(n1036), .B(A[335]), .Z(n1033) );
  XOR U1214 ( .A(n1036), .B(n1037), .Z(DIFF[335]) );
  XOR U1215 ( .A(B[335]), .B(A[335]), .Z(n1037) );
  AND U1216 ( .A(n1038), .B(n1039), .Z(n1036) );
  NANDN U1217 ( .A(B[334]), .B(n1040), .Z(n1039) );
  NANDN U1218 ( .A(A[334]), .B(n1041), .Z(n1040) );
  NANDN U1219 ( .A(n1041), .B(A[334]), .Z(n1038) );
  XOR U1220 ( .A(n1041), .B(n1042), .Z(DIFF[334]) );
  XOR U1221 ( .A(B[334]), .B(A[334]), .Z(n1042) );
  AND U1222 ( .A(n1043), .B(n1044), .Z(n1041) );
  NANDN U1223 ( .A(B[333]), .B(n1045), .Z(n1044) );
  NANDN U1224 ( .A(A[333]), .B(n1046), .Z(n1045) );
  NANDN U1225 ( .A(n1046), .B(A[333]), .Z(n1043) );
  XOR U1226 ( .A(n1046), .B(n1047), .Z(DIFF[333]) );
  XOR U1227 ( .A(B[333]), .B(A[333]), .Z(n1047) );
  AND U1228 ( .A(n1048), .B(n1049), .Z(n1046) );
  NANDN U1229 ( .A(B[332]), .B(n1050), .Z(n1049) );
  NANDN U1230 ( .A(A[332]), .B(n1051), .Z(n1050) );
  NANDN U1231 ( .A(n1051), .B(A[332]), .Z(n1048) );
  XOR U1232 ( .A(n1051), .B(n1052), .Z(DIFF[332]) );
  XOR U1233 ( .A(B[332]), .B(A[332]), .Z(n1052) );
  AND U1234 ( .A(n1053), .B(n1054), .Z(n1051) );
  NANDN U1235 ( .A(B[331]), .B(n1055), .Z(n1054) );
  NANDN U1236 ( .A(A[331]), .B(n1056), .Z(n1055) );
  NANDN U1237 ( .A(n1056), .B(A[331]), .Z(n1053) );
  XOR U1238 ( .A(n1056), .B(n1057), .Z(DIFF[331]) );
  XOR U1239 ( .A(B[331]), .B(A[331]), .Z(n1057) );
  AND U1240 ( .A(n1058), .B(n1059), .Z(n1056) );
  NANDN U1241 ( .A(B[330]), .B(n1060), .Z(n1059) );
  NANDN U1242 ( .A(A[330]), .B(n1061), .Z(n1060) );
  NANDN U1243 ( .A(n1061), .B(A[330]), .Z(n1058) );
  XOR U1244 ( .A(n1061), .B(n1062), .Z(DIFF[330]) );
  XOR U1245 ( .A(B[330]), .B(A[330]), .Z(n1062) );
  AND U1246 ( .A(n1063), .B(n1064), .Z(n1061) );
  NANDN U1247 ( .A(B[329]), .B(n1065), .Z(n1064) );
  NANDN U1248 ( .A(A[329]), .B(n1066), .Z(n1065) );
  NANDN U1249 ( .A(n1066), .B(A[329]), .Z(n1063) );
  XOR U1250 ( .A(n1067), .B(n1068), .Z(DIFF[32]) );
  XOR U1251 ( .A(B[32]), .B(A[32]), .Z(n1068) );
  XOR U1252 ( .A(n1066), .B(n1069), .Z(DIFF[329]) );
  XOR U1253 ( .A(B[329]), .B(A[329]), .Z(n1069) );
  AND U1254 ( .A(n1070), .B(n1071), .Z(n1066) );
  NANDN U1255 ( .A(B[328]), .B(n1072), .Z(n1071) );
  NANDN U1256 ( .A(A[328]), .B(n1073), .Z(n1072) );
  NANDN U1257 ( .A(n1073), .B(A[328]), .Z(n1070) );
  XOR U1258 ( .A(n1073), .B(n1074), .Z(DIFF[328]) );
  XOR U1259 ( .A(B[328]), .B(A[328]), .Z(n1074) );
  AND U1260 ( .A(n1075), .B(n1076), .Z(n1073) );
  NANDN U1261 ( .A(B[327]), .B(n1077), .Z(n1076) );
  NANDN U1262 ( .A(A[327]), .B(n1078), .Z(n1077) );
  NANDN U1263 ( .A(n1078), .B(A[327]), .Z(n1075) );
  XOR U1264 ( .A(n1078), .B(n1079), .Z(DIFF[327]) );
  XOR U1265 ( .A(B[327]), .B(A[327]), .Z(n1079) );
  AND U1266 ( .A(n1080), .B(n1081), .Z(n1078) );
  NANDN U1267 ( .A(B[326]), .B(n1082), .Z(n1081) );
  NANDN U1268 ( .A(A[326]), .B(n1083), .Z(n1082) );
  NANDN U1269 ( .A(n1083), .B(A[326]), .Z(n1080) );
  XOR U1270 ( .A(n1083), .B(n1084), .Z(DIFF[326]) );
  XOR U1271 ( .A(B[326]), .B(A[326]), .Z(n1084) );
  AND U1272 ( .A(n1085), .B(n1086), .Z(n1083) );
  NANDN U1273 ( .A(B[325]), .B(n1087), .Z(n1086) );
  NANDN U1274 ( .A(A[325]), .B(n1088), .Z(n1087) );
  NANDN U1275 ( .A(n1088), .B(A[325]), .Z(n1085) );
  XOR U1276 ( .A(n1088), .B(n1089), .Z(DIFF[325]) );
  XOR U1277 ( .A(B[325]), .B(A[325]), .Z(n1089) );
  AND U1278 ( .A(n1090), .B(n1091), .Z(n1088) );
  NANDN U1279 ( .A(B[324]), .B(n1092), .Z(n1091) );
  NANDN U1280 ( .A(A[324]), .B(n1093), .Z(n1092) );
  NANDN U1281 ( .A(n1093), .B(A[324]), .Z(n1090) );
  XOR U1282 ( .A(n1093), .B(n1094), .Z(DIFF[324]) );
  XOR U1283 ( .A(B[324]), .B(A[324]), .Z(n1094) );
  AND U1284 ( .A(n1095), .B(n1096), .Z(n1093) );
  NANDN U1285 ( .A(B[323]), .B(n1097), .Z(n1096) );
  NANDN U1286 ( .A(A[323]), .B(n1098), .Z(n1097) );
  NANDN U1287 ( .A(n1098), .B(A[323]), .Z(n1095) );
  XOR U1288 ( .A(n1098), .B(n1099), .Z(DIFF[323]) );
  XOR U1289 ( .A(B[323]), .B(A[323]), .Z(n1099) );
  AND U1290 ( .A(n1100), .B(n1101), .Z(n1098) );
  NANDN U1291 ( .A(B[322]), .B(n1102), .Z(n1101) );
  NANDN U1292 ( .A(A[322]), .B(n1103), .Z(n1102) );
  NANDN U1293 ( .A(n1103), .B(A[322]), .Z(n1100) );
  XOR U1294 ( .A(n1103), .B(n1104), .Z(DIFF[322]) );
  XOR U1295 ( .A(B[322]), .B(A[322]), .Z(n1104) );
  AND U1296 ( .A(n1105), .B(n1106), .Z(n1103) );
  NANDN U1297 ( .A(B[321]), .B(n1107), .Z(n1106) );
  NANDN U1298 ( .A(A[321]), .B(n1108), .Z(n1107) );
  NANDN U1299 ( .A(n1108), .B(A[321]), .Z(n1105) );
  XOR U1300 ( .A(n1108), .B(n1109), .Z(DIFF[321]) );
  XOR U1301 ( .A(B[321]), .B(A[321]), .Z(n1109) );
  AND U1302 ( .A(n1110), .B(n1111), .Z(n1108) );
  NANDN U1303 ( .A(B[320]), .B(n1112), .Z(n1111) );
  NANDN U1304 ( .A(A[320]), .B(n1113), .Z(n1112) );
  NANDN U1305 ( .A(n1113), .B(A[320]), .Z(n1110) );
  XOR U1306 ( .A(n1113), .B(n1114), .Z(DIFF[320]) );
  XOR U1307 ( .A(B[320]), .B(A[320]), .Z(n1114) );
  AND U1308 ( .A(n1115), .B(n1116), .Z(n1113) );
  NANDN U1309 ( .A(B[319]), .B(n1117), .Z(n1116) );
  NANDN U1310 ( .A(A[319]), .B(n1118), .Z(n1117) );
  NANDN U1311 ( .A(n1118), .B(A[319]), .Z(n1115) );
  XOR U1312 ( .A(n1119), .B(n1120), .Z(DIFF[31]) );
  XOR U1313 ( .A(B[31]), .B(A[31]), .Z(n1120) );
  XOR U1314 ( .A(n1118), .B(n1121), .Z(DIFF[319]) );
  XOR U1315 ( .A(B[319]), .B(A[319]), .Z(n1121) );
  AND U1316 ( .A(n1122), .B(n1123), .Z(n1118) );
  NANDN U1317 ( .A(B[318]), .B(n1124), .Z(n1123) );
  NANDN U1318 ( .A(A[318]), .B(n1125), .Z(n1124) );
  NANDN U1319 ( .A(n1125), .B(A[318]), .Z(n1122) );
  XOR U1320 ( .A(n1125), .B(n1126), .Z(DIFF[318]) );
  XOR U1321 ( .A(B[318]), .B(A[318]), .Z(n1126) );
  AND U1322 ( .A(n1127), .B(n1128), .Z(n1125) );
  NANDN U1323 ( .A(B[317]), .B(n1129), .Z(n1128) );
  NANDN U1324 ( .A(A[317]), .B(n1130), .Z(n1129) );
  NANDN U1325 ( .A(n1130), .B(A[317]), .Z(n1127) );
  XOR U1326 ( .A(n1130), .B(n1131), .Z(DIFF[317]) );
  XOR U1327 ( .A(B[317]), .B(A[317]), .Z(n1131) );
  AND U1328 ( .A(n1132), .B(n1133), .Z(n1130) );
  NANDN U1329 ( .A(B[316]), .B(n1134), .Z(n1133) );
  NANDN U1330 ( .A(A[316]), .B(n1135), .Z(n1134) );
  NANDN U1331 ( .A(n1135), .B(A[316]), .Z(n1132) );
  XOR U1332 ( .A(n1135), .B(n1136), .Z(DIFF[316]) );
  XOR U1333 ( .A(B[316]), .B(A[316]), .Z(n1136) );
  AND U1334 ( .A(n1137), .B(n1138), .Z(n1135) );
  NANDN U1335 ( .A(B[315]), .B(n1139), .Z(n1138) );
  NANDN U1336 ( .A(A[315]), .B(n1140), .Z(n1139) );
  NANDN U1337 ( .A(n1140), .B(A[315]), .Z(n1137) );
  XOR U1338 ( .A(n1140), .B(n1141), .Z(DIFF[315]) );
  XOR U1339 ( .A(B[315]), .B(A[315]), .Z(n1141) );
  AND U1340 ( .A(n1142), .B(n1143), .Z(n1140) );
  NANDN U1341 ( .A(B[314]), .B(n1144), .Z(n1143) );
  NANDN U1342 ( .A(A[314]), .B(n1145), .Z(n1144) );
  NANDN U1343 ( .A(n1145), .B(A[314]), .Z(n1142) );
  XOR U1344 ( .A(n1145), .B(n1146), .Z(DIFF[314]) );
  XOR U1345 ( .A(B[314]), .B(A[314]), .Z(n1146) );
  AND U1346 ( .A(n1147), .B(n1148), .Z(n1145) );
  NANDN U1347 ( .A(B[313]), .B(n1149), .Z(n1148) );
  NANDN U1348 ( .A(A[313]), .B(n1150), .Z(n1149) );
  NANDN U1349 ( .A(n1150), .B(A[313]), .Z(n1147) );
  XOR U1350 ( .A(n1150), .B(n1151), .Z(DIFF[313]) );
  XOR U1351 ( .A(B[313]), .B(A[313]), .Z(n1151) );
  AND U1352 ( .A(n1152), .B(n1153), .Z(n1150) );
  NANDN U1353 ( .A(B[312]), .B(n1154), .Z(n1153) );
  NANDN U1354 ( .A(A[312]), .B(n1155), .Z(n1154) );
  NANDN U1355 ( .A(n1155), .B(A[312]), .Z(n1152) );
  XOR U1356 ( .A(n1155), .B(n1156), .Z(DIFF[312]) );
  XOR U1357 ( .A(B[312]), .B(A[312]), .Z(n1156) );
  AND U1358 ( .A(n1157), .B(n1158), .Z(n1155) );
  NANDN U1359 ( .A(B[311]), .B(n1159), .Z(n1158) );
  NANDN U1360 ( .A(A[311]), .B(n1160), .Z(n1159) );
  NANDN U1361 ( .A(n1160), .B(A[311]), .Z(n1157) );
  XOR U1362 ( .A(n1160), .B(n1161), .Z(DIFF[311]) );
  XOR U1363 ( .A(B[311]), .B(A[311]), .Z(n1161) );
  AND U1364 ( .A(n1162), .B(n1163), .Z(n1160) );
  NANDN U1365 ( .A(B[310]), .B(n1164), .Z(n1163) );
  NANDN U1366 ( .A(A[310]), .B(n1165), .Z(n1164) );
  NANDN U1367 ( .A(n1165), .B(A[310]), .Z(n1162) );
  XOR U1368 ( .A(n1165), .B(n1166), .Z(DIFF[310]) );
  XOR U1369 ( .A(B[310]), .B(A[310]), .Z(n1166) );
  AND U1370 ( .A(n1167), .B(n1168), .Z(n1165) );
  NANDN U1371 ( .A(B[309]), .B(n1169), .Z(n1168) );
  NANDN U1372 ( .A(A[309]), .B(n1170), .Z(n1169) );
  NANDN U1373 ( .A(n1170), .B(A[309]), .Z(n1167) );
  XOR U1374 ( .A(n1171), .B(n1172), .Z(DIFF[30]) );
  XOR U1375 ( .A(B[30]), .B(A[30]), .Z(n1172) );
  XOR U1376 ( .A(n1170), .B(n1173), .Z(DIFF[309]) );
  XOR U1377 ( .A(B[309]), .B(A[309]), .Z(n1173) );
  AND U1378 ( .A(n1174), .B(n1175), .Z(n1170) );
  NANDN U1379 ( .A(B[308]), .B(n1176), .Z(n1175) );
  NANDN U1380 ( .A(A[308]), .B(n1177), .Z(n1176) );
  NANDN U1381 ( .A(n1177), .B(A[308]), .Z(n1174) );
  XOR U1382 ( .A(n1177), .B(n1178), .Z(DIFF[308]) );
  XOR U1383 ( .A(B[308]), .B(A[308]), .Z(n1178) );
  AND U1384 ( .A(n1179), .B(n1180), .Z(n1177) );
  NANDN U1385 ( .A(B[307]), .B(n1181), .Z(n1180) );
  NANDN U1386 ( .A(A[307]), .B(n1182), .Z(n1181) );
  NANDN U1387 ( .A(n1182), .B(A[307]), .Z(n1179) );
  XOR U1388 ( .A(n1182), .B(n1183), .Z(DIFF[307]) );
  XOR U1389 ( .A(B[307]), .B(A[307]), .Z(n1183) );
  AND U1390 ( .A(n1184), .B(n1185), .Z(n1182) );
  NANDN U1391 ( .A(B[306]), .B(n1186), .Z(n1185) );
  NANDN U1392 ( .A(A[306]), .B(n1187), .Z(n1186) );
  NANDN U1393 ( .A(n1187), .B(A[306]), .Z(n1184) );
  XOR U1394 ( .A(n1187), .B(n1188), .Z(DIFF[306]) );
  XOR U1395 ( .A(B[306]), .B(A[306]), .Z(n1188) );
  AND U1396 ( .A(n1189), .B(n1190), .Z(n1187) );
  NANDN U1397 ( .A(B[305]), .B(n1191), .Z(n1190) );
  NANDN U1398 ( .A(A[305]), .B(n1192), .Z(n1191) );
  NANDN U1399 ( .A(n1192), .B(A[305]), .Z(n1189) );
  XOR U1400 ( .A(n1192), .B(n1193), .Z(DIFF[305]) );
  XOR U1401 ( .A(B[305]), .B(A[305]), .Z(n1193) );
  AND U1402 ( .A(n1194), .B(n1195), .Z(n1192) );
  NANDN U1403 ( .A(B[304]), .B(n1196), .Z(n1195) );
  NANDN U1404 ( .A(A[304]), .B(n1197), .Z(n1196) );
  NANDN U1405 ( .A(n1197), .B(A[304]), .Z(n1194) );
  XOR U1406 ( .A(n1197), .B(n1198), .Z(DIFF[304]) );
  XOR U1407 ( .A(B[304]), .B(A[304]), .Z(n1198) );
  AND U1408 ( .A(n1199), .B(n1200), .Z(n1197) );
  NANDN U1409 ( .A(B[303]), .B(n1201), .Z(n1200) );
  NANDN U1410 ( .A(A[303]), .B(n1202), .Z(n1201) );
  NANDN U1411 ( .A(n1202), .B(A[303]), .Z(n1199) );
  XOR U1412 ( .A(n1202), .B(n1203), .Z(DIFF[303]) );
  XOR U1413 ( .A(B[303]), .B(A[303]), .Z(n1203) );
  AND U1414 ( .A(n1204), .B(n1205), .Z(n1202) );
  NANDN U1415 ( .A(B[302]), .B(n1206), .Z(n1205) );
  NANDN U1416 ( .A(A[302]), .B(n1207), .Z(n1206) );
  NANDN U1417 ( .A(n1207), .B(A[302]), .Z(n1204) );
  XOR U1418 ( .A(n1207), .B(n1208), .Z(DIFF[302]) );
  XOR U1419 ( .A(B[302]), .B(A[302]), .Z(n1208) );
  AND U1420 ( .A(n1209), .B(n1210), .Z(n1207) );
  NANDN U1421 ( .A(B[301]), .B(n1211), .Z(n1210) );
  NANDN U1422 ( .A(A[301]), .B(n1212), .Z(n1211) );
  NANDN U1423 ( .A(n1212), .B(A[301]), .Z(n1209) );
  XOR U1424 ( .A(n1212), .B(n1213), .Z(DIFF[301]) );
  XOR U1425 ( .A(B[301]), .B(A[301]), .Z(n1213) );
  AND U1426 ( .A(n1214), .B(n1215), .Z(n1212) );
  NANDN U1427 ( .A(B[300]), .B(n1216), .Z(n1215) );
  NANDN U1428 ( .A(A[300]), .B(n1217), .Z(n1216) );
  NANDN U1429 ( .A(n1217), .B(A[300]), .Z(n1214) );
  XOR U1430 ( .A(n1217), .B(n1218), .Z(DIFF[300]) );
  XOR U1431 ( .A(B[300]), .B(A[300]), .Z(n1218) );
  AND U1432 ( .A(n1219), .B(n1220), .Z(n1217) );
  NANDN U1433 ( .A(B[299]), .B(n1221), .Z(n1220) );
  NANDN U1434 ( .A(A[299]), .B(n1222), .Z(n1221) );
  NANDN U1435 ( .A(n1222), .B(A[299]), .Z(n1219) );
  XOR U1436 ( .A(n1223), .B(n1224), .Z(DIFF[2]) );
  XOR U1437 ( .A(B[2]), .B(A[2]), .Z(n1224) );
  XOR U1438 ( .A(n1225), .B(n1226), .Z(DIFF[29]) );
  XOR U1439 ( .A(B[29]), .B(A[29]), .Z(n1226) );
  XOR U1440 ( .A(n1222), .B(n1227), .Z(DIFF[299]) );
  XOR U1441 ( .A(B[299]), .B(A[299]), .Z(n1227) );
  AND U1442 ( .A(n1228), .B(n1229), .Z(n1222) );
  NANDN U1443 ( .A(B[298]), .B(n1230), .Z(n1229) );
  NANDN U1444 ( .A(A[298]), .B(n1231), .Z(n1230) );
  NANDN U1445 ( .A(n1231), .B(A[298]), .Z(n1228) );
  XOR U1446 ( .A(n1231), .B(n1232), .Z(DIFF[298]) );
  XOR U1447 ( .A(B[298]), .B(A[298]), .Z(n1232) );
  AND U1448 ( .A(n1233), .B(n1234), .Z(n1231) );
  NANDN U1449 ( .A(B[297]), .B(n1235), .Z(n1234) );
  NANDN U1450 ( .A(A[297]), .B(n1236), .Z(n1235) );
  NANDN U1451 ( .A(n1236), .B(A[297]), .Z(n1233) );
  XOR U1452 ( .A(n1236), .B(n1237), .Z(DIFF[297]) );
  XOR U1453 ( .A(B[297]), .B(A[297]), .Z(n1237) );
  AND U1454 ( .A(n1238), .B(n1239), .Z(n1236) );
  NANDN U1455 ( .A(B[296]), .B(n1240), .Z(n1239) );
  NANDN U1456 ( .A(A[296]), .B(n1241), .Z(n1240) );
  NANDN U1457 ( .A(n1241), .B(A[296]), .Z(n1238) );
  XOR U1458 ( .A(n1241), .B(n1242), .Z(DIFF[296]) );
  XOR U1459 ( .A(B[296]), .B(A[296]), .Z(n1242) );
  AND U1460 ( .A(n1243), .B(n1244), .Z(n1241) );
  NANDN U1461 ( .A(B[295]), .B(n1245), .Z(n1244) );
  NANDN U1462 ( .A(A[295]), .B(n1246), .Z(n1245) );
  NANDN U1463 ( .A(n1246), .B(A[295]), .Z(n1243) );
  XOR U1464 ( .A(n1246), .B(n1247), .Z(DIFF[295]) );
  XOR U1465 ( .A(B[295]), .B(A[295]), .Z(n1247) );
  AND U1466 ( .A(n1248), .B(n1249), .Z(n1246) );
  NANDN U1467 ( .A(B[294]), .B(n1250), .Z(n1249) );
  NANDN U1468 ( .A(A[294]), .B(n1251), .Z(n1250) );
  NANDN U1469 ( .A(n1251), .B(A[294]), .Z(n1248) );
  XOR U1470 ( .A(n1251), .B(n1252), .Z(DIFF[294]) );
  XOR U1471 ( .A(B[294]), .B(A[294]), .Z(n1252) );
  AND U1472 ( .A(n1253), .B(n1254), .Z(n1251) );
  NANDN U1473 ( .A(B[293]), .B(n1255), .Z(n1254) );
  NANDN U1474 ( .A(A[293]), .B(n1256), .Z(n1255) );
  NANDN U1475 ( .A(n1256), .B(A[293]), .Z(n1253) );
  XOR U1476 ( .A(n1256), .B(n1257), .Z(DIFF[293]) );
  XOR U1477 ( .A(B[293]), .B(A[293]), .Z(n1257) );
  AND U1478 ( .A(n1258), .B(n1259), .Z(n1256) );
  NANDN U1479 ( .A(B[292]), .B(n1260), .Z(n1259) );
  NANDN U1480 ( .A(A[292]), .B(n1261), .Z(n1260) );
  NANDN U1481 ( .A(n1261), .B(A[292]), .Z(n1258) );
  XOR U1482 ( .A(n1261), .B(n1262), .Z(DIFF[292]) );
  XOR U1483 ( .A(B[292]), .B(A[292]), .Z(n1262) );
  AND U1484 ( .A(n1263), .B(n1264), .Z(n1261) );
  NANDN U1485 ( .A(B[291]), .B(n1265), .Z(n1264) );
  NANDN U1486 ( .A(A[291]), .B(n1266), .Z(n1265) );
  NANDN U1487 ( .A(n1266), .B(A[291]), .Z(n1263) );
  XOR U1488 ( .A(n1266), .B(n1267), .Z(DIFF[291]) );
  XOR U1489 ( .A(B[291]), .B(A[291]), .Z(n1267) );
  AND U1490 ( .A(n1268), .B(n1269), .Z(n1266) );
  NANDN U1491 ( .A(B[290]), .B(n1270), .Z(n1269) );
  NANDN U1492 ( .A(A[290]), .B(n1271), .Z(n1270) );
  NANDN U1493 ( .A(n1271), .B(A[290]), .Z(n1268) );
  XOR U1494 ( .A(n1271), .B(n1272), .Z(DIFF[290]) );
  XOR U1495 ( .A(B[290]), .B(A[290]), .Z(n1272) );
  AND U1496 ( .A(n1273), .B(n1274), .Z(n1271) );
  NANDN U1497 ( .A(B[289]), .B(n1275), .Z(n1274) );
  NANDN U1498 ( .A(A[289]), .B(n1276), .Z(n1275) );
  NANDN U1499 ( .A(n1276), .B(A[289]), .Z(n1273) );
  XOR U1500 ( .A(n1277), .B(n1278), .Z(DIFF[28]) );
  XOR U1501 ( .A(B[28]), .B(A[28]), .Z(n1278) );
  XOR U1502 ( .A(n1276), .B(n1279), .Z(DIFF[289]) );
  XOR U1503 ( .A(B[289]), .B(A[289]), .Z(n1279) );
  AND U1504 ( .A(n1280), .B(n1281), .Z(n1276) );
  NANDN U1505 ( .A(B[288]), .B(n1282), .Z(n1281) );
  NANDN U1506 ( .A(A[288]), .B(n1283), .Z(n1282) );
  NANDN U1507 ( .A(n1283), .B(A[288]), .Z(n1280) );
  XOR U1508 ( .A(n1283), .B(n1284), .Z(DIFF[288]) );
  XOR U1509 ( .A(B[288]), .B(A[288]), .Z(n1284) );
  AND U1510 ( .A(n1285), .B(n1286), .Z(n1283) );
  NANDN U1511 ( .A(B[287]), .B(n1287), .Z(n1286) );
  NANDN U1512 ( .A(A[287]), .B(n1288), .Z(n1287) );
  NANDN U1513 ( .A(n1288), .B(A[287]), .Z(n1285) );
  XOR U1514 ( .A(n1288), .B(n1289), .Z(DIFF[287]) );
  XOR U1515 ( .A(B[287]), .B(A[287]), .Z(n1289) );
  AND U1516 ( .A(n1290), .B(n1291), .Z(n1288) );
  NANDN U1517 ( .A(B[286]), .B(n1292), .Z(n1291) );
  NANDN U1518 ( .A(A[286]), .B(n1293), .Z(n1292) );
  NANDN U1519 ( .A(n1293), .B(A[286]), .Z(n1290) );
  XOR U1520 ( .A(n1293), .B(n1294), .Z(DIFF[286]) );
  XOR U1521 ( .A(B[286]), .B(A[286]), .Z(n1294) );
  AND U1522 ( .A(n1295), .B(n1296), .Z(n1293) );
  NANDN U1523 ( .A(B[285]), .B(n1297), .Z(n1296) );
  NANDN U1524 ( .A(A[285]), .B(n1298), .Z(n1297) );
  NANDN U1525 ( .A(n1298), .B(A[285]), .Z(n1295) );
  XOR U1526 ( .A(n1298), .B(n1299), .Z(DIFF[285]) );
  XOR U1527 ( .A(B[285]), .B(A[285]), .Z(n1299) );
  AND U1528 ( .A(n1300), .B(n1301), .Z(n1298) );
  NANDN U1529 ( .A(B[284]), .B(n1302), .Z(n1301) );
  NANDN U1530 ( .A(A[284]), .B(n1303), .Z(n1302) );
  NANDN U1531 ( .A(n1303), .B(A[284]), .Z(n1300) );
  XOR U1532 ( .A(n1303), .B(n1304), .Z(DIFF[284]) );
  XOR U1533 ( .A(B[284]), .B(A[284]), .Z(n1304) );
  AND U1534 ( .A(n1305), .B(n1306), .Z(n1303) );
  NANDN U1535 ( .A(B[283]), .B(n1307), .Z(n1306) );
  NANDN U1536 ( .A(A[283]), .B(n1308), .Z(n1307) );
  NANDN U1537 ( .A(n1308), .B(A[283]), .Z(n1305) );
  XOR U1538 ( .A(n1308), .B(n1309), .Z(DIFF[283]) );
  XOR U1539 ( .A(B[283]), .B(A[283]), .Z(n1309) );
  AND U1540 ( .A(n1310), .B(n1311), .Z(n1308) );
  NANDN U1541 ( .A(B[282]), .B(n1312), .Z(n1311) );
  NANDN U1542 ( .A(A[282]), .B(n1313), .Z(n1312) );
  NANDN U1543 ( .A(n1313), .B(A[282]), .Z(n1310) );
  XOR U1544 ( .A(n1313), .B(n1314), .Z(DIFF[282]) );
  XOR U1545 ( .A(B[282]), .B(A[282]), .Z(n1314) );
  AND U1546 ( .A(n1315), .B(n1316), .Z(n1313) );
  NANDN U1547 ( .A(B[281]), .B(n1317), .Z(n1316) );
  NANDN U1548 ( .A(A[281]), .B(n1318), .Z(n1317) );
  NANDN U1549 ( .A(n1318), .B(A[281]), .Z(n1315) );
  XOR U1550 ( .A(n1318), .B(n1319), .Z(DIFF[281]) );
  XOR U1551 ( .A(B[281]), .B(A[281]), .Z(n1319) );
  AND U1552 ( .A(n1320), .B(n1321), .Z(n1318) );
  NANDN U1553 ( .A(B[280]), .B(n1322), .Z(n1321) );
  NANDN U1554 ( .A(A[280]), .B(n1323), .Z(n1322) );
  NANDN U1555 ( .A(n1323), .B(A[280]), .Z(n1320) );
  XOR U1556 ( .A(n1323), .B(n1324), .Z(DIFF[280]) );
  XOR U1557 ( .A(B[280]), .B(A[280]), .Z(n1324) );
  AND U1558 ( .A(n1325), .B(n1326), .Z(n1323) );
  NANDN U1559 ( .A(B[279]), .B(n1327), .Z(n1326) );
  NANDN U1560 ( .A(A[279]), .B(n1328), .Z(n1327) );
  NANDN U1561 ( .A(n1328), .B(A[279]), .Z(n1325) );
  XOR U1562 ( .A(n1329), .B(n1330), .Z(DIFF[27]) );
  XOR U1563 ( .A(B[27]), .B(A[27]), .Z(n1330) );
  XOR U1564 ( .A(n1328), .B(n1331), .Z(DIFF[279]) );
  XOR U1565 ( .A(B[279]), .B(A[279]), .Z(n1331) );
  AND U1566 ( .A(n1332), .B(n1333), .Z(n1328) );
  NANDN U1567 ( .A(B[278]), .B(n1334), .Z(n1333) );
  NANDN U1568 ( .A(A[278]), .B(n1335), .Z(n1334) );
  NANDN U1569 ( .A(n1335), .B(A[278]), .Z(n1332) );
  XOR U1570 ( .A(n1335), .B(n1336), .Z(DIFF[278]) );
  XOR U1571 ( .A(B[278]), .B(A[278]), .Z(n1336) );
  AND U1572 ( .A(n1337), .B(n1338), .Z(n1335) );
  NANDN U1573 ( .A(B[277]), .B(n1339), .Z(n1338) );
  NANDN U1574 ( .A(A[277]), .B(n1340), .Z(n1339) );
  NANDN U1575 ( .A(n1340), .B(A[277]), .Z(n1337) );
  XOR U1576 ( .A(n1340), .B(n1341), .Z(DIFF[277]) );
  XOR U1577 ( .A(B[277]), .B(A[277]), .Z(n1341) );
  AND U1578 ( .A(n1342), .B(n1343), .Z(n1340) );
  NANDN U1579 ( .A(B[276]), .B(n1344), .Z(n1343) );
  NANDN U1580 ( .A(A[276]), .B(n1345), .Z(n1344) );
  NANDN U1581 ( .A(n1345), .B(A[276]), .Z(n1342) );
  XOR U1582 ( .A(n1345), .B(n1346), .Z(DIFF[276]) );
  XOR U1583 ( .A(B[276]), .B(A[276]), .Z(n1346) );
  AND U1584 ( .A(n1347), .B(n1348), .Z(n1345) );
  NANDN U1585 ( .A(B[275]), .B(n1349), .Z(n1348) );
  NANDN U1586 ( .A(A[275]), .B(n1350), .Z(n1349) );
  NANDN U1587 ( .A(n1350), .B(A[275]), .Z(n1347) );
  XOR U1588 ( .A(n1350), .B(n1351), .Z(DIFF[275]) );
  XOR U1589 ( .A(B[275]), .B(A[275]), .Z(n1351) );
  AND U1590 ( .A(n1352), .B(n1353), .Z(n1350) );
  NANDN U1591 ( .A(B[274]), .B(n1354), .Z(n1353) );
  NANDN U1592 ( .A(A[274]), .B(n1355), .Z(n1354) );
  NANDN U1593 ( .A(n1355), .B(A[274]), .Z(n1352) );
  XOR U1594 ( .A(n1355), .B(n1356), .Z(DIFF[274]) );
  XOR U1595 ( .A(B[274]), .B(A[274]), .Z(n1356) );
  AND U1596 ( .A(n1357), .B(n1358), .Z(n1355) );
  NANDN U1597 ( .A(B[273]), .B(n1359), .Z(n1358) );
  NANDN U1598 ( .A(A[273]), .B(n1360), .Z(n1359) );
  NANDN U1599 ( .A(n1360), .B(A[273]), .Z(n1357) );
  XOR U1600 ( .A(n1360), .B(n1361), .Z(DIFF[273]) );
  XOR U1601 ( .A(B[273]), .B(A[273]), .Z(n1361) );
  AND U1602 ( .A(n1362), .B(n1363), .Z(n1360) );
  NANDN U1603 ( .A(B[272]), .B(n1364), .Z(n1363) );
  NANDN U1604 ( .A(A[272]), .B(n1365), .Z(n1364) );
  NANDN U1605 ( .A(n1365), .B(A[272]), .Z(n1362) );
  XOR U1606 ( .A(n1365), .B(n1366), .Z(DIFF[272]) );
  XOR U1607 ( .A(B[272]), .B(A[272]), .Z(n1366) );
  AND U1608 ( .A(n1367), .B(n1368), .Z(n1365) );
  NANDN U1609 ( .A(B[271]), .B(n1369), .Z(n1368) );
  NANDN U1610 ( .A(A[271]), .B(n1370), .Z(n1369) );
  NANDN U1611 ( .A(n1370), .B(A[271]), .Z(n1367) );
  XOR U1612 ( .A(n1370), .B(n1371), .Z(DIFF[271]) );
  XOR U1613 ( .A(B[271]), .B(A[271]), .Z(n1371) );
  AND U1614 ( .A(n1372), .B(n1373), .Z(n1370) );
  NANDN U1615 ( .A(B[270]), .B(n1374), .Z(n1373) );
  NANDN U1616 ( .A(A[270]), .B(n1375), .Z(n1374) );
  NANDN U1617 ( .A(n1375), .B(A[270]), .Z(n1372) );
  XOR U1618 ( .A(n1375), .B(n1376), .Z(DIFF[270]) );
  XOR U1619 ( .A(B[270]), .B(A[270]), .Z(n1376) );
  AND U1620 ( .A(n1377), .B(n1378), .Z(n1375) );
  NANDN U1621 ( .A(B[269]), .B(n1379), .Z(n1378) );
  NANDN U1622 ( .A(A[269]), .B(n1380), .Z(n1379) );
  NANDN U1623 ( .A(n1380), .B(A[269]), .Z(n1377) );
  XOR U1624 ( .A(n1381), .B(n1382), .Z(DIFF[26]) );
  XOR U1625 ( .A(B[26]), .B(A[26]), .Z(n1382) );
  XOR U1626 ( .A(n1380), .B(n1383), .Z(DIFF[269]) );
  XOR U1627 ( .A(B[269]), .B(A[269]), .Z(n1383) );
  AND U1628 ( .A(n1384), .B(n1385), .Z(n1380) );
  NANDN U1629 ( .A(B[268]), .B(n1386), .Z(n1385) );
  NANDN U1630 ( .A(A[268]), .B(n1387), .Z(n1386) );
  NANDN U1631 ( .A(n1387), .B(A[268]), .Z(n1384) );
  XOR U1632 ( .A(n1387), .B(n1388), .Z(DIFF[268]) );
  XOR U1633 ( .A(B[268]), .B(A[268]), .Z(n1388) );
  AND U1634 ( .A(n1389), .B(n1390), .Z(n1387) );
  NANDN U1635 ( .A(B[267]), .B(n1391), .Z(n1390) );
  NANDN U1636 ( .A(A[267]), .B(n1392), .Z(n1391) );
  NANDN U1637 ( .A(n1392), .B(A[267]), .Z(n1389) );
  XOR U1638 ( .A(n1392), .B(n1393), .Z(DIFF[267]) );
  XOR U1639 ( .A(B[267]), .B(A[267]), .Z(n1393) );
  AND U1640 ( .A(n1394), .B(n1395), .Z(n1392) );
  NANDN U1641 ( .A(B[266]), .B(n1396), .Z(n1395) );
  NANDN U1642 ( .A(A[266]), .B(n1397), .Z(n1396) );
  NANDN U1643 ( .A(n1397), .B(A[266]), .Z(n1394) );
  XOR U1644 ( .A(n1397), .B(n1398), .Z(DIFF[266]) );
  XOR U1645 ( .A(B[266]), .B(A[266]), .Z(n1398) );
  AND U1646 ( .A(n1399), .B(n1400), .Z(n1397) );
  NANDN U1647 ( .A(B[265]), .B(n1401), .Z(n1400) );
  NANDN U1648 ( .A(A[265]), .B(n1402), .Z(n1401) );
  NANDN U1649 ( .A(n1402), .B(A[265]), .Z(n1399) );
  XOR U1650 ( .A(n1402), .B(n1403), .Z(DIFF[265]) );
  XOR U1651 ( .A(B[265]), .B(A[265]), .Z(n1403) );
  AND U1652 ( .A(n1404), .B(n1405), .Z(n1402) );
  NANDN U1653 ( .A(B[264]), .B(n1406), .Z(n1405) );
  NANDN U1654 ( .A(A[264]), .B(n1407), .Z(n1406) );
  NANDN U1655 ( .A(n1407), .B(A[264]), .Z(n1404) );
  XOR U1656 ( .A(n1407), .B(n1408), .Z(DIFF[264]) );
  XOR U1657 ( .A(B[264]), .B(A[264]), .Z(n1408) );
  AND U1658 ( .A(n1409), .B(n1410), .Z(n1407) );
  NANDN U1659 ( .A(B[263]), .B(n1411), .Z(n1410) );
  NANDN U1660 ( .A(A[263]), .B(n1412), .Z(n1411) );
  NANDN U1661 ( .A(n1412), .B(A[263]), .Z(n1409) );
  XOR U1662 ( .A(n1412), .B(n1413), .Z(DIFF[263]) );
  XOR U1663 ( .A(B[263]), .B(A[263]), .Z(n1413) );
  AND U1664 ( .A(n1414), .B(n1415), .Z(n1412) );
  NANDN U1665 ( .A(B[262]), .B(n1416), .Z(n1415) );
  NANDN U1666 ( .A(A[262]), .B(n1417), .Z(n1416) );
  NANDN U1667 ( .A(n1417), .B(A[262]), .Z(n1414) );
  XOR U1668 ( .A(n1417), .B(n1418), .Z(DIFF[262]) );
  XOR U1669 ( .A(B[262]), .B(A[262]), .Z(n1418) );
  AND U1670 ( .A(n1419), .B(n1420), .Z(n1417) );
  NANDN U1671 ( .A(B[261]), .B(n1421), .Z(n1420) );
  NANDN U1672 ( .A(A[261]), .B(n1422), .Z(n1421) );
  NANDN U1673 ( .A(n1422), .B(A[261]), .Z(n1419) );
  XOR U1674 ( .A(n1422), .B(n1423), .Z(DIFF[261]) );
  XOR U1675 ( .A(B[261]), .B(A[261]), .Z(n1423) );
  AND U1676 ( .A(n1424), .B(n1425), .Z(n1422) );
  NANDN U1677 ( .A(B[260]), .B(n1426), .Z(n1425) );
  NANDN U1678 ( .A(A[260]), .B(n1427), .Z(n1426) );
  NANDN U1679 ( .A(n1427), .B(A[260]), .Z(n1424) );
  XOR U1680 ( .A(n1427), .B(n1428), .Z(DIFF[260]) );
  XOR U1681 ( .A(B[260]), .B(A[260]), .Z(n1428) );
  AND U1682 ( .A(n1429), .B(n1430), .Z(n1427) );
  NANDN U1683 ( .A(B[259]), .B(n1431), .Z(n1430) );
  NANDN U1684 ( .A(A[259]), .B(n1432), .Z(n1431) );
  NANDN U1685 ( .A(n1432), .B(A[259]), .Z(n1429) );
  XOR U1686 ( .A(n1433), .B(n1434), .Z(DIFF[25]) );
  XOR U1687 ( .A(B[25]), .B(A[25]), .Z(n1434) );
  XOR U1688 ( .A(n1432), .B(n1435), .Z(DIFF[259]) );
  XOR U1689 ( .A(B[259]), .B(A[259]), .Z(n1435) );
  AND U1690 ( .A(n1436), .B(n1437), .Z(n1432) );
  NANDN U1691 ( .A(B[258]), .B(n1438), .Z(n1437) );
  NANDN U1692 ( .A(A[258]), .B(n1439), .Z(n1438) );
  NANDN U1693 ( .A(n1439), .B(A[258]), .Z(n1436) );
  XOR U1694 ( .A(n1439), .B(n1440), .Z(DIFF[258]) );
  XOR U1695 ( .A(B[258]), .B(A[258]), .Z(n1440) );
  AND U1696 ( .A(n1441), .B(n1442), .Z(n1439) );
  NANDN U1697 ( .A(B[257]), .B(n1443), .Z(n1442) );
  NANDN U1698 ( .A(A[257]), .B(n1444), .Z(n1443) );
  NANDN U1699 ( .A(n1444), .B(A[257]), .Z(n1441) );
  XOR U1700 ( .A(n1444), .B(n1445), .Z(DIFF[257]) );
  XOR U1701 ( .A(B[257]), .B(A[257]), .Z(n1445) );
  AND U1702 ( .A(n1446), .B(n1447), .Z(n1444) );
  NANDN U1703 ( .A(B[256]), .B(n1448), .Z(n1447) );
  NANDN U1704 ( .A(A[256]), .B(n1449), .Z(n1448) );
  NANDN U1705 ( .A(n1449), .B(A[256]), .Z(n1446) );
  XOR U1706 ( .A(n1449), .B(n1450), .Z(DIFF[256]) );
  XOR U1707 ( .A(B[256]), .B(A[256]), .Z(n1450) );
  AND U1708 ( .A(n1451), .B(n1452), .Z(n1449) );
  NANDN U1709 ( .A(B[255]), .B(n1453), .Z(n1452) );
  NANDN U1710 ( .A(A[255]), .B(n1454), .Z(n1453) );
  NANDN U1711 ( .A(n1454), .B(A[255]), .Z(n1451) );
  XOR U1712 ( .A(n1454), .B(n1455), .Z(DIFF[255]) );
  XOR U1713 ( .A(B[255]), .B(A[255]), .Z(n1455) );
  AND U1714 ( .A(n1456), .B(n1457), .Z(n1454) );
  NANDN U1715 ( .A(B[254]), .B(n1458), .Z(n1457) );
  NANDN U1716 ( .A(A[254]), .B(n1459), .Z(n1458) );
  NANDN U1717 ( .A(n1459), .B(A[254]), .Z(n1456) );
  XOR U1718 ( .A(n1459), .B(n1460), .Z(DIFF[254]) );
  XOR U1719 ( .A(B[254]), .B(A[254]), .Z(n1460) );
  AND U1720 ( .A(n1461), .B(n1462), .Z(n1459) );
  NANDN U1721 ( .A(B[253]), .B(n1463), .Z(n1462) );
  NANDN U1722 ( .A(A[253]), .B(n1464), .Z(n1463) );
  NANDN U1723 ( .A(n1464), .B(A[253]), .Z(n1461) );
  XOR U1724 ( .A(n1464), .B(n1465), .Z(DIFF[253]) );
  XOR U1725 ( .A(B[253]), .B(A[253]), .Z(n1465) );
  AND U1726 ( .A(n1466), .B(n1467), .Z(n1464) );
  NANDN U1727 ( .A(B[252]), .B(n1468), .Z(n1467) );
  NANDN U1728 ( .A(A[252]), .B(n1469), .Z(n1468) );
  NANDN U1729 ( .A(n1469), .B(A[252]), .Z(n1466) );
  XOR U1730 ( .A(n1469), .B(n1470), .Z(DIFF[252]) );
  XOR U1731 ( .A(B[252]), .B(A[252]), .Z(n1470) );
  AND U1732 ( .A(n1471), .B(n1472), .Z(n1469) );
  NANDN U1733 ( .A(B[251]), .B(n1473), .Z(n1472) );
  NANDN U1734 ( .A(A[251]), .B(n1474), .Z(n1473) );
  NANDN U1735 ( .A(n1474), .B(A[251]), .Z(n1471) );
  XOR U1736 ( .A(n1474), .B(n1475), .Z(DIFF[251]) );
  XOR U1737 ( .A(B[251]), .B(A[251]), .Z(n1475) );
  AND U1738 ( .A(n1476), .B(n1477), .Z(n1474) );
  NANDN U1739 ( .A(B[250]), .B(n1478), .Z(n1477) );
  NANDN U1740 ( .A(A[250]), .B(n1479), .Z(n1478) );
  NANDN U1741 ( .A(n1479), .B(A[250]), .Z(n1476) );
  XOR U1742 ( .A(n1479), .B(n1480), .Z(DIFF[250]) );
  XOR U1743 ( .A(B[250]), .B(A[250]), .Z(n1480) );
  AND U1744 ( .A(n1481), .B(n1482), .Z(n1479) );
  NANDN U1745 ( .A(B[249]), .B(n1483), .Z(n1482) );
  NANDN U1746 ( .A(A[249]), .B(n1484), .Z(n1483) );
  NANDN U1747 ( .A(n1484), .B(A[249]), .Z(n1481) );
  XOR U1748 ( .A(n1485), .B(n1486), .Z(DIFF[24]) );
  XOR U1749 ( .A(B[24]), .B(A[24]), .Z(n1486) );
  XOR U1750 ( .A(n1484), .B(n1487), .Z(DIFF[249]) );
  XOR U1751 ( .A(B[249]), .B(A[249]), .Z(n1487) );
  AND U1752 ( .A(n1488), .B(n1489), .Z(n1484) );
  NANDN U1753 ( .A(B[248]), .B(n1490), .Z(n1489) );
  NANDN U1754 ( .A(A[248]), .B(n1491), .Z(n1490) );
  NANDN U1755 ( .A(n1491), .B(A[248]), .Z(n1488) );
  XOR U1756 ( .A(n1491), .B(n1492), .Z(DIFF[248]) );
  XOR U1757 ( .A(B[248]), .B(A[248]), .Z(n1492) );
  AND U1758 ( .A(n1493), .B(n1494), .Z(n1491) );
  NANDN U1759 ( .A(B[247]), .B(n1495), .Z(n1494) );
  NANDN U1760 ( .A(A[247]), .B(n1496), .Z(n1495) );
  NANDN U1761 ( .A(n1496), .B(A[247]), .Z(n1493) );
  XOR U1762 ( .A(n1496), .B(n1497), .Z(DIFF[247]) );
  XOR U1763 ( .A(B[247]), .B(A[247]), .Z(n1497) );
  AND U1764 ( .A(n1498), .B(n1499), .Z(n1496) );
  NANDN U1765 ( .A(B[246]), .B(n1500), .Z(n1499) );
  NANDN U1766 ( .A(A[246]), .B(n1501), .Z(n1500) );
  NANDN U1767 ( .A(n1501), .B(A[246]), .Z(n1498) );
  XOR U1768 ( .A(n1501), .B(n1502), .Z(DIFF[246]) );
  XOR U1769 ( .A(B[246]), .B(A[246]), .Z(n1502) );
  AND U1770 ( .A(n1503), .B(n1504), .Z(n1501) );
  NANDN U1771 ( .A(B[245]), .B(n1505), .Z(n1504) );
  NANDN U1772 ( .A(A[245]), .B(n1506), .Z(n1505) );
  NANDN U1773 ( .A(n1506), .B(A[245]), .Z(n1503) );
  XOR U1774 ( .A(n1506), .B(n1507), .Z(DIFF[245]) );
  XOR U1775 ( .A(B[245]), .B(A[245]), .Z(n1507) );
  AND U1776 ( .A(n1508), .B(n1509), .Z(n1506) );
  NANDN U1777 ( .A(B[244]), .B(n1510), .Z(n1509) );
  NANDN U1778 ( .A(A[244]), .B(n1511), .Z(n1510) );
  NANDN U1779 ( .A(n1511), .B(A[244]), .Z(n1508) );
  XOR U1780 ( .A(n1511), .B(n1512), .Z(DIFF[244]) );
  XOR U1781 ( .A(B[244]), .B(A[244]), .Z(n1512) );
  AND U1782 ( .A(n1513), .B(n1514), .Z(n1511) );
  NANDN U1783 ( .A(B[243]), .B(n1515), .Z(n1514) );
  NANDN U1784 ( .A(A[243]), .B(n1516), .Z(n1515) );
  NANDN U1785 ( .A(n1516), .B(A[243]), .Z(n1513) );
  XOR U1786 ( .A(n1516), .B(n1517), .Z(DIFF[243]) );
  XOR U1787 ( .A(B[243]), .B(A[243]), .Z(n1517) );
  AND U1788 ( .A(n1518), .B(n1519), .Z(n1516) );
  NANDN U1789 ( .A(B[242]), .B(n1520), .Z(n1519) );
  NANDN U1790 ( .A(A[242]), .B(n1521), .Z(n1520) );
  NANDN U1791 ( .A(n1521), .B(A[242]), .Z(n1518) );
  XOR U1792 ( .A(n1521), .B(n1522), .Z(DIFF[242]) );
  XOR U1793 ( .A(B[242]), .B(A[242]), .Z(n1522) );
  AND U1794 ( .A(n1523), .B(n1524), .Z(n1521) );
  NANDN U1795 ( .A(B[241]), .B(n1525), .Z(n1524) );
  NANDN U1796 ( .A(A[241]), .B(n1526), .Z(n1525) );
  NANDN U1797 ( .A(n1526), .B(A[241]), .Z(n1523) );
  XOR U1798 ( .A(n1526), .B(n1527), .Z(DIFF[241]) );
  XOR U1799 ( .A(B[241]), .B(A[241]), .Z(n1527) );
  AND U1800 ( .A(n1528), .B(n1529), .Z(n1526) );
  NANDN U1801 ( .A(B[240]), .B(n1530), .Z(n1529) );
  NANDN U1802 ( .A(A[240]), .B(n1531), .Z(n1530) );
  NANDN U1803 ( .A(n1531), .B(A[240]), .Z(n1528) );
  XOR U1804 ( .A(n1531), .B(n1532), .Z(DIFF[240]) );
  XOR U1805 ( .A(B[240]), .B(A[240]), .Z(n1532) );
  AND U1806 ( .A(n1533), .B(n1534), .Z(n1531) );
  NANDN U1807 ( .A(B[239]), .B(n1535), .Z(n1534) );
  NANDN U1808 ( .A(A[239]), .B(n1536), .Z(n1535) );
  NANDN U1809 ( .A(n1536), .B(A[239]), .Z(n1533) );
  XOR U1810 ( .A(n1537), .B(n1538), .Z(DIFF[23]) );
  XOR U1811 ( .A(B[23]), .B(A[23]), .Z(n1538) );
  XOR U1812 ( .A(n1536), .B(n1539), .Z(DIFF[239]) );
  XOR U1813 ( .A(B[239]), .B(A[239]), .Z(n1539) );
  AND U1814 ( .A(n1540), .B(n1541), .Z(n1536) );
  NANDN U1815 ( .A(B[238]), .B(n1542), .Z(n1541) );
  NANDN U1816 ( .A(A[238]), .B(n1543), .Z(n1542) );
  NANDN U1817 ( .A(n1543), .B(A[238]), .Z(n1540) );
  XOR U1818 ( .A(n1543), .B(n1544), .Z(DIFF[238]) );
  XOR U1819 ( .A(B[238]), .B(A[238]), .Z(n1544) );
  AND U1820 ( .A(n1545), .B(n1546), .Z(n1543) );
  NANDN U1821 ( .A(B[237]), .B(n1547), .Z(n1546) );
  NANDN U1822 ( .A(A[237]), .B(n1548), .Z(n1547) );
  NANDN U1823 ( .A(n1548), .B(A[237]), .Z(n1545) );
  XOR U1824 ( .A(n1548), .B(n1549), .Z(DIFF[237]) );
  XOR U1825 ( .A(B[237]), .B(A[237]), .Z(n1549) );
  AND U1826 ( .A(n1550), .B(n1551), .Z(n1548) );
  NANDN U1827 ( .A(B[236]), .B(n1552), .Z(n1551) );
  NANDN U1828 ( .A(A[236]), .B(n1553), .Z(n1552) );
  NANDN U1829 ( .A(n1553), .B(A[236]), .Z(n1550) );
  XOR U1830 ( .A(n1553), .B(n1554), .Z(DIFF[236]) );
  XOR U1831 ( .A(B[236]), .B(A[236]), .Z(n1554) );
  AND U1832 ( .A(n1555), .B(n1556), .Z(n1553) );
  NANDN U1833 ( .A(B[235]), .B(n1557), .Z(n1556) );
  NANDN U1834 ( .A(A[235]), .B(n1558), .Z(n1557) );
  NANDN U1835 ( .A(n1558), .B(A[235]), .Z(n1555) );
  XOR U1836 ( .A(n1558), .B(n1559), .Z(DIFF[235]) );
  XOR U1837 ( .A(B[235]), .B(A[235]), .Z(n1559) );
  AND U1838 ( .A(n1560), .B(n1561), .Z(n1558) );
  NANDN U1839 ( .A(B[234]), .B(n1562), .Z(n1561) );
  NANDN U1840 ( .A(A[234]), .B(n1563), .Z(n1562) );
  NANDN U1841 ( .A(n1563), .B(A[234]), .Z(n1560) );
  XOR U1842 ( .A(n1563), .B(n1564), .Z(DIFF[234]) );
  XOR U1843 ( .A(B[234]), .B(A[234]), .Z(n1564) );
  AND U1844 ( .A(n1565), .B(n1566), .Z(n1563) );
  NANDN U1845 ( .A(B[233]), .B(n1567), .Z(n1566) );
  NANDN U1846 ( .A(A[233]), .B(n1568), .Z(n1567) );
  NANDN U1847 ( .A(n1568), .B(A[233]), .Z(n1565) );
  XOR U1848 ( .A(n1568), .B(n1569), .Z(DIFF[233]) );
  XOR U1849 ( .A(B[233]), .B(A[233]), .Z(n1569) );
  AND U1850 ( .A(n1570), .B(n1571), .Z(n1568) );
  NANDN U1851 ( .A(B[232]), .B(n1572), .Z(n1571) );
  NANDN U1852 ( .A(A[232]), .B(n1573), .Z(n1572) );
  NANDN U1853 ( .A(n1573), .B(A[232]), .Z(n1570) );
  XOR U1854 ( .A(n1573), .B(n1574), .Z(DIFF[232]) );
  XOR U1855 ( .A(B[232]), .B(A[232]), .Z(n1574) );
  AND U1856 ( .A(n1575), .B(n1576), .Z(n1573) );
  NANDN U1857 ( .A(B[231]), .B(n1577), .Z(n1576) );
  NANDN U1858 ( .A(A[231]), .B(n1578), .Z(n1577) );
  NANDN U1859 ( .A(n1578), .B(A[231]), .Z(n1575) );
  XOR U1860 ( .A(n1578), .B(n1579), .Z(DIFF[231]) );
  XOR U1861 ( .A(B[231]), .B(A[231]), .Z(n1579) );
  AND U1862 ( .A(n1580), .B(n1581), .Z(n1578) );
  NANDN U1863 ( .A(B[230]), .B(n1582), .Z(n1581) );
  NANDN U1864 ( .A(A[230]), .B(n1583), .Z(n1582) );
  NANDN U1865 ( .A(n1583), .B(A[230]), .Z(n1580) );
  XOR U1866 ( .A(n1583), .B(n1584), .Z(DIFF[230]) );
  XOR U1867 ( .A(B[230]), .B(A[230]), .Z(n1584) );
  AND U1868 ( .A(n1585), .B(n1586), .Z(n1583) );
  NANDN U1869 ( .A(B[229]), .B(n1587), .Z(n1586) );
  NANDN U1870 ( .A(A[229]), .B(n1588), .Z(n1587) );
  NANDN U1871 ( .A(n1588), .B(A[229]), .Z(n1585) );
  XOR U1872 ( .A(n1589), .B(n1590), .Z(DIFF[22]) );
  XOR U1873 ( .A(B[22]), .B(A[22]), .Z(n1590) );
  XOR U1874 ( .A(n1588), .B(n1591), .Z(DIFF[229]) );
  XOR U1875 ( .A(B[229]), .B(A[229]), .Z(n1591) );
  AND U1876 ( .A(n1592), .B(n1593), .Z(n1588) );
  NANDN U1877 ( .A(B[228]), .B(n1594), .Z(n1593) );
  NANDN U1878 ( .A(A[228]), .B(n1595), .Z(n1594) );
  NANDN U1879 ( .A(n1595), .B(A[228]), .Z(n1592) );
  XOR U1880 ( .A(n1595), .B(n1596), .Z(DIFF[228]) );
  XOR U1881 ( .A(B[228]), .B(A[228]), .Z(n1596) );
  AND U1882 ( .A(n1597), .B(n1598), .Z(n1595) );
  NANDN U1883 ( .A(B[227]), .B(n1599), .Z(n1598) );
  NANDN U1884 ( .A(A[227]), .B(n1600), .Z(n1599) );
  NANDN U1885 ( .A(n1600), .B(A[227]), .Z(n1597) );
  XOR U1886 ( .A(n1600), .B(n1601), .Z(DIFF[227]) );
  XOR U1887 ( .A(B[227]), .B(A[227]), .Z(n1601) );
  AND U1888 ( .A(n1602), .B(n1603), .Z(n1600) );
  NANDN U1889 ( .A(B[226]), .B(n1604), .Z(n1603) );
  NANDN U1890 ( .A(A[226]), .B(n1605), .Z(n1604) );
  NANDN U1891 ( .A(n1605), .B(A[226]), .Z(n1602) );
  XOR U1892 ( .A(n1605), .B(n1606), .Z(DIFF[226]) );
  XOR U1893 ( .A(B[226]), .B(A[226]), .Z(n1606) );
  AND U1894 ( .A(n1607), .B(n1608), .Z(n1605) );
  NANDN U1895 ( .A(B[225]), .B(n1609), .Z(n1608) );
  NANDN U1896 ( .A(A[225]), .B(n1610), .Z(n1609) );
  NANDN U1897 ( .A(n1610), .B(A[225]), .Z(n1607) );
  XOR U1898 ( .A(n1610), .B(n1611), .Z(DIFF[225]) );
  XOR U1899 ( .A(B[225]), .B(A[225]), .Z(n1611) );
  AND U1900 ( .A(n1612), .B(n1613), .Z(n1610) );
  NANDN U1901 ( .A(B[224]), .B(n1614), .Z(n1613) );
  NANDN U1902 ( .A(A[224]), .B(n1615), .Z(n1614) );
  NANDN U1903 ( .A(n1615), .B(A[224]), .Z(n1612) );
  XOR U1904 ( .A(n1615), .B(n1616), .Z(DIFF[224]) );
  XOR U1905 ( .A(B[224]), .B(A[224]), .Z(n1616) );
  AND U1906 ( .A(n1617), .B(n1618), .Z(n1615) );
  NANDN U1907 ( .A(B[223]), .B(n1619), .Z(n1618) );
  NANDN U1908 ( .A(A[223]), .B(n1620), .Z(n1619) );
  NANDN U1909 ( .A(n1620), .B(A[223]), .Z(n1617) );
  XOR U1910 ( .A(n1620), .B(n1621), .Z(DIFF[223]) );
  XOR U1911 ( .A(B[223]), .B(A[223]), .Z(n1621) );
  AND U1912 ( .A(n1622), .B(n1623), .Z(n1620) );
  NANDN U1913 ( .A(B[222]), .B(n1624), .Z(n1623) );
  NANDN U1914 ( .A(A[222]), .B(n1625), .Z(n1624) );
  NANDN U1915 ( .A(n1625), .B(A[222]), .Z(n1622) );
  XOR U1916 ( .A(n1625), .B(n1626), .Z(DIFF[222]) );
  XOR U1917 ( .A(B[222]), .B(A[222]), .Z(n1626) );
  AND U1918 ( .A(n1627), .B(n1628), .Z(n1625) );
  NANDN U1919 ( .A(B[221]), .B(n1629), .Z(n1628) );
  NANDN U1920 ( .A(A[221]), .B(n1630), .Z(n1629) );
  NANDN U1921 ( .A(n1630), .B(A[221]), .Z(n1627) );
  XOR U1922 ( .A(n1630), .B(n1631), .Z(DIFF[221]) );
  XOR U1923 ( .A(B[221]), .B(A[221]), .Z(n1631) );
  AND U1924 ( .A(n1632), .B(n1633), .Z(n1630) );
  NANDN U1925 ( .A(B[220]), .B(n1634), .Z(n1633) );
  NANDN U1926 ( .A(A[220]), .B(n1635), .Z(n1634) );
  NANDN U1927 ( .A(n1635), .B(A[220]), .Z(n1632) );
  XOR U1928 ( .A(n1635), .B(n1636), .Z(DIFF[220]) );
  XOR U1929 ( .A(B[220]), .B(A[220]), .Z(n1636) );
  AND U1930 ( .A(n1637), .B(n1638), .Z(n1635) );
  NANDN U1931 ( .A(B[219]), .B(n1639), .Z(n1638) );
  NANDN U1932 ( .A(A[219]), .B(n1640), .Z(n1639) );
  NANDN U1933 ( .A(n1640), .B(A[219]), .Z(n1637) );
  XOR U1934 ( .A(n1641), .B(n1642), .Z(DIFF[21]) );
  XOR U1935 ( .A(B[21]), .B(A[21]), .Z(n1642) );
  XOR U1936 ( .A(n1640), .B(n1643), .Z(DIFF[219]) );
  XOR U1937 ( .A(B[219]), .B(A[219]), .Z(n1643) );
  AND U1938 ( .A(n1644), .B(n1645), .Z(n1640) );
  NANDN U1939 ( .A(B[218]), .B(n1646), .Z(n1645) );
  NANDN U1940 ( .A(A[218]), .B(n1647), .Z(n1646) );
  NANDN U1941 ( .A(n1647), .B(A[218]), .Z(n1644) );
  XOR U1942 ( .A(n1647), .B(n1648), .Z(DIFF[218]) );
  XOR U1943 ( .A(B[218]), .B(A[218]), .Z(n1648) );
  AND U1944 ( .A(n1649), .B(n1650), .Z(n1647) );
  NANDN U1945 ( .A(B[217]), .B(n1651), .Z(n1650) );
  NANDN U1946 ( .A(A[217]), .B(n1652), .Z(n1651) );
  NANDN U1947 ( .A(n1652), .B(A[217]), .Z(n1649) );
  XOR U1948 ( .A(n1652), .B(n1653), .Z(DIFF[217]) );
  XOR U1949 ( .A(B[217]), .B(A[217]), .Z(n1653) );
  AND U1950 ( .A(n1654), .B(n1655), .Z(n1652) );
  NANDN U1951 ( .A(B[216]), .B(n1656), .Z(n1655) );
  NANDN U1952 ( .A(A[216]), .B(n1657), .Z(n1656) );
  NANDN U1953 ( .A(n1657), .B(A[216]), .Z(n1654) );
  XOR U1954 ( .A(n1657), .B(n1658), .Z(DIFF[216]) );
  XOR U1955 ( .A(B[216]), .B(A[216]), .Z(n1658) );
  AND U1956 ( .A(n1659), .B(n1660), .Z(n1657) );
  NANDN U1957 ( .A(B[215]), .B(n1661), .Z(n1660) );
  NANDN U1958 ( .A(A[215]), .B(n1662), .Z(n1661) );
  NANDN U1959 ( .A(n1662), .B(A[215]), .Z(n1659) );
  XOR U1960 ( .A(n1662), .B(n1663), .Z(DIFF[215]) );
  XOR U1961 ( .A(B[215]), .B(A[215]), .Z(n1663) );
  AND U1962 ( .A(n1664), .B(n1665), .Z(n1662) );
  NANDN U1963 ( .A(B[214]), .B(n1666), .Z(n1665) );
  NANDN U1964 ( .A(A[214]), .B(n1667), .Z(n1666) );
  NANDN U1965 ( .A(n1667), .B(A[214]), .Z(n1664) );
  XOR U1966 ( .A(n1667), .B(n1668), .Z(DIFF[214]) );
  XOR U1967 ( .A(B[214]), .B(A[214]), .Z(n1668) );
  AND U1968 ( .A(n1669), .B(n1670), .Z(n1667) );
  NANDN U1969 ( .A(B[213]), .B(n1671), .Z(n1670) );
  NANDN U1970 ( .A(A[213]), .B(n1672), .Z(n1671) );
  NANDN U1971 ( .A(n1672), .B(A[213]), .Z(n1669) );
  XOR U1972 ( .A(n1672), .B(n1673), .Z(DIFF[213]) );
  XOR U1973 ( .A(B[213]), .B(A[213]), .Z(n1673) );
  AND U1974 ( .A(n1674), .B(n1675), .Z(n1672) );
  NANDN U1975 ( .A(B[212]), .B(n1676), .Z(n1675) );
  NANDN U1976 ( .A(A[212]), .B(n1677), .Z(n1676) );
  NANDN U1977 ( .A(n1677), .B(A[212]), .Z(n1674) );
  XOR U1978 ( .A(n1677), .B(n1678), .Z(DIFF[212]) );
  XOR U1979 ( .A(B[212]), .B(A[212]), .Z(n1678) );
  AND U1980 ( .A(n1679), .B(n1680), .Z(n1677) );
  NANDN U1981 ( .A(B[211]), .B(n1681), .Z(n1680) );
  NANDN U1982 ( .A(A[211]), .B(n1682), .Z(n1681) );
  NANDN U1983 ( .A(n1682), .B(A[211]), .Z(n1679) );
  XOR U1984 ( .A(n1682), .B(n1683), .Z(DIFF[211]) );
  XOR U1985 ( .A(B[211]), .B(A[211]), .Z(n1683) );
  AND U1986 ( .A(n1684), .B(n1685), .Z(n1682) );
  NANDN U1987 ( .A(B[210]), .B(n1686), .Z(n1685) );
  NANDN U1988 ( .A(A[210]), .B(n1687), .Z(n1686) );
  NANDN U1989 ( .A(n1687), .B(A[210]), .Z(n1684) );
  XOR U1990 ( .A(n1687), .B(n1688), .Z(DIFF[210]) );
  XOR U1991 ( .A(B[210]), .B(A[210]), .Z(n1688) );
  AND U1992 ( .A(n1689), .B(n1690), .Z(n1687) );
  NANDN U1993 ( .A(B[209]), .B(n1691), .Z(n1690) );
  NANDN U1994 ( .A(A[209]), .B(n1692), .Z(n1691) );
  NANDN U1995 ( .A(n1692), .B(A[209]), .Z(n1689) );
  XOR U1996 ( .A(n1693), .B(n1694), .Z(DIFF[20]) );
  XOR U1997 ( .A(B[20]), .B(A[20]), .Z(n1694) );
  XOR U1998 ( .A(n1692), .B(n1695), .Z(DIFF[209]) );
  XOR U1999 ( .A(B[209]), .B(A[209]), .Z(n1695) );
  AND U2000 ( .A(n1696), .B(n1697), .Z(n1692) );
  NANDN U2001 ( .A(B[208]), .B(n1698), .Z(n1697) );
  NANDN U2002 ( .A(A[208]), .B(n1699), .Z(n1698) );
  NANDN U2003 ( .A(n1699), .B(A[208]), .Z(n1696) );
  XOR U2004 ( .A(n1699), .B(n1700), .Z(DIFF[208]) );
  XOR U2005 ( .A(B[208]), .B(A[208]), .Z(n1700) );
  AND U2006 ( .A(n1701), .B(n1702), .Z(n1699) );
  NANDN U2007 ( .A(B[207]), .B(n1703), .Z(n1702) );
  NANDN U2008 ( .A(A[207]), .B(n1704), .Z(n1703) );
  NANDN U2009 ( .A(n1704), .B(A[207]), .Z(n1701) );
  XOR U2010 ( .A(n1704), .B(n1705), .Z(DIFF[207]) );
  XOR U2011 ( .A(B[207]), .B(A[207]), .Z(n1705) );
  AND U2012 ( .A(n1706), .B(n1707), .Z(n1704) );
  NANDN U2013 ( .A(B[206]), .B(n1708), .Z(n1707) );
  NANDN U2014 ( .A(A[206]), .B(n1709), .Z(n1708) );
  NANDN U2015 ( .A(n1709), .B(A[206]), .Z(n1706) );
  XOR U2016 ( .A(n1709), .B(n1710), .Z(DIFF[206]) );
  XOR U2017 ( .A(B[206]), .B(A[206]), .Z(n1710) );
  AND U2018 ( .A(n1711), .B(n1712), .Z(n1709) );
  NANDN U2019 ( .A(B[205]), .B(n1713), .Z(n1712) );
  NANDN U2020 ( .A(A[205]), .B(n1714), .Z(n1713) );
  NANDN U2021 ( .A(n1714), .B(A[205]), .Z(n1711) );
  XOR U2022 ( .A(n1714), .B(n1715), .Z(DIFF[205]) );
  XOR U2023 ( .A(B[205]), .B(A[205]), .Z(n1715) );
  AND U2024 ( .A(n1716), .B(n1717), .Z(n1714) );
  NANDN U2025 ( .A(B[204]), .B(n1718), .Z(n1717) );
  NANDN U2026 ( .A(A[204]), .B(n1719), .Z(n1718) );
  NANDN U2027 ( .A(n1719), .B(A[204]), .Z(n1716) );
  XOR U2028 ( .A(n1719), .B(n1720), .Z(DIFF[204]) );
  XOR U2029 ( .A(B[204]), .B(A[204]), .Z(n1720) );
  AND U2030 ( .A(n1721), .B(n1722), .Z(n1719) );
  NANDN U2031 ( .A(B[203]), .B(n1723), .Z(n1722) );
  NANDN U2032 ( .A(A[203]), .B(n1724), .Z(n1723) );
  NANDN U2033 ( .A(n1724), .B(A[203]), .Z(n1721) );
  XOR U2034 ( .A(n1724), .B(n1725), .Z(DIFF[203]) );
  XOR U2035 ( .A(B[203]), .B(A[203]), .Z(n1725) );
  AND U2036 ( .A(n1726), .B(n1727), .Z(n1724) );
  NANDN U2037 ( .A(B[202]), .B(n1728), .Z(n1727) );
  NANDN U2038 ( .A(A[202]), .B(n1729), .Z(n1728) );
  NANDN U2039 ( .A(n1729), .B(A[202]), .Z(n1726) );
  XOR U2040 ( .A(n1729), .B(n1730), .Z(DIFF[202]) );
  XOR U2041 ( .A(B[202]), .B(A[202]), .Z(n1730) );
  AND U2042 ( .A(n1731), .B(n1732), .Z(n1729) );
  NANDN U2043 ( .A(B[201]), .B(n1733), .Z(n1732) );
  NANDN U2044 ( .A(A[201]), .B(n1734), .Z(n1733) );
  NANDN U2045 ( .A(n1734), .B(A[201]), .Z(n1731) );
  XOR U2046 ( .A(n1734), .B(n1735), .Z(DIFF[201]) );
  XOR U2047 ( .A(B[201]), .B(A[201]), .Z(n1735) );
  AND U2048 ( .A(n1736), .B(n1737), .Z(n1734) );
  NANDN U2049 ( .A(B[200]), .B(n1738), .Z(n1737) );
  NANDN U2050 ( .A(A[200]), .B(n1739), .Z(n1738) );
  NANDN U2051 ( .A(n1739), .B(A[200]), .Z(n1736) );
  XOR U2052 ( .A(n1739), .B(n1740), .Z(DIFF[200]) );
  XOR U2053 ( .A(B[200]), .B(A[200]), .Z(n1740) );
  AND U2054 ( .A(n1741), .B(n1742), .Z(n1739) );
  NANDN U2055 ( .A(B[199]), .B(n1743), .Z(n1742) );
  NANDN U2056 ( .A(A[199]), .B(n1744), .Z(n1743) );
  NANDN U2057 ( .A(n1744), .B(A[199]), .Z(n1741) );
  XOR U2058 ( .A(n1), .B(n1745), .Z(DIFF[1]) );
  XOR U2059 ( .A(B[1]), .B(A[1]), .Z(n1745) );
  XOR U2060 ( .A(n1746), .B(n1747), .Z(DIFF[19]) );
  XOR U2061 ( .A(B[19]), .B(A[19]), .Z(n1747) );
  XOR U2062 ( .A(n1744), .B(n1748), .Z(DIFF[199]) );
  XOR U2063 ( .A(B[199]), .B(A[199]), .Z(n1748) );
  AND U2064 ( .A(n1749), .B(n1750), .Z(n1744) );
  NANDN U2065 ( .A(B[198]), .B(n1751), .Z(n1750) );
  NANDN U2066 ( .A(A[198]), .B(n1752), .Z(n1751) );
  NANDN U2067 ( .A(n1752), .B(A[198]), .Z(n1749) );
  XOR U2068 ( .A(n1752), .B(n1753), .Z(DIFF[198]) );
  XOR U2069 ( .A(B[198]), .B(A[198]), .Z(n1753) );
  AND U2070 ( .A(n1754), .B(n1755), .Z(n1752) );
  NANDN U2071 ( .A(B[197]), .B(n1756), .Z(n1755) );
  NANDN U2072 ( .A(A[197]), .B(n1757), .Z(n1756) );
  NANDN U2073 ( .A(n1757), .B(A[197]), .Z(n1754) );
  XOR U2074 ( .A(n1757), .B(n1758), .Z(DIFF[197]) );
  XOR U2075 ( .A(B[197]), .B(A[197]), .Z(n1758) );
  AND U2076 ( .A(n1759), .B(n1760), .Z(n1757) );
  NANDN U2077 ( .A(B[196]), .B(n1761), .Z(n1760) );
  NANDN U2078 ( .A(A[196]), .B(n1762), .Z(n1761) );
  NANDN U2079 ( .A(n1762), .B(A[196]), .Z(n1759) );
  XOR U2080 ( .A(n1762), .B(n1763), .Z(DIFF[196]) );
  XOR U2081 ( .A(B[196]), .B(A[196]), .Z(n1763) );
  AND U2082 ( .A(n1764), .B(n1765), .Z(n1762) );
  NANDN U2083 ( .A(B[195]), .B(n1766), .Z(n1765) );
  NANDN U2084 ( .A(A[195]), .B(n1767), .Z(n1766) );
  NANDN U2085 ( .A(n1767), .B(A[195]), .Z(n1764) );
  XOR U2086 ( .A(n1767), .B(n1768), .Z(DIFF[195]) );
  XOR U2087 ( .A(B[195]), .B(A[195]), .Z(n1768) );
  AND U2088 ( .A(n1769), .B(n1770), .Z(n1767) );
  NANDN U2089 ( .A(B[194]), .B(n1771), .Z(n1770) );
  NANDN U2090 ( .A(A[194]), .B(n1772), .Z(n1771) );
  NANDN U2091 ( .A(n1772), .B(A[194]), .Z(n1769) );
  XOR U2092 ( .A(n1772), .B(n1773), .Z(DIFF[194]) );
  XOR U2093 ( .A(B[194]), .B(A[194]), .Z(n1773) );
  AND U2094 ( .A(n1774), .B(n1775), .Z(n1772) );
  NANDN U2095 ( .A(B[193]), .B(n1776), .Z(n1775) );
  NANDN U2096 ( .A(A[193]), .B(n1777), .Z(n1776) );
  NANDN U2097 ( .A(n1777), .B(A[193]), .Z(n1774) );
  XOR U2098 ( .A(n1777), .B(n1778), .Z(DIFF[193]) );
  XOR U2099 ( .A(B[193]), .B(A[193]), .Z(n1778) );
  AND U2100 ( .A(n1779), .B(n1780), .Z(n1777) );
  NANDN U2101 ( .A(B[192]), .B(n1781), .Z(n1780) );
  NANDN U2102 ( .A(A[192]), .B(n1782), .Z(n1781) );
  NANDN U2103 ( .A(n1782), .B(A[192]), .Z(n1779) );
  XOR U2104 ( .A(n1782), .B(n1783), .Z(DIFF[192]) );
  XOR U2105 ( .A(B[192]), .B(A[192]), .Z(n1783) );
  AND U2106 ( .A(n1784), .B(n1785), .Z(n1782) );
  NANDN U2107 ( .A(B[191]), .B(n1786), .Z(n1785) );
  NANDN U2108 ( .A(A[191]), .B(n1787), .Z(n1786) );
  NANDN U2109 ( .A(n1787), .B(A[191]), .Z(n1784) );
  XOR U2110 ( .A(n1787), .B(n1788), .Z(DIFF[191]) );
  XOR U2111 ( .A(B[191]), .B(A[191]), .Z(n1788) );
  AND U2112 ( .A(n1789), .B(n1790), .Z(n1787) );
  NANDN U2113 ( .A(B[190]), .B(n1791), .Z(n1790) );
  NANDN U2114 ( .A(A[190]), .B(n1792), .Z(n1791) );
  NANDN U2115 ( .A(n1792), .B(A[190]), .Z(n1789) );
  XOR U2116 ( .A(n1792), .B(n1793), .Z(DIFF[190]) );
  XOR U2117 ( .A(B[190]), .B(A[190]), .Z(n1793) );
  AND U2118 ( .A(n1794), .B(n1795), .Z(n1792) );
  NANDN U2119 ( .A(B[189]), .B(n1796), .Z(n1795) );
  NANDN U2120 ( .A(A[189]), .B(n1797), .Z(n1796) );
  NANDN U2121 ( .A(n1797), .B(A[189]), .Z(n1794) );
  XOR U2122 ( .A(n1798), .B(n1799), .Z(DIFF[18]) );
  XOR U2123 ( .A(B[18]), .B(A[18]), .Z(n1799) );
  XOR U2124 ( .A(n1797), .B(n1800), .Z(DIFF[189]) );
  XOR U2125 ( .A(B[189]), .B(A[189]), .Z(n1800) );
  AND U2126 ( .A(n1801), .B(n1802), .Z(n1797) );
  NANDN U2127 ( .A(B[188]), .B(n1803), .Z(n1802) );
  NANDN U2128 ( .A(A[188]), .B(n1804), .Z(n1803) );
  NANDN U2129 ( .A(n1804), .B(A[188]), .Z(n1801) );
  XOR U2130 ( .A(n1804), .B(n1805), .Z(DIFF[188]) );
  XOR U2131 ( .A(B[188]), .B(A[188]), .Z(n1805) );
  AND U2132 ( .A(n1806), .B(n1807), .Z(n1804) );
  NANDN U2133 ( .A(B[187]), .B(n1808), .Z(n1807) );
  NANDN U2134 ( .A(A[187]), .B(n1809), .Z(n1808) );
  NANDN U2135 ( .A(n1809), .B(A[187]), .Z(n1806) );
  XOR U2136 ( .A(n1809), .B(n1810), .Z(DIFF[187]) );
  XOR U2137 ( .A(B[187]), .B(A[187]), .Z(n1810) );
  AND U2138 ( .A(n1811), .B(n1812), .Z(n1809) );
  NANDN U2139 ( .A(B[186]), .B(n1813), .Z(n1812) );
  NANDN U2140 ( .A(A[186]), .B(n1814), .Z(n1813) );
  NANDN U2141 ( .A(n1814), .B(A[186]), .Z(n1811) );
  XOR U2142 ( .A(n1814), .B(n1815), .Z(DIFF[186]) );
  XOR U2143 ( .A(B[186]), .B(A[186]), .Z(n1815) );
  AND U2144 ( .A(n1816), .B(n1817), .Z(n1814) );
  NANDN U2145 ( .A(B[185]), .B(n1818), .Z(n1817) );
  NANDN U2146 ( .A(A[185]), .B(n1819), .Z(n1818) );
  NANDN U2147 ( .A(n1819), .B(A[185]), .Z(n1816) );
  XOR U2148 ( .A(n1819), .B(n1820), .Z(DIFF[185]) );
  XOR U2149 ( .A(B[185]), .B(A[185]), .Z(n1820) );
  AND U2150 ( .A(n1821), .B(n1822), .Z(n1819) );
  NANDN U2151 ( .A(B[184]), .B(n1823), .Z(n1822) );
  NANDN U2152 ( .A(A[184]), .B(n1824), .Z(n1823) );
  NANDN U2153 ( .A(n1824), .B(A[184]), .Z(n1821) );
  XOR U2154 ( .A(n1824), .B(n1825), .Z(DIFF[184]) );
  XOR U2155 ( .A(B[184]), .B(A[184]), .Z(n1825) );
  AND U2156 ( .A(n1826), .B(n1827), .Z(n1824) );
  NANDN U2157 ( .A(B[183]), .B(n1828), .Z(n1827) );
  NANDN U2158 ( .A(A[183]), .B(n1829), .Z(n1828) );
  NANDN U2159 ( .A(n1829), .B(A[183]), .Z(n1826) );
  XOR U2160 ( .A(n1829), .B(n1830), .Z(DIFF[183]) );
  XOR U2161 ( .A(B[183]), .B(A[183]), .Z(n1830) );
  AND U2162 ( .A(n1831), .B(n1832), .Z(n1829) );
  NANDN U2163 ( .A(B[182]), .B(n1833), .Z(n1832) );
  NANDN U2164 ( .A(A[182]), .B(n1834), .Z(n1833) );
  NANDN U2165 ( .A(n1834), .B(A[182]), .Z(n1831) );
  XOR U2166 ( .A(n1834), .B(n1835), .Z(DIFF[182]) );
  XOR U2167 ( .A(B[182]), .B(A[182]), .Z(n1835) );
  AND U2168 ( .A(n1836), .B(n1837), .Z(n1834) );
  NANDN U2169 ( .A(B[181]), .B(n1838), .Z(n1837) );
  NANDN U2170 ( .A(A[181]), .B(n1839), .Z(n1838) );
  NANDN U2171 ( .A(n1839), .B(A[181]), .Z(n1836) );
  XOR U2172 ( .A(n1839), .B(n1840), .Z(DIFF[181]) );
  XOR U2173 ( .A(B[181]), .B(A[181]), .Z(n1840) );
  AND U2174 ( .A(n1841), .B(n1842), .Z(n1839) );
  NANDN U2175 ( .A(B[180]), .B(n1843), .Z(n1842) );
  NANDN U2176 ( .A(A[180]), .B(n1844), .Z(n1843) );
  NANDN U2177 ( .A(n1844), .B(A[180]), .Z(n1841) );
  XOR U2178 ( .A(n1844), .B(n1845), .Z(DIFF[180]) );
  XOR U2179 ( .A(B[180]), .B(A[180]), .Z(n1845) );
  AND U2180 ( .A(n1846), .B(n1847), .Z(n1844) );
  NANDN U2181 ( .A(B[179]), .B(n1848), .Z(n1847) );
  NANDN U2182 ( .A(A[179]), .B(n1849), .Z(n1848) );
  NANDN U2183 ( .A(n1849), .B(A[179]), .Z(n1846) );
  XOR U2184 ( .A(n1850), .B(n1851), .Z(DIFF[17]) );
  XOR U2185 ( .A(B[17]), .B(A[17]), .Z(n1851) );
  XOR U2186 ( .A(n1849), .B(n1852), .Z(DIFF[179]) );
  XOR U2187 ( .A(B[179]), .B(A[179]), .Z(n1852) );
  AND U2188 ( .A(n1853), .B(n1854), .Z(n1849) );
  NANDN U2189 ( .A(B[178]), .B(n1855), .Z(n1854) );
  NANDN U2190 ( .A(A[178]), .B(n1856), .Z(n1855) );
  NANDN U2191 ( .A(n1856), .B(A[178]), .Z(n1853) );
  XOR U2192 ( .A(n1856), .B(n1857), .Z(DIFF[178]) );
  XOR U2193 ( .A(B[178]), .B(A[178]), .Z(n1857) );
  AND U2194 ( .A(n1858), .B(n1859), .Z(n1856) );
  NANDN U2195 ( .A(B[177]), .B(n1860), .Z(n1859) );
  NANDN U2196 ( .A(A[177]), .B(n1861), .Z(n1860) );
  NANDN U2197 ( .A(n1861), .B(A[177]), .Z(n1858) );
  XOR U2198 ( .A(n1861), .B(n1862), .Z(DIFF[177]) );
  XOR U2199 ( .A(B[177]), .B(A[177]), .Z(n1862) );
  AND U2200 ( .A(n1863), .B(n1864), .Z(n1861) );
  NANDN U2201 ( .A(B[176]), .B(n1865), .Z(n1864) );
  NANDN U2202 ( .A(A[176]), .B(n1866), .Z(n1865) );
  NANDN U2203 ( .A(n1866), .B(A[176]), .Z(n1863) );
  XOR U2204 ( .A(n1866), .B(n1867), .Z(DIFF[176]) );
  XOR U2205 ( .A(B[176]), .B(A[176]), .Z(n1867) );
  AND U2206 ( .A(n1868), .B(n1869), .Z(n1866) );
  NANDN U2207 ( .A(B[175]), .B(n1870), .Z(n1869) );
  NANDN U2208 ( .A(A[175]), .B(n1871), .Z(n1870) );
  NANDN U2209 ( .A(n1871), .B(A[175]), .Z(n1868) );
  XOR U2210 ( .A(n1871), .B(n1872), .Z(DIFF[175]) );
  XOR U2211 ( .A(B[175]), .B(A[175]), .Z(n1872) );
  AND U2212 ( .A(n1873), .B(n1874), .Z(n1871) );
  NANDN U2213 ( .A(B[174]), .B(n1875), .Z(n1874) );
  NANDN U2214 ( .A(A[174]), .B(n1876), .Z(n1875) );
  NANDN U2215 ( .A(n1876), .B(A[174]), .Z(n1873) );
  XOR U2216 ( .A(n1876), .B(n1877), .Z(DIFF[174]) );
  XOR U2217 ( .A(B[174]), .B(A[174]), .Z(n1877) );
  AND U2218 ( .A(n1878), .B(n1879), .Z(n1876) );
  NANDN U2219 ( .A(B[173]), .B(n1880), .Z(n1879) );
  NANDN U2220 ( .A(A[173]), .B(n1881), .Z(n1880) );
  NANDN U2221 ( .A(n1881), .B(A[173]), .Z(n1878) );
  XOR U2222 ( .A(n1881), .B(n1882), .Z(DIFF[173]) );
  XOR U2223 ( .A(B[173]), .B(A[173]), .Z(n1882) );
  AND U2224 ( .A(n1883), .B(n1884), .Z(n1881) );
  NANDN U2225 ( .A(B[172]), .B(n1885), .Z(n1884) );
  NANDN U2226 ( .A(A[172]), .B(n1886), .Z(n1885) );
  NANDN U2227 ( .A(n1886), .B(A[172]), .Z(n1883) );
  XOR U2228 ( .A(n1886), .B(n1887), .Z(DIFF[172]) );
  XOR U2229 ( .A(B[172]), .B(A[172]), .Z(n1887) );
  AND U2230 ( .A(n1888), .B(n1889), .Z(n1886) );
  NANDN U2231 ( .A(B[171]), .B(n1890), .Z(n1889) );
  NANDN U2232 ( .A(A[171]), .B(n1891), .Z(n1890) );
  NANDN U2233 ( .A(n1891), .B(A[171]), .Z(n1888) );
  XOR U2234 ( .A(n1891), .B(n1892), .Z(DIFF[171]) );
  XOR U2235 ( .A(B[171]), .B(A[171]), .Z(n1892) );
  AND U2236 ( .A(n1893), .B(n1894), .Z(n1891) );
  NANDN U2237 ( .A(B[170]), .B(n1895), .Z(n1894) );
  NANDN U2238 ( .A(A[170]), .B(n1896), .Z(n1895) );
  NANDN U2239 ( .A(n1896), .B(A[170]), .Z(n1893) );
  XOR U2240 ( .A(n1896), .B(n1897), .Z(DIFF[170]) );
  XOR U2241 ( .A(B[170]), .B(A[170]), .Z(n1897) );
  AND U2242 ( .A(n1898), .B(n1899), .Z(n1896) );
  NANDN U2243 ( .A(B[169]), .B(n1900), .Z(n1899) );
  NANDN U2244 ( .A(A[169]), .B(n1901), .Z(n1900) );
  NANDN U2245 ( .A(n1901), .B(A[169]), .Z(n1898) );
  XOR U2246 ( .A(n1902), .B(n1903), .Z(DIFF[16]) );
  XOR U2247 ( .A(B[16]), .B(A[16]), .Z(n1903) );
  XOR U2248 ( .A(n1901), .B(n1904), .Z(DIFF[169]) );
  XOR U2249 ( .A(B[169]), .B(A[169]), .Z(n1904) );
  AND U2250 ( .A(n1905), .B(n1906), .Z(n1901) );
  NANDN U2251 ( .A(B[168]), .B(n1907), .Z(n1906) );
  NANDN U2252 ( .A(A[168]), .B(n1908), .Z(n1907) );
  NANDN U2253 ( .A(n1908), .B(A[168]), .Z(n1905) );
  XOR U2254 ( .A(n1908), .B(n1909), .Z(DIFF[168]) );
  XOR U2255 ( .A(B[168]), .B(A[168]), .Z(n1909) );
  AND U2256 ( .A(n1910), .B(n1911), .Z(n1908) );
  NANDN U2257 ( .A(B[167]), .B(n1912), .Z(n1911) );
  NANDN U2258 ( .A(A[167]), .B(n1913), .Z(n1912) );
  NANDN U2259 ( .A(n1913), .B(A[167]), .Z(n1910) );
  XOR U2260 ( .A(n1913), .B(n1914), .Z(DIFF[167]) );
  XOR U2261 ( .A(B[167]), .B(A[167]), .Z(n1914) );
  AND U2262 ( .A(n1915), .B(n1916), .Z(n1913) );
  NANDN U2263 ( .A(B[166]), .B(n1917), .Z(n1916) );
  NANDN U2264 ( .A(A[166]), .B(n1918), .Z(n1917) );
  NANDN U2265 ( .A(n1918), .B(A[166]), .Z(n1915) );
  XOR U2266 ( .A(n1918), .B(n1919), .Z(DIFF[166]) );
  XOR U2267 ( .A(B[166]), .B(A[166]), .Z(n1919) );
  AND U2268 ( .A(n1920), .B(n1921), .Z(n1918) );
  NANDN U2269 ( .A(B[165]), .B(n1922), .Z(n1921) );
  NANDN U2270 ( .A(A[165]), .B(n1923), .Z(n1922) );
  NANDN U2271 ( .A(n1923), .B(A[165]), .Z(n1920) );
  XOR U2272 ( .A(n1923), .B(n1924), .Z(DIFF[165]) );
  XOR U2273 ( .A(B[165]), .B(A[165]), .Z(n1924) );
  AND U2274 ( .A(n1925), .B(n1926), .Z(n1923) );
  NANDN U2275 ( .A(B[164]), .B(n1927), .Z(n1926) );
  NANDN U2276 ( .A(A[164]), .B(n1928), .Z(n1927) );
  NANDN U2277 ( .A(n1928), .B(A[164]), .Z(n1925) );
  XOR U2278 ( .A(n1928), .B(n1929), .Z(DIFF[164]) );
  XOR U2279 ( .A(B[164]), .B(A[164]), .Z(n1929) );
  AND U2280 ( .A(n1930), .B(n1931), .Z(n1928) );
  NANDN U2281 ( .A(B[163]), .B(n1932), .Z(n1931) );
  NANDN U2282 ( .A(A[163]), .B(n1933), .Z(n1932) );
  NANDN U2283 ( .A(n1933), .B(A[163]), .Z(n1930) );
  XOR U2284 ( .A(n1933), .B(n1934), .Z(DIFF[163]) );
  XOR U2285 ( .A(B[163]), .B(A[163]), .Z(n1934) );
  AND U2286 ( .A(n1935), .B(n1936), .Z(n1933) );
  NANDN U2287 ( .A(B[162]), .B(n1937), .Z(n1936) );
  NANDN U2288 ( .A(A[162]), .B(n1938), .Z(n1937) );
  NANDN U2289 ( .A(n1938), .B(A[162]), .Z(n1935) );
  XOR U2290 ( .A(n1938), .B(n1939), .Z(DIFF[162]) );
  XOR U2291 ( .A(B[162]), .B(A[162]), .Z(n1939) );
  AND U2292 ( .A(n1940), .B(n1941), .Z(n1938) );
  NANDN U2293 ( .A(B[161]), .B(n1942), .Z(n1941) );
  NANDN U2294 ( .A(A[161]), .B(n1943), .Z(n1942) );
  NANDN U2295 ( .A(n1943), .B(A[161]), .Z(n1940) );
  XOR U2296 ( .A(n1943), .B(n1944), .Z(DIFF[161]) );
  XOR U2297 ( .A(B[161]), .B(A[161]), .Z(n1944) );
  AND U2298 ( .A(n1945), .B(n1946), .Z(n1943) );
  NANDN U2299 ( .A(B[160]), .B(n1947), .Z(n1946) );
  NANDN U2300 ( .A(A[160]), .B(n1948), .Z(n1947) );
  NANDN U2301 ( .A(n1948), .B(A[160]), .Z(n1945) );
  XOR U2302 ( .A(n1948), .B(n1949), .Z(DIFF[160]) );
  XOR U2303 ( .A(B[160]), .B(A[160]), .Z(n1949) );
  AND U2304 ( .A(n1950), .B(n1951), .Z(n1948) );
  NANDN U2305 ( .A(B[159]), .B(n1952), .Z(n1951) );
  NANDN U2306 ( .A(A[159]), .B(n1953), .Z(n1952) );
  NANDN U2307 ( .A(n1953), .B(A[159]), .Z(n1950) );
  XOR U2308 ( .A(n1954), .B(n1955), .Z(DIFF[15]) );
  XOR U2309 ( .A(B[15]), .B(A[15]), .Z(n1955) );
  XOR U2310 ( .A(n1953), .B(n1956), .Z(DIFF[159]) );
  XOR U2311 ( .A(B[159]), .B(A[159]), .Z(n1956) );
  AND U2312 ( .A(n1957), .B(n1958), .Z(n1953) );
  NANDN U2313 ( .A(B[158]), .B(n1959), .Z(n1958) );
  NANDN U2314 ( .A(A[158]), .B(n1960), .Z(n1959) );
  NANDN U2315 ( .A(n1960), .B(A[158]), .Z(n1957) );
  XOR U2316 ( .A(n1960), .B(n1961), .Z(DIFF[158]) );
  XOR U2317 ( .A(B[158]), .B(A[158]), .Z(n1961) );
  AND U2318 ( .A(n1962), .B(n1963), .Z(n1960) );
  NANDN U2319 ( .A(B[157]), .B(n1964), .Z(n1963) );
  NANDN U2320 ( .A(A[157]), .B(n1965), .Z(n1964) );
  NANDN U2321 ( .A(n1965), .B(A[157]), .Z(n1962) );
  XOR U2322 ( .A(n1965), .B(n1966), .Z(DIFF[157]) );
  XOR U2323 ( .A(B[157]), .B(A[157]), .Z(n1966) );
  AND U2324 ( .A(n1967), .B(n1968), .Z(n1965) );
  NANDN U2325 ( .A(B[156]), .B(n1969), .Z(n1968) );
  NANDN U2326 ( .A(A[156]), .B(n1970), .Z(n1969) );
  NANDN U2327 ( .A(n1970), .B(A[156]), .Z(n1967) );
  XOR U2328 ( .A(n1970), .B(n1971), .Z(DIFF[156]) );
  XOR U2329 ( .A(B[156]), .B(A[156]), .Z(n1971) );
  AND U2330 ( .A(n1972), .B(n1973), .Z(n1970) );
  NANDN U2331 ( .A(B[155]), .B(n1974), .Z(n1973) );
  NANDN U2332 ( .A(A[155]), .B(n1975), .Z(n1974) );
  NANDN U2333 ( .A(n1975), .B(A[155]), .Z(n1972) );
  XOR U2334 ( .A(n1975), .B(n1976), .Z(DIFF[155]) );
  XOR U2335 ( .A(B[155]), .B(A[155]), .Z(n1976) );
  AND U2336 ( .A(n1977), .B(n1978), .Z(n1975) );
  NANDN U2337 ( .A(B[154]), .B(n1979), .Z(n1978) );
  NANDN U2338 ( .A(A[154]), .B(n1980), .Z(n1979) );
  NANDN U2339 ( .A(n1980), .B(A[154]), .Z(n1977) );
  XOR U2340 ( .A(n1980), .B(n1981), .Z(DIFF[154]) );
  XOR U2341 ( .A(B[154]), .B(A[154]), .Z(n1981) );
  AND U2342 ( .A(n1982), .B(n1983), .Z(n1980) );
  NANDN U2343 ( .A(B[153]), .B(n1984), .Z(n1983) );
  NANDN U2344 ( .A(A[153]), .B(n1985), .Z(n1984) );
  NANDN U2345 ( .A(n1985), .B(A[153]), .Z(n1982) );
  XOR U2346 ( .A(n1985), .B(n1986), .Z(DIFF[153]) );
  XOR U2347 ( .A(B[153]), .B(A[153]), .Z(n1986) );
  AND U2348 ( .A(n1987), .B(n1988), .Z(n1985) );
  NANDN U2349 ( .A(B[152]), .B(n1989), .Z(n1988) );
  NANDN U2350 ( .A(A[152]), .B(n1990), .Z(n1989) );
  NANDN U2351 ( .A(n1990), .B(A[152]), .Z(n1987) );
  XOR U2352 ( .A(n1990), .B(n1991), .Z(DIFF[152]) );
  XOR U2353 ( .A(B[152]), .B(A[152]), .Z(n1991) );
  AND U2354 ( .A(n1992), .B(n1993), .Z(n1990) );
  NANDN U2355 ( .A(B[151]), .B(n1994), .Z(n1993) );
  NANDN U2356 ( .A(A[151]), .B(n1995), .Z(n1994) );
  NANDN U2357 ( .A(n1995), .B(A[151]), .Z(n1992) );
  XOR U2358 ( .A(n1995), .B(n1996), .Z(DIFF[151]) );
  XOR U2359 ( .A(B[151]), .B(A[151]), .Z(n1996) );
  AND U2360 ( .A(n1997), .B(n1998), .Z(n1995) );
  NANDN U2361 ( .A(B[150]), .B(n1999), .Z(n1998) );
  NANDN U2362 ( .A(A[150]), .B(n2000), .Z(n1999) );
  NANDN U2363 ( .A(n2000), .B(A[150]), .Z(n1997) );
  XOR U2364 ( .A(n2000), .B(n2001), .Z(DIFF[150]) );
  XOR U2365 ( .A(B[150]), .B(A[150]), .Z(n2001) );
  AND U2366 ( .A(n2002), .B(n2003), .Z(n2000) );
  NANDN U2367 ( .A(B[149]), .B(n2004), .Z(n2003) );
  NANDN U2368 ( .A(A[149]), .B(n2005), .Z(n2004) );
  NANDN U2369 ( .A(n2005), .B(A[149]), .Z(n2002) );
  XOR U2370 ( .A(n2006), .B(n2007), .Z(DIFF[14]) );
  XOR U2371 ( .A(B[14]), .B(A[14]), .Z(n2007) );
  XOR U2372 ( .A(n2005), .B(n2008), .Z(DIFF[149]) );
  XOR U2373 ( .A(B[149]), .B(A[149]), .Z(n2008) );
  AND U2374 ( .A(n2009), .B(n2010), .Z(n2005) );
  NANDN U2375 ( .A(B[148]), .B(n2011), .Z(n2010) );
  NANDN U2376 ( .A(A[148]), .B(n2012), .Z(n2011) );
  NANDN U2377 ( .A(n2012), .B(A[148]), .Z(n2009) );
  XOR U2378 ( .A(n2012), .B(n2013), .Z(DIFF[148]) );
  XOR U2379 ( .A(B[148]), .B(A[148]), .Z(n2013) );
  AND U2380 ( .A(n2014), .B(n2015), .Z(n2012) );
  NANDN U2381 ( .A(B[147]), .B(n2016), .Z(n2015) );
  NANDN U2382 ( .A(A[147]), .B(n2017), .Z(n2016) );
  NANDN U2383 ( .A(n2017), .B(A[147]), .Z(n2014) );
  XOR U2384 ( .A(n2017), .B(n2018), .Z(DIFF[147]) );
  XOR U2385 ( .A(B[147]), .B(A[147]), .Z(n2018) );
  AND U2386 ( .A(n2019), .B(n2020), .Z(n2017) );
  NANDN U2387 ( .A(B[146]), .B(n2021), .Z(n2020) );
  NANDN U2388 ( .A(A[146]), .B(n2022), .Z(n2021) );
  NANDN U2389 ( .A(n2022), .B(A[146]), .Z(n2019) );
  XOR U2390 ( .A(n2022), .B(n2023), .Z(DIFF[146]) );
  XOR U2391 ( .A(B[146]), .B(A[146]), .Z(n2023) );
  AND U2392 ( .A(n2024), .B(n2025), .Z(n2022) );
  NANDN U2393 ( .A(B[145]), .B(n2026), .Z(n2025) );
  NANDN U2394 ( .A(A[145]), .B(n2027), .Z(n2026) );
  NANDN U2395 ( .A(n2027), .B(A[145]), .Z(n2024) );
  XOR U2396 ( .A(n2027), .B(n2028), .Z(DIFF[145]) );
  XOR U2397 ( .A(B[145]), .B(A[145]), .Z(n2028) );
  AND U2398 ( .A(n2029), .B(n2030), .Z(n2027) );
  NANDN U2399 ( .A(B[144]), .B(n2031), .Z(n2030) );
  NANDN U2400 ( .A(A[144]), .B(n2032), .Z(n2031) );
  NANDN U2401 ( .A(n2032), .B(A[144]), .Z(n2029) );
  XOR U2402 ( .A(n2032), .B(n2033), .Z(DIFF[144]) );
  XOR U2403 ( .A(B[144]), .B(A[144]), .Z(n2033) );
  AND U2404 ( .A(n2034), .B(n2035), .Z(n2032) );
  NANDN U2405 ( .A(B[143]), .B(n2036), .Z(n2035) );
  NANDN U2406 ( .A(A[143]), .B(n2037), .Z(n2036) );
  NANDN U2407 ( .A(n2037), .B(A[143]), .Z(n2034) );
  XOR U2408 ( .A(n2037), .B(n2038), .Z(DIFF[143]) );
  XOR U2409 ( .A(B[143]), .B(A[143]), .Z(n2038) );
  AND U2410 ( .A(n2039), .B(n2040), .Z(n2037) );
  NANDN U2411 ( .A(B[142]), .B(n2041), .Z(n2040) );
  NANDN U2412 ( .A(A[142]), .B(n2042), .Z(n2041) );
  NANDN U2413 ( .A(n2042), .B(A[142]), .Z(n2039) );
  XOR U2414 ( .A(n2042), .B(n2043), .Z(DIFF[142]) );
  XOR U2415 ( .A(B[142]), .B(A[142]), .Z(n2043) );
  AND U2416 ( .A(n2044), .B(n2045), .Z(n2042) );
  NANDN U2417 ( .A(B[141]), .B(n2046), .Z(n2045) );
  NANDN U2418 ( .A(A[141]), .B(n2047), .Z(n2046) );
  NANDN U2419 ( .A(n2047), .B(A[141]), .Z(n2044) );
  XOR U2420 ( .A(n2047), .B(n2048), .Z(DIFF[141]) );
  XOR U2421 ( .A(B[141]), .B(A[141]), .Z(n2048) );
  AND U2422 ( .A(n2049), .B(n2050), .Z(n2047) );
  NANDN U2423 ( .A(B[140]), .B(n2051), .Z(n2050) );
  NANDN U2424 ( .A(A[140]), .B(n2052), .Z(n2051) );
  NANDN U2425 ( .A(n2052), .B(A[140]), .Z(n2049) );
  XOR U2426 ( .A(n2052), .B(n2053), .Z(DIFF[140]) );
  XOR U2427 ( .A(B[140]), .B(A[140]), .Z(n2053) );
  AND U2428 ( .A(n2054), .B(n2055), .Z(n2052) );
  NANDN U2429 ( .A(B[139]), .B(n2056), .Z(n2055) );
  NANDN U2430 ( .A(A[139]), .B(n2057), .Z(n2056) );
  NANDN U2431 ( .A(n2057), .B(A[139]), .Z(n2054) );
  XOR U2432 ( .A(n2058), .B(n2059), .Z(DIFF[13]) );
  XOR U2433 ( .A(B[13]), .B(A[13]), .Z(n2059) );
  XOR U2434 ( .A(n2057), .B(n2060), .Z(DIFF[139]) );
  XOR U2435 ( .A(B[139]), .B(A[139]), .Z(n2060) );
  AND U2436 ( .A(n2061), .B(n2062), .Z(n2057) );
  NANDN U2437 ( .A(B[138]), .B(n2063), .Z(n2062) );
  NANDN U2438 ( .A(A[138]), .B(n2064), .Z(n2063) );
  NANDN U2439 ( .A(n2064), .B(A[138]), .Z(n2061) );
  XOR U2440 ( .A(n2064), .B(n2065), .Z(DIFF[138]) );
  XOR U2441 ( .A(B[138]), .B(A[138]), .Z(n2065) );
  AND U2442 ( .A(n2066), .B(n2067), .Z(n2064) );
  NANDN U2443 ( .A(B[137]), .B(n2068), .Z(n2067) );
  NANDN U2444 ( .A(A[137]), .B(n2069), .Z(n2068) );
  NANDN U2445 ( .A(n2069), .B(A[137]), .Z(n2066) );
  XOR U2446 ( .A(n2069), .B(n2070), .Z(DIFF[137]) );
  XOR U2447 ( .A(B[137]), .B(A[137]), .Z(n2070) );
  AND U2448 ( .A(n2071), .B(n2072), .Z(n2069) );
  NANDN U2449 ( .A(B[136]), .B(n2073), .Z(n2072) );
  NANDN U2450 ( .A(A[136]), .B(n2074), .Z(n2073) );
  NANDN U2451 ( .A(n2074), .B(A[136]), .Z(n2071) );
  XOR U2452 ( .A(n2074), .B(n2075), .Z(DIFF[136]) );
  XOR U2453 ( .A(B[136]), .B(A[136]), .Z(n2075) );
  AND U2454 ( .A(n2076), .B(n2077), .Z(n2074) );
  NANDN U2455 ( .A(B[135]), .B(n2078), .Z(n2077) );
  NANDN U2456 ( .A(A[135]), .B(n2079), .Z(n2078) );
  NANDN U2457 ( .A(n2079), .B(A[135]), .Z(n2076) );
  XOR U2458 ( .A(n2079), .B(n2080), .Z(DIFF[135]) );
  XOR U2459 ( .A(B[135]), .B(A[135]), .Z(n2080) );
  AND U2460 ( .A(n2081), .B(n2082), .Z(n2079) );
  NANDN U2461 ( .A(B[134]), .B(n2083), .Z(n2082) );
  NANDN U2462 ( .A(A[134]), .B(n2084), .Z(n2083) );
  NANDN U2463 ( .A(n2084), .B(A[134]), .Z(n2081) );
  XOR U2464 ( .A(n2084), .B(n2085), .Z(DIFF[134]) );
  XOR U2465 ( .A(B[134]), .B(A[134]), .Z(n2085) );
  AND U2466 ( .A(n2086), .B(n2087), .Z(n2084) );
  NANDN U2467 ( .A(B[133]), .B(n2088), .Z(n2087) );
  NANDN U2468 ( .A(A[133]), .B(n2089), .Z(n2088) );
  NANDN U2469 ( .A(n2089), .B(A[133]), .Z(n2086) );
  XOR U2470 ( .A(n2089), .B(n2090), .Z(DIFF[133]) );
  XOR U2471 ( .A(B[133]), .B(A[133]), .Z(n2090) );
  AND U2472 ( .A(n2091), .B(n2092), .Z(n2089) );
  NANDN U2473 ( .A(B[132]), .B(n2093), .Z(n2092) );
  NANDN U2474 ( .A(A[132]), .B(n2094), .Z(n2093) );
  NANDN U2475 ( .A(n2094), .B(A[132]), .Z(n2091) );
  XOR U2476 ( .A(n2094), .B(n2095), .Z(DIFF[132]) );
  XOR U2477 ( .A(B[132]), .B(A[132]), .Z(n2095) );
  AND U2478 ( .A(n2096), .B(n2097), .Z(n2094) );
  NANDN U2479 ( .A(B[131]), .B(n2098), .Z(n2097) );
  NANDN U2480 ( .A(A[131]), .B(n2099), .Z(n2098) );
  NANDN U2481 ( .A(n2099), .B(A[131]), .Z(n2096) );
  XOR U2482 ( .A(n2099), .B(n2100), .Z(DIFF[131]) );
  XOR U2483 ( .A(B[131]), .B(A[131]), .Z(n2100) );
  AND U2484 ( .A(n2101), .B(n2102), .Z(n2099) );
  NANDN U2485 ( .A(B[130]), .B(n2103), .Z(n2102) );
  NANDN U2486 ( .A(A[130]), .B(n2104), .Z(n2103) );
  NANDN U2487 ( .A(n2104), .B(A[130]), .Z(n2101) );
  XOR U2488 ( .A(n2104), .B(n2105), .Z(DIFF[130]) );
  XOR U2489 ( .A(B[130]), .B(A[130]), .Z(n2105) );
  AND U2490 ( .A(n2106), .B(n2107), .Z(n2104) );
  NANDN U2491 ( .A(B[129]), .B(n2108), .Z(n2107) );
  NANDN U2492 ( .A(A[129]), .B(n2109), .Z(n2108) );
  NANDN U2493 ( .A(n2109), .B(A[129]), .Z(n2106) );
  XOR U2494 ( .A(n2110), .B(n2111), .Z(DIFF[12]) );
  XOR U2495 ( .A(B[12]), .B(A[12]), .Z(n2111) );
  XOR U2496 ( .A(n2109), .B(n2112), .Z(DIFF[129]) );
  XOR U2497 ( .A(B[129]), .B(A[129]), .Z(n2112) );
  AND U2498 ( .A(n2113), .B(n2114), .Z(n2109) );
  NANDN U2499 ( .A(B[128]), .B(n2115), .Z(n2114) );
  NANDN U2500 ( .A(A[128]), .B(n2116), .Z(n2115) );
  NANDN U2501 ( .A(n2116), .B(A[128]), .Z(n2113) );
  XOR U2502 ( .A(n2116), .B(n2117), .Z(DIFF[128]) );
  XOR U2503 ( .A(B[128]), .B(A[128]), .Z(n2117) );
  AND U2504 ( .A(n2118), .B(n2119), .Z(n2116) );
  NANDN U2505 ( .A(B[127]), .B(n2120), .Z(n2119) );
  NANDN U2506 ( .A(A[127]), .B(n2121), .Z(n2120) );
  NANDN U2507 ( .A(n2121), .B(A[127]), .Z(n2118) );
  XOR U2508 ( .A(n2121), .B(n2122), .Z(DIFF[127]) );
  XOR U2509 ( .A(B[127]), .B(A[127]), .Z(n2122) );
  AND U2510 ( .A(n2123), .B(n2124), .Z(n2121) );
  NANDN U2511 ( .A(B[126]), .B(n2125), .Z(n2124) );
  NANDN U2512 ( .A(A[126]), .B(n2126), .Z(n2125) );
  NANDN U2513 ( .A(n2126), .B(A[126]), .Z(n2123) );
  XOR U2514 ( .A(n2126), .B(n2127), .Z(DIFF[126]) );
  XOR U2515 ( .A(B[126]), .B(A[126]), .Z(n2127) );
  AND U2516 ( .A(n2128), .B(n2129), .Z(n2126) );
  NANDN U2517 ( .A(B[125]), .B(n2130), .Z(n2129) );
  NANDN U2518 ( .A(A[125]), .B(n2131), .Z(n2130) );
  NANDN U2519 ( .A(n2131), .B(A[125]), .Z(n2128) );
  XOR U2520 ( .A(n2131), .B(n2132), .Z(DIFF[125]) );
  XOR U2521 ( .A(B[125]), .B(A[125]), .Z(n2132) );
  AND U2522 ( .A(n2133), .B(n2134), .Z(n2131) );
  NANDN U2523 ( .A(B[124]), .B(n2135), .Z(n2134) );
  NANDN U2524 ( .A(A[124]), .B(n2136), .Z(n2135) );
  NANDN U2525 ( .A(n2136), .B(A[124]), .Z(n2133) );
  XOR U2526 ( .A(n2136), .B(n2137), .Z(DIFF[124]) );
  XOR U2527 ( .A(B[124]), .B(A[124]), .Z(n2137) );
  AND U2528 ( .A(n2138), .B(n2139), .Z(n2136) );
  NANDN U2529 ( .A(B[123]), .B(n2140), .Z(n2139) );
  NANDN U2530 ( .A(A[123]), .B(n2141), .Z(n2140) );
  NANDN U2531 ( .A(n2141), .B(A[123]), .Z(n2138) );
  XOR U2532 ( .A(n2141), .B(n2142), .Z(DIFF[123]) );
  XOR U2533 ( .A(B[123]), .B(A[123]), .Z(n2142) );
  AND U2534 ( .A(n2143), .B(n2144), .Z(n2141) );
  NANDN U2535 ( .A(B[122]), .B(n2145), .Z(n2144) );
  NANDN U2536 ( .A(A[122]), .B(n2146), .Z(n2145) );
  NANDN U2537 ( .A(n2146), .B(A[122]), .Z(n2143) );
  XOR U2538 ( .A(n2146), .B(n2147), .Z(DIFF[122]) );
  XOR U2539 ( .A(B[122]), .B(A[122]), .Z(n2147) );
  AND U2540 ( .A(n2148), .B(n2149), .Z(n2146) );
  NANDN U2541 ( .A(B[121]), .B(n2150), .Z(n2149) );
  NANDN U2542 ( .A(A[121]), .B(n2151), .Z(n2150) );
  NANDN U2543 ( .A(n2151), .B(A[121]), .Z(n2148) );
  XOR U2544 ( .A(n2151), .B(n2152), .Z(DIFF[121]) );
  XOR U2545 ( .A(B[121]), .B(A[121]), .Z(n2152) );
  AND U2546 ( .A(n2153), .B(n2154), .Z(n2151) );
  NANDN U2547 ( .A(B[120]), .B(n2155), .Z(n2154) );
  NANDN U2548 ( .A(A[120]), .B(n2156), .Z(n2155) );
  NANDN U2549 ( .A(n2156), .B(A[120]), .Z(n2153) );
  XOR U2550 ( .A(n2156), .B(n2157), .Z(DIFF[120]) );
  XOR U2551 ( .A(B[120]), .B(A[120]), .Z(n2157) );
  AND U2552 ( .A(n2158), .B(n2159), .Z(n2156) );
  NANDN U2553 ( .A(B[119]), .B(n2160), .Z(n2159) );
  NANDN U2554 ( .A(A[119]), .B(n2161), .Z(n2160) );
  NANDN U2555 ( .A(n2161), .B(A[119]), .Z(n2158) );
  XOR U2556 ( .A(n2162), .B(n2163), .Z(DIFF[11]) );
  XOR U2557 ( .A(B[11]), .B(A[11]), .Z(n2163) );
  XOR U2558 ( .A(n2161), .B(n2164), .Z(DIFF[119]) );
  XOR U2559 ( .A(B[119]), .B(A[119]), .Z(n2164) );
  AND U2560 ( .A(n2165), .B(n2166), .Z(n2161) );
  NANDN U2561 ( .A(B[118]), .B(n2167), .Z(n2166) );
  NANDN U2562 ( .A(A[118]), .B(n2168), .Z(n2167) );
  NANDN U2563 ( .A(n2168), .B(A[118]), .Z(n2165) );
  XOR U2564 ( .A(n2168), .B(n2169), .Z(DIFF[118]) );
  XOR U2565 ( .A(B[118]), .B(A[118]), .Z(n2169) );
  AND U2566 ( .A(n2170), .B(n2171), .Z(n2168) );
  NANDN U2567 ( .A(B[117]), .B(n2172), .Z(n2171) );
  NANDN U2568 ( .A(A[117]), .B(n2173), .Z(n2172) );
  NANDN U2569 ( .A(n2173), .B(A[117]), .Z(n2170) );
  XOR U2570 ( .A(n2173), .B(n2174), .Z(DIFF[117]) );
  XOR U2571 ( .A(B[117]), .B(A[117]), .Z(n2174) );
  AND U2572 ( .A(n2175), .B(n2176), .Z(n2173) );
  NANDN U2573 ( .A(B[116]), .B(n2177), .Z(n2176) );
  NANDN U2574 ( .A(A[116]), .B(n2178), .Z(n2177) );
  NANDN U2575 ( .A(n2178), .B(A[116]), .Z(n2175) );
  XOR U2576 ( .A(n2178), .B(n2179), .Z(DIFF[116]) );
  XOR U2577 ( .A(B[116]), .B(A[116]), .Z(n2179) );
  AND U2578 ( .A(n2180), .B(n2181), .Z(n2178) );
  NANDN U2579 ( .A(B[115]), .B(n2182), .Z(n2181) );
  NANDN U2580 ( .A(A[115]), .B(n2183), .Z(n2182) );
  NANDN U2581 ( .A(n2183), .B(A[115]), .Z(n2180) );
  XOR U2582 ( .A(n2183), .B(n2184), .Z(DIFF[115]) );
  XOR U2583 ( .A(B[115]), .B(A[115]), .Z(n2184) );
  AND U2584 ( .A(n2185), .B(n2186), .Z(n2183) );
  NANDN U2585 ( .A(B[114]), .B(n2187), .Z(n2186) );
  NANDN U2586 ( .A(A[114]), .B(n2188), .Z(n2187) );
  NANDN U2587 ( .A(n2188), .B(A[114]), .Z(n2185) );
  XOR U2588 ( .A(n2188), .B(n2189), .Z(DIFF[114]) );
  XOR U2589 ( .A(B[114]), .B(A[114]), .Z(n2189) );
  AND U2590 ( .A(n2190), .B(n2191), .Z(n2188) );
  NANDN U2591 ( .A(B[113]), .B(n2192), .Z(n2191) );
  NANDN U2592 ( .A(A[113]), .B(n2193), .Z(n2192) );
  NANDN U2593 ( .A(n2193), .B(A[113]), .Z(n2190) );
  XOR U2594 ( .A(n2193), .B(n2194), .Z(DIFF[113]) );
  XOR U2595 ( .A(B[113]), .B(A[113]), .Z(n2194) );
  AND U2596 ( .A(n2195), .B(n2196), .Z(n2193) );
  NANDN U2597 ( .A(B[112]), .B(n2197), .Z(n2196) );
  NANDN U2598 ( .A(A[112]), .B(n2198), .Z(n2197) );
  NANDN U2599 ( .A(n2198), .B(A[112]), .Z(n2195) );
  XOR U2600 ( .A(n2198), .B(n2199), .Z(DIFF[112]) );
  XOR U2601 ( .A(B[112]), .B(A[112]), .Z(n2199) );
  AND U2602 ( .A(n2200), .B(n2201), .Z(n2198) );
  NANDN U2603 ( .A(B[111]), .B(n2202), .Z(n2201) );
  NANDN U2604 ( .A(A[111]), .B(n2203), .Z(n2202) );
  NANDN U2605 ( .A(n2203), .B(A[111]), .Z(n2200) );
  XOR U2606 ( .A(n2203), .B(n2204), .Z(DIFF[111]) );
  XOR U2607 ( .A(B[111]), .B(A[111]), .Z(n2204) );
  AND U2608 ( .A(n2205), .B(n2206), .Z(n2203) );
  NANDN U2609 ( .A(B[110]), .B(n2207), .Z(n2206) );
  NANDN U2610 ( .A(A[110]), .B(n2208), .Z(n2207) );
  NANDN U2611 ( .A(n2208), .B(A[110]), .Z(n2205) );
  XOR U2612 ( .A(n2208), .B(n2209), .Z(DIFF[110]) );
  XOR U2613 ( .A(B[110]), .B(A[110]), .Z(n2209) );
  AND U2614 ( .A(n2210), .B(n2211), .Z(n2208) );
  NANDN U2615 ( .A(B[109]), .B(n2212), .Z(n2211) );
  NANDN U2616 ( .A(A[109]), .B(n2213), .Z(n2212) );
  NANDN U2617 ( .A(n2213), .B(A[109]), .Z(n2210) );
  XOR U2618 ( .A(n2214), .B(n2215), .Z(DIFF[10]) );
  XOR U2619 ( .A(B[10]), .B(A[10]), .Z(n2215) );
  XOR U2620 ( .A(n2213), .B(n2216), .Z(DIFF[109]) );
  XOR U2621 ( .A(B[109]), .B(A[109]), .Z(n2216) );
  AND U2622 ( .A(n2217), .B(n2218), .Z(n2213) );
  NANDN U2623 ( .A(B[108]), .B(n2219), .Z(n2218) );
  NANDN U2624 ( .A(A[108]), .B(n2220), .Z(n2219) );
  NANDN U2625 ( .A(n2220), .B(A[108]), .Z(n2217) );
  XOR U2626 ( .A(n2220), .B(n2221), .Z(DIFF[108]) );
  XOR U2627 ( .A(B[108]), .B(A[108]), .Z(n2221) );
  AND U2628 ( .A(n2222), .B(n2223), .Z(n2220) );
  NANDN U2629 ( .A(B[107]), .B(n2224), .Z(n2223) );
  NANDN U2630 ( .A(A[107]), .B(n2225), .Z(n2224) );
  NANDN U2631 ( .A(n2225), .B(A[107]), .Z(n2222) );
  XOR U2632 ( .A(n2225), .B(n2226), .Z(DIFF[107]) );
  XOR U2633 ( .A(B[107]), .B(A[107]), .Z(n2226) );
  AND U2634 ( .A(n2227), .B(n2228), .Z(n2225) );
  NANDN U2635 ( .A(B[106]), .B(n2229), .Z(n2228) );
  NANDN U2636 ( .A(A[106]), .B(n2230), .Z(n2229) );
  NANDN U2637 ( .A(n2230), .B(A[106]), .Z(n2227) );
  XOR U2638 ( .A(n2230), .B(n2231), .Z(DIFF[106]) );
  XOR U2639 ( .A(B[106]), .B(A[106]), .Z(n2231) );
  AND U2640 ( .A(n2232), .B(n2233), .Z(n2230) );
  NANDN U2641 ( .A(B[105]), .B(n2234), .Z(n2233) );
  NANDN U2642 ( .A(A[105]), .B(n2235), .Z(n2234) );
  NANDN U2643 ( .A(n2235), .B(A[105]), .Z(n2232) );
  XOR U2644 ( .A(n2235), .B(n2236), .Z(DIFF[105]) );
  XOR U2645 ( .A(B[105]), .B(A[105]), .Z(n2236) );
  AND U2646 ( .A(n2237), .B(n2238), .Z(n2235) );
  NANDN U2647 ( .A(B[104]), .B(n2239), .Z(n2238) );
  NANDN U2648 ( .A(A[104]), .B(n2240), .Z(n2239) );
  NANDN U2649 ( .A(n2240), .B(A[104]), .Z(n2237) );
  XOR U2650 ( .A(n2240), .B(n2241), .Z(DIFF[104]) );
  XOR U2651 ( .A(B[104]), .B(A[104]), .Z(n2241) );
  AND U2652 ( .A(n2242), .B(n2243), .Z(n2240) );
  NANDN U2653 ( .A(B[103]), .B(n2244), .Z(n2243) );
  NANDN U2654 ( .A(A[103]), .B(n2245), .Z(n2244) );
  NANDN U2655 ( .A(n2245), .B(A[103]), .Z(n2242) );
  XOR U2656 ( .A(n2245), .B(n2246), .Z(DIFF[103]) );
  XOR U2657 ( .A(B[103]), .B(A[103]), .Z(n2246) );
  AND U2658 ( .A(n2247), .B(n2248), .Z(n2245) );
  NANDN U2659 ( .A(B[102]), .B(n2249), .Z(n2248) );
  NANDN U2660 ( .A(A[102]), .B(n2250), .Z(n2249) );
  NANDN U2661 ( .A(n2250), .B(A[102]), .Z(n2247) );
  XOR U2662 ( .A(n2250), .B(n2251), .Z(DIFF[102]) );
  XOR U2663 ( .A(B[102]), .B(A[102]), .Z(n2251) );
  AND U2664 ( .A(n2252), .B(n2253), .Z(n2250) );
  NANDN U2665 ( .A(B[101]), .B(n2254), .Z(n2253) );
  NANDN U2666 ( .A(A[101]), .B(n2255), .Z(n2254) );
  NANDN U2667 ( .A(n2255), .B(A[101]), .Z(n2252) );
  XOR U2668 ( .A(n2255), .B(n2256), .Z(DIFF[101]) );
  XOR U2669 ( .A(B[101]), .B(A[101]), .Z(n2256) );
  AND U2670 ( .A(n2257), .B(n2258), .Z(n2255) );
  NANDN U2671 ( .A(B[100]), .B(n2259), .Z(n2258) );
  NANDN U2672 ( .A(A[100]), .B(n2260), .Z(n2259) );
  NANDN U2673 ( .A(n2260), .B(A[100]), .Z(n2257) );
  XOR U2674 ( .A(n2260), .B(n2261), .Z(DIFF[100]) );
  XOR U2675 ( .A(B[100]), .B(A[100]), .Z(n2261) );
  AND U2676 ( .A(n2262), .B(n2263), .Z(n2260) );
  NANDN U2677 ( .A(B[99]), .B(n2264), .Z(n2263) );
  OR U2678 ( .A(n5), .B(A[99]), .Z(n2264) );
  NAND U2679 ( .A(A[99]), .B(n5), .Z(n2262) );
  NAND U2680 ( .A(n2265), .B(n2266), .Z(n5) );
  NANDN U2681 ( .A(B[98]), .B(n2267), .Z(n2266) );
  NANDN U2682 ( .A(A[98]), .B(n7), .Z(n2267) );
  NANDN U2683 ( .A(n7), .B(A[98]), .Z(n2265) );
  AND U2684 ( .A(n2268), .B(n2269), .Z(n7) );
  NANDN U2685 ( .A(B[97]), .B(n2270), .Z(n2269) );
  NANDN U2686 ( .A(A[97]), .B(n9), .Z(n2270) );
  NANDN U2687 ( .A(n9), .B(A[97]), .Z(n2268) );
  AND U2688 ( .A(n2271), .B(n2272), .Z(n9) );
  NANDN U2689 ( .A(B[96]), .B(n2273), .Z(n2272) );
  NANDN U2690 ( .A(A[96]), .B(n11), .Z(n2273) );
  NANDN U2691 ( .A(n11), .B(A[96]), .Z(n2271) );
  AND U2692 ( .A(n2274), .B(n2275), .Z(n11) );
  NANDN U2693 ( .A(B[95]), .B(n2276), .Z(n2275) );
  NANDN U2694 ( .A(A[95]), .B(n13), .Z(n2276) );
  NANDN U2695 ( .A(n13), .B(A[95]), .Z(n2274) );
  AND U2696 ( .A(n2277), .B(n2278), .Z(n13) );
  NANDN U2697 ( .A(B[94]), .B(n2279), .Z(n2278) );
  NANDN U2698 ( .A(A[94]), .B(n15), .Z(n2279) );
  NANDN U2699 ( .A(n15), .B(A[94]), .Z(n2277) );
  AND U2700 ( .A(n2280), .B(n2281), .Z(n15) );
  NANDN U2701 ( .A(B[93]), .B(n2282), .Z(n2281) );
  NANDN U2702 ( .A(A[93]), .B(n17), .Z(n2282) );
  NANDN U2703 ( .A(n17), .B(A[93]), .Z(n2280) );
  AND U2704 ( .A(n2283), .B(n2284), .Z(n17) );
  NANDN U2705 ( .A(B[92]), .B(n2285), .Z(n2284) );
  NANDN U2706 ( .A(A[92]), .B(n19), .Z(n2285) );
  NANDN U2707 ( .A(n19), .B(A[92]), .Z(n2283) );
  AND U2708 ( .A(n2286), .B(n2287), .Z(n19) );
  NANDN U2709 ( .A(B[91]), .B(n2288), .Z(n2287) );
  NANDN U2710 ( .A(A[91]), .B(n21), .Z(n2288) );
  NANDN U2711 ( .A(n21), .B(A[91]), .Z(n2286) );
  AND U2712 ( .A(n2289), .B(n2290), .Z(n21) );
  NANDN U2713 ( .A(B[90]), .B(n2291), .Z(n2290) );
  NANDN U2714 ( .A(A[90]), .B(n23), .Z(n2291) );
  NANDN U2715 ( .A(n23), .B(A[90]), .Z(n2289) );
  AND U2716 ( .A(n2292), .B(n2293), .Z(n23) );
  NANDN U2717 ( .A(B[89]), .B(n2294), .Z(n2293) );
  NANDN U2718 ( .A(A[89]), .B(n27), .Z(n2294) );
  NANDN U2719 ( .A(n27), .B(A[89]), .Z(n2292) );
  AND U2720 ( .A(n2295), .B(n2296), .Z(n27) );
  NANDN U2721 ( .A(B[88]), .B(n2297), .Z(n2296) );
  NANDN U2722 ( .A(A[88]), .B(n29), .Z(n2297) );
  NANDN U2723 ( .A(n29), .B(A[88]), .Z(n2295) );
  AND U2724 ( .A(n2298), .B(n2299), .Z(n29) );
  NANDN U2725 ( .A(B[87]), .B(n2300), .Z(n2299) );
  NANDN U2726 ( .A(A[87]), .B(n31), .Z(n2300) );
  NANDN U2727 ( .A(n31), .B(A[87]), .Z(n2298) );
  AND U2728 ( .A(n2301), .B(n2302), .Z(n31) );
  NANDN U2729 ( .A(B[86]), .B(n2303), .Z(n2302) );
  NANDN U2730 ( .A(A[86]), .B(n33), .Z(n2303) );
  NANDN U2731 ( .A(n33), .B(A[86]), .Z(n2301) );
  AND U2732 ( .A(n2304), .B(n2305), .Z(n33) );
  NANDN U2733 ( .A(B[85]), .B(n2306), .Z(n2305) );
  NANDN U2734 ( .A(A[85]), .B(n35), .Z(n2306) );
  NANDN U2735 ( .A(n35), .B(A[85]), .Z(n2304) );
  AND U2736 ( .A(n2307), .B(n2308), .Z(n35) );
  NANDN U2737 ( .A(B[84]), .B(n2309), .Z(n2308) );
  NANDN U2738 ( .A(A[84]), .B(n37), .Z(n2309) );
  NANDN U2739 ( .A(n37), .B(A[84]), .Z(n2307) );
  AND U2740 ( .A(n2310), .B(n2311), .Z(n37) );
  NANDN U2741 ( .A(B[83]), .B(n2312), .Z(n2311) );
  NANDN U2742 ( .A(A[83]), .B(n39), .Z(n2312) );
  NANDN U2743 ( .A(n39), .B(A[83]), .Z(n2310) );
  AND U2744 ( .A(n2313), .B(n2314), .Z(n39) );
  NANDN U2745 ( .A(B[82]), .B(n2315), .Z(n2314) );
  NANDN U2746 ( .A(A[82]), .B(n41), .Z(n2315) );
  NANDN U2747 ( .A(n41), .B(A[82]), .Z(n2313) );
  AND U2748 ( .A(n2316), .B(n2317), .Z(n41) );
  NANDN U2749 ( .A(B[81]), .B(n2318), .Z(n2317) );
  NANDN U2750 ( .A(A[81]), .B(n43), .Z(n2318) );
  NANDN U2751 ( .A(n43), .B(A[81]), .Z(n2316) );
  AND U2752 ( .A(n2319), .B(n2320), .Z(n43) );
  NANDN U2753 ( .A(B[80]), .B(n2321), .Z(n2320) );
  NANDN U2754 ( .A(A[80]), .B(n45), .Z(n2321) );
  NANDN U2755 ( .A(n45), .B(A[80]), .Z(n2319) );
  AND U2756 ( .A(n2322), .B(n2323), .Z(n45) );
  NANDN U2757 ( .A(B[79]), .B(n2324), .Z(n2323) );
  NANDN U2758 ( .A(A[79]), .B(n49), .Z(n2324) );
  NANDN U2759 ( .A(n49), .B(A[79]), .Z(n2322) );
  AND U2760 ( .A(n2325), .B(n2326), .Z(n49) );
  NANDN U2761 ( .A(B[78]), .B(n2327), .Z(n2326) );
  NANDN U2762 ( .A(A[78]), .B(n51), .Z(n2327) );
  NANDN U2763 ( .A(n51), .B(A[78]), .Z(n2325) );
  AND U2764 ( .A(n2328), .B(n2329), .Z(n51) );
  NANDN U2765 ( .A(B[77]), .B(n2330), .Z(n2329) );
  NANDN U2766 ( .A(A[77]), .B(n53), .Z(n2330) );
  NANDN U2767 ( .A(n53), .B(A[77]), .Z(n2328) );
  AND U2768 ( .A(n2331), .B(n2332), .Z(n53) );
  NANDN U2769 ( .A(B[76]), .B(n2333), .Z(n2332) );
  NANDN U2770 ( .A(A[76]), .B(n55), .Z(n2333) );
  NANDN U2771 ( .A(n55), .B(A[76]), .Z(n2331) );
  AND U2772 ( .A(n2334), .B(n2335), .Z(n55) );
  NANDN U2773 ( .A(B[75]), .B(n2336), .Z(n2335) );
  NANDN U2774 ( .A(A[75]), .B(n57), .Z(n2336) );
  NANDN U2775 ( .A(n57), .B(A[75]), .Z(n2334) );
  AND U2776 ( .A(n2337), .B(n2338), .Z(n57) );
  NANDN U2777 ( .A(B[74]), .B(n2339), .Z(n2338) );
  NANDN U2778 ( .A(A[74]), .B(n59), .Z(n2339) );
  NANDN U2779 ( .A(n59), .B(A[74]), .Z(n2337) );
  AND U2780 ( .A(n2340), .B(n2341), .Z(n59) );
  NANDN U2781 ( .A(B[73]), .B(n2342), .Z(n2341) );
  NANDN U2782 ( .A(A[73]), .B(n61), .Z(n2342) );
  NANDN U2783 ( .A(n61), .B(A[73]), .Z(n2340) );
  AND U2784 ( .A(n2343), .B(n2344), .Z(n61) );
  NANDN U2785 ( .A(B[72]), .B(n2345), .Z(n2344) );
  NANDN U2786 ( .A(A[72]), .B(n63), .Z(n2345) );
  NANDN U2787 ( .A(n63), .B(A[72]), .Z(n2343) );
  AND U2788 ( .A(n2346), .B(n2347), .Z(n63) );
  NANDN U2789 ( .A(B[71]), .B(n2348), .Z(n2347) );
  NANDN U2790 ( .A(A[71]), .B(n65), .Z(n2348) );
  NANDN U2791 ( .A(n65), .B(A[71]), .Z(n2346) );
  AND U2792 ( .A(n2349), .B(n2350), .Z(n65) );
  NANDN U2793 ( .A(B[70]), .B(n2351), .Z(n2350) );
  NANDN U2794 ( .A(A[70]), .B(n67), .Z(n2351) );
  NANDN U2795 ( .A(n67), .B(A[70]), .Z(n2349) );
  AND U2796 ( .A(n2352), .B(n2353), .Z(n67) );
  NANDN U2797 ( .A(B[69]), .B(n2354), .Z(n2353) );
  NANDN U2798 ( .A(A[69]), .B(n71), .Z(n2354) );
  NANDN U2799 ( .A(n71), .B(A[69]), .Z(n2352) );
  AND U2800 ( .A(n2355), .B(n2356), .Z(n71) );
  NANDN U2801 ( .A(B[68]), .B(n2357), .Z(n2356) );
  NANDN U2802 ( .A(A[68]), .B(n73), .Z(n2357) );
  NANDN U2803 ( .A(n73), .B(A[68]), .Z(n2355) );
  AND U2804 ( .A(n2358), .B(n2359), .Z(n73) );
  NANDN U2805 ( .A(B[67]), .B(n2360), .Z(n2359) );
  NANDN U2806 ( .A(A[67]), .B(n75), .Z(n2360) );
  NANDN U2807 ( .A(n75), .B(A[67]), .Z(n2358) );
  AND U2808 ( .A(n2361), .B(n2362), .Z(n75) );
  NANDN U2809 ( .A(B[66]), .B(n2363), .Z(n2362) );
  NANDN U2810 ( .A(A[66]), .B(n77), .Z(n2363) );
  NANDN U2811 ( .A(n77), .B(A[66]), .Z(n2361) );
  AND U2812 ( .A(n2364), .B(n2365), .Z(n77) );
  NANDN U2813 ( .A(B[65]), .B(n2366), .Z(n2365) );
  NANDN U2814 ( .A(A[65]), .B(n79), .Z(n2366) );
  NANDN U2815 ( .A(n79), .B(A[65]), .Z(n2364) );
  AND U2816 ( .A(n2367), .B(n2368), .Z(n79) );
  NANDN U2817 ( .A(B[64]), .B(n2369), .Z(n2368) );
  NANDN U2818 ( .A(A[64]), .B(n81), .Z(n2369) );
  NANDN U2819 ( .A(n81), .B(A[64]), .Z(n2367) );
  AND U2820 ( .A(n2370), .B(n2371), .Z(n81) );
  NANDN U2821 ( .A(B[63]), .B(n2372), .Z(n2371) );
  NANDN U2822 ( .A(A[63]), .B(n83), .Z(n2372) );
  NANDN U2823 ( .A(n83), .B(A[63]), .Z(n2370) );
  AND U2824 ( .A(n2373), .B(n2374), .Z(n83) );
  NANDN U2825 ( .A(B[62]), .B(n2375), .Z(n2374) );
  NANDN U2826 ( .A(A[62]), .B(n85), .Z(n2375) );
  NANDN U2827 ( .A(n85), .B(A[62]), .Z(n2373) );
  AND U2828 ( .A(n2376), .B(n2377), .Z(n85) );
  NANDN U2829 ( .A(B[61]), .B(n2378), .Z(n2377) );
  NANDN U2830 ( .A(A[61]), .B(n87), .Z(n2378) );
  NANDN U2831 ( .A(n87), .B(A[61]), .Z(n2376) );
  AND U2832 ( .A(n2379), .B(n2380), .Z(n87) );
  NANDN U2833 ( .A(B[60]), .B(n2381), .Z(n2380) );
  NANDN U2834 ( .A(A[60]), .B(n89), .Z(n2381) );
  NANDN U2835 ( .A(n89), .B(A[60]), .Z(n2379) );
  AND U2836 ( .A(n2382), .B(n2383), .Z(n89) );
  NANDN U2837 ( .A(B[59]), .B(n2384), .Z(n2383) );
  NANDN U2838 ( .A(A[59]), .B(n93), .Z(n2384) );
  NANDN U2839 ( .A(n93), .B(A[59]), .Z(n2382) );
  AND U2840 ( .A(n2385), .B(n2386), .Z(n93) );
  NANDN U2841 ( .A(B[58]), .B(n2387), .Z(n2386) );
  NANDN U2842 ( .A(A[58]), .B(n95), .Z(n2387) );
  NANDN U2843 ( .A(n95), .B(A[58]), .Z(n2385) );
  AND U2844 ( .A(n2388), .B(n2389), .Z(n95) );
  NANDN U2845 ( .A(B[57]), .B(n2390), .Z(n2389) );
  NANDN U2846 ( .A(A[57]), .B(n97), .Z(n2390) );
  NANDN U2847 ( .A(n97), .B(A[57]), .Z(n2388) );
  AND U2848 ( .A(n2391), .B(n2392), .Z(n97) );
  NANDN U2849 ( .A(B[56]), .B(n2393), .Z(n2392) );
  NANDN U2850 ( .A(A[56]), .B(n99), .Z(n2393) );
  NANDN U2851 ( .A(n99), .B(A[56]), .Z(n2391) );
  AND U2852 ( .A(n2394), .B(n2395), .Z(n99) );
  NANDN U2853 ( .A(B[55]), .B(n2396), .Z(n2395) );
  NANDN U2854 ( .A(A[55]), .B(n101), .Z(n2396) );
  NANDN U2855 ( .A(n101), .B(A[55]), .Z(n2394) );
  AND U2856 ( .A(n2397), .B(n2398), .Z(n101) );
  NANDN U2857 ( .A(B[54]), .B(n2399), .Z(n2398) );
  NANDN U2858 ( .A(A[54]), .B(n103), .Z(n2399) );
  NANDN U2859 ( .A(n103), .B(A[54]), .Z(n2397) );
  AND U2860 ( .A(n2400), .B(n2401), .Z(n103) );
  NANDN U2861 ( .A(B[53]), .B(n2402), .Z(n2401) );
  NANDN U2862 ( .A(A[53]), .B(n105), .Z(n2402) );
  NANDN U2863 ( .A(n105), .B(A[53]), .Z(n2400) );
  AND U2864 ( .A(n2403), .B(n2404), .Z(n105) );
  NANDN U2865 ( .A(B[52]), .B(n2405), .Z(n2404) );
  NANDN U2866 ( .A(A[52]), .B(n107), .Z(n2405) );
  NANDN U2867 ( .A(n107), .B(A[52]), .Z(n2403) );
  AND U2868 ( .A(n2406), .B(n2407), .Z(n107) );
  NANDN U2869 ( .A(B[51]), .B(n2408), .Z(n2407) );
  NANDN U2870 ( .A(A[51]), .B(n109), .Z(n2408) );
  NANDN U2871 ( .A(n109), .B(A[51]), .Z(n2406) );
  AND U2872 ( .A(n2409), .B(n2410), .Z(n109) );
  NANDN U2873 ( .A(B[50]), .B(n2411), .Z(n2410) );
  NANDN U2874 ( .A(A[50]), .B(n127), .Z(n2411) );
  NANDN U2875 ( .A(n127), .B(A[50]), .Z(n2409) );
  AND U2876 ( .A(n2412), .B(n2413), .Z(n127) );
  NANDN U2877 ( .A(B[49]), .B(n2414), .Z(n2413) );
  NANDN U2878 ( .A(A[49]), .B(n181), .Z(n2414) );
  NANDN U2879 ( .A(n181), .B(A[49]), .Z(n2412) );
  AND U2880 ( .A(n2415), .B(n2416), .Z(n181) );
  NANDN U2881 ( .A(B[48]), .B(n2417), .Z(n2416) );
  NANDN U2882 ( .A(A[48]), .B(n233), .Z(n2417) );
  NANDN U2883 ( .A(n233), .B(A[48]), .Z(n2415) );
  AND U2884 ( .A(n2418), .B(n2419), .Z(n233) );
  NANDN U2885 ( .A(B[47]), .B(n2420), .Z(n2419) );
  NANDN U2886 ( .A(A[47]), .B(n285), .Z(n2420) );
  NANDN U2887 ( .A(n285), .B(A[47]), .Z(n2418) );
  AND U2888 ( .A(n2421), .B(n2422), .Z(n285) );
  NANDN U2889 ( .A(B[46]), .B(n2423), .Z(n2422) );
  NANDN U2890 ( .A(A[46]), .B(n337), .Z(n2423) );
  NANDN U2891 ( .A(n337), .B(A[46]), .Z(n2421) );
  AND U2892 ( .A(n2424), .B(n2425), .Z(n337) );
  NANDN U2893 ( .A(B[45]), .B(n2426), .Z(n2425) );
  NANDN U2894 ( .A(A[45]), .B(n389), .Z(n2426) );
  NANDN U2895 ( .A(n389), .B(A[45]), .Z(n2424) );
  AND U2896 ( .A(n2427), .B(n2428), .Z(n389) );
  NANDN U2897 ( .A(B[44]), .B(n2429), .Z(n2428) );
  NANDN U2898 ( .A(A[44]), .B(n441), .Z(n2429) );
  NANDN U2899 ( .A(n441), .B(A[44]), .Z(n2427) );
  AND U2900 ( .A(n2430), .B(n2431), .Z(n441) );
  NANDN U2901 ( .A(B[43]), .B(n2432), .Z(n2431) );
  NANDN U2902 ( .A(A[43]), .B(n493), .Z(n2432) );
  NANDN U2903 ( .A(n493), .B(A[43]), .Z(n2430) );
  AND U2904 ( .A(n2433), .B(n2434), .Z(n493) );
  NANDN U2905 ( .A(B[42]), .B(n2435), .Z(n2434) );
  NANDN U2906 ( .A(A[42]), .B(n545), .Z(n2435) );
  NANDN U2907 ( .A(n545), .B(A[42]), .Z(n2433) );
  AND U2908 ( .A(n2436), .B(n2437), .Z(n545) );
  NANDN U2909 ( .A(B[41]), .B(n2438), .Z(n2437) );
  NANDN U2910 ( .A(A[41]), .B(n597), .Z(n2438) );
  NANDN U2911 ( .A(n597), .B(A[41]), .Z(n2436) );
  AND U2912 ( .A(n2439), .B(n2440), .Z(n597) );
  NANDN U2913 ( .A(B[40]), .B(n2441), .Z(n2440) );
  NANDN U2914 ( .A(A[40]), .B(n649), .Z(n2441) );
  NANDN U2915 ( .A(n649), .B(A[40]), .Z(n2439) );
  AND U2916 ( .A(n2442), .B(n2443), .Z(n649) );
  NANDN U2917 ( .A(B[39]), .B(n2444), .Z(n2443) );
  NANDN U2918 ( .A(A[39]), .B(n703), .Z(n2444) );
  NANDN U2919 ( .A(n703), .B(A[39]), .Z(n2442) );
  AND U2920 ( .A(n2445), .B(n2446), .Z(n703) );
  NANDN U2921 ( .A(B[38]), .B(n2447), .Z(n2446) );
  NANDN U2922 ( .A(A[38]), .B(n755), .Z(n2447) );
  NANDN U2923 ( .A(n755), .B(A[38]), .Z(n2445) );
  AND U2924 ( .A(n2448), .B(n2449), .Z(n755) );
  NANDN U2925 ( .A(B[37]), .B(n2450), .Z(n2449) );
  NANDN U2926 ( .A(A[37]), .B(n807), .Z(n2450) );
  NANDN U2927 ( .A(n807), .B(A[37]), .Z(n2448) );
  AND U2928 ( .A(n2451), .B(n2452), .Z(n807) );
  NANDN U2929 ( .A(B[36]), .B(n2453), .Z(n2452) );
  NANDN U2930 ( .A(A[36]), .B(n859), .Z(n2453) );
  NANDN U2931 ( .A(n859), .B(A[36]), .Z(n2451) );
  AND U2932 ( .A(n2454), .B(n2455), .Z(n859) );
  NANDN U2933 ( .A(B[35]), .B(n2456), .Z(n2455) );
  NANDN U2934 ( .A(A[35]), .B(n911), .Z(n2456) );
  NANDN U2935 ( .A(n911), .B(A[35]), .Z(n2454) );
  AND U2936 ( .A(n2457), .B(n2458), .Z(n911) );
  NANDN U2937 ( .A(B[34]), .B(n2459), .Z(n2458) );
  NANDN U2938 ( .A(A[34]), .B(n963), .Z(n2459) );
  NANDN U2939 ( .A(n963), .B(A[34]), .Z(n2457) );
  AND U2940 ( .A(n2460), .B(n2461), .Z(n963) );
  NANDN U2941 ( .A(B[33]), .B(n2462), .Z(n2461) );
  NANDN U2942 ( .A(A[33]), .B(n1015), .Z(n2462) );
  NANDN U2943 ( .A(n1015), .B(A[33]), .Z(n2460) );
  AND U2944 ( .A(n2463), .B(n2464), .Z(n1015) );
  NANDN U2945 ( .A(B[32]), .B(n2465), .Z(n2464) );
  NANDN U2946 ( .A(A[32]), .B(n1067), .Z(n2465) );
  NANDN U2947 ( .A(n1067), .B(A[32]), .Z(n2463) );
  AND U2948 ( .A(n2466), .B(n2467), .Z(n1067) );
  NANDN U2949 ( .A(B[31]), .B(n2468), .Z(n2467) );
  NANDN U2950 ( .A(A[31]), .B(n1119), .Z(n2468) );
  NANDN U2951 ( .A(n1119), .B(A[31]), .Z(n2466) );
  AND U2952 ( .A(n2469), .B(n2470), .Z(n1119) );
  NANDN U2953 ( .A(B[30]), .B(n2471), .Z(n2470) );
  NANDN U2954 ( .A(A[30]), .B(n1171), .Z(n2471) );
  NANDN U2955 ( .A(n1171), .B(A[30]), .Z(n2469) );
  AND U2956 ( .A(n2472), .B(n2473), .Z(n1171) );
  NANDN U2957 ( .A(B[29]), .B(n2474), .Z(n2473) );
  NANDN U2958 ( .A(A[29]), .B(n1225), .Z(n2474) );
  NANDN U2959 ( .A(n1225), .B(A[29]), .Z(n2472) );
  AND U2960 ( .A(n2475), .B(n2476), .Z(n1225) );
  NANDN U2961 ( .A(B[28]), .B(n2477), .Z(n2476) );
  NANDN U2962 ( .A(A[28]), .B(n1277), .Z(n2477) );
  NANDN U2963 ( .A(n1277), .B(A[28]), .Z(n2475) );
  AND U2964 ( .A(n2478), .B(n2479), .Z(n1277) );
  NANDN U2965 ( .A(B[27]), .B(n2480), .Z(n2479) );
  NANDN U2966 ( .A(A[27]), .B(n1329), .Z(n2480) );
  NANDN U2967 ( .A(n1329), .B(A[27]), .Z(n2478) );
  AND U2968 ( .A(n2481), .B(n2482), .Z(n1329) );
  NANDN U2969 ( .A(B[26]), .B(n2483), .Z(n2482) );
  NANDN U2970 ( .A(A[26]), .B(n1381), .Z(n2483) );
  NANDN U2971 ( .A(n1381), .B(A[26]), .Z(n2481) );
  AND U2972 ( .A(n2484), .B(n2485), .Z(n1381) );
  NANDN U2973 ( .A(B[25]), .B(n2486), .Z(n2485) );
  NANDN U2974 ( .A(A[25]), .B(n1433), .Z(n2486) );
  NANDN U2975 ( .A(n1433), .B(A[25]), .Z(n2484) );
  AND U2976 ( .A(n2487), .B(n2488), .Z(n1433) );
  NANDN U2977 ( .A(B[24]), .B(n2489), .Z(n2488) );
  NANDN U2978 ( .A(A[24]), .B(n1485), .Z(n2489) );
  NANDN U2979 ( .A(n1485), .B(A[24]), .Z(n2487) );
  AND U2980 ( .A(n2490), .B(n2491), .Z(n1485) );
  NANDN U2981 ( .A(B[23]), .B(n2492), .Z(n2491) );
  NANDN U2982 ( .A(A[23]), .B(n1537), .Z(n2492) );
  NANDN U2983 ( .A(n1537), .B(A[23]), .Z(n2490) );
  AND U2984 ( .A(n2493), .B(n2494), .Z(n1537) );
  NANDN U2985 ( .A(B[22]), .B(n2495), .Z(n2494) );
  NANDN U2986 ( .A(A[22]), .B(n1589), .Z(n2495) );
  NANDN U2987 ( .A(n1589), .B(A[22]), .Z(n2493) );
  AND U2988 ( .A(n2496), .B(n2497), .Z(n1589) );
  NANDN U2989 ( .A(B[21]), .B(n2498), .Z(n2497) );
  NANDN U2990 ( .A(A[21]), .B(n1641), .Z(n2498) );
  NANDN U2991 ( .A(n1641), .B(A[21]), .Z(n2496) );
  AND U2992 ( .A(n2499), .B(n2500), .Z(n1641) );
  NANDN U2993 ( .A(B[20]), .B(n2501), .Z(n2500) );
  NANDN U2994 ( .A(A[20]), .B(n1693), .Z(n2501) );
  NANDN U2995 ( .A(n1693), .B(A[20]), .Z(n2499) );
  AND U2996 ( .A(n2502), .B(n2503), .Z(n1693) );
  NANDN U2997 ( .A(B[19]), .B(n2504), .Z(n2503) );
  NANDN U2998 ( .A(A[19]), .B(n1746), .Z(n2504) );
  NANDN U2999 ( .A(n1746), .B(A[19]), .Z(n2502) );
  AND U3000 ( .A(n2505), .B(n2506), .Z(n1746) );
  NANDN U3001 ( .A(B[18]), .B(n2507), .Z(n2506) );
  NANDN U3002 ( .A(A[18]), .B(n1798), .Z(n2507) );
  NANDN U3003 ( .A(n1798), .B(A[18]), .Z(n2505) );
  AND U3004 ( .A(n2508), .B(n2509), .Z(n1798) );
  NANDN U3005 ( .A(B[17]), .B(n2510), .Z(n2509) );
  NANDN U3006 ( .A(A[17]), .B(n1850), .Z(n2510) );
  NANDN U3007 ( .A(n1850), .B(A[17]), .Z(n2508) );
  AND U3008 ( .A(n2511), .B(n2512), .Z(n1850) );
  NANDN U3009 ( .A(B[16]), .B(n2513), .Z(n2512) );
  NANDN U3010 ( .A(A[16]), .B(n1902), .Z(n2513) );
  NANDN U3011 ( .A(n1902), .B(A[16]), .Z(n2511) );
  AND U3012 ( .A(n2514), .B(n2515), .Z(n1902) );
  NANDN U3013 ( .A(B[15]), .B(n2516), .Z(n2515) );
  NANDN U3014 ( .A(A[15]), .B(n1954), .Z(n2516) );
  NANDN U3015 ( .A(n1954), .B(A[15]), .Z(n2514) );
  AND U3016 ( .A(n2517), .B(n2518), .Z(n1954) );
  NANDN U3017 ( .A(B[14]), .B(n2519), .Z(n2518) );
  NANDN U3018 ( .A(A[14]), .B(n2006), .Z(n2519) );
  NANDN U3019 ( .A(n2006), .B(A[14]), .Z(n2517) );
  AND U3020 ( .A(n2520), .B(n2521), .Z(n2006) );
  NANDN U3021 ( .A(B[13]), .B(n2522), .Z(n2521) );
  NANDN U3022 ( .A(A[13]), .B(n2058), .Z(n2522) );
  NANDN U3023 ( .A(n2058), .B(A[13]), .Z(n2520) );
  AND U3024 ( .A(n2523), .B(n2524), .Z(n2058) );
  NANDN U3025 ( .A(B[12]), .B(n2525), .Z(n2524) );
  NANDN U3026 ( .A(A[12]), .B(n2110), .Z(n2525) );
  NANDN U3027 ( .A(n2110), .B(A[12]), .Z(n2523) );
  AND U3028 ( .A(n2526), .B(n2527), .Z(n2110) );
  NANDN U3029 ( .A(B[11]), .B(n2528), .Z(n2527) );
  NANDN U3030 ( .A(A[11]), .B(n2162), .Z(n2528) );
  NANDN U3031 ( .A(n2162), .B(A[11]), .Z(n2526) );
  AND U3032 ( .A(n2529), .B(n2530), .Z(n2162) );
  NANDN U3033 ( .A(B[10]), .B(n2531), .Z(n2530) );
  NANDN U3034 ( .A(A[10]), .B(n2214), .Z(n2531) );
  NANDN U3035 ( .A(n2214), .B(A[10]), .Z(n2529) );
  AND U3036 ( .A(n2532), .B(n2533), .Z(n2214) );
  NANDN U3037 ( .A(B[9]), .B(n2534), .Z(n2533) );
  OR U3038 ( .A(n3), .B(A[9]), .Z(n2534) );
  NAND U3039 ( .A(A[9]), .B(n3), .Z(n2532) );
  NAND U3040 ( .A(n2535), .B(n2536), .Z(n3) );
  NANDN U3041 ( .A(B[8]), .B(n2537), .Z(n2536) );
  NANDN U3042 ( .A(A[8]), .B(n25), .Z(n2537) );
  NANDN U3043 ( .A(n25), .B(A[8]), .Z(n2535) );
  AND U3044 ( .A(n2538), .B(n2539), .Z(n25) );
  NANDN U3045 ( .A(B[7]), .B(n2540), .Z(n2539) );
  NANDN U3046 ( .A(A[7]), .B(n47), .Z(n2540) );
  NANDN U3047 ( .A(n47), .B(A[7]), .Z(n2538) );
  AND U3048 ( .A(n2541), .B(n2542), .Z(n47) );
  NANDN U3049 ( .A(B[6]), .B(n2543), .Z(n2542) );
  NANDN U3050 ( .A(A[6]), .B(n69), .Z(n2543) );
  NANDN U3051 ( .A(n69), .B(A[6]), .Z(n2541) );
  AND U3052 ( .A(n2544), .B(n2545), .Z(n69) );
  NANDN U3053 ( .A(B[5]), .B(n2546), .Z(n2545) );
  NANDN U3054 ( .A(A[5]), .B(n91), .Z(n2546) );
  NANDN U3055 ( .A(n91), .B(A[5]), .Z(n2544) );
  AND U3056 ( .A(n2547), .B(n2548), .Z(n91) );
  NANDN U3057 ( .A(B[4]), .B(n2549), .Z(n2548) );
  NANDN U3058 ( .A(A[4]), .B(n179), .Z(n2549) );
  NANDN U3059 ( .A(n179), .B(A[4]), .Z(n2547) );
  AND U3060 ( .A(n2550), .B(n2551), .Z(n179) );
  NANDN U3061 ( .A(B[3]), .B(n2552), .Z(n2551) );
  NANDN U3062 ( .A(A[3]), .B(n701), .Z(n2552) );
  NANDN U3063 ( .A(n701), .B(A[3]), .Z(n2550) );
  AND U3064 ( .A(n2553), .B(n2554), .Z(n701) );
  NANDN U3065 ( .A(B[2]), .B(n2555), .Z(n2554) );
  NANDN U3066 ( .A(A[2]), .B(n1223), .Z(n2555) );
  NANDN U3067 ( .A(n1223), .B(A[2]), .Z(n2553) );
  AND U3068 ( .A(n2556), .B(n2557), .Z(n1223) );
  NANDN U3069 ( .A(B[1]), .B(n2558), .Z(n2557) );
  NAND U3070 ( .A(n1), .B(n2), .Z(n2558) );
  NAND U3071 ( .A(A[1]), .B(n2559), .Z(n2556) );
  NAND U3072 ( .A(n2559), .B(n2560), .Z(DIFF[0]) );
  NANDN U3073 ( .A(B[0]), .B(A[0]), .Z(n2560) );
  NANDN U3074 ( .A(A[0]), .B(B[0]), .Z(n2559) );
endmodule


module modmult_step_N512_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [511:0] A;
  input [0:0] B;
  output [512:0] PRODUCT;
  input TC;


  AND U2 ( .A(A[511]), .B(B[0]), .Z(PRODUCT[511]) );
  AND U3 ( .A(A[510]), .B(B[0]), .Z(PRODUCT[510]) );
  AND U4 ( .A(A[509]), .B(B[0]), .Z(PRODUCT[509]) );
  AND U5 ( .A(A[508]), .B(B[0]), .Z(PRODUCT[508]) );
  AND U6 ( .A(A[507]), .B(B[0]), .Z(PRODUCT[507]) );
  AND U7 ( .A(A[506]), .B(B[0]), .Z(PRODUCT[506]) );
  AND U8 ( .A(A[505]), .B(B[0]), .Z(PRODUCT[505]) );
  AND U9 ( .A(A[504]), .B(B[0]), .Z(PRODUCT[504]) );
  AND U10 ( .A(A[503]), .B(B[0]), .Z(PRODUCT[503]) );
  AND U11 ( .A(A[502]), .B(B[0]), .Z(PRODUCT[502]) );
  AND U12 ( .A(A[501]), .B(B[0]), .Z(PRODUCT[501]) );
  AND U13 ( .A(A[500]), .B(B[0]), .Z(PRODUCT[500]) );
  AND U14 ( .A(A[499]), .B(B[0]), .Z(PRODUCT[499]) );
  AND U15 ( .A(A[498]), .B(B[0]), .Z(PRODUCT[498]) );
  AND U16 ( .A(A[497]), .B(B[0]), .Z(PRODUCT[497]) );
  AND U17 ( .A(A[496]), .B(B[0]), .Z(PRODUCT[496]) );
  AND U18 ( .A(A[495]), .B(B[0]), .Z(PRODUCT[495]) );
  AND U19 ( .A(A[494]), .B(B[0]), .Z(PRODUCT[494]) );
  AND U20 ( .A(A[493]), .B(B[0]), .Z(PRODUCT[493]) );
  AND U21 ( .A(A[492]), .B(B[0]), .Z(PRODUCT[492]) );
  AND U22 ( .A(A[491]), .B(B[0]), .Z(PRODUCT[491]) );
  AND U23 ( .A(A[490]), .B(B[0]), .Z(PRODUCT[490]) );
  AND U24 ( .A(A[489]), .B(B[0]), .Z(PRODUCT[489]) );
  AND U25 ( .A(A[488]), .B(B[0]), .Z(PRODUCT[488]) );
  AND U26 ( .A(A[487]), .B(B[0]), .Z(PRODUCT[487]) );
  AND U27 ( .A(A[486]), .B(B[0]), .Z(PRODUCT[486]) );
  AND U28 ( .A(A[485]), .B(B[0]), .Z(PRODUCT[485]) );
  AND U29 ( .A(A[484]), .B(B[0]), .Z(PRODUCT[484]) );
  AND U30 ( .A(A[483]), .B(B[0]), .Z(PRODUCT[483]) );
  AND U31 ( .A(A[482]), .B(B[0]), .Z(PRODUCT[482]) );
  AND U32 ( .A(A[481]), .B(B[0]), .Z(PRODUCT[481]) );
  AND U33 ( .A(A[480]), .B(B[0]), .Z(PRODUCT[480]) );
  AND U34 ( .A(A[479]), .B(B[0]), .Z(PRODUCT[479]) );
  AND U35 ( .A(A[478]), .B(B[0]), .Z(PRODUCT[478]) );
  AND U36 ( .A(A[477]), .B(B[0]), .Z(PRODUCT[477]) );
  AND U37 ( .A(A[476]), .B(B[0]), .Z(PRODUCT[476]) );
  AND U38 ( .A(A[475]), .B(B[0]), .Z(PRODUCT[475]) );
  AND U39 ( .A(A[474]), .B(B[0]), .Z(PRODUCT[474]) );
  AND U40 ( .A(A[473]), .B(B[0]), .Z(PRODUCT[473]) );
  AND U41 ( .A(A[472]), .B(B[0]), .Z(PRODUCT[472]) );
  AND U42 ( .A(A[471]), .B(B[0]), .Z(PRODUCT[471]) );
  AND U43 ( .A(A[470]), .B(B[0]), .Z(PRODUCT[470]) );
  AND U44 ( .A(A[469]), .B(B[0]), .Z(PRODUCT[469]) );
  AND U45 ( .A(A[468]), .B(B[0]), .Z(PRODUCT[468]) );
  AND U46 ( .A(A[467]), .B(B[0]), .Z(PRODUCT[467]) );
  AND U47 ( .A(A[466]), .B(B[0]), .Z(PRODUCT[466]) );
  AND U48 ( .A(A[465]), .B(B[0]), .Z(PRODUCT[465]) );
  AND U49 ( .A(A[464]), .B(B[0]), .Z(PRODUCT[464]) );
  AND U50 ( .A(A[463]), .B(B[0]), .Z(PRODUCT[463]) );
  AND U51 ( .A(A[462]), .B(B[0]), .Z(PRODUCT[462]) );
  AND U52 ( .A(A[461]), .B(B[0]), .Z(PRODUCT[461]) );
  AND U53 ( .A(A[460]), .B(B[0]), .Z(PRODUCT[460]) );
  AND U54 ( .A(A[459]), .B(B[0]), .Z(PRODUCT[459]) );
  AND U55 ( .A(A[458]), .B(B[0]), .Z(PRODUCT[458]) );
  AND U56 ( .A(A[457]), .B(B[0]), .Z(PRODUCT[457]) );
  AND U57 ( .A(A[456]), .B(B[0]), .Z(PRODUCT[456]) );
  AND U58 ( .A(A[455]), .B(B[0]), .Z(PRODUCT[455]) );
  AND U59 ( .A(A[454]), .B(B[0]), .Z(PRODUCT[454]) );
  AND U60 ( .A(A[453]), .B(B[0]), .Z(PRODUCT[453]) );
  AND U61 ( .A(A[452]), .B(B[0]), .Z(PRODUCT[452]) );
  AND U62 ( .A(A[451]), .B(B[0]), .Z(PRODUCT[451]) );
  AND U63 ( .A(A[450]), .B(B[0]), .Z(PRODUCT[450]) );
  AND U64 ( .A(A[449]), .B(B[0]), .Z(PRODUCT[449]) );
  AND U65 ( .A(A[448]), .B(B[0]), .Z(PRODUCT[448]) );
  AND U66 ( .A(A[447]), .B(B[0]), .Z(PRODUCT[447]) );
  AND U67 ( .A(A[446]), .B(B[0]), .Z(PRODUCT[446]) );
  AND U68 ( .A(A[445]), .B(B[0]), .Z(PRODUCT[445]) );
  AND U69 ( .A(A[444]), .B(B[0]), .Z(PRODUCT[444]) );
  AND U70 ( .A(A[443]), .B(B[0]), .Z(PRODUCT[443]) );
  AND U71 ( .A(A[442]), .B(B[0]), .Z(PRODUCT[442]) );
  AND U72 ( .A(A[441]), .B(B[0]), .Z(PRODUCT[441]) );
  AND U73 ( .A(A[440]), .B(B[0]), .Z(PRODUCT[440]) );
  AND U74 ( .A(A[439]), .B(B[0]), .Z(PRODUCT[439]) );
  AND U75 ( .A(A[438]), .B(B[0]), .Z(PRODUCT[438]) );
  AND U76 ( .A(A[437]), .B(B[0]), .Z(PRODUCT[437]) );
  AND U77 ( .A(A[436]), .B(B[0]), .Z(PRODUCT[436]) );
  AND U78 ( .A(A[435]), .B(B[0]), .Z(PRODUCT[435]) );
  AND U79 ( .A(A[434]), .B(B[0]), .Z(PRODUCT[434]) );
  AND U80 ( .A(A[433]), .B(B[0]), .Z(PRODUCT[433]) );
  AND U81 ( .A(A[432]), .B(B[0]), .Z(PRODUCT[432]) );
  AND U82 ( .A(A[431]), .B(B[0]), .Z(PRODUCT[431]) );
  AND U83 ( .A(A[430]), .B(B[0]), .Z(PRODUCT[430]) );
  AND U84 ( .A(A[429]), .B(B[0]), .Z(PRODUCT[429]) );
  AND U85 ( .A(A[428]), .B(B[0]), .Z(PRODUCT[428]) );
  AND U86 ( .A(A[427]), .B(B[0]), .Z(PRODUCT[427]) );
  AND U87 ( .A(A[426]), .B(B[0]), .Z(PRODUCT[426]) );
  AND U88 ( .A(A[425]), .B(B[0]), .Z(PRODUCT[425]) );
  AND U89 ( .A(A[424]), .B(B[0]), .Z(PRODUCT[424]) );
  AND U90 ( .A(A[423]), .B(B[0]), .Z(PRODUCT[423]) );
  AND U91 ( .A(A[422]), .B(B[0]), .Z(PRODUCT[422]) );
  AND U92 ( .A(A[421]), .B(B[0]), .Z(PRODUCT[421]) );
  AND U93 ( .A(A[420]), .B(B[0]), .Z(PRODUCT[420]) );
  AND U94 ( .A(A[419]), .B(B[0]), .Z(PRODUCT[419]) );
  AND U95 ( .A(A[418]), .B(B[0]), .Z(PRODUCT[418]) );
  AND U96 ( .A(A[417]), .B(B[0]), .Z(PRODUCT[417]) );
  AND U97 ( .A(A[416]), .B(B[0]), .Z(PRODUCT[416]) );
  AND U98 ( .A(A[415]), .B(B[0]), .Z(PRODUCT[415]) );
  AND U99 ( .A(A[414]), .B(B[0]), .Z(PRODUCT[414]) );
  AND U100 ( .A(A[413]), .B(B[0]), .Z(PRODUCT[413]) );
  AND U101 ( .A(A[412]), .B(B[0]), .Z(PRODUCT[412]) );
  AND U102 ( .A(A[411]), .B(B[0]), .Z(PRODUCT[411]) );
  AND U103 ( .A(A[410]), .B(B[0]), .Z(PRODUCT[410]) );
  AND U104 ( .A(A[409]), .B(B[0]), .Z(PRODUCT[409]) );
  AND U105 ( .A(A[408]), .B(B[0]), .Z(PRODUCT[408]) );
  AND U106 ( .A(A[407]), .B(B[0]), .Z(PRODUCT[407]) );
  AND U107 ( .A(A[406]), .B(B[0]), .Z(PRODUCT[406]) );
  AND U108 ( .A(A[405]), .B(B[0]), .Z(PRODUCT[405]) );
  AND U109 ( .A(A[404]), .B(B[0]), .Z(PRODUCT[404]) );
  AND U110 ( .A(A[403]), .B(B[0]), .Z(PRODUCT[403]) );
  AND U111 ( .A(A[402]), .B(B[0]), .Z(PRODUCT[402]) );
  AND U112 ( .A(A[401]), .B(B[0]), .Z(PRODUCT[401]) );
  AND U113 ( .A(A[400]), .B(B[0]), .Z(PRODUCT[400]) );
  AND U114 ( .A(A[399]), .B(B[0]), .Z(PRODUCT[399]) );
  AND U115 ( .A(A[398]), .B(B[0]), .Z(PRODUCT[398]) );
  AND U116 ( .A(A[397]), .B(B[0]), .Z(PRODUCT[397]) );
  AND U117 ( .A(A[396]), .B(B[0]), .Z(PRODUCT[396]) );
  AND U118 ( .A(A[395]), .B(B[0]), .Z(PRODUCT[395]) );
  AND U119 ( .A(A[394]), .B(B[0]), .Z(PRODUCT[394]) );
  AND U120 ( .A(A[393]), .B(B[0]), .Z(PRODUCT[393]) );
  AND U121 ( .A(A[392]), .B(B[0]), .Z(PRODUCT[392]) );
  AND U122 ( .A(A[391]), .B(B[0]), .Z(PRODUCT[391]) );
  AND U123 ( .A(A[390]), .B(B[0]), .Z(PRODUCT[390]) );
  AND U124 ( .A(A[389]), .B(B[0]), .Z(PRODUCT[389]) );
  AND U125 ( .A(A[388]), .B(B[0]), .Z(PRODUCT[388]) );
  AND U126 ( .A(A[387]), .B(B[0]), .Z(PRODUCT[387]) );
  AND U127 ( .A(A[386]), .B(B[0]), .Z(PRODUCT[386]) );
  AND U128 ( .A(A[385]), .B(B[0]), .Z(PRODUCT[385]) );
  AND U129 ( .A(A[384]), .B(B[0]), .Z(PRODUCT[384]) );
  AND U130 ( .A(A[383]), .B(B[0]), .Z(PRODUCT[383]) );
  AND U131 ( .A(A[382]), .B(B[0]), .Z(PRODUCT[382]) );
  AND U132 ( .A(A[381]), .B(B[0]), .Z(PRODUCT[381]) );
  AND U133 ( .A(A[380]), .B(B[0]), .Z(PRODUCT[380]) );
  AND U134 ( .A(A[379]), .B(B[0]), .Z(PRODUCT[379]) );
  AND U135 ( .A(A[378]), .B(B[0]), .Z(PRODUCT[378]) );
  AND U136 ( .A(A[377]), .B(B[0]), .Z(PRODUCT[377]) );
  AND U137 ( .A(A[376]), .B(B[0]), .Z(PRODUCT[376]) );
  AND U138 ( .A(A[375]), .B(B[0]), .Z(PRODUCT[375]) );
  AND U139 ( .A(A[374]), .B(B[0]), .Z(PRODUCT[374]) );
  AND U140 ( .A(A[373]), .B(B[0]), .Z(PRODUCT[373]) );
  AND U141 ( .A(A[372]), .B(B[0]), .Z(PRODUCT[372]) );
  AND U142 ( .A(A[371]), .B(B[0]), .Z(PRODUCT[371]) );
  AND U143 ( .A(A[370]), .B(B[0]), .Z(PRODUCT[370]) );
  AND U144 ( .A(A[369]), .B(B[0]), .Z(PRODUCT[369]) );
  AND U145 ( .A(A[368]), .B(B[0]), .Z(PRODUCT[368]) );
  AND U146 ( .A(A[367]), .B(B[0]), .Z(PRODUCT[367]) );
  AND U147 ( .A(A[366]), .B(B[0]), .Z(PRODUCT[366]) );
  AND U148 ( .A(A[365]), .B(B[0]), .Z(PRODUCT[365]) );
  AND U149 ( .A(A[364]), .B(B[0]), .Z(PRODUCT[364]) );
  AND U150 ( .A(A[363]), .B(B[0]), .Z(PRODUCT[363]) );
  AND U151 ( .A(A[362]), .B(B[0]), .Z(PRODUCT[362]) );
  AND U152 ( .A(A[361]), .B(B[0]), .Z(PRODUCT[361]) );
  AND U153 ( .A(A[360]), .B(B[0]), .Z(PRODUCT[360]) );
  AND U154 ( .A(A[359]), .B(B[0]), .Z(PRODUCT[359]) );
  AND U155 ( .A(A[358]), .B(B[0]), .Z(PRODUCT[358]) );
  AND U156 ( .A(A[357]), .B(B[0]), .Z(PRODUCT[357]) );
  AND U157 ( .A(A[356]), .B(B[0]), .Z(PRODUCT[356]) );
  AND U158 ( .A(A[355]), .B(B[0]), .Z(PRODUCT[355]) );
  AND U159 ( .A(A[354]), .B(B[0]), .Z(PRODUCT[354]) );
  AND U160 ( .A(A[353]), .B(B[0]), .Z(PRODUCT[353]) );
  AND U161 ( .A(A[352]), .B(B[0]), .Z(PRODUCT[352]) );
  AND U162 ( .A(A[351]), .B(B[0]), .Z(PRODUCT[351]) );
  AND U163 ( .A(A[350]), .B(B[0]), .Z(PRODUCT[350]) );
  AND U164 ( .A(A[349]), .B(B[0]), .Z(PRODUCT[349]) );
  AND U165 ( .A(A[348]), .B(B[0]), .Z(PRODUCT[348]) );
  AND U166 ( .A(A[347]), .B(B[0]), .Z(PRODUCT[347]) );
  AND U167 ( .A(A[346]), .B(B[0]), .Z(PRODUCT[346]) );
  AND U168 ( .A(A[345]), .B(B[0]), .Z(PRODUCT[345]) );
  AND U169 ( .A(A[344]), .B(B[0]), .Z(PRODUCT[344]) );
  AND U170 ( .A(A[343]), .B(B[0]), .Z(PRODUCT[343]) );
  AND U171 ( .A(A[342]), .B(B[0]), .Z(PRODUCT[342]) );
  AND U172 ( .A(A[341]), .B(B[0]), .Z(PRODUCT[341]) );
  AND U173 ( .A(A[340]), .B(B[0]), .Z(PRODUCT[340]) );
  AND U174 ( .A(A[339]), .B(B[0]), .Z(PRODUCT[339]) );
  AND U175 ( .A(A[338]), .B(B[0]), .Z(PRODUCT[338]) );
  AND U176 ( .A(A[337]), .B(B[0]), .Z(PRODUCT[337]) );
  AND U177 ( .A(A[336]), .B(B[0]), .Z(PRODUCT[336]) );
  AND U178 ( .A(A[335]), .B(B[0]), .Z(PRODUCT[335]) );
  AND U179 ( .A(A[334]), .B(B[0]), .Z(PRODUCT[334]) );
  AND U180 ( .A(A[333]), .B(B[0]), .Z(PRODUCT[333]) );
  AND U181 ( .A(A[332]), .B(B[0]), .Z(PRODUCT[332]) );
  AND U182 ( .A(A[331]), .B(B[0]), .Z(PRODUCT[331]) );
  AND U183 ( .A(A[330]), .B(B[0]), .Z(PRODUCT[330]) );
  AND U184 ( .A(A[329]), .B(B[0]), .Z(PRODUCT[329]) );
  AND U185 ( .A(A[328]), .B(B[0]), .Z(PRODUCT[328]) );
  AND U186 ( .A(A[327]), .B(B[0]), .Z(PRODUCT[327]) );
  AND U187 ( .A(A[326]), .B(B[0]), .Z(PRODUCT[326]) );
  AND U188 ( .A(A[325]), .B(B[0]), .Z(PRODUCT[325]) );
  AND U189 ( .A(A[324]), .B(B[0]), .Z(PRODUCT[324]) );
  AND U190 ( .A(A[323]), .B(B[0]), .Z(PRODUCT[323]) );
  AND U191 ( .A(A[322]), .B(B[0]), .Z(PRODUCT[322]) );
  AND U192 ( .A(A[321]), .B(B[0]), .Z(PRODUCT[321]) );
  AND U193 ( .A(A[320]), .B(B[0]), .Z(PRODUCT[320]) );
  AND U194 ( .A(A[319]), .B(B[0]), .Z(PRODUCT[319]) );
  AND U195 ( .A(A[318]), .B(B[0]), .Z(PRODUCT[318]) );
  AND U196 ( .A(A[317]), .B(B[0]), .Z(PRODUCT[317]) );
  AND U197 ( .A(A[316]), .B(B[0]), .Z(PRODUCT[316]) );
  AND U198 ( .A(A[315]), .B(B[0]), .Z(PRODUCT[315]) );
  AND U199 ( .A(A[314]), .B(B[0]), .Z(PRODUCT[314]) );
  AND U200 ( .A(A[313]), .B(B[0]), .Z(PRODUCT[313]) );
  AND U201 ( .A(A[312]), .B(B[0]), .Z(PRODUCT[312]) );
  AND U202 ( .A(A[311]), .B(B[0]), .Z(PRODUCT[311]) );
  AND U203 ( .A(A[310]), .B(B[0]), .Z(PRODUCT[310]) );
  AND U204 ( .A(A[309]), .B(B[0]), .Z(PRODUCT[309]) );
  AND U205 ( .A(A[308]), .B(B[0]), .Z(PRODUCT[308]) );
  AND U206 ( .A(A[307]), .B(B[0]), .Z(PRODUCT[307]) );
  AND U207 ( .A(A[306]), .B(B[0]), .Z(PRODUCT[306]) );
  AND U208 ( .A(A[305]), .B(B[0]), .Z(PRODUCT[305]) );
  AND U209 ( .A(A[304]), .B(B[0]), .Z(PRODUCT[304]) );
  AND U210 ( .A(A[303]), .B(B[0]), .Z(PRODUCT[303]) );
  AND U211 ( .A(A[302]), .B(B[0]), .Z(PRODUCT[302]) );
  AND U212 ( .A(A[301]), .B(B[0]), .Z(PRODUCT[301]) );
  AND U213 ( .A(A[300]), .B(B[0]), .Z(PRODUCT[300]) );
  AND U214 ( .A(A[299]), .B(B[0]), .Z(PRODUCT[299]) );
  AND U215 ( .A(A[298]), .B(B[0]), .Z(PRODUCT[298]) );
  AND U216 ( .A(A[297]), .B(B[0]), .Z(PRODUCT[297]) );
  AND U217 ( .A(A[296]), .B(B[0]), .Z(PRODUCT[296]) );
  AND U218 ( .A(A[295]), .B(B[0]), .Z(PRODUCT[295]) );
  AND U219 ( .A(A[294]), .B(B[0]), .Z(PRODUCT[294]) );
  AND U220 ( .A(A[293]), .B(B[0]), .Z(PRODUCT[293]) );
  AND U221 ( .A(A[292]), .B(B[0]), .Z(PRODUCT[292]) );
  AND U222 ( .A(A[291]), .B(B[0]), .Z(PRODUCT[291]) );
  AND U223 ( .A(A[290]), .B(B[0]), .Z(PRODUCT[290]) );
  AND U224 ( .A(A[289]), .B(B[0]), .Z(PRODUCT[289]) );
  AND U225 ( .A(A[288]), .B(B[0]), .Z(PRODUCT[288]) );
  AND U226 ( .A(A[287]), .B(B[0]), .Z(PRODUCT[287]) );
  AND U227 ( .A(A[286]), .B(B[0]), .Z(PRODUCT[286]) );
  AND U228 ( .A(A[285]), .B(B[0]), .Z(PRODUCT[285]) );
  AND U229 ( .A(A[284]), .B(B[0]), .Z(PRODUCT[284]) );
  AND U230 ( .A(A[283]), .B(B[0]), .Z(PRODUCT[283]) );
  AND U231 ( .A(A[282]), .B(B[0]), .Z(PRODUCT[282]) );
  AND U232 ( .A(A[281]), .B(B[0]), .Z(PRODUCT[281]) );
  AND U233 ( .A(A[280]), .B(B[0]), .Z(PRODUCT[280]) );
  AND U234 ( .A(A[279]), .B(B[0]), .Z(PRODUCT[279]) );
  AND U235 ( .A(A[278]), .B(B[0]), .Z(PRODUCT[278]) );
  AND U236 ( .A(A[277]), .B(B[0]), .Z(PRODUCT[277]) );
  AND U237 ( .A(A[276]), .B(B[0]), .Z(PRODUCT[276]) );
  AND U238 ( .A(A[275]), .B(B[0]), .Z(PRODUCT[275]) );
  AND U239 ( .A(A[274]), .B(B[0]), .Z(PRODUCT[274]) );
  AND U240 ( .A(A[273]), .B(B[0]), .Z(PRODUCT[273]) );
  AND U241 ( .A(A[272]), .B(B[0]), .Z(PRODUCT[272]) );
  AND U242 ( .A(A[271]), .B(B[0]), .Z(PRODUCT[271]) );
  AND U243 ( .A(A[270]), .B(B[0]), .Z(PRODUCT[270]) );
  AND U244 ( .A(A[269]), .B(B[0]), .Z(PRODUCT[269]) );
  AND U245 ( .A(A[268]), .B(B[0]), .Z(PRODUCT[268]) );
  AND U246 ( .A(A[267]), .B(B[0]), .Z(PRODUCT[267]) );
  AND U247 ( .A(A[266]), .B(B[0]), .Z(PRODUCT[266]) );
  AND U248 ( .A(A[265]), .B(B[0]), .Z(PRODUCT[265]) );
  AND U249 ( .A(A[264]), .B(B[0]), .Z(PRODUCT[264]) );
  AND U250 ( .A(A[263]), .B(B[0]), .Z(PRODUCT[263]) );
  AND U251 ( .A(A[262]), .B(B[0]), .Z(PRODUCT[262]) );
  AND U252 ( .A(A[261]), .B(B[0]), .Z(PRODUCT[261]) );
  AND U253 ( .A(A[260]), .B(B[0]), .Z(PRODUCT[260]) );
  AND U254 ( .A(A[259]), .B(B[0]), .Z(PRODUCT[259]) );
  AND U255 ( .A(A[258]), .B(B[0]), .Z(PRODUCT[258]) );
  AND U256 ( .A(A[257]), .B(B[0]), .Z(PRODUCT[257]) );
  AND U257 ( .A(A[256]), .B(B[0]), .Z(PRODUCT[256]) );
  AND U258 ( .A(A[255]), .B(B[0]), .Z(PRODUCT[255]) );
  AND U259 ( .A(A[254]), .B(B[0]), .Z(PRODUCT[254]) );
  AND U260 ( .A(A[253]), .B(B[0]), .Z(PRODUCT[253]) );
  AND U261 ( .A(A[252]), .B(B[0]), .Z(PRODUCT[252]) );
  AND U262 ( .A(A[251]), .B(B[0]), .Z(PRODUCT[251]) );
  AND U263 ( .A(A[250]), .B(B[0]), .Z(PRODUCT[250]) );
  AND U264 ( .A(A[249]), .B(B[0]), .Z(PRODUCT[249]) );
  AND U265 ( .A(A[248]), .B(B[0]), .Z(PRODUCT[248]) );
  AND U266 ( .A(A[247]), .B(B[0]), .Z(PRODUCT[247]) );
  AND U267 ( .A(A[246]), .B(B[0]), .Z(PRODUCT[246]) );
  AND U268 ( .A(A[245]), .B(B[0]), .Z(PRODUCT[245]) );
  AND U269 ( .A(A[244]), .B(B[0]), .Z(PRODUCT[244]) );
  AND U270 ( .A(A[243]), .B(B[0]), .Z(PRODUCT[243]) );
  AND U271 ( .A(A[242]), .B(B[0]), .Z(PRODUCT[242]) );
  AND U272 ( .A(A[241]), .B(B[0]), .Z(PRODUCT[241]) );
  AND U273 ( .A(A[240]), .B(B[0]), .Z(PRODUCT[240]) );
  AND U274 ( .A(A[239]), .B(B[0]), .Z(PRODUCT[239]) );
  AND U275 ( .A(A[238]), .B(B[0]), .Z(PRODUCT[238]) );
  AND U276 ( .A(A[237]), .B(B[0]), .Z(PRODUCT[237]) );
  AND U277 ( .A(A[236]), .B(B[0]), .Z(PRODUCT[236]) );
  AND U278 ( .A(A[235]), .B(B[0]), .Z(PRODUCT[235]) );
  AND U279 ( .A(A[234]), .B(B[0]), .Z(PRODUCT[234]) );
  AND U280 ( .A(A[233]), .B(B[0]), .Z(PRODUCT[233]) );
  AND U281 ( .A(A[232]), .B(B[0]), .Z(PRODUCT[232]) );
  AND U282 ( .A(A[231]), .B(B[0]), .Z(PRODUCT[231]) );
  AND U283 ( .A(A[230]), .B(B[0]), .Z(PRODUCT[230]) );
  AND U284 ( .A(A[229]), .B(B[0]), .Z(PRODUCT[229]) );
  AND U285 ( .A(A[228]), .B(B[0]), .Z(PRODUCT[228]) );
  AND U286 ( .A(A[227]), .B(B[0]), .Z(PRODUCT[227]) );
  AND U287 ( .A(A[226]), .B(B[0]), .Z(PRODUCT[226]) );
  AND U288 ( .A(A[225]), .B(B[0]), .Z(PRODUCT[225]) );
  AND U289 ( .A(A[224]), .B(B[0]), .Z(PRODUCT[224]) );
  AND U290 ( .A(A[223]), .B(B[0]), .Z(PRODUCT[223]) );
  AND U291 ( .A(A[222]), .B(B[0]), .Z(PRODUCT[222]) );
  AND U292 ( .A(A[221]), .B(B[0]), .Z(PRODUCT[221]) );
  AND U293 ( .A(A[220]), .B(B[0]), .Z(PRODUCT[220]) );
  AND U294 ( .A(A[219]), .B(B[0]), .Z(PRODUCT[219]) );
  AND U295 ( .A(A[218]), .B(B[0]), .Z(PRODUCT[218]) );
  AND U296 ( .A(A[217]), .B(B[0]), .Z(PRODUCT[217]) );
  AND U297 ( .A(A[216]), .B(B[0]), .Z(PRODUCT[216]) );
  AND U298 ( .A(A[215]), .B(B[0]), .Z(PRODUCT[215]) );
  AND U299 ( .A(A[214]), .B(B[0]), .Z(PRODUCT[214]) );
  AND U300 ( .A(A[213]), .B(B[0]), .Z(PRODUCT[213]) );
  AND U301 ( .A(A[212]), .B(B[0]), .Z(PRODUCT[212]) );
  AND U302 ( .A(A[211]), .B(B[0]), .Z(PRODUCT[211]) );
  AND U303 ( .A(A[210]), .B(B[0]), .Z(PRODUCT[210]) );
  AND U304 ( .A(A[209]), .B(B[0]), .Z(PRODUCT[209]) );
  AND U305 ( .A(A[208]), .B(B[0]), .Z(PRODUCT[208]) );
  AND U306 ( .A(A[207]), .B(B[0]), .Z(PRODUCT[207]) );
  AND U307 ( .A(A[206]), .B(B[0]), .Z(PRODUCT[206]) );
  AND U308 ( .A(A[205]), .B(B[0]), .Z(PRODUCT[205]) );
  AND U309 ( .A(A[204]), .B(B[0]), .Z(PRODUCT[204]) );
  AND U310 ( .A(A[203]), .B(B[0]), .Z(PRODUCT[203]) );
  AND U311 ( .A(A[202]), .B(B[0]), .Z(PRODUCT[202]) );
  AND U312 ( .A(A[201]), .B(B[0]), .Z(PRODUCT[201]) );
  AND U313 ( .A(A[200]), .B(B[0]), .Z(PRODUCT[200]) );
  AND U314 ( .A(A[199]), .B(B[0]), .Z(PRODUCT[199]) );
  AND U315 ( .A(A[198]), .B(B[0]), .Z(PRODUCT[198]) );
  AND U316 ( .A(A[197]), .B(B[0]), .Z(PRODUCT[197]) );
  AND U317 ( .A(A[196]), .B(B[0]), .Z(PRODUCT[196]) );
  AND U318 ( .A(A[195]), .B(B[0]), .Z(PRODUCT[195]) );
  AND U319 ( .A(A[194]), .B(B[0]), .Z(PRODUCT[194]) );
  AND U320 ( .A(A[193]), .B(B[0]), .Z(PRODUCT[193]) );
  AND U321 ( .A(A[192]), .B(B[0]), .Z(PRODUCT[192]) );
  AND U322 ( .A(A[191]), .B(B[0]), .Z(PRODUCT[191]) );
  AND U323 ( .A(A[190]), .B(B[0]), .Z(PRODUCT[190]) );
  AND U324 ( .A(A[189]), .B(B[0]), .Z(PRODUCT[189]) );
  AND U325 ( .A(A[188]), .B(B[0]), .Z(PRODUCT[188]) );
  AND U326 ( .A(A[187]), .B(B[0]), .Z(PRODUCT[187]) );
  AND U327 ( .A(A[186]), .B(B[0]), .Z(PRODUCT[186]) );
  AND U328 ( .A(A[185]), .B(B[0]), .Z(PRODUCT[185]) );
  AND U329 ( .A(A[184]), .B(B[0]), .Z(PRODUCT[184]) );
  AND U330 ( .A(A[183]), .B(B[0]), .Z(PRODUCT[183]) );
  AND U331 ( .A(A[182]), .B(B[0]), .Z(PRODUCT[182]) );
  AND U332 ( .A(A[181]), .B(B[0]), .Z(PRODUCT[181]) );
  AND U333 ( .A(A[180]), .B(B[0]), .Z(PRODUCT[180]) );
  AND U334 ( .A(A[179]), .B(B[0]), .Z(PRODUCT[179]) );
  AND U335 ( .A(A[178]), .B(B[0]), .Z(PRODUCT[178]) );
  AND U336 ( .A(A[177]), .B(B[0]), .Z(PRODUCT[177]) );
  AND U337 ( .A(A[176]), .B(B[0]), .Z(PRODUCT[176]) );
  AND U338 ( .A(A[175]), .B(B[0]), .Z(PRODUCT[175]) );
  AND U339 ( .A(A[174]), .B(B[0]), .Z(PRODUCT[174]) );
  AND U340 ( .A(A[173]), .B(B[0]), .Z(PRODUCT[173]) );
  AND U341 ( .A(A[172]), .B(B[0]), .Z(PRODUCT[172]) );
  AND U342 ( .A(A[171]), .B(B[0]), .Z(PRODUCT[171]) );
  AND U343 ( .A(A[170]), .B(B[0]), .Z(PRODUCT[170]) );
  AND U344 ( .A(A[169]), .B(B[0]), .Z(PRODUCT[169]) );
  AND U345 ( .A(A[168]), .B(B[0]), .Z(PRODUCT[168]) );
  AND U346 ( .A(A[167]), .B(B[0]), .Z(PRODUCT[167]) );
  AND U347 ( .A(A[166]), .B(B[0]), .Z(PRODUCT[166]) );
  AND U348 ( .A(A[165]), .B(B[0]), .Z(PRODUCT[165]) );
  AND U349 ( .A(A[164]), .B(B[0]), .Z(PRODUCT[164]) );
  AND U350 ( .A(A[163]), .B(B[0]), .Z(PRODUCT[163]) );
  AND U351 ( .A(A[162]), .B(B[0]), .Z(PRODUCT[162]) );
  AND U352 ( .A(A[161]), .B(B[0]), .Z(PRODUCT[161]) );
  AND U353 ( .A(A[160]), .B(B[0]), .Z(PRODUCT[160]) );
  AND U354 ( .A(A[159]), .B(B[0]), .Z(PRODUCT[159]) );
  AND U355 ( .A(A[158]), .B(B[0]), .Z(PRODUCT[158]) );
  AND U356 ( .A(A[157]), .B(B[0]), .Z(PRODUCT[157]) );
  AND U357 ( .A(A[156]), .B(B[0]), .Z(PRODUCT[156]) );
  AND U358 ( .A(A[155]), .B(B[0]), .Z(PRODUCT[155]) );
  AND U359 ( .A(A[154]), .B(B[0]), .Z(PRODUCT[154]) );
  AND U360 ( .A(A[153]), .B(B[0]), .Z(PRODUCT[153]) );
  AND U361 ( .A(A[152]), .B(B[0]), .Z(PRODUCT[152]) );
  AND U362 ( .A(A[151]), .B(B[0]), .Z(PRODUCT[151]) );
  AND U363 ( .A(A[150]), .B(B[0]), .Z(PRODUCT[150]) );
  AND U364 ( .A(A[149]), .B(B[0]), .Z(PRODUCT[149]) );
  AND U365 ( .A(A[148]), .B(B[0]), .Z(PRODUCT[148]) );
  AND U366 ( .A(A[147]), .B(B[0]), .Z(PRODUCT[147]) );
  AND U367 ( .A(A[146]), .B(B[0]), .Z(PRODUCT[146]) );
  AND U368 ( .A(A[145]), .B(B[0]), .Z(PRODUCT[145]) );
  AND U369 ( .A(A[144]), .B(B[0]), .Z(PRODUCT[144]) );
  AND U370 ( .A(A[143]), .B(B[0]), .Z(PRODUCT[143]) );
  AND U371 ( .A(A[142]), .B(B[0]), .Z(PRODUCT[142]) );
  AND U372 ( .A(A[141]), .B(B[0]), .Z(PRODUCT[141]) );
  AND U373 ( .A(A[140]), .B(B[0]), .Z(PRODUCT[140]) );
  AND U374 ( .A(A[139]), .B(B[0]), .Z(PRODUCT[139]) );
  AND U375 ( .A(A[138]), .B(B[0]), .Z(PRODUCT[138]) );
  AND U376 ( .A(A[137]), .B(B[0]), .Z(PRODUCT[137]) );
  AND U377 ( .A(A[136]), .B(B[0]), .Z(PRODUCT[136]) );
  AND U378 ( .A(A[135]), .B(B[0]), .Z(PRODUCT[135]) );
  AND U379 ( .A(A[134]), .B(B[0]), .Z(PRODUCT[134]) );
  AND U380 ( .A(A[133]), .B(B[0]), .Z(PRODUCT[133]) );
  AND U381 ( .A(A[132]), .B(B[0]), .Z(PRODUCT[132]) );
  AND U382 ( .A(A[131]), .B(B[0]), .Z(PRODUCT[131]) );
  AND U383 ( .A(A[130]), .B(B[0]), .Z(PRODUCT[130]) );
  AND U384 ( .A(A[129]), .B(B[0]), .Z(PRODUCT[129]) );
  AND U385 ( .A(A[128]), .B(B[0]), .Z(PRODUCT[128]) );
  AND U386 ( .A(A[127]), .B(B[0]), .Z(PRODUCT[127]) );
  AND U387 ( .A(A[126]), .B(B[0]), .Z(PRODUCT[126]) );
  AND U388 ( .A(A[125]), .B(B[0]), .Z(PRODUCT[125]) );
  AND U389 ( .A(A[124]), .B(B[0]), .Z(PRODUCT[124]) );
  AND U390 ( .A(A[123]), .B(B[0]), .Z(PRODUCT[123]) );
  AND U391 ( .A(A[122]), .B(B[0]), .Z(PRODUCT[122]) );
  AND U392 ( .A(A[121]), .B(B[0]), .Z(PRODUCT[121]) );
  AND U393 ( .A(A[120]), .B(B[0]), .Z(PRODUCT[120]) );
  AND U394 ( .A(A[119]), .B(B[0]), .Z(PRODUCT[119]) );
  AND U395 ( .A(A[118]), .B(B[0]), .Z(PRODUCT[118]) );
  AND U396 ( .A(A[117]), .B(B[0]), .Z(PRODUCT[117]) );
  AND U397 ( .A(A[116]), .B(B[0]), .Z(PRODUCT[116]) );
  AND U398 ( .A(A[115]), .B(B[0]), .Z(PRODUCT[115]) );
  AND U399 ( .A(A[114]), .B(B[0]), .Z(PRODUCT[114]) );
  AND U400 ( .A(A[113]), .B(B[0]), .Z(PRODUCT[113]) );
  AND U401 ( .A(A[112]), .B(B[0]), .Z(PRODUCT[112]) );
  AND U402 ( .A(A[111]), .B(B[0]), .Z(PRODUCT[111]) );
  AND U403 ( .A(A[110]), .B(B[0]), .Z(PRODUCT[110]) );
  AND U404 ( .A(A[109]), .B(B[0]), .Z(PRODUCT[109]) );
  AND U405 ( .A(A[108]), .B(B[0]), .Z(PRODUCT[108]) );
  AND U406 ( .A(A[107]), .B(B[0]), .Z(PRODUCT[107]) );
  AND U407 ( .A(A[106]), .B(B[0]), .Z(PRODUCT[106]) );
  AND U408 ( .A(A[105]), .B(B[0]), .Z(PRODUCT[105]) );
  AND U409 ( .A(A[104]), .B(B[0]), .Z(PRODUCT[104]) );
  AND U410 ( .A(A[103]), .B(B[0]), .Z(PRODUCT[103]) );
  AND U411 ( .A(A[102]), .B(B[0]), .Z(PRODUCT[102]) );
  AND U412 ( .A(A[101]), .B(B[0]), .Z(PRODUCT[101]) );
  AND U413 ( .A(A[100]), .B(B[0]), .Z(PRODUCT[100]) );
  AND U414 ( .A(A[99]), .B(B[0]), .Z(PRODUCT[99]) );
  AND U415 ( .A(A[98]), .B(B[0]), .Z(PRODUCT[98]) );
  AND U416 ( .A(A[97]), .B(B[0]), .Z(PRODUCT[97]) );
  AND U417 ( .A(A[96]), .B(B[0]), .Z(PRODUCT[96]) );
  AND U418 ( .A(A[95]), .B(B[0]), .Z(PRODUCT[95]) );
  AND U419 ( .A(A[94]), .B(B[0]), .Z(PRODUCT[94]) );
  AND U420 ( .A(A[93]), .B(B[0]), .Z(PRODUCT[93]) );
  AND U421 ( .A(A[92]), .B(B[0]), .Z(PRODUCT[92]) );
  AND U422 ( .A(A[91]), .B(B[0]), .Z(PRODUCT[91]) );
  AND U423 ( .A(A[90]), .B(B[0]), .Z(PRODUCT[90]) );
  AND U424 ( .A(A[89]), .B(B[0]), .Z(PRODUCT[89]) );
  AND U425 ( .A(A[88]), .B(B[0]), .Z(PRODUCT[88]) );
  AND U426 ( .A(A[87]), .B(B[0]), .Z(PRODUCT[87]) );
  AND U427 ( .A(A[86]), .B(B[0]), .Z(PRODUCT[86]) );
  AND U428 ( .A(A[85]), .B(B[0]), .Z(PRODUCT[85]) );
  AND U429 ( .A(A[84]), .B(B[0]), .Z(PRODUCT[84]) );
  AND U430 ( .A(A[83]), .B(B[0]), .Z(PRODUCT[83]) );
  AND U431 ( .A(A[82]), .B(B[0]), .Z(PRODUCT[82]) );
  AND U432 ( .A(A[81]), .B(B[0]), .Z(PRODUCT[81]) );
  AND U433 ( .A(A[80]), .B(B[0]), .Z(PRODUCT[80]) );
  AND U434 ( .A(A[79]), .B(B[0]), .Z(PRODUCT[79]) );
  AND U435 ( .A(A[78]), .B(B[0]), .Z(PRODUCT[78]) );
  AND U436 ( .A(A[77]), .B(B[0]), .Z(PRODUCT[77]) );
  AND U437 ( .A(A[76]), .B(B[0]), .Z(PRODUCT[76]) );
  AND U438 ( .A(A[75]), .B(B[0]), .Z(PRODUCT[75]) );
  AND U439 ( .A(A[74]), .B(B[0]), .Z(PRODUCT[74]) );
  AND U440 ( .A(A[73]), .B(B[0]), .Z(PRODUCT[73]) );
  AND U441 ( .A(A[72]), .B(B[0]), .Z(PRODUCT[72]) );
  AND U442 ( .A(A[71]), .B(B[0]), .Z(PRODUCT[71]) );
  AND U443 ( .A(A[70]), .B(B[0]), .Z(PRODUCT[70]) );
  AND U444 ( .A(A[69]), .B(B[0]), .Z(PRODUCT[69]) );
  AND U445 ( .A(A[68]), .B(B[0]), .Z(PRODUCT[68]) );
  AND U446 ( .A(A[67]), .B(B[0]), .Z(PRODUCT[67]) );
  AND U447 ( .A(A[66]), .B(B[0]), .Z(PRODUCT[66]) );
  AND U448 ( .A(A[65]), .B(B[0]), .Z(PRODUCT[65]) );
  AND U449 ( .A(A[64]), .B(B[0]), .Z(PRODUCT[64]) );
  AND U450 ( .A(A[63]), .B(B[0]), .Z(PRODUCT[63]) );
  AND U451 ( .A(A[62]), .B(B[0]), .Z(PRODUCT[62]) );
  AND U452 ( .A(A[61]), .B(B[0]), .Z(PRODUCT[61]) );
  AND U453 ( .A(A[60]), .B(B[0]), .Z(PRODUCT[60]) );
  AND U454 ( .A(A[59]), .B(B[0]), .Z(PRODUCT[59]) );
  AND U455 ( .A(A[58]), .B(B[0]), .Z(PRODUCT[58]) );
  AND U456 ( .A(A[57]), .B(B[0]), .Z(PRODUCT[57]) );
  AND U457 ( .A(A[56]), .B(B[0]), .Z(PRODUCT[56]) );
  AND U458 ( .A(A[55]), .B(B[0]), .Z(PRODUCT[55]) );
  AND U459 ( .A(A[54]), .B(B[0]), .Z(PRODUCT[54]) );
  AND U460 ( .A(A[53]), .B(B[0]), .Z(PRODUCT[53]) );
  AND U461 ( .A(A[52]), .B(B[0]), .Z(PRODUCT[52]) );
  AND U462 ( .A(A[51]), .B(B[0]), .Z(PRODUCT[51]) );
  AND U463 ( .A(A[50]), .B(B[0]), .Z(PRODUCT[50]) );
  AND U464 ( .A(A[49]), .B(B[0]), .Z(PRODUCT[49]) );
  AND U465 ( .A(A[48]), .B(B[0]), .Z(PRODUCT[48]) );
  AND U466 ( .A(A[47]), .B(B[0]), .Z(PRODUCT[47]) );
  AND U467 ( .A(A[46]), .B(B[0]), .Z(PRODUCT[46]) );
  AND U468 ( .A(A[45]), .B(B[0]), .Z(PRODUCT[45]) );
  AND U469 ( .A(A[44]), .B(B[0]), .Z(PRODUCT[44]) );
  AND U470 ( .A(A[43]), .B(B[0]), .Z(PRODUCT[43]) );
  AND U471 ( .A(A[42]), .B(B[0]), .Z(PRODUCT[42]) );
  AND U472 ( .A(A[41]), .B(B[0]), .Z(PRODUCT[41]) );
  AND U473 ( .A(A[40]), .B(B[0]), .Z(PRODUCT[40]) );
  AND U474 ( .A(A[39]), .B(B[0]), .Z(PRODUCT[39]) );
  AND U475 ( .A(A[38]), .B(B[0]), .Z(PRODUCT[38]) );
  AND U476 ( .A(A[37]), .B(B[0]), .Z(PRODUCT[37]) );
  AND U477 ( .A(A[36]), .B(B[0]), .Z(PRODUCT[36]) );
  AND U478 ( .A(A[35]), .B(B[0]), .Z(PRODUCT[35]) );
  AND U479 ( .A(A[34]), .B(B[0]), .Z(PRODUCT[34]) );
  AND U480 ( .A(A[33]), .B(B[0]), .Z(PRODUCT[33]) );
  AND U481 ( .A(A[32]), .B(B[0]), .Z(PRODUCT[32]) );
  AND U482 ( .A(A[31]), .B(B[0]), .Z(PRODUCT[31]) );
  AND U483 ( .A(A[30]), .B(B[0]), .Z(PRODUCT[30]) );
  AND U484 ( .A(A[29]), .B(B[0]), .Z(PRODUCT[29]) );
  AND U485 ( .A(A[28]), .B(B[0]), .Z(PRODUCT[28]) );
  AND U486 ( .A(A[27]), .B(B[0]), .Z(PRODUCT[27]) );
  AND U487 ( .A(A[26]), .B(B[0]), .Z(PRODUCT[26]) );
  AND U488 ( .A(A[25]), .B(B[0]), .Z(PRODUCT[25]) );
  AND U489 ( .A(A[24]), .B(B[0]), .Z(PRODUCT[24]) );
  AND U490 ( .A(A[23]), .B(B[0]), .Z(PRODUCT[23]) );
  AND U491 ( .A(A[22]), .B(B[0]), .Z(PRODUCT[22]) );
  AND U492 ( .A(A[21]), .B(B[0]), .Z(PRODUCT[21]) );
  AND U493 ( .A(A[20]), .B(B[0]), .Z(PRODUCT[20]) );
  AND U494 ( .A(A[19]), .B(B[0]), .Z(PRODUCT[19]) );
  AND U495 ( .A(A[18]), .B(B[0]), .Z(PRODUCT[18]) );
  AND U496 ( .A(A[17]), .B(B[0]), .Z(PRODUCT[17]) );
  AND U497 ( .A(A[16]), .B(B[0]), .Z(PRODUCT[16]) );
  AND U498 ( .A(A[15]), .B(B[0]), .Z(PRODUCT[15]) );
  AND U499 ( .A(A[14]), .B(B[0]), .Z(PRODUCT[14]) );
  AND U500 ( .A(A[13]), .B(B[0]), .Z(PRODUCT[13]) );
  AND U501 ( .A(A[12]), .B(B[0]), .Z(PRODUCT[12]) );
  AND U502 ( .A(A[11]), .B(B[0]), .Z(PRODUCT[11]) );
  AND U503 ( .A(A[10]), .B(B[0]), .Z(PRODUCT[10]) );
  AND U504 ( .A(B[0]), .B(A[9]), .Z(PRODUCT[9]) );
  AND U505 ( .A(A[8]), .B(B[0]), .Z(PRODUCT[8]) );
  AND U506 ( .A(A[7]), .B(B[0]), .Z(PRODUCT[7]) );
  AND U507 ( .A(A[6]), .B(B[0]), .Z(PRODUCT[6]) );
  AND U508 ( .A(A[5]), .B(B[0]), .Z(PRODUCT[5]) );
  AND U509 ( .A(A[4]), .B(B[0]), .Z(PRODUCT[4]) );
  AND U510 ( .A(A[3]), .B(B[0]), .Z(PRODUCT[3]) );
  AND U511 ( .A(A[2]), .B(B[0]), .Z(PRODUCT[2]) );
  AND U512 ( .A(A[1]), .B(B[0]), .Z(PRODUCT[1]) );
  AND U513 ( .A(A[0]), .B(B[0]), .Z(PRODUCT[0]) );
endmodule


module modmult_step_N512_DW01_cmp2_0 ( A, B, LEQ, TC, LT_LE, GE_GT );
  input [513:0] A;
  input [513:0] B;
  input LEQ, TC;
  output LT_LE, GE_GT;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046;

  NAND U1 ( .A(n1), .B(n2), .Z(LT_LE) );
  NOR U2 ( .A(B[513]), .B(B[512]), .Z(n2) );
  AND U3 ( .A(n3), .B(n4), .Z(n1) );
  NAND U4 ( .A(n5), .B(n6), .Z(n4) );
  NANDN U5 ( .A(B[511]), .B(A[511]), .Z(n6) );
  NAND U6 ( .A(n7), .B(n8), .Z(n5) );
  NANDN U7 ( .A(A[510]), .B(B[510]), .Z(n8) );
  NAND U8 ( .A(n9), .B(n10), .Z(n7) );
  NANDN U9 ( .A(B[510]), .B(A[510]), .Z(n10) );
  AND U10 ( .A(n11), .B(n12), .Z(n9) );
  NAND U11 ( .A(n13), .B(n14), .Z(n12) );
  NANDN U12 ( .A(A[509]), .B(B[509]), .Z(n14) );
  AND U13 ( .A(n15), .B(n16), .Z(n13) );
  NANDN U14 ( .A(A[508]), .B(B[508]), .Z(n16) );
  NAND U15 ( .A(n17), .B(n18), .Z(n15) );
  NANDN U16 ( .A(B[508]), .B(A[508]), .Z(n18) );
  AND U17 ( .A(n19), .B(n20), .Z(n17) );
  NAND U18 ( .A(n21), .B(n22), .Z(n20) );
  NANDN U19 ( .A(A[507]), .B(B[507]), .Z(n22) );
  AND U20 ( .A(n23), .B(n24), .Z(n21) );
  NANDN U21 ( .A(A[506]), .B(B[506]), .Z(n24) );
  NAND U22 ( .A(n25), .B(n26), .Z(n23) );
  NANDN U23 ( .A(B[506]), .B(A[506]), .Z(n26) );
  AND U24 ( .A(n27), .B(n28), .Z(n25) );
  NAND U25 ( .A(n29), .B(n30), .Z(n28) );
  NANDN U26 ( .A(A[505]), .B(B[505]), .Z(n30) );
  AND U27 ( .A(n31), .B(n32), .Z(n29) );
  NANDN U28 ( .A(A[504]), .B(B[504]), .Z(n32) );
  NAND U29 ( .A(n33), .B(n34), .Z(n31) );
  NANDN U30 ( .A(B[504]), .B(A[504]), .Z(n34) );
  AND U31 ( .A(n35), .B(n36), .Z(n33) );
  NAND U32 ( .A(n37), .B(n38), .Z(n36) );
  NANDN U33 ( .A(A[503]), .B(B[503]), .Z(n38) );
  AND U34 ( .A(n39), .B(n40), .Z(n37) );
  NANDN U35 ( .A(A[502]), .B(B[502]), .Z(n40) );
  NAND U36 ( .A(n41), .B(n42), .Z(n39) );
  NANDN U37 ( .A(B[502]), .B(A[502]), .Z(n42) );
  AND U38 ( .A(n43), .B(n44), .Z(n41) );
  NAND U39 ( .A(n45), .B(n46), .Z(n44) );
  NANDN U40 ( .A(A[501]), .B(B[501]), .Z(n46) );
  AND U41 ( .A(n47), .B(n48), .Z(n45) );
  NANDN U42 ( .A(A[500]), .B(B[500]), .Z(n48) );
  NAND U43 ( .A(n49), .B(n50), .Z(n47) );
  NANDN U44 ( .A(B[500]), .B(A[500]), .Z(n50) );
  AND U45 ( .A(n51), .B(n52), .Z(n49) );
  NAND U46 ( .A(n53), .B(n54), .Z(n52) );
  NANDN U47 ( .A(A[499]), .B(B[499]), .Z(n54) );
  AND U48 ( .A(n55), .B(n56), .Z(n53) );
  NANDN U49 ( .A(A[498]), .B(B[498]), .Z(n56) );
  NAND U50 ( .A(n57), .B(n58), .Z(n55) );
  NANDN U51 ( .A(B[498]), .B(A[498]), .Z(n58) );
  AND U52 ( .A(n59), .B(n60), .Z(n57) );
  NAND U53 ( .A(n61), .B(n62), .Z(n60) );
  NANDN U54 ( .A(A[497]), .B(B[497]), .Z(n62) );
  AND U55 ( .A(n63), .B(n64), .Z(n61) );
  NANDN U56 ( .A(A[496]), .B(B[496]), .Z(n64) );
  NAND U57 ( .A(n65), .B(n66), .Z(n63) );
  NANDN U58 ( .A(B[496]), .B(A[496]), .Z(n66) );
  AND U59 ( .A(n67), .B(n68), .Z(n65) );
  NAND U60 ( .A(n69), .B(n70), .Z(n68) );
  NANDN U61 ( .A(A[495]), .B(B[495]), .Z(n70) );
  AND U62 ( .A(n71), .B(n72), .Z(n69) );
  NANDN U63 ( .A(A[494]), .B(B[494]), .Z(n72) );
  NAND U64 ( .A(n73), .B(n74), .Z(n71) );
  NANDN U65 ( .A(B[494]), .B(A[494]), .Z(n74) );
  AND U66 ( .A(n75), .B(n76), .Z(n73) );
  NAND U67 ( .A(n77), .B(n78), .Z(n76) );
  NANDN U68 ( .A(A[493]), .B(B[493]), .Z(n78) );
  AND U69 ( .A(n79), .B(n80), .Z(n77) );
  NANDN U70 ( .A(A[492]), .B(B[492]), .Z(n80) );
  NAND U71 ( .A(n81), .B(n82), .Z(n79) );
  NANDN U72 ( .A(B[492]), .B(A[492]), .Z(n82) );
  AND U73 ( .A(n83), .B(n84), .Z(n81) );
  NAND U74 ( .A(n85), .B(n86), .Z(n84) );
  NANDN U75 ( .A(A[491]), .B(B[491]), .Z(n86) );
  AND U76 ( .A(n87), .B(n88), .Z(n85) );
  NANDN U77 ( .A(A[490]), .B(B[490]), .Z(n88) );
  NAND U78 ( .A(n89), .B(n90), .Z(n87) );
  NANDN U79 ( .A(B[490]), .B(A[490]), .Z(n90) );
  AND U80 ( .A(n91), .B(n92), .Z(n89) );
  NAND U81 ( .A(n93), .B(n94), .Z(n92) );
  NANDN U82 ( .A(A[489]), .B(B[489]), .Z(n94) );
  AND U83 ( .A(n95), .B(n96), .Z(n93) );
  NANDN U84 ( .A(A[488]), .B(B[488]), .Z(n96) );
  NAND U85 ( .A(n97), .B(n98), .Z(n95) );
  NANDN U86 ( .A(B[488]), .B(A[488]), .Z(n98) );
  AND U87 ( .A(n99), .B(n100), .Z(n97) );
  NAND U88 ( .A(n101), .B(n102), .Z(n100) );
  NANDN U89 ( .A(A[487]), .B(B[487]), .Z(n102) );
  AND U90 ( .A(n103), .B(n104), .Z(n101) );
  NANDN U91 ( .A(A[486]), .B(B[486]), .Z(n104) );
  NAND U92 ( .A(n105), .B(n106), .Z(n103) );
  NANDN U93 ( .A(B[486]), .B(A[486]), .Z(n106) );
  AND U94 ( .A(n107), .B(n108), .Z(n105) );
  NAND U95 ( .A(n109), .B(n110), .Z(n108) );
  NANDN U96 ( .A(A[485]), .B(B[485]), .Z(n110) );
  AND U97 ( .A(n111), .B(n112), .Z(n109) );
  NANDN U98 ( .A(A[484]), .B(B[484]), .Z(n112) );
  NAND U99 ( .A(n113), .B(n114), .Z(n111) );
  NANDN U100 ( .A(B[484]), .B(A[484]), .Z(n114) );
  AND U101 ( .A(n115), .B(n116), .Z(n113) );
  NAND U102 ( .A(n117), .B(n118), .Z(n116) );
  NANDN U103 ( .A(A[483]), .B(B[483]), .Z(n118) );
  AND U104 ( .A(n119), .B(n120), .Z(n117) );
  NANDN U105 ( .A(A[482]), .B(B[482]), .Z(n120) );
  NAND U106 ( .A(n121), .B(n122), .Z(n119) );
  NANDN U107 ( .A(B[482]), .B(A[482]), .Z(n122) );
  AND U108 ( .A(n123), .B(n124), .Z(n121) );
  NAND U109 ( .A(n125), .B(n126), .Z(n124) );
  NANDN U110 ( .A(A[481]), .B(B[481]), .Z(n126) );
  AND U111 ( .A(n127), .B(n128), .Z(n125) );
  NANDN U112 ( .A(A[480]), .B(B[480]), .Z(n128) );
  NAND U113 ( .A(n129), .B(n130), .Z(n127) );
  NANDN U114 ( .A(B[480]), .B(A[480]), .Z(n130) );
  AND U115 ( .A(n131), .B(n132), .Z(n129) );
  NAND U116 ( .A(n133), .B(n134), .Z(n132) );
  NANDN U117 ( .A(A[479]), .B(B[479]), .Z(n134) );
  AND U118 ( .A(n135), .B(n136), .Z(n133) );
  NANDN U119 ( .A(A[478]), .B(B[478]), .Z(n136) );
  NAND U120 ( .A(n137), .B(n138), .Z(n135) );
  NANDN U121 ( .A(B[478]), .B(A[478]), .Z(n138) );
  AND U122 ( .A(n139), .B(n140), .Z(n137) );
  NAND U123 ( .A(n141), .B(n142), .Z(n140) );
  NANDN U124 ( .A(A[477]), .B(B[477]), .Z(n142) );
  AND U125 ( .A(n143), .B(n144), .Z(n141) );
  NANDN U126 ( .A(A[476]), .B(B[476]), .Z(n144) );
  NAND U127 ( .A(n145), .B(n146), .Z(n143) );
  NANDN U128 ( .A(B[476]), .B(A[476]), .Z(n146) );
  AND U129 ( .A(n147), .B(n148), .Z(n145) );
  NAND U130 ( .A(n149), .B(n150), .Z(n148) );
  NANDN U131 ( .A(A[475]), .B(B[475]), .Z(n150) );
  AND U132 ( .A(n151), .B(n152), .Z(n149) );
  NANDN U133 ( .A(A[474]), .B(B[474]), .Z(n152) );
  NAND U134 ( .A(n153), .B(n154), .Z(n151) );
  NANDN U135 ( .A(B[474]), .B(A[474]), .Z(n154) );
  AND U136 ( .A(n155), .B(n156), .Z(n153) );
  NAND U137 ( .A(n157), .B(n158), .Z(n156) );
  NANDN U138 ( .A(A[473]), .B(B[473]), .Z(n158) );
  AND U139 ( .A(n159), .B(n160), .Z(n157) );
  NANDN U140 ( .A(A[472]), .B(B[472]), .Z(n160) );
  NAND U141 ( .A(n161), .B(n162), .Z(n159) );
  NANDN U142 ( .A(B[472]), .B(A[472]), .Z(n162) );
  AND U143 ( .A(n163), .B(n164), .Z(n161) );
  NAND U144 ( .A(n165), .B(n166), .Z(n164) );
  NANDN U145 ( .A(A[471]), .B(B[471]), .Z(n166) );
  AND U146 ( .A(n167), .B(n168), .Z(n165) );
  NANDN U147 ( .A(A[470]), .B(B[470]), .Z(n168) );
  NAND U148 ( .A(n169), .B(n170), .Z(n167) );
  NANDN U149 ( .A(B[470]), .B(A[470]), .Z(n170) );
  AND U150 ( .A(n171), .B(n172), .Z(n169) );
  NAND U151 ( .A(n173), .B(n174), .Z(n172) );
  NANDN U152 ( .A(A[469]), .B(B[469]), .Z(n174) );
  AND U153 ( .A(n175), .B(n176), .Z(n173) );
  NANDN U154 ( .A(A[468]), .B(B[468]), .Z(n176) );
  NAND U155 ( .A(n177), .B(n178), .Z(n175) );
  NANDN U156 ( .A(B[468]), .B(A[468]), .Z(n178) );
  AND U157 ( .A(n179), .B(n180), .Z(n177) );
  NAND U158 ( .A(n181), .B(n182), .Z(n180) );
  NANDN U159 ( .A(A[467]), .B(B[467]), .Z(n182) );
  AND U160 ( .A(n183), .B(n184), .Z(n181) );
  NANDN U161 ( .A(A[466]), .B(B[466]), .Z(n184) );
  NAND U162 ( .A(n185), .B(n186), .Z(n183) );
  NANDN U163 ( .A(B[466]), .B(A[466]), .Z(n186) );
  AND U164 ( .A(n187), .B(n188), .Z(n185) );
  NAND U165 ( .A(n189), .B(n190), .Z(n188) );
  NANDN U166 ( .A(A[465]), .B(B[465]), .Z(n190) );
  AND U167 ( .A(n191), .B(n192), .Z(n189) );
  NANDN U168 ( .A(A[464]), .B(B[464]), .Z(n192) );
  NAND U169 ( .A(n193), .B(n194), .Z(n191) );
  NANDN U170 ( .A(B[464]), .B(A[464]), .Z(n194) );
  AND U171 ( .A(n195), .B(n196), .Z(n193) );
  NAND U172 ( .A(n197), .B(n198), .Z(n196) );
  NANDN U173 ( .A(A[463]), .B(B[463]), .Z(n198) );
  AND U174 ( .A(n199), .B(n200), .Z(n197) );
  NANDN U175 ( .A(A[462]), .B(B[462]), .Z(n200) );
  NAND U176 ( .A(n201), .B(n202), .Z(n199) );
  NANDN U177 ( .A(B[462]), .B(A[462]), .Z(n202) );
  AND U178 ( .A(n203), .B(n204), .Z(n201) );
  NAND U179 ( .A(n205), .B(n206), .Z(n204) );
  NANDN U180 ( .A(A[461]), .B(B[461]), .Z(n206) );
  AND U181 ( .A(n207), .B(n208), .Z(n205) );
  NANDN U182 ( .A(A[460]), .B(B[460]), .Z(n208) );
  NAND U183 ( .A(n209), .B(n210), .Z(n207) );
  NANDN U184 ( .A(B[460]), .B(A[460]), .Z(n210) );
  AND U185 ( .A(n211), .B(n212), .Z(n209) );
  NAND U186 ( .A(n213), .B(n214), .Z(n212) );
  NANDN U187 ( .A(A[459]), .B(B[459]), .Z(n214) );
  AND U188 ( .A(n215), .B(n216), .Z(n213) );
  NANDN U189 ( .A(A[458]), .B(B[458]), .Z(n216) );
  NAND U190 ( .A(n217), .B(n218), .Z(n215) );
  NANDN U191 ( .A(B[458]), .B(A[458]), .Z(n218) );
  AND U192 ( .A(n219), .B(n220), .Z(n217) );
  NAND U193 ( .A(n221), .B(n222), .Z(n220) );
  NANDN U194 ( .A(A[457]), .B(B[457]), .Z(n222) );
  AND U195 ( .A(n223), .B(n224), .Z(n221) );
  NANDN U196 ( .A(A[456]), .B(B[456]), .Z(n224) );
  NAND U197 ( .A(n225), .B(n226), .Z(n223) );
  NANDN U198 ( .A(B[456]), .B(A[456]), .Z(n226) );
  AND U199 ( .A(n227), .B(n228), .Z(n225) );
  NAND U200 ( .A(n229), .B(n230), .Z(n228) );
  NANDN U201 ( .A(A[455]), .B(B[455]), .Z(n230) );
  AND U202 ( .A(n231), .B(n232), .Z(n229) );
  NANDN U203 ( .A(A[454]), .B(B[454]), .Z(n232) );
  NAND U204 ( .A(n233), .B(n234), .Z(n231) );
  NANDN U205 ( .A(B[454]), .B(A[454]), .Z(n234) );
  AND U206 ( .A(n235), .B(n236), .Z(n233) );
  NAND U207 ( .A(n237), .B(n238), .Z(n236) );
  NANDN U208 ( .A(A[453]), .B(B[453]), .Z(n238) );
  AND U209 ( .A(n239), .B(n240), .Z(n237) );
  NANDN U210 ( .A(A[452]), .B(B[452]), .Z(n240) );
  NAND U211 ( .A(n241), .B(n242), .Z(n239) );
  NANDN U212 ( .A(B[452]), .B(A[452]), .Z(n242) );
  AND U213 ( .A(n243), .B(n244), .Z(n241) );
  NAND U214 ( .A(n245), .B(n246), .Z(n244) );
  NANDN U215 ( .A(A[451]), .B(B[451]), .Z(n246) );
  AND U216 ( .A(n247), .B(n248), .Z(n245) );
  NANDN U217 ( .A(A[450]), .B(B[450]), .Z(n248) );
  NAND U218 ( .A(n249), .B(n250), .Z(n247) );
  NANDN U219 ( .A(B[450]), .B(A[450]), .Z(n250) );
  AND U220 ( .A(n251), .B(n252), .Z(n249) );
  NAND U221 ( .A(n253), .B(n254), .Z(n252) );
  NANDN U222 ( .A(A[449]), .B(B[449]), .Z(n254) );
  AND U223 ( .A(n255), .B(n256), .Z(n253) );
  NANDN U224 ( .A(A[448]), .B(B[448]), .Z(n256) );
  NAND U225 ( .A(n257), .B(n258), .Z(n255) );
  NANDN U226 ( .A(B[448]), .B(A[448]), .Z(n258) );
  AND U227 ( .A(n259), .B(n260), .Z(n257) );
  NAND U228 ( .A(n261), .B(n262), .Z(n260) );
  NANDN U229 ( .A(A[447]), .B(B[447]), .Z(n262) );
  AND U230 ( .A(n263), .B(n264), .Z(n261) );
  NANDN U231 ( .A(A[446]), .B(B[446]), .Z(n264) );
  NAND U232 ( .A(n265), .B(n266), .Z(n263) );
  NANDN U233 ( .A(B[446]), .B(A[446]), .Z(n266) );
  AND U234 ( .A(n267), .B(n268), .Z(n265) );
  NAND U235 ( .A(n269), .B(n270), .Z(n268) );
  NANDN U236 ( .A(A[445]), .B(B[445]), .Z(n270) );
  AND U237 ( .A(n271), .B(n272), .Z(n269) );
  NANDN U238 ( .A(A[444]), .B(B[444]), .Z(n272) );
  NAND U239 ( .A(n273), .B(n274), .Z(n271) );
  NANDN U240 ( .A(B[444]), .B(A[444]), .Z(n274) );
  AND U241 ( .A(n275), .B(n276), .Z(n273) );
  NAND U242 ( .A(n277), .B(n278), .Z(n276) );
  NANDN U243 ( .A(A[443]), .B(B[443]), .Z(n278) );
  AND U244 ( .A(n279), .B(n280), .Z(n277) );
  NANDN U245 ( .A(A[442]), .B(B[442]), .Z(n280) );
  NAND U246 ( .A(n281), .B(n282), .Z(n279) );
  NANDN U247 ( .A(B[442]), .B(A[442]), .Z(n282) );
  AND U248 ( .A(n283), .B(n284), .Z(n281) );
  NAND U249 ( .A(n285), .B(n286), .Z(n284) );
  NANDN U250 ( .A(A[441]), .B(B[441]), .Z(n286) );
  AND U251 ( .A(n287), .B(n288), .Z(n285) );
  NANDN U252 ( .A(A[440]), .B(B[440]), .Z(n288) );
  NAND U253 ( .A(n289), .B(n290), .Z(n287) );
  NANDN U254 ( .A(B[440]), .B(A[440]), .Z(n290) );
  AND U255 ( .A(n291), .B(n292), .Z(n289) );
  NAND U256 ( .A(n293), .B(n294), .Z(n292) );
  NANDN U257 ( .A(A[439]), .B(B[439]), .Z(n294) );
  AND U258 ( .A(n295), .B(n296), .Z(n293) );
  NANDN U259 ( .A(A[438]), .B(B[438]), .Z(n296) );
  NAND U260 ( .A(n297), .B(n298), .Z(n295) );
  NANDN U261 ( .A(B[438]), .B(A[438]), .Z(n298) );
  AND U262 ( .A(n299), .B(n300), .Z(n297) );
  NAND U263 ( .A(n301), .B(n302), .Z(n300) );
  NANDN U264 ( .A(A[437]), .B(B[437]), .Z(n302) );
  AND U265 ( .A(n303), .B(n304), .Z(n301) );
  NANDN U266 ( .A(A[436]), .B(B[436]), .Z(n304) );
  NAND U267 ( .A(n305), .B(n306), .Z(n303) );
  NANDN U268 ( .A(B[436]), .B(A[436]), .Z(n306) );
  AND U269 ( .A(n307), .B(n308), .Z(n305) );
  NAND U270 ( .A(n309), .B(n310), .Z(n308) );
  NANDN U271 ( .A(A[435]), .B(B[435]), .Z(n310) );
  AND U272 ( .A(n311), .B(n312), .Z(n309) );
  NANDN U273 ( .A(A[434]), .B(B[434]), .Z(n312) );
  NAND U274 ( .A(n313), .B(n314), .Z(n311) );
  NANDN U275 ( .A(B[434]), .B(A[434]), .Z(n314) );
  AND U276 ( .A(n315), .B(n316), .Z(n313) );
  NAND U277 ( .A(n317), .B(n318), .Z(n316) );
  NANDN U278 ( .A(A[433]), .B(B[433]), .Z(n318) );
  AND U279 ( .A(n319), .B(n320), .Z(n317) );
  NANDN U280 ( .A(A[432]), .B(B[432]), .Z(n320) );
  NAND U281 ( .A(n321), .B(n322), .Z(n319) );
  NANDN U282 ( .A(B[432]), .B(A[432]), .Z(n322) );
  AND U283 ( .A(n323), .B(n324), .Z(n321) );
  NAND U284 ( .A(n325), .B(n326), .Z(n324) );
  NANDN U285 ( .A(A[431]), .B(B[431]), .Z(n326) );
  AND U286 ( .A(n327), .B(n328), .Z(n325) );
  NANDN U287 ( .A(A[430]), .B(B[430]), .Z(n328) );
  NAND U288 ( .A(n329), .B(n330), .Z(n327) );
  NANDN U289 ( .A(B[430]), .B(A[430]), .Z(n330) );
  AND U290 ( .A(n331), .B(n332), .Z(n329) );
  NAND U291 ( .A(n333), .B(n334), .Z(n332) );
  NANDN U292 ( .A(A[429]), .B(B[429]), .Z(n334) );
  AND U293 ( .A(n335), .B(n336), .Z(n333) );
  NANDN U294 ( .A(A[428]), .B(B[428]), .Z(n336) );
  NAND U295 ( .A(n337), .B(n338), .Z(n335) );
  NANDN U296 ( .A(B[428]), .B(A[428]), .Z(n338) );
  AND U297 ( .A(n339), .B(n340), .Z(n337) );
  NAND U298 ( .A(n341), .B(n342), .Z(n340) );
  NANDN U299 ( .A(A[427]), .B(B[427]), .Z(n342) );
  AND U300 ( .A(n343), .B(n344), .Z(n341) );
  NANDN U301 ( .A(A[426]), .B(B[426]), .Z(n344) );
  NAND U302 ( .A(n345), .B(n346), .Z(n343) );
  NANDN U303 ( .A(B[426]), .B(A[426]), .Z(n346) );
  AND U304 ( .A(n347), .B(n348), .Z(n345) );
  NAND U305 ( .A(n349), .B(n350), .Z(n348) );
  NANDN U306 ( .A(A[425]), .B(B[425]), .Z(n350) );
  AND U307 ( .A(n351), .B(n352), .Z(n349) );
  NANDN U308 ( .A(A[424]), .B(B[424]), .Z(n352) );
  NAND U309 ( .A(n353), .B(n354), .Z(n351) );
  NANDN U310 ( .A(B[424]), .B(A[424]), .Z(n354) );
  AND U311 ( .A(n355), .B(n356), .Z(n353) );
  NAND U312 ( .A(n357), .B(n358), .Z(n356) );
  NANDN U313 ( .A(A[423]), .B(B[423]), .Z(n358) );
  AND U314 ( .A(n359), .B(n360), .Z(n357) );
  NANDN U315 ( .A(A[422]), .B(B[422]), .Z(n360) );
  NAND U316 ( .A(n361), .B(n362), .Z(n359) );
  NANDN U317 ( .A(B[422]), .B(A[422]), .Z(n362) );
  AND U318 ( .A(n363), .B(n364), .Z(n361) );
  NAND U319 ( .A(n365), .B(n366), .Z(n364) );
  NANDN U320 ( .A(A[421]), .B(B[421]), .Z(n366) );
  AND U321 ( .A(n367), .B(n368), .Z(n365) );
  NANDN U322 ( .A(A[420]), .B(B[420]), .Z(n368) );
  NAND U323 ( .A(n369), .B(n370), .Z(n367) );
  NANDN U324 ( .A(B[420]), .B(A[420]), .Z(n370) );
  AND U325 ( .A(n371), .B(n372), .Z(n369) );
  NAND U326 ( .A(n373), .B(n374), .Z(n372) );
  NANDN U327 ( .A(A[419]), .B(B[419]), .Z(n374) );
  AND U328 ( .A(n375), .B(n376), .Z(n373) );
  NANDN U329 ( .A(A[418]), .B(B[418]), .Z(n376) );
  NAND U330 ( .A(n377), .B(n378), .Z(n375) );
  NANDN U331 ( .A(B[418]), .B(A[418]), .Z(n378) );
  AND U332 ( .A(n379), .B(n380), .Z(n377) );
  NAND U333 ( .A(n381), .B(n382), .Z(n380) );
  NANDN U334 ( .A(A[417]), .B(B[417]), .Z(n382) );
  AND U335 ( .A(n383), .B(n384), .Z(n381) );
  NANDN U336 ( .A(A[416]), .B(B[416]), .Z(n384) );
  NAND U337 ( .A(n385), .B(n386), .Z(n383) );
  NANDN U338 ( .A(B[416]), .B(A[416]), .Z(n386) );
  AND U339 ( .A(n387), .B(n388), .Z(n385) );
  NAND U340 ( .A(n389), .B(n390), .Z(n388) );
  NANDN U341 ( .A(A[415]), .B(B[415]), .Z(n390) );
  AND U342 ( .A(n391), .B(n392), .Z(n389) );
  NANDN U343 ( .A(A[414]), .B(B[414]), .Z(n392) );
  NAND U344 ( .A(n393), .B(n394), .Z(n391) );
  NANDN U345 ( .A(B[414]), .B(A[414]), .Z(n394) );
  AND U346 ( .A(n395), .B(n396), .Z(n393) );
  NAND U347 ( .A(n397), .B(n398), .Z(n396) );
  NANDN U348 ( .A(A[413]), .B(B[413]), .Z(n398) );
  AND U349 ( .A(n399), .B(n400), .Z(n397) );
  NANDN U350 ( .A(A[412]), .B(B[412]), .Z(n400) );
  NAND U351 ( .A(n401), .B(n402), .Z(n399) );
  NANDN U352 ( .A(B[412]), .B(A[412]), .Z(n402) );
  AND U353 ( .A(n403), .B(n404), .Z(n401) );
  NAND U354 ( .A(n405), .B(n406), .Z(n404) );
  NANDN U355 ( .A(A[411]), .B(B[411]), .Z(n406) );
  AND U356 ( .A(n407), .B(n408), .Z(n405) );
  NANDN U357 ( .A(A[410]), .B(B[410]), .Z(n408) );
  NAND U358 ( .A(n409), .B(n410), .Z(n407) );
  NANDN U359 ( .A(B[410]), .B(A[410]), .Z(n410) );
  AND U360 ( .A(n411), .B(n412), .Z(n409) );
  NAND U361 ( .A(n413), .B(n414), .Z(n412) );
  NANDN U362 ( .A(A[409]), .B(B[409]), .Z(n414) );
  AND U363 ( .A(n415), .B(n416), .Z(n413) );
  NANDN U364 ( .A(A[408]), .B(B[408]), .Z(n416) );
  NAND U365 ( .A(n417), .B(n418), .Z(n415) );
  NANDN U366 ( .A(B[408]), .B(A[408]), .Z(n418) );
  AND U367 ( .A(n419), .B(n420), .Z(n417) );
  NAND U368 ( .A(n421), .B(n422), .Z(n420) );
  NANDN U369 ( .A(A[407]), .B(B[407]), .Z(n422) );
  AND U370 ( .A(n423), .B(n424), .Z(n421) );
  NANDN U371 ( .A(A[406]), .B(B[406]), .Z(n424) );
  NAND U372 ( .A(n425), .B(n426), .Z(n423) );
  NANDN U373 ( .A(B[406]), .B(A[406]), .Z(n426) );
  AND U374 ( .A(n427), .B(n428), .Z(n425) );
  NAND U375 ( .A(n429), .B(n430), .Z(n428) );
  NANDN U376 ( .A(A[405]), .B(B[405]), .Z(n430) );
  AND U377 ( .A(n431), .B(n432), .Z(n429) );
  NANDN U378 ( .A(A[404]), .B(B[404]), .Z(n432) );
  NAND U379 ( .A(n433), .B(n434), .Z(n431) );
  NANDN U380 ( .A(B[404]), .B(A[404]), .Z(n434) );
  AND U381 ( .A(n435), .B(n436), .Z(n433) );
  NAND U382 ( .A(n437), .B(n438), .Z(n436) );
  NANDN U383 ( .A(A[403]), .B(B[403]), .Z(n438) );
  AND U384 ( .A(n439), .B(n440), .Z(n437) );
  NANDN U385 ( .A(A[402]), .B(B[402]), .Z(n440) );
  NAND U386 ( .A(n441), .B(n442), .Z(n439) );
  NANDN U387 ( .A(B[402]), .B(A[402]), .Z(n442) );
  AND U388 ( .A(n443), .B(n444), .Z(n441) );
  NAND U389 ( .A(n445), .B(n446), .Z(n444) );
  NANDN U390 ( .A(A[401]), .B(B[401]), .Z(n446) );
  AND U391 ( .A(n447), .B(n448), .Z(n445) );
  NANDN U392 ( .A(A[400]), .B(B[400]), .Z(n448) );
  NAND U393 ( .A(n449), .B(n450), .Z(n447) );
  NANDN U394 ( .A(B[400]), .B(A[400]), .Z(n450) );
  AND U395 ( .A(n451), .B(n452), .Z(n449) );
  NAND U396 ( .A(n453), .B(n454), .Z(n452) );
  NANDN U397 ( .A(A[399]), .B(B[399]), .Z(n454) );
  AND U398 ( .A(n455), .B(n456), .Z(n453) );
  NANDN U399 ( .A(A[398]), .B(B[398]), .Z(n456) );
  NAND U400 ( .A(n457), .B(n458), .Z(n455) );
  NANDN U401 ( .A(B[398]), .B(A[398]), .Z(n458) );
  AND U402 ( .A(n459), .B(n460), .Z(n457) );
  NAND U403 ( .A(n461), .B(n462), .Z(n460) );
  NANDN U404 ( .A(A[397]), .B(B[397]), .Z(n462) );
  AND U405 ( .A(n463), .B(n464), .Z(n461) );
  NANDN U406 ( .A(A[396]), .B(B[396]), .Z(n464) );
  NAND U407 ( .A(n465), .B(n466), .Z(n463) );
  NANDN U408 ( .A(B[396]), .B(A[396]), .Z(n466) );
  AND U409 ( .A(n467), .B(n468), .Z(n465) );
  NAND U410 ( .A(n469), .B(n470), .Z(n468) );
  NANDN U411 ( .A(A[395]), .B(B[395]), .Z(n470) );
  AND U412 ( .A(n471), .B(n472), .Z(n469) );
  NANDN U413 ( .A(A[394]), .B(B[394]), .Z(n472) );
  NAND U414 ( .A(n473), .B(n474), .Z(n471) );
  NANDN U415 ( .A(B[394]), .B(A[394]), .Z(n474) );
  AND U416 ( .A(n475), .B(n476), .Z(n473) );
  NAND U417 ( .A(n477), .B(n478), .Z(n476) );
  NANDN U418 ( .A(A[393]), .B(B[393]), .Z(n478) );
  AND U419 ( .A(n479), .B(n480), .Z(n477) );
  NANDN U420 ( .A(A[392]), .B(B[392]), .Z(n480) );
  NAND U421 ( .A(n481), .B(n482), .Z(n479) );
  NANDN U422 ( .A(B[392]), .B(A[392]), .Z(n482) );
  AND U423 ( .A(n483), .B(n484), .Z(n481) );
  NAND U424 ( .A(n485), .B(n486), .Z(n484) );
  NANDN U425 ( .A(A[391]), .B(B[391]), .Z(n486) );
  AND U426 ( .A(n487), .B(n488), .Z(n485) );
  NANDN U427 ( .A(A[390]), .B(B[390]), .Z(n488) );
  NAND U428 ( .A(n489), .B(n490), .Z(n487) );
  NANDN U429 ( .A(B[390]), .B(A[390]), .Z(n490) );
  AND U430 ( .A(n491), .B(n492), .Z(n489) );
  NAND U431 ( .A(n493), .B(n494), .Z(n492) );
  NANDN U432 ( .A(A[389]), .B(B[389]), .Z(n494) );
  AND U433 ( .A(n495), .B(n496), .Z(n493) );
  NANDN U434 ( .A(A[388]), .B(B[388]), .Z(n496) );
  NAND U435 ( .A(n497), .B(n498), .Z(n495) );
  NANDN U436 ( .A(B[388]), .B(A[388]), .Z(n498) );
  AND U437 ( .A(n499), .B(n500), .Z(n497) );
  NAND U438 ( .A(n501), .B(n502), .Z(n500) );
  NANDN U439 ( .A(A[387]), .B(B[387]), .Z(n502) );
  AND U440 ( .A(n503), .B(n504), .Z(n501) );
  NANDN U441 ( .A(A[386]), .B(B[386]), .Z(n504) );
  NAND U442 ( .A(n505), .B(n506), .Z(n503) );
  NANDN U443 ( .A(B[386]), .B(A[386]), .Z(n506) );
  AND U444 ( .A(n507), .B(n508), .Z(n505) );
  NAND U445 ( .A(n509), .B(n510), .Z(n508) );
  NANDN U446 ( .A(A[385]), .B(B[385]), .Z(n510) );
  AND U447 ( .A(n511), .B(n512), .Z(n509) );
  NANDN U448 ( .A(A[384]), .B(B[384]), .Z(n512) );
  NAND U449 ( .A(n513), .B(n514), .Z(n511) );
  NANDN U450 ( .A(B[384]), .B(A[384]), .Z(n514) );
  AND U451 ( .A(n515), .B(n516), .Z(n513) );
  NAND U452 ( .A(n517), .B(n518), .Z(n516) );
  NANDN U453 ( .A(A[383]), .B(B[383]), .Z(n518) );
  AND U454 ( .A(n519), .B(n520), .Z(n517) );
  NANDN U455 ( .A(A[382]), .B(B[382]), .Z(n520) );
  NAND U456 ( .A(n521), .B(n522), .Z(n519) );
  NANDN U457 ( .A(B[382]), .B(A[382]), .Z(n522) );
  AND U458 ( .A(n523), .B(n524), .Z(n521) );
  NAND U459 ( .A(n525), .B(n526), .Z(n524) );
  NANDN U460 ( .A(A[381]), .B(B[381]), .Z(n526) );
  AND U461 ( .A(n527), .B(n528), .Z(n525) );
  NANDN U462 ( .A(A[380]), .B(B[380]), .Z(n528) );
  NAND U463 ( .A(n529), .B(n530), .Z(n527) );
  NANDN U464 ( .A(B[380]), .B(A[380]), .Z(n530) );
  AND U465 ( .A(n531), .B(n532), .Z(n529) );
  NAND U466 ( .A(n533), .B(n534), .Z(n532) );
  NANDN U467 ( .A(A[379]), .B(B[379]), .Z(n534) );
  AND U468 ( .A(n535), .B(n536), .Z(n533) );
  NANDN U469 ( .A(A[378]), .B(B[378]), .Z(n536) );
  NAND U470 ( .A(n537), .B(n538), .Z(n535) );
  NANDN U471 ( .A(B[378]), .B(A[378]), .Z(n538) );
  AND U472 ( .A(n539), .B(n540), .Z(n537) );
  NAND U473 ( .A(n541), .B(n542), .Z(n540) );
  NANDN U474 ( .A(A[377]), .B(B[377]), .Z(n542) );
  AND U475 ( .A(n543), .B(n544), .Z(n541) );
  NANDN U476 ( .A(A[376]), .B(B[376]), .Z(n544) );
  NAND U477 ( .A(n545), .B(n546), .Z(n543) );
  NANDN U478 ( .A(B[376]), .B(A[376]), .Z(n546) );
  AND U479 ( .A(n547), .B(n548), .Z(n545) );
  NAND U480 ( .A(n549), .B(n550), .Z(n548) );
  NANDN U481 ( .A(A[375]), .B(B[375]), .Z(n550) );
  AND U482 ( .A(n551), .B(n552), .Z(n549) );
  NANDN U483 ( .A(A[374]), .B(B[374]), .Z(n552) );
  NAND U484 ( .A(n553), .B(n554), .Z(n551) );
  NANDN U485 ( .A(B[374]), .B(A[374]), .Z(n554) );
  AND U486 ( .A(n555), .B(n556), .Z(n553) );
  NAND U487 ( .A(n557), .B(n558), .Z(n556) );
  NANDN U488 ( .A(A[373]), .B(B[373]), .Z(n558) );
  AND U489 ( .A(n559), .B(n560), .Z(n557) );
  NANDN U490 ( .A(A[372]), .B(B[372]), .Z(n560) );
  NAND U491 ( .A(n561), .B(n562), .Z(n559) );
  NANDN U492 ( .A(B[372]), .B(A[372]), .Z(n562) );
  AND U493 ( .A(n563), .B(n564), .Z(n561) );
  NAND U494 ( .A(n565), .B(n566), .Z(n564) );
  NANDN U495 ( .A(A[371]), .B(B[371]), .Z(n566) );
  AND U496 ( .A(n567), .B(n568), .Z(n565) );
  NANDN U497 ( .A(A[370]), .B(B[370]), .Z(n568) );
  NAND U498 ( .A(n569), .B(n570), .Z(n567) );
  NANDN U499 ( .A(B[370]), .B(A[370]), .Z(n570) );
  AND U500 ( .A(n571), .B(n572), .Z(n569) );
  NAND U501 ( .A(n573), .B(n574), .Z(n572) );
  NANDN U502 ( .A(A[369]), .B(B[369]), .Z(n574) );
  AND U503 ( .A(n575), .B(n576), .Z(n573) );
  NANDN U504 ( .A(A[368]), .B(B[368]), .Z(n576) );
  NAND U505 ( .A(n577), .B(n578), .Z(n575) );
  NANDN U506 ( .A(B[368]), .B(A[368]), .Z(n578) );
  AND U507 ( .A(n579), .B(n580), .Z(n577) );
  NAND U508 ( .A(n581), .B(n582), .Z(n580) );
  NANDN U509 ( .A(A[367]), .B(B[367]), .Z(n582) );
  AND U510 ( .A(n583), .B(n584), .Z(n581) );
  NANDN U511 ( .A(A[366]), .B(B[366]), .Z(n584) );
  NAND U512 ( .A(n585), .B(n586), .Z(n583) );
  NANDN U513 ( .A(B[366]), .B(A[366]), .Z(n586) );
  AND U514 ( .A(n587), .B(n588), .Z(n585) );
  NAND U515 ( .A(n589), .B(n590), .Z(n588) );
  NANDN U516 ( .A(A[365]), .B(B[365]), .Z(n590) );
  AND U517 ( .A(n591), .B(n592), .Z(n589) );
  NANDN U518 ( .A(A[364]), .B(B[364]), .Z(n592) );
  NAND U519 ( .A(n593), .B(n594), .Z(n591) );
  NANDN U520 ( .A(B[364]), .B(A[364]), .Z(n594) );
  AND U521 ( .A(n595), .B(n596), .Z(n593) );
  NAND U522 ( .A(n597), .B(n598), .Z(n596) );
  NANDN U523 ( .A(A[363]), .B(B[363]), .Z(n598) );
  AND U524 ( .A(n599), .B(n600), .Z(n597) );
  NANDN U525 ( .A(A[362]), .B(B[362]), .Z(n600) );
  NAND U526 ( .A(n601), .B(n602), .Z(n599) );
  NANDN U527 ( .A(B[362]), .B(A[362]), .Z(n602) );
  AND U528 ( .A(n603), .B(n604), .Z(n601) );
  NAND U529 ( .A(n605), .B(n606), .Z(n604) );
  NANDN U530 ( .A(A[361]), .B(B[361]), .Z(n606) );
  AND U531 ( .A(n607), .B(n608), .Z(n605) );
  NANDN U532 ( .A(A[360]), .B(B[360]), .Z(n608) );
  NAND U533 ( .A(n609), .B(n610), .Z(n607) );
  NANDN U534 ( .A(B[360]), .B(A[360]), .Z(n610) );
  AND U535 ( .A(n611), .B(n612), .Z(n609) );
  NAND U536 ( .A(n613), .B(n614), .Z(n612) );
  NANDN U537 ( .A(A[359]), .B(B[359]), .Z(n614) );
  AND U538 ( .A(n615), .B(n616), .Z(n613) );
  NANDN U539 ( .A(A[358]), .B(B[358]), .Z(n616) );
  NAND U540 ( .A(n617), .B(n618), .Z(n615) );
  NANDN U541 ( .A(B[358]), .B(A[358]), .Z(n618) );
  AND U542 ( .A(n619), .B(n620), .Z(n617) );
  NAND U543 ( .A(n621), .B(n622), .Z(n620) );
  NANDN U544 ( .A(A[357]), .B(B[357]), .Z(n622) );
  AND U545 ( .A(n623), .B(n624), .Z(n621) );
  NANDN U546 ( .A(A[356]), .B(B[356]), .Z(n624) );
  NAND U547 ( .A(n625), .B(n626), .Z(n623) );
  NANDN U548 ( .A(B[356]), .B(A[356]), .Z(n626) );
  AND U549 ( .A(n627), .B(n628), .Z(n625) );
  NAND U550 ( .A(n629), .B(n630), .Z(n628) );
  NANDN U551 ( .A(A[355]), .B(B[355]), .Z(n630) );
  AND U552 ( .A(n631), .B(n632), .Z(n629) );
  NANDN U553 ( .A(A[354]), .B(B[354]), .Z(n632) );
  NAND U554 ( .A(n633), .B(n634), .Z(n631) );
  NANDN U555 ( .A(B[354]), .B(A[354]), .Z(n634) );
  AND U556 ( .A(n635), .B(n636), .Z(n633) );
  NAND U557 ( .A(n637), .B(n638), .Z(n636) );
  NANDN U558 ( .A(A[353]), .B(B[353]), .Z(n638) );
  AND U559 ( .A(n639), .B(n640), .Z(n637) );
  NANDN U560 ( .A(A[352]), .B(B[352]), .Z(n640) );
  NAND U561 ( .A(n641), .B(n642), .Z(n639) );
  NANDN U562 ( .A(B[352]), .B(A[352]), .Z(n642) );
  AND U563 ( .A(n643), .B(n644), .Z(n641) );
  NAND U564 ( .A(n645), .B(n646), .Z(n644) );
  NANDN U565 ( .A(A[351]), .B(B[351]), .Z(n646) );
  AND U566 ( .A(n647), .B(n648), .Z(n645) );
  NANDN U567 ( .A(A[350]), .B(B[350]), .Z(n648) );
  NAND U568 ( .A(n649), .B(n650), .Z(n647) );
  NANDN U569 ( .A(B[350]), .B(A[350]), .Z(n650) );
  AND U570 ( .A(n651), .B(n652), .Z(n649) );
  NAND U571 ( .A(n653), .B(n654), .Z(n652) );
  NANDN U572 ( .A(A[349]), .B(B[349]), .Z(n654) );
  AND U573 ( .A(n655), .B(n656), .Z(n653) );
  NANDN U574 ( .A(A[348]), .B(B[348]), .Z(n656) );
  NAND U575 ( .A(n657), .B(n658), .Z(n655) );
  NANDN U576 ( .A(B[348]), .B(A[348]), .Z(n658) );
  AND U577 ( .A(n659), .B(n660), .Z(n657) );
  NAND U578 ( .A(n661), .B(n662), .Z(n660) );
  NANDN U579 ( .A(A[347]), .B(B[347]), .Z(n662) );
  AND U580 ( .A(n663), .B(n664), .Z(n661) );
  NANDN U581 ( .A(A[346]), .B(B[346]), .Z(n664) );
  NAND U582 ( .A(n665), .B(n666), .Z(n663) );
  NANDN U583 ( .A(B[346]), .B(A[346]), .Z(n666) );
  AND U584 ( .A(n667), .B(n668), .Z(n665) );
  NAND U585 ( .A(n669), .B(n670), .Z(n668) );
  NANDN U586 ( .A(A[345]), .B(B[345]), .Z(n670) );
  AND U587 ( .A(n671), .B(n672), .Z(n669) );
  NANDN U588 ( .A(A[344]), .B(B[344]), .Z(n672) );
  NAND U589 ( .A(n673), .B(n674), .Z(n671) );
  NANDN U590 ( .A(B[344]), .B(A[344]), .Z(n674) );
  AND U591 ( .A(n675), .B(n676), .Z(n673) );
  NAND U592 ( .A(n677), .B(n678), .Z(n676) );
  NANDN U593 ( .A(A[343]), .B(B[343]), .Z(n678) );
  AND U594 ( .A(n679), .B(n680), .Z(n677) );
  NANDN U595 ( .A(A[342]), .B(B[342]), .Z(n680) );
  NAND U596 ( .A(n681), .B(n682), .Z(n679) );
  NANDN U597 ( .A(B[342]), .B(A[342]), .Z(n682) );
  AND U598 ( .A(n683), .B(n684), .Z(n681) );
  NAND U599 ( .A(n685), .B(n686), .Z(n684) );
  NANDN U600 ( .A(A[341]), .B(B[341]), .Z(n686) );
  AND U601 ( .A(n687), .B(n688), .Z(n685) );
  NANDN U602 ( .A(A[340]), .B(B[340]), .Z(n688) );
  NAND U603 ( .A(n689), .B(n690), .Z(n687) );
  NANDN U604 ( .A(B[340]), .B(A[340]), .Z(n690) );
  AND U605 ( .A(n691), .B(n692), .Z(n689) );
  NAND U606 ( .A(n693), .B(n694), .Z(n692) );
  NANDN U607 ( .A(A[339]), .B(B[339]), .Z(n694) );
  AND U608 ( .A(n695), .B(n696), .Z(n693) );
  NANDN U609 ( .A(A[338]), .B(B[338]), .Z(n696) );
  NAND U610 ( .A(n697), .B(n698), .Z(n695) );
  NANDN U611 ( .A(B[338]), .B(A[338]), .Z(n698) );
  AND U612 ( .A(n699), .B(n700), .Z(n697) );
  NAND U613 ( .A(n701), .B(n702), .Z(n700) );
  NANDN U614 ( .A(A[337]), .B(B[337]), .Z(n702) );
  AND U615 ( .A(n703), .B(n704), .Z(n701) );
  NANDN U616 ( .A(A[336]), .B(B[336]), .Z(n704) );
  NAND U617 ( .A(n705), .B(n706), .Z(n703) );
  NANDN U618 ( .A(B[336]), .B(A[336]), .Z(n706) );
  AND U619 ( .A(n707), .B(n708), .Z(n705) );
  NAND U620 ( .A(n709), .B(n710), .Z(n708) );
  NANDN U621 ( .A(A[335]), .B(B[335]), .Z(n710) );
  AND U622 ( .A(n711), .B(n712), .Z(n709) );
  NANDN U623 ( .A(A[334]), .B(B[334]), .Z(n712) );
  NAND U624 ( .A(n713), .B(n714), .Z(n711) );
  NANDN U625 ( .A(B[334]), .B(A[334]), .Z(n714) );
  AND U626 ( .A(n715), .B(n716), .Z(n713) );
  NAND U627 ( .A(n717), .B(n718), .Z(n716) );
  NANDN U628 ( .A(A[333]), .B(B[333]), .Z(n718) );
  AND U629 ( .A(n719), .B(n720), .Z(n717) );
  NANDN U630 ( .A(A[332]), .B(B[332]), .Z(n720) );
  NAND U631 ( .A(n721), .B(n722), .Z(n719) );
  NANDN U632 ( .A(B[332]), .B(A[332]), .Z(n722) );
  AND U633 ( .A(n723), .B(n724), .Z(n721) );
  NAND U634 ( .A(n725), .B(n726), .Z(n724) );
  NANDN U635 ( .A(A[331]), .B(B[331]), .Z(n726) );
  AND U636 ( .A(n727), .B(n728), .Z(n725) );
  NANDN U637 ( .A(A[330]), .B(B[330]), .Z(n728) );
  NAND U638 ( .A(n729), .B(n730), .Z(n727) );
  NANDN U639 ( .A(B[330]), .B(A[330]), .Z(n730) );
  AND U640 ( .A(n731), .B(n732), .Z(n729) );
  NAND U641 ( .A(n733), .B(n734), .Z(n732) );
  NANDN U642 ( .A(A[329]), .B(B[329]), .Z(n734) );
  AND U643 ( .A(n735), .B(n736), .Z(n733) );
  NANDN U644 ( .A(A[328]), .B(B[328]), .Z(n736) );
  NAND U645 ( .A(n737), .B(n738), .Z(n735) );
  NANDN U646 ( .A(B[328]), .B(A[328]), .Z(n738) );
  AND U647 ( .A(n739), .B(n740), .Z(n737) );
  NAND U648 ( .A(n741), .B(n742), .Z(n740) );
  NANDN U649 ( .A(A[327]), .B(B[327]), .Z(n742) );
  AND U650 ( .A(n743), .B(n744), .Z(n741) );
  NANDN U651 ( .A(A[326]), .B(B[326]), .Z(n744) );
  NAND U652 ( .A(n745), .B(n746), .Z(n743) );
  NANDN U653 ( .A(B[326]), .B(A[326]), .Z(n746) );
  AND U654 ( .A(n747), .B(n748), .Z(n745) );
  NAND U655 ( .A(n749), .B(n750), .Z(n748) );
  NANDN U656 ( .A(A[325]), .B(B[325]), .Z(n750) );
  AND U657 ( .A(n751), .B(n752), .Z(n749) );
  NANDN U658 ( .A(A[324]), .B(B[324]), .Z(n752) );
  NAND U659 ( .A(n753), .B(n754), .Z(n751) );
  NANDN U660 ( .A(B[324]), .B(A[324]), .Z(n754) );
  AND U661 ( .A(n755), .B(n756), .Z(n753) );
  NAND U662 ( .A(n757), .B(n758), .Z(n756) );
  NANDN U663 ( .A(A[323]), .B(B[323]), .Z(n758) );
  AND U664 ( .A(n759), .B(n760), .Z(n757) );
  NANDN U665 ( .A(A[322]), .B(B[322]), .Z(n760) );
  NAND U666 ( .A(n761), .B(n762), .Z(n759) );
  NANDN U667 ( .A(B[322]), .B(A[322]), .Z(n762) );
  AND U668 ( .A(n763), .B(n764), .Z(n761) );
  NAND U669 ( .A(n765), .B(n766), .Z(n764) );
  NANDN U670 ( .A(A[321]), .B(B[321]), .Z(n766) );
  AND U671 ( .A(n767), .B(n768), .Z(n765) );
  NANDN U672 ( .A(A[320]), .B(B[320]), .Z(n768) );
  NAND U673 ( .A(n769), .B(n770), .Z(n767) );
  NANDN U674 ( .A(B[320]), .B(A[320]), .Z(n770) );
  AND U675 ( .A(n771), .B(n772), .Z(n769) );
  NAND U676 ( .A(n773), .B(n774), .Z(n772) );
  NANDN U677 ( .A(A[319]), .B(B[319]), .Z(n774) );
  AND U678 ( .A(n775), .B(n776), .Z(n773) );
  NANDN U679 ( .A(A[318]), .B(B[318]), .Z(n776) );
  NAND U680 ( .A(n777), .B(n778), .Z(n775) );
  NANDN U681 ( .A(B[318]), .B(A[318]), .Z(n778) );
  AND U682 ( .A(n779), .B(n780), .Z(n777) );
  NAND U683 ( .A(n781), .B(n782), .Z(n780) );
  NANDN U684 ( .A(A[317]), .B(B[317]), .Z(n782) );
  AND U685 ( .A(n783), .B(n784), .Z(n781) );
  NANDN U686 ( .A(A[316]), .B(B[316]), .Z(n784) );
  NAND U687 ( .A(n785), .B(n786), .Z(n783) );
  NANDN U688 ( .A(B[316]), .B(A[316]), .Z(n786) );
  AND U689 ( .A(n787), .B(n788), .Z(n785) );
  NAND U690 ( .A(n789), .B(n790), .Z(n788) );
  NANDN U691 ( .A(A[315]), .B(B[315]), .Z(n790) );
  AND U692 ( .A(n791), .B(n792), .Z(n789) );
  NANDN U693 ( .A(A[314]), .B(B[314]), .Z(n792) );
  NAND U694 ( .A(n793), .B(n794), .Z(n791) );
  NANDN U695 ( .A(B[314]), .B(A[314]), .Z(n794) );
  AND U696 ( .A(n795), .B(n796), .Z(n793) );
  NAND U697 ( .A(n797), .B(n798), .Z(n796) );
  NANDN U698 ( .A(A[313]), .B(B[313]), .Z(n798) );
  AND U699 ( .A(n799), .B(n800), .Z(n797) );
  NANDN U700 ( .A(A[312]), .B(B[312]), .Z(n800) );
  NAND U701 ( .A(n801), .B(n802), .Z(n799) );
  NANDN U702 ( .A(B[312]), .B(A[312]), .Z(n802) );
  AND U703 ( .A(n803), .B(n804), .Z(n801) );
  NAND U704 ( .A(n805), .B(n806), .Z(n804) );
  NANDN U705 ( .A(A[311]), .B(B[311]), .Z(n806) );
  AND U706 ( .A(n807), .B(n808), .Z(n805) );
  NANDN U707 ( .A(A[310]), .B(B[310]), .Z(n808) );
  NAND U708 ( .A(n809), .B(n810), .Z(n807) );
  NANDN U709 ( .A(B[310]), .B(A[310]), .Z(n810) );
  AND U710 ( .A(n811), .B(n812), .Z(n809) );
  NAND U711 ( .A(n813), .B(n814), .Z(n812) );
  NANDN U712 ( .A(A[309]), .B(B[309]), .Z(n814) );
  AND U713 ( .A(n815), .B(n816), .Z(n813) );
  NANDN U714 ( .A(A[308]), .B(B[308]), .Z(n816) );
  NAND U715 ( .A(n817), .B(n818), .Z(n815) );
  NANDN U716 ( .A(B[308]), .B(A[308]), .Z(n818) );
  AND U717 ( .A(n819), .B(n820), .Z(n817) );
  NAND U718 ( .A(n821), .B(n822), .Z(n820) );
  NANDN U719 ( .A(A[307]), .B(B[307]), .Z(n822) );
  AND U720 ( .A(n823), .B(n824), .Z(n821) );
  NANDN U721 ( .A(A[306]), .B(B[306]), .Z(n824) );
  NAND U722 ( .A(n825), .B(n826), .Z(n823) );
  NANDN U723 ( .A(B[306]), .B(A[306]), .Z(n826) );
  AND U724 ( .A(n827), .B(n828), .Z(n825) );
  NAND U725 ( .A(n829), .B(n830), .Z(n828) );
  NANDN U726 ( .A(A[305]), .B(B[305]), .Z(n830) );
  AND U727 ( .A(n831), .B(n832), .Z(n829) );
  NANDN U728 ( .A(A[304]), .B(B[304]), .Z(n832) );
  NAND U729 ( .A(n833), .B(n834), .Z(n831) );
  NANDN U730 ( .A(B[304]), .B(A[304]), .Z(n834) );
  AND U731 ( .A(n835), .B(n836), .Z(n833) );
  NAND U732 ( .A(n837), .B(n838), .Z(n836) );
  NANDN U733 ( .A(A[303]), .B(B[303]), .Z(n838) );
  AND U734 ( .A(n839), .B(n840), .Z(n837) );
  NANDN U735 ( .A(A[302]), .B(B[302]), .Z(n840) );
  NAND U736 ( .A(n841), .B(n842), .Z(n839) );
  NANDN U737 ( .A(B[302]), .B(A[302]), .Z(n842) );
  AND U738 ( .A(n843), .B(n844), .Z(n841) );
  NAND U739 ( .A(n845), .B(n846), .Z(n844) );
  NANDN U740 ( .A(A[301]), .B(B[301]), .Z(n846) );
  AND U741 ( .A(n847), .B(n848), .Z(n845) );
  NANDN U742 ( .A(A[300]), .B(B[300]), .Z(n848) );
  NAND U743 ( .A(n849), .B(n850), .Z(n847) );
  NANDN U744 ( .A(B[300]), .B(A[300]), .Z(n850) );
  AND U745 ( .A(n851), .B(n852), .Z(n849) );
  NAND U746 ( .A(n853), .B(n854), .Z(n852) );
  NANDN U747 ( .A(A[299]), .B(B[299]), .Z(n854) );
  AND U748 ( .A(n855), .B(n856), .Z(n853) );
  NANDN U749 ( .A(A[298]), .B(B[298]), .Z(n856) );
  NAND U750 ( .A(n857), .B(n858), .Z(n855) );
  NANDN U751 ( .A(B[298]), .B(A[298]), .Z(n858) );
  AND U752 ( .A(n859), .B(n860), .Z(n857) );
  NAND U753 ( .A(n861), .B(n862), .Z(n860) );
  NANDN U754 ( .A(A[297]), .B(B[297]), .Z(n862) );
  AND U755 ( .A(n863), .B(n864), .Z(n861) );
  NANDN U756 ( .A(A[296]), .B(B[296]), .Z(n864) );
  NAND U757 ( .A(n865), .B(n866), .Z(n863) );
  NANDN U758 ( .A(B[296]), .B(A[296]), .Z(n866) );
  AND U759 ( .A(n867), .B(n868), .Z(n865) );
  NAND U760 ( .A(n869), .B(n870), .Z(n868) );
  NANDN U761 ( .A(A[295]), .B(B[295]), .Z(n870) );
  AND U762 ( .A(n871), .B(n872), .Z(n869) );
  NANDN U763 ( .A(A[294]), .B(B[294]), .Z(n872) );
  NAND U764 ( .A(n873), .B(n874), .Z(n871) );
  NANDN U765 ( .A(B[294]), .B(A[294]), .Z(n874) );
  AND U766 ( .A(n875), .B(n876), .Z(n873) );
  NAND U767 ( .A(n877), .B(n878), .Z(n876) );
  NANDN U768 ( .A(A[293]), .B(B[293]), .Z(n878) );
  AND U769 ( .A(n879), .B(n880), .Z(n877) );
  NANDN U770 ( .A(A[292]), .B(B[292]), .Z(n880) );
  NAND U771 ( .A(n881), .B(n882), .Z(n879) );
  NANDN U772 ( .A(B[292]), .B(A[292]), .Z(n882) );
  AND U773 ( .A(n883), .B(n884), .Z(n881) );
  NAND U774 ( .A(n885), .B(n886), .Z(n884) );
  NANDN U775 ( .A(A[291]), .B(B[291]), .Z(n886) );
  AND U776 ( .A(n887), .B(n888), .Z(n885) );
  NANDN U777 ( .A(A[290]), .B(B[290]), .Z(n888) );
  NAND U778 ( .A(n889), .B(n890), .Z(n887) );
  NANDN U779 ( .A(B[290]), .B(A[290]), .Z(n890) );
  AND U780 ( .A(n891), .B(n892), .Z(n889) );
  NAND U781 ( .A(n893), .B(n894), .Z(n892) );
  NANDN U782 ( .A(A[289]), .B(B[289]), .Z(n894) );
  AND U783 ( .A(n895), .B(n896), .Z(n893) );
  NANDN U784 ( .A(A[288]), .B(B[288]), .Z(n896) );
  NAND U785 ( .A(n897), .B(n898), .Z(n895) );
  NANDN U786 ( .A(B[288]), .B(A[288]), .Z(n898) );
  AND U787 ( .A(n899), .B(n900), .Z(n897) );
  NAND U788 ( .A(n901), .B(n902), .Z(n900) );
  NANDN U789 ( .A(A[287]), .B(B[287]), .Z(n902) );
  AND U790 ( .A(n903), .B(n904), .Z(n901) );
  NANDN U791 ( .A(A[286]), .B(B[286]), .Z(n904) );
  NAND U792 ( .A(n905), .B(n906), .Z(n903) );
  NANDN U793 ( .A(B[286]), .B(A[286]), .Z(n906) );
  AND U794 ( .A(n907), .B(n908), .Z(n905) );
  NAND U795 ( .A(n909), .B(n910), .Z(n908) );
  NANDN U796 ( .A(A[285]), .B(B[285]), .Z(n910) );
  AND U797 ( .A(n911), .B(n912), .Z(n909) );
  NANDN U798 ( .A(A[284]), .B(B[284]), .Z(n912) );
  NAND U799 ( .A(n913), .B(n914), .Z(n911) );
  NANDN U800 ( .A(B[284]), .B(A[284]), .Z(n914) );
  AND U801 ( .A(n915), .B(n916), .Z(n913) );
  NAND U802 ( .A(n917), .B(n918), .Z(n916) );
  NANDN U803 ( .A(A[283]), .B(B[283]), .Z(n918) );
  AND U804 ( .A(n919), .B(n920), .Z(n917) );
  NANDN U805 ( .A(A[282]), .B(B[282]), .Z(n920) );
  NAND U806 ( .A(n921), .B(n922), .Z(n919) );
  NANDN U807 ( .A(B[282]), .B(A[282]), .Z(n922) );
  AND U808 ( .A(n923), .B(n924), .Z(n921) );
  NAND U809 ( .A(n925), .B(n926), .Z(n924) );
  NANDN U810 ( .A(A[281]), .B(B[281]), .Z(n926) );
  AND U811 ( .A(n927), .B(n928), .Z(n925) );
  NANDN U812 ( .A(A[280]), .B(B[280]), .Z(n928) );
  NAND U813 ( .A(n929), .B(n930), .Z(n927) );
  NANDN U814 ( .A(B[280]), .B(A[280]), .Z(n930) );
  AND U815 ( .A(n931), .B(n932), .Z(n929) );
  NAND U816 ( .A(n933), .B(n934), .Z(n932) );
  NANDN U817 ( .A(A[279]), .B(B[279]), .Z(n934) );
  AND U818 ( .A(n935), .B(n936), .Z(n933) );
  NANDN U819 ( .A(A[278]), .B(B[278]), .Z(n936) );
  NAND U820 ( .A(n937), .B(n938), .Z(n935) );
  NANDN U821 ( .A(B[278]), .B(A[278]), .Z(n938) );
  AND U822 ( .A(n939), .B(n940), .Z(n937) );
  NAND U823 ( .A(n941), .B(n942), .Z(n940) );
  NANDN U824 ( .A(A[277]), .B(B[277]), .Z(n942) );
  AND U825 ( .A(n943), .B(n944), .Z(n941) );
  NANDN U826 ( .A(A[276]), .B(B[276]), .Z(n944) );
  NAND U827 ( .A(n945), .B(n946), .Z(n943) );
  NANDN U828 ( .A(B[276]), .B(A[276]), .Z(n946) );
  AND U829 ( .A(n947), .B(n948), .Z(n945) );
  NAND U830 ( .A(n949), .B(n950), .Z(n948) );
  NANDN U831 ( .A(A[275]), .B(B[275]), .Z(n950) );
  AND U832 ( .A(n951), .B(n952), .Z(n949) );
  NANDN U833 ( .A(A[274]), .B(B[274]), .Z(n952) );
  NAND U834 ( .A(n953), .B(n954), .Z(n951) );
  NANDN U835 ( .A(B[274]), .B(A[274]), .Z(n954) );
  AND U836 ( .A(n955), .B(n956), .Z(n953) );
  NAND U837 ( .A(n957), .B(n958), .Z(n956) );
  NANDN U838 ( .A(A[273]), .B(B[273]), .Z(n958) );
  AND U839 ( .A(n959), .B(n960), .Z(n957) );
  NANDN U840 ( .A(A[272]), .B(B[272]), .Z(n960) );
  NAND U841 ( .A(n961), .B(n962), .Z(n959) );
  NANDN U842 ( .A(B[272]), .B(A[272]), .Z(n962) );
  AND U843 ( .A(n963), .B(n964), .Z(n961) );
  NAND U844 ( .A(n965), .B(n966), .Z(n964) );
  NANDN U845 ( .A(A[271]), .B(B[271]), .Z(n966) );
  AND U846 ( .A(n967), .B(n968), .Z(n965) );
  NANDN U847 ( .A(A[270]), .B(B[270]), .Z(n968) );
  NAND U848 ( .A(n969), .B(n970), .Z(n967) );
  NANDN U849 ( .A(B[270]), .B(A[270]), .Z(n970) );
  AND U850 ( .A(n971), .B(n972), .Z(n969) );
  NAND U851 ( .A(n973), .B(n974), .Z(n972) );
  NANDN U852 ( .A(A[269]), .B(B[269]), .Z(n974) );
  AND U853 ( .A(n975), .B(n976), .Z(n973) );
  NANDN U854 ( .A(A[268]), .B(B[268]), .Z(n976) );
  NAND U855 ( .A(n977), .B(n978), .Z(n975) );
  NANDN U856 ( .A(B[268]), .B(A[268]), .Z(n978) );
  AND U857 ( .A(n979), .B(n980), .Z(n977) );
  NAND U858 ( .A(n981), .B(n982), .Z(n980) );
  NANDN U859 ( .A(A[267]), .B(B[267]), .Z(n982) );
  AND U860 ( .A(n983), .B(n984), .Z(n981) );
  NANDN U861 ( .A(A[266]), .B(B[266]), .Z(n984) );
  NAND U862 ( .A(n985), .B(n986), .Z(n983) );
  NANDN U863 ( .A(B[266]), .B(A[266]), .Z(n986) );
  AND U864 ( .A(n987), .B(n988), .Z(n985) );
  NAND U865 ( .A(n989), .B(n990), .Z(n988) );
  NANDN U866 ( .A(A[265]), .B(B[265]), .Z(n990) );
  AND U867 ( .A(n991), .B(n992), .Z(n989) );
  NANDN U868 ( .A(A[264]), .B(B[264]), .Z(n992) );
  NAND U869 ( .A(n993), .B(n994), .Z(n991) );
  NANDN U870 ( .A(B[264]), .B(A[264]), .Z(n994) );
  AND U871 ( .A(n995), .B(n996), .Z(n993) );
  NAND U872 ( .A(n997), .B(n998), .Z(n996) );
  NANDN U873 ( .A(A[263]), .B(B[263]), .Z(n998) );
  AND U874 ( .A(n999), .B(n1000), .Z(n997) );
  NANDN U875 ( .A(A[262]), .B(B[262]), .Z(n1000) );
  NAND U876 ( .A(n1001), .B(n1002), .Z(n999) );
  NANDN U877 ( .A(B[262]), .B(A[262]), .Z(n1002) );
  AND U878 ( .A(n1003), .B(n1004), .Z(n1001) );
  NAND U879 ( .A(n1005), .B(n1006), .Z(n1004) );
  NANDN U880 ( .A(A[261]), .B(B[261]), .Z(n1006) );
  AND U881 ( .A(n1007), .B(n1008), .Z(n1005) );
  NANDN U882 ( .A(A[260]), .B(B[260]), .Z(n1008) );
  NAND U883 ( .A(n1009), .B(n1010), .Z(n1007) );
  NANDN U884 ( .A(B[260]), .B(A[260]), .Z(n1010) );
  AND U885 ( .A(n1011), .B(n1012), .Z(n1009) );
  NAND U886 ( .A(n1013), .B(n1014), .Z(n1012) );
  NANDN U887 ( .A(A[259]), .B(B[259]), .Z(n1014) );
  AND U888 ( .A(n1015), .B(n1016), .Z(n1013) );
  NANDN U889 ( .A(A[258]), .B(B[258]), .Z(n1016) );
  NAND U890 ( .A(n1017), .B(n1018), .Z(n1015) );
  NANDN U891 ( .A(B[258]), .B(A[258]), .Z(n1018) );
  AND U892 ( .A(n1019), .B(n1020), .Z(n1017) );
  NAND U893 ( .A(n1021), .B(n1022), .Z(n1020) );
  NANDN U894 ( .A(A[257]), .B(B[257]), .Z(n1022) );
  AND U895 ( .A(n1023), .B(n1024), .Z(n1021) );
  NANDN U896 ( .A(A[256]), .B(B[256]), .Z(n1024) );
  NAND U897 ( .A(n1025), .B(n1026), .Z(n1023) );
  NANDN U898 ( .A(B[256]), .B(A[256]), .Z(n1026) );
  AND U899 ( .A(n1027), .B(n1028), .Z(n1025) );
  NAND U900 ( .A(n1029), .B(n1030), .Z(n1028) );
  NANDN U901 ( .A(A[255]), .B(B[255]), .Z(n1030) );
  AND U902 ( .A(n1031), .B(n1032), .Z(n1029) );
  NANDN U903 ( .A(A[254]), .B(B[254]), .Z(n1032) );
  NAND U904 ( .A(n1033), .B(n1034), .Z(n1031) );
  NANDN U905 ( .A(B[254]), .B(A[254]), .Z(n1034) );
  AND U906 ( .A(n1035), .B(n1036), .Z(n1033) );
  NAND U907 ( .A(n1037), .B(n1038), .Z(n1036) );
  NANDN U908 ( .A(A[253]), .B(B[253]), .Z(n1038) );
  AND U909 ( .A(n1039), .B(n1040), .Z(n1037) );
  NANDN U910 ( .A(A[252]), .B(B[252]), .Z(n1040) );
  NAND U911 ( .A(n1041), .B(n1042), .Z(n1039) );
  NANDN U912 ( .A(B[252]), .B(A[252]), .Z(n1042) );
  AND U913 ( .A(n1043), .B(n1044), .Z(n1041) );
  NAND U914 ( .A(n1045), .B(n1046), .Z(n1044) );
  NANDN U915 ( .A(A[251]), .B(B[251]), .Z(n1046) );
  AND U916 ( .A(n1047), .B(n1048), .Z(n1045) );
  NANDN U917 ( .A(A[250]), .B(B[250]), .Z(n1048) );
  NAND U918 ( .A(n1049), .B(n1050), .Z(n1047) );
  NANDN U919 ( .A(B[250]), .B(A[250]), .Z(n1050) );
  AND U920 ( .A(n1051), .B(n1052), .Z(n1049) );
  NAND U921 ( .A(n1053), .B(n1054), .Z(n1052) );
  NANDN U922 ( .A(A[249]), .B(B[249]), .Z(n1054) );
  AND U923 ( .A(n1055), .B(n1056), .Z(n1053) );
  NANDN U924 ( .A(A[248]), .B(B[248]), .Z(n1056) );
  NAND U925 ( .A(n1057), .B(n1058), .Z(n1055) );
  NANDN U926 ( .A(B[248]), .B(A[248]), .Z(n1058) );
  AND U927 ( .A(n1059), .B(n1060), .Z(n1057) );
  NAND U928 ( .A(n1061), .B(n1062), .Z(n1060) );
  NANDN U929 ( .A(A[247]), .B(B[247]), .Z(n1062) );
  AND U930 ( .A(n1063), .B(n1064), .Z(n1061) );
  NANDN U931 ( .A(A[246]), .B(B[246]), .Z(n1064) );
  NAND U932 ( .A(n1065), .B(n1066), .Z(n1063) );
  NANDN U933 ( .A(B[246]), .B(A[246]), .Z(n1066) );
  AND U934 ( .A(n1067), .B(n1068), .Z(n1065) );
  NAND U935 ( .A(n1069), .B(n1070), .Z(n1068) );
  NANDN U936 ( .A(A[245]), .B(B[245]), .Z(n1070) );
  AND U937 ( .A(n1071), .B(n1072), .Z(n1069) );
  NANDN U938 ( .A(A[244]), .B(B[244]), .Z(n1072) );
  NAND U939 ( .A(n1073), .B(n1074), .Z(n1071) );
  NANDN U940 ( .A(B[244]), .B(A[244]), .Z(n1074) );
  AND U941 ( .A(n1075), .B(n1076), .Z(n1073) );
  NAND U942 ( .A(n1077), .B(n1078), .Z(n1076) );
  NANDN U943 ( .A(A[243]), .B(B[243]), .Z(n1078) );
  AND U944 ( .A(n1079), .B(n1080), .Z(n1077) );
  NANDN U945 ( .A(A[242]), .B(B[242]), .Z(n1080) );
  NAND U946 ( .A(n1081), .B(n1082), .Z(n1079) );
  NANDN U947 ( .A(B[242]), .B(A[242]), .Z(n1082) );
  AND U948 ( .A(n1083), .B(n1084), .Z(n1081) );
  NAND U949 ( .A(n1085), .B(n1086), .Z(n1084) );
  NANDN U950 ( .A(A[241]), .B(B[241]), .Z(n1086) );
  AND U951 ( .A(n1087), .B(n1088), .Z(n1085) );
  NANDN U952 ( .A(A[240]), .B(B[240]), .Z(n1088) );
  NAND U953 ( .A(n1089), .B(n1090), .Z(n1087) );
  NANDN U954 ( .A(B[240]), .B(A[240]), .Z(n1090) );
  AND U955 ( .A(n1091), .B(n1092), .Z(n1089) );
  NAND U956 ( .A(n1093), .B(n1094), .Z(n1092) );
  NANDN U957 ( .A(A[239]), .B(B[239]), .Z(n1094) );
  AND U958 ( .A(n1095), .B(n1096), .Z(n1093) );
  NANDN U959 ( .A(A[238]), .B(B[238]), .Z(n1096) );
  NAND U960 ( .A(n1097), .B(n1098), .Z(n1095) );
  NANDN U961 ( .A(B[238]), .B(A[238]), .Z(n1098) );
  AND U962 ( .A(n1099), .B(n1100), .Z(n1097) );
  NAND U963 ( .A(n1101), .B(n1102), .Z(n1100) );
  NANDN U964 ( .A(A[237]), .B(B[237]), .Z(n1102) );
  AND U965 ( .A(n1103), .B(n1104), .Z(n1101) );
  NANDN U966 ( .A(A[236]), .B(B[236]), .Z(n1104) );
  NAND U967 ( .A(n1105), .B(n1106), .Z(n1103) );
  NANDN U968 ( .A(B[236]), .B(A[236]), .Z(n1106) );
  AND U969 ( .A(n1107), .B(n1108), .Z(n1105) );
  NAND U970 ( .A(n1109), .B(n1110), .Z(n1108) );
  NANDN U971 ( .A(A[235]), .B(B[235]), .Z(n1110) );
  AND U972 ( .A(n1111), .B(n1112), .Z(n1109) );
  NANDN U973 ( .A(A[234]), .B(B[234]), .Z(n1112) );
  NAND U974 ( .A(n1113), .B(n1114), .Z(n1111) );
  NANDN U975 ( .A(B[234]), .B(A[234]), .Z(n1114) );
  AND U976 ( .A(n1115), .B(n1116), .Z(n1113) );
  NAND U977 ( .A(n1117), .B(n1118), .Z(n1116) );
  NANDN U978 ( .A(A[233]), .B(B[233]), .Z(n1118) );
  AND U979 ( .A(n1119), .B(n1120), .Z(n1117) );
  NANDN U980 ( .A(A[232]), .B(B[232]), .Z(n1120) );
  NAND U981 ( .A(n1121), .B(n1122), .Z(n1119) );
  NANDN U982 ( .A(B[232]), .B(A[232]), .Z(n1122) );
  AND U983 ( .A(n1123), .B(n1124), .Z(n1121) );
  NAND U984 ( .A(n1125), .B(n1126), .Z(n1124) );
  NANDN U985 ( .A(A[231]), .B(B[231]), .Z(n1126) );
  AND U986 ( .A(n1127), .B(n1128), .Z(n1125) );
  NANDN U987 ( .A(A[230]), .B(B[230]), .Z(n1128) );
  NAND U988 ( .A(n1129), .B(n1130), .Z(n1127) );
  NANDN U989 ( .A(B[230]), .B(A[230]), .Z(n1130) );
  AND U990 ( .A(n1131), .B(n1132), .Z(n1129) );
  NAND U991 ( .A(n1133), .B(n1134), .Z(n1132) );
  NANDN U992 ( .A(A[229]), .B(B[229]), .Z(n1134) );
  AND U993 ( .A(n1135), .B(n1136), .Z(n1133) );
  NANDN U994 ( .A(A[228]), .B(B[228]), .Z(n1136) );
  NAND U995 ( .A(n1137), .B(n1138), .Z(n1135) );
  NANDN U996 ( .A(B[228]), .B(A[228]), .Z(n1138) );
  AND U997 ( .A(n1139), .B(n1140), .Z(n1137) );
  NAND U998 ( .A(n1141), .B(n1142), .Z(n1140) );
  NANDN U999 ( .A(A[227]), .B(B[227]), .Z(n1142) );
  AND U1000 ( .A(n1143), .B(n1144), .Z(n1141) );
  NANDN U1001 ( .A(A[226]), .B(B[226]), .Z(n1144) );
  NAND U1002 ( .A(n1145), .B(n1146), .Z(n1143) );
  NANDN U1003 ( .A(B[226]), .B(A[226]), .Z(n1146) );
  AND U1004 ( .A(n1147), .B(n1148), .Z(n1145) );
  NAND U1005 ( .A(n1149), .B(n1150), .Z(n1148) );
  NANDN U1006 ( .A(A[225]), .B(B[225]), .Z(n1150) );
  AND U1007 ( .A(n1151), .B(n1152), .Z(n1149) );
  NANDN U1008 ( .A(A[224]), .B(B[224]), .Z(n1152) );
  NAND U1009 ( .A(n1153), .B(n1154), .Z(n1151) );
  NANDN U1010 ( .A(B[224]), .B(A[224]), .Z(n1154) );
  AND U1011 ( .A(n1155), .B(n1156), .Z(n1153) );
  NAND U1012 ( .A(n1157), .B(n1158), .Z(n1156) );
  NANDN U1013 ( .A(A[223]), .B(B[223]), .Z(n1158) );
  AND U1014 ( .A(n1159), .B(n1160), .Z(n1157) );
  NANDN U1015 ( .A(A[222]), .B(B[222]), .Z(n1160) );
  NAND U1016 ( .A(n1161), .B(n1162), .Z(n1159) );
  NANDN U1017 ( .A(B[222]), .B(A[222]), .Z(n1162) );
  AND U1018 ( .A(n1163), .B(n1164), .Z(n1161) );
  NAND U1019 ( .A(n1165), .B(n1166), .Z(n1164) );
  NANDN U1020 ( .A(A[221]), .B(B[221]), .Z(n1166) );
  AND U1021 ( .A(n1167), .B(n1168), .Z(n1165) );
  NANDN U1022 ( .A(A[220]), .B(B[220]), .Z(n1168) );
  NAND U1023 ( .A(n1169), .B(n1170), .Z(n1167) );
  NANDN U1024 ( .A(B[220]), .B(A[220]), .Z(n1170) );
  AND U1025 ( .A(n1171), .B(n1172), .Z(n1169) );
  NAND U1026 ( .A(n1173), .B(n1174), .Z(n1172) );
  NANDN U1027 ( .A(A[219]), .B(B[219]), .Z(n1174) );
  AND U1028 ( .A(n1175), .B(n1176), .Z(n1173) );
  NANDN U1029 ( .A(A[218]), .B(B[218]), .Z(n1176) );
  NAND U1030 ( .A(n1177), .B(n1178), .Z(n1175) );
  NANDN U1031 ( .A(B[218]), .B(A[218]), .Z(n1178) );
  AND U1032 ( .A(n1179), .B(n1180), .Z(n1177) );
  NAND U1033 ( .A(n1181), .B(n1182), .Z(n1180) );
  NANDN U1034 ( .A(A[217]), .B(B[217]), .Z(n1182) );
  AND U1035 ( .A(n1183), .B(n1184), .Z(n1181) );
  NANDN U1036 ( .A(A[216]), .B(B[216]), .Z(n1184) );
  NAND U1037 ( .A(n1185), .B(n1186), .Z(n1183) );
  NANDN U1038 ( .A(B[216]), .B(A[216]), .Z(n1186) );
  AND U1039 ( .A(n1187), .B(n1188), .Z(n1185) );
  NAND U1040 ( .A(n1189), .B(n1190), .Z(n1188) );
  NANDN U1041 ( .A(A[215]), .B(B[215]), .Z(n1190) );
  AND U1042 ( .A(n1191), .B(n1192), .Z(n1189) );
  NANDN U1043 ( .A(A[214]), .B(B[214]), .Z(n1192) );
  NAND U1044 ( .A(n1193), .B(n1194), .Z(n1191) );
  NANDN U1045 ( .A(B[214]), .B(A[214]), .Z(n1194) );
  AND U1046 ( .A(n1195), .B(n1196), .Z(n1193) );
  NAND U1047 ( .A(n1197), .B(n1198), .Z(n1196) );
  NANDN U1048 ( .A(A[213]), .B(B[213]), .Z(n1198) );
  AND U1049 ( .A(n1199), .B(n1200), .Z(n1197) );
  NANDN U1050 ( .A(A[212]), .B(B[212]), .Z(n1200) );
  NAND U1051 ( .A(n1201), .B(n1202), .Z(n1199) );
  NANDN U1052 ( .A(B[212]), .B(A[212]), .Z(n1202) );
  AND U1053 ( .A(n1203), .B(n1204), .Z(n1201) );
  NAND U1054 ( .A(n1205), .B(n1206), .Z(n1204) );
  NANDN U1055 ( .A(A[211]), .B(B[211]), .Z(n1206) );
  AND U1056 ( .A(n1207), .B(n1208), .Z(n1205) );
  NANDN U1057 ( .A(A[210]), .B(B[210]), .Z(n1208) );
  NAND U1058 ( .A(n1209), .B(n1210), .Z(n1207) );
  NANDN U1059 ( .A(B[210]), .B(A[210]), .Z(n1210) );
  AND U1060 ( .A(n1211), .B(n1212), .Z(n1209) );
  NAND U1061 ( .A(n1213), .B(n1214), .Z(n1212) );
  NANDN U1062 ( .A(A[209]), .B(B[209]), .Z(n1214) );
  AND U1063 ( .A(n1215), .B(n1216), .Z(n1213) );
  NANDN U1064 ( .A(A[208]), .B(B[208]), .Z(n1216) );
  NAND U1065 ( .A(n1217), .B(n1218), .Z(n1215) );
  NANDN U1066 ( .A(B[208]), .B(A[208]), .Z(n1218) );
  AND U1067 ( .A(n1219), .B(n1220), .Z(n1217) );
  NAND U1068 ( .A(n1221), .B(n1222), .Z(n1220) );
  NANDN U1069 ( .A(A[207]), .B(B[207]), .Z(n1222) );
  AND U1070 ( .A(n1223), .B(n1224), .Z(n1221) );
  NANDN U1071 ( .A(A[206]), .B(B[206]), .Z(n1224) );
  NAND U1072 ( .A(n1225), .B(n1226), .Z(n1223) );
  NANDN U1073 ( .A(B[206]), .B(A[206]), .Z(n1226) );
  AND U1074 ( .A(n1227), .B(n1228), .Z(n1225) );
  NAND U1075 ( .A(n1229), .B(n1230), .Z(n1228) );
  NANDN U1076 ( .A(A[205]), .B(B[205]), .Z(n1230) );
  AND U1077 ( .A(n1231), .B(n1232), .Z(n1229) );
  NANDN U1078 ( .A(A[204]), .B(B[204]), .Z(n1232) );
  NAND U1079 ( .A(n1233), .B(n1234), .Z(n1231) );
  NANDN U1080 ( .A(B[204]), .B(A[204]), .Z(n1234) );
  AND U1081 ( .A(n1235), .B(n1236), .Z(n1233) );
  NAND U1082 ( .A(n1237), .B(n1238), .Z(n1236) );
  NANDN U1083 ( .A(A[203]), .B(B[203]), .Z(n1238) );
  AND U1084 ( .A(n1239), .B(n1240), .Z(n1237) );
  NANDN U1085 ( .A(A[202]), .B(B[202]), .Z(n1240) );
  NAND U1086 ( .A(n1241), .B(n1242), .Z(n1239) );
  NANDN U1087 ( .A(B[202]), .B(A[202]), .Z(n1242) );
  AND U1088 ( .A(n1243), .B(n1244), .Z(n1241) );
  NAND U1089 ( .A(n1245), .B(n1246), .Z(n1244) );
  NANDN U1090 ( .A(A[201]), .B(B[201]), .Z(n1246) );
  AND U1091 ( .A(n1247), .B(n1248), .Z(n1245) );
  NANDN U1092 ( .A(A[200]), .B(B[200]), .Z(n1248) );
  NAND U1093 ( .A(n1249), .B(n1250), .Z(n1247) );
  NANDN U1094 ( .A(B[200]), .B(A[200]), .Z(n1250) );
  AND U1095 ( .A(n1251), .B(n1252), .Z(n1249) );
  NAND U1096 ( .A(n1253), .B(n1254), .Z(n1252) );
  NANDN U1097 ( .A(A[199]), .B(B[199]), .Z(n1254) );
  AND U1098 ( .A(n1255), .B(n1256), .Z(n1253) );
  NANDN U1099 ( .A(A[198]), .B(B[198]), .Z(n1256) );
  NAND U1100 ( .A(n1257), .B(n1258), .Z(n1255) );
  NANDN U1101 ( .A(B[198]), .B(A[198]), .Z(n1258) );
  AND U1102 ( .A(n1259), .B(n1260), .Z(n1257) );
  NAND U1103 ( .A(n1261), .B(n1262), .Z(n1260) );
  NANDN U1104 ( .A(A[197]), .B(B[197]), .Z(n1262) );
  AND U1105 ( .A(n1263), .B(n1264), .Z(n1261) );
  NANDN U1106 ( .A(A[196]), .B(B[196]), .Z(n1264) );
  NAND U1107 ( .A(n1265), .B(n1266), .Z(n1263) );
  NANDN U1108 ( .A(B[196]), .B(A[196]), .Z(n1266) );
  AND U1109 ( .A(n1267), .B(n1268), .Z(n1265) );
  NAND U1110 ( .A(n1269), .B(n1270), .Z(n1268) );
  NANDN U1111 ( .A(A[195]), .B(B[195]), .Z(n1270) );
  AND U1112 ( .A(n1271), .B(n1272), .Z(n1269) );
  NANDN U1113 ( .A(A[194]), .B(B[194]), .Z(n1272) );
  NAND U1114 ( .A(n1273), .B(n1274), .Z(n1271) );
  NANDN U1115 ( .A(B[194]), .B(A[194]), .Z(n1274) );
  AND U1116 ( .A(n1275), .B(n1276), .Z(n1273) );
  NAND U1117 ( .A(n1277), .B(n1278), .Z(n1276) );
  NANDN U1118 ( .A(A[193]), .B(B[193]), .Z(n1278) );
  AND U1119 ( .A(n1279), .B(n1280), .Z(n1277) );
  NANDN U1120 ( .A(A[192]), .B(B[192]), .Z(n1280) );
  NAND U1121 ( .A(n1281), .B(n1282), .Z(n1279) );
  NANDN U1122 ( .A(B[192]), .B(A[192]), .Z(n1282) );
  AND U1123 ( .A(n1283), .B(n1284), .Z(n1281) );
  NAND U1124 ( .A(n1285), .B(n1286), .Z(n1284) );
  NANDN U1125 ( .A(A[191]), .B(B[191]), .Z(n1286) );
  AND U1126 ( .A(n1287), .B(n1288), .Z(n1285) );
  NANDN U1127 ( .A(A[190]), .B(B[190]), .Z(n1288) );
  NAND U1128 ( .A(n1289), .B(n1290), .Z(n1287) );
  NANDN U1129 ( .A(B[190]), .B(A[190]), .Z(n1290) );
  AND U1130 ( .A(n1291), .B(n1292), .Z(n1289) );
  NAND U1131 ( .A(n1293), .B(n1294), .Z(n1292) );
  NANDN U1132 ( .A(A[189]), .B(B[189]), .Z(n1294) );
  AND U1133 ( .A(n1295), .B(n1296), .Z(n1293) );
  NANDN U1134 ( .A(A[188]), .B(B[188]), .Z(n1296) );
  NAND U1135 ( .A(n1297), .B(n1298), .Z(n1295) );
  NANDN U1136 ( .A(B[188]), .B(A[188]), .Z(n1298) );
  AND U1137 ( .A(n1299), .B(n1300), .Z(n1297) );
  NAND U1138 ( .A(n1301), .B(n1302), .Z(n1300) );
  NANDN U1139 ( .A(A[187]), .B(B[187]), .Z(n1302) );
  AND U1140 ( .A(n1303), .B(n1304), .Z(n1301) );
  NANDN U1141 ( .A(A[186]), .B(B[186]), .Z(n1304) );
  NAND U1142 ( .A(n1305), .B(n1306), .Z(n1303) );
  NANDN U1143 ( .A(B[186]), .B(A[186]), .Z(n1306) );
  AND U1144 ( .A(n1307), .B(n1308), .Z(n1305) );
  NAND U1145 ( .A(n1309), .B(n1310), .Z(n1308) );
  NANDN U1146 ( .A(A[185]), .B(B[185]), .Z(n1310) );
  AND U1147 ( .A(n1311), .B(n1312), .Z(n1309) );
  NANDN U1148 ( .A(A[184]), .B(B[184]), .Z(n1312) );
  NAND U1149 ( .A(n1313), .B(n1314), .Z(n1311) );
  NANDN U1150 ( .A(B[184]), .B(A[184]), .Z(n1314) );
  AND U1151 ( .A(n1315), .B(n1316), .Z(n1313) );
  NAND U1152 ( .A(n1317), .B(n1318), .Z(n1316) );
  NANDN U1153 ( .A(A[183]), .B(B[183]), .Z(n1318) );
  AND U1154 ( .A(n1319), .B(n1320), .Z(n1317) );
  NANDN U1155 ( .A(A[182]), .B(B[182]), .Z(n1320) );
  NAND U1156 ( .A(n1321), .B(n1322), .Z(n1319) );
  NANDN U1157 ( .A(B[182]), .B(A[182]), .Z(n1322) );
  AND U1158 ( .A(n1323), .B(n1324), .Z(n1321) );
  NAND U1159 ( .A(n1325), .B(n1326), .Z(n1324) );
  NANDN U1160 ( .A(A[181]), .B(B[181]), .Z(n1326) );
  AND U1161 ( .A(n1327), .B(n1328), .Z(n1325) );
  NANDN U1162 ( .A(A[180]), .B(B[180]), .Z(n1328) );
  NAND U1163 ( .A(n1329), .B(n1330), .Z(n1327) );
  NANDN U1164 ( .A(B[180]), .B(A[180]), .Z(n1330) );
  AND U1165 ( .A(n1331), .B(n1332), .Z(n1329) );
  NAND U1166 ( .A(n1333), .B(n1334), .Z(n1332) );
  NANDN U1167 ( .A(A[179]), .B(B[179]), .Z(n1334) );
  AND U1168 ( .A(n1335), .B(n1336), .Z(n1333) );
  NANDN U1169 ( .A(A[178]), .B(B[178]), .Z(n1336) );
  NAND U1170 ( .A(n1337), .B(n1338), .Z(n1335) );
  NANDN U1171 ( .A(B[178]), .B(A[178]), .Z(n1338) );
  AND U1172 ( .A(n1339), .B(n1340), .Z(n1337) );
  NAND U1173 ( .A(n1341), .B(n1342), .Z(n1340) );
  NANDN U1174 ( .A(A[177]), .B(B[177]), .Z(n1342) );
  AND U1175 ( .A(n1343), .B(n1344), .Z(n1341) );
  NANDN U1176 ( .A(A[176]), .B(B[176]), .Z(n1344) );
  NAND U1177 ( .A(n1345), .B(n1346), .Z(n1343) );
  NANDN U1178 ( .A(B[176]), .B(A[176]), .Z(n1346) );
  AND U1179 ( .A(n1347), .B(n1348), .Z(n1345) );
  NAND U1180 ( .A(n1349), .B(n1350), .Z(n1348) );
  NANDN U1181 ( .A(A[175]), .B(B[175]), .Z(n1350) );
  AND U1182 ( .A(n1351), .B(n1352), .Z(n1349) );
  NANDN U1183 ( .A(A[174]), .B(B[174]), .Z(n1352) );
  NAND U1184 ( .A(n1353), .B(n1354), .Z(n1351) );
  NANDN U1185 ( .A(B[174]), .B(A[174]), .Z(n1354) );
  AND U1186 ( .A(n1355), .B(n1356), .Z(n1353) );
  NAND U1187 ( .A(n1357), .B(n1358), .Z(n1356) );
  NANDN U1188 ( .A(A[173]), .B(B[173]), .Z(n1358) );
  AND U1189 ( .A(n1359), .B(n1360), .Z(n1357) );
  NANDN U1190 ( .A(A[172]), .B(B[172]), .Z(n1360) );
  NAND U1191 ( .A(n1361), .B(n1362), .Z(n1359) );
  NANDN U1192 ( .A(B[172]), .B(A[172]), .Z(n1362) );
  AND U1193 ( .A(n1363), .B(n1364), .Z(n1361) );
  NAND U1194 ( .A(n1365), .B(n1366), .Z(n1364) );
  NANDN U1195 ( .A(A[171]), .B(B[171]), .Z(n1366) );
  AND U1196 ( .A(n1367), .B(n1368), .Z(n1365) );
  NANDN U1197 ( .A(A[170]), .B(B[170]), .Z(n1368) );
  NAND U1198 ( .A(n1369), .B(n1370), .Z(n1367) );
  NANDN U1199 ( .A(B[170]), .B(A[170]), .Z(n1370) );
  AND U1200 ( .A(n1371), .B(n1372), .Z(n1369) );
  NAND U1201 ( .A(n1373), .B(n1374), .Z(n1372) );
  NANDN U1202 ( .A(A[169]), .B(B[169]), .Z(n1374) );
  AND U1203 ( .A(n1375), .B(n1376), .Z(n1373) );
  NANDN U1204 ( .A(A[168]), .B(B[168]), .Z(n1376) );
  NAND U1205 ( .A(n1377), .B(n1378), .Z(n1375) );
  NANDN U1206 ( .A(B[168]), .B(A[168]), .Z(n1378) );
  AND U1207 ( .A(n1379), .B(n1380), .Z(n1377) );
  NAND U1208 ( .A(n1381), .B(n1382), .Z(n1380) );
  NANDN U1209 ( .A(A[167]), .B(B[167]), .Z(n1382) );
  AND U1210 ( .A(n1383), .B(n1384), .Z(n1381) );
  NANDN U1211 ( .A(A[166]), .B(B[166]), .Z(n1384) );
  NAND U1212 ( .A(n1385), .B(n1386), .Z(n1383) );
  NANDN U1213 ( .A(B[166]), .B(A[166]), .Z(n1386) );
  AND U1214 ( .A(n1387), .B(n1388), .Z(n1385) );
  NAND U1215 ( .A(n1389), .B(n1390), .Z(n1388) );
  NANDN U1216 ( .A(A[165]), .B(B[165]), .Z(n1390) );
  AND U1217 ( .A(n1391), .B(n1392), .Z(n1389) );
  NANDN U1218 ( .A(A[164]), .B(B[164]), .Z(n1392) );
  NAND U1219 ( .A(n1393), .B(n1394), .Z(n1391) );
  NANDN U1220 ( .A(B[164]), .B(A[164]), .Z(n1394) );
  AND U1221 ( .A(n1395), .B(n1396), .Z(n1393) );
  NAND U1222 ( .A(n1397), .B(n1398), .Z(n1396) );
  NANDN U1223 ( .A(A[163]), .B(B[163]), .Z(n1398) );
  AND U1224 ( .A(n1399), .B(n1400), .Z(n1397) );
  NANDN U1225 ( .A(A[162]), .B(B[162]), .Z(n1400) );
  NAND U1226 ( .A(n1401), .B(n1402), .Z(n1399) );
  NANDN U1227 ( .A(B[162]), .B(A[162]), .Z(n1402) );
  AND U1228 ( .A(n1403), .B(n1404), .Z(n1401) );
  NAND U1229 ( .A(n1405), .B(n1406), .Z(n1404) );
  NANDN U1230 ( .A(A[161]), .B(B[161]), .Z(n1406) );
  AND U1231 ( .A(n1407), .B(n1408), .Z(n1405) );
  NANDN U1232 ( .A(A[160]), .B(B[160]), .Z(n1408) );
  NAND U1233 ( .A(n1409), .B(n1410), .Z(n1407) );
  NANDN U1234 ( .A(B[160]), .B(A[160]), .Z(n1410) );
  AND U1235 ( .A(n1411), .B(n1412), .Z(n1409) );
  NAND U1236 ( .A(n1413), .B(n1414), .Z(n1412) );
  NANDN U1237 ( .A(A[159]), .B(B[159]), .Z(n1414) );
  AND U1238 ( .A(n1415), .B(n1416), .Z(n1413) );
  NANDN U1239 ( .A(A[158]), .B(B[158]), .Z(n1416) );
  NAND U1240 ( .A(n1417), .B(n1418), .Z(n1415) );
  NANDN U1241 ( .A(B[158]), .B(A[158]), .Z(n1418) );
  AND U1242 ( .A(n1419), .B(n1420), .Z(n1417) );
  NAND U1243 ( .A(n1421), .B(n1422), .Z(n1420) );
  NANDN U1244 ( .A(A[157]), .B(B[157]), .Z(n1422) );
  AND U1245 ( .A(n1423), .B(n1424), .Z(n1421) );
  NANDN U1246 ( .A(A[156]), .B(B[156]), .Z(n1424) );
  NAND U1247 ( .A(n1425), .B(n1426), .Z(n1423) );
  NANDN U1248 ( .A(B[156]), .B(A[156]), .Z(n1426) );
  AND U1249 ( .A(n1427), .B(n1428), .Z(n1425) );
  NAND U1250 ( .A(n1429), .B(n1430), .Z(n1428) );
  NANDN U1251 ( .A(A[155]), .B(B[155]), .Z(n1430) );
  AND U1252 ( .A(n1431), .B(n1432), .Z(n1429) );
  NANDN U1253 ( .A(A[154]), .B(B[154]), .Z(n1432) );
  NAND U1254 ( .A(n1433), .B(n1434), .Z(n1431) );
  NANDN U1255 ( .A(B[154]), .B(A[154]), .Z(n1434) );
  AND U1256 ( .A(n1435), .B(n1436), .Z(n1433) );
  NAND U1257 ( .A(n1437), .B(n1438), .Z(n1436) );
  NANDN U1258 ( .A(A[153]), .B(B[153]), .Z(n1438) );
  AND U1259 ( .A(n1439), .B(n1440), .Z(n1437) );
  NANDN U1260 ( .A(A[152]), .B(B[152]), .Z(n1440) );
  NAND U1261 ( .A(n1441), .B(n1442), .Z(n1439) );
  NANDN U1262 ( .A(B[152]), .B(A[152]), .Z(n1442) );
  AND U1263 ( .A(n1443), .B(n1444), .Z(n1441) );
  NAND U1264 ( .A(n1445), .B(n1446), .Z(n1444) );
  NANDN U1265 ( .A(A[151]), .B(B[151]), .Z(n1446) );
  AND U1266 ( .A(n1447), .B(n1448), .Z(n1445) );
  NANDN U1267 ( .A(A[150]), .B(B[150]), .Z(n1448) );
  NAND U1268 ( .A(n1449), .B(n1450), .Z(n1447) );
  NANDN U1269 ( .A(B[150]), .B(A[150]), .Z(n1450) );
  AND U1270 ( .A(n1451), .B(n1452), .Z(n1449) );
  NAND U1271 ( .A(n1453), .B(n1454), .Z(n1452) );
  NANDN U1272 ( .A(A[149]), .B(B[149]), .Z(n1454) );
  AND U1273 ( .A(n1455), .B(n1456), .Z(n1453) );
  NANDN U1274 ( .A(A[148]), .B(B[148]), .Z(n1456) );
  NAND U1275 ( .A(n1457), .B(n1458), .Z(n1455) );
  NANDN U1276 ( .A(B[148]), .B(A[148]), .Z(n1458) );
  AND U1277 ( .A(n1459), .B(n1460), .Z(n1457) );
  NAND U1278 ( .A(n1461), .B(n1462), .Z(n1460) );
  NANDN U1279 ( .A(A[147]), .B(B[147]), .Z(n1462) );
  AND U1280 ( .A(n1463), .B(n1464), .Z(n1461) );
  NANDN U1281 ( .A(A[146]), .B(B[146]), .Z(n1464) );
  NAND U1282 ( .A(n1465), .B(n1466), .Z(n1463) );
  NANDN U1283 ( .A(B[146]), .B(A[146]), .Z(n1466) );
  AND U1284 ( .A(n1467), .B(n1468), .Z(n1465) );
  NAND U1285 ( .A(n1469), .B(n1470), .Z(n1468) );
  NANDN U1286 ( .A(A[145]), .B(B[145]), .Z(n1470) );
  AND U1287 ( .A(n1471), .B(n1472), .Z(n1469) );
  NANDN U1288 ( .A(A[144]), .B(B[144]), .Z(n1472) );
  NAND U1289 ( .A(n1473), .B(n1474), .Z(n1471) );
  NANDN U1290 ( .A(B[144]), .B(A[144]), .Z(n1474) );
  AND U1291 ( .A(n1475), .B(n1476), .Z(n1473) );
  NAND U1292 ( .A(n1477), .B(n1478), .Z(n1476) );
  NANDN U1293 ( .A(A[143]), .B(B[143]), .Z(n1478) );
  AND U1294 ( .A(n1479), .B(n1480), .Z(n1477) );
  NANDN U1295 ( .A(A[142]), .B(B[142]), .Z(n1480) );
  NAND U1296 ( .A(n1481), .B(n1482), .Z(n1479) );
  NANDN U1297 ( .A(B[142]), .B(A[142]), .Z(n1482) );
  AND U1298 ( .A(n1483), .B(n1484), .Z(n1481) );
  NAND U1299 ( .A(n1485), .B(n1486), .Z(n1484) );
  NANDN U1300 ( .A(A[141]), .B(B[141]), .Z(n1486) );
  AND U1301 ( .A(n1487), .B(n1488), .Z(n1485) );
  NANDN U1302 ( .A(A[140]), .B(B[140]), .Z(n1488) );
  NAND U1303 ( .A(n1489), .B(n1490), .Z(n1487) );
  NANDN U1304 ( .A(B[140]), .B(A[140]), .Z(n1490) );
  AND U1305 ( .A(n1491), .B(n1492), .Z(n1489) );
  NAND U1306 ( .A(n1493), .B(n1494), .Z(n1492) );
  NANDN U1307 ( .A(A[139]), .B(B[139]), .Z(n1494) );
  AND U1308 ( .A(n1495), .B(n1496), .Z(n1493) );
  NANDN U1309 ( .A(A[138]), .B(B[138]), .Z(n1496) );
  NAND U1310 ( .A(n1497), .B(n1498), .Z(n1495) );
  NANDN U1311 ( .A(B[138]), .B(A[138]), .Z(n1498) );
  AND U1312 ( .A(n1499), .B(n1500), .Z(n1497) );
  NAND U1313 ( .A(n1501), .B(n1502), .Z(n1500) );
  NANDN U1314 ( .A(A[137]), .B(B[137]), .Z(n1502) );
  AND U1315 ( .A(n1503), .B(n1504), .Z(n1501) );
  NANDN U1316 ( .A(A[136]), .B(B[136]), .Z(n1504) );
  NAND U1317 ( .A(n1505), .B(n1506), .Z(n1503) );
  NANDN U1318 ( .A(B[136]), .B(A[136]), .Z(n1506) );
  AND U1319 ( .A(n1507), .B(n1508), .Z(n1505) );
  NAND U1320 ( .A(n1509), .B(n1510), .Z(n1508) );
  NANDN U1321 ( .A(A[135]), .B(B[135]), .Z(n1510) );
  AND U1322 ( .A(n1511), .B(n1512), .Z(n1509) );
  NANDN U1323 ( .A(A[134]), .B(B[134]), .Z(n1512) );
  NAND U1324 ( .A(n1513), .B(n1514), .Z(n1511) );
  NANDN U1325 ( .A(B[134]), .B(A[134]), .Z(n1514) );
  AND U1326 ( .A(n1515), .B(n1516), .Z(n1513) );
  NAND U1327 ( .A(n1517), .B(n1518), .Z(n1516) );
  NANDN U1328 ( .A(A[133]), .B(B[133]), .Z(n1518) );
  AND U1329 ( .A(n1519), .B(n1520), .Z(n1517) );
  NANDN U1330 ( .A(A[132]), .B(B[132]), .Z(n1520) );
  NAND U1331 ( .A(n1521), .B(n1522), .Z(n1519) );
  NANDN U1332 ( .A(B[132]), .B(A[132]), .Z(n1522) );
  AND U1333 ( .A(n1523), .B(n1524), .Z(n1521) );
  NAND U1334 ( .A(n1525), .B(n1526), .Z(n1524) );
  NANDN U1335 ( .A(A[131]), .B(B[131]), .Z(n1526) );
  AND U1336 ( .A(n1527), .B(n1528), .Z(n1525) );
  NANDN U1337 ( .A(A[130]), .B(B[130]), .Z(n1528) );
  NAND U1338 ( .A(n1529), .B(n1530), .Z(n1527) );
  NANDN U1339 ( .A(B[130]), .B(A[130]), .Z(n1530) );
  AND U1340 ( .A(n1531), .B(n1532), .Z(n1529) );
  NAND U1341 ( .A(n1533), .B(n1534), .Z(n1532) );
  NANDN U1342 ( .A(A[129]), .B(B[129]), .Z(n1534) );
  AND U1343 ( .A(n1535), .B(n1536), .Z(n1533) );
  NANDN U1344 ( .A(A[128]), .B(B[128]), .Z(n1536) );
  NAND U1345 ( .A(n1537), .B(n1538), .Z(n1535) );
  NANDN U1346 ( .A(B[128]), .B(A[128]), .Z(n1538) );
  AND U1347 ( .A(n1539), .B(n1540), .Z(n1537) );
  NAND U1348 ( .A(n1541), .B(n1542), .Z(n1540) );
  NANDN U1349 ( .A(A[127]), .B(B[127]), .Z(n1542) );
  AND U1350 ( .A(n1543), .B(n1544), .Z(n1541) );
  NANDN U1351 ( .A(A[126]), .B(B[126]), .Z(n1544) );
  NAND U1352 ( .A(n1545), .B(n1546), .Z(n1543) );
  NANDN U1353 ( .A(B[126]), .B(A[126]), .Z(n1546) );
  AND U1354 ( .A(n1547), .B(n1548), .Z(n1545) );
  NAND U1355 ( .A(n1549), .B(n1550), .Z(n1548) );
  NANDN U1356 ( .A(A[125]), .B(B[125]), .Z(n1550) );
  AND U1357 ( .A(n1551), .B(n1552), .Z(n1549) );
  NANDN U1358 ( .A(A[124]), .B(B[124]), .Z(n1552) );
  NAND U1359 ( .A(n1553), .B(n1554), .Z(n1551) );
  NANDN U1360 ( .A(B[124]), .B(A[124]), .Z(n1554) );
  AND U1361 ( .A(n1555), .B(n1556), .Z(n1553) );
  NAND U1362 ( .A(n1557), .B(n1558), .Z(n1556) );
  NANDN U1363 ( .A(A[123]), .B(B[123]), .Z(n1558) );
  AND U1364 ( .A(n1559), .B(n1560), .Z(n1557) );
  NANDN U1365 ( .A(A[122]), .B(B[122]), .Z(n1560) );
  NAND U1366 ( .A(n1561), .B(n1562), .Z(n1559) );
  NANDN U1367 ( .A(B[122]), .B(A[122]), .Z(n1562) );
  AND U1368 ( .A(n1563), .B(n1564), .Z(n1561) );
  NAND U1369 ( .A(n1565), .B(n1566), .Z(n1564) );
  NANDN U1370 ( .A(A[121]), .B(B[121]), .Z(n1566) );
  AND U1371 ( .A(n1567), .B(n1568), .Z(n1565) );
  NANDN U1372 ( .A(A[120]), .B(B[120]), .Z(n1568) );
  NAND U1373 ( .A(n1569), .B(n1570), .Z(n1567) );
  NANDN U1374 ( .A(B[120]), .B(A[120]), .Z(n1570) );
  AND U1375 ( .A(n1571), .B(n1572), .Z(n1569) );
  NAND U1376 ( .A(n1573), .B(n1574), .Z(n1572) );
  NANDN U1377 ( .A(A[119]), .B(B[119]), .Z(n1574) );
  AND U1378 ( .A(n1575), .B(n1576), .Z(n1573) );
  NANDN U1379 ( .A(A[118]), .B(B[118]), .Z(n1576) );
  NAND U1380 ( .A(n1577), .B(n1578), .Z(n1575) );
  NANDN U1381 ( .A(B[118]), .B(A[118]), .Z(n1578) );
  AND U1382 ( .A(n1579), .B(n1580), .Z(n1577) );
  NAND U1383 ( .A(n1581), .B(n1582), .Z(n1580) );
  NANDN U1384 ( .A(A[117]), .B(B[117]), .Z(n1582) );
  AND U1385 ( .A(n1583), .B(n1584), .Z(n1581) );
  NANDN U1386 ( .A(A[116]), .B(B[116]), .Z(n1584) );
  NAND U1387 ( .A(n1585), .B(n1586), .Z(n1583) );
  NANDN U1388 ( .A(B[116]), .B(A[116]), .Z(n1586) );
  AND U1389 ( .A(n1587), .B(n1588), .Z(n1585) );
  NAND U1390 ( .A(n1589), .B(n1590), .Z(n1588) );
  NANDN U1391 ( .A(A[115]), .B(B[115]), .Z(n1590) );
  AND U1392 ( .A(n1591), .B(n1592), .Z(n1589) );
  NANDN U1393 ( .A(A[114]), .B(B[114]), .Z(n1592) );
  NAND U1394 ( .A(n1593), .B(n1594), .Z(n1591) );
  NANDN U1395 ( .A(B[114]), .B(A[114]), .Z(n1594) );
  AND U1396 ( .A(n1595), .B(n1596), .Z(n1593) );
  NAND U1397 ( .A(n1597), .B(n1598), .Z(n1596) );
  NANDN U1398 ( .A(A[113]), .B(B[113]), .Z(n1598) );
  AND U1399 ( .A(n1599), .B(n1600), .Z(n1597) );
  NANDN U1400 ( .A(A[112]), .B(B[112]), .Z(n1600) );
  NAND U1401 ( .A(n1601), .B(n1602), .Z(n1599) );
  NANDN U1402 ( .A(B[112]), .B(A[112]), .Z(n1602) );
  AND U1403 ( .A(n1603), .B(n1604), .Z(n1601) );
  NAND U1404 ( .A(n1605), .B(n1606), .Z(n1604) );
  NANDN U1405 ( .A(A[111]), .B(B[111]), .Z(n1606) );
  AND U1406 ( .A(n1607), .B(n1608), .Z(n1605) );
  NANDN U1407 ( .A(A[110]), .B(B[110]), .Z(n1608) );
  NAND U1408 ( .A(n1609), .B(n1610), .Z(n1607) );
  NANDN U1409 ( .A(B[110]), .B(A[110]), .Z(n1610) );
  AND U1410 ( .A(n1611), .B(n1612), .Z(n1609) );
  NAND U1411 ( .A(n1613), .B(n1614), .Z(n1612) );
  NANDN U1412 ( .A(A[109]), .B(B[109]), .Z(n1614) );
  AND U1413 ( .A(n1615), .B(n1616), .Z(n1613) );
  NANDN U1414 ( .A(A[108]), .B(B[108]), .Z(n1616) );
  NAND U1415 ( .A(n1617), .B(n1618), .Z(n1615) );
  NANDN U1416 ( .A(B[108]), .B(A[108]), .Z(n1618) );
  AND U1417 ( .A(n1619), .B(n1620), .Z(n1617) );
  NAND U1418 ( .A(n1621), .B(n1622), .Z(n1620) );
  NANDN U1419 ( .A(A[107]), .B(B[107]), .Z(n1622) );
  AND U1420 ( .A(n1623), .B(n1624), .Z(n1621) );
  NANDN U1421 ( .A(A[106]), .B(B[106]), .Z(n1624) );
  NAND U1422 ( .A(n1625), .B(n1626), .Z(n1623) );
  NANDN U1423 ( .A(B[106]), .B(A[106]), .Z(n1626) );
  AND U1424 ( .A(n1627), .B(n1628), .Z(n1625) );
  NAND U1425 ( .A(n1629), .B(n1630), .Z(n1628) );
  NANDN U1426 ( .A(A[105]), .B(B[105]), .Z(n1630) );
  AND U1427 ( .A(n1631), .B(n1632), .Z(n1629) );
  NANDN U1428 ( .A(A[104]), .B(B[104]), .Z(n1632) );
  NAND U1429 ( .A(n1633), .B(n1634), .Z(n1631) );
  NANDN U1430 ( .A(B[104]), .B(A[104]), .Z(n1634) );
  AND U1431 ( .A(n1635), .B(n1636), .Z(n1633) );
  NAND U1432 ( .A(n1637), .B(n1638), .Z(n1636) );
  NANDN U1433 ( .A(A[103]), .B(B[103]), .Z(n1638) );
  AND U1434 ( .A(n1639), .B(n1640), .Z(n1637) );
  NANDN U1435 ( .A(A[102]), .B(B[102]), .Z(n1640) );
  NAND U1436 ( .A(n1641), .B(n1642), .Z(n1639) );
  NANDN U1437 ( .A(B[102]), .B(A[102]), .Z(n1642) );
  AND U1438 ( .A(n1643), .B(n1644), .Z(n1641) );
  NAND U1439 ( .A(n1645), .B(n1646), .Z(n1644) );
  NANDN U1440 ( .A(A[101]), .B(B[101]), .Z(n1646) );
  AND U1441 ( .A(n1647), .B(n1648), .Z(n1645) );
  NANDN U1442 ( .A(A[100]), .B(B[100]), .Z(n1648) );
  NAND U1443 ( .A(n1649), .B(n1650), .Z(n1647) );
  NANDN U1444 ( .A(B[99]), .B(A[99]), .Z(n1650) );
  AND U1445 ( .A(n1651), .B(n1652), .Z(n1649) );
  NAND U1446 ( .A(n1653), .B(n1654), .Z(n1652) );
  NANDN U1447 ( .A(A[99]), .B(B[99]), .Z(n1654) );
  AND U1448 ( .A(n1655), .B(n1656), .Z(n1653) );
  NANDN U1449 ( .A(A[98]), .B(B[98]), .Z(n1656) );
  NAND U1450 ( .A(n1657), .B(n1658), .Z(n1655) );
  NANDN U1451 ( .A(B[98]), .B(A[98]), .Z(n1658) );
  AND U1452 ( .A(n1659), .B(n1660), .Z(n1657) );
  NAND U1453 ( .A(n1661), .B(n1662), .Z(n1660) );
  NANDN U1454 ( .A(A[97]), .B(B[97]), .Z(n1662) );
  AND U1455 ( .A(n1663), .B(n1664), .Z(n1661) );
  NANDN U1456 ( .A(A[96]), .B(B[96]), .Z(n1664) );
  NAND U1457 ( .A(n1665), .B(n1666), .Z(n1663) );
  NANDN U1458 ( .A(B[96]), .B(A[96]), .Z(n1666) );
  AND U1459 ( .A(n1667), .B(n1668), .Z(n1665) );
  NAND U1460 ( .A(n1669), .B(n1670), .Z(n1668) );
  NANDN U1461 ( .A(A[95]), .B(B[95]), .Z(n1670) );
  AND U1462 ( .A(n1671), .B(n1672), .Z(n1669) );
  NANDN U1463 ( .A(A[94]), .B(B[94]), .Z(n1672) );
  NAND U1464 ( .A(n1673), .B(n1674), .Z(n1671) );
  NANDN U1465 ( .A(B[94]), .B(A[94]), .Z(n1674) );
  AND U1466 ( .A(n1675), .B(n1676), .Z(n1673) );
  NAND U1467 ( .A(n1677), .B(n1678), .Z(n1676) );
  NANDN U1468 ( .A(A[93]), .B(B[93]), .Z(n1678) );
  AND U1469 ( .A(n1679), .B(n1680), .Z(n1677) );
  NANDN U1470 ( .A(A[92]), .B(B[92]), .Z(n1680) );
  NAND U1471 ( .A(n1681), .B(n1682), .Z(n1679) );
  NANDN U1472 ( .A(B[92]), .B(A[92]), .Z(n1682) );
  AND U1473 ( .A(n1683), .B(n1684), .Z(n1681) );
  NAND U1474 ( .A(n1685), .B(n1686), .Z(n1684) );
  NANDN U1475 ( .A(A[91]), .B(B[91]), .Z(n1686) );
  AND U1476 ( .A(n1687), .B(n1688), .Z(n1685) );
  NANDN U1477 ( .A(A[90]), .B(B[90]), .Z(n1688) );
  NAND U1478 ( .A(n1689), .B(n1690), .Z(n1687) );
  NANDN U1479 ( .A(B[90]), .B(A[90]), .Z(n1690) );
  AND U1480 ( .A(n1691), .B(n1692), .Z(n1689) );
  NAND U1481 ( .A(n1693), .B(n1694), .Z(n1692) );
  NANDN U1482 ( .A(A[89]), .B(B[89]), .Z(n1694) );
  AND U1483 ( .A(n1695), .B(n1696), .Z(n1693) );
  NANDN U1484 ( .A(A[88]), .B(B[88]), .Z(n1696) );
  NAND U1485 ( .A(n1697), .B(n1698), .Z(n1695) );
  NANDN U1486 ( .A(B[88]), .B(A[88]), .Z(n1698) );
  AND U1487 ( .A(n1699), .B(n1700), .Z(n1697) );
  NAND U1488 ( .A(n1701), .B(n1702), .Z(n1700) );
  NANDN U1489 ( .A(A[87]), .B(B[87]), .Z(n1702) );
  AND U1490 ( .A(n1703), .B(n1704), .Z(n1701) );
  NANDN U1491 ( .A(A[86]), .B(B[86]), .Z(n1704) );
  NAND U1492 ( .A(n1705), .B(n1706), .Z(n1703) );
  NANDN U1493 ( .A(B[86]), .B(A[86]), .Z(n1706) );
  AND U1494 ( .A(n1707), .B(n1708), .Z(n1705) );
  NAND U1495 ( .A(n1709), .B(n1710), .Z(n1708) );
  NANDN U1496 ( .A(A[85]), .B(B[85]), .Z(n1710) );
  AND U1497 ( .A(n1711), .B(n1712), .Z(n1709) );
  NANDN U1498 ( .A(A[84]), .B(B[84]), .Z(n1712) );
  NAND U1499 ( .A(n1713), .B(n1714), .Z(n1711) );
  NANDN U1500 ( .A(B[84]), .B(A[84]), .Z(n1714) );
  AND U1501 ( .A(n1715), .B(n1716), .Z(n1713) );
  NAND U1502 ( .A(n1717), .B(n1718), .Z(n1716) );
  NANDN U1503 ( .A(A[83]), .B(B[83]), .Z(n1718) );
  AND U1504 ( .A(n1719), .B(n1720), .Z(n1717) );
  NANDN U1505 ( .A(A[82]), .B(B[82]), .Z(n1720) );
  NAND U1506 ( .A(n1721), .B(n1722), .Z(n1719) );
  NANDN U1507 ( .A(B[82]), .B(A[82]), .Z(n1722) );
  AND U1508 ( .A(n1723), .B(n1724), .Z(n1721) );
  NAND U1509 ( .A(n1725), .B(n1726), .Z(n1724) );
  NANDN U1510 ( .A(A[81]), .B(B[81]), .Z(n1726) );
  AND U1511 ( .A(n1727), .B(n1728), .Z(n1725) );
  NANDN U1512 ( .A(A[80]), .B(B[80]), .Z(n1728) );
  NAND U1513 ( .A(n1729), .B(n1730), .Z(n1727) );
  NANDN U1514 ( .A(B[80]), .B(A[80]), .Z(n1730) );
  AND U1515 ( .A(n1731), .B(n1732), .Z(n1729) );
  NAND U1516 ( .A(n1733), .B(n1734), .Z(n1732) );
  NANDN U1517 ( .A(A[79]), .B(B[79]), .Z(n1734) );
  AND U1518 ( .A(n1735), .B(n1736), .Z(n1733) );
  NANDN U1519 ( .A(A[78]), .B(B[78]), .Z(n1736) );
  NAND U1520 ( .A(n1737), .B(n1738), .Z(n1735) );
  NANDN U1521 ( .A(B[78]), .B(A[78]), .Z(n1738) );
  AND U1522 ( .A(n1739), .B(n1740), .Z(n1737) );
  NAND U1523 ( .A(n1741), .B(n1742), .Z(n1740) );
  NANDN U1524 ( .A(A[77]), .B(B[77]), .Z(n1742) );
  AND U1525 ( .A(n1743), .B(n1744), .Z(n1741) );
  NANDN U1526 ( .A(A[76]), .B(B[76]), .Z(n1744) );
  NAND U1527 ( .A(n1745), .B(n1746), .Z(n1743) );
  NANDN U1528 ( .A(B[76]), .B(A[76]), .Z(n1746) );
  AND U1529 ( .A(n1747), .B(n1748), .Z(n1745) );
  NAND U1530 ( .A(n1749), .B(n1750), .Z(n1748) );
  NANDN U1531 ( .A(A[75]), .B(B[75]), .Z(n1750) );
  AND U1532 ( .A(n1751), .B(n1752), .Z(n1749) );
  NANDN U1533 ( .A(A[74]), .B(B[74]), .Z(n1752) );
  NAND U1534 ( .A(n1753), .B(n1754), .Z(n1751) );
  NANDN U1535 ( .A(B[74]), .B(A[74]), .Z(n1754) );
  AND U1536 ( .A(n1755), .B(n1756), .Z(n1753) );
  NAND U1537 ( .A(n1757), .B(n1758), .Z(n1756) );
  NANDN U1538 ( .A(A[73]), .B(B[73]), .Z(n1758) );
  AND U1539 ( .A(n1759), .B(n1760), .Z(n1757) );
  NANDN U1540 ( .A(A[72]), .B(B[72]), .Z(n1760) );
  NAND U1541 ( .A(n1761), .B(n1762), .Z(n1759) );
  NANDN U1542 ( .A(B[72]), .B(A[72]), .Z(n1762) );
  AND U1543 ( .A(n1763), .B(n1764), .Z(n1761) );
  NAND U1544 ( .A(n1765), .B(n1766), .Z(n1764) );
  NANDN U1545 ( .A(A[71]), .B(B[71]), .Z(n1766) );
  AND U1546 ( .A(n1767), .B(n1768), .Z(n1765) );
  NANDN U1547 ( .A(A[70]), .B(B[70]), .Z(n1768) );
  NAND U1548 ( .A(n1769), .B(n1770), .Z(n1767) );
  NANDN U1549 ( .A(B[70]), .B(A[70]), .Z(n1770) );
  AND U1550 ( .A(n1771), .B(n1772), .Z(n1769) );
  NAND U1551 ( .A(n1773), .B(n1774), .Z(n1772) );
  NANDN U1552 ( .A(A[69]), .B(B[69]), .Z(n1774) );
  AND U1553 ( .A(n1775), .B(n1776), .Z(n1773) );
  NANDN U1554 ( .A(A[68]), .B(B[68]), .Z(n1776) );
  NAND U1555 ( .A(n1777), .B(n1778), .Z(n1775) );
  NANDN U1556 ( .A(B[68]), .B(A[68]), .Z(n1778) );
  AND U1557 ( .A(n1779), .B(n1780), .Z(n1777) );
  NAND U1558 ( .A(n1781), .B(n1782), .Z(n1780) );
  NANDN U1559 ( .A(A[67]), .B(B[67]), .Z(n1782) );
  AND U1560 ( .A(n1783), .B(n1784), .Z(n1781) );
  NANDN U1561 ( .A(A[66]), .B(B[66]), .Z(n1784) );
  NAND U1562 ( .A(n1785), .B(n1786), .Z(n1783) );
  NANDN U1563 ( .A(B[66]), .B(A[66]), .Z(n1786) );
  AND U1564 ( .A(n1787), .B(n1788), .Z(n1785) );
  NAND U1565 ( .A(n1789), .B(n1790), .Z(n1788) );
  NANDN U1566 ( .A(A[65]), .B(B[65]), .Z(n1790) );
  AND U1567 ( .A(n1791), .B(n1792), .Z(n1789) );
  NANDN U1568 ( .A(A[64]), .B(B[64]), .Z(n1792) );
  NAND U1569 ( .A(n1793), .B(n1794), .Z(n1791) );
  NANDN U1570 ( .A(B[64]), .B(A[64]), .Z(n1794) );
  AND U1571 ( .A(n1795), .B(n1796), .Z(n1793) );
  NAND U1572 ( .A(n1797), .B(n1798), .Z(n1796) );
  NANDN U1573 ( .A(A[63]), .B(B[63]), .Z(n1798) );
  AND U1574 ( .A(n1799), .B(n1800), .Z(n1797) );
  NANDN U1575 ( .A(A[62]), .B(B[62]), .Z(n1800) );
  NAND U1576 ( .A(n1801), .B(n1802), .Z(n1799) );
  NANDN U1577 ( .A(B[62]), .B(A[62]), .Z(n1802) );
  AND U1578 ( .A(n1803), .B(n1804), .Z(n1801) );
  NAND U1579 ( .A(n1805), .B(n1806), .Z(n1804) );
  NANDN U1580 ( .A(A[61]), .B(B[61]), .Z(n1806) );
  AND U1581 ( .A(n1807), .B(n1808), .Z(n1805) );
  NANDN U1582 ( .A(A[60]), .B(B[60]), .Z(n1808) );
  NAND U1583 ( .A(n1809), .B(n1810), .Z(n1807) );
  NANDN U1584 ( .A(B[60]), .B(A[60]), .Z(n1810) );
  AND U1585 ( .A(n1811), .B(n1812), .Z(n1809) );
  NAND U1586 ( .A(n1813), .B(n1814), .Z(n1812) );
  NANDN U1587 ( .A(A[59]), .B(B[59]), .Z(n1814) );
  AND U1588 ( .A(n1815), .B(n1816), .Z(n1813) );
  NANDN U1589 ( .A(A[58]), .B(B[58]), .Z(n1816) );
  NAND U1590 ( .A(n1817), .B(n1818), .Z(n1815) );
  NANDN U1591 ( .A(B[58]), .B(A[58]), .Z(n1818) );
  AND U1592 ( .A(n1819), .B(n1820), .Z(n1817) );
  NAND U1593 ( .A(n1821), .B(n1822), .Z(n1820) );
  NANDN U1594 ( .A(A[57]), .B(B[57]), .Z(n1822) );
  AND U1595 ( .A(n1823), .B(n1824), .Z(n1821) );
  NANDN U1596 ( .A(A[56]), .B(B[56]), .Z(n1824) );
  NAND U1597 ( .A(n1825), .B(n1826), .Z(n1823) );
  NANDN U1598 ( .A(B[56]), .B(A[56]), .Z(n1826) );
  AND U1599 ( .A(n1827), .B(n1828), .Z(n1825) );
  NAND U1600 ( .A(n1829), .B(n1830), .Z(n1828) );
  NANDN U1601 ( .A(A[55]), .B(B[55]), .Z(n1830) );
  AND U1602 ( .A(n1831), .B(n1832), .Z(n1829) );
  NANDN U1603 ( .A(A[54]), .B(B[54]), .Z(n1832) );
  NAND U1604 ( .A(n1833), .B(n1834), .Z(n1831) );
  NANDN U1605 ( .A(B[54]), .B(A[54]), .Z(n1834) );
  AND U1606 ( .A(n1835), .B(n1836), .Z(n1833) );
  NAND U1607 ( .A(n1837), .B(n1838), .Z(n1836) );
  NANDN U1608 ( .A(A[53]), .B(B[53]), .Z(n1838) );
  AND U1609 ( .A(n1839), .B(n1840), .Z(n1837) );
  NANDN U1610 ( .A(A[52]), .B(B[52]), .Z(n1840) );
  NAND U1611 ( .A(n1841), .B(n1842), .Z(n1839) );
  NANDN U1612 ( .A(B[52]), .B(A[52]), .Z(n1842) );
  AND U1613 ( .A(n1843), .B(n1844), .Z(n1841) );
  NAND U1614 ( .A(n1845), .B(n1846), .Z(n1844) );
  NANDN U1615 ( .A(A[51]), .B(B[51]), .Z(n1846) );
  AND U1616 ( .A(n1847), .B(n1848), .Z(n1845) );
  NANDN U1617 ( .A(A[50]), .B(B[50]), .Z(n1848) );
  NAND U1618 ( .A(n1849), .B(n1850), .Z(n1847) );
  NANDN U1619 ( .A(B[50]), .B(A[50]), .Z(n1850) );
  AND U1620 ( .A(n1851), .B(n1852), .Z(n1849) );
  NAND U1621 ( .A(n1853), .B(n1854), .Z(n1852) );
  NANDN U1622 ( .A(A[49]), .B(B[49]), .Z(n1854) );
  AND U1623 ( .A(n1855), .B(n1856), .Z(n1853) );
  NANDN U1624 ( .A(A[48]), .B(B[48]), .Z(n1856) );
  NAND U1625 ( .A(n1857), .B(n1858), .Z(n1855) );
  NANDN U1626 ( .A(B[48]), .B(A[48]), .Z(n1858) );
  AND U1627 ( .A(n1859), .B(n1860), .Z(n1857) );
  NAND U1628 ( .A(n1861), .B(n1862), .Z(n1860) );
  NANDN U1629 ( .A(A[47]), .B(B[47]), .Z(n1862) );
  AND U1630 ( .A(n1863), .B(n1864), .Z(n1861) );
  NANDN U1631 ( .A(A[46]), .B(B[46]), .Z(n1864) );
  NAND U1632 ( .A(n1865), .B(n1866), .Z(n1863) );
  NANDN U1633 ( .A(B[46]), .B(A[46]), .Z(n1866) );
  AND U1634 ( .A(n1867), .B(n1868), .Z(n1865) );
  NAND U1635 ( .A(n1869), .B(n1870), .Z(n1868) );
  NANDN U1636 ( .A(A[45]), .B(B[45]), .Z(n1870) );
  AND U1637 ( .A(n1871), .B(n1872), .Z(n1869) );
  NANDN U1638 ( .A(A[44]), .B(B[44]), .Z(n1872) );
  NAND U1639 ( .A(n1873), .B(n1874), .Z(n1871) );
  NANDN U1640 ( .A(B[44]), .B(A[44]), .Z(n1874) );
  AND U1641 ( .A(n1875), .B(n1876), .Z(n1873) );
  NAND U1642 ( .A(n1877), .B(n1878), .Z(n1876) );
  NANDN U1643 ( .A(A[43]), .B(B[43]), .Z(n1878) );
  AND U1644 ( .A(n1879), .B(n1880), .Z(n1877) );
  NANDN U1645 ( .A(A[42]), .B(B[42]), .Z(n1880) );
  NAND U1646 ( .A(n1881), .B(n1882), .Z(n1879) );
  NANDN U1647 ( .A(B[42]), .B(A[42]), .Z(n1882) );
  AND U1648 ( .A(n1883), .B(n1884), .Z(n1881) );
  NAND U1649 ( .A(n1885), .B(n1886), .Z(n1884) );
  NANDN U1650 ( .A(A[41]), .B(B[41]), .Z(n1886) );
  AND U1651 ( .A(n1887), .B(n1888), .Z(n1885) );
  NANDN U1652 ( .A(A[40]), .B(B[40]), .Z(n1888) );
  NAND U1653 ( .A(n1889), .B(n1890), .Z(n1887) );
  NANDN U1654 ( .A(B[40]), .B(A[40]), .Z(n1890) );
  AND U1655 ( .A(n1891), .B(n1892), .Z(n1889) );
  NAND U1656 ( .A(n1893), .B(n1894), .Z(n1892) );
  NANDN U1657 ( .A(A[39]), .B(B[39]), .Z(n1894) );
  AND U1658 ( .A(n1895), .B(n1896), .Z(n1893) );
  NANDN U1659 ( .A(A[38]), .B(B[38]), .Z(n1896) );
  NAND U1660 ( .A(n1897), .B(n1898), .Z(n1895) );
  NANDN U1661 ( .A(B[38]), .B(A[38]), .Z(n1898) );
  AND U1662 ( .A(n1899), .B(n1900), .Z(n1897) );
  NAND U1663 ( .A(n1901), .B(n1902), .Z(n1900) );
  NANDN U1664 ( .A(A[37]), .B(B[37]), .Z(n1902) );
  AND U1665 ( .A(n1903), .B(n1904), .Z(n1901) );
  NANDN U1666 ( .A(A[36]), .B(B[36]), .Z(n1904) );
  NAND U1667 ( .A(n1905), .B(n1906), .Z(n1903) );
  NANDN U1668 ( .A(B[36]), .B(A[36]), .Z(n1906) );
  AND U1669 ( .A(n1907), .B(n1908), .Z(n1905) );
  NAND U1670 ( .A(n1909), .B(n1910), .Z(n1908) );
  NANDN U1671 ( .A(A[35]), .B(B[35]), .Z(n1910) );
  AND U1672 ( .A(n1911), .B(n1912), .Z(n1909) );
  NANDN U1673 ( .A(A[34]), .B(B[34]), .Z(n1912) );
  NAND U1674 ( .A(n1913), .B(n1914), .Z(n1911) );
  NANDN U1675 ( .A(B[34]), .B(A[34]), .Z(n1914) );
  AND U1676 ( .A(n1915), .B(n1916), .Z(n1913) );
  NAND U1677 ( .A(n1917), .B(n1918), .Z(n1916) );
  NANDN U1678 ( .A(A[33]), .B(B[33]), .Z(n1918) );
  AND U1679 ( .A(n1919), .B(n1920), .Z(n1917) );
  NANDN U1680 ( .A(A[32]), .B(B[32]), .Z(n1920) );
  NAND U1681 ( .A(n1921), .B(n1922), .Z(n1919) );
  NANDN U1682 ( .A(B[32]), .B(A[32]), .Z(n1922) );
  AND U1683 ( .A(n1923), .B(n1924), .Z(n1921) );
  NAND U1684 ( .A(n1925), .B(n1926), .Z(n1924) );
  NANDN U1685 ( .A(A[31]), .B(B[31]), .Z(n1926) );
  AND U1686 ( .A(n1927), .B(n1928), .Z(n1925) );
  NANDN U1687 ( .A(A[30]), .B(B[30]), .Z(n1928) );
  NAND U1688 ( .A(n1929), .B(n1930), .Z(n1927) );
  NANDN U1689 ( .A(B[30]), .B(A[30]), .Z(n1930) );
  AND U1690 ( .A(n1931), .B(n1932), .Z(n1929) );
  NAND U1691 ( .A(n1933), .B(n1934), .Z(n1932) );
  NANDN U1692 ( .A(A[29]), .B(B[29]), .Z(n1934) );
  AND U1693 ( .A(n1935), .B(n1936), .Z(n1933) );
  NANDN U1694 ( .A(A[28]), .B(B[28]), .Z(n1936) );
  NAND U1695 ( .A(n1937), .B(n1938), .Z(n1935) );
  NANDN U1696 ( .A(B[28]), .B(A[28]), .Z(n1938) );
  AND U1697 ( .A(n1939), .B(n1940), .Z(n1937) );
  NAND U1698 ( .A(n1941), .B(n1942), .Z(n1940) );
  NANDN U1699 ( .A(A[27]), .B(B[27]), .Z(n1942) );
  AND U1700 ( .A(n1943), .B(n1944), .Z(n1941) );
  NANDN U1701 ( .A(A[26]), .B(B[26]), .Z(n1944) );
  NAND U1702 ( .A(n1945), .B(n1946), .Z(n1943) );
  NANDN U1703 ( .A(B[26]), .B(A[26]), .Z(n1946) );
  AND U1704 ( .A(n1947), .B(n1948), .Z(n1945) );
  NAND U1705 ( .A(n1949), .B(n1950), .Z(n1948) );
  NANDN U1706 ( .A(A[25]), .B(B[25]), .Z(n1950) );
  AND U1707 ( .A(n1951), .B(n1952), .Z(n1949) );
  NANDN U1708 ( .A(A[24]), .B(B[24]), .Z(n1952) );
  NAND U1709 ( .A(n1953), .B(n1954), .Z(n1951) );
  NANDN U1710 ( .A(B[24]), .B(A[24]), .Z(n1954) );
  AND U1711 ( .A(n1955), .B(n1956), .Z(n1953) );
  NAND U1712 ( .A(n1957), .B(n1958), .Z(n1956) );
  NANDN U1713 ( .A(A[23]), .B(B[23]), .Z(n1958) );
  AND U1714 ( .A(n1959), .B(n1960), .Z(n1957) );
  NANDN U1715 ( .A(A[22]), .B(B[22]), .Z(n1960) );
  NAND U1716 ( .A(n1961), .B(n1962), .Z(n1959) );
  NANDN U1717 ( .A(B[22]), .B(A[22]), .Z(n1962) );
  AND U1718 ( .A(n1963), .B(n1964), .Z(n1961) );
  NAND U1719 ( .A(n1965), .B(n1966), .Z(n1964) );
  NANDN U1720 ( .A(A[21]), .B(B[21]), .Z(n1966) );
  AND U1721 ( .A(n1967), .B(n1968), .Z(n1965) );
  NANDN U1722 ( .A(A[20]), .B(B[20]), .Z(n1968) );
  NAND U1723 ( .A(n1969), .B(n1970), .Z(n1967) );
  NANDN U1724 ( .A(B[20]), .B(A[20]), .Z(n1970) );
  AND U1725 ( .A(n1971), .B(n1972), .Z(n1969) );
  NAND U1726 ( .A(n1973), .B(n1974), .Z(n1972) );
  NANDN U1727 ( .A(A[19]), .B(B[19]), .Z(n1974) );
  AND U1728 ( .A(n1975), .B(n1976), .Z(n1973) );
  NANDN U1729 ( .A(A[18]), .B(B[18]), .Z(n1976) );
  NAND U1730 ( .A(n1977), .B(n1978), .Z(n1975) );
  NANDN U1731 ( .A(B[18]), .B(A[18]), .Z(n1978) );
  AND U1732 ( .A(n1979), .B(n1980), .Z(n1977) );
  NAND U1733 ( .A(n1981), .B(n1982), .Z(n1980) );
  NANDN U1734 ( .A(A[17]), .B(B[17]), .Z(n1982) );
  AND U1735 ( .A(n1983), .B(n1984), .Z(n1981) );
  NANDN U1736 ( .A(A[16]), .B(B[16]), .Z(n1984) );
  NAND U1737 ( .A(n1985), .B(n1986), .Z(n1983) );
  NANDN U1738 ( .A(B[16]), .B(A[16]), .Z(n1986) );
  AND U1739 ( .A(n1987), .B(n1988), .Z(n1985) );
  NAND U1740 ( .A(n1989), .B(n1990), .Z(n1988) );
  NANDN U1741 ( .A(A[15]), .B(B[15]), .Z(n1990) );
  AND U1742 ( .A(n1991), .B(n1992), .Z(n1989) );
  NANDN U1743 ( .A(A[14]), .B(B[14]), .Z(n1992) );
  NAND U1744 ( .A(n1993), .B(n1994), .Z(n1991) );
  NANDN U1745 ( .A(B[14]), .B(A[14]), .Z(n1994) );
  AND U1746 ( .A(n1995), .B(n1996), .Z(n1993) );
  NAND U1747 ( .A(n1997), .B(n1998), .Z(n1996) );
  NANDN U1748 ( .A(A[13]), .B(B[13]), .Z(n1998) );
  AND U1749 ( .A(n1999), .B(n2000), .Z(n1997) );
  NANDN U1750 ( .A(A[12]), .B(B[12]), .Z(n2000) );
  NAND U1751 ( .A(n2001), .B(n2002), .Z(n1999) );
  NANDN U1752 ( .A(B[12]), .B(A[12]), .Z(n2002) );
  AND U1753 ( .A(n2003), .B(n2004), .Z(n2001) );
  NAND U1754 ( .A(n2005), .B(n2006), .Z(n2004) );
  NANDN U1755 ( .A(A[11]), .B(B[11]), .Z(n2006) );
  AND U1756 ( .A(n2007), .B(n2008), .Z(n2005) );
  NANDN U1757 ( .A(A[10]), .B(B[10]), .Z(n2008) );
  NAND U1758 ( .A(n2009), .B(n2010), .Z(n2007) );
  NANDN U1759 ( .A(B[9]), .B(A[9]), .Z(n2010) );
  AND U1760 ( .A(n2011), .B(n2012), .Z(n2009) );
  NAND U1761 ( .A(n2013), .B(n2014), .Z(n2012) );
  NANDN U1762 ( .A(A[9]), .B(B[9]), .Z(n2014) );
  AND U1763 ( .A(n2015), .B(n2016), .Z(n2013) );
  NANDN U1764 ( .A(A[8]), .B(B[8]), .Z(n2016) );
  NAND U1765 ( .A(n2017), .B(n2018), .Z(n2015) );
  NANDN U1766 ( .A(B[8]), .B(A[8]), .Z(n2018) );
  AND U1767 ( .A(n2019), .B(n2020), .Z(n2017) );
  NAND U1768 ( .A(n2021), .B(n2022), .Z(n2020) );
  NANDN U1769 ( .A(A[7]), .B(B[7]), .Z(n2022) );
  AND U1770 ( .A(n2023), .B(n2024), .Z(n2021) );
  NANDN U1771 ( .A(A[6]), .B(B[6]), .Z(n2024) );
  NAND U1772 ( .A(n2025), .B(n2026), .Z(n2023) );
  NANDN U1773 ( .A(B[6]), .B(A[6]), .Z(n2026) );
  AND U1774 ( .A(n2027), .B(n2028), .Z(n2025) );
  NAND U1775 ( .A(n2029), .B(n2030), .Z(n2028) );
  NANDN U1776 ( .A(A[5]), .B(B[5]), .Z(n2030) );
  AND U1777 ( .A(n2031), .B(n2032), .Z(n2029) );
  NANDN U1778 ( .A(A[4]), .B(B[4]), .Z(n2032) );
  NAND U1779 ( .A(n2033), .B(n2034), .Z(n2031) );
  NANDN U1780 ( .A(B[4]), .B(A[4]), .Z(n2034) );
  AND U1781 ( .A(n2035), .B(n2036), .Z(n2033) );
  NAND U1782 ( .A(n2037), .B(n2038), .Z(n2036) );
  NANDN U1783 ( .A(A[3]), .B(B[3]), .Z(n2038) );
  AND U1784 ( .A(n2039), .B(n2040), .Z(n2037) );
  NANDN U1785 ( .A(A[2]), .B(B[2]), .Z(n2040) );
  NAND U1786 ( .A(n2041), .B(n2042), .Z(n2039) );
  NANDN U1787 ( .A(B[2]), .B(A[2]), .Z(n2042) );
  AND U1788 ( .A(n2043), .B(n2044), .Z(n2041) );
  NAND U1789 ( .A(n2045), .B(A[0]), .Z(n2044) );
  ANDN U1790 ( .B(n2046), .A(B[0]), .Z(n2045) );
  NANDN U1791 ( .A(A[1]), .B(B[1]), .Z(n2046) );
  NANDN U1792 ( .A(B[1]), .B(A[1]), .Z(n2043) );
  NANDN U1793 ( .A(B[3]), .B(A[3]), .Z(n2035) );
  NANDN U1794 ( .A(B[5]), .B(A[5]), .Z(n2027) );
  NANDN U1795 ( .A(B[7]), .B(A[7]), .Z(n2019) );
  NANDN U1796 ( .A(B[10]), .B(A[10]), .Z(n2011) );
  NANDN U1797 ( .A(B[11]), .B(A[11]), .Z(n2003) );
  NANDN U1798 ( .A(B[13]), .B(A[13]), .Z(n1995) );
  NANDN U1799 ( .A(B[15]), .B(A[15]), .Z(n1987) );
  NANDN U1800 ( .A(B[17]), .B(A[17]), .Z(n1979) );
  NANDN U1801 ( .A(B[19]), .B(A[19]), .Z(n1971) );
  NANDN U1802 ( .A(B[21]), .B(A[21]), .Z(n1963) );
  NANDN U1803 ( .A(B[23]), .B(A[23]), .Z(n1955) );
  NANDN U1804 ( .A(B[25]), .B(A[25]), .Z(n1947) );
  NANDN U1805 ( .A(B[27]), .B(A[27]), .Z(n1939) );
  NANDN U1806 ( .A(B[29]), .B(A[29]), .Z(n1931) );
  NANDN U1807 ( .A(B[31]), .B(A[31]), .Z(n1923) );
  NANDN U1808 ( .A(B[33]), .B(A[33]), .Z(n1915) );
  NANDN U1809 ( .A(B[35]), .B(A[35]), .Z(n1907) );
  NANDN U1810 ( .A(B[37]), .B(A[37]), .Z(n1899) );
  NANDN U1811 ( .A(B[39]), .B(A[39]), .Z(n1891) );
  NANDN U1812 ( .A(B[41]), .B(A[41]), .Z(n1883) );
  NANDN U1813 ( .A(B[43]), .B(A[43]), .Z(n1875) );
  NANDN U1814 ( .A(B[45]), .B(A[45]), .Z(n1867) );
  NANDN U1815 ( .A(B[47]), .B(A[47]), .Z(n1859) );
  NANDN U1816 ( .A(B[49]), .B(A[49]), .Z(n1851) );
  NANDN U1817 ( .A(B[51]), .B(A[51]), .Z(n1843) );
  NANDN U1818 ( .A(B[53]), .B(A[53]), .Z(n1835) );
  NANDN U1819 ( .A(B[55]), .B(A[55]), .Z(n1827) );
  NANDN U1820 ( .A(B[57]), .B(A[57]), .Z(n1819) );
  NANDN U1821 ( .A(B[59]), .B(A[59]), .Z(n1811) );
  NANDN U1822 ( .A(B[61]), .B(A[61]), .Z(n1803) );
  NANDN U1823 ( .A(B[63]), .B(A[63]), .Z(n1795) );
  NANDN U1824 ( .A(B[65]), .B(A[65]), .Z(n1787) );
  NANDN U1825 ( .A(B[67]), .B(A[67]), .Z(n1779) );
  NANDN U1826 ( .A(B[69]), .B(A[69]), .Z(n1771) );
  NANDN U1827 ( .A(B[71]), .B(A[71]), .Z(n1763) );
  NANDN U1828 ( .A(B[73]), .B(A[73]), .Z(n1755) );
  NANDN U1829 ( .A(B[75]), .B(A[75]), .Z(n1747) );
  NANDN U1830 ( .A(B[77]), .B(A[77]), .Z(n1739) );
  NANDN U1831 ( .A(B[79]), .B(A[79]), .Z(n1731) );
  NANDN U1832 ( .A(B[81]), .B(A[81]), .Z(n1723) );
  NANDN U1833 ( .A(B[83]), .B(A[83]), .Z(n1715) );
  NANDN U1834 ( .A(B[85]), .B(A[85]), .Z(n1707) );
  NANDN U1835 ( .A(B[87]), .B(A[87]), .Z(n1699) );
  NANDN U1836 ( .A(B[89]), .B(A[89]), .Z(n1691) );
  NANDN U1837 ( .A(B[91]), .B(A[91]), .Z(n1683) );
  NANDN U1838 ( .A(B[93]), .B(A[93]), .Z(n1675) );
  NANDN U1839 ( .A(B[95]), .B(A[95]), .Z(n1667) );
  NANDN U1840 ( .A(B[97]), .B(A[97]), .Z(n1659) );
  NANDN U1841 ( .A(B[100]), .B(A[100]), .Z(n1651) );
  NANDN U1842 ( .A(B[101]), .B(A[101]), .Z(n1643) );
  NANDN U1843 ( .A(B[103]), .B(A[103]), .Z(n1635) );
  NANDN U1844 ( .A(B[105]), .B(A[105]), .Z(n1627) );
  NANDN U1845 ( .A(B[107]), .B(A[107]), .Z(n1619) );
  NANDN U1846 ( .A(B[109]), .B(A[109]), .Z(n1611) );
  NANDN U1847 ( .A(B[111]), .B(A[111]), .Z(n1603) );
  NANDN U1848 ( .A(B[113]), .B(A[113]), .Z(n1595) );
  NANDN U1849 ( .A(B[115]), .B(A[115]), .Z(n1587) );
  NANDN U1850 ( .A(B[117]), .B(A[117]), .Z(n1579) );
  NANDN U1851 ( .A(B[119]), .B(A[119]), .Z(n1571) );
  NANDN U1852 ( .A(B[121]), .B(A[121]), .Z(n1563) );
  NANDN U1853 ( .A(B[123]), .B(A[123]), .Z(n1555) );
  NANDN U1854 ( .A(B[125]), .B(A[125]), .Z(n1547) );
  NANDN U1855 ( .A(B[127]), .B(A[127]), .Z(n1539) );
  NANDN U1856 ( .A(B[129]), .B(A[129]), .Z(n1531) );
  NANDN U1857 ( .A(B[131]), .B(A[131]), .Z(n1523) );
  NANDN U1858 ( .A(B[133]), .B(A[133]), .Z(n1515) );
  NANDN U1859 ( .A(B[135]), .B(A[135]), .Z(n1507) );
  NANDN U1860 ( .A(B[137]), .B(A[137]), .Z(n1499) );
  NANDN U1861 ( .A(B[139]), .B(A[139]), .Z(n1491) );
  NANDN U1862 ( .A(B[141]), .B(A[141]), .Z(n1483) );
  NANDN U1863 ( .A(B[143]), .B(A[143]), .Z(n1475) );
  NANDN U1864 ( .A(B[145]), .B(A[145]), .Z(n1467) );
  NANDN U1865 ( .A(B[147]), .B(A[147]), .Z(n1459) );
  NANDN U1866 ( .A(B[149]), .B(A[149]), .Z(n1451) );
  NANDN U1867 ( .A(B[151]), .B(A[151]), .Z(n1443) );
  NANDN U1868 ( .A(B[153]), .B(A[153]), .Z(n1435) );
  NANDN U1869 ( .A(B[155]), .B(A[155]), .Z(n1427) );
  NANDN U1870 ( .A(B[157]), .B(A[157]), .Z(n1419) );
  NANDN U1871 ( .A(B[159]), .B(A[159]), .Z(n1411) );
  NANDN U1872 ( .A(B[161]), .B(A[161]), .Z(n1403) );
  NANDN U1873 ( .A(B[163]), .B(A[163]), .Z(n1395) );
  NANDN U1874 ( .A(B[165]), .B(A[165]), .Z(n1387) );
  NANDN U1875 ( .A(B[167]), .B(A[167]), .Z(n1379) );
  NANDN U1876 ( .A(B[169]), .B(A[169]), .Z(n1371) );
  NANDN U1877 ( .A(B[171]), .B(A[171]), .Z(n1363) );
  NANDN U1878 ( .A(B[173]), .B(A[173]), .Z(n1355) );
  NANDN U1879 ( .A(B[175]), .B(A[175]), .Z(n1347) );
  NANDN U1880 ( .A(B[177]), .B(A[177]), .Z(n1339) );
  NANDN U1881 ( .A(B[179]), .B(A[179]), .Z(n1331) );
  NANDN U1882 ( .A(B[181]), .B(A[181]), .Z(n1323) );
  NANDN U1883 ( .A(B[183]), .B(A[183]), .Z(n1315) );
  NANDN U1884 ( .A(B[185]), .B(A[185]), .Z(n1307) );
  NANDN U1885 ( .A(B[187]), .B(A[187]), .Z(n1299) );
  NANDN U1886 ( .A(B[189]), .B(A[189]), .Z(n1291) );
  NANDN U1887 ( .A(B[191]), .B(A[191]), .Z(n1283) );
  NANDN U1888 ( .A(B[193]), .B(A[193]), .Z(n1275) );
  NANDN U1889 ( .A(B[195]), .B(A[195]), .Z(n1267) );
  NANDN U1890 ( .A(B[197]), .B(A[197]), .Z(n1259) );
  NANDN U1891 ( .A(B[199]), .B(A[199]), .Z(n1251) );
  NANDN U1892 ( .A(B[201]), .B(A[201]), .Z(n1243) );
  NANDN U1893 ( .A(B[203]), .B(A[203]), .Z(n1235) );
  NANDN U1894 ( .A(B[205]), .B(A[205]), .Z(n1227) );
  NANDN U1895 ( .A(B[207]), .B(A[207]), .Z(n1219) );
  NANDN U1896 ( .A(B[209]), .B(A[209]), .Z(n1211) );
  NANDN U1897 ( .A(B[211]), .B(A[211]), .Z(n1203) );
  NANDN U1898 ( .A(B[213]), .B(A[213]), .Z(n1195) );
  NANDN U1899 ( .A(B[215]), .B(A[215]), .Z(n1187) );
  NANDN U1900 ( .A(B[217]), .B(A[217]), .Z(n1179) );
  NANDN U1901 ( .A(B[219]), .B(A[219]), .Z(n1171) );
  NANDN U1902 ( .A(B[221]), .B(A[221]), .Z(n1163) );
  NANDN U1903 ( .A(B[223]), .B(A[223]), .Z(n1155) );
  NANDN U1904 ( .A(B[225]), .B(A[225]), .Z(n1147) );
  NANDN U1905 ( .A(B[227]), .B(A[227]), .Z(n1139) );
  NANDN U1906 ( .A(B[229]), .B(A[229]), .Z(n1131) );
  NANDN U1907 ( .A(B[231]), .B(A[231]), .Z(n1123) );
  NANDN U1908 ( .A(B[233]), .B(A[233]), .Z(n1115) );
  NANDN U1909 ( .A(B[235]), .B(A[235]), .Z(n1107) );
  NANDN U1910 ( .A(B[237]), .B(A[237]), .Z(n1099) );
  NANDN U1911 ( .A(B[239]), .B(A[239]), .Z(n1091) );
  NANDN U1912 ( .A(B[241]), .B(A[241]), .Z(n1083) );
  NANDN U1913 ( .A(B[243]), .B(A[243]), .Z(n1075) );
  NANDN U1914 ( .A(B[245]), .B(A[245]), .Z(n1067) );
  NANDN U1915 ( .A(B[247]), .B(A[247]), .Z(n1059) );
  NANDN U1916 ( .A(B[249]), .B(A[249]), .Z(n1051) );
  NANDN U1917 ( .A(B[251]), .B(A[251]), .Z(n1043) );
  NANDN U1918 ( .A(B[253]), .B(A[253]), .Z(n1035) );
  NANDN U1919 ( .A(B[255]), .B(A[255]), .Z(n1027) );
  NANDN U1920 ( .A(B[257]), .B(A[257]), .Z(n1019) );
  NANDN U1921 ( .A(B[259]), .B(A[259]), .Z(n1011) );
  NANDN U1922 ( .A(B[261]), .B(A[261]), .Z(n1003) );
  NANDN U1923 ( .A(B[263]), .B(A[263]), .Z(n995) );
  NANDN U1924 ( .A(B[265]), .B(A[265]), .Z(n987) );
  NANDN U1925 ( .A(B[267]), .B(A[267]), .Z(n979) );
  NANDN U1926 ( .A(B[269]), .B(A[269]), .Z(n971) );
  NANDN U1927 ( .A(B[271]), .B(A[271]), .Z(n963) );
  NANDN U1928 ( .A(B[273]), .B(A[273]), .Z(n955) );
  NANDN U1929 ( .A(B[275]), .B(A[275]), .Z(n947) );
  NANDN U1930 ( .A(B[277]), .B(A[277]), .Z(n939) );
  NANDN U1931 ( .A(B[279]), .B(A[279]), .Z(n931) );
  NANDN U1932 ( .A(B[281]), .B(A[281]), .Z(n923) );
  NANDN U1933 ( .A(B[283]), .B(A[283]), .Z(n915) );
  NANDN U1934 ( .A(B[285]), .B(A[285]), .Z(n907) );
  NANDN U1935 ( .A(B[287]), .B(A[287]), .Z(n899) );
  NANDN U1936 ( .A(B[289]), .B(A[289]), .Z(n891) );
  NANDN U1937 ( .A(B[291]), .B(A[291]), .Z(n883) );
  NANDN U1938 ( .A(B[293]), .B(A[293]), .Z(n875) );
  NANDN U1939 ( .A(B[295]), .B(A[295]), .Z(n867) );
  NANDN U1940 ( .A(B[297]), .B(A[297]), .Z(n859) );
  NANDN U1941 ( .A(B[299]), .B(A[299]), .Z(n851) );
  NANDN U1942 ( .A(B[301]), .B(A[301]), .Z(n843) );
  NANDN U1943 ( .A(B[303]), .B(A[303]), .Z(n835) );
  NANDN U1944 ( .A(B[305]), .B(A[305]), .Z(n827) );
  NANDN U1945 ( .A(B[307]), .B(A[307]), .Z(n819) );
  NANDN U1946 ( .A(B[309]), .B(A[309]), .Z(n811) );
  NANDN U1947 ( .A(B[311]), .B(A[311]), .Z(n803) );
  NANDN U1948 ( .A(B[313]), .B(A[313]), .Z(n795) );
  NANDN U1949 ( .A(B[315]), .B(A[315]), .Z(n787) );
  NANDN U1950 ( .A(B[317]), .B(A[317]), .Z(n779) );
  NANDN U1951 ( .A(B[319]), .B(A[319]), .Z(n771) );
  NANDN U1952 ( .A(B[321]), .B(A[321]), .Z(n763) );
  NANDN U1953 ( .A(B[323]), .B(A[323]), .Z(n755) );
  NANDN U1954 ( .A(B[325]), .B(A[325]), .Z(n747) );
  NANDN U1955 ( .A(B[327]), .B(A[327]), .Z(n739) );
  NANDN U1956 ( .A(B[329]), .B(A[329]), .Z(n731) );
  NANDN U1957 ( .A(B[331]), .B(A[331]), .Z(n723) );
  NANDN U1958 ( .A(B[333]), .B(A[333]), .Z(n715) );
  NANDN U1959 ( .A(B[335]), .B(A[335]), .Z(n707) );
  NANDN U1960 ( .A(B[337]), .B(A[337]), .Z(n699) );
  NANDN U1961 ( .A(B[339]), .B(A[339]), .Z(n691) );
  NANDN U1962 ( .A(B[341]), .B(A[341]), .Z(n683) );
  NANDN U1963 ( .A(B[343]), .B(A[343]), .Z(n675) );
  NANDN U1964 ( .A(B[345]), .B(A[345]), .Z(n667) );
  NANDN U1965 ( .A(B[347]), .B(A[347]), .Z(n659) );
  NANDN U1966 ( .A(B[349]), .B(A[349]), .Z(n651) );
  NANDN U1967 ( .A(B[351]), .B(A[351]), .Z(n643) );
  NANDN U1968 ( .A(B[353]), .B(A[353]), .Z(n635) );
  NANDN U1969 ( .A(B[355]), .B(A[355]), .Z(n627) );
  NANDN U1970 ( .A(B[357]), .B(A[357]), .Z(n619) );
  NANDN U1971 ( .A(B[359]), .B(A[359]), .Z(n611) );
  NANDN U1972 ( .A(B[361]), .B(A[361]), .Z(n603) );
  NANDN U1973 ( .A(B[363]), .B(A[363]), .Z(n595) );
  NANDN U1974 ( .A(B[365]), .B(A[365]), .Z(n587) );
  NANDN U1975 ( .A(B[367]), .B(A[367]), .Z(n579) );
  NANDN U1976 ( .A(B[369]), .B(A[369]), .Z(n571) );
  NANDN U1977 ( .A(B[371]), .B(A[371]), .Z(n563) );
  NANDN U1978 ( .A(B[373]), .B(A[373]), .Z(n555) );
  NANDN U1979 ( .A(B[375]), .B(A[375]), .Z(n547) );
  NANDN U1980 ( .A(B[377]), .B(A[377]), .Z(n539) );
  NANDN U1981 ( .A(B[379]), .B(A[379]), .Z(n531) );
  NANDN U1982 ( .A(B[381]), .B(A[381]), .Z(n523) );
  NANDN U1983 ( .A(B[383]), .B(A[383]), .Z(n515) );
  NANDN U1984 ( .A(B[385]), .B(A[385]), .Z(n507) );
  NANDN U1985 ( .A(B[387]), .B(A[387]), .Z(n499) );
  NANDN U1986 ( .A(B[389]), .B(A[389]), .Z(n491) );
  NANDN U1987 ( .A(B[391]), .B(A[391]), .Z(n483) );
  NANDN U1988 ( .A(B[393]), .B(A[393]), .Z(n475) );
  NANDN U1989 ( .A(B[395]), .B(A[395]), .Z(n467) );
  NANDN U1990 ( .A(B[397]), .B(A[397]), .Z(n459) );
  NANDN U1991 ( .A(B[399]), .B(A[399]), .Z(n451) );
  NANDN U1992 ( .A(B[401]), .B(A[401]), .Z(n443) );
  NANDN U1993 ( .A(B[403]), .B(A[403]), .Z(n435) );
  NANDN U1994 ( .A(B[405]), .B(A[405]), .Z(n427) );
  NANDN U1995 ( .A(B[407]), .B(A[407]), .Z(n419) );
  NANDN U1996 ( .A(B[409]), .B(A[409]), .Z(n411) );
  NANDN U1997 ( .A(B[411]), .B(A[411]), .Z(n403) );
  NANDN U1998 ( .A(B[413]), .B(A[413]), .Z(n395) );
  NANDN U1999 ( .A(B[415]), .B(A[415]), .Z(n387) );
  NANDN U2000 ( .A(B[417]), .B(A[417]), .Z(n379) );
  NANDN U2001 ( .A(B[419]), .B(A[419]), .Z(n371) );
  NANDN U2002 ( .A(B[421]), .B(A[421]), .Z(n363) );
  NANDN U2003 ( .A(B[423]), .B(A[423]), .Z(n355) );
  NANDN U2004 ( .A(B[425]), .B(A[425]), .Z(n347) );
  NANDN U2005 ( .A(B[427]), .B(A[427]), .Z(n339) );
  NANDN U2006 ( .A(B[429]), .B(A[429]), .Z(n331) );
  NANDN U2007 ( .A(B[431]), .B(A[431]), .Z(n323) );
  NANDN U2008 ( .A(B[433]), .B(A[433]), .Z(n315) );
  NANDN U2009 ( .A(B[435]), .B(A[435]), .Z(n307) );
  NANDN U2010 ( .A(B[437]), .B(A[437]), .Z(n299) );
  NANDN U2011 ( .A(B[439]), .B(A[439]), .Z(n291) );
  NANDN U2012 ( .A(B[441]), .B(A[441]), .Z(n283) );
  NANDN U2013 ( .A(B[443]), .B(A[443]), .Z(n275) );
  NANDN U2014 ( .A(B[445]), .B(A[445]), .Z(n267) );
  NANDN U2015 ( .A(B[447]), .B(A[447]), .Z(n259) );
  NANDN U2016 ( .A(B[449]), .B(A[449]), .Z(n251) );
  NANDN U2017 ( .A(B[451]), .B(A[451]), .Z(n243) );
  NANDN U2018 ( .A(B[453]), .B(A[453]), .Z(n235) );
  NANDN U2019 ( .A(B[455]), .B(A[455]), .Z(n227) );
  NANDN U2020 ( .A(B[457]), .B(A[457]), .Z(n219) );
  NANDN U2021 ( .A(B[459]), .B(A[459]), .Z(n211) );
  NANDN U2022 ( .A(B[461]), .B(A[461]), .Z(n203) );
  NANDN U2023 ( .A(B[463]), .B(A[463]), .Z(n195) );
  NANDN U2024 ( .A(B[465]), .B(A[465]), .Z(n187) );
  NANDN U2025 ( .A(B[467]), .B(A[467]), .Z(n179) );
  NANDN U2026 ( .A(B[469]), .B(A[469]), .Z(n171) );
  NANDN U2027 ( .A(B[471]), .B(A[471]), .Z(n163) );
  NANDN U2028 ( .A(B[473]), .B(A[473]), .Z(n155) );
  NANDN U2029 ( .A(B[475]), .B(A[475]), .Z(n147) );
  NANDN U2030 ( .A(B[477]), .B(A[477]), .Z(n139) );
  NANDN U2031 ( .A(B[479]), .B(A[479]), .Z(n131) );
  NANDN U2032 ( .A(B[481]), .B(A[481]), .Z(n123) );
  NANDN U2033 ( .A(B[483]), .B(A[483]), .Z(n115) );
  NANDN U2034 ( .A(B[485]), .B(A[485]), .Z(n107) );
  NANDN U2035 ( .A(B[487]), .B(A[487]), .Z(n99) );
  NANDN U2036 ( .A(B[489]), .B(A[489]), .Z(n91) );
  NANDN U2037 ( .A(B[491]), .B(A[491]), .Z(n83) );
  NANDN U2038 ( .A(B[493]), .B(A[493]), .Z(n75) );
  NANDN U2039 ( .A(B[495]), .B(A[495]), .Z(n67) );
  NANDN U2040 ( .A(B[497]), .B(A[497]), .Z(n59) );
  NANDN U2041 ( .A(B[499]), .B(A[499]), .Z(n51) );
  NANDN U2042 ( .A(B[501]), .B(A[501]), .Z(n43) );
  NANDN U2043 ( .A(B[503]), .B(A[503]), .Z(n35) );
  NANDN U2044 ( .A(B[505]), .B(A[505]), .Z(n27) );
  NANDN U2045 ( .A(B[507]), .B(A[507]), .Z(n19) );
  NANDN U2046 ( .A(B[509]), .B(A[509]), .Z(n11) );
  NANDN U2047 ( .A(A[511]), .B(B[511]), .Z(n3) );
endmodule


module modmult_step_N512_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [513:0] A;
  input [513:0] B;
  output [513:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560;

  IV U1 ( .A(A[1]), .Z(n1) );
  IV U2 ( .A(n2559), .Z(n2) );
  XNOR U3 ( .A(n3), .B(n4), .Z(DIFF[9]) );
  XOR U4 ( .A(B[9]), .B(A[9]), .Z(n4) );
  XNOR U5 ( .A(n5), .B(n6), .Z(DIFF[99]) );
  XOR U6 ( .A(B[99]), .B(A[99]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(DIFF[98]) );
  XOR U8 ( .A(B[98]), .B(A[98]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(DIFF[97]) );
  XOR U10 ( .A(B[97]), .B(A[97]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(DIFF[96]) );
  XOR U12 ( .A(B[96]), .B(A[96]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(DIFF[95]) );
  XOR U14 ( .A(B[95]), .B(A[95]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(DIFF[94]) );
  XOR U16 ( .A(B[94]), .B(A[94]), .Z(n16) );
  XOR U17 ( .A(n17), .B(n18), .Z(DIFF[93]) );
  XOR U18 ( .A(B[93]), .B(A[93]), .Z(n18) );
  XOR U19 ( .A(n19), .B(n20), .Z(DIFF[92]) );
  XOR U20 ( .A(B[92]), .B(A[92]), .Z(n20) );
  XOR U21 ( .A(n21), .B(n22), .Z(DIFF[91]) );
  XOR U22 ( .A(B[91]), .B(A[91]), .Z(n22) );
  XOR U23 ( .A(n23), .B(n24), .Z(DIFF[90]) );
  XOR U24 ( .A(B[90]), .B(A[90]), .Z(n24) );
  XOR U25 ( .A(n25), .B(n26), .Z(DIFF[8]) );
  XOR U26 ( .A(B[8]), .B(A[8]), .Z(n26) );
  XOR U27 ( .A(n27), .B(n28), .Z(DIFF[89]) );
  XOR U28 ( .A(B[89]), .B(A[89]), .Z(n28) );
  XOR U29 ( .A(n29), .B(n30), .Z(DIFF[88]) );
  XOR U30 ( .A(B[88]), .B(A[88]), .Z(n30) );
  XOR U31 ( .A(n31), .B(n32), .Z(DIFF[87]) );
  XOR U32 ( .A(B[87]), .B(A[87]), .Z(n32) );
  XOR U33 ( .A(n33), .B(n34), .Z(DIFF[86]) );
  XOR U34 ( .A(B[86]), .B(A[86]), .Z(n34) );
  XOR U35 ( .A(n35), .B(n36), .Z(DIFF[85]) );
  XOR U36 ( .A(B[85]), .B(A[85]), .Z(n36) );
  XOR U37 ( .A(n37), .B(n38), .Z(DIFF[84]) );
  XOR U38 ( .A(B[84]), .B(A[84]), .Z(n38) );
  XOR U39 ( .A(n39), .B(n40), .Z(DIFF[83]) );
  XOR U40 ( .A(B[83]), .B(A[83]), .Z(n40) );
  XOR U41 ( .A(n41), .B(n42), .Z(DIFF[82]) );
  XOR U42 ( .A(B[82]), .B(A[82]), .Z(n42) );
  XOR U43 ( .A(n43), .B(n44), .Z(DIFF[81]) );
  XOR U44 ( .A(B[81]), .B(A[81]), .Z(n44) );
  XOR U45 ( .A(n45), .B(n46), .Z(DIFF[80]) );
  XOR U46 ( .A(B[80]), .B(A[80]), .Z(n46) );
  XOR U47 ( .A(n47), .B(n48), .Z(DIFF[7]) );
  XOR U48 ( .A(B[7]), .B(A[7]), .Z(n48) );
  XOR U49 ( .A(n49), .B(n50), .Z(DIFF[79]) );
  XOR U50 ( .A(B[79]), .B(A[79]), .Z(n50) );
  XOR U51 ( .A(n51), .B(n52), .Z(DIFF[78]) );
  XOR U52 ( .A(B[78]), .B(A[78]), .Z(n52) );
  XOR U53 ( .A(n53), .B(n54), .Z(DIFF[77]) );
  XOR U54 ( .A(B[77]), .B(A[77]), .Z(n54) );
  XOR U55 ( .A(n55), .B(n56), .Z(DIFF[76]) );
  XOR U56 ( .A(B[76]), .B(A[76]), .Z(n56) );
  XOR U57 ( .A(n57), .B(n58), .Z(DIFF[75]) );
  XOR U58 ( .A(B[75]), .B(A[75]), .Z(n58) );
  XOR U59 ( .A(n59), .B(n60), .Z(DIFF[74]) );
  XOR U60 ( .A(B[74]), .B(A[74]), .Z(n60) );
  XOR U61 ( .A(n61), .B(n62), .Z(DIFF[73]) );
  XOR U62 ( .A(B[73]), .B(A[73]), .Z(n62) );
  XOR U63 ( .A(n63), .B(n64), .Z(DIFF[72]) );
  XOR U64 ( .A(B[72]), .B(A[72]), .Z(n64) );
  XOR U65 ( .A(n65), .B(n66), .Z(DIFF[71]) );
  XOR U66 ( .A(B[71]), .B(A[71]), .Z(n66) );
  XOR U67 ( .A(n67), .B(n68), .Z(DIFF[70]) );
  XOR U68 ( .A(B[70]), .B(A[70]), .Z(n68) );
  XOR U69 ( .A(n69), .B(n70), .Z(DIFF[6]) );
  XOR U70 ( .A(B[6]), .B(A[6]), .Z(n70) );
  XOR U71 ( .A(n71), .B(n72), .Z(DIFF[69]) );
  XOR U72 ( .A(B[69]), .B(A[69]), .Z(n72) );
  XOR U73 ( .A(n73), .B(n74), .Z(DIFF[68]) );
  XOR U74 ( .A(B[68]), .B(A[68]), .Z(n74) );
  XOR U75 ( .A(n75), .B(n76), .Z(DIFF[67]) );
  XOR U76 ( .A(B[67]), .B(A[67]), .Z(n76) );
  XOR U77 ( .A(n77), .B(n78), .Z(DIFF[66]) );
  XOR U78 ( .A(B[66]), .B(A[66]), .Z(n78) );
  XOR U79 ( .A(n79), .B(n80), .Z(DIFF[65]) );
  XOR U80 ( .A(B[65]), .B(A[65]), .Z(n80) );
  XOR U81 ( .A(n81), .B(n82), .Z(DIFF[64]) );
  XOR U82 ( .A(B[64]), .B(A[64]), .Z(n82) );
  XOR U83 ( .A(n83), .B(n84), .Z(DIFF[63]) );
  XOR U84 ( .A(B[63]), .B(A[63]), .Z(n84) );
  XOR U85 ( .A(n85), .B(n86), .Z(DIFF[62]) );
  XOR U86 ( .A(B[62]), .B(A[62]), .Z(n86) );
  XOR U87 ( .A(n87), .B(n88), .Z(DIFF[61]) );
  XOR U88 ( .A(B[61]), .B(A[61]), .Z(n88) );
  XOR U89 ( .A(n89), .B(n90), .Z(DIFF[60]) );
  XOR U90 ( .A(B[60]), .B(A[60]), .Z(n90) );
  XOR U91 ( .A(n91), .B(n92), .Z(DIFF[5]) );
  XOR U92 ( .A(B[5]), .B(A[5]), .Z(n92) );
  XOR U93 ( .A(n93), .B(n94), .Z(DIFF[59]) );
  XOR U94 ( .A(B[59]), .B(A[59]), .Z(n94) );
  XOR U95 ( .A(n95), .B(n96), .Z(DIFF[58]) );
  XOR U96 ( .A(B[58]), .B(A[58]), .Z(n96) );
  XOR U97 ( .A(n97), .B(n98), .Z(DIFF[57]) );
  XOR U98 ( .A(B[57]), .B(A[57]), .Z(n98) );
  XOR U99 ( .A(n99), .B(n100), .Z(DIFF[56]) );
  XOR U100 ( .A(B[56]), .B(A[56]), .Z(n100) );
  XOR U101 ( .A(n101), .B(n102), .Z(DIFF[55]) );
  XOR U102 ( .A(B[55]), .B(A[55]), .Z(n102) );
  XOR U103 ( .A(n103), .B(n104), .Z(DIFF[54]) );
  XOR U104 ( .A(B[54]), .B(A[54]), .Z(n104) );
  XOR U105 ( .A(n105), .B(n106), .Z(DIFF[53]) );
  XOR U106 ( .A(B[53]), .B(A[53]), .Z(n106) );
  XOR U107 ( .A(n107), .B(n108), .Z(DIFF[52]) );
  XOR U108 ( .A(B[52]), .B(A[52]), .Z(n108) );
  XOR U109 ( .A(n109), .B(n110), .Z(DIFF[51]) );
  XOR U110 ( .A(B[51]), .B(A[51]), .Z(n110) );
  XOR U111 ( .A(A[513]), .B(n111), .Z(DIFF[513]) );
  ANDN U112 ( .B(n112), .A(A[512]), .Z(n111) );
  XOR U113 ( .A(A[512]), .B(n112), .Z(DIFF[512]) );
  AND U114 ( .A(n113), .B(n114), .Z(n112) );
  NANDN U115 ( .A(B[511]), .B(n115), .Z(n114) );
  NANDN U116 ( .A(A[511]), .B(n116), .Z(n115) );
  NANDN U117 ( .A(n116), .B(A[511]), .Z(n113) );
  XOR U118 ( .A(n116), .B(n117), .Z(DIFF[511]) );
  XOR U119 ( .A(B[511]), .B(A[511]), .Z(n117) );
  AND U120 ( .A(n118), .B(n119), .Z(n116) );
  NANDN U121 ( .A(B[510]), .B(n120), .Z(n119) );
  NANDN U122 ( .A(A[510]), .B(n121), .Z(n120) );
  NANDN U123 ( .A(n121), .B(A[510]), .Z(n118) );
  XOR U124 ( .A(n121), .B(n122), .Z(DIFF[510]) );
  XOR U125 ( .A(B[510]), .B(A[510]), .Z(n122) );
  AND U126 ( .A(n123), .B(n124), .Z(n121) );
  NANDN U127 ( .A(B[509]), .B(n125), .Z(n124) );
  NANDN U128 ( .A(A[509]), .B(n126), .Z(n125) );
  NANDN U129 ( .A(n126), .B(A[509]), .Z(n123) );
  XOR U130 ( .A(n127), .B(n128), .Z(DIFF[50]) );
  XOR U131 ( .A(B[50]), .B(A[50]), .Z(n128) );
  XOR U132 ( .A(n126), .B(n129), .Z(DIFF[509]) );
  XOR U133 ( .A(B[509]), .B(A[509]), .Z(n129) );
  AND U134 ( .A(n130), .B(n131), .Z(n126) );
  NANDN U135 ( .A(B[508]), .B(n132), .Z(n131) );
  NANDN U136 ( .A(A[508]), .B(n133), .Z(n132) );
  NANDN U137 ( .A(n133), .B(A[508]), .Z(n130) );
  XOR U138 ( .A(n133), .B(n134), .Z(DIFF[508]) );
  XOR U139 ( .A(B[508]), .B(A[508]), .Z(n134) );
  AND U140 ( .A(n135), .B(n136), .Z(n133) );
  NANDN U141 ( .A(B[507]), .B(n137), .Z(n136) );
  NANDN U142 ( .A(A[507]), .B(n138), .Z(n137) );
  NANDN U143 ( .A(n138), .B(A[507]), .Z(n135) );
  XOR U144 ( .A(n138), .B(n139), .Z(DIFF[507]) );
  XOR U145 ( .A(B[507]), .B(A[507]), .Z(n139) );
  AND U146 ( .A(n140), .B(n141), .Z(n138) );
  NANDN U147 ( .A(B[506]), .B(n142), .Z(n141) );
  NANDN U148 ( .A(A[506]), .B(n143), .Z(n142) );
  NANDN U149 ( .A(n143), .B(A[506]), .Z(n140) );
  XOR U150 ( .A(n143), .B(n144), .Z(DIFF[506]) );
  XOR U151 ( .A(B[506]), .B(A[506]), .Z(n144) );
  AND U152 ( .A(n145), .B(n146), .Z(n143) );
  NANDN U153 ( .A(B[505]), .B(n147), .Z(n146) );
  NANDN U154 ( .A(A[505]), .B(n148), .Z(n147) );
  NANDN U155 ( .A(n148), .B(A[505]), .Z(n145) );
  XOR U156 ( .A(n148), .B(n149), .Z(DIFF[505]) );
  XOR U157 ( .A(B[505]), .B(A[505]), .Z(n149) );
  AND U158 ( .A(n150), .B(n151), .Z(n148) );
  NANDN U159 ( .A(B[504]), .B(n152), .Z(n151) );
  NANDN U160 ( .A(A[504]), .B(n153), .Z(n152) );
  NANDN U161 ( .A(n153), .B(A[504]), .Z(n150) );
  XOR U162 ( .A(n153), .B(n154), .Z(DIFF[504]) );
  XOR U163 ( .A(B[504]), .B(A[504]), .Z(n154) );
  AND U164 ( .A(n155), .B(n156), .Z(n153) );
  NANDN U165 ( .A(B[503]), .B(n157), .Z(n156) );
  NANDN U166 ( .A(A[503]), .B(n158), .Z(n157) );
  NANDN U167 ( .A(n158), .B(A[503]), .Z(n155) );
  XOR U168 ( .A(n158), .B(n159), .Z(DIFF[503]) );
  XOR U169 ( .A(B[503]), .B(A[503]), .Z(n159) );
  AND U170 ( .A(n160), .B(n161), .Z(n158) );
  NANDN U171 ( .A(B[502]), .B(n162), .Z(n161) );
  NANDN U172 ( .A(A[502]), .B(n163), .Z(n162) );
  NANDN U173 ( .A(n163), .B(A[502]), .Z(n160) );
  XOR U174 ( .A(n163), .B(n164), .Z(DIFF[502]) );
  XOR U175 ( .A(B[502]), .B(A[502]), .Z(n164) );
  AND U176 ( .A(n165), .B(n166), .Z(n163) );
  NANDN U177 ( .A(B[501]), .B(n167), .Z(n166) );
  NANDN U178 ( .A(A[501]), .B(n168), .Z(n167) );
  NANDN U179 ( .A(n168), .B(A[501]), .Z(n165) );
  XOR U180 ( .A(n168), .B(n169), .Z(DIFF[501]) );
  XOR U181 ( .A(B[501]), .B(A[501]), .Z(n169) );
  AND U182 ( .A(n170), .B(n171), .Z(n168) );
  NANDN U183 ( .A(B[500]), .B(n172), .Z(n171) );
  NANDN U184 ( .A(A[500]), .B(n173), .Z(n172) );
  NANDN U185 ( .A(n173), .B(A[500]), .Z(n170) );
  XOR U186 ( .A(n173), .B(n174), .Z(DIFF[500]) );
  XOR U187 ( .A(B[500]), .B(A[500]), .Z(n174) );
  AND U188 ( .A(n175), .B(n176), .Z(n173) );
  NANDN U189 ( .A(B[499]), .B(n177), .Z(n176) );
  NANDN U190 ( .A(A[499]), .B(n178), .Z(n177) );
  NANDN U191 ( .A(n178), .B(A[499]), .Z(n175) );
  XOR U192 ( .A(n179), .B(n180), .Z(DIFF[4]) );
  XOR U193 ( .A(B[4]), .B(A[4]), .Z(n180) );
  XOR U194 ( .A(n181), .B(n182), .Z(DIFF[49]) );
  XOR U195 ( .A(B[49]), .B(A[49]), .Z(n182) );
  XOR U196 ( .A(n178), .B(n183), .Z(DIFF[499]) );
  XOR U197 ( .A(B[499]), .B(A[499]), .Z(n183) );
  AND U198 ( .A(n184), .B(n185), .Z(n178) );
  NANDN U199 ( .A(B[498]), .B(n186), .Z(n185) );
  NANDN U200 ( .A(A[498]), .B(n187), .Z(n186) );
  NANDN U201 ( .A(n187), .B(A[498]), .Z(n184) );
  XOR U202 ( .A(n187), .B(n188), .Z(DIFF[498]) );
  XOR U203 ( .A(B[498]), .B(A[498]), .Z(n188) );
  AND U204 ( .A(n189), .B(n190), .Z(n187) );
  NANDN U205 ( .A(B[497]), .B(n191), .Z(n190) );
  NANDN U206 ( .A(A[497]), .B(n192), .Z(n191) );
  NANDN U207 ( .A(n192), .B(A[497]), .Z(n189) );
  XOR U208 ( .A(n192), .B(n193), .Z(DIFF[497]) );
  XOR U209 ( .A(B[497]), .B(A[497]), .Z(n193) );
  AND U210 ( .A(n194), .B(n195), .Z(n192) );
  NANDN U211 ( .A(B[496]), .B(n196), .Z(n195) );
  NANDN U212 ( .A(A[496]), .B(n197), .Z(n196) );
  NANDN U213 ( .A(n197), .B(A[496]), .Z(n194) );
  XOR U214 ( .A(n197), .B(n198), .Z(DIFF[496]) );
  XOR U215 ( .A(B[496]), .B(A[496]), .Z(n198) );
  AND U216 ( .A(n199), .B(n200), .Z(n197) );
  NANDN U217 ( .A(B[495]), .B(n201), .Z(n200) );
  NANDN U218 ( .A(A[495]), .B(n202), .Z(n201) );
  NANDN U219 ( .A(n202), .B(A[495]), .Z(n199) );
  XOR U220 ( .A(n202), .B(n203), .Z(DIFF[495]) );
  XOR U221 ( .A(B[495]), .B(A[495]), .Z(n203) );
  AND U222 ( .A(n204), .B(n205), .Z(n202) );
  NANDN U223 ( .A(B[494]), .B(n206), .Z(n205) );
  NANDN U224 ( .A(A[494]), .B(n207), .Z(n206) );
  NANDN U225 ( .A(n207), .B(A[494]), .Z(n204) );
  XOR U226 ( .A(n207), .B(n208), .Z(DIFF[494]) );
  XOR U227 ( .A(B[494]), .B(A[494]), .Z(n208) );
  AND U228 ( .A(n209), .B(n210), .Z(n207) );
  NANDN U229 ( .A(B[493]), .B(n211), .Z(n210) );
  NANDN U230 ( .A(A[493]), .B(n212), .Z(n211) );
  NANDN U231 ( .A(n212), .B(A[493]), .Z(n209) );
  XOR U232 ( .A(n212), .B(n213), .Z(DIFF[493]) );
  XOR U233 ( .A(B[493]), .B(A[493]), .Z(n213) );
  AND U234 ( .A(n214), .B(n215), .Z(n212) );
  NANDN U235 ( .A(B[492]), .B(n216), .Z(n215) );
  NANDN U236 ( .A(A[492]), .B(n217), .Z(n216) );
  NANDN U237 ( .A(n217), .B(A[492]), .Z(n214) );
  XOR U238 ( .A(n217), .B(n218), .Z(DIFF[492]) );
  XOR U239 ( .A(B[492]), .B(A[492]), .Z(n218) );
  AND U240 ( .A(n219), .B(n220), .Z(n217) );
  NANDN U241 ( .A(B[491]), .B(n221), .Z(n220) );
  NANDN U242 ( .A(A[491]), .B(n222), .Z(n221) );
  NANDN U243 ( .A(n222), .B(A[491]), .Z(n219) );
  XOR U244 ( .A(n222), .B(n223), .Z(DIFF[491]) );
  XOR U245 ( .A(B[491]), .B(A[491]), .Z(n223) );
  AND U246 ( .A(n224), .B(n225), .Z(n222) );
  NANDN U247 ( .A(B[490]), .B(n226), .Z(n225) );
  NANDN U248 ( .A(A[490]), .B(n227), .Z(n226) );
  NANDN U249 ( .A(n227), .B(A[490]), .Z(n224) );
  XOR U250 ( .A(n227), .B(n228), .Z(DIFF[490]) );
  XOR U251 ( .A(B[490]), .B(A[490]), .Z(n228) );
  AND U252 ( .A(n229), .B(n230), .Z(n227) );
  NANDN U253 ( .A(B[489]), .B(n231), .Z(n230) );
  NANDN U254 ( .A(A[489]), .B(n232), .Z(n231) );
  NANDN U255 ( .A(n232), .B(A[489]), .Z(n229) );
  XOR U256 ( .A(n233), .B(n234), .Z(DIFF[48]) );
  XOR U257 ( .A(B[48]), .B(A[48]), .Z(n234) );
  XOR U258 ( .A(n232), .B(n235), .Z(DIFF[489]) );
  XOR U259 ( .A(B[489]), .B(A[489]), .Z(n235) );
  AND U260 ( .A(n236), .B(n237), .Z(n232) );
  NANDN U261 ( .A(B[488]), .B(n238), .Z(n237) );
  NANDN U262 ( .A(A[488]), .B(n239), .Z(n238) );
  NANDN U263 ( .A(n239), .B(A[488]), .Z(n236) );
  XOR U264 ( .A(n239), .B(n240), .Z(DIFF[488]) );
  XOR U265 ( .A(B[488]), .B(A[488]), .Z(n240) );
  AND U266 ( .A(n241), .B(n242), .Z(n239) );
  NANDN U267 ( .A(B[487]), .B(n243), .Z(n242) );
  NANDN U268 ( .A(A[487]), .B(n244), .Z(n243) );
  NANDN U269 ( .A(n244), .B(A[487]), .Z(n241) );
  XOR U270 ( .A(n244), .B(n245), .Z(DIFF[487]) );
  XOR U271 ( .A(B[487]), .B(A[487]), .Z(n245) );
  AND U272 ( .A(n246), .B(n247), .Z(n244) );
  NANDN U273 ( .A(B[486]), .B(n248), .Z(n247) );
  NANDN U274 ( .A(A[486]), .B(n249), .Z(n248) );
  NANDN U275 ( .A(n249), .B(A[486]), .Z(n246) );
  XOR U276 ( .A(n249), .B(n250), .Z(DIFF[486]) );
  XOR U277 ( .A(B[486]), .B(A[486]), .Z(n250) );
  AND U278 ( .A(n251), .B(n252), .Z(n249) );
  NANDN U279 ( .A(B[485]), .B(n253), .Z(n252) );
  NANDN U280 ( .A(A[485]), .B(n254), .Z(n253) );
  NANDN U281 ( .A(n254), .B(A[485]), .Z(n251) );
  XOR U282 ( .A(n254), .B(n255), .Z(DIFF[485]) );
  XOR U283 ( .A(B[485]), .B(A[485]), .Z(n255) );
  AND U284 ( .A(n256), .B(n257), .Z(n254) );
  NANDN U285 ( .A(B[484]), .B(n258), .Z(n257) );
  NANDN U286 ( .A(A[484]), .B(n259), .Z(n258) );
  NANDN U287 ( .A(n259), .B(A[484]), .Z(n256) );
  XOR U288 ( .A(n259), .B(n260), .Z(DIFF[484]) );
  XOR U289 ( .A(B[484]), .B(A[484]), .Z(n260) );
  AND U290 ( .A(n261), .B(n262), .Z(n259) );
  NANDN U291 ( .A(B[483]), .B(n263), .Z(n262) );
  NANDN U292 ( .A(A[483]), .B(n264), .Z(n263) );
  NANDN U293 ( .A(n264), .B(A[483]), .Z(n261) );
  XOR U294 ( .A(n264), .B(n265), .Z(DIFF[483]) );
  XOR U295 ( .A(B[483]), .B(A[483]), .Z(n265) );
  AND U296 ( .A(n266), .B(n267), .Z(n264) );
  NANDN U297 ( .A(B[482]), .B(n268), .Z(n267) );
  NANDN U298 ( .A(A[482]), .B(n269), .Z(n268) );
  NANDN U299 ( .A(n269), .B(A[482]), .Z(n266) );
  XOR U300 ( .A(n269), .B(n270), .Z(DIFF[482]) );
  XOR U301 ( .A(B[482]), .B(A[482]), .Z(n270) );
  AND U302 ( .A(n271), .B(n272), .Z(n269) );
  NANDN U303 ( .A(B[481]), .B(n273), .Z(n272) );
  NANDN U304 ( .A(A[481]), .B(n274), .Z(n273) );
  NANDN U305 ( .A(n274), .B(A[481]), .Z(n271) );
  XOR U306 ( .A(n274), .B(n275), .Z(DIFF[481]) );
  XOR U307 ( .A(B[481]), .B(A[481]), .Z(n275) );
  AND U308 ( .A(n276), .B(n277), .Z(n274) );
  NANDN U309 ( .A(B[480]), .B(n278), .Z(n277) );
  NANDN U310 ( .A(A[480]), .B(n279), .Z(n278) );
  NANDN U311 ( .A(n279), .B(A[480]), .Z(n276) );
  XOR U312 ( .A(n279), .B(n280), .Z(DIFF[480]) );
  XOR U313 ( .A(B[480]), .B(A[480]), .Z(n280) );
  AND U314 ( .A(n281), .B(n282), .Z(n279) );
  NANDN U315 ( .A(B[479]), .B(n283), .Z(n282) );
  NANDN U316 ( .A(A[479]), .B(n284), .Z(n283) );
  NANDN U317 ( .A(n284), .B(A[479]), .Z(n281) );
  XOR U318 ( .A(n285), .B(n286), .Z(DIFF[47]) );
  XOR U319 ( .A(B[47]), .B(A[47]), .Z(n286) );
  XOR U320 ( .A(n284), .B(n287), .Z(DIFF[479]) );
  XOR U321 ( .A(B[479]), .B(A[479]), .Z(n287) );
  AND U322 ( .A(n288), .B(n289), .Z(n284) );
  NANDN U323 ( .A(B[478]), .B(n290), .Z(n289) );
  NANDN U324 ( .A(A[478]), .B(n291), .Z(n290) );
  NANDN U325 ( .A(n291), .B(A[478]), .Z(n288) );
  XOR U326 ( .A(n291), .B(n292), .Z(DIFF[478]) );
  XOR U327 ( .A(B[478]), .B(A[478]), .Z(n292) );
  AND U328 ( .A(n293), .B(n294), .Z(n291) );
  NANDN U329 ( .A(B[477]), .B(n295), .Z(n294) );
  NANDN U330 ( .A(A[477]), .B(n296), .Z(n295) );
  NANDN U331 ( .A(n296), .B(A[477]), .Z(n293) );
  XOR U332 ( .A(n296), .B(n297), .Z(DIFF[477]) );
  XOR U333 ( .A(B[477]), .B(A[477]), .Z(n297) );
  AND U334 ( .A(n298), .B(n299), .Z(n296) );
  NANDN U335 ( .A(B[476]), .B(n300), .Z(n299) );
  NANDN U336 ( .A(A[476]), .B(n301), .Z(n300) );
  NANDN U337 ( .A(n301), .B(A[476]), .Z(n298) );
  XOR U338 ( .A(n301), .B(n302), .Z(DIFF[476]) );
  XOR U339 ( .A(B[476]), .B(A[476]), .Z(n302) );
  AND U340 ( .A(n303), .B(n304), .Z(n301) );
  NANDN U341 ( .A(B[475]), .B(n305), .Z(n304) );
  NANDN U342 ( .A(A[475]), .B(n306), .Z(n305) );
  NANDN U343 ( .A(n306), .B(A[475]), .Z(n303) );
  XOR U344 ( .A(n306), .B(n307), .Z(DIFF[475]) );
  XOR U345 ( .A(B[475]), .B(A[475]), .Z(n307) );
  AND U346 ( .A(n308), .B(n309), .Z(n306) );
  NANDN U347 ( .A(B[474]), .B(n310), .Z(n309) );
  NANDN U348 ( .A(A[474]), .B(n311), .Z(n310) );
  NANDN U349 ( .A(n311), .B(A[474]), .Z(n308) );
  XOR U350 ( .A(n311), .B(n312), .Z(DIFF[474]) );
  XOR U351 ( .A(B[474]), .B(A[474]), .Z(n312) );
  AND U352 ( .A(n313), .B(n314), .Z(n311) );
  NANDN U353 ( .A(B[473]), .B(n315), .Z(n314) );
  NANDN U354 ( .A(A[473]), .B(n316), .Z(n315) );
  NANDN U355 ( .A(n316), .B(A[473]), .Z(n313) );
  XOR U356 ( .A(n316), .B(n317), .Z(DIFF[473]) );
  XOR U357 ( .A(B[473]), .B(A[473]), .Z(n317) );
  AND U358 ( .A(n318), .B(n319), .Z(n316) );
  NANDN U359 ( .A(B[472]), .B(n320), .Z(n319) );
  NANDN U360 ( .A(A[472]), .B(n321), .Z(n320) );
  NANDN U361 ( .A(n321), .B(A[472]), .Z(n318) );
  XOR U362 ( .A(n321), .B(n322), .Z(DIFF[472]) );
  XOR U363 ( .A(B[472]), .B(A[472]), .Z(n322) );
  AND U364 ( .A(n323), .B(n324), .Z(n321) );
  NANDN U365 ( .A(B[471]), .B(n325), .Z(n324) );
  NANDN U366 ( .A(A[471]), .B(n326), .Z(n325) );
  NANDN U367 ( .A(n326), .B(A[471]), .Z(n323) );
  XOR U368 ( .A(n326), .B(n327), .Z(DIFF[471]) );
  XOR U369 ( .A(B[471]), .B(A[471]), .Z(n327) );
  AND U370 ( .A(n328), .B(n329), .Z(n326) );
  NANDN U371 ( .A(B[470]), .B(n330), .Z(n329) );
  NANDN U372 ( .A(A[470]), .B(n331), .Z(n330) );
  NANDN U373 ( .A(n331), .B(A[470]), .Z(n328) );
  XOR U374 ( .A(n331), .B(n332), .Z(DIFF[470]) );
  XOR U375 ( .A(B[470]), .B(A[470]), .Z(n332) );
  AND U376 ( .A(n333), .B(n334), .Z(n331) );
  NANDN U377 ( .A(B[469]), .B(n335), .Z(n334) );
  NANDN U378 ( .A(A[469]), .B(n336), .Z(n335) );
  NANDN U379 ( .A(n336), .B(A[469]), .Z(n333) );
  XOR U380 ( .A(n337), .B(n338), .Z(DIFF[46]) );
  XOR U381 ( .A(B[46]), .B(A[46]), .Z(n338) );
  XOR U382 ( .A(n336), .B(n339), .Z(DIFF[469]) );
  XOR U383 ( .A(B[469]), .B(A[469]), .Z(n339) );
  AND U384 ( .A(n340), .B(n341), .Z(n336) );
  NANDN U385 ( .A(B[468]), .B(n342), .Z(n341) );
  NANDN U386 ( .A(A[468]), .B(n343), .Z(n342) );
  NANDN U387 ( .A(n343), .B(A[468]), .Z(n340) );
  XOR U388 ( .A(n343), .B(n344), .Z(DIFF[468]) );
  XOR U389 ( .A(B[468]), .B(A[468]), .Z(n344) );
  AND U390 ( .A(n345), .B(n346), .Z(n343) );
  NANDN U391 ( .A(B[467]), .B(n347), .Z(n346) );
  NANDN U392 ( .A(A[467]), .B(n348), .Z(n347) );
  NANDN U393 ( .A(n348), .B(A[467]), .Z(n345) );
  XOR U394 ( .A(n348), .B(n349), .Z(DIFF[467]) );
  XOR U395 ( .A(B[467]), .B(A[467]), .Z(n349) );
  AND U396 ( .A(n350), .B(n351), .Z(n348) );
  NANDN U397 ( .A(B[466]), .B(n352), .Z(n351) );
  NANDN U398 ( .A(A[466]), .B(n353), .Z(n352) );
  NANDN U399 ( .A(n353), .B(A[466]), .Z(n350) );
  XOR U400 ( .A(n353), .B(n354), .Z(DIFF[466]) );
  XOR U401 ( .A(B[466]), .B(A[466]), .Z(n354) );
  AND U402 ( .A(n355), .B(n356), .Z(n353) );
  NANDN U403 ( .A(B[465]), .B(n357), .Z(n356) );
  NANDN U404 ( .A(A[465]), .B(n358), .Z(n357) );
  NANDN U405 ( .A(n358), .B(A[465]), .Z(n355) );
  XOR U406 ( .A(n358), .B(n359), .Z(DIFF[465]) );
  XOR U407 ( .A(B[465]), .B(A[465]), .Z(n359) );
  AND U408 ( .A(n360), .B(n361), .Z(n358) );
  NANDN U409 ( .A(B[464]), .B(n362), .Z(n361) );
  NANDN U410 ( .A(A[464]), .B(n363), .Z(n362) );
  NANDN U411 ( .A(n363), .B(A[464]), .Z(n360) );
  XOR U412 ( .A(n363), .B(n364), .Z(DIFF[464]) );
  XOR U413 ( .A(B[464]), .B(A[464]), .Z(n364) );
  AND U414 ( .A(n365), .B(n366), .Z(n363) );
  NANDN U415 ( .A(B[463]), .B(n367), .Z(n366) );
  NANDN U416 ( .A(A[463]), .B(n368), .Z(n367) );
  NANDN U417 ( .A(n368), .B(A[463]), .Z(n365) );
  XOR U418 ( .A(n368), .B(n369), .Z(DIFF[463]) );
  XOR U419 ( .A(B[463]), .B(A[463]), .Z(n369) );
  AND U420 ( .A(n370), .B(n371), .Z(n368) );
  NANDN U421 ( .A(B[462]), .B(n372), .Z(n371) );
  NANDN U422 ( .A(A[462]), .B(n373), .Z(n372) );
  NANDN U423 ( .A(n373), .B(A[462]), .Z(n370) );
  XOR U424 ( .A(n373), .B(n374), .Z(DIFF[462]) );
  XOR U425 ( .A(B[462]), .B(A[462]), .Z(n374) );
  AND U426 ( .A(n375), .B(n376), .Z(n373) );
  NANDN U427 ( .A(B[461]), .B(n377), .Z(n376) );
  NANDN U428 ( .A(A[461]), .B(n378), .Z(n377) );
  NANDN U429 ( .A(n378), .B(A[461]), .Z(n375) );
  XOR U430 ( .A(n378), .B(n379), .Z(DIFF[461]) );
  XOR U431 ( .A(B[461]), .B(A[461]), .Z(n379) );
  AND U432 ( .A(n380), .B(n381), .Z(n378) );
  NANDN U433 ( .A(B[460]), .B(n382), .Z(n381) );
  NANDN U434 ( .A(A[460]), .B(n383), .Z(n382) );
  NANDN U435 ( .A(n383), .B(A[460]), .Z(n380) );
  XOR U436 ( .A(n383), .B(n384), .Z(DIFF[460]) );
  XOR U437 ( .A(B[460]), .B(A[460]), .Z(n384) );
  AND U438 ( .A(n385), .B(n386), .Z(n383) );
  NANDN U439 ( .A(B[459]), .B(n387), .Z(n386) );
  NANDN U440 ( .A(A[459]), .B(n388), .Z(n387) );
  NANDN U441 ( .A(n388), .B(A[459]), .Z(n385) );
  XOR U442 ( .A(n389), .B(n390), .Z(DIFF[45]) );
  XOR U443 ( .A(B[45]), .B(A[45]), .Z(n390) );
  XOR U444 ( .A(n388), .B(n391), .Z(DIFF[459]) );
  XOR U445 ( .A(B[459]), .B(A[459]), .Z(n391) );
  AND U446 ( .A(n392), .B(n393), .Z(n388) );
  NANDN U447 ( .A(B[458]), .B(n394), .Z(n393) );
  NANDN U448 ( .A(A[458]), .B(n395), .Z(n394) );
  NANDN U449 ( .A(n395), .B(A[458]), .Z(n392) );
  XOR U450 ( .A(n395), .B(n396), .Z(DIFF[458]) );
  XOR U451 ( .A(B[458]), .B(A[458]), .Z(n396) );
  AND U452 ( .A(n397), .B(n398), .Z(n395) );
  NANDN U453 ( .A(B[457]), .B(n399), .Z(n398) );
  NANDN U454 ( .A(A[457]), .B(n400), .Z(n399) );
  NANDN U455 ( .A(n400), .B(A[457]), .Z(n397) );
  XOR U456 ( .A(n400), .B(n401), .Z(DIFF[457]) );
  XOR U457 ( .A(B[457]), .B(A[457]), .Z(n401) );
  AND U458 ( .A(n402), .B(n403), .Z(n400) );
  NANDN U459 ( .A(B[456]), .B(n404), .Z(n403) );
  NANDN U460 ( .A(A[456]), .B(n405), .Z(n404) );
  NANDN U461 ( .A(n405), .B(A[456]), .Z(n402) );
  XOR U462 ( .A(n405), .B(n406), .Z(DIFF[456]) );
  XOR U463 ( .A(B[456]), .B(A[456]), .Z(n406) );
  AND U464 ( .A(n407), .B(n408), .Z(n405) );
  NANDN U465 ( .A(B[455]), .B(n409), .Z(n408) );
  NANDN U466 ( .A(A[455]), .B(n410), .Z(n409) );
  NANDN U467 ( .A(n410), .B(A[455]), .Z(n407) );
  XOR U468 ( .A(n410), .B(n411), .Z(DIFF[455]) );
  XOR U469 ( .A(B[455]), .B(A[455]), .Z(n411) );
  AND U470 ( .A(n412), .B(n413), .Z(n410) );
  NANDN U471 ( .A(B[454]), .B(n414), .Z(n413) );
  NANDN U472 ( .A(A[454]), .B(n415), .Z(n414) );
  NANDN U473 ( .A(n415), .B(A[454]), .Z(n412) );
  XOR U474 ( .A(n415), .B(n416), .Z(DIFF[454]) );
  XOR U475 ( .A(B[454]), .B(A[454]), .Z(n416) );
  AND U476 ( .A(n417), .B(n418), .Z(n415) );
  NANDN U477 ( .A(B[453]), .B(n419), .Z(n418) );
  NANDN U478 ( .A(A[453]), .B(n420), .Z(n419) );
  NANDN U479 ( .A(n420), .B(A[453]), .Z(n417) );
  XOR U480 ( .A(n420), .B(n421), .Z(DIFF[453]) );
  XOR U481 ( .A(B[453]), .B(A[453]), .Z(n421) );
  AND U482 ( .A(n422), .B(n423), .Z(n420) );
  NANDN U483 ( .A(B[452]), .B(n424), .Z(n423) );
  NANDN U484 ( .A(A[452]), .B(n425), .Z(n424) );
  NANDN U485 ( .A(n425), .B(A[452]), .Z(n422) );
  XOR U486 ( .A(n425), .B(n426), .Z(DIFF[452]) );
  XOR U487 ( .A(B[452]), .B(A[452]), .Z(n426) );
  AND U488 ( .A(n427), .B(n428), .Z(n425) );
  NANDN U489 ( .A(B[451]), .B(n429), .Z(n428) );
  NANDN U490 ( .A(A[451]), .B(n430), .Z(n429) );
  NANDN U491 ( .A(n430), .B(A[451]), .Z(n427) );
  XOR U492 ( .A(n430), .B(n431), .Z(DIFF[451]) );
  XOR U493 ( .A(B[451]), .B(A[451]), .Z(n431) );
  AND U494 ( .A(n432), .B(n433), .Z(n430) );
  NANDN U495 ( .A(B[450]), .B(n434), .Z(n433) );
  NANDN U496 ( .A(A[450]), .B(n435), .Z(n434) );
  NANDN U497 ( .A(n435), .B(A[450]), .Z(n432) );
  XOR U498 ( .A(n435), .B(n436), .Z(DIFF[450]) );
  XOR U499 ( .A(B[450]), .B(A[450]), .Z(n436) );
  AND U500 ( .A(n437), .B(n438), .Z(n435) );
  NANDN U501 ( .A(B[449]), .B(n439), .Z(n438) );
  NANDN U502 ( .A(A[449]), .B(n440), .Z(n439) );
  NANDN U503 ( .A(n440), .B(A[449]), .Z(n437) );
  XOR U504 ( .A(n441), .B(n442), .Z(DIFF[44]) );
  XOR U505 ( .A(B[44]), .B(A[44]), .Z(n442) );
  XOR U506 ( .A(n440), .B(n443), .Z(DIFF[449]) );
  XOR U507 ( .A(B[449]), .B(A[449]), .Z(n443) );
  AND U508 ( .A(n444), .B(n445), .Z(n440) );
  NANDN U509 ( .A(B[448]), .B(n446), .Z(n445) );
  NANDN U510 ( .A(A[448]), .B(n447), .Z(n446) );
  NANDN U511 ( .A(n447), .B(A[448]), .Z(n444) );
  XOR U512 ( .A(n447), .B(n448), .Z(DIFF[448]) );
  XOR U513 ( .A(B[448]), .B(A[448]), .Z(n448) );
  AND U514 ( .A(n449), .B(n450), .Z(n447) );
  NANDN U515 ( .A(B[447]), .B(n451), .Z(n450) );
  NANDN U516 ( .A(A[447]), .B(n452), .Z(n451) );
  NANDN U517 ( .A(n452), .B(A[447]), .Z(n449) );
  XOR U518 ( .A(n452), .B(n453), .Z(DIFF[447]) );
  XOR U519 ( .A(B[447]), .B(A[447]), .Z(n453) );
  AND U520 ( .A(n454), .B(n455), .Z(n452) );
  NANDN U521 ( .A(B[446]), .B(n456), .Z(n455) );
  NANDN U522 ( .A(A[446]), .B(n457), .Z(n456) );
  NANDN U523 ( .A(n457), .B(A[446]), .Z(n454) );
  XOR U524 ( .A(n457), .B(n458), .Z(DIFF[446]) );
  XOR U525 ( .A(B[446]), .B(A[446]), .Z(n458) );
  AND U526 ( .A(n459), .B(n460), .Z(n457) );
  NANDN U527 ( .A(B[445]), .B(n461), .Z(n460) );
  NANDN U528 ( .A(A[445]), .B(n462), .Z(n461) );
  NANDN U529 ( .A(n462), .B(A[445]), .Z(n459) );
  XOR U530 ( .A(n462), .B(n463), .Z(DIFF[445]) );
  XOR U531 ( .A(B[445]), .B(A[445]), .Z(n463) );
  AND U532 ( .A(n464), .B(n465), .Z(n462) );
  NANDN U533 ( .A(B[444]), .B(n466), .Z(n465) );
  NANDN U534 ( .A(A[444]), .B(n467), .Z(n466) );
  NANDN U535 ( .A(n467), .B(A[444]), .Z(n464) );
  XOR U536 ( .A(n467), .B(n468), .Z(DIFF[444]) );
  XOR U537 ( .A(B[444]), .B(A[444]), .Z(n468) );
  AND U538 ( .A(n469), .B(n470), .Z(n467) );
  NANDN U539 ( .A(B[443]), .B(n471), .Z(n470) );
  NANDN U540 ( .A(A[443]), .B(n472), .Z(n471) );
  NANDN U541 ( .A(n472), .B(A[443]), .Z(n469) );
  XOR U542 ( .A(n472), .B(n473), .Z(DIFF[443]) );
  XOR U543 ( .A(B[443]), .B(A[443]), .Z(n473) );
  AND U544 ( .A(n474), .B(n475), .Z(n472) );
  NANDN U545 ( .A(B[442]), .B(n476), .Z(n475) );
  NANDN U546 ( .A(A[442]), .B(n477), .Z(n476) );
  NANDN U547 ( .A(n477), .B(A[442]), .Z(n474) );
  XOR U548 ( .A(n477), .B(n478), .Z(DIFF[442]) );
  XOR U549 ( .A(B[442]), .B(A[442]), .Z(n478) );
  AND U550 ( .A(n479), .B(n480), .Z(n477) );
  NANDN U551 ( .A(B[441]), .B(n481), .Z(n480) );
  NANDN U552 ( .A(A[441]), .B(n482), .Z(n481) );
  NANDN U553 ( .A(n482), .B(A[441]), .Z(n479) );
  XOR U554 ( .A(n482), .B(n483), .Z(DIFF[441]) );
  XOR U555 ( .A(B[441]), .B(A[441]), .Z(n483) );
  AND U556 ( .A(n484), .B(n485), .Z(n482) );
  NANDN U557 ( .A(B[440]), .B(n486), .Z(n485) );
  NANDN U558 ( .A(A[440]), .B(n487), .Z(n486) );
  NANDN U559 ( .A(n487), .B(A[440]), .Z(n484) );
  XOR U560 ( .A(n487), .B(n488), .Z(DIFF[440]) );
  XOR U561 ( .A(B[440]), .B(A[440]), .Z(n488) );
  AND U562 ( .A(n489), .B(n490), .Z(n487) );
  NANDN U563 ( .A(B[439]), .B(n491), .Z(n490) );
  NANDN U564 ( .A(A[439]), .B(n492), .Z(n491) );
  NANDN U565 ( .A(n492), .B(A[439]), .Z(n489) );
  XOR U566 ( .A(n493), .B(n494), .Z(DIFF[43]) );
  XOR U567 ( .A(B[43]), .B(A[43]), .Z(n494) );
  XOR U568 ( .A(n492), .B(n495), .Z(DIFF[439]) );
  XOR U569 ( .A(B[439]), .B(A[439]), .Z(n495) );
  AND U570 ( .A(n496), .B(n497), .Z(n492) );
  NANDN U571 ( .A(B[438]), .B(n498), .Z(n497) );
  NANDN U572 ( .A(A[438]), .B(n499), .Z(n498) );
  NANDN U573 ( .A(n499), .B(A[438]), .Z(n496) );
  XOR U574 ( .A(n499), .B(n500), .Z(DIFF[438]) );
  XOR U575 ( .A(B[438]), .B(A[438]), .Z(n500) );
  AND U576 ( .A(n501), .B(n502), .Z(n499) );
  NANDN U577 ( .A(B[437]), .B(n503), .Z(n502) );
  NANDN U578 ( .A(A[437]), .B(n504), .Z(n503) );
  NANDN U579 ( .A(n504), .B(A[437]), .Z(n501) );
  XOR U580 ( .A(n504), .B(n505), .Z(DIFF[437]) );
  XOR U581 ( .A(B[437]), .B(A[437]), .Z(n505) );
  AND U582 ( .A(n506), .B(n507), .Z(n504) );
  NANDN U583 ( .A(B[436]), .B(n508), .Z(n507) );
  NANDN U584 ( .A(A[436]), .B(n509), .Z(n508) );
  NANDN U585 ( .A(n509), .B(A[436]), .Z(n506) );
  XOR U586 ( .A(n509), .B(n510), .Z(DIFF[436]) );
  XOR U587 ( .A(B[436]), .B(A[436]), .Z(n510) );
  AND U588 ( .A(n511), .B(n512), .Z(n509) );
  NANDN U589 ( .A(B[435]), .B(n513), .Z(n512) );
  NANDN U590 ( .A(A[435]), .B(n514), .Z(n513) );
  NANDN U591 ( .A(n514), .B(A[435]), .Z(n511) );
  XOR U592 ( .A(n514), .B(n515), .Z(DIFF[435]) );
  XOR U593 ( .A(B[435]), .B(A[435]), .Z(n515) );
  AND U594 ( .A(n516), .B(n517), .Z(n514) );
  NANDN U595 ( .A(B[434]), .B(n518), .Z(n517) );
  NANDN U596 ( .A(A[434]), .B(n519), .Z(n518) );
  NANDN U597 ( .A(n519), .B(A[434]), .Z(n516) );
  XOR U598 ( .A(n519), .B(n520), .Z(DIFF[434]) );
  XOR U599 ( .A(B[434]), .B(A[434]), .Z(n520) );
  AND U600 ( .A(n521), .B(n522), .Z(n519) );
  NANDN U601 ( .A(B[433]), .B(n523), .Z(n522) );
  NANDN U602 ( .A(A[433]), .B(n524), .Z(n523) );
  NANDN U603 ( .A(n524), .B(A[433]), .Z(n521) );
  XOR U604 ( .A(n524), .B(n525), .Z(DIFF[433]) );
  XOR U605 ( .A(B[433]), .B(A[433]), .Z(n525) );
  AND U606 ( .A(n526), .B(n527), .Z(n524) );
  NANDN U607 ( .A(B[432]), .B(n528), .Z(n527) );
  NANDN U608 ( .A(A[432]), .B(n529), .Z(n528) );
  NANDN U609 ( .A(n529), .B(A[432]), .Z(n526) );
  XOR U610 ( .A(n529), .B(n530), .Z(DIFF[432]) );
  XOR U611 ( .A(B[432]), .B(A[432]), .Z(n530) );
  AND U612 ( .A(n531), .B(n532), .Z(n529) );
  NANDN U613 ( .A(B[431]), .B(n533), .Z(n532) );
  NANDN U614 ( .A(A[431]), .B(n534), .Z(n533) );
  NANDN U615 ( .A(n534), .B(A[431]), .Z(n531) );
  XOR U616 ( .A(n534), .B(n535), .Z(DIFF[431]) );
  XOR U617 ( .A(B[431]), .B(A[431]), .Z(n535) );
  AND U618 ( .A(n536), .B(n537), .Z(n534) );
  NANDN U619 ( .A(B[430]), .B(n538), .Z(n537) );
  NANDN U620 ( .A(A[430]), .B(n539), .Z(n538) );
  NANDN U621 ( .A(n539), .B(A[430]), .Z(n536) );
  XOR U622 ( .A(n539), .B(n540), .Z(DIFF[430]) );
  XOR U623 ( .A(B[430]), .B(A[430]), .Z(n540) );
  AND U624 ( .A(n541), .B(n542), .Z(n539) );
  NANDN U625 ( .A(B[429]), .B(n543), .Z(n542) );
  NANDN U626 ( .A(A[429]), .B(n544), .Z(n543) );
  NANDN U627 ( .A(n544), .B(A[429]), .Z(n541) );
  XOR U628 ( .A(n545), .B(n546), .Z(DIFF[42]) );
  XOR U629 ( .A(B[42]), .B(A[42]), .Z(n546) );
  XOR U630 ( .A(n544), .B(n547), .Z(DIFF[429]) );
  XOR U631 ( .A(B[429]), .B(A[429]), .Z(n547) );
  AND U632 ( .A(n548), .B(n549), .Z(n544) );
  NANDN U633 ( .A(B[428]), .B(n550), .Z(n549) );
  NANDN U634 ( .A(A[428]), .B(n551), .Z(n550) );
  NANDN U635 ( .A(n551), .B(A[428]), .Z(n548) );
  XOR U636 ( .A(n551), .B(n552), .Z(DIFF[428]) );
  XOR U637 ( .A(B[428]), .B(A[428]), .Z(n552) );
  AND U638 ( .A(n553), .B(n554), .Z(n551) );
  NANDN U639 ( .A(B[427]), .B(n555), .Z(n554) );
  NANDN U640 ( .A(A[427]), .B(n556), .Z(n555) );
  NANDN U641 ( .A(n556), .B(A[427]), .Z(n553) );
  XOR U642 ( .A(n556), .B(n557), .Z(DIFF[427]) );
  XOR U643 ( .A(B[427]), .B(A[427]), .Z(n557) );
  AND U644 ( .A(n558), .B(n559), .Z(n556) );
  NANDN U645 ( .A(B[426]), .B(n560), .Z(n559) );
  NANDN U646 ( .A(A[426]), .B(n561), .Z(n560) );
  NANDN U647 ( .A(n561), .B(A[426]), .Z(n558) );
  XOR U648 ( .A(n561), .B(n562), .Z(DIFF[426]) );
  XOR U649 ( .A(B[426]), .B(A[426]), .Z(n562) );
  AND U650 ( .A(n563), .B(n564), .Z(n561) );
  NANDN U651 ( .A(B[425]), .B(n565), .Z(n564) );
  NANDN U652 ( .A(A[425]), .B(n566), .Z(n565) );
  NANDN U653 ( .A(n566), .B(A[425]), .Z(n563) );
  XOR U654 ( .A(n566), .B(n567), .Z(DIFF[425]) );
  XOR U655 ( .A(B[425]), .B(A[425]), .Z(n567) );
  AND U656 ( .A(n568), .B(n569), .Z(n566) );
  NANDN U657 ( .A(B[424]), .B(n570), .Z(n569) );
  NANDN U658 ( .A(A[424]), .B(n571), .Z(n570) );
  NANDN U659 ( .A(n571), .B(A[424]), .Z(n568) );
  XOR U660 ( .A(n571), .B(n572), .Z(DIFF[424]) );
  XOR U661 ( .A(B[424]), .B(A[424]), .Z(n572) );
  AND U662 ( .A(n573), .B(n574), .Z(n571) );
  NANDN U663 ( .A(B[423]), .B(n575), .Z(n574) );
  NANDN U664 ( .A(A[423]), .B(n576), .Z(n575) );
  NANDN U665 ( .A(n576), .B(A[423]), .Z(n573) );
  XOR U666 ( .A(n576), .B(n577), .Z(DIFF[423]) );
  XOR U667 ( .A(B[423]), .B(A[423]), .Z(n577) );
  AND U668 ( .A(n578), .B(n579), .Z(n576) );
  NANDN U669 ( .A(B[422]), .B(n580), .Z(n579) );
  NANDN U670 ( .A(A[422]), .B(n581), .Z(n580) );
  NANDN U671 ( .A(n581), .B(A[422]), .Z(n578) );
  XOR U672 ( .A(n581), .B(n582), .Z(DIFF[422]) );
  XOR U673 ( .A(B[422]), .B(A[422]), .Z(n582) );
  AND U674 ( .A(n583), .B(n584), .Z(n581) );
  NANDN U675 ( .A(B[421]), .B(n585), .Z(n584) );
  NANDN U676 ( .A(A[421]), .B(n586), .Z(n585) );
  NANDN U677 ( .A(n586), .B(A[421]), .Z(n583) );
  XOR U678 ( .A(n586), .B(n587), .Z(DIFF[421]) );
  XOR U679 ( .A(B[421]), .B(A[421]), .Z(n587) );
  AND U680 ( .A(n588), .B(n589), .Z(n586) );
  NANDN U681 ( .A(B[420]), .B(n590), .Z(n589) );
  NANDN U682 ( .A(A[420]), .B(n591), .Z(n590) );
  NANDN U683 ( .A(n591), .B(A[420]), .Z(n588) );
  XOR U684 ( .A(n591), .B(n592), .Z(DIFF[420]) );
  XOR U685 ( .A(B[420]), .B(A[420]), .Z(n592) );
  AND U686 ( .A(n593), .B(n594), .Z(n591) );
  NANDN U687 ( .A(B[419]), .B(n595), .Z(n594) );
  NANDN U688 ( .A(A[419]), .B(n596), .Z(n595) );
  NANDN U689 ( .A(n596), .B(A[419]), .Z(n593) );
  XOR U690 ( .A(n597), .B(n598), .Z(DIFF[41]) );
  XOR U691 ( .A(B[41]), .B(A[41]), .Z(n598) );
  XOR U692 ( .A(n596), .B(n599), .Z(DIFF[419]) );
  XOR U693 ( .A(B[419]), .B(A[419]), .Z(n599) );
  AND U694 ( .A(n600), .B(n601), .Z(n596) );
  NANDN U695 ( .A(B[418]), .B(n602), .Z(n601) );
  NANDN U696 ( .A(A[418]), .B(n603), .Z(n602) );
  NANDN U697 ( .A(n603), .B(A[418]), .Z(n600) );
  XOR U698 ( .A(n603), .B(n604), .Z(DIFF[418]) );
  XOR U699 ( .A(B[418]), .B(A[418]), .Z(n604) );
  AND U700 ( .A(n605), .B(n606), .Z(n603) );
  NANDN U701 ( .A(B[417]), .B(n607), .Z(n606) );
  NANDN U702 ( .A(A[417]), .B(n608), .Z(n607) );
  NANDN U703 ( .A(n608), .B(A[417]), .Z(n605) );
  XOR U704 ( .A(n608), .B(n609), .Z(DIFF[417]) );
  XOR U705 ( .A(B[417]), .B(A[417]), .Z(n609) );
  AND U706 ( .A(n610), .B(n611), .Z(n608) );
  NANDN U707 ( .A(B[416]), .B(n612), .Z(n611) );
  NANDN U708 ( .A(A[416]), .B(n613), .Z(n612) );
  NANDN U709 ( .A(n613), .B(A[416]), .Z(n610) );
  XOR U710 ( .A(n613), .B(n614), .Z(DIFF[416]) );
  XOR U711 ( .A(B[416]), .B(A[416]), .Z(n614) );
  AND U712 ( .A(n615), .B(n616), .Z(n613) );
  NANDN U713 ( .A(B[415]), .B(n617), .Z(n616) );
  NANDN U714 ( .A(A[415]), .B(n618), .Z(n617) );
  NANDN U715 ( .A(n618), .B(A[415]), .Z(n615) );
  XOR U716 ( .A(n618), .B(n619), .Z(DIFF[415]) );
  XOR U717 ( .A(B[415]), .B(A[415]), .Z(n619) );
  AND U718 ( .A(n620), .B(n621), .Z(n618) );
  NANDN U719 ( .A(B[414]), .B(n622), .Z(n621) );
  NANDN U720 ( .A(A[414]), .B(n623), .Z(n622) );
  NANDN U721 ( .A(n623), .B(A[414]), .Z(n620) );
  XOR U722 ( .A(n623), .B(n624), .Z(DIFF[414]) );
  XOR U723 ( .A(B[414]), .B(A[414]), .Z(n624) );
  AND U724 ( .A(n625), .B(n626), .Z(n623) );
  NANDN U725 ( .A(B[413]), .B(n627), .Z(n626) );
  NANDN U726 ( .A(A[413]), .B(n628), .Z(n627) );
  NANDN U727 ( .A(n628), .B(A[413]), .Z(n625) );
  XOR U728 ( .A(n628), .B(n629), .Z(DIFF[413]) );
  XOR U729 ( .A(B[413]), .B(A[413]), .Z(n629) );
  AND U730 ( .A(n630), .B(n631), .Z(n628) );
  NANDN U731 ( .A(B[412]), .B(n632), .Z(n631) );
  NANDN U732 ( .A(A[412]), .B(n633), .Z(n632) );
  NANDN U733 ( .A(n633), .B(A[412]), .Z(n630) );
  XOR U734 ( .A(n633), .B(n634), .Z(DIFF[412]) );
  XOR U735 ( .A(B[412]), .B(A[412]), .Z(n634) );
  AND U736 ( .A(n635), .B(n636), .Z(n633) );
  NANDN U737 ( .A(B[411]), .B(n637), .Z(n636) );
  NANDN U738 ( .A(A[411]), .B(n638), .Z(n637) );
  NANDN U739 ( .A(n638), .B(A[411]), .Z(n635) );
  XOR U740 ( .A(n638), .B(n639), .Z(DIFF[411]) );
  XOR U741 ( .A(B[411]), .B(A[411]), .Z(n639) );
  AND U742 ( .A(n640), .B(n641), .Z(n638) );
  NANDN U743 ( .A(B[410]), .B(n642), .Z(n641) );
  NANDN U744 ( .A(A[410]), .B(n643), .Z(n642) );
  NANDN U745 ( .A(n643), .B(A[410]), .Z(n640) );
  XOR U746 ( .A(n643), .B(n644), .Z(DIFF[410]) );
  XOR U747 ( .A(B[410]), .B(A[410]), .Z(n644) );
  AND U748 ( .A(n645), .B(n646), .Z(n643) );
  NANDN U749 ( .A(B[409]), .B(n647), .Z(n646) );
  NANDN U750 ( .A(A[409]), .B(n648), .Z(n647) );
  NANDN U751 ( .A(n648), .B(A[409]), .Z(n645) );
  XOR U752 ( .A(n649), .B(n650), .Z(DIFF[40]) );
  XOR U753 ( .A(B[40]), .B(A[40]), .Z(n650) );
  XOR U754 ( .A(n648), .B(n651), .Z(DIFF[409]) );
  XOR U755 ( .A(B[409]), .B(A[409]), .Z(n651) );
  AND U756 ( .A(n652), .B(n653), .Z(n648) );
  NANDN U757 ( .A(B[408]), .B(n654), .Z(n653) );
  NANDN U758 ( .A(A[408]), .B(n655), .Z(n654) );
  NANDN U759 ( .A(n655), .B(A[408]), .Z(n652) );
  XOR U760 ( .A(n655), .B(n656), .Z(DIFF[408]) );
  XOR U761 ( .A(B[408]), .B(A[408]), .Z(n656) );
  AND U762 ( .A(n657), .B(n658), .Z(n655) );
  NANDN U763 ( .A(B[407]), .B(n659), .Z(n658) );
  NANDN U764 ( .A(A[407]), .B(n660), .Z(n659) );
  NANDN U765 ( .A(n660), .B(A[407]), .Z(n657) );
  XOR U766 ( .A(n660), .B(n661), .Z(DIFF[407]) );
  XOR U767 ( .A(B[407]), .B(A[407]), .Z(n661) );
  AND U768 ( .A(n662), .B(n663), .Z(n660) );
  NANDN U769 ( .A(B[406]), .B(n664), .Z(n663) );
  NANDN U770 ( .A(A[406]), .B(n665), .Z(n664) );
  NANDN U771 ( .A(n665), .B(A[406]), .Z(n662) );
  XOR U772 ( .A(n665), .B(n666), .Z(DIFF[406]) );
  XOR U773 ( .A(B[406]), .B(A[406]), .Z(n666) );
  AND U774 ( .A(n667), .B(n668), .Z(n665) );
  NANDN U775 ( .A(B[405]), .B(n669), .Z(n668) );
  NANDN U776 ( .A(A[405]), .B(n670), .Z(n669) );
  NANDN U777 ( .A(n670), .B(A[405]), .Z(n667) );
  XOR U778 ( .A(n670), .B(n671), .Z(DIFF[405]) );
  XOR U779 ( .A(B[405]), .B(A[405]), .Z(n671) );
  AND U780 ( .A(n672), .B(n673), .Z(n670) );
  NANDN U781 ( .A(B[404]), .B(n674), .Z(n673) );
  NANDN U782 ( .A(A[404]), .B(n675), .Z(n674) );
  NANDN U783 ( .A(n675), .B(A[404]), .Z(n672) );
  XOR U784 ( .A(n675), .B(n676), .Z(DIFF[404]) );
  XOR U785 ( .A(B[404]), .B(A[404]), .Z(n676) );
  AND U786 ( .A(n677), .B(n678), .Z(n675) );
  NANDN U787 ( .A(B[403]), .B(n679), .Z(n678) );
  NANDN U788 ( .A(A[403]), .B(n680), .Z(n679) );
  NANDN U789 ( .A(n680), .B(A[403]), .Z(n677) );
  XOR U790 ( .A(n680), .B(n681), .Z(DIFF[403]) );
  XOR U791 ( .A(B[403]), .B(A[403]), .Z(n681) );
  AND U792 ( .A(n682), .B(n683), .Z(n680) );
  NANDN U793 ( .A(B[402]), .B(n684), .Z(n683) );
  NANDN U794 ( .A(A[402]), .B(n685), .Z(n684) );
  NANDN U795 ( .A(n685), .B(A[402]), .Z(n682) );
  XOR U796 ( .A(n685), .B(n686), .Z(DIFF[402]) );
  XOR U797 ( .A(B[402]), .B(A[402]), .Z(n686) );
  AND U798 ( .A(n687), .B(n688), .Z(n685) );
  NANDN U799 ( .A(B[401]), .B(n689), .Z(n688) );
  NANDN U800 ( .A(A[401]), .B(n690), .Z(n689) );
  NANDN U801 ( .A(n690), .B(A[401]), .Z(n687) );
  XOR U802 ( .A(n690), .B(n691), .Z(DIFF[401]) );
  XOR U803 ( .A(B[401]), .B(A[401]), .Z(n691) );
  AND U804 ( .A(n692), .B(n693), .Z(n690) );
  NANDN U805 ( .A(B[400]), .B(n694), .Z(n693) );
  NANDN U806 ( .A(A[400]), .B(n695), .Z(n694) );
  NANDN U807 ( .A(n695), .B(A[400]), .Z(n692) );
  XOR U808 ( .A(n695), .B(n696), .Z(DIFF[400]) );
  XOR U809 ( .A(B[400]), .B(A[400]), .Z(n696) );
  AND U810 ( .A(n697), .B(n698), .Z(n695) );
  NANDN U811 ( .A(B[399]), .B(n699), .Z(n698) );
  NANDN U812 ( .A(A[399]), .B(n700), .Z(n699) );
  NANDN U813 ( .A(n700), .B(A[399]), .Z(n697) );
  XOR U814 ( .A(n701), .B(n702), .Z(DIFF[3]) );
  XOR U815 ( .A(B[3]), .B(A[3]), .Z(n702) );
  XOR U816 ( .A(n703), .B(n704), .Z(DIFF[39]) );
  XOR U817 ( .A(B[39]), .B(A[39]), .Z(n704) );
  XOR U818 ( .A(n700), .B(n705), .Z(DIFF[399]) );
  XOR U819 ( .A(B[399]), .B(A[399]), .Z(n705) );
  AND U820 ( .A(n706), .B(n707), .Z(n700) );
  NANDN U821 ( .A(B[398]), .B(n708), .Z(n707) );
  NANDN U822 ( .A(A[398]), .B(n709), .Z(n708) );
  NANDN U823 ( .A(n709), .B(A[398]), .Z(n706) );
  XOR U824 ( .A(n709), .B(n710), .Z(DIFF[398]) );
  XOR U825 ( .A(B[398]), .B(A[398]), .Z(n710) );
  AND U826 ( .A(n711), .B(n712), .Z(n709) );
  NANDN U827 ( .A(B[397]), .B(n713), .Z(n712) );
  NANDN U828 ( .A(A[397]), .B(n714), .Z(n713) );
  NANDN U829 ( .A(n714), .B(A[397]), .Z(n711) );
  XOR U830 ( .A(n714), .B(n715), .Z(DIFF[397]) );
  XOR U831 ( .A(B[397]), .B(A[397]), .Z(n715) );
  AND U832 ( .A(n716), .B(n717), .Z(n714) );
  NANDN U833 ( .A(B[396]), .B(n718), .Z(n717) );
  NANDN U834 ( .A(A[396]), .B(n719), .Z(n718) );
  NANDN U835 ( .A(n719), .B(A[396]), .Z(n716) );
  XOR U836 ( .A(n719), .B(n720), .Z(DIFF[396]) );
  XOR U837 ( .A(B[396]), .B(A[396]), .Z(n720) );
  AND U838 ( .A(n721), .B(n722), .Z(n719) );
  NANDN U839 ( .A(B[395]), .B(n723), .Z(n722) );
  NANDN U840 ( .A(A[395]), .B(n724), .Z(n723) );
  NANDN U841 ( .A(n724), .B(A[395]), .Z(n721) );
  XOR U842 ( .A(n724), .B(n725), .Z(DIFF[395]) );
  XOR U843 ( .A(B[395]), .B(A[395]), .Z(n725) );
  AND U844 ( .A(n726), .B(n727), .Z(n724) );
  NANDN U845 ( .A(B[394]), .B(n728), .Z(n727) );
  NANDN U846 ( .A(A[394]), .B(n729), .Z(n728) );
  NANDN U847 ( .A(n729), .B(A[394]), .Z(n726) );
  XOR U848 ( .A(n729), .B(n730), .Z(DIFF[394]) );
  XOR U849 ( .A(B[394]), .B(A[394]), .Z(n730) );
  AND U850 ( .A(n731), .B(n732), .Z(n729) );
  NANDN U851 ( .A(B[393]), .B(n733), .Z(n732) );
  NANDN U852 ( .A(A[393]), .B(n734), .Z(n733) );
  NANDN U853 ( .A(n734), .B(A[393]), .Z(n731) );
  XOR U854 ( .A(n734), .B(n735), .Z(DIFF[393]) );
  XOR U855 ( .A(B[393]), .B(A[393]), .Z(n735) );
  AND U856 ( .A(n736), .B(n737), .Z(n734) );
  NANDN U857 ( .A(B[392]), .B(n738), .Z(n737) );
  NANDN U858 ( .A(A[392]), .B(n739), .Z(n738) );
  NANDN U859 ( .A(n739), .B(A[392]), .Z(n736) );
  XOR U860 ( .A(n739), .B(n740), .Z(DIFF[392]) );
  XOR U861 ( .A(B[392]), .B(A[392]), .Z(n740) );
  AND U862 ( .A(n741), .B(n742), .Z(n739) );
  NANDN U863 ( .A(B[391]), .B(n743), .Z(n742) );
  NANDN U864 ( .A(A[391]), .B(n744), .Z(n743) );
  NANDN U865 ( .A(n744), .B(A[391]), .Z(n741) );
  XOR U866 ( .A(n744), .B(n745), .Z(DIFF[391]) );
  XOR U867 ( .A(B[391]), .B(A[391]), .Z(n745) );
  AND U868 ( .A(n746), .B(n747), .Z(n744) );
  NANDN U869 ( .A(B[390]), .B(n748), .Z(n747) );
  NANDN U870 ( .A(A[390]), .B(n749), .Z(n748) );
  NANDN U871 ( .A(n749), .B(A[390]), .Z(n746) );
  XOR U872 ( .A(n749), .B(n750), .Z(DIFF[390]) );
  XOR U873 ( .A(B[390]), .B(A[390]), .Z(n750) );
  AND U874 ( .A(n751), .B(n752), .Z(n749) );
  NANDN U875 ( .A(B[389]), .B(n753), .Z(n752) );
  NANDN U876 ( .A(A[389]), .B(n754), .Z(n753) );
  NANDN U877 ( .A(n754), .B(A[389]), .Z(n751) );
  XOR U878 ( .A(n755), .B(n756), .Z(DIFF[38]) );
  XOR U879 ( .A(B[38]), .B(A[38]), .Z(n756) );
  XOR U880 ( .A(n754), .B(n757), .Z(DIFF[389]) );
  XOR U881 ( .A(B[389]), .B(A[389]), .Z(n757) );
  AND U882 ( .A(n758), .B(n759), .Z(n754) );
  NANDN U883 ( .A(B[388]), .B(n760), .Z(n759) );
  NANDN U884 ( .A(A[388]), .B(n761), .Z(n760) );
  NANDN U885 ( .A(n761), .B(A[388]), .Z(n758) );
  XOR U886 ( .A(n761), .B(n762), .Z(DIFF[388]) );
  XOR U887 ( .A(B[388]), .B(A[388]), .Z(n762) );
  AND U888 ( .A(n763), .B(n764), .Z(n761) );
  NANDN U889 ( .A(B[387]), .B(n765), .Z(n764) );
  NANDN U890 ( .A(A[387]), .B(n766), .Z(n765) );
  NANDN U891 ( .A(n766), .B(A[387]), .Z(n763) );
  XOR U892 ( .A(n766), .B(n767), .Z(DIFF[387]) );
  XOR U893 ( .A(B[387]), .B(A[387]), .Z(n767) );
  AND U894 ( .A(n768), .B(n769), .Z(n766) );
  NANDN U895 ( .A(B[386]), .B(n770), .Z(n769) );
  NANDN U896 ( .A(A[386]), .B(n771), .Z(n770) );
  NANDN U897 ( .A(n771), .B(A[386]), .Z(n768) );
  XOR U898 ( .A(n771), .B(n772), .Z(DIFF[386]) );
  XOR U899 ( .A(B[386]), .B(A[386]), .Z(n772) );
  AND U900 ( .A(n773), .B(n774), .Z(n771) );
  NANDN U901 ( .A(B[385]), .B(n775), .Z(n774) );
  NANDN U902 ( .A(A[385]), .B(n776), .Z(n775) );
  NANDN U903 ( .A(n776), .B(A[385]), .Z(n773) );
  XOR U904 ( .A(n776), .B(n777), .Z(DIFF[385]) );
  XOR U905 ( .A(B[385]), .B(A[385]), .Z(n777) );
  AND U906 ( .A(n778), .B(n779), .Z(n776) );
  NANDN U907 ( .A(B[384]), .B(n780), .Z(n779) );
  NANDN U908 ( .A(A[384]), .B(n781), .Z(n780) );
  NANDN U909 ( .A(n781), .B(A[384]), .Z(n778) );
  XOR U910 ( .A(n781), .B(n782), .Z(DIFF[384]) );
  XOR U911 ( .A(B[384]), .B(A[384]), .Z(n782) );
  AND U912 ( .A(n783), .B(n784), .Z(n781) );
  NANDN U913 ( .A(B[383]), .B(n785), .Z(n784) );
  NANDN U914 ( .A(A[383]), .B(n786), .Z(n785) );
  NANDN U915 ( .A(n786), .B(A[383]), .Z(n783) );
  XOR U916 ( .A(n786), .B(n787), .Z(DIFF[383]) );
  XOR U917 ( .A(B[383]), .B(A[383]), .Z(n787) );
  AND U918 ( .A(n788), .B(n789), .Z(n786) );
  NANDN U919 ( .A(B[382]), .B(n790), .Z(n789) );
  NANDN U920 ( .A(A[382]), .B(n791), .Z(n790) );
  NANDN U921 ( .A(n791), .B(A[382]), .Z(n788) );
  XOR U922 ( .A(n791), .B(n792), .Z(DIFF[382]) );
  XOR U923 ( .A(B[382]), .B(A[382]), .Z(n792) );
  AND U924 ( .A(n793), .B(n794), .Z(n791) );
  NANDN U925 ( .A(B[381]), .B(n795), .Z(n794) );
  NANDN U926 ( .A(A[381]), .B(n796), .Z(n795) );
  NANDN U927 ( .A(n796), .B(A[381]), .Z(n793) );
  XOR U928 ( .A(n796), .B(n797), .Z(DIFF[381]) );
  XOR U929 ( .A(B[381]), .B(A[381]), .Z(n797) );
  AND U930 ( .A(n798), .B(n799), .Z(n796) );
  NANDN U931 ( .A(B[380]), .B(n800), .Z(n799) );
  NANDN U932 ( .A(A[380]), .B(n801), .Z(n800) );
  NANDN U933 ( .A(n801), .B(A[380]), .Z(n798) );
  XOR U934 ( .A(n801), .B(n802), .Z(DIFF[380]) );
  XOR U935 ( .A(B[380]), .B(A[380]), .Z(n802) );
  AND U936 ( .A(n803), .B(n804), .Z(n801) );
  NANDN U937 ( .A(B[379]), .B(n805), .Z(n804) );
  NANDN U938 ( .A(A[379]), .B(n806), .Z(n805) );
  NANDN U939 ( .A(n806), .B(A[379]), .Z(n803) );
  XOR U940 ( .A(n807), .B(n808), .Z(DIFF[37]) );
  XOR U941 ( .A(B[37]), .B(A[37]), .Z(n808) );
  XOR U942 ( .A(n806), .B(n809), .Z(DIFF[379]) );
  XOR U943 ( .A(B[379]), .B(A[379]), .Z(n809) );
  AND U944 ( .A(n810), .B(n811), .Z(n806) );
  NANDN U945 ( .A(B[378]), .B(n812), .Z(n811) );
  NANDN U946 ( .A(A[378]), .B(n813), .Z(n812) );
  NANDN U947 ( .A(n813), .B(A[378]), .Z(n810) );
  XOR U948 ( .A(n813), .B(n814), .Z(DIFF[378]) );
  XOR U949 ( .A(B[378]), .B(A[378]), .Z(n814) );
  AND U950 ( .A(n815), .B(n816), .Z(n813) );
  NANDN U951 ( .A(B[377]), .B(n817), .Z(n816) );
  NANDN U952 ( .A(A[377]), .B(n818), .Z(n817) );
  NANDN U953 ( .A(n818), .B(A[377]), .Z(n815) );
  XOR U954 ( .A(n818), .B(n819), .Z(DIFF[377]) );
  XOR U955 ( .A(B[377]), .B(A[377]), .Z(n819) );
  AND U956 ( .A(n820), .B(n821), .Z(n818) );
  NANDN U957 ( .A(B[376]), .B(n822), .Z(n821) );
  NANDN U958 ( .A(A[376]), .B(n823), .Z(n822) );
  NANDN U959 ( .A(n823), .B(A[376]), .Z(n820) );
  XOR U960 ( .A(n823), .B(n824), .Z(DIFF[376]) );
  XOR U961 ( .A(B[376]), .B(A[376]), .Z(n824) );
  AND U962 ( .A(n825), .B(n826), .Z(n823) );
  NANDN U963 ( .A(B[375]), .B(n827), .Z(n826) );
  NANDN U964 ( .A(A[375]), .B(n828), .Z(n827) );
  NANDN U965 ( .A(n828), .B(A[375]), .Z(n825) );
  XOR U966 ( .A(n828), .B(n829), .Z(DIFF[375]) );
  XOR U967 ( .A(B[375]), .B(A[375]), .Z(n829) );
  AND U968 ( .A(n830), .B(n831), .Z(n828) );
  NANDN U969 ( .A(B[374]), .B(n832), .Z(n831) );
  NANDN U970 ( .A(A[374]), .B(n833), .Z(n832) );
  NANDN U971 ( .A(n833), .B(A[374]), .Z(n830) );
  XOR U972 ( .A(n833), .B(n834), .Z(DIFF[374]) );
  XOR U973 ( .A(B[374]), .B(A[374]), .Z(n834) );
  AND U974 ( .A(n835), .B(n836), .Z(n833) );
  NANDN U975 ( .A(B[373]), .B(n837), .Z(n836) );
  NANDN U976 ( .A(A[373]), .B(n838), .Z(n837) );
  NANDN U977 ( .A(n838), .B(A[373]), .Z(n835) );
  XOR U978 ( .A(n838), .B(n839), .Z(DIFF[373]) );
  XOR U979 ( .A(B[373]), .B(A[373]), .Z(n839) );
  AND U980 ( .A(n840), .B(n841), .Z(n838) );
  NANDN U981 ( .A(B[372]), .B(n842), .Z(n841) );
  NANDN U982 ( .A(A[372]), .B(n843), .Z(n842) );
  NANDN U983 ( .A(n843), .B(A[372]), .Z(n840) );
  XOR U984 ( .A(n843), .B(n844), .Z(DIFF[372]) );
  XOR U985 ( .A(B[372]), .B(A[372]), .Z(n844) );
  AND U986 ( .A(n845), .B(n846), .Z(n843) );
  NANDN U987 ( .A(B[371]), .B(n847), .Z(n846) );
  NANDN U988 ( .A(A[371]), .B(n848), .Z(n847) );
  NANDN U989 ( .A(n848), .B(A[371]), .Z(n845) );
  XOR U990 ( .A(n848), .B(n849), .Z(DIFF[371]) );
  XOR U991 ( .A(B[371]), .B(A[371]), .Z(n849) );
  AND U992 ( .A(n850), .B(n851), .Z(n848) );
  NANDN U993 ( .A(B[370]), .B(n852), .Z(n851) );
  NANDN U994 ( .A(A[370]), .B(n853), .Z(n852) );
  NANDN U995 ( .A(n853), .B(A[370]), .Z(n850) );
  XOR U996 ( .A(n853), .B(n854), .Z(DIFF[370]) );
  XOR U997 ( .A(B[370]), .B(A[370]), .Z(n854) );
  AND U998 ( .A(n855), .B(n856), .Z(n853) );
  NANDN U999 ( .A(B[369]), .B(n857), .Z(n856) );
  NANDN U1000 ( .A(A[369]), .B(n858), .Z(n857) );
  NANDN U1001 ( .A(n858), .B(A[369]), .Z(n855) );
  XOR U1002 ( .A(n859), .B(n860), .Z(DIFF[36]) );
  XOR U1003 ( .A(B[36]), .B(A[36]), .Z(n860) );
  XOR U1004 ( .A(n858), .B(n861), .Z(DIFF[369]) );
  XOR U1005 ( .A(B[369]), .B(A[369]), .Z(n861) );
  AND U1006 ( .A(n862), .B(n863), .Z(n858) );
  NANDN U1007 ( .A(B[368]), .B(n864), .Z(n863) );
  NANDN U1008 ( .A(A[368]), .B(n865), .Z(n864) );
  NANDN U1009 ( .A(n865), .B(A[368]), .Z(n862) );
  XOR U1010 ( .A(n865), .B(n866), .Z(DIFF[368]) );
  XOR U1011 ( .A(B[368]), .B(A[368]), .Z(n866) );
  AND U1012 ( .A(n867), .B(n868), .Z(n865) );
  NANDN U1013 ( .A(B[367]), .B(n869), .Z(n868) );
  NANDN U1014 ( .A(A[367]), .B(n870), .Z(n869) );
  NANDN U1015 ( .A(n870), .B(A[367]), .Z(n867) );
  XOR U1016 ( .A(n870), .B(n871), .Z(DIFF[367]) );
  XOR U1017 ( .A(B[367]), .B(A[367]), .Z(n871) );
  AND U1018 ( .A(n872), .B(n873), .Z(n870) );
  NANDN U1019 ( .A(B[366]), .B(n874), .Z(n873) );
  NANDN U1020 ( .A(A[366]), .B(n875), .Z(n874) );
  NANDN U1021 ( .A(n875), .B(A[366]), .Z(n872) );
  XOR U1022 ( .A(n875), .B(n876), .Z(DIFF[366]) );
  XOR U1023 ( .A(B[366]), .B(A[366]), .Z(n876) );
  AND U1024 ( .A(n877), .B(n878), .Z(n875) );
  NANDN U1025 ( .A(B[365]), .B(n879), .Z(n878) );
  NANDN U1026 ( .A(A[365]), .B(n880), .Z(n879) );
  NANDN U1027 ( .A(n880), .B(A[365]), .Z(n877) );
  XOR U1028 ( .A(n880), .B(n881), .Z(DIFF[365]) );
  XOR U1029 ( .A(B[365]), .B(A[365]), .Z(n881) );
  AND U1030 ( .A(n882), .B(n883), .Z(n880) );
  NANDN U1031 ( .A(B[364]), .B(n884), .Z(n883) );
  NANDN U1032 ( .A(A[364]), .B(n885), .Z(n884) );
  NANDN U1033 ( .A(n885), .B(A[364]), .Z(n882) );
  XOR U1034 ( .A(n885), .B(n886), .Z(DIFF[364]) );
  XOR U1035 ( .A(B[364]), .B(A[364]), .Z(n886) );
  AND U1036 ( .A(n887), .B(n888), .Z(n885) );
  NANDN U1037 ( .A(B[363]), .B(n889), .Z(n888) );
  NANDN U1038 ( .A(A[363]), .B(n890), .Z(n889) );
  NANDN U1039 ( .A(n890), .B(A[363]), .Z(n887) );
  XOR U1040 ( .A(n890), .B(n891), .Z(DIFF[363]) );
  XOR U1041 ( .A(B[363]), .B(A[363]), .Z(n891) );
  AND U1042 ( .A(n892), .B(n893), .Z(n890) );
  NANDN U1043 ( .A(B[362]), .B(n894), .Z(n893) );
  NANDN U1044 ( .A(A[362]), .B(n895), .Z(n894) );
  NANDN U1045 ( .A(n895), .B(A[362]), .Z(n892) );
  XOR U1046 ( .A(n895), .B(n896), .Z(DIFF[362]) );
  XOR U1047 ( .A(B[362]), .B(A[362]), .Z(n896) );
  AND U1048 ( .A(n897), .B(n898), .Z(n895) );
  NANDN U1049 ( .A(B[361]), .B(n899), .Z(n898) );
  NANDN U1050 ( .A(A[361]), .B(n900), .Z(n899) );
  NANDN U1051 ( .A(n900), .B(A[361]), .Z(n897) );
  XOR U1052 ( .A(n900), .B(n901), .Z(DIFF[361]) );
  XOR U1053 ( .A(B[361]), .B(A[361]), .Z(n901) );
  AND U1054 ( .A(n902), .B(n903), .Z(n900) );
  NANDN U1055 ( .A(B[360]), .B(n904), .Z(n903) );
  NANDN U1056 ( .A(A[360]), .B(n905), .Z(n904) );
  NANDN U1057 ( .A(n905), .B(A[360]), .Z(n902) );
  XOR U1058 ( .A(n905), .B(n906), .Z(DIFF[360]) );
  XOR U1059 ( .A(B[360]), .B(A[360]), .Z(n906) );
  AND U1060 ( .A(n907), .B(n908), .Z(n905) );
  NANDN U1061 ( .A(B[359]), .B(n909), .Z(n908) );
  NANDN U1062 ( .A(A[359]), .B(n910), .Z(n909) );
  NANDN U1063 ( .A(n910), .B(A[359]), .Z(n907) );
  XOR U1064 ( .A(n911), .B(n912), .Z(DIFF[35]) );
  XOR U1065 ( .A(B[35]), .B(A[35]), .Z(n912) );
  XOR U1066 ( .A(n910), .B(n913), .Z(DIFF[359]) );
  XOR U1067 ( .A(B[359]), .B(A[359]), .Z(n913) );
  AND U1068 ( .A(n914), .B(n915), .Z(n910) );
  NANDN U1069 ( .A(B[358]), .B(n916), .Z(n915) );
  NANDN U1070 ( .A(A[358]), .B(n917), .Z(n916) );
  NANDN U1071 ( .A(n917), .B(A[358]), .Z(n914) );
  XOR U1072 ( .A(n917), .B(n918), .Z(DIFF[358]) );
  XOR U1073 ( .A(B[358]), .B(A[358]), .Z(n918) );
  AND U1074 ( .A(n919), .B(n920), .Z(n917) );
  NANDN U1075 ( .A(B[357]), .B(n921), .Z(n920) );
  NANDN U1076 ( .A(A[357]), .B(n922), .Z(n921) );
  NANDN U1077 ( .A(n922), .B(A[357]), .Z(n919) );
  XOR U1078 ( .A(n922), .B(n923), .Z(DIFF[357]) );
  XOR U1079 ( .A(B[357]), .B(A[357]), .Z(n923) );
  AND U1080 ( .A(n924), .B(n925), .Z(n922) );
  NANDN U1081 ( .A(B[356]), .B(n926), .Z(n925) );
  NANDN U1082 ( .A(A[356]), .B(n927), .Z(n926) );
  NANDN U1083 ( .A(n927), .B(A[356]), .Z(n924) );
  XOR U1084 ( .A(n927), .B(n928), .Z(DIFF[356]) );
  XOR U1085 ( .A(B[356]), .B(A[356]), .Z(n928) );
  AND U1086 ( .A(n929), .B(n930), .Z(n927) );
  NANDN U1087 ( .A(B[355]), .B(n931), .Z(n930) );
  NANDN U1088 ( .A(A[355]), .B(n932), .Z(n931) );
  NANDN U1089 ( .A(n932), .B(A[355]), .Z(n929) );
  XOR U1090 ( .A(n932), .B(n933), .Z(DIFF[355]) );
  XOR U1091 ( .A(B[355]), .B(A[355]), .Z(n933) );
  AND U1092 ( .A(n934), .B(n935), .Z(n932) );
  NANDN U1093 ( .A(B[354]), .B(n936), .Z(n935) );
  NANDN U1094 ( .A(A[354]), .B(n937), .Z(n936) );
  NANDN U1095 ( .A(n937), .B(A[354]), .Z(n934) );
  XOR U1096 ( .A(n937), .B(n938), .Z(DIFF[354]) );
  XOR U1097 ( .A(B[354]), .B(A[354]), .Z(n938) );
  AND U1098 ( .A(n939), .B(n940), .Z(n937) );
  NANDN U1099 ( .A(B[353]), .B(n941), .Z(n940) );
  NANDN U1100 ( .A(A[353]), .B(n942), .Z(n941) );
  NANDN U1101 ( .A(n942), .B(A[353]), .Z(n939) );
  XOR U1102 ( .A(n942), .B(n943), .Z(DIFF[353]) );
  XOR U1103 ( .A(B[353]), .B(A[353]), .Z(n943) );
  AND U1104 ( .A(n944), .B(n945), .Z(n942) );
  NANDN U1105 ( .A(B[352]), .B(n946), .Z(n945) );
  NANDN U1106 ( .A(A[352]), .B(n947), .Z(n946) );
  NANDN U1107 ( .A(n947), .B(A[352]), .Z(n944) );
  XOR U1108 ( .A(n947), .B(n948), .Z(DIFF[352]) );
  XOR U1109 ( .A(B[352]), .B(A[352]), .Z(n948) );
  AND U1110 ( .A(n949), .B(n950), .Z(n947) );
  NANDN U1111 ( .A(B[351]), .B(n951), .Z(n950) );
  NANDN U1112 ( .A(A[351]), .B(n952), .Z(n951) );
  NANDN U1113 ( .A(n952), .B(A[351]), .Z(n949) );
  XOR U1114 ( .A(n952), .B(n953), .Z(DIFF[351]) );
  XOR U1115 ( .A(B[351]), .B(A[351]), .Z(n953) );
  AND U1116 ( .A(n954), .B(n955), .Z(n952) );
  NANDN U1117 ( .A(B[350]), .B(n956), .Z(n955) );
  NANDN U1118 ( .A(A[350]), .B(n957), .Z(n956) );
  NANDN U1119 ( .A(n957), .B(A[350]), .Z(n954) );
  XOR U1120 ( .A(n957), .B(n958), .Z(DIFF[350]) );
  XOR U1121 ( .A(B[350]), .B(A[350]), .Z(n958) );
  AND U1122 ( .A(n959), .B(n960), .Z(n957) );
  NANDN U1123 ( .A(B[349]), .B(n961), .Z(n960) );
  NANDN U1124 ( .A(A[349]), .B(n962), .Z(n961) );
  NANDN U1125 ( .A(n962), .B(A[349]), .Z(n959) );
  XOR U1126 ( .A(n963), .B(n964), .Z(DIFF[34]) );
  XOR U1127 ( .A(B[34]), .B(A[34]), .Z(n964) );
  XOR U1128 ( .A(n962), .B(n965), .Z(DIFF[349]) );
  XOR U1129 ( .A(B[349]), .B(A[349]), .Z(n965) );
  AND U1130 ( .A(n966), .B(n967), .Z(n962) );
  NANDN U1131 ( .A(B[348]), .B(n968), .Z(n967) );
  NANDN U1132 ( .A(A[348]), .B(n969), .Z(n968) );
  NANDN U1133 ( .A(n969), .B(A[348]), .Z(n966) );
  XOR U1134 ( .A(n969), .B(n970), .Z(DIFF[348]) );
  XOR U1135 ( .A(B[348]), .B(A[348]), .Z(n970) );
  AND U1136 ( .A(n971), .B(n972), .Z(n969) );
  NANDN U1137 ( .A(B[347]), .B(n973), .Z(n972) );
  NANDN U1138 ( .A(A[347]), .B(n974), .Z(n973) );
  NANDN U1139 ( .A(n974), .B(A[347]), .Z(n971) );
  XOR U1140 ( .A(n974), .B(n975), .Z(DIFF[347]) );
  XOR U1141 ( .A(B[347]), .B(A[347]), .Z(n975) );
  AND U1142 ( .A(n976), .B(n977), .Z(n974) );
  NANDN U1143 ( .A(B[346]), .B(n978), .Z(n977) );
  NANDN U1144 ( .A(A[346]), .B(n979), .Z(n978) );
  NANDN U1145 ( .A(n979), .B(A[346]), .Z(n976) );
  XOR U1146 ( .A(n979), .B(n980), .Z(DIFF[346]) );
  XOR U1147 ( .A(B[346]), .B(A[346]), .Z(n980) );
  AND U1148 ( .A(n981), .B(n982), .Z(n979) );
  NANDN U1149 ( .A(B[345]), .B(n983), .Z(n982) );
  NANDN U1150 ( .A(A[345]), .B(n984), .Z(n983) );
  NANDN U1151 ( .A(n984), .B(A[345]), .Z(n981) );
  XOR U1152 ( .A(n984), .B(n985), .Z(DIFF[345]) );
  XOR U1153 ( .A(B[345]), .B(A[345]), .Z(n985) );
  AND U1154 ( .A(n986), .B(n987), .Z(n984) );
  NANDN U1155 ( .A(B[344]), .B(n988), .Z(n987) );
  NANDN U1156 ( .A(A[344]), .B(n989), .Z(n988) );
  NANDN U1157 ( .A(n989), .B(A[344]), .Z(n986) );
  XOR U1158 ( .A(n989), .B(n990), .Z(DIFF[344]) );
  XOR U1159 ( .A(B[344]), .B(A[344]), .Z(n990) );
  AND U1160 ( .A(n991), .B(n992), .Z(n989) );
  NANDN U1161 ( .A(B[343]), .B(n993), .Z(n992) );
  NANDN U1162 ( .A(A[343]), .B(n994), .Z(n993) );
  NANDN U1163 ( .A(n994), .B(A[343]), .Z(n991) );
  XOR U1164 ( .A(n994), .B(n995), .Z(DIFF[343]) );
  XOR U1165 ( .A(B[343]), .B(A[343]), .Z(n995) );
  AND U1166 ( .A(n996), .B(n997), .Z(n994) );
  NANDN U1167 ( .A(B[342]), .B(n998), .Z(n997) );
  NANDN U1168 ( .A(A[342]), .B(n999), .Z(n998) );
  NANDN U1169 ( .A(n999), .B(A[342]), .Z(n996) );
  XOR U1170 ( .A(n999), .B(n1000), .Z(DIFF[342]) );
  XOR U1171 ( .A(B[342]), .B(A[342]), .Z(n1000) );
  AND U1172 ( .A(n1001), .B(n1002), .Z(n999) );
  NANDN U1173 ( .A(B[341]), .B(n1003), .Z(n1002) );
  NANDN U1174 ( .A(A[341]), .B(n1004), .Z(n1003) );
  NANDN U1175 ( .A(n1004), .B(A[341]), .Z(n1001) );
  XOR U1176 ( .A(n1004), .B(n1005), .Z(DIFF[341]) );
  XOR U1177 ( .A(B[341]), .B(A[341]), .Z(n1005) );
  AND U1178 ( .A(n1006), .B(n1007), .Z(n1004) );
  NANDN U1179 ( .A(B[340]), .B(n1008), .Z(n1007) );
  NANDN U1180 ( .A(A[340]), .B(n1009), .Z(n1008) );
  NANDN U1181 ( .A(n1009), .B(A[340]), .Z(n1006) );
  XOR U1182 ( .A(n1009), .B(n1010), .Z(DIFF[340]) );
  XOR U1183 ( .A(B[340]), .B(A[340]), .Z(n1010) );
  AND U1184 ( .A(n1011), .B(n1012), .Z(n1009) );
  NANDN U1185 ( .A(B[339]), .B(n1013), .Z(n1012) );
  NANDN U1186 ( .A(A[339]), .B(n1014), .Z(n1013) );
  NANDN U1187 ( .A(n1014), .B(A[339]), .Z(n1011) );
  XOR U1188 ( .A(n1015), .B(n1016), .Z(DIFF[33]) );
  XOR U1189 ( .A(B[33]), .B(A[33]), .Z(n1016) );
  XOR U1190 ( .A(n1014), .B(n1017), .Z(DIFF[339]) );
  XOR U1191 ( .A(B[339]), .B(A[339]), .Z(n1017) );
  AND U1192 ( .A(n1018), .B(n1019), .Z(n1014) );
  NANDN U1193 ( .A(B[338]), .B(n1020), .Z(n1019) );
  NANDN U1194 ( .A(A[338]), .B(n1021), .Z(n1020) );
  NANDN U1195 ( .A(n1021), .B(A[338]), .Z(n1018) );
  XOR U1196 ( .A(n1021), .B(n1022), .Z(DIFF[338]) );
  XOR U1197 ( .A(B[338]), .B(A[338]), .Z(n1022) );
  AND U1198 ( .A(n1023), .B(n1024), .Z(n1021) );
  NANDN U1199 ( .A(B[337]), .B(n1025), .Z(n1024) );
  NANDN U1200 ( .A(A[337]), .B(n1026), .Z(n1025) );
  NANDN U1201 ( .A(n1026), .B(A[337]), .Z(n1023) );
  XOR U1202 ( .A(n1026), .B(n1027), .Z(DIFF[337]) );
  XOR U1203 ( .A(B[337]), .B(A[337]), .Z(n1027) );
  AND U1204 ( .A(n1028), .B(n1029), .Z(n1026) );
  NANDN U1205 ( .A(B[336]), .B(n1030), .Z(n1029) );
  NANDN U1206 ( .A(A[336]), .B(n1031), .Z(n1030) );
  NANDN U1207 ( .A(n1031), .B(A[336]), .Z(n1028) );
  XOR U1208 ( .A(n1031), .B(n1032), .Z(DIFF[336]) );
  XOR U1209 ( .A(B[336]), .B(A[336]), .Z(n1032) );
  AND U1210 ( .A(n1033), .B(n1034), .Z(n1031) );
  NANDN U1211 ( .A(B[335]), .B(n1035), .Z(n1034) );
  NANDN U1212 ( .A(A[335]), .B(n1036), .Z(n1035) );
  NANDN U1213 ( .A(n1036), .B(A[335]), .Z(n1033) );
  XOR U1214 ( .A(n1036), .B(n1037), .Z(DIFF[335]) );
  XOR U1215 ( .A(B[335]), .B(A[335]), .Z(n1037) );
  AND U1216 ( .A(n1038), .B(n1039), .Z(n1036) );
  NANDN U1217 ( .A(B[334]), .B(n1040), .Z(n1039) );
  NANDN U1218 ( .A(A[334]), .B(n1041), .Z(n1040) );
  NANDN U1219 ( .A(n1041), .B(A[334]), .Z(n1038) );
  XOR U1220 ( .A(n1041), .B(n1042), .Z(DIFF[334]) );
  XOR U1221 ( .A(B[334]), .B(A[334]), .Z(n1042) );
  AND U1222 ( .A(n1043), .B(n1044), .Z(n1041) );
  NANDN U1223 ( .A(B[333]), .B(n1045), .Z(n1044) );
  NANDN U1224 ( .A(A[333]), .B(n1046), .Z(n1045) );
  NANDN U1225 ( .A(n1046), .B(A[333]), .Z(n1043) );
  XOR U1226 ( .A(n1046), .B(n1047), .Z(DIFF[333]) );
  XOR U1227 ( .A(B[333]), .B(A[333]), .Z(n1047) );
  AND U1228 ( .A(n1048), .B(n1049), .Z(n1046) );
  NANDN U1229 ( .A(B[332]), .B(n1050), .Z(n1049) );
  NANDN U1230 ( .A(A[332]), .B(n1051), .Z(n1050) );
  NANDN U1231 ( .A(n1051), .B(A[332]), .Z(n1048) );
  XOR U1232 ( .A(n1051), .B(n1052), .Z(DIFF[332]) );
  XOR U1233 ( .A(B[332]), .B(A[332]), .Z(n1052) );
  AND U1234 ( .A(n1053), .B(n1054), .Z(n1051) );
  NANDN U1235 ( .A(B[331]), .B(n1055), .Z(n1054) );
  NANDN U1236 ( .A(A[331]), .B(n1056), .Z(n1055) );
  NANDN U1237 ( .A(n1056), .B(A[331]), .Z(n1053) );
  XOR U1238 ( .A(n1056), .B(n1057), .Z(DIFF[331]) );
  XOR U1239 ( .A(B[331]), .B(A[331]), .Z(n1057) );
  AND U1240 ( .A(n1058), .B(n1059), .Z(n1056) );
  NANDN U1241 ( .A(B[330]), .B(n1060), .Z(n1059) );
  NANDN U1242 ( .A(A[330]), .B(n1061), .Z(n1060) );
  NANDN U1243 ( .A(n1061), .B(A[330]), .Z(n1058) );
  XOR U1244 ( .A(n1061), .B(n1062), .Z(DIFF[330]) );
  XOR U1245 ( .A(B[330]), .B(A[330]), .Z(n1062) );
  AND U1246 ( .A(n1063), .B(n1064), .Z(n1061) );
  NANDN U1247 ( .A(B[329]), .B(n1065), .Z(n1064) );
  NANDN U1248 ( .A(A[329]), .B(n1066), .Z(n1065) );
  NANDN U1249 ( .A(n1066), .B(A[329]), .Z(n1063) );
  XOR U1250 ( .A(n1067), .B(n1068), .Z(DIFF[32]) );
  XOR U1251 ( .A(B[32]), .B(A[32]), .Z(n1068) );
  XOR U1252 ( .A(n1066), .B(n1069), .Z(DIFF[329]) );
  XOR U1253 ( .A(B[329]), .B(A[329]), .Z(n1069) );
  AND U1254 ( .A(n1070), .B(n1071), .Z(n1066) );
  NANDN U1255 ( .A(B[328]), .B(n1072), .Z(n1071) );
  NANDN U1256 ( .A(A[328]), .B(n1073), .Z(n1072) );
  NANDN U1257 ( .A(n1073), .B(A[328]), .Z(n1070) );
  XOR U1258 ( .A(n1073), .B(n1074), .Z(DIFF[328]) );
  XOR U1259 ( .A(B[328]), .B(A[328]), .Z(n1074) );
  AND U1260 ( .A(n1075), .B(n1076), .Z(n1073) );
  NANDN U1261 ( .A(B[327]), .B(n1077), .Z(n1076) );
  NANDN U1262 ( .A(A[327]), .B(n1078), .Z(n1077) );
  NANDN U1263 ( .A(n1078), .B(A[327]), .Z(n1075) );
  XOR U1264 ( .A(n1078), .B(n1079), .Z(DIFF[327]) );
  XOR U1265 ( .A(B[327]), .B(A[327]), .Z(n1079) );
  AND U1266 ( .A(n1080), .B(n1081), .Z(n1078) );
  NANDN U1267 ( .A(B[326]), .B(n1082), .Z(n1081) );
  NANDN U1268 ( .A(A[326]), .B(n1083), .Z(n1082) );
  NANDN U1269 ( .A(n1083), .B(A[326]), .Z(n1080) );
  XOR U1270 ( .A(n1083), .B(n1084), .Z(DIFF[326]) );
  XOR U1271 ( .A(B[326]), .B(A[326]), .Z(n1084) );
  AND U1272 ( .A(n1085), .B(n1086), .Z(n1083) );
  NANDN U1273 ( .A(B[325]), .B(n1087), .Z(n1086) );
  NANDN U1274 ( .A(A[325]), .B(n1088), .Z(n1087) );
  NANDN U1275 ( .A(n1088), .B(A[325]), .Z(n1085) );
  XOR U1276 ( .A(n1088), .B(n1089), .Z(DIFF[325]) );
  XOR U1277 ( .A(B[325]), .B(A[325]), .Z(n1089) );
  AND U1278 ( .A(n1090), .B(n1091), .Z(n1088) );
  NANDN U1279 ( .A(B[324]), .B(n1092), .Z(n1091) );
  NANDN U1280 ( .A(A[324]), .B(n1093), .Z(n1092) );
  NANDN U1281 ( .A(n1093), .B(A[324]), .Z(n1090) );
  XOR U1282 ( .A(n1093), .B(n1094), .Z(DIFF[324]) );
  XOR U1283 ( .A(B[324]), .B(A[324]), .Z(n1094) );
  AND U1284 ( .A(n1095), .B(n1096), .Z(n1093) );
  NANDN U1285 ( .A(B[323]), .B(n1097), .Z(n1096) );
  NANDN U1286 ( .A(A[323]), .B(n1098), .Z(n1097) );
  NANDN U1287 ( .A(n1098), .B(A[323]), .Z(n1095) );
  XOR U1288 ( .A(n1098), .B(n1099), .Z(DIFF[323]) );
  XOR U1289 ( .A(B[323]), .B(A[323]), .Z(n1099) );
  AND U1290 ( .A(n1100), .B(n1101), .Z(n1098) );
  NANDN U1291 ( .A(B[322]), .B(n1102), .Z(n1101) );
  NANDN U1292 ( .A(A[322]), .B(n1103), .Z(n1102) );
  NANDN U1293 ( .A(n1103), .B(A[322]), .Z(n1100) );
  XOR U1294 ( .A(n1103), .B(n1104), .Z(DIFF[322]) );
  XOR U1295 ( .A(B[322]), .B(A[322]), .Z(n1104) );
  AND U1296 ( .A(n1105), .B(n1106), .Z(n1103) );
  NANDN U1297 ( .A(B[321]), .B(n1107), .Z(n1106) );
  NANDN U1298 ( .A(A[321]), .B(n1108), .Z(n1107) );
  NANDN U1299 ( .A(n1108), .B(A[321]), .Z(n1105) );
  XOR U1300 ( .A(n1108), .B(n1109), .Z(DIFF[321]) );
  XOR U1301 ( .A(B[321]), .B(A[321]), .Z(n1109) );
  AND U1302 ( .A(n1110), .B(n1111), .Z(n1108) );
  NANDN U1303 ( .A(B[320]), .B(n1112), .Z(n1111) );
  NANDN U1304 ( .A(A[320]), .B(n1113), .Z(n1112) );
  NANDN U1305 ( .A(n1113), .B(A[320]), .Z(n1110) );
  XOR U1306 ( .A(n1113), .B(n1114), .Z(DIFF[320]) );
  XOR U1307 ( .A(B[320]), .B(A[320]), .Z(n1114) );
  AND U1308 ( .A(n1115), .B(n1116), .Z(n1113) );
  NANDN U1309 ( .A(B[319]), .B(n1117), .Z(n1116) );
  NANDN U1310 ( .A(A[319]), .B(n1118), .Z(n1117) );
  NANDN U1311 ( .A(n1118), .B(A[319]), .Z(n1115) );
  XOR U1312 ( .A(n1119), .B(n1120), .Z(DIFF[31]) );
  XOR U1313 ( .A(B[31]), .B(A[31]), .Z(n1120) );
  XOR U1314 ( .A(n1118), .B(n1121), .Z(DIFF[319]) );
  XOR U1315 ( .A(B[319]), .B(A[319]), .Z(n1121) );
  AND U1316 ( .A(n1122), .B(n1123), .Z(n1118) );
  NANDN U1317 ( .A(B[318]), .B(n1124), .Z(n1123) );
  NANDN U1318 ( .A(A[318]), .B(n1125), .Z(n1124) );
  NANDN U1319 ( .A(n1125), .B(A[318]), .Z(n1122) );
  XOR U1320 ( .A(n1125), .B(n1126), .Z(DIFF[318]) );
  XOR U1321 ( .A(B[318]), .B(A[318]), .Z(n1126) );
  AND U1322 ( .A(n1127), .B(n1128), .Z(n1125) );
  NANDN U1323 ( .A(B[317]), .B(n1129), .Z(n1128) );
  NANDN U1324 ( .A(A[317]), .B(n1130), .Z(n1129) );
  NANDN U1325 ( .A(n1130), .B(A[317]), .Z(n1127) );
  XOR U1326 ( .A(n1130), .B(n1131), .Z(DIFF[317]) );
  XOR U1327 ( .A(B[317]), .B(A[317]), .Z(n1131) );
  AND U1328 ( .A(n1132), .B(n1133), .Z(n1130) );
  NANDN U1329 ( .A(B[316]), .B(n1134), .Z(n1133) );
  NANDN U1330 ( .A(A[316]), .B(n1135), .Z(n1134) );
  NANDN U1331 ( .A(n1135), .B(A[316]), .Z(n1132) );
  XOR U1332 ( .A(n1135), .B(n1136), .Z(DIFF[316]) );
  XOR U1333 ( .A(B[316]), .B(A[316]), .Z(n1136) );
  AND U1334 ( .A(n1137), .B(n1138), .Z(n1135) );
  NANDN U1335 ( .A(B[315]), .B(n1139), .Z(n1138) );
  NANDN U1336 ( .A(A[315]), .B(n1140), .Z(n1139) );
  NANDN U1337 ( .A(n1140), .B(A[315]), .Z(n1137) );
  XOR U1338 ( .A(n1140), .B(n1141), .Z(DIFF[315]) );
  XOR U1339 ( .A(B[315]), .B(A[315]), .Z(n1141) );
  AND U1340 ( .A(n1142), .B(n1143), .Z(n1140) );
  NANDN U1341 ( .A(B[314]), .B(n1144), .Z(n1143) );
  NANDN U1342 ( .A(A[314]), .B(n1145), .Z(n1144) );
  NANDN U1343 ( .A(n1145), .B(A[314]), .Z(n1142) );
  XOR U1344 ( .A(n1145), .B(n1146), .Z(DIFF[314]) );
  XOR U1345 ( .A(B[314]), .B(A[314]), .Z(n1146) );
  AND U1346 ( .A(n1147), .B(n1148), .Z(n1145) );
  NANDN U1347 ( .A(B[313]), .B(n1149), .Z(n1148) );
  NANDN U1348 ( .A(A[313]), .B(n1150), .Z(n1149) );
  NANDN U1349 ( .A(n1150), .B(A[313]), .Z(n1147) );
  XOR U1350 ( .A(n1150), .B(n1151), .Z(DIFF[313]) );
  XOR U1351 ( .A(B[313]), .B(A[313]), .Z(n1151) );
  AND U1352 ( .A(n1152), .B(n1153), .Z(n1150) );
  NANDN U1353 ( .A(B[312]), .B(n1154), .Z(n1153) );
  NANDN U1354 ( .A(A[312]), .B(n1155), .Z(n1154) );
  NANDN U1355 ( .A(n1155), .B(A[312]), .Z(n1152) );
  XOR U1356 ( .A(n1155), .B(n1156), .Z(DIFF[312]) );
  XOR U1357 ( .A(B[312]), .B(A[312]), .Z(n1156) );
  AND U1358 ( .A(n1157), .B(n1158), .Z(n1155) );
  NANDN U1359 ( .A(B[311]), .B(n1159), .Z(n1158) );
  NANDN U1360 ( .A(A[311]), .B(n1160), .Z(n1159) );
  NANDN U1361 ( .A(n1160), .B(A[311]), .Z(n1157) );
  XOR U1362 ( .A(n1160), .B(n1161), .Z(DIFF[311]) );
  XOR U1363 ( .A(B[311]), .B(A[311]), .Z(n1161) );
  AND U1364 ( .A(n1162), .B(n1163), .Z(n1160) );
  NANDN U1365 ( .A(B[310]), .B(n1164), .Z(n1163) );
  NANDN U1366 ( .A(A[310]), .B(n1165), .Z(n1164) );
  NANDN U1367 ( .A(n1165), .B(A[310]), .Z(n1162) );
  XOR U1368 ( .A(n1165), .B(n1166), .Z(DIFF[310]) );
  XOR U1369 ( .A(B[310]), .B(A[310]), .Z(n1166) );
  AND U1370 ( .A(n1167), .B(n1168), .Z(n1165) );
  NANDN U1371 ( .A(B[309]), .B(n1169), .Z(n1168) );
  NANDN U1372 ( .A(A[309]), .B(n1170), .Z(n1169) );
  NANDN U1373 ( .A(n1170), .B(A[309]), .Z(n1167) );
  XOR U1374 ( .A(n1171), .B(n1172), .Z(DIFF[30]) );
  XOR U1375 ( .A(B[30]), .B(A[30]), .Z(n1172) );
  XOR U1376 ( .A(n1170), .B(n1173), .Z(DIFF[309]) );
  XOR U1377 ( .A(B[309]), .B(A[309]), .Z(n1173) );
  AND U1378 ( .A(n1174), .B(n1175), .Z(n1170) );
  NANDN U1379 ( .A(B[308]), .B(n1176), .Z(n1175) );
  NANDN U1380 ( .A(A[308]), .B(n1177), .Z(n1176) );
  NANDN U1381 ( .A(n1177), .B(A[308]), .Z(n1174) );
  XOR U1382 ( .A(n1177), .B(n1178), .Z(DIFF[308]) );
  XOR U1383 ( .A(B[308]), .B(A[308]), .Z(n1178) );
  AND U1384 ( .A(n1179), .B(n1180), .Z(n1177) );
  NANDN U1385 ( .A(B[307]), .B(n1181), .Z(n1180) );
  NANDN U1386 ( .A(A[307]), .B(n1182), .Z(n1181) );
  NANDN U1387 ( .A(n1182), .B(A[307]), .Z(n1179) );
  XOR U1388 ( .A(n1182), .B(n1183), .Z(DIFF[307]) );
  XOR U1389 ( .A(B[307]), .B(A[307]), .Z(n1183) );
  AND U1390 ( .A(n1184), .B(n1185), .Z(n1182) );
  NANDN U1391 ( .A(B[306]), .B(n1186), .Z(n1185) );
  NANDN U1392 ( .A(A[306]), .B(n1187), .Z(n1186) );
  NANDN U1393 ( .A(n1187), .B(A[306]), .Z(n1184) );
  XOR U1394 ( .A(n1187), .B(n1188), .Z(DIFF[306]) );
  XOR U1395 ( .A(B[306]), .B(A[306]), .Z(n1188) );
  AND U1396 ( .A(n1189), .B(n1190), .Z(n1187) );
  NANDN U1397 ( .A(B[305]), .B(n1191), .Z(n1190) );
  NANDN U1398 ( .A(A[305]), .B(n1192), .Z(n1191) );
  NANDN U1399 ( .A(n1192), .B(A[305]), .Z(n1189) );
  XOR U1400 ( .A(n1192), .B(n1193), .Z(DIFF[305]) );
  XOR U1401 ( .A(B[305]), .B(A[305]), .Z(n1193) );
  AND U1402 ( .A(n1194), .B(n1195), .Z(n1192) );
  NANDN U1403 ( .A(B[304]), .B(n1196), .Z(n1195) );
  NANDN U1404 ( .A(A[304]), .B(n1197), .Z(n1196) );
  NANDN U1405 ( .A(n1197), .B(A[304]), .Z(n1194) );
  XOR U1406 ( .A(n1197), .B(n1198), .Z(DIFF[304]) );
  XOR U1407 ( .A(B[304]), .B(A[304]), .Z(n1198) );
  AND U1408 ( .A(n1199), .B(n1200), .Z(n1197) );
  NANDN U1409 ( .A(B[303]), .B(n1201), .Z(n1200) );
  NANDN U1410 ( .A(A[303]), .B(n1202), .Z(n1201) );
  NANDN U1411 ( .A(n1202), .B(A[303]), .Z(n1199) );
  XOR U1412 ( .A(n1202), .B(n1203), .Z(DIFF[303]) );
  XOR U1413 ( .A(B[303]), .B(A[303]), .Z(n1203) );
  AND U1414 ( .A(n1204), .B(n1205), .Z(n1202) );
  NANDN U1415 ( .A(B[302]), .B(n1206), .Z(n1205) );
  NANDN U1416 ( .A(A[302]), .B(n1207), .Z(n1206) );
  NANDN U1417 ( .A(n1207), .B(A[302]), .Z(n1204) );
  XOR U1418 ( .A(n1207), .B(n1208), .Z(DIFF[302]) );
  XOR U1419 ( .A(B[302]), .B(A[302]), .Z(n1208) );
  AND U1420 ( .A(n1209), .B(n1210), .Z(n1207) );
  NANDN U1421 ( .A(B[301]), .B(n1211), .Z(n1210) );
  NANDN U1422 ( .A(A[301]), .B(n1212), .Z(n1211) );
  NANDN U1423 ( .A(n1212), .B(A[301]), .Z(n1209) );
  XOR U1424 ( .A(n1212), .B(n1213), .Z(DIFF[301]) );
  XOR U1425 ( .A(B[301]), .B(A[301]), .Z(n1213) );
  AND U1426 ( .A(n1214), .B(n1215), .Z(n1212) );
  NANDN U1427 ( .A(B[300]), .B(n1216), .Z(n1215) );
  NANDN U1428 ( .A(A[300]), .B(n1217), .Z(n1216) );
  NANDN U1429 ( .A(n1217), .B(A[300]), .Z(n1214) );
  XOR U1430 ( .A(n1217), .B(n1218), .Z(DIFF[300]) );
  XOR U1431 ( .A(B[300]), .B(A[300]), .Z(n1218) );
  AND U1432 ( .A(n1219), .B(n1220), .Z(n1217) );
  NANDN U1433 ( .A(B[299]), .B(n1221), .Z(n1220) );
  NANDN U1434 ( .A(A[299]), .B(n1222), .Z(n1221) );
  NANDN U1435 ( .A(n1222), .B(A[299]), .Z(n1219) );
  XOR U1436 ( .A(n1223), .B(n1224), .Z(DIFF[2]) );
  XOR U1437 ( .A(B[2]), .B(A[2]), .Z(n1224) );
  XOR U1438 ( .A(n1225), .B(n1226), .Z(DIFF[29]) );
  XOR U1439 ( .A(B[29]), .B(A[29]), .Z(n1226) );
  XOR U1440 ( .A(n1222), .B(n1227), .Z(DIFF[299]) );
  XOR U1441 ( .A(B[299]), .B(A[299]), .Z(n1227) );
  AND U1442 ( .A(n1228), .B(n1229), .Z(n1222) );
  NANDN U1443 ( .A(B[298]), .B(n1230), .Z(n1229) );
  NANDN U1444 ( .A(A[298]), .B(n1231), .Z(n1230) );
  NANDN U1445 ( .A(n1231), .B(A[298]), .Z(n1228) );
  XOR U1446 ( .A(n1231), .B(n1232), .Z(DIFF[298]) );
  XOR U1447 ( .A(B[298]), .B(A[298]), .Z(n1232) );
  AND U1448 ( .A(n1233), .B(n1234), .Z(n1231) );
  NANDN U1449 ( .A(B[297]), .B(n1235), .Z(n1234) );
  NANDN U1450 ( .A(A[297]), .B(n1236), .Z(n1235) );
  NANDN U1451 ( .A(n1236), .B(A[297]), .Z(n1233) );
  XOR U1452 ( .A(n1236), .B(n1237), .Z(DIFF[297]) );
  XOR U1453 ( .A(B[297]), .B(A[297]), .Z(n1237) );
  AND U1454 ( .A(n1238), .B(n1239), .Z(n1236) );
  NANDN U1455 ( .A(B[296]), .B(n1240), .Z(n1239) );
  NANDN U1456 ( .A(A[296]), .B(n1241), .Z(n1240) );
  NANDN U1457 ( .A(n1241), .B(A[296]), .Z(n1238) );
  XOR U1458 ( .A(n1241), .B(n1242), .Z(DIFF[296]) );
  XOR U1459 ( .A(B[296]), .B(A[296]), .Z(n1242) );
  AND U1460 ( .A(n1243), .B(n1244), .Z(n1241) );
  NANDN U1461 ( .A(B[295]), .B(n1245), .Z(n1244) );
  NANDN U1462 ( .A(A[295]), .B(n1246), .Z(n1245) );
  NANDN U1463 ( .A(n1246), .B(A[295]), .Z(n1243) );
  XOR U1464 ( .A(n1246), .B(n1247), .Z(DIFF[295]) );
  XOR U1465 ( .A(B[295]), .B(A[295]), .Z(n1247) );
  AND U1466 ( .A(n1248), .B(n1249), .Z(n1246) );
  NANDN U1467 ( .A(B[294]), .B(n1250), .Z(n1249) );
  NANDN U1468 ( .A(A[294]), .B(n1251), .Z(n1250) );
  NANDN U1469 ( .A(n1251), .B(A[294]), .Z(n1248) );
  XOR U1470 ( .A(n1251), .B(n1252), .Z(DIFF[294]) );
  XOR U1471 ( .A(B[294]), .B(A[294]), .Z(n1252) );
  AND U1472 ( .A(n1253), .B(n1254), .Z(n1251) );
  NANDN U1473 ( .A(B[293]), .B(n1255), .Z(n1254) );
  NANDN U1474 ( .A(A[293]), .B(n1256), .Z(n1255) );
  NANDN U1475 ( .A(n1256), .B(A[293]), .Z(n1253) );
  XOR U1476 ( .A(n1256), .B(n1257), .Z(DIFF[293]) );
  XOR U1477 ( .A(B[293]), .B(A[293]), .Z(n1257) );
  AND U1478 ( .A(n1258), .B(n1259), .Z(n1256) );
  NANDN U1479 ( .A(B[292]), .B(n1260), .Z(n1259) );
  NANDN U1480 ( .A(A[292]), .B(n1261), .Z(n1260) );
  NANDN U1481 ( .A(n1261), .B(A[292]), .Z(n1258) );
  XOR U1482 ( .A(n1261), .B(n1262), .Z(DIFF[292]) );
  XOR U1483 ( .A(B[292]), .B(A[292]), .Z(n1262) );
  AND U1484 ( .A(n1263), .B(n1264), .Z(n1261) );
  NANDN U1485 ( .A(B[291]), .B(n1265), .Z(n1264) );
  NANDN U1486 ( .A(A[291]), .B(n1266), .Z(n1265) );
  NANDN U1487 ( .A(n1266), .B(A[291]), .Z(n1263) );
  XOR U1488 ( .A(n1266), .B(n1267), .Z(DIFF[291]) );
  XOR U1489 ( .A(B[291]), .B(A[291]), .Z(n1267) );
  AND U1490 ( .A(n1268), .B(n1269), .Z(n1266) );
  NANDN U1491 ( .A(B[290]), .B(n1270), .Z(n1269) );
  NANDN U1492 ( .A(A[290]), .B(n1271), .Z(n1270) );
  NANDN U1493 ( .A(n1271), .B(A[290]), .Z(n1268) );
  XOR U1494 ( .A(n1271), .B(n1272), .Z(DIFF[290]) );
  XOR U1495 ( .A(B[290]), .B(A[290]), .Z(n1272) );
  AND U1496 ( .A(n1273), .B(n1274), .Z(n1271) );
  NANDN U1497 ( .A(B[289]), .B(n1275), .Z(n1274) );
  NANDN U1498 ( .A(A[289]), .B(n1276), .Z(n1275) );
  NANDN U1499 ( .A(n1276), .B(A[289]), .Z(n1273) );
  XOR U1500 ( .A(n1277), .B(n1278), .Z(DIFF[28]) );
  XOR U1501 ( .A(B[28]), .B(A[28]), .Z(n1278) );
  XOR U1502 ( .A(n1276), .B(n1279), .Z(DIFF[289]) );
  XOR U1503 ( .A(B[289]), .B(A[289]), .Z(n1279) );
  AND U1504 ( .A(n1280), .B(n1281), .Z(n1276) );
  NANDN U1505 ( .A(B[288]), .B(n1282), .Z(n1281) );
  NANDN U1506 ( .A(A[288]), .B(n1283), .Z(n1282) );
  NANDN U1507 ( .A(n1283), .B(A[288]), .Z(n1280) );
  XOR U1508 ( .A(n1283), .B(n1284), .Z(DIFF[288]) );
  XOR U1509 ( .A(B[288]), .B(A[288]), .Z(n1284) );
  AND U1510 ( .A(n1285), .B(n1286), .Z(n1283) );
  NANDN U1511 ( .A(B[287]), .B(n1287), .Z(n1286) );
  NANDN U1512 ( .A(A[287]), .B(n1288), .Z(n1287) );
  NANDN U1513 ( .A(n1288), .B(A[287]), .Z(n1285) );
  XOR U1514 ( .A(n1288), .B(n1289), .Z(DIFF[287]) );
  XOR U1515 ( .A(B[287]), .B(A[287]), .Z(n1289) );
  AND U1516 ( .A(n1290), .B(n1291), .Z(n1288) );
  NANDN U1517 ( .A(B[286]), .B(n1292), .Z(n1291) );
  NANDN U1518 ( .A(A[286]), .B(n1293), .Z(n1292) );
  NANDN U1519 ( .A(n1293), .B(A[286]), .Z(n1290) );
  XOR U1520 ( .A(n1293), .B(n1294), .Z(DIFF[286]) );
  XOR U1521 ( .A(B[286]), .B(A[286]), .Z(n1294) );
  AND U1522 ( .A(n1295), .B(n1296), .Z(n1293) );
  NANDN U1523 ( .A(B[285]), .B(n1297), .Z(n1296) );
  NANDN U1524 ( .A(A[285]), .B(n1298), .Z(n1297) );
  NANDN U1525 ( .A(n1298), .B(A[285]), .Z(n1295) );
  XOR U1526 ( .A(n1298), .B(n1299), .Z(DIFF[285]) );
  XOR U1527 ( .A(B[285]), .B(A[285]), .Z(n1299) );
  AND U1528 ( .A(n1300), .B(n1301), .Z(n1298) );
  NANDN U1529 ( .A(B[284]), .B(n1302), .Z(n1301) );
  NANDN U1530 ( .A(A[284]), .B(n1303), .Z(n1302) );
  NANDN U1531 ( .A(n1303), .B(A[284]), .Z(n1300) );
  XOR U1532 ( .A(n1303), .B(n1304), .Z(DIFF[284]) );
  XOR U1533 ( .A(B[284]), .B(A[284]), .Z(n1304) );
  AND U1534 ( .A(n1305), .B(n1306), .Z(n1303) );
  NANDN U1535 ( .A(B[283]), .B(n1307), .Z(n1306) );
  NANDN U1536 ( .A(A[283]), .B(n1308), .Z(n1307) );
  NANDN U1537 ( .A(n1308), .B(A[283]), .Z(n1305) );
  XOR U1538 ( .A(n1308), .B(n1309), .Z(DIFF[283]) );
  XOR U1539 ( .A(B[283]), .B(A[283]), .Z(n1309) );
  AND U1540 ( .A(n1310), .B(n1311), .Z(n1308) );
  NANDN U1541 ( .A(B[282]), .B(n1312), .Z(n1311) );
  NANDN U1542 ( .A(A[282]), .B(n1313), .Z(n1312) );
  NANDN U1543 ( .A(n1313), .B(A[282]), .Z(n1310) );
  XOR U1544 ( .A(n1313), .B(n1314), .Z(DIFF[282]) );
  XOR U1545 ( .A(B[282]), .B(A[282]), .Z(n1314) );
  AND U1546 ( .A(n1315), .B(n1316), .Z(n1313) );
  NANDN U1547 ( .A(B[281]), .B(n1317), .Z(n1316) );
  NANDN U1548 ( .A(A[281]), .B(n1318), .Z(n1317) );
  NANDN U1549 ( .A(n1318), .B(A[281]), .Z(n1315) );
  XOR U1550 ( .A(n1318), .B(n1319), .Z(DIFF[281]) );
  XOR U1551 ( .A(B[281]), .B(A[281]), .Z(n1319) );
  AND U1552 ( .A(n1320), .B(n1321), .Z(n1318) );
  NANDN U1553 ( .A(B[280]), .B(n1322), .Z(n1321) );
  NANDN U1554 ( .A(A[280]), .B(n1323), .Z(n1322) );
  NANDN U1555 ( .A(n1323), .B(A[280]), .Z(n1320) );
  XOR U1556 ( .A(n1323), .B(n1324), .Z(DIFF[280]) );
  XOR U1557 ( .A(B[280]), .B(A[280]), .Z(n1324) );
  AND U1558 ( .A(n1325), .B(n1326), .Z(n1323) );
  NANDN U1559 ( .A(B[279]), .B(n1327), .Z(n1326) );
  NANDN U1560 ( .A(A[279]), .B(n1328), .Z(n1327) );
  NANDN U1561 ( .A(n1328), .B(A[279]), .Z(n1325) );
  XOR U1562 ( .A(n1329), .B(n1330), .Z(DIFF[27]) );
  XOR U1563 ( .A(B[27]), .B(A[27]), .Z(n1330) );
  XOR U1564 ( .A(n1328), .B(n1331), .Z(DIFF[279]) );
  XOR U1565 ( .A(B[279]), .B(A[279]), .Z(n1331) );
  AND U1566 ( .A(n1332), .B(n1333), .Z(n1328) );
  NANDN U1567 ( .A(B[278]), .B(n1334), .Z(n1333) );
  NANDN U1568 ( .A(A[278]), .B(n1335), .Z(n1334) );
  NANDN U1569 ( .A(n1335), .B(A[278]), .Z(n1332) );
  XOR U1570 ( .A(n1335), .B(n1336), .Z(DIFF[278]) );
  XOR U1571 ( .A(B[278]), .B(A[278]), .Z(n1336) );
  AND U1572 ( .A(n1337), .B(n1338), .Z(n1335) );
  NANDN U1573 ( .A(B[277]), .B(n1339), .Z(n1338) );
  NANDN U1574 ( .A(A[277]), .B(n1340), .Z(n1339) );
  NANDN U1575 ( .A(n1340), .B(A[277]), .Z(n1337) );
  XOR U1576 ( .A(n1340), .B(n1341), .Z(DIFF[277]) );
  XOR U1577 ( .A(B[277]), .B(A[277]), .Z(n1341) );
  AND U1578 ( .A(n1342), .B(n1343), .Z(n1340) );
  NANDN U1579 ( .A(B[276]), .B(n1344), .Z(n1343) );
  NANDN U1580 ( .A(A[276]), .B(n1345), .Z(n1344) );
  NANDN U1581 ( .A(n1345), .B(A[276]), .Z(n1342) );
  XOR U1582 ( .A(n1345), .B(n1346), .Z(DIFF[276]) );
  XOR U1583 ( .A(B[276]), .B(A[276]), .Z(n1346) );
  AND U1584 ( .A(n1347), .B(n1348), .Z(n1345) );
  NANDN U1585 ( .A(B[275]), .B(n1349), .Z(n1348) );
  NANDN U1586 ( .A(A[275]), .B(n1350), .Z(n1349) );
  NANDN U1587 ( .A(n1350), .B(A[275]), .Z(n1347) );
  XOR U1588 ( .A(n1350), .B(n1351), .Z(DIFF[275]) );
  XOR U1589 ( .A(B[275]), .B(A[275]), .Z(n1351) );
  AND U1590 ( .A(n1352), .B(n1353), .Z(n1350) );
  NANDN U1591 ( .A(B[274]), .B(n1354), .Z(n1353) );
  NANDN U1592 ( .A(A[274]), .B(n1355), .Z(n1354) );
  NANDN U1593 ( .A(n1355), .B(A[274]), .Z(n1352) );
  XOR U1594 ( .A(n1355), .B(n1356), .Z(DIFF[274]) );
  XOR U1595 ( .A(B[274]), .B(A[274]), .Z(n1356) );
  AND U1596 ( .A(n1357), .B(n1358), .Z(n1355) );
  NANDN U1597 ( .A(B[273]), .B(n1359), .Z(n1358) );
  NANDN U1598 ( .A(A[273]), .B(n1360), .Z(n1359) );
  NANDN U1599 ( .A(n1360), .B(A[273]), .Z(n1357) );
  XOR U1600 ( .A(n1360), .B(n1361), .Z(DIFF[273]) );
  XOR U1601 ( .A(B[273]), .B(A[273]), .Z(n1361) );
  AND U1602 ( .A(n1362), .B(n1363), .Z(n1360) );
  NANDN U1603 ( .A(B[272]), .B(n1364), .Z(n1363) );
  NANDN U1604 ( .A(A[272]), .B(n1365), .Z(n1364) );
  NANDN U1605 ( .A(n1365), .B(A[272]), .Z(n1362) );
  XOR U1606 ( .A(n1365), .B(n1366), .Z(DIFF[272]) );
  XOR U1607 ( .A(B[272]), .B(A[272]), .Z(n1366) );
  AND U1608 ( .A(n1367), .B(n1368), .Z(n1365) );
  NANDN U1609 ( .A(B[271]), .B(n1369), .Z(n1368) );
  NANDN U1610 ( .A(A[271]), .B(n1370), .Z(n1369) );
  NANDN U1611 ( .A(n1370), .B(A[271]), .Z(n1367) );
  XOR U1612 ( .A(n1370), .B(n1371), .Z(DIFF[271]) );
  XOR U1613 ( .A(B[271]), .B(A[271]), .Z(n1371) );
  AND U1614 ( .A(n1372), .B(n1373), .Z(n1370) );
  NANDN U1615 ( .A(B[270]), .B(n1374), .Z(n1373) );
  NANDN U1616 ( .A(A[270]), .B(n1375), .Z(n1374) );
  NANDN U1617 ( .A(n1375), .B(A[270]), .Z(n1372) );
  XOR U1618 ( .A(n1375), .B(n1376), .Z(DIFF[270]) );
  XOR U1619 ( .A(B[270]), .B(A[270]), .Z(n1376) );
  AND U1620 ( .A(n1377), .B(n1378), .Z(n1375) );
  NANDN U1621 ( .A(B[269]), .B(n1379), .Z(n1378) );
  NANDN U1622 ( .A(A[269]), .B(n1380), .Z(n1379) );
  NANDN U1623 ( .A(n1380), .B(A[269]), .Z(n1377) );
  XOR U1624 ( .A(n1381), .B(n1382), .Z(DIFF[26]) );
  XOR U1625 ( .A(B[26]), .B(A[26]), .Z(n1382) );
  XOR U1626 ( .A(n1380), .B(n1383), .Z(DIFF[269]) );
  XOR U1627 ( .A(B[269]), .B(A[269]), .Z(n1383) );
  AND U1628 ( .A(n1384), .B(n1385), .Z(n1380) );
  NANDN U1629 ( .A(B[268]), .B(n1386), .Z(n1385) );
  NANDN U1630 ( .A(A[268]), .B(n1387), .Z(n1386) );
  NANDN U1631 ( .A(n1387), .B(A[268]), .Z(n1384) );
  XOR U1632 ( .A(n1387), .B(n1388), .Z(DIFF[268]) );
  XOR U1633 ( .A(B[268]), .B(A[268]), .Z(n1388) );
  AND U1634 ( .A(n1389), .B(n1390), .Z(n1387) );
  NANDN U1635 ( .A(B[267]), .B(n1391), .Z(n1390) );
  NANDN U1636 ( .A(A[267]), .B(n1392), .Z(n1391) );
  NANDN U1637 ( .A(n1392), .B(A[267]), .Z(n1389) );
  XOR U1638 ( .A(n1392), .B(n1393), .Z(DIFF[267]) );
  XOR U1639 ( .A(B[267]), .B(A[267]), .Z(n1393) );
  AND U1640 ( .A(n1394), .B(n1395), .Z(n1392) );
  NANDN U1641 ( .A(B[266]), .B(n1396), .Z(n1395) );
  NANDN U1642 ( .A(A[266]), .B(n1397), .Z(n1396) );
  NANDN U1643 ( .A(n1397), .B(A[266]), .Z(n1394) );
  XOR U1644 ( .A(n1397), .B(n1398), .Z(DIFF[266]) );
  XOR U1645 ( .A(B[266]), .B(A[266]), .Z(n1398) );
  AND U1646 ( .A(n1399), .B(n1400), .Z(n1397) );
  NANDN U1647 ( .A(B[265]), .B(n1401), .Z(n1400) );
  NANDN U1648 ( .A(A[265]), .B(n1402), .Z(n1401) );
  NANDN U1649 ( .A(n1402), .B(A[265]), .Z(n1399) );
  XOR U1650 ( .A(n1402), .B(n1403), .Z(DIFF[265]) );
  XOR U1651 ( .A(B[265]), .B(A[265]), .Z(n1403) );
  AND U1652 ( .A(n1404), .B(n1405), .Z(n1402) );
  NANDN U1653 ( .A(B[264]), .B(n1406), .Z(n1405) );
  NANDN U1654 ( .A(A[264]), .B(n1407), .Z(n1406) );
  NANDN U1655 ( .A(n1407), .B(A[264]), .Z(n1404) );
  XOR U1656 ( .A(n1407), .B(n1408), .Z(DIFF[264]) );
  XOR U1657 ( .A(B[264]), .B(A[264]), .Z(n1408) );
  AND U1658 ( .A(n1409), .B(n1410), .Z(n1407) );
  NANDN U1659 ( .A(B[263]), .B(n1411), .Z(n1410) );
  NANDN U1660 ( .A(A[263]), .B(n1412), .Z(n1411) );
  NANDN U1661 ( .A(n1412), .B(A[263]), .Z(n1409) );
  XOR U1662 ( .A(n1412), .B(n1413), .Z(DIFF[263]) );
  XOR U1663 ( .A(B[263]), .B(A[263]), .Z(n1413) );
  AND U1664 ( .A(n1414), .B(n1415), .Z(n1412) );
  NANDN U1665 ( .A(B[262]), .B(n1416), .Z(n1415) );
  NANDN U1666 ( .A(A[262]), .B(n1417), .Z(n1416) );
  NANDN U1667 ( .A(n1417), .B(A[262]), .Z(n1414) );
  XOR U1668 ( .A(n1417), .B(n1418), .Z(DIFF[262]) );
  XOR U1669 ( .A(B[262]), .B(A[262]), .Z(n1418) );
  AND U1670 ( .A(n1419), .B(n1420), .Z(n1417) );
  NANDN U1671 ( .A(B[261]), .B(n1421), .Z(n1420) );
  NANDN U1672 ( .A(A[261]), .B(n1422), .Z(n1421) );
  NANDN U1673 ( .A(n1422), .B(A[261]), .Z(n1419) );
  XOR U1674 ( .A(n1422), .B(n1423), .Z(DIFF[261]) );
  XOR U1675 ( .A(B[261]), .B(A[261]), .Z(n1423) );
  AND U1676 ( .A(n1424), .B(n1425), .Z(n1422) );
  NANDN U1677 ( .A(B[260]), .B(n1426), .Z(n1425) );
  NANDN U1678 ( .A(A[260]), .B(n1427), .Z(n1426) );
  NANDN U1679 ( .A(n1427), .B(A[260]), .Z(n1424) );
  XOR U1680 ( .A(n1427), .B(n1428), .Z(DIFF[260]) );
  XOR U1681 ( .A(B[260]), .B(A[260]), .Z(n1428) );
  AND U1682 ( .A(n1429), .B(n1430), .Z(n1427) );
  NANDN U1683 ( .A(B[259]), .B(n1431), .Z(n1430) );
  NANDN U1684 ( .A(A[259]), .B(n1432), .Z(n1431) );
  NANDN U1685 ( .A(n1432), .B(A[259]), .Z(n1429) );
  XOR U1686 ( .A(n1433), .B(n1434), .Z(DIFF[25]) );
  XOR U1687 ( .A(B[25]), .B(A[25]), .Z(n1434) );
  XOR U1688 ( .A(n1432), .B(n1435), .Z(DIFF[259]) );
  XOR U1689 ( .A(B[259]), .B(A[259]), .Z(n1435) );
  AND U1690 ( .A(n1436), .B(n1437), .Z(n1432) );
  NANDN U1691 ( .A(B[258]), .B(n1438), .Z(n1437) );
  NANDN U1692 ( .A(A[258]), .B(n1439), .Z(n1438) );
  NANDN U1693 ( .A(n1439), .B(A[258]), .Z(n1436) );
  XOR U1694 ( .A(n1439), .B(n1440), .Z(DIFF[258]) );
  XOR U1695 ( .A(B[258]), .B(A[258]), .Z(n1440) );
  AND U1696 ( .A(n1441), .B(n1442), .Z(n1439) );
  NANDN U1697 ( .A(B[257]), .B(n1443), .Z(n1442) );
  NANDN U1698 ( .A(A[257]), .B(n1444), .Z(n1443) );
  NANDN U1699 ( .A(n1444), .B(A[257]), .Z(n1441) );
  XOR U1700 ( .A(n1444), .B(n1445), .Z(DIFF[257]) );
  XOR U1701 ( .A(B[257]), .B(A[257]), .Z(n1445) );
  AND U1702 ( .A(n1446), .B(n1447), .Z(n1444) );
  NANDN U1703 ( .A(B[256]), .B(n1448), .Z(n1447) );
  NANDN U1704 ( .A(A[256]), .B(n1449), .Z(n1448) );
  NANDN U1705 ( .A(n1449), .B(A[256]), .Z(n1446) );
  XOR U1706 ( .A(n1449), .B(n1450), .Z(DIFF[256]) );
  XOR U1707 ( .A(B[256]), .B(A[256]), .Z(n1450) );
  AND U1708 ( .A(n1451), .B(n1452), .Z(n1449) );
  NANDN U1709 ( .A(B[255]), .B(n1453), .Z(n1452) );
  NANDN U1710 ( .A(A[255]), .B(n1454), .Z(n1453) );
  NANDN U1711 ( .A(n1454), .B(A[255]), .Z(n1451) );
  XOR U1712 ( .A(n1454), .B(n1455), .Z(DIFF[255]) );
  XOR U1713 ( .A(B[255]), .B(A[255]), .Z(n1455) );
  AND U1714 ( .A(n1456), .B(n1457), .Z(n1454) );
  NANDN U1715 ( .A(B[254]), .B(n1458), .Z(n1457) );
  NANDN U1716 ( .A(A[254]), .B(n1459), .Z(n1458) );
  NANDN U1717 ( .A(n1459), .B(A[254]), .Z(n1456) );
  XOR U1718 ( .A(n1459), .B(n1460), .Z(DIFF[254]) );
  XOR U1719 ( .A(B[254]), .B(A[254]), .Z(n1460) );
  AND U1720 ( .A(n1461), .B(n1462), .Z(n1459) );
  NANDN U1721 ( .A(B[253]), .B(n1463), .Z(n1462) );
  NANDN U1722 ( .A(A[253]), .B(n1464), .Z(n1463) );
  NANDN U1723 ( .A(n1464), .B(A[253]), .Z(n1461) );
  XOR U1724 ( .A(n1464), .B(n1465), .Z(DIFF[253]) );
  XOR U1725 ( .A(B[253]), .B(A[253]), .Z(n1465) );
  AND U1726 ( .A(n1466), .B(n1467), .Z(n1464) );
  NANDN U1727 ( .A(B[252]), .B(n1468), .Z(n1467) );
  NANDN U1728 ( .A(A[252]), .B(n1469), .Z(n1468) );
  NANDN U1729 ( .A(n1469), .B(A[252]), .Z(n1466) );
  XOR U1730 ( .A(n1469), .B(n1470), .Z(DIFF[252]) );
  XOR U1731 ( .A(B[252]), .B(A[252]), .Z(n1470) );
  AND U1732 ( .A(n1471), .B(n1472), .Z(n1469) );
  NANDN U1733 ( .A(B[251]), .B(n1473), .Z(n1472) );
  NANDN U1734 ( .A(A[251]), .B(n1474), .Z(n1473) );
  NANDN U1735 ( .A(n1474), .B(A[251]), .Z(n1471) );
  XOR U1736 ( .A(n1474), .B(n1475), .Z(DIFF[251]) );
  XOR U1737 ( .A(B[251]), .B(A[251]), .Z(n1475) );
  AND U1738 ( .A(n1476), .B(n1477), .Z(n1474) );
  NANDN U1739 ( .A(B[250]), .B(n1478), .Z(n1477) );
  NANDN U1740 ( .A(A[250]), .B(n1479), .Z(n1478) );
  NANDN U1741 ( .A(n1479), .B(A[250]), .Z(n1476) );
  XOR U1742 ( .A(n1479), .B(n1480), .Z(DIFF[250]) );
  XOR U1743 ( .A(B[250]), .B(A[250]), .Z(n1480) );
  AND U1744 ( .A(n1481), .B(n1482), .Z(n1479) );
  NANDN U1745 ( .A(B[249]), .B(n1483), .Z(n1482) );
  NANDN U1746 ( .A(A[249]), .B(n1484), .Z(n1483) );
  NANDN U1747 ( .A(n1484), .B(A[249]), .Z(n1481) );
  XOR U1748 ( .A(n1485), .B(n1486), .Z(DIFF[24]) );
  XOR U1749 ( .A(B[24]), .B(A[24]), .Z(n1486) );
  XOR U1750 ( .A(n1484), .B(n1487), .Z(DIFF[249]) );
  XOR U1751 ( .A(B[249]), .B(A[249]), .Z(n1487) );
  AND U1752 ( .A(n1488), .B(n1489), .Z(n1484) );
  NANDN U1753 ( .A(B[248]), .B(n1490), .Z(n1489) );
  NANDN U1754 ( .A(A[248]), .B(n1491), .Z(n1490) );
  NANDN U1755 ( .A(n1491), .B(A[248]), .Z(n1488) );
  XOR U1756 ( .A(n1491), .B(n1492), .Z(DIFF[248]) );
  XOR U1757 ( .A(B[248]), .B(A[248]), .Z(n1492) );
  AND U1758 ( .A(n1493), .B(n1494), .Z(n1491) );
  NANDN U1759 ( .A(B[247]), .B(n1495), .Z(n1494) );
  NANDN U1760 ( .A(A[247]), .B(n1496), .Z(n1495) );
  NANDN U1761 ( .A(n1496), .B(A[247]), .Z(n1493) );
  XOR U1762 ( .A(n1496), .B(n1497), .Z(DIFF[247]) );
  XOR U1763 ( .A(B[247]), .B(A[247]), .Z(n1497) );
  AND U1764 ( .A(n1498), .B(n1499), .Z(n1496) );
  NANDN U1765 ( .A(B[246]), .B(n1500), .Z(n1499) );
  NANDN U1766 ( .A(A[246]), .B(n1501), .Z(n1500) );
  NANDN U1767 ( .A(n1501), .B(A[246]), .Z(n1498) );
  XOR U1768 ( .A(n1501), .B(n1502), .Z(DIFF[246]) );
  XOR U1769 ( .A(B[246]), .B(A[246]), .Z(n1502) );
  AND U1770 ( .A(n1503), .B(n1504), .Z(n1501) );
  NANDN U1771 ( .A(B[245]), .B(n1505), .Z(n1504) );
  NANDN U1772 ( .A(A[245]), .B(n1506), .Z(n1505) );
  NANDN U1773 ( .A(n1506), .B(A[245]), .Z(n1503) );
  XOR U1774 ( .A(n1506), .B(n1507), .Z(DIFF[245]) );
  XOR U1775 ( .A(B[245]), .B(A[245]), .Z(n1507) );
  AND U1776 ( .A(n1508), .B(n1509), .Z(n1506) );
  NANDN U1777 ( .A(B[244]), .B(n1510), .Z(n1509) );
  NANDN U1778 ( .A(A[244]), .B(n1511), .Z(n1510) );
  NANDN U1779 ( .A(n1511), .B(A[244]), .Z(n1508) );
  XOR U1780 ( .A(n1511), .B(n1512), .Z(DIFF[244]) );
  XOR U1781 ( .A(B[244]), .B(A[244]), .Z(n1512) );
  AND U1782 ( .A(n1513), .B(n1514), .Z(n1511) );
  NANDN U1783 ( .A(B[243]), .B(n1515), .Z(n1514) );
  NANDN U1784 ( .A(A[243]), .B(n1516), .Z(n1515) );
  NANDN U1785 ( .A(n1516), .B(A[243]), .Z(n1513) );
  XOR U1786 ( .A(n1516), .B(n1517), .Z(DIFF[243]) );
  XOR U1787 ( .A(B[243]), .B(A[243]), .Z(n1517) );
  AND U1788 ( .A(n1518), .B(n1519), .Z(n1516) );
  NANDN U1789 ( .A(B[242]), .B(n1520), .Z(n1519) );
  NANDN U1790 ( .A(A[242]), .B(n1521), .Z(n1520) );
  NANDN U1791 ( .A(n1521), .B(A[242]), .Z(n1518) );
  XOR U1792 ( .A(n1521), .B(n1522), .Z(DIFF[242]) );
  XOR U1793 ( .A(B[242]), .B(A[242]), .Z(n1522) );
  AND U1794 ( .A(n1523), .B(n1524), .Z(n1521) );
  NANDN U1795 ( .A(B[241]), .B(n1525), .Z(n1524) );
  NANDN U1796 ( .A(A[241]), .B(n1526), .Z(n1525) );
  NANDN U1797 ( .A(n1526), .B(A[241]), .Z(n1523) );
  XOR U1798 ( .A(n1526), .B(n1527), .Z(DIFF[241]) );
  XOR U1799 ( .A(B[241]), .B(A[241]), .Z(n1527) );
  AND U1800 ( .A(n1528), .B(n1529), .Z(n1526) );
  NANDN U1801 ( .A(B[240]), .B(n1530), .Z(n1529) );
  NANDN U1802 ( .A(A[240]), .B(n1531), .Z(n1530) );
  NANDN U1803 ( .A(n1531), .B(A[240]), .Z(n1528) );
  XOR U1804 ( .A(n1531), .B(n1532), .Z(DIFF[240]) );
  XOR U1805 ( .A(B[240]), .B(A[240]), .Z(n1532) );
  AND U1806 ( .A(n1533), .B(n1534), .Z(n1531) );
  NANDN U1807 ( .A(B[239]), .B(n1535), .Z(n1534) );
  NANDN U1808 ( .A(A[239]), .B(n1536), .Z(n1535) );
  NANDN U1809 ( .A(n1536), .B(A[239]), .Z(n1533) );
  XOR U1810 ( .A(n1537), .B(n1538), .Z(DIFF[23]) );
  XOR U1811 ( .A(B[23]), .B(A[23]), .Z(n1538) );
  XOR U1812 ( .A(n1536), .B(n1539), .Z(DIFF[239]) );
  XOR U1813 ( .A(B[239]), .B(A[239]), .Z(n1539) );
  AND U1814 ( .A(n1540), .B(n1541), .Z(n1536) );
  NANDN U1815 ( .A(B[238]), .B(n1542), .Z(n1541) );
  NANDN U1816 ( .A(A[238]), .B(n1543), .Z(n1542) );
  NANDN U1817 ( .A(n1543), .B(A[238]), .Z(n1540) );
  XOR U1818 ( .A(n1543), .B(n1544), .Z(DIFF[238]) );
  XOR U1819 ( .A(B[238]), .B(A[238]), .Z(n1544) );
  AND U1820 ( .A(n1545), .B(n1546), .Z(n1543) );
  NANDN U1821 ( .A(B[237]), .B(n1547), .Z(n1546) );
  NANDN U1822 ( .A(A[237]), .B(n1548), .Z(n1547) );
  NANDN U1823 ( .A(n1548), .B(A[237]), .Z(n1545) );
  XOR U1824 ( .A(n1548), .B(n1549), .Z(DIFF[237]) );
  XOR U1825 ( .A(B[237]), .B(A[237]), .Z(n1549) );
  AND U1826 ( .A(n1550), .B(n1551), .Z(n1548) );
  NANDN U1827 ( .A(B[236]), .B(n1552), .Z(n1551) );
  NANDN U1828 ( .A(A[236]), .B(n1553), .Z(n1552) );
  NANDN U1829 ( .A(n1553), .B(A[236]), .Z(n1550) );
  XOR U1830 ( .A(n1553), .B(n1554), .Z(DIFF[236]) );
  XOR U1831 ( .A(B[236]), .B(A[236]), .Z(n1554) );
  AND U1832 ( .A(n1555), .B(n1556), .Z(n1553) );
  NANDN U1833 ( .A(B[235]), .B(n1557), .Z(n1556) );
  NANDN U1834 ( .A(A[235]), .B(n1558), .Z(n1557) );
  NANDN U1835 ( .A(n1558), .B(A[235]), .Z(n1555) );
  XOR U1836 ( .A(n1558), .B(n1559), .Z(DIFF[235]) );
  XOR U1837 ( .A(B[235]), .B(A[235]), .Z(n1559) );
  AND U1838 ( .A(n1560), .B(n1561), .Z(n1558) );
  NANDN U1839 ( .A(B[234]), .B(n1562), .Z(n1561) );
  NANDN U1840 ( .A(A[234]), .B(n1563), .Z(n1562) );
  NANDN U1841 ( .A(n1563), .B(A[234]), .Z(n1560) );
  XOR U1842 ( .A(n1563), .B(n1564), .Z(DIFF[234]) );
  XOR U1843 ( .A(B[234]), .B(A[234]), .Z(n1564) );
  AND U1844 ( .A(n1565), .B(n1566), .Z(n1563) );
  NANDN U1845 ( .A(B[233]), .B(n1567), .Z(n1566) );
  NANDN U1846 ( .A(A[233]), .B(n1568), .Z(n1567) );
  NANDN U1847 ( .A(n1568), .B(A[233]), .Z(n1565) );
  XOR U1848 ( .A(n1568), .B(n1569), .Z(DIFF[233]) );
  XOR U1849 ( .A(B[233]), .B(A[233]), .Z(n1569) );
  AND U1850 ( .A(n1570), .B(n1571), .Z(n1568) );
  NANDN U1851 ( .A(B[232]), .B(n1572), .Z(n1571) );
  NANDN U1852 ( .A(A[232]), .B(n1573), .Z(n1572) );
  NANDN U1853 ( .A(n1573), .B(A[232]), .Z(n1570) );
  XOR U1854 ( .A(n1573), .B(n1574), .Z(DIFF[232]) );
  XOR U1855 ( .A(B[232]), .B(A[232]), .Z(n1574) );
  AND U1856 ( .A(n1575), .B(n1576), .Z(n1573) );
  NANDN U1857 ( .A(B[231]), .B(n1577), .Z(n1576) );
  NANDN U1858 ( .A(A[231]), .B(n1578), .Z(n1577) );
  NANDN U1859 ( .A(n1578), .B(A[231]), .Z(n1575) );
  XOR U1860 ( .A(n1578), .B(n1579), .Z(DIFF[231]) );
  XOR U1861 ( .A(B[231]), .B(A[231]), .Z(n1579) );
  AND U1862 ( .A(n1580), .B(n1581), .Z(n1578) );
  NANDN U1863 ( .A(B[230]), .B(n1582), .Z(n1581) );
  NANDN U1864 ( .A(A[230]), .B(n1583), .Z(n1582) );
  NANDN U1865 ( .A(n1583), .B(A[230]), .Z(n1580) );
  XOR U1866 ( .A(n1583), .B(n1584), .Z(DIFF[230]) );
  XOR U1867 ( .A(B[230]), .B(A[230]), .Z(n1584) );
  AND U1868 ( .A(n1585), .B(n1586), .Z(n1583) );
  NANDN U1869 ( .A(B[229]), .B(n1587), .Z(n1586) );
  NANDN U1870 ( .A(A[229]), .B(n1588), .Z(n1587) );
  NANDN U1871 ( .A(n1588), .B(A[229]), .Z(n1585) );
  XOR U1872 ( .A(n1589), .B(n1590), .Z(DIFF[22]) );
  XOR U1873 ( .A(B[22]), .B(A[22]), .Z(n1590) );
  XOR U1874 ( .A(n1588), .B(n1591), .Z(DIFF[229]) );
  XOR U1875 ( .A(B[229]), .B(A[229]), .Z(n1591) );
  AND U1876 ( .A(n1592), .B(n1593), .Z(n1588) );
  NANDN U1877 ( .A(B[228]), .B(n1594), .Z(n1593) );
  NANDN U1878 ( .A(A[228]), .B(n1595), .Z(n1594) );
  NANDN U1879 ( .A(n1595), .B(A[228]), .Z(n1592) );
  XOR U1880 ( .A(n1595), .B(n1596), .Z(DIFF[228]) );
  XOR U1881 ( .A(B[228]), .B(A[228]), .Z(n1596) );
  AND U1882 ( .A(n1597), .B(n1598), .Z(n1595) );
  NANDN U1883 ( .A(B[227]), .B(n1599), .Z(n1598) );
  NANDN U1884 ( .A(A[227]), .B(n1600), .Z(n1599) );
  NANDN U1885 ( .A(n1600), .B(A[227]), .Z(n1597) );
  XOR U1886 ( .A(n1600), .B(n1601), .Z(DIFF[227]) );
  XOR U1887 ( .A(B[227]), .B(A[227]), .Z(n1601) );
  AND U1888 ( .A(n1602), .B(n1603), .Z(n1600) );
  NANDN U1889 ( .A(B[226]), .B(n1604), .Z(n1603) );
  NANDN U1890 ( .A(A[226]), .B(n1605), .Z(n1604) );
  NANDN U1891 ( .A(n1605), .B(A[226]), .Z(n1602) );
  XOR U1892 ( .A(n1605), .B(n1606), .Z(DIFF[226]) );
  XOR U1893 ( .A(B[226]), .B(A[226]), .Z(n1606) );
  AND U1894 ( .A(n1607), .B(n1608), .Z(n1605) );
  NANDN U1895 ( .A(B[225]), .B(n1609), .Z(n1608) );
  NANDN U1896 ( .A(A[225]), .B(n1610), .Z(n1609) );
  NANDN U1897 ( .A(n1610), .B(A[225]), .Z(n1607) );
  XOR U1898 ( .A(n1610), .B(n1611), .Z(DIFF[225]) );
  XOR U1899 ( .A(B[225]), .B(A[225]), .Z(n1611) );
  AND U1900 ( .A(n1612), .B(n1613), .Z(n1610) );
  NANDN U1901 ( .A(B[224]), .B(n1614), .Z(n1613) );
  NANDN U1902 ( .A(A[224]), .B(n1615), .Z(n1614) );
  NANDN U1903 ( .A(n1615), .B(A[224]), .Z(n1612) );
  XOR U1904 ( .A(n1615), .B(n1616), .Z(DIFF[224]) );
  XOR U1905 ( .A(B[224]), .B(A[224]), .Z(n1616) );
  AND U1906 ( .A(n1617), .B(n1618), .Z(n1615) );
  NANDN U1907 ( .A(B[223]), .B(n1619), .Z(n1618) );
  NANDN U1908 ( .A(A[223]), .B(n1620), .Z(n1619) );
  NANDN U1909 ( .A(n1620), .B(A[223]), .Z(n1617) );
  XOR U1910 ( .A(n1620), .B(n1621), .Z(DIFF[223]) );
  XOR U1911 ( .A(B[223]), .B(A[223]), .Z(n1621) );
  AND U1912 ( .A(n1622), .B(n1623), .Z(n1620) );
  NANDN U1913 ( .A(B[222]), .B(n1624), .Z(n1623) );
  NANDN U1914 ( .A(A[222]), .B(n1625), .Z(n1624) );
  NANDN U1915 ( .A(n1625), .B(A[222]), .Z(n1622) );
  XOR U1916 ( .A(n1625), .B(n1626), .Z(DIFF[222]) );
  XOR U1917 ( .A(B[222]), .B(A[222]), .Z(n1626) );
  AND U1918 ( .A(n1627), .B(n1628), .Z(n1625) );
  NANDN U1919 ( .A(B[221]), .B(n1629), .Z(n1628) );
  NANDN U1920 ( .A(A[221]), .B(n1630), .Z(n1629) );
  NANDN U1921 ( .A(n1630), .B(A[221]), .Z(n1627) );
  XOR U1922 ( .A(n1630), .B(n1631), .Z(DIFF[221]) );
  XOR U1923 ( .A(B[221]), .B(A[221]), .Z(n1631) );
  AND U1924 ( .A(n1632), .B(n1633), .Z(n1630) );
  NANDN U1925 ( .A(B[220]), .B(n1634), .Z(n1633) );
  NANDN U1926 ( .A(A[220]), .B(n1635), .Z(n1634) );
  NANDN U1927 ( .A(n1635), .B(A[220]), .Z(n1632) );
  XOR U1928 ( .A(n1635), .B(n1636), .Z(DIFF[220]) );
  XOR U1929 ( .A(B[220]), .B(A[220]), .Z(n1636) );
  AND U1930 ( .A(n1637), .B(n1638), .Z(n1635) );
  NANDN U1931 ( .A(B[219]), .B(n1639), .Z(n1638) );
  NANDN U1932 ( .A(A[219]), .B(n1640), .Z(n1639) );
  NANDN U1933 ( .A(n1640), .B(A[219]), .Z(n1637) );
  XOR U1934 ( .A(n1641), .B(n1642), .Z(DIFF[21]) );
  XOR U1935 ( .A(B[21]), .B(A[21]), .Z(n1642) );
  XOR U1936 ( .A(n1640), .B(n1643), .Z(DIFF[219]) );
  XOR U1937 ( .A(B[219]), .B(A[219]), .Z(n1643) );
  AND U1938 ( .A(n1644), .B(n1645), .Z(n1640) );
  NANDN U1939 ( .A(B[218]), .B(n1646), .Z(n1645) );
  NANDN U1940 ( .A(A[218]), .B(n1647), .Z(n1646) );
  NANDN U1941 ( .A(n1647), .B(A[218]), .Z(n1644) );
  XOR U1942 ( .A(n1647), .B(n1648), .Z(DIFF[218]) );
  XOR U1943 ( .A(B[218]), .B(A[218]), .Z(n1648) );
  AND U1944 ( .A(n1649), .B(n1650), .Z(n1647) );
  NANDN U1945 ( .A(B[217]), .B(n1651), .Z(n1650) );
  NANDN U1946 ( .A(A[217]), .B(n1652), .Z(n1651) );
  NANDN U1947 ( .A(n1652), .B(A[217]), .Z(n1649) );
  XOR U1948 ( .A(n1652), .B(n1653), .Z(DIFF[217]) );
  XOR U1949 ( .A(B[217]), .B(A[217]), .Z(n1653) );
  AND U1950 ( .A(n1654), .B(n1655), .Z(n1652) );
  NANDN U1951 ( .A(B[216]), .B(n1656), .Z(n1655) );
  NANDN U1952 ( .A(A[216]), .B(n1657), .Z(n1656) );
  NANDN U1953 ( .A(n1657), .B(A[216]), .Z(n1654) );
  XOR U1954 ( .A(n1657), .B(n1658), .Z(DIFF[216]) );
  XOR U1955 ( .A(B[216]), .B(A[216]), .Z(n1658) );
  AND U1956 ( .A(n1659), .B(n1660), .Z(n1657) );
  NANDN U1957 ( .A(B[215]), .B(n1661), .Z(n1660) );
  NANDN U1958 ( .A(A[215]), .B(n1662), .Z(n1661) );
  NANDN U1959 ( .A(n1662), .B(A[215]), .Z(n1659) );
  XOR U1960 ( .A(n1662), .B(n1663), .Z(DIFF[215]) );
  XOR U1961 ( .A(B[215]), .B(A[215]), .Z(n1663) );
  AND U1962 ( .A(n1664), .B(n1665), .Z(n1662) );
  NANDN U1963 ( .A(B[214]), .B(n1666), .Z(n1665) );
  NANDN U1964 ( .A(A[214]), .B(n1667), .Z(n1666) );
  NANDN U1965 ( .A(n1667), .B(A[214]), .Z(n1664) );
  XOR U1966 ( .A(n1667), .B(n1668), .Z(DIFF[214]) );
  XOR U1967 ( .A(B[214]), .B(A[214]), .Z(n1668) );
  AND U1968 ( .A(n1669), .B(n1670), .Z(n1667) );
  NANDN U1969 ( .A(B[213]), .B(n1671), .Z(n1670) );
  NANDN U1970 ( .A(A[213]), .B(n1672), .Z(n1671) );
  NANDN U1971 ( .A(n1672), .B(A[213]), .Z(n1669) );
  XOR U1972 ( .A(n1672), .B(n1673), .Z(DIFF[213]) );
  XOR U1973 ( .A(B[213]), .B(A[213]), .Z(n1673) );
  AND U1974 ( .A(n1674), .B(n1675), .Z(n1672) );
  NANDN U1975 ( .A(B[212]), .B(n1676), .Z(n1675) );
  NANDN U1976 ( .A(A[212]), .B(n1677), .Z(n1676) );
  NANDN U1977 ( .A(n1677), .B(A[212]), .Z(n1674) );
  XOR U1978 ( .A(n1677), .B(n1678), .Z(DIFF[212]) );
  XOR U1979 ( .A(B[212]), .B(A[212]), .Z(n1678) );
  AND U1980 ( .A(n1679), .B(n1680), .Z(n1677) );
  NANDN U1981 ( .A(B[211]), .B(n1681), .Z(n1680) );
  NANDN U1982 ( .A(A[211]), .B(n1682), .Z(n1681) );
  NANDN U1983 ( .A(n1682), .B(A[211]), .Z(n1679) );
  XOR U1984 ( .A(n1682), .B(n1683), .Z(DIFF[211]) );
  XOR U1985 ( .A(B[211]), .B(A[211]), .Z(n1683) );
  AND U1986 ( .A(n1684), .B(n1685), .Z(n1682) );
  NANDN U1987 ( .A(B[210]), .B(n1686), .Z(n1685) );
  NANDN U1988 ( .A(A[210]), .B(n1687), .Z(n1686) );
  NANDN U1989 ( .A(n1687), .B(A[210]), .Z(n1684) );
  XOR U1990 ( .A(n1687), .B(n1688), .Z(DIFF[210]) );
  XOR U1991 ( .A(B[210]), .B(A[210]), .Z(n1688) );
  AND U1992 ( .A(n1689), .B(n1690), .Z(n1687) );
  NANDN U1993 ( .A(B[209]), .B(n1691), .Z(n1690) );
  NANDN U1994 ( .A(A[209]), .B(n1692), .Z(n1691) );
  NANDN U1995 ( .A(n1692), .B(A[209]), .Z(n1689) );
  XOR U1996 ( .A(n1693), .B(n1694), .Z(DIFF[20]) );
  XOR U1997 ( .A(B[20]), .B(A[20]), .Z(n1694) );
  XOR U1998 ( .A(n1692), .B(n1695), .Z(DIFF[209]) );
  XOR U1999 ( .A(B[209]), .B(A[209]), .Z(n1695) );
  AND U2000 ( .A(n1696), .B(n1697), .Z(n1692) );
  NANDN U2001 ( .A(B[208]), .B(n1698), .Z(n1697) );
  NANDN U2002 ( .A(A[208]), .B(n1699), .Z(n1698) );
  NANDN U2003 ( .A(n1699), .B(A[208]), .Z(n1696) );
  XOR U2004 ( .A(n1699), .B(n1700), .Z(DIFF[208]) );
  XOR U2005 ( .A(B[208]), .B(A[208]), .Z(n1700) );
  AND U2006 ( .A(n1701), .B(n1702), .Z(n1699) );
  NANDN U2007 ( .A(B[207]), .B(n1703), .Z(n1702) );
  NANDN U2008 ( .A(A[207]), .B(n1704), .Z(n1703) );
  NANDN U2009 ( .A(n1704), .B(A[207]), .Z(n1701) );
  XOR U2010 ( .A(n1704), .B(n1705), .Z(DIFF[207]) );
  XOR U2011 ( .A(B[207]), .B(A[207]), .Z(n1705) );
  AND U2012 ( .A(n1706), .B(n1707), .Z(n1704) );
  NANDN U2013 ( .A(B[206]), .B(n1708), .Z(n1707) );
  NANDN U2014 ( .A(A[206]), .B(n1709), .Z(n1708) );
  NANDN U2015 ( .A(n1709), .B(A[206]), .Z(n1706) );
  XOR U2016 ( .A(n1709), .B(n1710), .Z(DIFF[206]) );
  XOR U2017 ( .A(B[206]), .B(A[206]), .Z(n1710) );
  AND U2018 ( .A(n1711), .B(n1712), .Z(n1709) );
  NANDN U2019 ( .A(B[205]), .B(n1713), .Z(n1712) );
  NANDN U2020 ( .A(A[205]), .B(n1714), .Z(n1713) );
  NANDN U2021 ( .A(n1714), .B(A[205]), .Z(n1711) );
  XOR U2022 ( .A(n1714), .B(n1715), .Z(DIFF[205]) );
  XOR U2023 ( .A(B[205]), .B(A[205]), .Z(n1715) );
  AND U2024 ( .A(n1716), .B(n1717), .Z(n1714) );
  NANDN U2025 ( .A(B[204]), .B(n1718), .Z(n1717) );
  NANDN U2026 ( .A(A[204]), .B(n1719), .Z(n1718) );
  NANDN U2027 ( .A(n1719), .B(A[204]), .Z(n1716) );
  XOR U2028 ( .A(n1719), .B(n1720), .Z(DIFF[204]) );
  XOR U2029 ( .A(B[204]), .B(A[204]), .Z(n1720) );
  AND U2030 ( .A(n1721), .B(n1722), .Z(n1719) );
  NANDN U2031 ( .A(B[203]), .B(n1723), .Z(n1722) );
  NANDN U2032 ( .A(A[203]), .B(n1724), .Z(n1723) );
  NANDN U2033 ( .A(n1724), .B(A[203]), .Z(n1721) );
  XOR U2034 ( .A(n1724), .B(n1725), .Z(DIFF[203]) );
  XOR U2035 ( .A(B[203]), .B(A[203]), .Z(n1725) );
  AND U2036 ( .A(n1726), .B(n1727), .Z(n1724) );
  NANDN U2037 ( .A(B[202]), .B(n1728), .Z(n1727) );
  NANDN U2038 ( .A(A[202]), .B(n1729), .Z(n1728) );
  NANDN U2039 ( .A(n1729), .B(A[202]), .Z(n1726) );
  XOR U2040 ( .A(n1729), .B(n1730), .Z(DIFF[202]) );
  XOR U2041 ( .A(B[202]), .B(A[202]), .Z(n1730) );
  AND U2042 ( .A(n1731), .B(n1732), .Z(n1729) );
  NANDN U2043 ( .A(B[201]), .B(n1733), .Z(n1732) );
  NANDN U2044 ( .A(A[201]), .B(n1734), .Z(n1733) );
  NANDN U2045 ( .A(n1734), .B(A[201]), .Z(n1731) );
  XOR U2046 ( .A(n1734), .B(n1735), .Z(DIFF[201]) );
  XOR U2047 ( .A(B[201]), .B(A[201]), .Z(n1735) );
  AND U2048 ( .A(n1736), .B(n1737), .Z(n1734) );
  NANDN U2049 ( .A(B[200]), .B(n1738), .Z(n1737) );
  NANDN U2050 ( .A(A[200]), .B(n1739), .Z(n1738) );
  NANDN U2051 ( .A(n1739), .B(A[200]), .Z(n1736) );
  XOR U2052 ( .A(n1739), .B(n1740), .Z(DIFF[200]) );
  XOR U2053 ( .A(B[200]), .B(A[200]), .Z(n1740) );
  AND U2054 ( .A(n1741), .B(n1742), .Z(n1739) );
  NANDN U2055 ( .A(B[199]), .B(n1743), .Z(n1742) );
  NANDN U2056 ( .A(A[199]), .B(n1744), .Z(n1743) );
  NANDN U2057 ( .A(n1744), .B(A[199]), .Z(n1741) );
  XOR U2058 ( .A(n2), .B(n1745), .Z(DIFF[1]) );
  XOR U2059 ( .A(B[1]), .B(A[1]), .Z(n1745) );
  XOR U2060 ( .A(n1746), .B(n1747), .Z(DIFF[19]) );
  XOR U2061 ( .A(B[19]), .B(A[19]), .Z(n1747) );
  XOR U2062 ( .A(n1744), .B(n1748), .Z(DIFF[199]) );
  XOR U2063 ( .A(B[199]), .B(A[199]), .Z(n1748) );
  AND U2064 ( .A(n1749), .B(n1750), .Z(n1744) );
  NANDN U2065 ( .A(B[198]), .B(n1751), .Z(n1750) );
  NANDN U2066 ( .A(A[198]), .B(n1752), .Z(n1751) );
  NANDN U2067 ( .A(n1752), .B(A[198]), .Z(n1749) );
  XOR U2068 ( .A(n1752), .B(n1753), .Z(DIFF[198]) );
  XOR U2069 ( .A(B[198]), .B(A[198]), .Z(n1753) );
  AND U2070 ( .A(n1754), .B(n1755), .Z(n1752) );
  NANDN U2071 ( .A(B[197]), .B(n1756), .Z(n1755) );
  NANDN U2072 ( .A(A[197]), .B(n1757), .Z(n1756) );
  NANDN U2073 ( .A(n1757), .B(A[197]), .Z(n1754) );
  XOR U2074 ( .A(n1757), .B(n1758), .Z(DIFF[197]) );
  XOR U2075 ( .A(B[197]), .B(A[197]), .Z(n1758) );
  AND U2076 ( .A(n1759), .B(n1760), .Z(n1757) );
  NANDN U2077 ( .A(B[196]), .B(n1761), .Z(n1760) );
  NANDN U2078 ( .A(A[196]), .B(n1762), .Z(n1761) );
  NANDN U2079 ( .A(n1762), .B(A[196]), .Z(n1759) );
  XOR U2080 ( .A(n1762), .B(n1763), .Z(DIFF[196]) );
  XOR U2081 ( .A(B[196]), .B(A[196]), .Z(n1763) );
  AND U2082 ( .A(n1764), .B(n1765), .Z(n1762) );
  NANDN U2083 ( .A(B[195]), .B(n1766), .Z(n1765) );
  NANDN U2084 ( .A(A[195]), .B(n1767), .Z(n1766) );
  NANDN U2085 ( .A(n1767), .B(A[195]), .Z(n1764) );
  XOR U2086 ( .A(n1767), .B(n1768), .Z(DIFF[195]) );
  XOR U2087 ( .A(B[195]), .B(A[195]), .Z(n1768) );
  AND U2088 ( .A(n1769), .B(n1770), .Z(n1767) );
  NANDN U2089 ( .A(B[194]), .B(n1771), .Z(n1770) );
  NANDN U2090 ( .A(A[194]), .B(n1772), .Z(n1771) );
  NANDN U2091 ( .A(n1772), .B(A[194]), .Z(n1769) );
  XOR U2092 ( .A(n1772), .B(n1773), .Z(DIFF[194]) );
  XOR U2093 ( .A(B[194]), .B(A[194]), .Z(n1773) );
  AND U2094 ( .A(n1774), .B(n1775), .Z(n1772) );
  NANDN U2095 ( .A(B[193]), .B(n1776), .Z(n1775) );
  NANDN U2096 ( .A(A[193]), .B(n1777), .Z(n1776) );
  NANDN U2097 ( .A(n1777), .B(A[193]), .Z(n1774) );
  XOR U2098 ( .A(n1777), .B(n1778), .Z(DIFF[193]) );
  XOR U2099 ( .A(B[193]), .B(A[193]), .Z(n1778) );
  AND U2100 ( .A(n1779), .B(n1780), .Z(n1777) );
  NANDN U2101 ( .A(B[192]), .B(n1781), .Z(n1780) );
  NANDN U2102 ( .A(A[192]), .B(n1782), .Z(n1781) );
  NANDN U2103 ( .A(n1782), .B(A[192]), .Z(n1779) );
  XOR U2104 ( .A(n1782), .B(n1783), .Z(DIFF[192]) );
  XOR U2105 ( .A(B[192]), .B(A[192]), .Z(n1783) );
  AND U2106 ( .A(n1784), .B(n1785), .Z(n1782) );
  NANDN U2107 ( .A(B[191]), .B(n1786), .Z(n1785) );
  NANDN U2108 ( .A(A[191]), .B(n1787), .Z(n1786) );
  NANDN U2109 ( .A(n1787), .B(A[191]), .Z(n1784) );
  XOR U2110 ( .A(n1787), .B(n1788), .Z(DIFF[191]) );
  XOR U2111 ( .A(B[191]), .B(A[191]), .Z(n1788) );
  AND U2112 ( .A(n1789), .B(n1790), .Z(n1787) );
  NANDN U2113 ( .A(B[190]), .B(n1791), .Z(n1790) );
  NANDN U2114 ( .A(A[190]), .B(n1792), .Z(n1791) );
  NANDN U2115 ( .A(n1792), .B(A[190]), .Z(n1789) );
  XOR U2116 ( .A(n1792), .B(n1793), .Z(DIFF[190]) );
  XOR U2117 ( .A(B[190]), .B(A[190]), .Z(n1793) );
  AND U2118 ( .A(n1794), .B(n1795), .Z(n1792) );
  NANDN U2119 ( .A(B[189]), .B(n1796), .Z(n1795) );
  NANDN U2120 ( .A(A[189]), .B(n1797), .Z(n1796) );
  NANDN U2121 ( .A(n1797), .B(A[189]), .Z(n1794) );
  XOR U2122 ( .A(n1798), .B(n1799), .Z(DIFF[18]) );
  XOR U2123 ( .A(B[18]), .B(A[18]), .Z(n1799) );
  XOR U2124 ( .A(n1797), .B(n1800), .Z(DIFF[189]) );
  XOR U2125 ( .A(B[189]), .B(A[189]), .Z(n1800) );
  AND U2126 ( .A(n1801), .B(n1802), .Z(n1797) );
  NANDN U2127 ( .A(B[188]), .B(n1803), .Z(n1802) );
  NANDN U2128 ( .A(A[188]), .B(n1804), .Z(n1803) );
  NANDN U2129 ( .A(n1804), .B(A[188]), .Z(n1801) );
  XOR U2130 ( .A(n1804), .B(n1805), .Z(DIFF[188]) );
  XOR U2131 ( .A(B[188]), .B(A[188]), .Z(n1805) );
  AND U2132 ( .A(n1806), .B(n1807), .Z(n1804) );
  NANDN U2133 ( .A(B[187]), .B(n1808), .Z(n1807) );
  NANDN U2134 ( .A(A[187]), .B(n1809), .Z(n1808) );
  NANDN U2135 ( .A(n1809), .B(A[187]), .Z(n1806) );
  XOR U2136 ( .A(n1809), .B(n1810), .Z(DIFF[187]) );
  XOR U2137 ( .A(B[187]), .B(A[187]), .Z(n1810) );
  AND U2138 ( .A(n1811), .B(n1812), .Z(n1809) );
  NANDN U2139 ( .A(B[186]), .B(n1813), .Z(n1812) );
  NANDN U2140 ( .A(A[186]), .B(n1814), .Z(n1813) );
  NANDN U2141 ( .A(n1814), .B(A[186]), .Z(n1811) );
  XOR U2142 ( .A(n1814), .B(n1815), .Z(DIFF[186]) );
  XOR U2143 ( .A(B[186]), .B(A[186]), .Z(n1815) );
  AND U2144 ( .A(n1816), .B(n1817), .Z(n1814) );
  NANDN U2145 ( .A(B[185]), .B(n1818), .Z(n1817) );
  NANDN U2146 ( .A(A[185]), .B(n1819), .Z(n1818) );
  NANDN U2147 ( .A(n1819), .B(A[185]), .Z(n1816) );
  XOR U2148 ( .A(n1819), .B(n1820), .Z(DIFF[185]) );
  XOR U2149 ( .A(B[185]), .B(A[185]), .Z(n1820) );
  AND U2150 ( .A(n1821), .B(n1822), .Z(n1819) );
  NANDN U2151 ( .A(B[184]), .B(n1823), .Z(n1822) );
  NANDN U2152 ( .A(A[184]), .B(n1824), .Z(n1823) );
  NANDN U2153 ( .A(n1824), .B(A[184]), .Z(n1821) );
  XOR U2154 ( .A(n1824), .B(n1825), .Z(DIFF[184]) );
  XOR U2155 ( .A(B[184]), .B(A[184]), .Z(n1825) );
  AND U2156 ( .A(n1826), .B(n1827), .Z(n1824) );
  NANDN U2157 ( .A(B[183]), .B(n1828), .Z(n1827) );
  NANDN U2158 ( .A(A[183]), .B(n1829), .Z(n1828) );
  NANDN U2159 ( .A(n1829), .B(A[183]), .Z(n1826) );
  XOR U2160 ( .A(n1829), .B(n1830), .Z(DIFF[183]) );
  XOR U2161 ( .A(B[183]), .B(A[183]), .Z(n1830) );
  AND U2162 ( .A(n1831), .B(n1832), .Z(n1829) );
  NANDN U2163 ( .A(B[182]), .B(n1833), .Z(n1832) );
  NANDN U2164 ( .A(A[182]), .B(n1834), .Z(n1833) );
  NANDN U2165 ( .A(n1834), .B(A[182]), .Z(n1831) );
  XOR U2166 ( .A(n1834), .B(n1835), .Z(DIFF[182]) );
  XOR U2167 ( .A(B[182]), .B(A[182]), .Z(n1835) );
  AND U2168 ( .A(n1836), .B(n1837), .Z(n1834) );
  NANDN U2169 ( .A(B[181]), .B(n1838), .Z(n1837) );
  NANDN U2170 ( .A(A[181]), .B(n1839), .Z(n1838) );
  NANDN U2171 ( .A(n1839), .B(A[181]), .Z(n1836) );
  XOR U2172 ( .A(n1839), .B(n1840), .Z(DIFF[181]) );
  XOR U2173 ( .A(B[181]), .B(A[181]), .Z(n1840) );
  AND U2174 ( .A(n1841), .B(n1842), .Z(n1839) );
  NANDN U2175 ( .A(B[180]), .B(n1843), .Z(n1842) );
  NANDN U2176 ( .A(A[180]), .B(n1844), .Z(n1843) );
  NANDN U2177 ( .A(n1844), .B(A[180]), .Z(n1841) );
  XOR U2178 ( .A(n1844), .B(n1845), .Z(DIFF[180]) );
  XOR U2179 ( .A(B[180]), .B(A[180]), .Z(n1845) );
  AND U2180 ( .A(n1846), .B(n1847), .Z(n1844) );
  NANDN U2181 ( .A(B[179]), .B(n1848), .Z(n1847) );
  NANDN U2182 ( .A(A[179]), .B(n1849), .Z(n1848) );
  NANDN U2183 ( .A(n1849), .B(A[179]), .Z(n1846) );
  XOR U2184 ( .A(n1850), .B(n1851), .Z(DIFF[17]) );
  XOR U2185 ( .A(B[17]), .B(A[17]), .Z(n1851) );
  XOR U2186 ( .A(n1849), .B(n1852), .Z(DIFF[179]) );
  XOR U2187 ( .A(B[179]), .B(A[179]), .Z(n1852) );
  AND U2188 ( .A(n1853), .B(n1854), .Z(n1849) );
  NANDN U2189 ( .A(B[178]), .B(n1855), .Z(n1854) );
  NANDN U2190 ( .A(A[178]), .B(n1856), .Z(n1855) );
  NANDN U2191 ( .A(n1856), .B(A[178]), .Z(n1853) );
  XOR U2192 ( .A(n1856), .B(n1857), .Z(DIFF[178]) );
  XOR U2193 ( .A(B[178]), .B(A[178]), .Z(n1857) );
  AND U2194 ( .A(n1858), .B(n1859), .Z(n1856) );
  NANDN U2195 ( .A(B[177]), .B(n1860), .Z(n1859) );
  NANDN U2196 ( .A(A[177]), .B(n1861), .Z(n1860) );
  NANDN U2197 ( .A(n1861), .B(A[177]), .Z(n1858) );
  XOR U2198 ( .A(n1861), .B(n1862), .Z(DIFF[177]) );
  XOR U2199 ( .A(B[177]), .B(A[177]), .Z(n1862) );
  AND U2200 ( .A(n1863), .B(n1864), .Z(n1861) );
  NANDN U2201 ( .A(B[176]), .B(n1865), .Z(n1864) );
  NANDN U2202 ( .A(A[176]), .B(n1866), .Z(n1865) );
  NANDN U2203 ( .A(n1866), .B(A[176]), .Z(n1863) );
  XOR U2204 ( .A(n1866), .B(n1867), .Z(DIFF[176]) );
  XOR U2205 ( .A(B[176]), .B(A[176]), .Z(n1867) );
  AND U2206 ( .A(n1868), .B(n1869), .Z(n1866) );
  NANDN U2207 ( .A(B[175]), .B(n1870), .Z(n1869) );
  NANDN U2208 ( .A(A[175]), .B(n1871), .Z(n1870) );
  NANDN U2209 ( .A(n1871), .B(A[175]), .Z(n1868) );
  XOR U2210 ( .A(n1871), .B(n1872), .Z(DIFF[175]) );
  XOR U2211 ( .A(B[175]), .B(A[175]), .Z(n1872) );
  AND U2212 ( .A(n1873), .B(n1874), .Z(n1871) );
  NANDN U2213 ( .A(B[174]), .B(n1875), .Z(n1874) );
  NANDN U2214 ( .A(A[174]), .B(n1876), .Z(n1875) );
  NANDN U2215 ( .A(n1876), .B(A[174]), .Z(n1873) );
  XOR U2216 ( .A(n1876), .B(n1877), .Z(DIFF[174]) );
  XOR U2217 ( .A(B[174]), .B(A[174]), .Z(n1877) );
  AND U2218 ( .A(n1878), .B(n1879), .Z(n1876) );
  NANDN U2219 ( .A(B[173]), .B(n1880), .Z(n1879) );
  NANDN U2220 ( .A(A[173]), .B(n1881), .Z(n1880) );
  NANDN U2221 ( .A(n1881), .B(A[173]), .Z(n1878) );
  XOR U2222 ( .A(n1881), .B(n1882), .Z(DIFF[173]) );
  XOR U2223 ( .A(B[173]), .B(A[173]), .Z(n1882) );
  AND U2224 ( .A(n1883), .B(n1884), .Z(n1881) );
  NANDN U2225 ( .A(B[172]), .B(n1885), .Z(n1884) );
  NANDN U2226 ( .A(A[172]), .B(n1886), .Z(n1885) );
  NANDN U2227 ( .A(n1886), .B(A[172]), .Z(n1883) );
  XOR U2228 ( .A(n1886), .B(n1887), .Z(DIFF[172]) );
  XOR U2229 ( .A(B[172]), .B(A[172]), .Z(n1887) );
  AND U2230 ( .A(n1888), .B(n1889), .Z(n1886) );
  NANDN U2231 ( .A(B[171]), .B(n1890), .Z(n1889) );
  NANDN U2232 ( .A(A[171]), .B(n1891), .Z(n1890) );
  NANDN U2233 ( .A(n1891), .B(A[171]), .Z(n1888) );
  XOR U2234 ( .A(n1891), .B(n1892), .Z(DIFF[171]) );
  XOR U2235 ( .A(B[171]), .B(A[171]), .Z(n1892) );
  AND U2236 ( .A(n1893), .B(n1894), .Z(n1891) );
  NANDN U2237 ( .A(B[170]), .B(n1895), .Z(n1894) );
  NANDN U2238 ( .A(A[170]), .B(n1896), .Z(n1895) );
  NANDN U2239 ( .A(n1896), .B(A[170]), .Z(n1893) );
  XOR U2240 ( .A(n1896), .B(n1897), .Z(DIFF[170]) );
  XOR U2241 ( .A(B[170]), .B(A[170]), .Z(n1897) );
  AND U2242 ( .A(n1898), .B(n1899), .Z(n1896) );
  NANDN U2243 ( .A(B[169]), .B(n1900), .Z(n1899) );
  NANDN U2244 ( .A(A[169]), .B(n1901), .Z(n1900) );
  NANDN U2245 ( .A(n1901), .B(A[169]), .Z(n1898) );
  XOR U2246 ( .A(n1902), .B(n1903), .Z(DIFF[16]) );
  XOR U2247 ( .A(B[16]), .B(A[16]), .Z(n1903) );
  XOR U2248 ( .A(n1901), .B(n1904), .Z(DIFF[169]) );
  XOR U2249 ( .A(B[169]), .B(A[169]), .Z(n1904) );
  AND U2250 ( .A(n1905), .B(n1906), .Z(n1901) );
  NANDN U2251 ( .A(B[168]), .B(n1907), .Z(n1906) );
  NANDN U2252 ( .A(A[168]), .B(n1908), .Z(n1907) );
  NANDN U2253 ( .A(n1908), .B(A[168]), .Z(n1905) );
  XOR U2254 ( .A(n1908), .B(n1909), .Z(DIFF[168]) );
  XOR U2255 ( .A(B[168]), .B(A[168]), .Z(n1909) );
  AND U2256 ( .A(n1910), .B(n1911), .Z(n1908) );
  NANDN U2257 ( .A(B[167]), .B(n1912), .Z(n1911) );
  NANDN U2258 ( .A(A[167]), .B(n1913), .Z(n1912) );
  NANDN U2259 ( .A(n1913), .B(A[167]), .Z(n1910) );
  XOR U2260 ( .A(n1913), .B(n1914), .Z(DIFF[167]) );
  XOR U2261 ( .A(B[167]), .B(A[167]), .Z(n1914) );
  AND U2262 ( .A(n1915), .B(n1916), .Z(n1913) );
  NANDN U2263 ( .A(B[166]), .B(n1917), .Z(n1916) );
  NANDN U2264 ( .A(A[166]), .B(n1918), .Z(n1917) );
  NANDN U2265 ( .A(n1918), .B(A[166]), .Z(n1915) );
  XOR U2266 ( .A(n1918), .B(n1919), .Z(DIFF[166]) );
  XOR U2267 ( .A(B[166]), .B(A[166]), .Z(n1919) );
  AND U2268 ( .A(n1920), .B(n1921), .Z(n1918) );
  NANDN U2269 ( .A(B[165]), .B(n1922), .Z(n1921) );
  NANDN U2270 ( .A(A[165]), .B(n1923), .Z(n1922) );
  NANDN U2271 ( .A(n1923), .B(A[165]), .Z(n1920) );
  XOR U2272 ( .A(n1923), .B(n1924), .Z(DIFF[165]) );
  XOR U2273 ( .A(B[165]), .B(A[165]), .Z(n1924) );
  AND U2274 ( .A(n1925), .B(n1926), .Z(n1923) );
  NANDN U2275 ( .A(B[164]), .B(n1927), .Z(n1926) );
  NANDN U2276 ( .A(A[164]), .B(n1928), .Z(n1927) );
  NANDN U2277 ( .A(n1928), .B(A[164]), .Z(n1925) );
  XOR U2278 ( .A(n1928), .B(n1929), .Z(DIFF[164]) );
  XOR U2279 ( .A(B[164]), .B(A[164]), .Z(n1929) );
  AND U2280 ( .A(n1930), .B(n1931), .Z(n1928) );
  NANDN U2281 ( .A(B[163]), .B(n1932), .Z(n1931) );
  NANDN U2282 ( .A(A[163]), .B(n1933), .Z(n1932) );
  NANDN U2283 ( .A(n1933), .B(A[163]), .Z(n1930) );
  XOR U2284 ( .A(n1933), .B(n1934), .Z(DIFF[163]) );
  XOR U2285 ( .A(B[163]), .B(A[163]), .Z(n1934) );
  AND U2286 ( .A(n1935), .B(n1936), .Z(n1933) );
  NANDN U2287 ( .A(B[162]), .B(n1937), .Z(n1936) );
  NANDN U2288 ( .A(A[162]), .B(n1938), .Z(n1937) );
  NANDN U2289 ( .A(n1938), .B(A[162]), .Z(n1935) );
  XOR U2290 ( .A(n1938), .B(n1939), .Z(DIFF[162]) );
  XOR U2291 ( .A(B[162]), .B(A[162]), .Z(n1939) );
  AND U2292 ( .A(n1940), .B(n1941), .Z(n1938) );
  NANDN U2293 ( .A(B[161]), .B(n1942), .Z(n1941) );
  NANDN U2294 ( .A(A[161]), .B(n1943), .Z(n1942) );
  NANDN U2295 ( .A(n1943), .B(A[161]), .Z(n1940) );
  XOR U2296 ( .A(n1943), .B(n1944), .Z(DIFF[161]) );
  XOR U2297 ( .A(B[161]), .B(A[161]), .Z(n1944) );
  AND U2298 ( .A(n1945), .B(n1946), .Z(n1943) );
  NANDN U2299 ( .A(B[160]), .B(n1947), .Z(n1946) );
  NANDN U2300 ( .A(A[160]), .B(n1948), .Z(n1947) );
  NANDN U2301 ( .A(n1948), .B(A[160]), .Z(n1945) );
  XOR U2302 ( .A(n1948), .B(n1949), .Z(DIFF[160]) );
  XOR U2303 ( .A(B[160]), .B(A[160]), .Z(n1949) );
  AND U2304 ( .A(n1950), .B(n1951), .Z(n1948) );
  NANDN U2305 ( .A(B[159]), .B(n1952), .Z(n1951) );
  NANDN U2306 ( .A(A[159]), .B(n1953), .Z(n1952) );
  NANDN U2307 ( .A(n1953), .B(A[159]), .Z(n1950) );
  XOR U2308 ( .A(n1954), .B(n1955), .Z(DIFF[15]) );
  XOR U2309 ( .A(B[15]), .B(A[15]), .Z(n1955) );
  XOR U2310 ( .A(n1953), .B(n1956), .Z(DIFF[159]) );
  XOR U2311 ( .A(B[159]), .B(A[159]), .Z(n1956) );
  AND U2312 ( .A(n1957), .B(n1958), .Z(n1953) );
  NANDN U2313 ( .A(B[158]), .B(n1959), .Z(n1958) );
  NANDN U2314 ( .A(A[158]), .B(n1960), .Z(n1959) );
  NANDN U2315 ( .A(n1960), .B(A[158]), .Z(n1957) );
  XOR U2316 ( .A(n1960), .B(n1961), .Z(DIFF[158]) );
  XOR U2317 ( .A(B[158]), .B(A[158]), .Z(n1961) );
  AND U2318 ( .A(n1962), .B(n1963), .Z(n1960) );
  NANDN U2319 ( .A(B[157]), .B(n1964), .Z(n1963) );
  NANDN U2320 ( .A(A[157]), .B(n1965), .Z(n1964) );
  NANDN U2321 ( .A(n1965), .B(A[157]), .Z(n1962) );
  XOR U2322 ( .A(n1965), .B(n1966), .Z(DIFF[157]) );
  XOR U2323 ( .A(B[157]), .B(A[157]), .Z(n1966) );
  AND U2324 ( .A(n1967), .B(n1968), .Z(n1965) );
  NANDN U2325 ( .A(B[156]), .B(n1969), .Z(n1968) );
  NANDN U2326 ( .A(A[156]), .B(n1970), .Z(n1969) );
  NANDN U2327 ( .A(n1970), .B(A[156]), .Z(n1967) );
  XOR U2328 ( .A(n1970), .B(n1971), .Z(DIFF[156]) );
  XOR U2329 ( .A(B[156]), .B(A[156]), .Z(n1971) );
  AND U2330 ( .A(n1972), .B(n1973), .Z(n1970) );
  NANDN U2331 ( .A(B[155]), .B(n1974), .Z(n1973) );
  NANDN U2332 ( .A(A[155]), .B(n1975), .Z(n1974) );
  NANDN U2333 ( .A(n1975), .B(A[155]), .Z(n1972) );
  XOR U2334 ( .A(n1975), .B(n1976), .Z(DIFF[155]) );
  XOR U2335 ( .A(B[155]), .B(A[155]), .Z(n1976) );
  AND U2336 ( .A(n1977), .B(n1978), .Z(n1975) );
  NANDN U2337 ( .A(B[154]), .B(n1979), .Z(n1978) );
  NANDN U2338 ( .A(A[154]), .B(n1980), .Z(n1979) );
  NANDN U2339 ( .A(n1980), .B(A[154]), .Z(n1977) );
  XOR U2340 ( .A(n1980), .B(n1981), .Z(DIFF[154]) );
  XOR U2341 ( .A(B[154]), .B(A[154]), .Z(n1981) );
  AND U2342 ( .A(n1982), .B(n1983), .Z(n1980) );
  NANDN U2343 ( .A(B[153]), .B(n1984), .Z(n1983) );
  NANDN U2344 ( .A(A[153]), .B(n1985), .Z(n1984) );
  NANDN U2345 ( .A(n1985), .B(A[153]), .Z(n1982) );
  XOR U2346 ( .A(n1985), .B(n1986), .Z(DIFF[153]) );
  XOR U2347 ( .A(B[153]), .B(A[153]), .Z(n1986) );
  AND U2348 ( .A(n1987), .B(n1988), .Z(n1985) );
  NANDN U2349 ( .A(B[152]), .B(n1989), .Z(n1988) );
  NANDN U2350 ( .A(A[152]), .B(n1990), .Z(n1989) );
  NANDN U2351 ( .A(n1990), .B(A[152]), .Z(n1987) );
  XOR U2352 ( .A(n1990), .B(n1991), .Z(DIFF[152]) );
  XOR U2353 ( .A(B[152]), .B(A[152]), .Z(n1991) );
  AND U2354 ( .A(n1992), .B(n1993), .Z(n1990) );
  NANDN U2355 ( .A(B[151]), .B(n1994), .Z(n1993) );
  NANDN U2356 ( .A(A[151]), .B(n1995), .Z(n1994) );
  NANDN U2357 ( .A(n1995), .B(A[151]), .Z(n1992) );
  XOR U2358 ( .A(n1995), .B(n1996), .Z(DIFF[151]) );
  XOR U2359 ( .A(B[151]), .B(A[151]), .Z(n1996) );
  AND U2360 ( .A(n1997), .B(n1998), .Z(n1995) );
  NANDN U2361 ( .A(B[150]), .B(n1999), .Z(n1998) );
  NANDN U2362 ( .A(A[150]), .B(n2000), .Z(n1999) );
  NANDN U2363 ( .A(n2000), .B(A[150]), .Z(n1997) );
  XOR U2364 ( .A(n2000), .B(n2001), .Z(DIFF[150]) );
  XOR U2365 ( .A(B[150]), .B(A[150]), .Z(n2001) );
  AND U2366 ( .A(n2002), .B(n2003), .Z(n2000) );
  NANDN U2367 ( .A(B[149]), .B(n2004), .Z(n2003) );
  NANDN U2368 ( .A(A[149]), .B(n2005), .Z(n2004) );
  NANDN U2369 ( .A(n2005), .B(A[149]), .Z(n2002) );
  XOR U2370 ( .A(n2006), .B(n2007), .Z(DIFF[14]) );
  XOR U2371 ( .A(B[14]), .B(A[14]), .Z(n2007) );
  XOR U2372 ( .A(n2005), .B(n2008), .Z(DIFF[149]) );
  XOR U2373 ( .A(B[149]), .B(A[149]), .Z(n2008) );
  AND U2374 ( .A(n2009), .B(n2010), .Z(n2005) );
  NANDN U2375 ( .A(B[148]), .B(n2011), .Z(n2010) );
  NANDN U2376 ( .A(A[148]), .B(n2012), .Z(n2011) );
  NANDN U2377 ( .A(n2012), .B(A[148]), .Z(n2009) );
  XOR U2378 ( .A(n2012), .B(n2013), .Z(DIFF[148]) );
  XOR U2379 ( .A(B[148]), .B(A[148]), .Z(n2013) );
  AND U2380 ( .A(n2014), .B(n2015), .Z(n2012) );
  NANDN U2381 ( .A(B[147]), .B(n2016), .Z(n2015) );
  NANDN U2382 ( .A(A[147]), .B(n2017), .Z(n2016) );
  NANDN U2383 ( .A(n2017), .B(A[147]), .Z(n2014) );
  XOR U2384 ( .A(n2017), .B(n2018), .Z(DIFF[147]) );
  XOR U2385 ( .A(B[147]), .B(A[147]), .Z(n2018) );
  AND U2386 ( .A(n2019), .B(n2020), .Z(n2017) );
  NANDN U2387 ( .A(B[146]), .B(n2021), .Z(n2020) );
  NANDN U2388 ( .A(A[146]), .B(n2022), .Z(n2021) );
  NANDN U2389 ( .A(n2022), .B(A[146]), .Z(n2019) );
  XOR U2390 ( .A(n2022), .B(n2023), .Z(DIFF[146]) );
  XOR U2391 ( .A(B[146]), .B(A[146]), .Z(n2023) );
  AND U2392 ( .A(n2024), .B(n2025), .Z(n2022) );
  NANDN U2393 ( .A(B[145]), .B(n2026), .Z(n2025) );
  NANDN U2394 ( .A(A[145]), .B(n2027), .Z(n2026) );
  NANDN U2395 ( .A(n2027), .B(A[145]), .Z(n2024) );
  XOR U2396 ( .A(n2027), .B(n2028), .Z(DIFF[145]) );
  XOR U2397 ( .A(B[145]), .B(A[145]), .Z(n2028) );
  AND U2398 ( .A(n2029), .B(n2030), .Z(n2027) );
  NANDN U2399 ( .A(B[144]), .B(n2031), .Z(n2030) );
  NANDN U2400 ( .A(A[144]), .B(n2032), .Z(n2031) );
  NANDN U2401 ( .A(n2032), .B(A[144]), .Z(n2029) );
  XOR U2402 ( .A(n2032), .B(n2033), .Z(DIFF[144]) );
  XOR U2403 ( .A(B[144]), .B(A[144]), .Z(n2033) );
  AND U2404 ( .A(n2034), .B(n2035), .Z(n2032) );
  NANDN U2405 ( .A(B[143]), .B(n2036), .Z(n2035) );
  NANDN U2406 ( .A(A[143]), .B(n2037), .Z(n2036) );
  NANDN U2407 ( .A(n2037), .B(A[143]), .Z(n2034) );
  XOR U2408 ( .A(n2037), .B(n2038), .Z(DIFF[143]) );
  XOR U2409 ( .A(B[143]), .B(A[143]), .Z(n2038) );
  AND U2410 ( .A(n2039), .B(n2040), .Z(n2037) );
  NANDN U2411 ( .A(B[142]), .B(n2041), .Z(n2040) );
  NANDN U2412 ( .A(A[142]), .B(n2042), .Z(n2041) );
  NANDN U2413 ( .A(n2042), .B(A[142]), .Z(n2039) );
  XOR U2414 ( .A(n2042), .B(n2043), .Z(DIFF[142]) );
  XOR U2415 ( .A(B[142]), .B(A[142]), .Z(n2043) );
  AND U2416 ( .A(n2044), .B(n2045), .Z(n2042) );
  NANDN U2417 ( .A(B[141]), .B(n2046), .Z(n2045) );
  NANDN U2418 ( .A(A[141]), .B(n2047), .Z(n2046) );
  NANDN U2419 ( .A(n2047), .B(A[141]), .Z(n2044) );
  XOR U2420 ( .A(n2047), .B(n2048), .Z(DIFF[141]) );
  XOR U2421 ( .A(B[141]), .B(A[141]), .Z(n2048) );
  AND U2422 ( .A(n2049), .B(n2050), .Z(n2047) );
  NANDN U2423 ( .A(B[140]), .B(n2051), .Z(n2050) );
  NANDN U2424 ( .A(A[140]), .B(n2052), .Z(n2051) );
  NANDN U2425 ( .A(n2052), .B(A[140]), .Z(n2049) );
  XOR U2426 ( .A(n2052), .B(n2053), .Z(DIFF[140]) );
  XOR U2427 ( .A(B[140]), .B(A[140]), .Z(n2053) );
  AND U2428 ( .A(n2054), .B(n2055), .Z(n2052) );
  NANDN U2429 ( .A(B[139]), .B(n2056), .Z(n2055) );
  NANDN U2430 ( .A(A[139]), .B(n2057), .Z(n2056) );
  NANDN U2431 ( .A(n2057), .B(A[139]), .Z(n2054) );
  XOR U2432 ( .A(n2058), .B(n2059), .Z(DIFF[13]) );
  XOR U2433 ( .A(B[13]), .B(A[13]), .Z(n2059) );
  XOR U2434 ( .A(n2057), .B(n2060), .Z(DIFF[139]) );
  XOR U2435 ( .A(B[139]), .B(A[139]), .Z(n2060) );
  AND U2436 ( .A(n2061), .B(n2062), .Z(n2057) );
  NANDN U2437 ( .A(B[138]), .B(n2063), .Z(n2062) );
  NANDN U2438 ( .A(A[138]), .B(n2064), .Z(n2063) );
  NANDN U2439 ( .A(n2064), .B(A[138]), .Z(n2061) );
  XOR U2440 ( .A(n2064), .B(n2065), .Z(DIFF[138]) );
  XOR U2441 ( .A(B[138]), .B(A[138]), .Z(n2065) );
  AND U2442 ( .A(n2066), .B(n2067), .Z(n2064) );
  NANDN U2443 ( .A(B[137]), .B(n2068), .Z(n2067) );
  NANDN U2444 ( .A(A[137]), .B(n2069), .Z(n2068) );
  NANDN U2445 ( .A(n2069), .B(A[137]), .Z(n2066) );
  XOR U2446 ( .A(n2069), .B(n2070), .Z(DIFF[137]) );
  XOR U2447 ( .A(B[137]), .B(A[137]), .Z(n2070) );
  AND U2448 ( .A(n2071), .B(n2072), .Z(n2069) );
  NANDN U2449 ( .A(B[136]), .B(n2073), .Z(n2072) );
  NANDN U2450 ( .A(A[136]), .B(n2074), .Z(n2073) );
  NANDN U2451 ( .A(n2074), .B(A[136]), .Z(n2071) );
  XOR U2452 ( .A(n2074), .B(n2075), .Z(DIFF[136]) );
  XOR U2453 ( .A(B[136]), .B(A[136]), .Z(n2075) );
  AND U2454 ( .A(n2076), .B(n2077), .Z(n2074) );
  NANDN U2455 ( .A(B[135]), .B(n2078), .Z(n2077) );
  NANDN U2456 ( .A(A[135]), .B(n2079), .Z(n2078) );
  NANDN U2457 ( .A(n2079), .B(A[135]), .Z(n2076) );
  XOR U2458 ( .A(n2079), .B(n2080), .Z(DIFF[135]) );
  XOR U2459 ( .A(B[135]), .B(A[135]), .Z(n2080) );
  AND U2460 ( .A(n2081), .B(n2082), .Z(n2079) );
  NANDN U2461 ( .A(B[134]), .B(n2083), .Z(n2082) );
  NANDN U2462 ( .A(A[134]), .B(n2084), .Z(n2083) );
  NANDN U2463 ( .A(n2084), .B(A[134]), .Z(n2081) );
  XOR U2464 ( .A(n2084), .B(n2085), .Z(DIFF[134]) );
  XOR U2465 ( .A(B[134]), .B(A[134]), .Z(n2085) );
  AND U2466 ( .A(n2086), .B(n2087), .Z(n2084) );
  NANDN U2467 ( .A(B[133]), .B(n2088), .Z(n2087) );
  NANDN U2468 ( .A(A[133]), .B(n2089), .Z(n2088) );
  NANDN U2469 ( .A(n2089), .B(A[133]), .Z(n2086) );
  XOR U2470 ( .A(n2089), .B(n2090), .Z(DIFF[133]) );
  XOR U2471 ( .A(B[133]), .B(A[133]), .Z(n2090) );
  AND U2472 ( .A(n2091), .B(n2092), .Z(n2089) );
  NANDN U2473 ( .A(B[132]), .B(n2093), .Z(n2092) );
  NANDN U2474 ( .A(A[132]), .B(n2094), .Z(n2093) );
  NANDN U2475 ( .A(n2094), .B(A[132]), .Z(n2091) );
  XOR U2476 ( .A(n2094), .B(n2095), .Z(DIFF[132]) );
  XOR U2477 ( .A(B[132]), .B(A[132]), .Z(n2095) );
  AND U2478 ( .A(n2096), .B(n2097), .Z(n2094) );
  NANDN U2479 ( .A(B[131]), .B(n2098), .Z(n2097) );
  NANDN U2480 ( .A(A[131]), .B(n2099), .Z(n2098) );
  NANDN U2481 ( .A(n2099), .B(A[131]), .Z(n2096) );
  XOR U2482 ( .A(n2099), .B(n2100), .Z(DIFF[131]) );
  XOR U2483 ( .A(B[131]), .B(A[131]), .Z(n2100) );
  AND U2484 ( .A(n2101), .B(n2102), .Z(n2099) );
  NANDN U2485 ( .A(B[130]), .B(n2103), .Z(n2102) );
  NANDN U2486 ( .A(A[130]), .B(n2104), .Z(n2103) );
  NANDN U2487 ( .A(n2104), .B(A[130]), .Z(n2101) );
  XOR U2488 ( .A(n2104), .B(n2105), .Z(DIFF[130]) );
  XOR U2489 ( .A(B[130]), .B(A[130]), .Z(n2105) );
  AND U2490 ( .A(n2106), .B(n2107), .Z(n2104) );
  NANDN U2491 ( .A(B[129]), .B(n2108), .Z(n2107) );
  NANDN U2492 ( .A(A[129]), .B(n2109), .Z(n2108) );
  NANDN U2493 ( .A(n2109), .B(A[129]), .Z(n2106) );
  XOR U2494 ( .A(n2110), .B(n2111), .Z(DIFF[12]) );
  XOR U2495 ( .A(B[12]), .B(A[12]), .Z(n2111) );
  XOR U2496 ( .A(n2109), .B(n2112), .Z(DIFF[129]) );
  XOR U2497 ( .A(B[129]), .B(A[129]), .Z(n2112) );
  AND U2498 ( .A(n2113), .B(n2114), .Z(n2109) );
  NANDN U2499 ( .A(B[128]), .B(n2115), .Z(n2114) );
  NANDN U2500 ( .A(A[128]), .B(n2116), .Z(n2115) );
  NANDN U2501 ( .A(n2116), .B(A[128]), .Z(n2113) );
  XOR U2502 ( .A(n2116), .B(n2117), .Z(DIFF[128]) );
  XOR U2503 ( .A(B[128]), .B(A[128]), .Z(n2117) );
  AND U2504 ( .A(n2118), .B(n2119), .Z(n2116) );
  NANDN U2505 ( .A(B[127]), .B(n2120), .Z(n2119) );
  NANDN U2506 ( .A(A[127]), .B(n2121), .Z(n2120) );
  NANDN U2507 ( .A(n2121), .B(A[127]), .Z(n2118) );
  XOR U2508 ( .A(n2121), .B(n2122), .Z(DIFF[127]) );
  XOR U2509 ( .A(B[127]), .B(A[127]), .Z(n2122) );
  AND U2510 ( .A(n2123), .B(n2124), .Z(n2121) );
  NANDN U2511 ( .A(B[126]), .B(n2125), .Z(n2124) );
  NANDN U2512 ( .A(A[126]), .B(n2126), .Z(n2125) );
  NANDN U2513 ( .A(n2126), .B(A[126]), .Z(n2123) );
  XOR U2514 ( .A(n2126), .B(n2127), .Z(DIFF[126]) );
  XOR U2515 ( .A(B[126]), .B(A[126]), .Z(n2127) );
  AND U2516 ( .A(n2128), .B(n2129), .Z(n2126) );
  NANDN U2517 ( .A(B[125]), .B(n2130), .Z(n2129) );
  NANDN U2518 ( .A(A[125]), .B(n2131), .Z(n2130) );
  NANDN U2519 ( .A(n2131), .B(A[125]), .Z(n2128) );
  XOR U2520 ( .A(n2131), .B(n2132), .Z(DIFF[125]) );
  XOR U2521 ( .A(B[125]), .B(A[125]), .Z(n2132) );
  AND U2522 ( .A(n2133), .B(n2134), .Z(n2131) );
  NANDN U2523 ( .A(B[124]), .B(n2135), .Z(n2134) );
  NANDN U2524 ( .A(A[124]), .B(n2136), .Z(n2135) );
  NANDN U2525 ( .A(n2136), .B(A[124]), .Z(n2133) );
  XOR U2526 ( .A(n2136), .B(n2137), .Z(DIFF[124]) );
  XOR U2527 ( .A(B[124]), .B(A[124]), .Z(n2137) );
  AND U2528 ( .A(n2138), .B(n2139), .Z(n2136) );
  NANDN U2529 ( .A(B[123]), .B(n2140), .Z(n2139) );
  NANDN U2530 ( .A(A[123]), .B(n2141), .Z(n2140) );
  NANDN U2531 ( .A(n2141), .B(A[123]), .Z(n2138) );
  XOR U2532 ( .A(n2141), .B(n2142), .Z(DIFF[123]) );
  XOR U2533 ( .A(B[123]), .B(A[123]), .Z(n2142) );
  AND U2534 ( .A(n2143), .B(n2144), .Z(n2141) );
  NANDN U2535 ( .A(B[122]), .B(n2145), .Z(n2144) );
  NANDN U2536 ( .A(A[122]), .B(n2146), .Z(n2145) );
  NANDN U2537 ( .A(n2146), .B(A[122]), .Z(n2143) );
  XOR U2538 ( .A(n2146), .B(n2147), .Z(DIFF[122]) );
  XOR U2539 ( .A(B[122]), .B(A[122]), .Z(n2147) );
  AND U2540 ( .A(n2148), .B(n2149), .Z(n2146) );
  NANDN U2541 ( .A(B[121]), .B(n2150), .Z(n2149) );
  NANDN U2542 ( .A(A[121]), .B(n2151), .Z(n2150) );
  NANDN U2543 ( .A(n2151), .B(A[121]), .Z(n2148) );
  XOR U2544 ( .A(n2151), .B(n2152), .Z(DIFF[121]) );
  XOR U2545 ( .A(B[121]), .B(A[121]), .Z(n2152) );
  AND U2546 ( .A(n2153), .B(n2154), .Z(n2151) );
  NANDN U2547 ( .A(B[120]), .B(n2155), .Z(n2154) );
  NANDN U2548 ( .A(A[120]), .B(n2156), .Z(n2155) );
  NANDN U2549 ( .A(n2156), .B(A[120]), .Z(n2153) );
  XOR U2550 ( .A(n2156), .B(n2157), .Z(DIFF[120]) );
  XOR U2551 ( .A(B[120]), .B(A[120]), .Z(n2157) );
  AND U2552 ( .A(n2158), .B(n2159), .Z(n2156) );
  NANDN U2553 ( .A(B[119]), .B(n2160), .Z(n2159) );
  NANDN U2554 ( .A(A[119]), .B(n2161), .Z(n2160) );
  NANDN U2555 ( .A(n2161), .B(A[119]), .Z(n2158) );
  XOR U2556 ( .A(n2162), .B(n2163), .Z(DIFF[11]) );
  XOR U2557 ( .A(B[11]), .B(A[11]), .Z(n2163) );
  XOR U2558 ( .A(n2161), .B(n2164), .Z(DIFF[119]) );
  XOR U2559 ( .A(B[119]), .B(A[119]), .Z(n2164) );
  AND U2560 ( .A(n2165), .B(n2166), .Z(n2161) );
  NANDN U2561 ( .A(B[118]), .B(n2167), .Z(n2166) );
  NANDN U2562 ( .A(A[118]), .B(n2168), .Z(n2167) );
  NANDN U2563 ( .A(n2168), .B(A[118]), .Z(n2165) );
  XOR U2564 ( .A(n2168), .B(n2169), .Z(DIFF[118]) );
  XOR U2565 ( .A(B[118]), .B(A[118]), .Z(n2169) );
  AND U2566 ( .A(n2170), .B(n2171), .Z(n2168) );
  NANDN U2567 ( .A(B[117]), .B(n2172), .Z(n2171) );
  NANDN U2568 ( .A(A[117]), .B(n2173), .Z(n2172) );
  NANDN U2569 ( .A(n2173), .B(A[117]), .Z(n2170) );
  XOR U2570 ( .A(n2173), .B(n2174), .Z(DIFF[117]) );
  XOR U2571 ( .A(B[117]), .B(A[117]), .Z(n2174) );
  AND U2572 ( .A(n2175), .B(n2176), .Z(n2173) );
  NANDN U2573 ( .A(B[116]), .B(n2177), .Z(n2176) );
  NANDN U2574 ( .A(A[116]), .B(n2178), .Z(n2177) );
  NANDN U2575 ( .A(n2178), .B(A[116]), .Z(n2175) );
  XOR U2576 ( .A(n2178), .B(n2179), .Z(DIFF[116]) );
  XOR U2577 ( .A(B[116]), .B(A[116]), .Z(n2179) );
  AND U2578 ( .A(n2180), .B(n2181), .Z(n2178) );
  NANDN U2579 ( .A(B[115]), .B(n2182), .Z(n2181) );
  NANDN U2580 ( .A(A[115]), .B(n2183), .Z(n2182) );
  NANDN U2581 ( .A(n2183), .B(A[115]), .Z(n2180) );
  XOR U2582 ( .A(n2183), .B(n2184), .Z(DIFF[115]) );
  XOR U2583 ( .A(B[115]), .B(A[115]), .Z(n2184) );
  AND U2584 ( .A(n2185), .B(n2186), .Z(n2183) );
  NANDN U2585 ( .A(B[114]), .B(n2187), .Z(n2186) );
  NANDN U2586 ( .A(A[114]), .B(n2188), .Z(n2187) );
  NANDN U2587 ( .A(n2188), .B(A[114]), .Z(n2185) );
  XOR U2588 ( .A(n2188), .B(n2189), .Z(DIFF[114]) );
  XOR U2589 ( .A(B[114]), .B(A[114]), .Z(n2189) );
  AND U2590 ( .A(n2190), .B(n2191), .Z(n2188) );
  NANDN U2591 ( .A(B[113]), .B(n2192), .Z(n2191) );
  NANDN U2592 ( .A(A[113]), .B(n2193), .Z(n2192) );
  NANDN U2593 ( .A(n2193), .B(A[113]), .Z(n2190) );
  XOR U2594 ( .A(n2193), .B(n2194), .Z(DIFF[113]) );
  XOR U2595 ( .A(B[113]), .B(A[113]), .Z(n2194) );
  AND U2596 ( .A(n2195), .B(n2196), .Z(n2193) );
  NANDN U2597 ( .A(B[112]), .B(n2197), .Z(n2196) );
  NANDN U2598 ( .A(A[112]), .B(n2198), .Z(n2197) );
  NANDN U2599 ( .A(n2198), .B(A[112]), .Z(n2195) );
  XOR U2600 ( .A(n2198), .B(n2199), .Z(DIFF[112]) );
  XOR U2601 ( .A(B[112]), .B(A[112]), .Z(n2199) );
  AND U2602 ( .A(n2200), .B(n2201), .Z(n2198) );
  NANDN U2603 ( .A(B[111]), .B(n2202), .Z(n2201) );
  NANDN U2604 ( .A(A[111]), .B(n2203), .Z(n2202) );
  NANDN U2605 ( .A(n2203), .B(A[111]), .Z(n2200) );
  XOR U2606 ( .A(n2203), .B(n2204), .Z(DIFF[111]) );
  XOR U2607 ( .A(B[111]), .B(A[111]), .Z(n2204) );
  AND U2608 ( .A(n2205), .B(n2206), .Z(n2203) );
  NANDN U2609 ( .A(B[110]), .B(n2207), .Z(n2206) );
  NANDN U2610 ( .A(A[110]), .B(n2208), .Z(n2207) );
  NANDN U2611 ( .A(n2208), .B(A[110]), .Z(n2205) );
  XOR U2612 ( .A(n2208), .B(n2209), .Z(DIFF[110]) );
  XOR U2613 ( .A(B[110]), .B(A[110]), .Z(n2209) );
  AND U2614 ( .A(n2210), .B(n2211), .Z(n2208) );
  NANDN U2615 ( .A(B[109]), .B(n2212), .Z(n2211) );
  NANDN U2616 ( .A(A[109]), .B(n2213), .Z(n2212) );
  NANDN U2617 ( .A(n2213), .B(A[109]), .Z(n2210) );
  XOR U2618 ( .A(n2214), .B(n2215), .Z(DIFF[10]) );
  XOR U2619 ( .A(B[10]), .B(A[10]), .Z(n2215) );
  XOR U2620 ( .A(n2213), .B(n2216), .Z(DIFF[109]) );
  XOR U2621 ( .A(B[109]), .B(A[109]), .Z(n2216) );
  AND U2622 ( .A(n2217), .B(n2218), .Z(n2213) );
  NANDN U2623 ( .A(B[108]), .B(n2219), .Z(n2218) );
  NANDN U2624 ( .A(A[108]), .B(n2220), .Z(n2219) );
  NANDN U2625 ( .A(n2220), .B(A[108]), .Z(n2217) );
  XOR U2626 ( .A(n2220), .B(n2221), .Z(DIFF[108]) );
  XOR U2627 ( .A(B[108]), .B(A[108]), .Z(n2221) );
  AND U2628 ( .A(n2222), .B(n2223), .Z(n2220) );
  NANDN U2629 ( .A(B[107]), .B(n2224), .Z(n2223) );
  NANDN U2630 ( .A(A[107]), .B(n2225), .Z(n2224) );
  NANDN U2631 ( .A(n2225), .B(A[107]), .Z(n2222) );
  XOR U2632 ( .A(n2225), .B(n2226), .Z(DIFF[107]) );
  XOR U2633 ( .A(B[107]), .B(A[107]), .Z(n2226) );
  AND U2634 ( .A(n2227), .B(n2228), .Z(n2225) );
  NANDN U2635 ( .A(B[106]), .B(n2229), .Z(n2228) );
  NANDN U2636 ( .A(A[106]), .B(n2230), .Z(n2229) );
  NANDN U2637 ( .A(n2230), .B(A[106]), .Z(n2227) );
  XOR U2638 ( .A(n2230), .B(n2231), .Z(DIFF[106]) );
  XOR U2639 ( .A(B[106]), .B(A[106]), .Z(n2231) );
  AND U2640 ( .A(n2232), .B(n2233), .Z(n2230) );
  NANDN U2641 ( .A(B[105]), .B(n2234), .Z(n2233) );
  NANDN U2642 ( .A(A[105]), .B(n2235), .Z(n2234) );
  NANDN U2643 ( .A(n2235), .B(A[105]), .Z(n2232) );
  XOR U2644 ( .A(n2235), .B(n2236), .Z(DIFF[105]) );
  XOR U2645 ( .A(B[105]), .B(A[105]), .Z(n2236) );
  AND U2646 ( .A(n2237), .B(n2238), .Z(n2235) );
  NANDN U2647 ( .A(B[104]), .B(n2239), .Z(n2238) );
  NANDN U2648 ( .A(A[104]), .B(n2240), .Z(n2239) );
  NANDN U2649 ( .A(n2240), .B(A[104]), .Z(n2237) );
  XOR U2650 ( .A(n2240), .B(n2241), .Z(DIFF[104]) );
  XOR U2651 ( .A(B[104]), .B(A[104]), .Z(n2241) );
  AND U2652 ( .A(n2242), .B(n2243), .Z(n2240) );
  NANDN U2653 ( .A(B[103]), .B(n2244), .Z(n2243) );
  NANDN U2654 ( .A(A[103]), .B(n2245), .Z(n2244) );
  NANDN U2655 ( .A(n2245), .B(A[103]), .Z(n2242) );
  XOR U2656 ( .A(n2245), .B(n2246), .Z(DIFF[103]) );
  XOR U2657 ( .A(B[103]), .B(A[103]), .Z(n2246) );
  AND U2658 ( .A(n2247), .B(n2248), .Z(n2245) );
  NANDN U2659 ( .A(B[102]), .B(n2249), .Z(n2248) );
  NANDN U2660 ( .A(A[102]), .B(n2250), .Z(n2249) );
  NANDN U2661 ( .A(n2250), .B(A[102]), .Z(n2247) );
  XOR U2662 ( .A(n2250), .B(n2251), .Z(DIFF[102]) );
  XOR U2663 ( .A(B[102]), .B(A[102]), .Z(n2251) );
  AND U2664 ( .A(n2252), .B(n2253), .Z(n2250) );
  NANDN U2665 ( .A(B[101]), .B(n2254), .Z(n2253) );
  NANDN U2666 ( .A(A[101]), .B(n2255), .Z(n2254) );
  NANDN U2667 ( .A(n2255), .B(A[101]), .Z(n2252) );
  XOR U2668 ( .A(n2255), .B(n2256), .Z(DIFF[101]) );
  XOR U2669 ( .A(B[101]), .B(A[101]), .Z(n2256) );
  AND U2670 ( .A(n2257), .B(n2258), .Z(n2255) );
  NANDN U2671 ( .A(B[100]), .B(n2259), .Z(n2258) );
  NANDN U2672 ( .A(A[100]), .B(n2260), .Z(n2259) );
  NANDN U2673 ( .A(n2260), .B(A[100]), .Z(n2257) );
  XOR U2674 ( .A(n2260), .B(n2261), .Z(DIFF[100]) );
  XOR U2675 ( .A(B[100]), .B(A[100]), .Z(n2261) );
  AND U2676 ( .A(n2262), .B(n2263), .Z(n2260) );
  NANDN U2677 ( .A(B[99]), .B(n2264), .Z(n2263) );
  OR U2678 ( .A(n5), .B(A[99]), .Z(n2264) );
  NAND U2679 ( .A(A[99]), .B(n5), .Z(n2262) );
  NAND U2680 ( .A(n2265), .B(n2266), .Z(n5) );
  NANDN U2681 ( .A(B[98]), .B(n2267), .Z(n2266) );
  NANDN U2682 ( .A(A[98]), .B(n7), .Z(n2267) );
  NANDN U2683 ( .A(n7), .B(A[98]), .Z(n2265) );
  AND U2684 ( .A(n2268), .B(n2269), .Z(n7) );
  NANDN U2685 ( .A(B[97]), .B(n2270), .Z(n2269) );
  NANDN U2686 ( .A(A[97]), .B(n9), .Z(n2270) );
  NANDN U2687 ( .A(n9), .B(A[97]), .Z(n2268) );
  AND U2688 ( .A(n2271), .B(n2272), .Z(n9) );
  NANDN U2689 ( .A(B[96]), .B(n2273), .Z(n2272) );
  NANDN U2690 ( .A(A[96]), .B(n11), .Z(n2273) );
  NANDN U2691 ( .A(n11), .B(A[96]), .Z(n2271) );
  AND U2692 ( .A(n2274), .B(n2275), .Z(n11) );
  NANDN U2693 ( .A(B[95]), .B(n2276), .Z(n2275) );
  NANDN U2694 ( .A(A[95]), .B(n13), .Z(n2276) );
  NANDN U2695 ( .A(n13), .B(A[95]), .Z(n2274) );
  AND U2696 ( .A(n2277), .B(n2278), .Z(n13) );
  NANDN U2697 ( .A(B[94]), .B(n2279), .Z(n2278) );
  NANDN U2698 ( .A(A[94]), .B(n15), .Z(n2279) );
  NANDN U2699 ( .A(n15), .B(A[94]), .Z(n2277) );
  AND U2700 ( .A(n2280), .B(n2281), .Z(n15) );
  NANDN U2701 ( .A(B[93]), .B(n2282), .Z(n2281) );
  NANDN U2702 ( .A(A[93]), .B(n17), .Z(n2282) );
  NANDN U2703 ( .A(n17), .B(A[93]), .Z(n2280) );
  AND U2704 ( .A(n2283), .B(n2284), .Z(n17) );
  NANDN U2705 ( .A(B[92]), .B(n2285), .Z(n2284) );
  NANDN U2706 ( .A(A[92]), .B(n19), .Z(n2285) );
  NANDN U2707 ( .A(n19), .B(A[92]), .Z(n2283) );
  AND U2708 ( .A(n2286), .B(n2287), .Z(n19) );
  NANDN U2709 ( .A(B[91]), .B(n2288), .Z(n2287) );
  NANDN U2710 ( .A(A[91]), .B(n21), .Z(n2288) );
  NANDN U2711 ( .A(n21), .B(A[91]), .Z(n2286) );
  AND U2712 ( .A(n2289), .B(n2290), .Z(n21) );
  NANDN U2713 ( .A(B[90]), .B(n2291), .Z(n2290) );
  NANDN U2714 ( .A(A[90]), .B(n23), .Z(n2291) );
  NANDN U2715 ( .A(n23), .B(A[90]), .Z(n2289) );
  AND U2716 ( .A(n2292), .B(n2293), .Z(n23) );
  NANDN U2717 ( .A(B[89]), .B(n2294), .Z(n2293) );
  NANDN U2718 ( .A(A[89]), .B(n27), .Z(n2294) );
  NANDN U2719 ( .A(n27), .B(A[89]), .Z(n2292) );
  AND U2720 ( .A(n2295), .B(n2296), .Z(n27) );
  NANDN U2721 ( .A(B[88]), .B(n2297), .Z(n2296) );
  NANDN U2722 ( .A(A[88]), .B(n29), .Z(n2297) );
  NANDN U2723 ( .A(n29), .B(A[88]), .Z(n2295) );
  AND U2724 ( .A(n2298), .B(n2299), .Z(n29) );
  NANDN U2725 ( .A(B[87]), .B(n2300), .Z(n2299) );
  NANDN U2726 ( .A(A[87]), .B(n31), .Z(n2300) );
  NANDN U2727 ( .A(n31), .B(A[87]), .Z(n2298) );
  AND U2728 ( .A(n2301), .B(n2302), .Z(n31) );
  NANDN U2729 ( .A(B[86]), .B(n2303), .Z(n2302) );
  NANDN U2730 ( .A(A[86]), .B(n33), .Z(n2303) );
  NANDN U2731 ( .A(n33), .B(A[86]), .Z(n2301) );
  AND U2732 ( .A(n2304), .B(n2305), .Z(n33) );
  NANDN U2733 ( .A(B[85]), .B(n2306), .Z(n2305) );
  NANDN U2734 ( .A(A[85]), .B(n35), .Z(n2306) );
  NANDN U2735 ( .A(n35), .B(A[85]), .Z(n2304) );
  AND U2736 ( .A(n2307), .B(n2308), .Z(n35) );
  NANDN U2737 ( .A(B[84]), .B(n2309), .Z(n2308) );
  NANDN U2738 ( .A(A[84]), .B(n37), .Z(n2309) );
  NANDN U2739 ( .A(n37), .B(A[84]), .Z(n2307) );
  AND U2740 ( .A(n2310), .B(n2311), .Z(n37) );
  NANDN U2741 ( .A(B[83]), .B(n2312), .Z(n2311) );
  NANDN U2742 ( .A(A[83]), .B(n39), .Z(n2312) );
  NANDN U2743 ( .A(n39), .B(A[83]), .Z(n2310) );
  AND U2744 ( .A(n2313), .B(n2314), .Z(n39) );
  NANDN U2745 ( .A(B[82]), .B(n2315), .Z(n2314) );
  NANDN U2746 ( .A(A[82]), .B(n41), .Z(n2315) );
  NANDN U2747 ( .A(n41), .B(A[82]), .Z(n2313) );
  AND U2748 ( .A(n2316), .B(n2317), .Z(n41) );
  NANDN U2749 ( .A(B[81]), .B(n2318), .Z(n2317) );
  NANDN U2750 ( .A(A[81]), .B(n43), .Z(n2318) );
  NANDN U2751 ( .A(n43), .B(A[81]), .Z(n2316) );
  AND U2752 ( .A(n2319), .B(n2320), .Z(n43) );
  NANDN U2753 ( .A(B[80]), .B(n2321), .Z(n2320) );
  NANDN U2754 ( .A(A[80]), .B(n45), .Z(n2321) );
  NANDN U2755 ( .A(n45), .B(A[80]), .Z(n2319) );
  AND U2756 ( .A(n2322), .B(n2323), .Z(n45) );
  NANDN U2757 ( .A(B[79]), .B(n2324), .Z(n2323) );
  NANDN U2758 ( .A(A[79]), .B(n49), .Z(n2324) );
  NANDN U2759 ( .A(n49), .B(A[79]), .Z(n2322) );
  AND U2760 ( .A(n2325), .B(n2326), .Z(n49) );
  NANDN U2761 ( .A(B[78]), .B(n2327), .Z(n2326) );
  NANDN U2762 ( .A(A[78]), .B(n51), .Z(n2327) );
  NANDN U2763 ( .A(n51), .B(A[78]), .Z(n2325) );
  AND U2764 ( .A(n2328), .B(n2329), .Z(n51) );
  NANDN U2765 ( .A(B[77]), .B(n2330), .Z(n2329) );
  NANDN U2766 ( .A(A[77]), .B(n53), .Z(n2330) );
  NANDN U2767 ( .A(n53), .B(A[77]), .Z(n2328) );
  AND U2768 ( .A(n2331), .B(n2332), .Z(n53) );
  NANDN U2769 ( .A(B[76]), .B(n2333), .Z(n2332) );
  NANDN U2770 ( .A(A[76]), .B(n55), .Z(n2333) );
  NANDN U2771 ( .A(n55), .B(A[76]), .Z(n2331) );
  AND U2772 ( .A(n2334), .B(n2335), .Z(n55) );
  NANDN U2773 ( .A(B[75]), .B(n2336), .Z(n2335) );
  NANDN U2774 ( .A(A[75]), .B(n57), .Z(n2336) );
  NANDN U2775 ( .A(n57), .B(A[75]), .Z(n2334) );
  AND U2776 ( .A(n2337), .B(n2338), .Z(n57) );
  NANDN U2777 ( .A(B[74]), .B(n2339), .Z(n2338) );
  NANDN U2778 ( .A(A[74]), .B(n59), .Z(n2339) );
  NANDN U2779 ( .A(n59), .B(A[74]), .Z(n2337) );
  AND U2780 ( .A(n2340), .B(n2341), .Z(n59) );
  NANDN U2781 ( .A(B[73]), .B(n2342), .Z(n2341) );
  NANDN U2782 ( .A(A[73]), .B(n61), .Z(n2342) );
  NANDN U2783 ( .A(n61), .B(A[73]), .Z(n2340) );
  AND U2784 ( .A(n2343), .B(n2344), .Z(n61) );
  NANDN U2785 ( .A(B[72]), .B(n2345), .Z(n2344) );
  NANDN U2786 ( .A(A[72]), .B(n63), .Z(n2345) );
  NANDN U2787 ( .A(n63), .B(A[72]), .Z(n2343) );
  AND U2788 ( .A(n2346), .B(n2347), .Z(n63) );
  NANDN U2789 ( .A(B[71]), .B(n2348), .Z(n2347) );
  NANDN U2790 ( .A(A[71]), .B(n65), .Z(n2348) );
  NANDN U2791 ( .A(n65), .B(A[71]), .Z(n2346) );
  AND U2792 ( .A(n2349), .B(n2350), .Z(n65) );
  NANDN U2793 ( .A(B[70]), .B(n2351), .Z(n2350) );
  NANDN U2794 ( .A(A[70]), .B(n67), .Z(n2351) );
  NANDN U2795 ( .A(n67), .B(A[70]), .Z(n2349) );
  AND U2796 ( .A(n2352), .B(n2353), .Z(n67) );
  NANDN U2797 ( .A(B[69]), .B(n2354), .Z(n2353) );
  NANDN U2798 ( .A(A[69]), .B(n71), .Z(n2354) );
  NANDN U2799 ( .A(n71), .B(A[69]), .Z(n2352) );
  AND U2800 ( .A(n2355), .B(n2356), .Z(n71) );
  NANDN U2801 ( .A(B[68]), .B(n2357), .Z(n2356) );
  NANDN U2802 ( .A(A[68]), .B(n73), .Z(n2357) );
  NANDN U2803 ( .A(n73), .B(A[68]), .Z(n2355) );
  AND U2804 ( .A(n2358), .B(n2359), .Z(n73) );
  NANDN U2805 ( .A(B[67]), .B(n2360), .Z(n2359) );
  NANDN U2806 ( .A(A[67]), .B(n75), .Z(n2360) );
  NANDN U2807 ( .A(n75), .B(A[67]), .Z(n2358) );
  AND U2808 ( .A(n2361), .B(n2362), .Z(n75) );
  NANDN U2809 ( .A(B[66]), .B(n2363), .Z(n2362) );
  NANDN U2810 ( .A(A[66]), .B(n77), .Z(n2363) );
  NANDN U2811 ( .A(n77), .B(A[66]), .Z(n2361) );
  AND U2812 ( .A(n2364), .B(n2365), .Z(n77) );
  NANDN U2813 ( .A(B[65]), .B(n2366), .Z(n2365) );
  NANDN U2814 ( .A(A[65]), .B(n79), .Z(n2366) );
  NANDN U2815 ( .A(n79), .B(A[65]), .Z(n2364) );
  AND U2816 ( .A(n2367), .B(n2368), .Z(n79) );
  NANDN U2817 ( .A(B[64]), .B(n2369), .Z(n2368) );
  NANDN U2818 ( .A(A[64]), .B(n81), .Z(n2369) );
  NANDN U2819 ( .A(n81), .B(A[64]), .Z(n2367) );
  AND U2820 ( .A(n2370), .B(n2371), .Z(n81) );
  NANDN U2821 ( .A(B[63]), .B(n2372), .Z(n2371) );
  NANDN U2822 ( .A(A[63]), .B(n83), .Z(n2372) );
  NANDN U2823 ( .A(n83), .B(A[63]), .Z(n2370) );
  AND U2824 ( .A(n2373), .B(n2374), .Z(n83) );
  NANDN U2825 ( .A(B[62]), .B(n2375), .Z(n2374) );
  NANDN U2826 ( .A(A[62]), .B(n85), .Z(n2375) );
  NANDN U2827 ( .A(n85), .B(A[62]), .Z(n2373) );
  AND U2828 ( .A(n2376), .B(n2377), .Z(n85) );
  NANDN U2829 ( .A(B[61]), .B(n2378), .Z(n2377) );
  NANDN U2830 ( .A(A[61]), .B(n87), .Z(n2378) );
  NANDN U2831 ( .A(n87), .B(A[61]), .Z(n2376) );
  AND U2832 ( .A(n2379), .B(n2380), .Z(n87) );
  NANDN U2833 ( .A(B[60]), .B(n2381), .Z(n2380) );
  NANDN U2834 ( .A(A[60]), .B(n89), .Z(n2381) );
  NANDN U2835 ( .A(n89), .B(A[60]), .Z(n2379) );
  AND U2836 ( .A(n2382), .B(n2383), .Z(n89) );
  NANDN U2837 ( .A(B[59]), .B(n2384), .Z(n2383) );
  NANDN U2838 ( .A(A[59]), .B(n93), .Z(n2384) );
  NANDN U2839 ( .A(n93), .B(A[59]), .Z(n2382) );
  AND U2840 ( .A(n2385), .B(n2386), .Z(n93) );
  NANDN U2841 ( .A(B[58]), .B(n2387), .Z(n2386) );
  NANDN U2842 ( .A(A[58]), .B(n95), .Z(n2387) );
  NANDN U2843 ( .A(n95), .B(A[58]), .Z(n2385) );
  AND U2844 ( .A(n2388), .B(n2389), .Z(n95) );
  NANDN U2845 ( .A(B[57]), .B(n2390), .Z(n2389) );
  NANDN U2846 ( .A(A[57]), .B(n97), .Z(n2390) );
  NANDN U2847 ( .A(n97), .B(A[57]), .Z(n2388) );
  AND U2848 ( .A(n2391), .B(n2392), .Z(n97) );
  NANDN U2849 ( .A(B[56]), .B(n2393), .Z(n2392) );
  NANDN U2850 ( .A(A[56]), .B(n99), .Z(n2393) );
  NANDN U2851 ( .A(n99), .B(A[56]), .Z(n2391) );
  AND U2852 ( .A(n2394), .B(n2395), .Z(n99) );
  NANDN U2853 ( .A(B[55]), .B(n2396), .Z(n2395) );
  NANDN U2854 ( .A(A[55]), .B(n101), .Z(n2396) );
  NANDN U2855 ( .A(n101), .B(A[55]), .Z(n2394) );
  AND U2856 ( .A(n2397), .B(n2398), .Z(n101) );
  NANDN U2857 ( .A(B[54]), .B(n2399), .Z(n2398) );
  NANDN U2858 ( .A(A[54]), .B(n103), .Z(n2399) );
  NANDN U2859 ( .A(n103), .B(A[54]), .Z(n2397) );
  AND U2860 ( .A(n2400), .B(n2401), .Z(n103) );
  NANDN U2861 ( .A(B[53]), .B(n2402), .Z(n2401) );
  NANDN U2862 ( .A(A[53]), .B(n105), .Z(n2402) );
  NANDN U2863 ( .A(n105), .B(A[53]), .Z(n2400) );
  AND U2864 ( .A(n2403), .B(n2404), .Z(n105) );
  NANDN U2865 ( .A(B[52]), .B(n2405), .Z(n2404) );
  NANDN U2866 ( .A(A[52]), .B(n107), .Z(n2405) );
  NANDN U2867 ( .A(n107), .B(A[52]), .Z(n2403) );
  AND U2868 ( .A(n2406), .B(n2407), .Z(n107) );
  NANDN U2869 ( .A(B[51]), .B(n2408), .Z(n2407) );
  NANDN U2870 ( .A(A[51]), .B(n109), .Z(n2408) );
  NANDN U2871 ( .A(n109), .B(A[51]), .Z(n2406) );
  AND U2872 ( .A(n2409), .B(n2410), .Z(n109) );
  NANDN U2873 ( .A(B[50]), .B(n2411), .Z(n2410) );
  NANDN U2874 ( .A(A[50]), .B(n127), .Z(n2411) );
  NANDN U2875 ( .A(n127), .B(A[50]), .Z(n2409) );
  AND U2876 ( .A(n2412), .B(n2413), .Z(n127) );
  NANDN U2877 ( .A(B[49]), .B(n2414), .Z(n2413) );
  NANDN U2878 ( .A(A[49]), .B(n181), .Z(n2414) );
  NANDN U2879 ( .A(n181), .B(A[49]), .Z(n2412) );
  AND U2880 ( .A(n2415), .B(n2416), .Z(n181) );
  NANDN U2881 ( .A(B[48]), .B(n2417), .Z(n2416) );
  NANDN U2882 ( .A(A[48]), .B(n233), .Z(n2417) );
  NANDN U2883 ( .A(n233), .B(A[48]), .Z(n2415) );
  AND U2884 ( .A(n2418), .B(n2419), .Z(n233) );
  NANDN U2885 ( .A(B[47]), .B(n2420), .Z(n2419) );
  NANDN U2886 ( .A(A[47]), .B(n285), .Z(n2420) );
  NANDN U2887 ( .A(n285), .B(A[47]), .Z(n2418) );
  AND U2888 ( .A(n2421), .B(n2422), .Z(n285) );
  NANDN U2889 ( .A(B[46]), .B(n2423), .Z(n2422) );
  NANDN U2890 ( .A(A[46]), .B(n337), .Z(n2423) );
  NANDN U2891 ( .A(n337), .B(A[46]), .Z(n2421) );
  AND U2892 ( .A(n2424), .B(n2425), .Z(n337) );
  NANDN U2893 ( .A(B[45]), .B(n2426), .Z(n2425) );
  NANDN U2894 ( .A(A[45]), .B(n389), .Z(n2426) );
  NANDN U2895 ( .A(n389), .B(A[45]), .Z(n2424) );
  AND U2896 ( .A(n2427), .B(n2428), .Z(n389) );
  NANDN U2897 ( .A(B[44]), .B(n2429), .Z(n2428) );
  NANDN U2898 ( .A(A[44]), .B(n441), .Z(n2429) );
  NANDN U2899 ( .A(n441), .B(A[44]), .Z(n2427) );
  AND U2900 ( .A(n2430), .B(n2431), .Z(n441) );
  NANDN U2901 ( .A(B[43]), .B(n2432), .Z(n2431) );
  NANDN U2902 ( .A(A[43]), .B(n493), .Z(n2432) );
  NANDN U2903 ( .A(n493), .B(A[43]), .Z(n2430) );
  AND U2904 ( .A(n2433), .B(n2434), .Z(n493) );
  NANDN U2905 ( .A(B[42]), .B(n2435), .Z(n2434) );
  NANDN U2906 ( .A(A[42]), .B(n545), .Z(n2435) );
  NANDN U2907 ( .A(n545), .B(A[42]), .Z(n2433) );
  AND U2908 ( .A(n2436), .B(n2437), .Z(n545) );
  NANDN U2909 ( .A(B[41]), .B(n2438), .Z(n2437) );
  NANDN U2910 ( .A(A[41]), .B(n597), .Z(n2438) );
  NANDN U2911 ( .A(n597), .B(A[41]), .Z(n2436) );
  AND U2912 ( .A(n2439), .B(n2440), .Z(n597) );
  NANDN U2913 ( .A(B[40]), .B(n2441), .Z(n2440) );
  NANDN U2914 ( .A(A[40]), .B(n649), .Z(n2441) );
  NANDN U2915 ( .A(n649), .B(A[40]), .Z(n2439) );
  AND U2916 ( .A(n2442), .B(n2443), .Z(n649) );
  NANDN U2917 ( .A(B[39]), .B(n2444), .Z(n2443) );
  NANDN U2918 ( .A(A[39]), .B(n703), .Z(n2444) );
  NANDN U2919 ( .A(n703), .B(A[39]), .Z(n2442) );
  AND U2920 ( .A(n2445), .B(n2446), .Z(n703) );
  NANDN U2921 ( .A(B[38]), .B(n2447), .Z(n2446) );
  NANDN U2922 ( .A(A[38]), .B(n755), .Z(n2447) );
  NANDN U2923 ( .A(n755), .B(A[38]), .Z(n2445) );
  AND U2924 ( .A(n2448), .B(n2449), .Z(n755) );
  NANDN U2925 ( .A(B[37]), .B(n2450), .Z(n2449) );
  NANDN U2926 ( .A(A[37]), .B(n807), .Z(n2450) );
  NANDN U2927 ( .A(n807), .B(A[37]), .Z(n2448) );
  AND U2928 ( .A(n2451), .B(n2452), .Z(n807) );
  NANDN U2929 ( .A(B[36]), .B(n2453), .Z(n2452) );
  NANDN U2930 ( .A(A[36]), .B(n859), .Z(n2453) );
  NANDN U2931 ( .A(n859), .B(A[36]), .Z(n2451) );
  AND U2932 ( .A(n2454), .B(n2455), .Z(n859) );
  NANDN U2933 ( .A(B[35]), .B(n2456), .Z(n2455) );
  NANDN U2934 ( .A(A[35]), .B(n911), .Z(n2456) );
  NANDN U2935 ( .A(n911), .B(A[35]), .Z(n2454) );
  AND U2936 ( .A(n2457), .B(n2458), .Z(n911) );
  NANDN U2937 ( .A(B[34]), .B(n2459), .Z(n2458) );
  NANDN U2938 ( .A(A[34]), .B(n963), .Z(n2459) );
  NANDN U2939 ( .A(n963), .B(A[34]), .Z(n2457) );
  AND U2940 ( .A(n2460), .B(n2461), .Z(n963) );
  NANDN U2941 ( .A(B[33]), .B(n2462), .Z(n2461) );
  NANDN U2942 ( .A(A[33]), .B(n1015), .Z(n2462) );
  NANDN U2943 ( .A(n1015), .B(A[33]), .Z(n2460) );
  AND U2944 ( .A(n2463), .B(n2464), .Z(n1015) );
  NANDN U2945 ( .A(B[32]), .B(n2465), .Z(n2464) );
  NANDN U2946 ( .A(A[32]), .B(n1067), .Z(n2465) );
  NANDN U2947 ( .A(n1067), .B(A[32]), .Z(n2463) );
  AND U2948 ( .A(n2466), .B(n2467), .Z(n1067) );
  NANDN U2949 ( .A(B[31]), .B(n2468), .Z(n2467) );
  NANDN U2950 ( .A(A[31]), .B(n1119), .Z(n2468) );
  NANDN U2951 ( .A(n1119), .B(A[31]), .Z(n2466) );
  AND U2952 ( .A(n2469), .B(n2470), .Z(n1119) );
  NANDN U2953 ( .A(B[30]), .B(n2471), .Z(n2470) );
  NANDN U2954 ( .A(A[30]), .B(n1171), .Z(n2471) );
  NANDN U2955 ( .A(n1171), .B(A[30]), .Z(n2469) );
  AND U2956 ( .A(n2472), .B(n2473), .Z(n1171) );
  NANDN U2957 ( .A(B[29]), .B(n2474), .Z(n2473) );
  NANDN U2958 ( .A(A[29]), .B(n1225), .Z(n2474) );
  NANDN U2959 ( .A(n1225), .B(A[29]), .Z(n2472) );
  AND U2960 ( .A(n2475), .B(n2476), .Z(n1225) );
  NANDN U2961 ( .A(B[28]), .B(n2477), .Z(n2476) );
  NANDN U2962 ( .A(A[28]), .B(n1277), .Z(n2477) );
  NANDN U2963 ( .A(n1277), .B(A[28]), .Z(n2475) );
  AND U2964 ( .A(n2478), .B(n2479), .Z(n1277) );
  NANDN U2965 ( .A(B[27]), .B(n2480), .Z(n2479) );
  NANDN U2966 ( .A(A[27]), .B(n1329), .Z(n2480) );
  NANDN U2967 ( .A(n1329), .B(A[27]), .Z(n2478) );
  AND U2968 ( .A(n2481), .B(n2482), .Z(n1329) );
  NANDN U2969 ( .A(B[26]), .B(n2483), .Z(n2482) );
  NANDN U2970 ( .A(A[26]), .B(n1381), .Z(n2483) );
  NANDN U2971 ( .A(n1381), .B(A[26]), .Z(n2481) );
  AND U2972 ( .A(n2484), .B(n2485), .Z(n1381) );
  NANDN U2973 ( .A(B[25]), .B(n2486), .Z(n2485) );
  NANDN U2974 ( .A(A[25]), .B(n1433), .Z(n2486) );
  NANDN U2975 ( .A(n1433), .B(A[25]), .Z(n2484) );
  AND U2976 ( .A(n2487), .B(n2488), .Z(n1433) );
  NANDN U2977 ( .A(B[24]), .B(n2489), .Z(n2488) );
  NANDN U2978 ( .A(A[24]), .B(n1485), .Z(n2489) );
  NANDN U2979 ( .A(n1485), .B(A[24]), .Z(n2487) );
  AND U2980 ( .A(n2490), .B(n2491), .Z(n1485) );
  NANDN U2981 ( .A(B[23]), .B(n2492), .Z(n2491) );
  NANDN U2982 ( .A(A[23]), .B(n1537), .Z(n2492) );
  NANDN U2983 ( .A(n1537), .B(A[23]), .Z(n2490) );
  AND U2984 ( .A(n2493), .B(n2494), .Z(n1537) );
  NANDN U2985 ( .A(B[22]), .B(n2495), .Z(n2494) );
  NANDN U2986 ( .A(A[22]), .B(n1589), .Z(n2495) );
  NANDN U2987 ( .A(n1589), .B(A[22]), .Z(n2493) );
  AND U2988 ( .A(n2496), .B(n2497), .Z(n1589) );
  NANDN U2989 ( .A(B[21]), .B(n2498), .Z(n2497) );
  NANDN U2990 ( .A(A[21]), .B(n1641), .Z(n2498) );
  NANDN U2991 ( .A(n1641), .B(A[21]), .Z(n2496) );
  AND U2992 ( .A(n2499), .B(n2500), .Z(n1641) );
  NANDN U2993 ( .A(B[20]), .B(n2501), .Z(n2500) );
  NANDN U2994 ( .A(A[20]), .B(n1693), .Z(n2501) );
  NANDN U2995 ( .A(n1693), .B(A[20]), .Z(n2499) );
  AND U2996 ( .A(n2502), .B(n2503), .Z(n1693) );
  NANDN U2997 ( .A(B[19]), .B(n2504), .Z(n2503) );
  NANDN U2998 ( .A(A[19]), .B(n1746), .Z(n2504) );
  NANDN U2999 ( .A(n1746), .B(A[19]), .Z(n2502) );
  AND U3000 ( .A(n2505), .B(n2506), .Z(n1746) );
  NANDN U3001 ( .A(B[18]), .B(n2507), .Z(n2506) );
  NANDN U3002 ( .A(A[18]), .B(n1798), .Z(n2507) );
  NANDN U3003 ( .A(n1798), .B(A[18]), .Z(n2505) );
  AND U3004 ( .A(n2508), .B(n2509), .Z(n1798) );
  NANDN U3005 ( .A(B[17]), .B(n2510), .Z(n2509) );
  NANDN U3006 ( .A(A[17]), .B(n1850), .Z(n2510) );
  NANDN U3007 ( .A(n1850), .B(A[17]), .Z(n2508) );
  AND U3008 ( .A(n2511), .B(n2512), .Z(n1850) );
  NANDN U3009 ( .A(B[16]), .B(n2513), .Z(n2512) );
  NANDN U3010 ( .A(A[16]), .B(n1902), .Z(n2513) );
  NANDN U3011 ( .A(n1902), .B(A[16]), .Z(n2511) );
  AND U3012 ( .A(n2514), .B(n2515), .Z(n1902) );
  NANDN U3013 ( .A(B[15]), .B(n2516), .Z(n2515) );
  NANDN U3014 ( .A(A[15]), .B(n1954), .Z(n2516) );
  NANDN U3015 ( .A(n1954), .B(A[15]), .Z(n2514) );
  AND U3016 ( .A(n2517), .B(n2518), .Z(n1954) );
  NANDN U3017 ( .A(B[14]), .B(n2519), .Z(n2518) );
  NANDN U3018 ( .A(A[14]), .B(n2006), .Z(n2519) );
  NANDN U3019 ( .A(n2006), .B(A[14]), .Z(n2517) );
  AND U3020 ( .A(n2520), .B(n2521), .Z(n2006) );
  NANDN U3021 ( .A(B[13]), .B(n2522), .Z(n2521) );
  NANDN U3022 ( .A(A[13]), .B(n2058), .Z(n2522) );
  NANDN U3023 ( .A(n2058), .B(A[13]), .Z(n2520) );
  AND U3024 ( .A(n2523), .B(n2524), .Z(n2058) );
  NANDN U3025 ( .A(B[12]), .B(n2525), .Z(n2524) );
  NANDN U3026 ( .A(A[12]), .B(n2110), .Z(n2525) );
  NANDN U3027 ( .A(n2110), .B(A[12]), .Z(n2523) );
  AND U3028 ( .A(n2526), .B(n2527), .Z(n2110) );
  NANDN U3029 ( .A(B[11]), .B(n2528), .Z(n2527) );
  NANDN U3030 ( .A(A[11]), .B(n2162), .Z(n2528) );
  NANDN U3031 ( .A(n2162), .B(A[11]), .Z(n2526) );
  AND U3032 ( .A(n2529), .B(n2530), .Z(n2162) );
  NANDN U3033 ( .A(B[10]), .B(n2531), .Z(n2530) );
  NANDN U3034 ( .A(A[10]), .B(n2214), .Z(n2531) );
  NANDN U3035 ( .A(n2214), .B(A[10]), .Z(n2529) );
  AND U3036 ( .A(n2532), .B(n2533), .Z(n2214) );
  NANDN U3037 ( .A(B[9]), .B(n2534), .Z(n2533) );
  OR U3038 ( .A(n3), .B(A[9]), .Z(n2534) );
  NAND U3039 ( .A(A[9]), .B(n3), .Z(n2532) );
  NAND U3040 ( .A(n2535), .B(n2536), .Z(n3) );
  NANDN U3041 ( .A(B[8]), .B(n2537), .Z(n2536) );
  NANDN U3042 ( .A(A[8]), .B(n25), .Z(n2537) );
  NANDN U3043 ( .A(n25), .B(A[8]), .Z(n2535) );
  AND U3044 ( .A(n2538), .B(n2539), .Z(n25) );
  NANDN U3045 ( .A(B[7]), .B(n2540), .Z(n2539) );
  NANDN U3046 ( .A(A[7]), .B(n47), .Z(n2540) );
  NANDN U3047 ( .A(n47), .B(A[7]), .Z(n2538) );
  AND U3048 ( .A(n2541), .B(n2542), .Z(n47) );
  NANDN U3049 ( .A(B[6]), .B(n2543), .Z(n2542) );
  NANDN U3050 ( .A(A[6]), .B(n69), .Z(n2543) );
  NANDN U3051 ( .A(n69), .B(A[6]), .Z(n2541) );
  AND U3052 ( .A(n2544), .B(n2545), .Z(n69) );
  NANDN U3053 ( .A(B[5]), .B(n2546), .Z(n2545) );
  NANDN U3054 ( .A(A[5]), .B(n91), .Z(n2546) );
  NANDN U3055 ( .A(n91), .B(A[5]), .Z(n2544) );
  AND U3056 ( .A(n2547), .B(n2548), .Z(n91) );
  NANDN U3057 ( .A(B[4]), .B(n2549), .Z(n2548) );
  NANDN U3058 ( .A(A[4]), .B(n179), .Z(n2549) );
  NANDN U3059 ( .A(n179), .B(A[4]), .Z(n2547) );
  AND U3060 ( .A(n2550), .B(n2551), .Z(n179) );
  NANDN U3061 ( .A(B[3]), .B(n2552), .Z(n2551) );
  NANDN U3062 ( .A(A[3]), .B(n701), .Z(n2552) );
  NANDN U3063 ( .A(n701), .B(A[3]), .Z(n2550) );
  AND U3064 ( .A(n2553), .B(n2554), .Z(n701) );
  NANDN U3065 ( .A(B[2]), .B(n2555), .Z(n2554) );
  NANDN U3066 ( .A(A[2]), .B(n1223), .Z(n2555) );
  NANDN U3067 ( .A(n1223), .B(A[2]), .Z(n2553) );
  AND U3068 ( .A(n2556), .B(n2557), .Z(n1223) );
  NANDN U3069 ( .A(B[1]), .B(n2558), .Z(n2557) );
  NAND U3070 ( .A(n2), .B(n1), .Z(n2558) );
  NAND U3071 ( .A(A[1]), .B(n2559), .Z(n2556) );
  NAND U3072 ( .A(n2559), .B(n2560), .Z(DIFF[0]) );
  NANDN U3073 ( .A(B[0]), .B(A[0]), .Z(n2560) );
  NANDN U3074 ( .A(A[0]), .B(B[0]), .Z(n2559) );
endmodule


module modmult_step_N512_DW01_cmp2_1 ( A, B, LEQ, TC, LT_LE, GE_GT );
  input [513:0] A;
  input [513:0] B;
  input LEQ, TC;
  output LT_LE, GE_GT;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046;

  NAND U1 ( .A(n1), .B(n2), .Z(LT_LE) );
  NOR U2 ( .A(B[513]), .B(B[512]), .Z(n2) );
  AND U3 ( .A(n3), .B(n4), .Z(n1) );
  NAND U4 ( .A(n5), .B(n6), .Z(n4) );
  NANDN U5 ( .A(B[511]), .B(A[511]), .Z(n6) );
  NAND U6 ( .A(n7), .B(n8), .Z(n5) );
  NANDN U7 ( .A(A[510]), .B(B[510]), .Z(n8) );
  NAND U8 ( .A(n9), .B(n10), .Z(n7) );
  NANDN U9 ( .A(B[510]), .B(A[510]), .Z(n10) );
  AND U10 ( .A(n11), .B(n12), .Z(n9) );
  NAND U11 ( .A(n13), .B(n14), .Z(n12) );
  NANDN U12 ( .A(A[509]), .B(B[509]), .Z(n14) );
  AND U13 ( .A(n15), .B(n16), .Z(n13) );
  NANDN U14 ( .A(A[508]), .B(B[508]), .Z(n16) );
  NAND U15 ( .A(n17), .B(n18), .Z(n15) );
  NANDN U16 ( .A(B[508]), .B(A[508]), .Z(n18) );
  AND U17 ( .A(n19), .B(n20), .Z(n17) );
  NAND U18 ( .A(n21), .B(n22), .Z(n20) );
  NANDN U19 ( .A(A[507]), .B(B[507]), .Z(n22) );
  AND U20 ( .A(n23), .B(n24), .Z(n21) );
  NANDN U21 ( .A(A[506]), .B(B[506]), .Z(n24) );
  NAND U22 ( .A(n25), .B(n26), .Z(n23) );
  NANDN U23 ( .A(B[506]), .B(A[506]), .Z(n26) );
  AND U24 ( .A(n27), .B(n28), .Z(n25) );
  NAND U25 ( .A(n29), .B(n30), .Z(n28) );
  NANDN U26 ( .A(A[505]), .B(B[505]), .Z(n30) );
  AND U27 ( .A(n31), .B(n32), .Z(n29) );
  NANDN U28 ( .A(A[504]), .B(B[504]), .Z(n32) );
  NAND U29 ( .A(n33), .B(n34), .Z(n31) );
  NANDN U30 ( .A(B[504]), .B(A[504]), .Z(n34) );
  AND U31 ( .A(n35), .B(n36), .Z(n33) );
  NAND U32 ( .A(n37), .B(n38), .Z(n36) );
  NANDN U33 ( .A(A[503]), .B(B[503]), .Z(n38) );
  AND U34 ( .A(n39), .B(n40), .Z(n37) );
  NANDN U35 ( .A(A[502]), .B(B[502]), .Z(n40) );
  NAND U36 ( .A(n41), .B(n42), .Z(n39) );
  NANDN U37 ( .A(B[502]), .B(A[502]), .Z(n42) );
  AND U38 ( .A(n43), .B(n44), .Z(n41) );
  NAND U39 ( .A(n45), .B(n46), .Z(n44) );
  NANDN U40 ( .A(A[501]), .B(B[501]), .Z(n46) );
  AND U41 ( .A(n47), .B(n48), .Z(n45) );
  NANDN U42 ( .A(A[500]), .B(B[500]), .Z(n48) );
  NAND U43 ( .A(n49), .B(n50), .Z(n47) );
  NANDN U44 ( .A(B[500]), .B(A[500]), .Z(n50) );
  AND U45 ( .A(n51), .B(n52), .Z(n49) );
  NAND U46 ( .A(n53), .B(n54), .Z(n52) );
  NANDN U47 ( .A(A[499]), .B(B[499]), .Z(n54) );
  AND U48 ( .A(n55), .B(n56), .Z(n53) );
  NANDN U49 ( .A(A[498]), .B(B[498]), .Z(n56) );
  NAND U50 ( .A(n57), .B(n58), .Z(n55) );
  NANDN U51 ( .A(B[498]), .B(A[498]), .Z(n58) );
  AND U52 ( .A(n59), .B(n60), .Z(n57) );
  NAND U53 ( .A(n61), .B(n62), .Z(n60) );
  NANDN U54 ( .A(A[497]), .B(B[497]), .Z(n62) );
  AND U55 ( .A(n63), .B(n64), .Z(n61) );
  NANDN U56 ( .A(A[496]), .B(B[496]), .Z(n64) );
  NAND U57 ( .A(n65), .B(n66), .Z(n63) );
  NANDN U58 ( .A(B[496]), .B(A[496]), .Z(n66) );
  AND U59 ( .A(n67), .B(n68), .Z(n65) );
  NAND U60 ( .A(n69), .B(n70), .Z(n68) );
  NANDN U61 ( .A(A[495]), .B(B[495]), .Z(n70) );
  AND U62 ( .A(n71), .B(n72), .Z(n69) );
  NANDN U63 ( .A(A[494]), .B(B[494]), .Z(n72) );
  NAND U64 ( .A(n73), .B(n74), .Z(n71) );
  NANDN U65 ( .A(B[494]), .B(A[494]), .Z(n74) );
  AND U66 ( .A(n75), .B(n76), .Z(n73) );
  NAND U67 ( .A(n77), .B(n78), .Z(n76) );
  NANDN U68 ( .A(A[493]), .B(B[493]), .Z(n78) );
  AND U69 ( .A(n79), .B(n80), .Z(n77) );
  NANDN U70 ( .A(A[492]), .B(B[492]), .Z(n80) );
  NAND U71 ( .A(n81), .B(n82), .Z(n79) );
  NANDN U72 ( .A(B[492]), .B(A[492]), .Z(n82) );
  AND U73 ( .A(n83), .B(n84), .Z(n81) );
  NAND U74 ( .A(n85), .B(n86), .Z(n84) );
  NANDN U75 ( .A(A[491]), .B(B[491]), .Z(n86) );
  AND U76 ( .A(n87), .B(n88), .Z(n85) );
  NANDN U77 ( .A(A[490]), .B(B[490]), .Z(n88) );
  NAND U78 ( .A(n89), .B(n90), .Z(n87) );
  NANDN U79 ( .A(B[490]), .B(A[490]), .Z(n90) );
  AND U80 ( .A(n91), .B(n92), .Z(n89) );
  NAND U81 ( .A(n93), .B(n94), .Z(n92) );
  NANDN U82 ( .A(A[489]), .B(B[489]), .Z(n94) );
  AND U83 ( .A(n95), .B(n96), .Z(n93) );
  NANDN U84 ( .A(A[488]), .B(B[488]), .Z(n96) );
  NAND U85 ( .A(n97), .B(n98), .Z(n95) );
  NANDN U86 ( .A(B[488]), .B(A[488]), .Z(n98) );
  AND U87 ( .A(n99), .B(n100), .Z(n97) );
  NAND U88 ( .A(n101), .B(n102), .Z(n100) );
  NANDN U89 ( .A(A[487]), .B(B[487]), .Z(n102) );
  AND U90 ( .A(n103), .B(n104), .Z(n101) );
  NANDN U91 ( .A(A[486]), .B(B[486]), .Z(n104) );
  NAND U92 ( .A(n105), .B(n106), .Z(n103) );
  NANDN U93 ( .A(B[486]), .B(A[486]), .Z(n106) );
  AND U94 ( .A(n107), .B(n108), .Z(n105) );
  NAND U95 ( .A(n109), .B(n110), .Z(n108) );
  NANDN U96 ( .A(A[485]), .B(B[485]), .Z(n110) );
  AND U97 ( .A(n111), .B(n112), .Z(n109) );
  NANDN U98 ( .A(A[484]), .B(B[484]), .Z(n112) );
  NAND U99 ( .A(n113), .B(n114), .Z(n111) );
  NANDN U100 ( .A(B[484]), .B(A[484]), .Z(n114) );
  AND U101 ( .A(n115), .B(n116), .Z(n113) );
  NAND U102 ( .A(n117), .B(n118), .Z(n116) );
  NANDN U103 ( .A(A[483]), .B(B[483]), .Z(n118) );
  AND U104 ( .A(n119), .B(n120), .Z(n117) );
  NANDN U105 ( .A(A[482]), .B(B[482]), .Z(n120) );
  NAND U106 ( .A(n121), .B(n122), .Z(n119) );
  NANDN U107 ( .A(B[482]), .B(A[482]), .Z(n122) );
  AND U108 ( .A(n123), .B(n124), .Z(n121) );
  NAND U109 ( .A(n125), .B(n126), .Z(n124) );
  NANDN U110 ( .A(A[481]), .B(B[481]), .Z(n126) );
  AND U111 ( .A(n127), .B(n128), .Z(n125) );
  NANDN U112 ( .A(A[480]), .B(B[480]), .Z(n128) );
  NAND U113 ( .A(n129), .B(n130), .Z(n127) );
  NANDN U114 ( .A(B[480]), .B(A[480]), .Z(n130) );
  AND U115 ( .A(n131), .B(n132), .Z(n129) );
  NAND U116 ( .A(n133), .B(n134), .Z(n132) );
  NANDN U117 ( .A(A[479]), .B(B[479]), .Z(n134) );
  AND U118 ( .A(n135), .B(n136), .Z(n133) );
  NANDN U119 ( .A(A[478]), .B(B[478]), .Z(n136) );
  NAND U120 ( .A(n137), .B(n138), .Z(n135) );
  NANDN U121 ( .A(B[478]), .B(A[478]), .Z(n138) );
  AND U122 ( .A(n139), .B(n140), .Z(n137) );
  NAND U123 ( .A(n141), .B(n142), .Z(n140) );
  NANDN U124 ( .A(A[477]), .B(B[477]), .Z(n142) );
  AND U125 ( .A(n143), .B(n144), .Z(n141) );
  NANDN U126 ( .A(A[476]), .B(B[476]), .Z(n144) );
  NAND U127 ( .A(n145), .B(n146), .Z(n143) );
  NANDN U128 ( .A(B[476]), .B(A[476]), .Z(n146) );
  AND U129 ( .A(n147), .B(n148), .Z(n145) );
  NAND U130 ( .A(n149), .B(n150), .Z(n148) );
  NANDN U131 ( .A(A[475]), .B(B[475]), .Z(n150) );
  AND U132 ( .A(n151), .B(n152), .Z(n149) );
  NANDN U133 ( .A(A[474]), .B(B[474]), .Z(n152) );
  NAND U134 ( .A(n153), .B(n154), .Z(n151) );
  NANDN U135 ( .A(B[474]), .B(A[474]), .Z(n154) );
  AND U136 ( .A(n155), .B(n156), .Z(n153) );
  NAND U137 ( .A(n157), .B(n158), .Z(n156) );
  NANDN U138 ( .A(A[473]), .B(B[473]), .Z(n158) );
  AND U139 ( .A(n159), .B(n160), .Z(n157) );
  NANDN U140 ( .A(A[472]), .B(B[472]), .Z(n160) );
  NAND U141 ( .A(n161), .B(n162), .Z(n159) );
  NANDN U142 ( .A(B[472]), .B(A[472]), .Z(n162) );
  AND U143 ( .A(n163), .B(n164), .Z(n161) );
  NAND U144 ( .A(n165), .B(n166), .Z(n164) );
  NANDN U145 ( .A(A[471]), .B(B[471]), .Z(n166) );
  AND U146 ( .A(n167), .B(n168), .Z(n165) );
  NANDN U147 ( .A(A[470]), .B(B[470]), .Z(n168) );
  NAND U148 ( .A(n169), .B(n170), .Z(n167) );
  NANDN U149 ( .A(B[470]), .B(A[470]), .Z(n170) );
  AND U150 ( .A(n171), .B(n172), .Z(n169) );
  NAND U151 ( .A(n173), .B(n174), .Z(n172) );
  NANDN U152 ( .A(A[469]), .B(B[469]), .Z(n174) );
  AND U153 ( .A(n175), .B(n176), .Z(n173) );
  NANDN U154 ( .A(A[468]), .B(B[468]), .Z(n176) );
  NAND U155 ( .A(n177), .B(n178), .Z(n175) );
  NANDN U156 ( .A(B[468]), .B(A[468]), .Z(n178) );
  AND U157 ( .A(n179), .B(n180), .Z(n177) );
  NAND U158 ( .A(n181), .B(n182), .Z(n180) );
  NANDN U159 ( .A(A[467]), .B(B[467]), .Z(n182) );
  AND U160 ( .A(n183), .B(n184), .Z(n181) );
  NANDN U161 ( .A(A[466]), .B(B[466]), .Z(n184) );
  NAND U162 ( .A(n185), .B(n186), .Z(n183) );
  NANDN U163 ( .A(B[466]), .B(A[466]), .Z(n186) );
  AND U164 ( .A(n187), .B(n188), .Z(n185) );
  NAND U165 ( .A(n189), .B(n190), .Z(n188) );
  NANDN U166 ( .A(A[465]), .B(B[465]), .Z(n190) );
  AND U167 ( .A(n191), .B(n192), .Z(n189) );
  NANDN U168 ( .A(A[464]), .B(B[464]), .Z(n192) );
  NAND U169 ( .A(n193), .B(n194), .Z(n191) );
  NANDN U170 ( .A(B[464]), .B(A[464]), .Z(n194) );
  AND U171 ( .A(n195), .B(n196), .Z(n193) );
  NAND U172 ( .A(n197), .B(n198), .Z(n196) );
  NANDN U173 ( .A(A[463]), .B(B[463]), .Z(n198) );
  AND U174 ( .A(n199), .B(n200), .Z(n197) );
  NANDN U175 ( .A(A[462]), .B(B[462]), .Z(n200) );
  NAND U176 ( .A(n201), .B(n202), .Z(n199) );
  NANDN U177 ( .A(B[462]), .B(A[462]), .Z(n202) );
  AND U178 ( .A(n203), .B(n204), .Z(n201) );
  NAND U179 ( .A(n205), .B(n206), .Z(n204) );
  NANDN U180 ( .A(A[461]), .B(B[461]), .Z(n206) );
  AND U181 ( .A(n207), .B(n208), .Z(n205) );
  NANDN U182 ( .A(A[460]), .B(B[460]), .Z(n208) );
  NAND U183 ( .A(n209), .B(n210), .Z(n207) );
  NANDN U184 ( .A(B[460]), .B(A[460]), .Z(n210) );
  AND U185 ( .A(n211), .B(n212), .Z(n209) );
  NAND U186 ( .A(n213), .B(n214), .Z(n212) );
  NANDN U187 ( .A(A[459]), .B(B[459]), .Z(n214) );
  AND U188 ( .A(n215), .B(n216), .Z(n213) );
  NANDN U189 ( .A(A[458]), .B(B[458]), .Z(n216) );
  NAND U190 ( .A(n217), .B(n218), .Z(n215) );
  NANDN U191 ( .A(B[458]), .B(A[458]), .Z(n218) );
  AND U192 ( .A(n219), .B(n220), .Z(n217) );
  NAND U193 ( .A(n221), .B(n222), .Z(n220) );
  NANDN U194 ( .A(A[457]), .B(B[457]), .Z(n222) );
  AND U195 ( .A(n223), .B(n224), .Z(n221) );
  NANDN U196 ( .A(A[456]), .B(B[456]), .Z(n224) );
  NAND U197 ( .A(n225), .B(n226), .Z(n223) );
  NANDN U198 ( .A(B[456]), .B(A[456]), .Z(n226) );
  AND U199 ( .A(n227), .B(n228), .Z(n225) );
  NAND U200 ( .A(n229), .B(n230), .Z(n228) );
  NANDN U201 ( .A(A[455]), .B(B[455]), .Z(n230) );
  AND U202 ( .A(n231), .B(n232), .Z(n229) );
  NANDN U203 ( .A(A[454]), .B(B[454]), .Z(n232) );
  NAND U204 ( .A(n233), .B(n234), .Z(n231) );
  NANDN U205 ( .A(B[454]), .B(A[454]), .Z(n234) );
  AND U206 ( .A(n235), .B(n236), .Z(n233) );
  NAND U207 ( .A(n237), .B(n238), .Z(n236) );
  NANDN U208 ( .A(A[453]), .B(B[453]), .Z(n238) );
  AND U209 ( .A(n239), .B(n240), .Z(n237) );
  NANDN U210 ( .A(A[452]), .B(B[452]), .Z(n240) );
  NAND U211 ( .A(n241), .B(n242), .Z(n239) );
  NANDN U212 ( .A(B[452]), .B(A[452]), .Z(n242) );
  AND U213 ( .A(n243), .B(n244), .Z(n241) );
  NAND U214 ( .A(n245), .B(n246), .Z(n244) );
  NANDN U215 ( .A(A[451]), .B(B[451]), .Z(n246) );
  AND U216 ( .A(n247), .B(n248), .Z(n245) );
  NANDN U217 ( .A(A[450]), .B(B[450]), .Z(n248) );
  NAND U218 ( .A(n249), .B(n250), .Z(n247) );
  NANDN U219 ( .A(B[450]), .B(A[450]), .Z(n250) );
  AND U220 ( .A(n251), .B(n252), .Z(n249) );
  NAND U221 ( .A(n253), .B(n254), .Z(n252) );
  NANDN U222 ( .A(A[449]), .B(B[449]), .Z(n254) );
  AND U223 ( .A(n255), .B(n256), .Z(n253) );
  NANDN U224 ( .A(A[448]), .B(B[448]), .Z(n256) );
  NAND U225 ( .A(n257), .B(n258), .Z(n255) );
  NANDN U226 ( .A(B[448]), .B(A[448]), .Z(n258) );
  AND U227 ( .A(n259), .B(n260), .Z(n257) );
  NAND U228 ( .A(n261), .B(n262), .Z(n260) );
  NANDN U229 ( .A(A[447]), .B(B[447]), .Z(n262) );
  AND U230 ( .A(n263), .B(n264), .Z(n261) );
  NANDN U231 ( .A(A[446]), .B(B[446]), .Z(n264) );
  NAND U232 ( .A(n265), .B(n266), .Z(n263) );
  NANDN U233 ( .A(B[446]), .B(A[446]), .Z(n266) );
  AND U234 ( .A(n267), .B(n268), .Z(n265) );
  NAND U235 ( .A(n269), .B(n270), .Z(n268) );
  NANDN U236 ( .A(A[445]), .B(B[445]), .Z(n270) );
  AND U237 ( .A(n271), .B(n272), .Z(n269) );
  NANDN U238 ( .A(A[444]), .B(B[444]), .Z(n272) );
  NAND U239 ( .A(n273), .B(n274), .Z(n271) );
  NANDN U240 ( .A(B[444]), .B(A[444]), .Z(n274) );
  AND U241 ( .A(n275), .B(n276), .Z(n273) );
  NAND U242 ( .A(n277), .B(n278), .Z(n276) );
  NANDN U243 ( .A(A[443]), .B(B[443]), .Z(n278) );
  AND U244 ( .A(n279), .B(n280), .Z(n277) );
  NANDN U245 ( .A(A[442]), .B(B[442]), .Z(n280) );
  NAND U246 ( .A(n281), .B(n282), .Z(n279) );
  NANDN U247 ( .A(B[442]), .B(A[442]), .Z(n282) );
  AND U248 ( .A(n283), .B(n284), .Z(n281) );
  NAND U249 ( .A(n285), .B(n286), .Z(n284) );
  NANDN U250 ( .A(A[441]), .B(B[441]), .Z(n286) );
  AND U251 ( .A(n287), .B(n288), .Z(n285) );
  NANDN U252 ( .A(A[440]), .B(B[440]), .Z(n288) );
  NAND U253 ( .A(n289), .B(n290), .Z(n287) );
  NANDN U254 ( .A(B[440]), .B(A[440]), .Z(n290) );
  AND U255 ( .A(n291), .B(n292), .Z(n289) );
  NAND U256 ( .A(n293), .B(n294), .Z(n292) );
  NANDN U257 ( .A(A[439]), .B(B[439]), .Z(n294) );
  AND U258 ( .A(n295), .B(n296), .Z(n293) );
  NANDN U259 ( .A(A[438]), .B(B[438]), .Z(n296) );
  NAND U260 ( .A(n297), .B(n298), .Z(n295) );
  NANDN U261 ( .A(B[438]), .B(A[438]), .Z(n298) );
  AND U262 ( .A(n299), .B(n300), .Z(n297) );
  NAND U263 ( .A(n301), .B(n302), .Z(n300) );
  NANDN U264 ( .A(A[437]), .B(B[437]), .Z(n302) );
  AND U265 ( .A(n303), .B(n304), .Z(n301) );
  NANDN U266 ( .A(A[436]), .B(B[436]), .Z(n304) );
  NAND U267 ( .A(n305), .B(n306), .Z(n303) );
  NANDN U268 ( .A(B[436]), .B(A[436]), .Z(n306) );
  AND U269 ( .A(n307), .B(n308), .Z(n305) );
  NAND U270 ( .A(n309), .B(n310), .Z(n308) );
  NANDN U271 ( .A(A[435]), .B(B[435]), .Z(n310) );
  AND U272 ( .A(n311), .B(n312), .Z(n309) );
  NANDN U273 ( .A(A[434]), .B(B[434]), .Z(n312) );
  NAND U274 ( .A(n313), .B(n314), .Z(n311) );
  NANDN U275 ( .A(B[434]), .B(A[434]), .Z(n314) );
  AND U276 ( .A(n315), .B(n316), .Z(n313) );
  NAND U277 ( .A(n317), .B(n318), .Z(n316) );
  NANDN U278 ( .A(A[433]), .B(B[433]), .Z(n318) );
  AND U279 ( .A(n319), .B(n320), .Z(n317) );
  NANDN U280 ( .A(A[432]), .B(B[432]), .Z(n320) );
  NAND U281 ( .A(n321), .B(n322), .Z(n319) );
  NANDN U282 ( .A(B[432]), .B(A[432]), .Z(n322) );
  AND U283 ( .A(n323), .B(n324), .Z(n321) );
  NAND U284 ( .A(n325), .B(n326), .Z(n324) );
  NANDN U285 ( .A(A[431]), .B(B[431]), .Z(n326) );
  AND U286 ( .A(n327), .B(n328), .Z(n325) );
  NANDN U287 ( .A(A[430]), .B(B[430]), .Z(n328) );
  NAND U288 ( .A(n329), .B(n330), .Z(n327) );
  NANDN U289 ( .A(B[430]), .B(A[430]), .Z(n330) );
  AND U290 ( .A(n331), .B(n332), .Z(n329) );
  NAND U291 ( .A(n333), .B(n334), .Z(n332) );
  NANDN U292 ( .A(A[429]), .B(B[429]), .Z(n334) );
  AND U293 ( .A(n335), .B(n336), .Z(n333) );
  NANDN U294 ( .A(A[428]), .B(B[428]), .Z(n336) );
  NAND U295 ( .A(n337), .B(n338), .Z(n335) );
  NANDN U296 ( .A(B[428]), .B(A[428]), .Z(n338) );
  AND U297 ( .A(n339), .B(n340), .Z(n337) );
  NAND U298 ( .A(n341), .B(n342), .Z(n340) );
  NANDN U299 ( .A(A[427]), .B(B[427]), .Z(n342) );
  AND U300 ( .A(n343), .B(n344), .Z(n341) );
  NANDN U301 ( .A(A[426]), .B(B[426]), .Z(n344) );
  NAND U302 ( .A(n345), .B(n346), .Z(n343) );
  NANDN U303 ( .A(B[426]), .B(A[426]), .Z(n346) );
  AND U304 ( .A(n347), .B(n348), .Z(n345) );
  NAND U305 ( .A(n349), .B(n350), .Z(n348) );
  NANDN U306 ( .A(A[425]), .B(B[425]), .Z(n350) );
  AND U307 ( .A(n351), .B(n352), .Z(n349) );
  NANDN U308 ( .A(A[424]), .B(B[424]), .Z(n352) );
  NAND U309 ( .A(n353), .B(n354), .Z(n351) );
  NANDN U310 ( .A(B[424]), .B(A[424]), .Z(n354) );
  AND U311 ( .A(n355), .B(n356), .Z(n353) );
  NAND U312 ( .A(n357), .B(n358), .Z(n356) );
  NANDN U313 ( .A(A[423]), .B(B[423]), .Z(n358) );
  AND U314 ( .A(n359), .B(n360), .Z(n357) );
  NANDN U315 ( .A(A[422]), .B(B[422]), .Z(n360) );
  NAND U316 ( .A(n361), .B(n362), .Z(n359) );
  NANDN U317 ( .A(B[422]), .B(A[422]), .Z(n362) );
  AND U318 ( .A(n363), .B(n364), .Z(n361) );
  NAND U319 ( .A(n365), .B(n366), .Z(n364) );
  NANDN U320 ( .A(A[421]), .B(B[421]), .Z(n366) );
  AND U321 ( .A(n367), .B(n368), .Z(n365) );
  NANDN U322 ( .A(A[420]), .B(B[420]), .Z(n368) );
  NAND U323 ( .A(n369), .B(n370), .Z(n367) );
  NANDN U324 ( .A(B[420]), .B(A[420]), .Z(n370) );
  AND U325 ( .A(n371), .B(n372), .Z(n369) );
  NAND U326 ( .A(n373), .B(n374), .Z(n372) );
  NANDN U327 ( .A(A[419]), .B(B[419]), .Z(n374) );
  AND U328 ( .A(n375), .B(n376), .Z(n373) );
  NANDN U329 ( .A(A[418]), .B(B[418]), .Z(n376) );
  NAND U330 ( .A(n377), .B(n378), .Z(n375) );
  NANDN U331 ( .A(B[418]), .B(A[418]), .Z(n378) );
  AND U332 ( .A(n379), .B(n380), .Z(n377) );
  NAND U333 ( .A(n381), .B(n382), .Z(n380) );
  NANDN U334 ( .A(A[417]), .B(B[417]), .Z(n382) );
  AND U335 ( .A(n383), .B(n384), .Z(n381) );
  NANDN U336 ( .A(A[416]), .B(B[416]), .Z(n384) );
  NAND U337 ( .A(n385), .B(n386), .Z(n383) );
  NANDN U338 ( .A(B[416]), .B(A[416]), .Z(n386) );
  AND U339 ( .A(n387), .B(n388), .Z(n385) );
  NAND U340 ( .A(n389), .B(n390), .Z(n388) );
  NANDN U341 ( .A(A[415]), .B(B[415]), .Z(n390) );
  AND U342 ( .A(n391), .B(n392), .Z(n389) );
  NANDN U343 ( .A(A[414]), .B(B[414]), .Z(n392) );
  NAND U344 ( .A(n393), .B(n394), .Z(n391) );
  NANDN U345 ( .A(B[414]), .B(A[414]), .Z(n394) );
  AND U346 ( .A(n395), .B(n396), .Z(n393) );
  NAND U347 ( .A(n397), .B(n398), .Z(n396) );
  NANDN U348 ( .A(A[413]), .B(B[413]), .Z(n398) );
  AND U349 ( .A(n399), .B(n400), .Z(n397) );
  NANDN U350 ( .A(A[412]), .B(B[412]), .Z(n400) );
  NAND U351 ( .A(n401), .B(n402), .Z(n399) );
  NANDN U352 ( .A(B[412]), .B(A[412]), .Z(n402) );
  AND U353 ( .A(n403), .B(n404), .Z(n401) );
  NAND U354 ( .A(n405), .B(n406), .Z(n404) );
  NANDN U355 ( .A(A[411]), .B(B[411]), .Z(n406) );
  AND U356 ( .A(n407), .B(n408), .Z(n405) );
  NANDN U357 ( .A(A[410]), .B(B[410]), .Z(n408) );
  NAND U358 ( .A(n409), .B(n410), .Z(n407) );
  NANDN U359 ( .A(B[410]), .B(A[410]), .Z(n410) );
  AND U360 ( .A(n411), .B(n412), .Z(n409) );
  NAND U361 ( .A(n413), .B(n414), .Z(n412) );
  NANDN U362 ( .A(A[409]), .B(B[409]), .Z(n414) );
  AND U363 ( .A(n415), .B(n416), .Z(n413) );
  NANDN U364 ( .A(A[408]), .B(B[408]), .Z(n416) );
  NAND U365 ( .A(n417), .B(n418), .Z(n415) );
  NANDN U366 ( .A(B[408]), .B(A[408]), .Z(n418) );
  AND U367 ( .A(n419), .B(n420), .Z(n417) );
  NAND U368 ( .A(n421), .B(n422), .Z(n420) );
  NANDN U369 ( .A(A[407]), .B(B[407]), .Z(n422) );
  AND U370 ( .A(n423), .B(n424), .Z(n421) );
  NANDN U371 ( .A(A[406]), .B(B[406]), .Z(n424) );
  NAND U372 ( .A(n425), .B(n426), .Z(n423) );
  NANDN U373 ( .A(B[406]), .B(A[406]), .Z(n426) );
  AND U374 ( .A(n427), .B(n428), .Z(n425) );
  NAND U375 ( .A(n429), .B(n430), .Z(n428) );
  NANDN U376 ( .A(A[405]), .B(B[405]), .Z(n430) );
  AND U377 ( .A(n431), .B(n432), .Z(n429) );
  NANDN U378 ( .A(A[404]), .B(B[404]), .Z(n432) );
  NAND U379 ( .A(n433), .B(n434), .Z(n431) );
  NANDN U380 ( .A(B[404]), .B(A[404]), .Z(n434) );
  AND U381 ( .A(n435), .B(n436), .Z(n433) );
  NAND U382 ( .A(n437), .B(n438), .Z(n436) );
  NANDN U383 ( .A(A[403]), .B(B[403]), .Z(n438) );
  AND U384 ( .A(n439), .B(n440), .Z(n437) );
  NANDN U385 ( .A(A[402]), .B(B[402]), .Z(n440) );
  NAND U386 ( .A(n441), .B(n442), .Z(n439) );
  NANDN U387 ( .A(B[402]), .B(A[402]), .Z(n442) );
  AND U388 ( .A(n443), .B(n444), .Z(n441) );
  NAND U389 ( .A(n445), .B(n446), .Z(n444) );
  NANDN U390 ( .A(A[401]), .B(B[401]), .Z(n446) );
  AND U391 ( .A(n447), .B(n448), .Z(n445) );
  NANDN U392 ( .A(A[400]), .B(B[400]), .Z(n448) );
  NAND U393 ( .A(n449), .B(n450), .Z(n447) );
  NANDN U394 ( .A(B[400]), .B(A[400]), .Z(n450) );
  AND U395 ( .A(n451), .B(n452), .Z(n449) );
  NAND U396 ( .A(n453), .B(n454), .Z(n452) );
  NANDN U397 ( .A(A[399]), .B(B[399]), .Z(n454) );
  AND U398 ( .A(n455), .B(n456), .Z(n453) );
  NANDN U399 ( .A(A[398]), .B(B[398]), .Z(n456) );
  NAND U400 ( .A(n457), .B(n458), .Z(n455) );
  NANDN U401 ( .A(B[398]), .B(A[398]), .Z(n458) );
  AND U402 ( .A(n459), .B(n460), .Z(n457) );
  NAND U403 ( .A(n461), .B(n462), .Z(n460) );
  NANDN U404 ( .A(A[397]), .B(B[397]), .Z(n462) );
  AND U405 ( .A(n463), .B(n464), .Z(n461) );
  NANDN U406 ( .A(A[396]), .B(B[396]), .Z(n464) );
  NAND U407 ( .A(n465), .B(n466), .Z(n463) );
  NANDN U408 ( .A(B[396]), .B(A[396]), .Z(n466) );
  AND U409 ( .A(n467), .B(n468), .Z(n465) );
  NAND U410 ( .A(n469), .B(n470), .Z(n468) );
  NANDN U411 ( .A(A[395]), .B(B[395]), .Z(n470) );
  AND U412 ( .A(n471), .B(n472), .Z(n469) );
  NANDN U413 ( .A(A[394]), .B(B[394]), .Z(n472) );
  NAND U414 ( .A(n473), .B(n474), .Z(n471) );
  NANDN U415 ( .A(B[394]), .B(A[394]), .Z(n474) );
  AND U416 ( .A(n475), .B(n476), .Z(n473) );
  NAND U417 ( .A(n477), .B(n478), .Z(n476) );
  NANDN U418 ( .A(A[393]), .B(B[393]), .Z(n478) );
  AND U419 ( .A(n479), .B(n480), .Z(n477) );
  NANDN U420 ( .A(A[392]), .B(B[392]), .Z(n480) );
  NAND U421 ( .A(n481), .B(n482), .Z(n479) );
  NANDN U422 ( .A(B[392]), .B(A[392]), .Z(n482) );
  AND U423 ( .A(n483), .B(n484), .Z(n481) );
  NAND U424 ( .A(n485), .B(n486), .Z(n484) );
  NANDN U425 ( .A(A[391]), .B(B[391]), .Z(n486) );
  AND U426 ( .A(n487), .B(n488), .Z(n485) );
  NANDN U427 ( .A(A[390]), .B(B[390]), .Z(n488) );
  NAND U428 ( .A(n489), .B(n490), .Z(n487) );
  NANDN U429 ( .A(B[390]), .B(A[390]), .Z(n490) );
  AND U430 ( .A(n491), .B(n492), .Z(n489) );
  NAND U431 ( .A(n493), .B(n494), .Z(n492) );
  NANDN U432 ( .A(A[389]), .B(B[389]), .Z(n494) );
  AND U433 ( .A(n495), .B(n496), .Z(n493) );
  NANDN U434 ( .A(A[388]), .B(B[388]), .Z(n496) );
  NAND U435 ( .A(n497), .B(n498), .Z(n495) );
  NANDN U436 ( .A(B[388]), .B(A[388]), .Z(n498) );
  AND U437 ( .A(n499), .B(n500), .Z(n497) );
  NAND U438 ( .A(n501), .B(n502), .Z(n500) );
  NANDN U439 ( .A(A[387]), .B(B[387]), .Z(n502) );
  AND U440 ( .A(n503), .B(n504), .Z(n501) );
  NANDN U441 ( .A(A[386]), .B(B[386]), .Z(n504) );
  NAND U442 ( .A(n505), .B(n506), .Z(n503) );
  NANDN U443 ( .A(B[386]), .B(A[386]), .Z(n506) );
  AND U444 ( .A(n507), .B(n508), .Z(n505) );
  NAND U445 ( .A(n509), .B(n510), .Z(n508) );
  NANDN U446 ( .A(A[385]), .B(B[385]), .Z(n510) );
  AND U447 ( .A(n511), .B(n512), .Z(n509) );
  NANDN U448 ( .A(A[384]), .B(B[384]), .Z(n512) );
  NAND U449 ( .A(n513), .B(n514), .Z(n511) );
  NANDN U450 ( .A(B[384]), .B(A[384]), .Z(n514) );
  AND U451 ( .A(n515), .B(n516), .Z(n513) );
  NAND U452 ( .A(n517), .B(n518), .Z(n516) );
  NANDN U453 ( .A(A[383]), .B(B[383]), .Z(n518) );
  AND U454 ( .A(n519), .B(n520), .Z(n517) );
  NANDN U455 ( .A(A[382]), .B(B[382]), .Z(n520) );
  NAND U456 ( .A(n521), .B(n522), .Z(n519) );
  NANDN U457 ( .A(B[382]), .B(A[382]), .Z(n522) );
  AND U458 ( .A(n523), .B(n524), .Z(n521) );
  NAND U459 ( .A(n525), .B(n526), .Z(n524) );
  NANDN U460 ( .A(A[381]), .B(B[381]), .Z(n526) );
  AND U461 ( .A(n527), .B(n528), .Z(n525) );
  NANDN U462 ( .A(A[380]), .B(B[380]), .Z(n528) );
  NAND U463 ( .A(n529), .B(n530), .Z(n527) );
  NANDN U464 ( .A(B[380]), .B(A[380]), .Z(n530) );
  AND U465 ( .A(n531), .B(n532), .Z(n529) );
  NAND U466 ( .A(n533), .B(n534), .Z(n532) );
  NANDN U467 ( .A(A[379]), .B(B[379]), .Z(n534) );
  AND U468 ( .A(n535), .B(n536), .Z(n533) );
  NANDN U469 ( .A(A[378]), .B(B[378]), .Z(n536) );
  NAND U470 ( .A(n537), .B(n538), .Z(n535) );
  NANDN U471 ( .A(B[378]), .B(A[378]), .Z(n538) );
  AND U472 ( .A(n539), .B(n540), .Z(n537) );
  NAND U473 ( .A(n541), .B(n542), .Z(n540) );
  NANDN U474 ( .A(A[377]), .B(B[377]), .Z(n542) );
  AND U475 ( .A(n543), .B(n544), .Z(n541) );
  NANDN U476 ( .A(A[376]), .B(B[376]), .Z(n544) );
  NAND U477 ( .A(n545), .B(n546), .Z(n543) );
  NANDN U478 ( .A(B[376]), .B(A[376]), .Z(n546) );
  AND U479 ( .A(n547), .B(n548), .Z(n545) );
  NAND U480 ( .A(n549), .B(n550), .Z(n548) );
  NANDN U481 ( .A(A[375]), .B(B[375]), .Z(n550) );
  AND U482 ( .A(n551), .B(n552), .Z(n549) );
  NANDN U483 ( .A(A[374]), .B(B[374]), .Z(n552) );
  NAND U484 ( .A(n553), .B(n554), .Z(n551) );
  NANDN U485 ( .A(B[374]), .B(A[374]), .Z(n554) );
  AND U486 ( .A(n555), .B(n556), .Z(n553) );
  NAND U487 ( .A(n557), .B(n558), .Z(n556) );
  NANDN U488 ( .A(A[373]), .B(B[373]), .Z(n558) );
  AND U489 ( .A(n559), .B(n560), .Z(n557) );
  NANDN U490 ( .A(A[372]), .B(B[372]), .Z(n560) );
  NAND U491 ( .A(n561), .B(n562), .Z(n559) );
  NANDN U492 ( .A(B[372]), .B(A[372]), .Z(n562) );
  AND U493 ( .A(n563), .B(n564), .Z(n561) );
  NAND U494 ( .A(n565), .B(n566), .Z(n564) );
  NANDN U495 ( .A(A[371]), .B(B[371]), .Z(n566) );
  AND U496 ( .A(n567), .B(n568), .Z(n565) );
  NANDN U497 ( .A(A[370]), .B(B[370]), .Z(n568) );
  NAND U498 ( .A(n569), .B(n570), .Z(n567) );
  NANDN U499 ( .A(B[370]), .B(A[370]), .Z(n570) );
  AND U500 ( .A(n571), .B(n572), .Z(n569) );
  NAND U501 ( .A(n573), .B(n574), .Z(n572) );
  NANDN U502 ( .A(A[369]), .B(B[369]), .Z(n574) );
  AND U503 ( .A(n575), .B(n576), .Z(n573) );
  NANDN U504 ( .A(A[368]), .B(B[368]), .Z(n576) );
  NAND U505 ( .A(n577), .B(n578), .Z(n575) );
  NANDN U506 ( .A(B[368]), .B(A[368]), .Z(n578) );
  AND U507 ( .A(n579), .B(n580), .Z(n577) );
  NAND U508 ( .A(n581), .B(n582), .Z(n580) );
  NANDN U509 ( .A(A[367]), .B(B[367]), .Z(n582) );
  AND U510 ( .A(n583), .B(n584), .Z(n581) );
  NANDN U511 ( .A(A[366]), .B(B[366]), .Z(n584) );
  NAND U512 ( .A(n585), .B(n586), .Z(n583) );
  NANDN U513 ( .A(B[366]), .B(A[366]), .Z(n586) );
  AND U514 ( .A(n587), .B(n588), .Z(n585) );
  NAND U515 ( .A(n589), .B(n590), .Z(n588) );
  NANDN U516 ( .A(A[365]), .B(B[365]), .Z(n590) );
  AND U517 ( .A(n591), .B(n592), .Z(n589) );
  NANDN U518 ( .A(A[364]), .B(B[364]), .Z(n592) );
  NAND U519 ( .A(n593), .B(n594), .Z(n591) );
  NANDN U520 ( .A(B[364]), .B(A[364]), .Z(n594) );
  AND U521 ( .A(n595), .B(n596), .Z(n593) );
  NAND U522 ( .A(n597), .B(n598), .Z(n596) );
  NANDN U523 ( .A(A[363]), .B(B[363]), .Z(n598) );
  AND U524 ( .A(n599), .B(n600), .Z(n597) );
  NANDN U525 ( .A(A[362]), .B(B[362]), .Z(n600) );
  NAND U526 ( .A(n601), .B(n602), .Z(n599) );
  NANDN U527 ( .A(B[362]), .B(A[362]), .Z(n602) );
  AND U528 ( .A(n603), .B(n604), .Z(n601) );
  NAND U529 ( .A(n605), .B(n606), .Z(n604) );
  NANDN U530 ( .A(A[361]), .B(B[361]), .Z(n606) );
  AND U531 ( .A(n607), .B(n608), .Z(n605) );
  NANDN U532 ( .A(A[360]), .B(B[360]), .Z(n608) );
  NAND U533 ( .A(n609), .B(n610), .Z(n607) );
  NANDN U534 ( .A(B[360]), .B(A[360]), .Z(n610) );
  AND U535 ( .A(n611), .B(n612), .Z(n609) );
  NAND U536 ( .A(n613), .B(n614), .Z(n612) );
  NANDN U537 ( .A(A[359]), .B(B[359]), .Z(n614) );
  AND U538 ( .A(n615), .B(n616), .Z(n613) );
  NANDN U539 ( .A(A[358]), .B(B[358]), .Z(n616) );
  NAND U540 ( .A(n617), .B(n618), .Z(n615) );
  NANDN U541 ( .A(B[358]), .B(A[358]), .Z(n618) );
  AND U542 ( .A(n619), .B(n620), .Z(n617) );
  NAND U543 ( .A(n621), .B(n622), .Z(n620) );
  NANDN U544 ( .A(A[357]), .B(B[357]), .Z(n622) );
  AND U545 ( .A(n623), .B(n624), .Z(n621) );
  NANDN U546 ( .A(A[356]), .B(B[356]), .Z(n624) );
  NAND U547 ( .A(n625), .B(n626), .Z(n623) );
  NANDN U548 ( .A(B[356]), .B(A[356]), .Z(n626) );
  AND U549 ( .A(n627), .B(n628), .Z(n625) );
  NAND U550 ( .A(n629), .B(n630), .Z(n628) );
  NANDN U551 ( .A(A[355]), .B(B[355]), .Z(n630) );
  AND U552 ( .A(n631), .B(n632), .Z(n629) );
  NANDN U553 ( .A(A[354]), .B(B[354]), .Z(n632) );
  NAND U554 ( .A(n633), .B(n634), .Z(n631) );
  NANDN U555 ( .A(B[354]), .B(A[354]), .Z(n634) );
  AND U556 ( .A(n635), .B(n636), .Z(n633) );
  NAND U557 ( .A(n637), .B(n638), .Z(n636) );
  NANDN U558 ( .A(A[353]), .B(B[353]), .Z(n638) );
  AND U559 ( .A(n639), .B(n640), .Z(n637) );
  NANDN U560 ( .A(A[352]), .B(B[352]), .Z(n640) );
  NAND U561 ( .A(n641), .B(n642), .Z(n639) );
  NANDN U562 ( .A(B[352]), .B(A[352]), .Z(n642) );
  AND U563 ( .A(n643), .B(n644), .Z(n641) );
  NAND U564 ( .A(n645), .B(n646), .Z(n644) );
  NANDN U565 ( .A(A[351]), .B(B[351]), .Z(n646) );
  AND U566 ( .A(n647), .B(n648), .Z(n645) );
  NANDN U567 ( .A(A[350]), .B(B[350]), .Z(n648) );
  NAND U568 ( .A(n649), .B(n650), .Z(n647) );
  NANDN U569 ( .A(B[350]), .B(A[350]), .Z(n650) );
  AND U570 ( .A(n651), .B(n652), .Z(n649) );
  NAND U571 ( .A(n653), .B(n654), .Z(n652) );
  NANDN U572 ( .A(A[349]), .B(B[349]), .Z(n654) );
  AND U573 ( .A(n655), .B(n656), .Z(n653) );
  NANDN U574 ( .A(A[348]), .B(B[348]), .Z(n656) );
  NAND U575 ( .A(n657), .B(n658), .Z(n655) );
  NANDN U576 ( .A(B[348]), .B(A[348]), .Z(n658) );
  AND U577 ( .A(n659), .B(n660), .Z(n657) );
  NAND U578 ( .A(n661), .B(n662), .Z(n660) );
  NANDN U579 ( .A(A[347]), .B(B[347]), .Z(n662) );
  AND U580 ( .A(n663), .B(n664), .Z(n661) );
  NANDN U581 ( .A(A[346]), .B(B[346]), .Z(n664) );
  NAND U582 ( .A(n665), .B(n666), .Z(n663) );
  NANDN U583 ( .A(B[346]), .B(A[346]), .Z(n666) );
  AND U584 ( .A(n667), .B(n668), .Z(n665) );
  NAND U585 ( .A(n669), .B(n670), .Z(n668) );
  NANDN U586 ( .A(A[345]), .B(B[345]), .Z(n670) );
  AND U587 ( .A(n671), .B(n672), .Z(n669) );
  NANDN U588 ( .A(A[344]), .B(B[344]), .Z(n672) );
  NAND U589 ( .A(n673), .B(n674), .Z(n671) );
  NANDN U590 ( .A(B[344]), .B(A[344]), .Z(n674) );
  AND U591 ( .A(n675), .B(n676), .Z(n673) );
  NAND U592 ( .A(n677), .B(n678), .Z(n676) );
  NANDN U593 ( .A(A[343]), .B(B[343]), .Z(n678) );
  AND U594 ( .A(n679), .B(n680), .Z(n677) );
  NANDN U595 ( .A(A[342]), .B(B[342]), .Z(n680) );
  NAND U596 ( .A(n681), .B(n682), .Z(n679) );
  NANDN U597 ( .A(B[342]), .B(A[342]), .Z(n682) );
  AND U598 ( .A(n683), .B(n684), .Z(n681) );
  NAND U599 ( .A(n685), .B(n686), .Z(n684) );
  NANDN U600 ( .A(A[341]), .B(B[341]), .Z(n686) );
  AND U601 ( .A(n687), .B(n688), .Z(n685) );
  NANDN U602 ( .A(A[340]), .B(B[340]), .Z(n688) );
  NAND U603 ( .A(n689), .B(n690), .Z(n687) );
  NANDN U604 ( .A(B[340]), .B(A[340]), .Z(n690) );
  AND U605 ( .A(n691), .B(n692), .Z(n689) );
  NAND U606 ( .A(n693), .B(n694), .Z(n692) );
  NANDN U607 ( .A(A[339]), .B(B[339]), .Z(n694) );
  AND U608 ( .A(n695), .B(n696), .Z(n693) );
  NANDN U609 ( .A(A[338]), .B(B[338]), .Z(n696) );
  NAND U610 ( .A(n697), .B(n698), .Z(n695) );
  NANDN U611 ( .A(B[338]), .B(A[338]), .Z(n698) );
  AND U612 ( .A(n699), .B(n700), .Z(n697) );
  NAND U613 ( .A(n701), .B(n702), .Z(n700) );
  NANDN U614 ( .A(A[337]), .B(B[337]), .Z(n702) );
  AND U615 ( .A(n703), .B(n704), .Z(n701) );
  NANDN U616 ( .A(A[336]), .B(B[336]), .Z(n704) );
  NAND U617 ( .A(n705), .B(n706), .Z(n703) );
  NANDN U618 ( .A(B[336]), .B(A[336]), .Z(n706) );
  AND U619 ( .A(n707), .B(n708), .Z(n705) );
  NAND U620 ( .A(n709), .B(n710), .Z(n708) );
  NANDN U621 ( .A(A[335]), .B(B[335]), .Z(n710) );
  AND U622 ( .A(n711), .B(n712), .Z(n709) );
  NANDN U623 ( .A(A[334]), .B(B[334]), .Z(n712) );
  NAND U624 ( .A(n713), .B(n714), .Z(n711) );
  NANDN U625 ( .A(B[334]), .B(A[334]), .Z(n714) );
  AND U626 ( .A(n715), .B(n716), .Z(n713) );
  NAND U627 ( .A(n717), .B(n718), .Z(n716) );
  NANDN U628 ( .A(A[333]), .B(B[333]), .Z(n718) );
  AND U629 ( .A(n719), .B(n720), .Z(n717) );
  NANDN U630 ( .A(A[332]), .B(B[332]), .Z(n720) );
  NAND U631 ( .A(n721), .B(n722), .Z(n719) );
  NANDN U632 ( .A(B[332]), .B(A[332]), .Z(n722) );
  AND U633 ( .A(n723), .B(n724), .Z(n721) );
  NAND U634 ( .A(n725), .B(n726), .Z(n724) );
  NANDN U635 ( .A(A[331]), .B(B[331]), .Z(n726) );
  AND U636 ( .A(n727), .B(n728), .Z(n725) );
  NANDN U637 ( .A(A[330]), .B(B[330]), .Z(n728) );
  NAND U638 ( .A(n729), .B(n730), .Z(n727) );
  NANDN U639 ( .A(B[330]), .B(A[330]), .Z(n730) );
  AND U640 ( .A(n731), .B(n732), .Z(n729) );
  NAND U641 ( .A(n733), .B(n734), .Z(n732) );
  NANDN U642 ( .A(A[329]), .B(B[329]), .Z(n734) );
  AND U643 ( .A(n735), .B(n736), .Z(n733) );
  NANDN U644 ( .A(A[328]), .B(B[328]), .Z(n736) );
  NAND U645 ( .A(n737), .B(n738), .Z(n735) );
  NANDN U646 ( .A(B[328]), .B(A[328]), .Z(n738) );
  AND U647 ( .A(n739), .B(n740), .Z(n737) );
  NAND U648 ( .A(n741), .B(n742), .Z(n740) );
  NANDN U649 ( .A(A[327]), .B(B[327]), .Z(n742) );
  AND U650 ( .A(n743), .B(n744), .Z(n741) );
  NANDN U651 ( .A(A[326]), .B(B[326]), .Z(n744) );
  NAND U652 ( .A(n745), .B(n746), .Z(n743) );
  NANDN U653 ( .A(B[326]), .B(A[326]), .Z(n746) );
  AND U654 ( .A(n747), .B(n748), .Z(n745) );
  NAND U655 ( .A(n749), .B(n750), .Z(n748) );
  NANDN U656 ( .A(A[325]), .B(B[325]), .Z(n750) );
  AND U657 ( .A(n751), .B(n752), .Z(n749) );
  NANDN U658 ( .A(A[324]), .B(B[324]), .Z(n752) );
  NAND U659 ( .A(n753), .B(n754), .Z(n751) );
  NANDN U660 ( .A(B[324]), .B(A[324]), .Z(n754) );
  AND U661 ( .A(n755), .B(n756), .Z(n753) );
  NAND U662 ( .A(n757), .B(n758), .Z(n756) );
  NANDN U663 ( .A(A[323]), .B(B[323]), .Z(n758) );
  AND U664 ( .A(n759), .B(n760), .Z(n757) );
  NANDN U665 ( .A(A[322]), .B(B[322]), .Z(n760) );
  NAND U666 ( .A(n761), .B(n762), .Z(n759) );
  NANDN U667 ( .A(B[322]), .B(A[322]), .Z(n762) );
  AND U668 ( .A(n763), .B(n764), .Z(n761) );
  NAND U669 ( .A(n765), .B(n766), .Z(n764) );
  NANDN U670 ( .A(A[321]), .B(B[321]), .Z(n766) );
  AND U671 ( .A(n767), .B(n768), .Z(n765) );
  NANDN U672 ( .A(A[320]), .B(B[320]), .Z(n768) );
  NAND U673 ( .A(n769), .B(n770), .Z(n767) );
  NANDN U674 ( .A(B[320]), .B(A[320]), .Z(n770) );
  AND U675 ( .A(n771), .B(n772), .Z(n769) );
  NAND U676 ( .A(n773), .B(n774), .Z(n772) );
  NANDN U677 ( .A(A[319]), .B(B[319]), .Z(n774) );
  AND U678 ( .A(n775), .B(n776), .Z(n773) );
  NANDN U679 ( .A(A[318]), .B(B[318]), .Z(n776) );
  NAND U680 ( .A(n777), .B(n778), .Z(n775) );
  NANDN U681 ( .A(B[318]), .B(A[318]), .Z(n778) );
  AND U682 ( .A(n779), .B(n780), .Z(n777) );
  NAND U683 ( .A(n781), .B(n782), .Z(n780) );
  NANDN U684 ( .A(A[317]), .B(B[317]), .Z(n782) );
  AND U685 ( .A(n783), .B(n784), .Z(n781) );
  NANDN U686 ( .A(A[316]), .B(B[316]), .Z(n784) );
  NAND U687 ( .A(n785), .B(n786), .Z(n783) );
  NANDN U688 ( .A(B[316]), .B(A[316]), .Z(n786) );
  AND U689 ( .A(n787), .B(n788), .Z(n785) );
  NAND U690 ( .A(n789), .B(n790), .Z(n788) );
  NANDN U691 ( .A(A[315]), .B(B[315]), .Z(n790) );
  AND U692 ( .A(n791), .B(n792), .Z(n789) );
  NANDN U693 ( .A(A[314]), .B(B[314]), .Z(n792) );
  NAND U694 ( .A(n793), .B(n794), .Z(n791) );
  NANDN U695 ( .A(B[314]), .B(A[314]), .Z(n794) );
  AND U696 ( .A(n795), .B(n796), .Z(n793) );
  NAND U697 ( .A(n797), .B(n798), .Z(n796) );
  NANDN U698 ( .A(A[313]), .B(B[313]), .Z(n798) );
  AND U699 ( .A(n799), .B(n800), .Z(n797) );
  NANDN U700 ( .A(A[312]), .B(B[312]), .Z(n800) );
  NAND U701 ( .A(n801), .B(n802), .Z(n799) );
  NANDN U702 ( .A(B[312]), .B(A[312]), .Z(n802) );
  AND U703 ( .A(n803), .B(n804), .Z(n801) );
  NAND U704 ( .A(n805), .B(n806), .Z(n804) );
  NANDN U705 ( .A(A[311]), .B(B[311]), .Z(n806) );
  AND U706 ( .A(n807), .B(n808), .Z(n805) );
  NANDN U707 ( .A(A[310]), .B(B[310]), .Z(n808) );
  NAND U708 ( .A(n809), .B(n810), .Z(n807) );
  NANDN U709 ( .A(B[310]), .B(A[310]), .Z(n810) );
  AND U710 ( .A(n811), .B(n812), .Z(n809) );
  NAND U711 ( .A(n813), .B(n814), .Z(n812) );
  NANDN U712 ( .A(A[309]), .B(B[309]), .Z(n814) );
  AND U713 ( .A(n815), .B(n816), .Z(n813) );
  NANDN U714 ( .A(A[308]), .B(B[308]), .Z(n816) );
  NAND U715 ( .A(n817), .B(n818), .Z(n815) );
  NANDN U716 ( .A(B[308]), .B(A[308]), .Z(n818) );
  AND U717 ( .A(n819), .B(n820), .Z(n817) );
  NAND U718 ( .A(n821), .B(n822), .Z(n820) );
  NANDN U719 ( .A(A[307]), .B(B[307]), .Z(n822) );
  AND U720 ( .A(n823), .B(n824), .Z(n821) );
  NANDN U721 ( .A(A[306]), .B(B[306]), .Z(n824) );
  NAND U722 ( .A(n825), .B(n826), .Z(n823) );
  NANDN U723 ( .A(B[306]), .B(A[306]), .Z(n826) );
  AND U724 ( .A(n827), .B(n828), .Z(n825) );
  NAND U725 ( .A(n829), .B(n830), .Z(n828) );
  NANDN U726 ( .A(A[305]), .B(B[305]), .Z(n830) );
  AND U727 ( .A(n831), .B(n832), .Z(n829) );
  NANDN U728 ( .A(A[304]), .B(B[304]), .Z(n832) );
  NAND U729 ( .A(n833), .B(n834), .Z(n831) );
  NANDN U730 ( .A(B[304]), .B(A[304]), .Z(n834) );
  AND U731 ( .A(n835), .B(n836), .Z(n833) );
  NAND U732 ( .A(n837), .B(n838), .Z(n836) );
  NANDN U733 ( .A(A[303]), .B(B[303]), .Z(n838) );
  AND U734 ( .A(n839), .B(n840), .Z(n837) );
  NANDN U735 ( .A(A[302]), .B(B[302]), .Z(n840) );
  NAND U736 ( .A(n841), .B(n842), .Z(n839) );
  NANDN U737 ( .A(B[302]), .B(A[302]), .Z(n842) );
  AND U738 ( .A(n843), .B(n844), .Z(n841) );
  NAND U739 ( .A(n845), .B(n846), .Z(n844) );
  NANDN U740 ( .A(A[301]), .B(B[301]), .Z(n846) );
  AND U741 ( .A(n847), .B(n848), .Z(n845) );
  NANDN U742 ( .A(A[300]), .B(B[300]), .Z(n848) );
  NAND U743 ( .A(n849), .B(n850), .Z(n847) );
  NANDN U744 ( .A(B[300]), .B(A[300]), .Z(n850) );
  AND U745 ( .A(n851), .B(n852), .Z(n849) );
  NAND U746 ( .A(n853), .B(n854), .Z(n852) );
  NANDN U747 ( .A(A[299]), .B(B[299]), .Z(n854) );
  AND U748 ( .A(n855), .B(n856), .Z(n853) );
  NANDN U749 ( .A(A[298]), .B(B[298]), .Z(n856) );
  NAND U750 ( .A(n857), .B(n858), .Z(n855) );
  NANDN U751 ( .A(B[298]), .B(A[298]), .Z(n858) );
  AND U752 ( .A(n859), .B(n860), .Z(n857) );
  NAND U753 ( .A(n861), .B(n862), .Z(n860) );
  NANDN U754 ( .A(A[297]), .B(B[297]), .Z(n862) );
  AND U755 ( .A(n863), .B(n864), .Z(n861) );
  NANDN U756 ( .A(A[296]), .B(B[296]), .Z(n864) );
  NAND U757 ( .A(n865), .B(n866), .Z(n863) );
  NANDN U758 ( .A(B[296]), .B(A[296]), .Z(n866) );
  AND U759 ( .A(n867), .B(n868), .Z(n865) );
  NAND U760 ( .A(n869), .B(n870), .Z(n868) );
  NANDN U761 ( .A(A[295]), .B(B[295]), .Z(n870) );
  AND U762 ( .A(n871), .B(n872), .Z(n869) );
  NANDN U763 ( .A(A[294]), .B(B[294]), .Z(n872) );
  NAND U764 ( .A(n873), .B(n874), .Z(n871) );
  NANDN U765 ( .A(B[294]), .B(A[294]), .Z(n874) );
  AND U766 ( .A(n875), .B(n876), .Z(n873) );
  NAND U767 ( .A(n877), .B(n878), .Z(n876) );
  NANDN U768 ( .A(A[293]), .B(B[293]), .Z(n878) );
  AND U769 ( .A(n879), .B(n880), .Z(n877) );
  NANDN U770 ( .A(A[292]), .B(B[292]), .Z(n880) );
  NAND U771 ( .A(n881), .B(n882), .Z(n879) );
  NANDN U772 ( .A(B[292]), .B(A[292]), .Z(n882) );
  AND U773 ( .A(n883), .B(n884), .Z(n881) );
  NAND U774 ( .A(n885), .B(n886), .Z(n884) );
  NANDN U775 ( .A(A[291]), .B(B[291]), .Z(n886) );
  AND U776 ( .A(n887), .B(n888), .Z(n885) );
  NANDN U777 ( .A(A[290]), .B(B[290]), .Z(n888) );
  NAND U778 ( .A(n889), .B(n890), .Z(n887) );
  NANDN U779 ( .A(B[290]), .B(A[290]), .Z(n890) );
  AND U780 ( .A(n891), .B(n892), .Z(n889) );
  NAND U781 ( .A(n893), .B(n894), .Z(n892) );
  NANDN U782 ( .A(A[289]), .B(B[289]), .Z(n894) );
  AND U783 ( .A(n895), .B(n896), .Z(n893) );
  NANDN U784 ( .A(A[288]), .B(B[288]), .Z(n896) );
  NAND U785 ( .A(n897), .B(n898), .Z(n895) );
  NANDN U786 ( .A(B[288]), .B(A[288]), .Z(n898) );
  AND U787 ( .A(n899), .B(n900), .Z(n897) );
  NAND U788 ( .A(n901), .B(n902), .Z(n900) );
  NANDN U789 ( .A(A[287]), .B(B[287]), .Z(n902) );
  AND U790 ( .A(n903), .B(n904), .Z(n901) );
  NANDN U791 ( .A(A[286]), .B(B[286]), .Z(n904) );
  NAND U792 ( .A(n905), .B(n906), .Z(n903) );
  NANDN U793 ( .A(B[286]), .B(A[286]), .Z(n906) );
  AND U794 ( .A(n907), .B(n908), .Z(n905) );
  NAND U795 ( .A(n909), .B(n910), .Z(n908) );
  NANDN U796 ( .A(A[285]), .B(B[285]), .Z(n910) );
  AND U797 ( .A(n911), .B(n912), .Z(n909) );
  NANDN U798 ( .A(A[284]), .B(B[284]), .Z(n912) );
  NAND U799 ( .A(n913), .B(n914), .Z(n911) );
  NANDN U800 ( .A(B[284]), .B(A[284]), .Z(n914) );
  AND U801 ( .A(n915), .B(n916), .Z(n913) );
  NAND U802 ( .A(n917), .B(n918), .Z(n916) );
  NANDN U803 ( .A(A[283]), .B(B[283]), .Z(n918) );
  AND U804 ( .A(n919), .B(n920), .Z(n917) );
  NANDN U805 ( .A(A[282]), .B(B[282]), .Z(n920) );
  NAND U806 ( .A(n921), .B(n922), .Z(n919) );
  NANDN U807 ( .A(B[282]), .B(A[282]), .Z(n922) );
  AND U808 ( .A(n923), .B(n924), .Z(n921) );
  NAND U809 ( .A(n925), .B(n926), .Z(n924) );
  NANDN U810 ( .A(A[281]), .B(B[281]), .Z(n926) );
  AND U811 ( .A(n927), .B(n928), .Z(n925) );
  NANDN U812 ( .A(A[280]), .B(B[280]), .Z(n928) );
  NAND U813 ( .A(n929), .B(n930), .Z(n927) );
  NANDN U814 ( .A(B[280]), .B(A[280]), .Z(n930) );
  AND U815 ( .A(n931), .B(n932), .Z(n929) );
  NAND U816 ( .A(n933), .B(n934), .Z(n932) );
  NANDN U817 ( .A(A[279]), .B(B[279]), .Z(n934) );
  AND U818 ( .A(n935), .B(n936), .Z(n933) );
  NANDN U819 ( .A(A[278]), .B(B[278]), .Z(n936) );
  NAND U820 ( .A(n937), .B(n938), .Z(n935) );
  NANDN U821 ( .A(B[278]), .B(A[278]), .Z(n938) );
  AND U822 ( .A(n939), .B(n940), .Z(n937) );
  NAND U823 ( .A(n941), .B(n942), .Z(n940) );
  NANDN U824 ( .A(A[277]), .B(B[277]), .Z(n942) );
  AND U825 ( .A(n943), .B(n944), .Z(n941) );
  NANDN U826 ( .A(A[276]), .B(B[276]), .Z(n944) );
  NAND U827 ( .A(n945), .B(n946), .Z(n943) );
  NANDN U828 ( .A(B[276]), .B(A[276]), .Z(n946) );
  AND U829 ( .A(n947), .B(n948), .Z(n945) );
  NAND U830 ( .A(n949), .B(n950), .Z(n948) );
  NANDN U831 ( .A(A[275]), .B(B[275]), .Z(n950) );
  AND U832 ( .A(n951), .B(n952), .Z(n949) );
  NANDN U833 ( .A(A[274]), .B(B[274]), .Z(n952) );
  NAND U834 ( .A(n953), .B(n954), .Z(n951) );
  NANDN U835 ( .A(B[274]), .B(A[274]), .Z(n954) );
  AND U836 ( .A(n955), .B(n956), .Z(n953) );
  NAND U837 ( .A(n957), .B(n958), .Z(n956) );
  NANDN U838 ( .A(A[273]), .B(B[273]), .Z(n958) );
  AND U839 ( .A(n959), .B(n960), .Z(n957) );
  NANDN U840 ( .A(A[272]), .B(B[272]), .Z(n960) );
  NAND U841 ( .A(n961), .B(n962), .Z(n959) );
  NANDN U842 ( .A(B[272]), .B(A[272]), .Z(n962) );
  AND U843 ( .A(n963), .B(n964), .Z(n961) );
  NAND U844 ( .A(n965), .B(n966), .Z(n964) );
  NANDN U845 ( .A(A[271]), .B(B[271]), .Z(n966) );
  AND U846 ( .A(n967), .B(n968), .Z(n965) );
  NANDN U847 ( .A(A[270]), .B(B[270]), .Z(n968) );
  NAND U848 ( .A(n969), .B(n970), .Z(n967) );
  NANDN U849 ( .A(B[270]), .B(A[270]), .Z(n970) );
  AND U850 ( .A(n971), .B(n972), .Z(n969) );
  NAND U851 ( .A(n973), .B(n974), .Z(n972) );
  NANDN U852 ( .A(A[269]), .B(B[269]), .Z(n974) );
  AND U853 ( .A(n975), .B(n976), .Z(n973) );
  NANDN U854 ( .A(A[268]), .B(B[268]), .Z(n976) );
  NAND U855 ( .A(n977), .B(n978), .Z(n975) );
  NANDN U856 ( .A(B[268]), .B(A[268]), .Z(n978) );
  AND U857 ( .A(n979), .B(n980), .Z(n977) );
  NAND U858 ( .A(n981), .B(n982), .Z(n980) );
  NANDN U859 ( .A(A[267]), .B(B[267]), .Z(n982) );
  AND U860 ( .A(n983), .B(n984), .Z(n981) );
  NANDN U861 ( .A(A[266]), .B(B[266]), .Z(n984) );
  NAND U862 ( .A(n985), .B(n986), .Z(n983) );
  NANDN U863 ( .A(B[266]), .B(A[266]), .Z(n986) );
  AND U864 ( .A(n987), .B(n988), .Z(n985) );
  NAND U865 ( .A(n989), .B(n990), .Z(n988) );
  NANDN U866 ( .A(A[265]), .B(B[265]), .Z(n990) );
  AND U867 ( .A(n991), .B(n992), .Z(n989) );
  NANDN U868 ( .A(A[264]), .B(B[264]), .Z(n992) );
  NAND U869 ( .A(n993), .B(n994), .Z(n991) );
  NANDN U870 ( .A(B[264]), .B(A[264]), .Z(n994) );
  AND U871 ( .A(n995), .B(n996), .Z(n993) );
  NAND U872 ( .A(n997), .B(n998), .Z(n996) );
  NANDN U873 ( .A(A[263]), .B(B[263]), .Z(n998) );
  AND U874 ( .A(n999), .B(n1000), .Z(n997) );
  NANDN U875 ( .A(A[262]), .B(B[262]), .Z(n1000) );
  NAND U876 ( .A(n1001), .B(n1002), .Z(n999) );
  NANDN U877 ( .A(B[262]), .B(A[262]), .Z(n1002) );
  AND U878 ( .A(n1003), .B(n1004), .Z(n1001) );
  NAND U879 ( .A(n1005), .B(n1006), .Z(n1004) );
  NANDN U880 ( .A(A[261]), .B(B[261]), .Z(n1006) );
  AND U881 ( .A(n1007), .B(n1008), .Z(n1005) );
  NANDN U882 ( .A(A[260]), .B(B[260]), .Z(n1008) );
  NAND U883 ( .A(n1009), .B(n1010), .Z(n1007) );
  NANDN U884 ( .A(B[260]), .B(A[260]), .Z(n1010) );
  AND U885 ( .A(n1011), .B(n1012), .Z(n1009) );
  NAND U886 ( .A(n1013), .B(n1014), .Z(n1012) );
  NANDN U887 ( .A(A[259]), .B(B[259]), .Z(n1014) );
  AND U888 ( .A(n1015), .B(n1016), .Z(n1013) );
  NANDN U889 ( .A(A[258]), .B(B[258]), .Z(n1016) );
  NAND U890 ( .A(n1017), .B(n1018), .Z(n1015) );
  NANDN U891 ( .A(B[258]), .B(A[258]), .Z(n1018) );
  AND U892 ( .A(n1019), .B(n1020), .Z(n1017) );
  NAND U893 ( .A(n1021), .B(n1022), .Z(n1020) );
  NANDN U894 ( .A(A[257]), .B(B[257]), .Z(n1022) );
  AND U895 ( .A(n1023), .B(n1024), .Z(n1021) );
  NANDN U896 ( .A(A[256]), .B(B[256]), .Z(n1024) );
  NAND U897 ( .A(n1025), .B(n1026), .Z(n1023) );
  NANDN U898 ( .A(B[256]), .B(A[256]), .Z(n1026) );
  AND U899 ( .A(n1027), .B(n1028), .Z(n1025) );
  NAND U900 ( .A(n1029), .B(n1030), .Z(n1028) );
  NANDN U901 ( .A(A[255]), .B(B[255]), .Z(n1030) );
  AND U902 ( .A(n1031), .B(n1032), .Z(n1029) );
  NANDN U903 ( .A(A[254]), .B(B[254]), .Z(n1032) );
  NAND U904 ( .A(n1033), .B(n1034), .Z(n1031) );
  NANDN U905 ( .A(B[254]), .B(A[254]), .Z(n1034) );
  AND U906 ( .A(n1035), .B(n1036), .Z(n1033) );
  NAND U907 ( .A(n1037), .B(n1038), .Z(n1036) );
  NANDN U908 ( .A(A[253]), .B(B[253]), .Z(n1038) );
  AND U909 ( .A(n1039), .B(n1040), .Z(n1037) );
  NANDN U910 ( .A(A[252]), .B(B[252]), .Z(n1040) );
  NAND U911 ( .A(n1041), .B(n1042), .Z(n1039) );
  NANDN U912 ( .A(B[252]), .B(A[252]), .Z(n1042) );
  AND U913 ( .A(n1043), .B(n1044), .Z(n1041) );
  NAND U914 ( .A(n1045), .B(n1046), .Z(n1044) );
  NANDN U915 ( .A(A[251]), .B(B[251]), .Z(n1046) );
  AND U916 ( .A(n1047), .B(n1048), .Z(n1045) );
  NANDN U917 ( .A(A[250]), .B(B[250]), .Z(n1048) );
  NAND U918 ( .A(n1049), .B(n1050), .Z(n1047) );
  NANDN U919 ( .A(B[250]), .B(A[250]), .Z(n1050) );
  AND U920 ( .A(n1051), .B(n1052), .Z(n1049) );
  NAND U921 ( .A(n1053), .B(n1054), .Z(n1052) );
  NANDN U922 ( .A(A[249]), .B(B[249]), .Z(n1054) );
  AND U923 ( .A(n1055), .B(n1056), .Z(n1053) );
  NANDN U924 ( .A(A[248]), .B(B[248]), .Z(n1056) );
  NAND U925 ( .A(n1057), .B(n1058), .Z(n1055) );
  NANDN U926 ( .A(B[248]), .B(A[248]), .Z(n1058) );
  AND U927 ( .A(n1059), .B(n1060), .Z(n1057) );
  NAND U928 ( .A(n1061), .B(n1062), .Z(n1060) );
  NANDN U929 ( .A(A[247]), .B(B[247]), .Z(n1062) );
  AND U930 ( .A(n1063), .B(n1064), .Z(n1061) );
  NANDN U931 ( .A(A[246]), .B(B[246]), .Z(n1064) );
  NAND U932 ( .A(n1065), .B(n1066), .Z(n1063) );
  NANDN U933 ( .A(B[246]), .B(A[246]), .Z(n1066) );
  AND U934 ( .A(n1067), .B(n1068), .Z(n1065) );
  NAND U935 ( .A(n1069), .B(n1070), .Z(n1068) );
  NANDN U936 ( .A(A[245]), .B(B[245]), .Z(n1070) );
  AND U937 ( .A(n1071), .B(n1072), .Z(n1069) );
  NANDN U938 ( .A(A[244]), .B(B[244]), .Z(n1072) );
  NAND U939 ( .A(n1073), .B(n1074), .Z(n1071) );
  NANDN U940 ( .A(B[244]), .B(A[244]), .Z(n1074) );
  AND U941 ( .A(n1075), .B(n1076), .Z(n1073) );
  NAND U942 ( .A(n1077), .B(n1078), .Z(n1076) );
  NANDN U943 ( .A(A[243]), .B(B[243]), .Z(n1078) );
  AND U944 ( .A(n1079), .B(n1080), .Z(n1077) );
  NANDN U945 ( .A(A[242]), .B(B[242]), .Z(n1080) );
  NAND U946 ( .A(n1081), .B(n1082), .Z(n1079) );
  NANDN U947 ( .A(B[242]), .B(A[242]), .Z(n1082) );
  AND U948 ( .A(n1083), .B(n1084), .Z(n1081) );
  NAND U949 ( .A(n1085), .B(n1086), .Z(n1084) );
  NANDN U950 ( .A(A[241]), .B(B[241]), .Z(n1086) );
  AND U951 ( .A(n1087), .B(n1088), .Z(n1085) );
  NANDN U952 ( .A(A[240]), .B(B[240]), .Z(n1088) );
  NAND U953 ( .A(n1089), .B(n1090), .Z(n1087) );
  NANDN U954 ( .A(B[240]), .B(A[240]), .Z(n1090) );
  AND U955 ( .A(n1091), .B(n1092), .Z(n1089) );
  NAND U956 ( .A(n1093), .B(n1094), .Z(n1092) );
  NANDN U957 ( .A(A[239]), .B(B[239]), .Z(n1094) );
  AND U958 ( .A(n1095), .B(n1096), .Z(n1093) );
  NANDN U959 ( .A(A[238]), .B(B[238]), .Z(n1096) );
  NAND U960 ( .A(n1097), .B(n1098), .Z(n1095) );
  NANDN U961 ( .A(B[238]), .B(A[238]), .Z(n1098) );
  AND U962 ( .A(n1099), .B(n1100), .Z(n1097) );
  NAND U963 ( .A(n1101), .B(n1102), .Z(n1100) );
  NANDN U964 ( .A(A[237]), .B(B[237]), .Z(n1102) );
  AND U965 ( .A(n1103), .B(n1104), .Z(n1101) );
  NANDN U966 ( .A(A[236]), .B(B[236]), .Z(n1104) );
  NAND U967 ( .A(n1105), .B(n1106), .Z(n1103) );
  NANDN U968 ( .A(B[236]), .B(A[236]), .Z(n1106) );
  AND U969 ( .A(n1107), .B(n1108), .Z(n1105) );
  NAND U970 ( .A(n1109), .B(n1110), .Z(n1108) );
  NANDN U971 ( .A(A[235]), .B(B[235]), .Z(n1110) );
  AND U972 ( .A(n1111), .B(n1112), .Z(n1109) );
  NANDN U973 ( .A(A[234]), .B(B[234]), .Z(n1112) );
  NAND U974 ( .A(n1113), .B(n1114), .Z(n1111) );
  NANDN U975 ( .A(B[234]), .B(A[234]), .Z(n1114) );
  AND U976 ( .A(n1115), .B(n1116), .Z(n1113) );
  NAND U977 ( .A(n1117), .B(n1118), .Z(n1116) );
  NANDN U978 ( .A(A[233]), .B(B[233]), .Z(n1118) );
  AND U979 ( .A(n1119), .B(n1120), .Z(n1117) );
  NANDN U980 ( .A(A[232]), .B(B[232]), .Z(n1120) );
  NAND U981 ( .A(n1121), .B(n1122), .Z(n1119) );
  NANDN U982 ( .A(B[232]), .B(A[232]), .Z(n1122) );
  AND U983 ( .A(n1123), .B(n1124), .Z(n1121) );
  NAND U984 ( .A(n1125), .B(n1126), .Z(n1124) );
  NANDN U985 ( .A(A[231]), .B(B[231]), .Z(n1126) );
  AND U986 ( .A(n1127), .B(n1128), .Z(n1125) );
  NANDN U987 ( .A(A[230]), .B(B[230]), .Z(n1128) );
  NAND U988 ( .A(n1129), .B(n1130), .Z(n1127) );
  NANDN U989 ( .A(B[230]), .B(A[230]), .Z(n1130) );
  AND U990 ( .A(n1131), .B(n1132), .Z(n1129) );
  NAND U991 ( .A(n1133), .B(n1134), .Z(n1132) );
  NANDN U992 ( .A(A[229]), .B(B[229]), .Z(n1134) );
  AND U993 ( .A(n1135), .B(n1136), .Z(n1133) );
  NANDN U994 ( .A(A[228]), .B(B[228]), .Z(n1136) );
  NAND U995 ( .A(n1137), .B(n1138), .Z(n1135) );
  NANDN U996 ( .A(B[228]), .B(A[228]), .Z(n1138) );
  AND U997 ( .A(n1139), .B(n1140), .Z(n1137) );
  NAND U998 ( .A(n1141), .B(n1142), .Z(n1140) );
  NANDN U999 ( .A(A[227]), .B(B[227]), .Z(n1142) );
  AND U1000 ( .A(n1143), .B(n1144), .Z(n1141) );
  NANDN U1001 ( .A(A[226]), .B(B[226]), .Z(n1144) );
  NAND U1002 ( .A(n1145), .B(n1146), .Z(n1143) );
  NANDN U1003 ( .A(B[226]), .B(A[226]), .Z(n1146) );
  AND U1004 ( .A(n1147), .B(n1148), .Z(n1145) );
  NAND U1005 ( .A(n1149), .B(n1150), .Z(n1148) );
  NANDN U1006 ( .A(A[225]), .B(B[225]), .Z(n1150) );
  AND U1007 ( .A(n1151), .B(n1152), .Z(n1149) );
  NANDN U1008 ( .A(A[224]), .B(B[224]), .Z(n1152) );
  NAND U1009 ( .A(n1153), .B(n1154), .Z(n1151) );
  NANDN U1010 ( .A(B[224]), .B(A[224]), .Z(n1154) );
  AND U1011 ( .A(n1155), .B(n1156), .Z(n1153) );
  NAND U1012 ( .A(n1157), .B(n1158), .Z(n1156) );
  NANDN U1013 ( .A(A[223]), .B(B[223]), .Z(n1158) );
  AND U1014 ( .A(n1159), .B(n1160), .Z(n1157) );
  NANDN U1015 ( .A(A[222]), .B(B[222]), .Z(n1160) );
  NAND U1016 ( .A(n1161), .B(n1162), .Z(n1159) );
  NANDN U1017 ( .A(B[222]), .B(A[222]), .Z(n1162) );
  AND U1018 ( .A(n1163), .B(n1164), .Z(n1161) );
  NAND U1019 ( .A(n1165), .B(n1166), .Z(n1164) );
  NANDN U1020 ( .A(A[221]), .B(B[221]), .Z(n1166) );
  AND U1021 ( .A(n1167), .B(n1168), .Z(n1165) );
  NANDN U1022 ( .A(A[220]), .B(B[220]), .Z(n1168) );
  NAND U1023 ( .A(n1169), .B(n1170), .Z(n1167) );
  NANDN U1024 ( .A(B[220]), .B(A[220]), .Z(n1170) );
  AND U1025 ( .A(n1171), .B(n1172), .Z(n1169) );
  NAND U1026 ( .A(n1173), .B(n1174), .Z(n1172) );
  NANDN U1027 ( .A(A[219]), .B(B[219]), .Z(n1174) );
  AND U1028 ( .A(n1175), .B(n1176), .Z(n1173) );
  NANDN U1029 ( .A(A[218]), .B(B[218]), .Z(n1176) );
  NAND U1030 ( .A(n1177), .B(n1178), .Z(n1175) );
  NANDN U1031 ( .A(B[218]), .B(A[218]), .Z(n1178) );
  AND U1032 ( .A(n1179), .B(n1180), .Z(n1177) );
  NAND U1033 ( .A(n1181), .B(n1182), .Z(n1180) );
  NANDN U1034 ( .A(A[217]), .B(B[217]), .Z(n1182) );
  AND U1035 ( .A(n1183), .B(n1184), .Z(n1181) );
  NANDN U1036 ( .A(A[216]), .B(B[216]), .Z(n1184) );
  NAND U1037 ( .A(n1185), .B(n1186), .Z(n1183) );
  NANDN U1038 ( .A(B[216]), .B(A[216]), .Z(n1186) );
  AND U1039 ( .A(n1187), .B(n1188), .Z(n1185) );
  NAND U1040 ( .A(n1189), .B(n1190), .Z(n1188) );
  NANDN U1041 ( .A(A[215]), .B(B[215]), .Z(n1190) );
  AND U1042 ( .A(n1191), .B(n1192), .Z(n1189) );
  NANDN U1043 ( .A(A[214]), .B(B[214]), .Z(n1192) );
  NAND U1044 ( .A(n1193), .B(n1194), .Z(n1191) );
  NANDN U1045 ( .A(B[214]), .B(A[214]), .Z(n1194) );
  AND U1046 ( .A(n1195), .B(n1196), .Z(n1193) );
  NAND U1047 ( .A(n1197), .B(n1198), .Z(n1196) );
  NANDN U1048 ( .A(A[213]), .B(B[213]), .Z(n1198) );
  AND U1049 ( .A(n1199), .B(n1200), .Z(n1197) );
  NANDN U1050 ( .A(A[212]), .B(B[212]), .Z(n1200) );
  NAND U1051 ( .A(n1201), .B(n1202), .Z(n1199) );
  NANDN U1052 ( .A(B[212]), .B(A[212]), .Z(n1202) );
  AND U1053 ( .A(n1203), .B(n1204), .Z(n1201) );
  NAND U1054 ( .A(n1205), .B(n1206), .Z(n1204) );
  NANDN U1055 ( .A(A[211]), .B(B[211]), .Z(n1206) );
  AND U1056 ( .A(n1207), .B(n1208), .Z(n1205) );
  NANDN U1057 ( .A(A[210]), .B(B[210]), .Z(n1208) );
  NAND U1058 ( .A(n1209), .B(n1210), .Z(n1207) );
  NANDN U1059 ( .A(B[210]), .B(A[210]), .Z(n1210) );
  AND U1060 ( .A(n1211), .B(n1212), .Z(n1209) );
  NAND U1061 ( .A(n1213), .B(n1214), .Z(n1212) );
  NANDN U1062 ( .A(A[209]), .B(B[209]), .Z(n1214) );
  AND U1063 ( .A(n1215), .B(n1216), .Z(n1213) );
  NANDN U1064 ( .A(A[208]), .B(B[208]), .Z(n1216) );
  NAND U1065 ( .A(n1217), .B(n1218), .Z(n1215) );
  NANDN U1066 ( .A(B[208]), .B(A[208]), .Z(n1218) );
  AND U1067 ( .A(n1219), .B(n1220), .Z(n1217) );
  NAND U1068 ( .A(n1221), .B(n1222), .Z(n1220) );
  NANDN U1069 ( .A(A[207]), .B(B[207]), .Z(n1222) );
  AND U1070 ( .A(n1223), .B(n1224), .Z(n1221) );
  NANDN U1071 ( .A(A[206]), .B(B[206]), .Z(n1224) );
  NAND U1072 ( .A(n1225), .B(n1226), .Z(n1223) );
  NANDN U1073 ( .A(B[206]), .B(A[206]), .Z(n1226) );
  AND U1074 ( .A(n1227), .B(n1228), .Z(n1225) );
  NAND U1075 ( .A(n1229), .B(n1230), .Z(n1228) );
  NANDN U1076 ( .A(A[205]), .B(B[205]), .Z(n1230) );
  AND U1077 ( .A(n1231), .B(n1232), .Z(n1229) );
  NANDN U1078 ( .A(A[204]), .B(B[204]), .Z(n1232) );
  NAND U1079 ( .A(n1233), .B(n1234), .Z(n1231) );
  NANDN U1080 ( .A(B[204]), .B(A[204]), .Z(n1234) );
  AND U1081 ( .A(n1235), .B(n1236), .Z(n1233) );
  NAND U1082 ( .A(n1237), .B(n1238), .Z(n1236) );
  NANDN U1083 ( .A(A[203]), .B(B[203]), .Z(n1238) );
  AND U1084 ( .A(n1239), .B(n1240), .Z(n1237) );
  NANDN U1085 ( .A(A[202]), .B(B[202]), .Z(n1240) );
  NAND U1086 ( .A(n1241), .B(n1242), .Z(n1239) );
  NANDN U1087 ( .A(B[202]), .B(A[202]), .Z(n1242) );
  AND U1088 ( .A(n1243), .B(n1244), .Z(n1241) );
  NAND U1089 ( .A(n1245), .B(n1246), .Z(n1244) );
  NANDN U1090 ( .A(A[201]), .B(B[201]), .Z(n1246) );
  AND U1091 ( .A(n1247), .B(n1248), .Z(n1245) );
  NANDN U1092 ( .A(A[200]), .B(B[200]), .Z(n1248) );
  NAND U1093 ( .A(n1249), .B(n1250), .Z(n1247) );
  NANDN U1094 ( .A(B[200]), .B(A[200]), .Z(n1250) );
  AND U1095 ( .A(n1251), .B(n1252), .Z(n1249) );
  NAND U1096 ( .A(n1253), .B(n1254), .Z(n1252) );
  NANDN U1097 ( .A(A[199]), .B(B[199]), .Z(n1254) );
  AND U1098 ( .A(n1255), .B(n1256), .Z(n1253) );
  NANDN U1099 ( .A(A[198]), .B(B[198]), .Z(n1256) );
  NAND U1100 ( .A(n1257), .B(n1258), .Z(n1255) );
  NANDN U1101 ( .A(B[198]), .B(A[198]), .Z(n1258) );
  AND U1102 ( .A(n1259), .B(n1260), .Z(n1257) );
  NAND U1103 ( .A(n1261), .B(n1262), .Z(n1260) );
  NANDN U1104 ( .A(A[197]), .B(B[197]), .Z(n1262) );
  AND U1105 ( .A(n1263), .B(n1264), .Z(n1261) );
  NANDN U1106 ( .A(A[196]), .B(B[196]), .Z(n1264) );
  NAND U1107 ( .A(n1265), .B(n1266), .Z(n1263) );
  NANDN U1108 ( .A(B[196]), .B(A[196]), .Z(n1266) );
  AND U1109 ( .A(n1267), .B(n1268), .Z(n1265) );
  NAND U1110 ( .A(n1269), .B(n1270), .Z(n1268) );
  NANDN U1111 ( .A(A[195]), .B(B[195]), .Z(n1270) );
  AND U1112 ( .A(n1271), .B(n1272), .Z(n1269) );
  NANDN U1113 ( .A(A[194]), .B(B[194]), .Z(n1272) );
  NAND U1114 ( .A(n1273), .B(n1274), .Z(n1271) );
  NANDN U1115 ( .A(B[194]), .B(A[194]), .Z(n1274) );
  AND U1116 ( .A(n1275), .B(n1276), .Z(n1273) );
  NAND U1117 ( .A(n1277), .B(n1278), .Z(n1276) );
  NANDN U1118 ( .A(A[193]), .B(B[193]), .Z(n1278) );
  AND U1119 ( .A(n1279), .B(n1280), .Z(n1277) );
  NANDN U1120 ( .A(A[192]), .B(B[192]), .Z(n1280) );
  NAND U1121 ( .A(n1281), .B(n1282), .Z(n1279) );
  NANDN U1122 ( .A(B[192]), .B(A[192]), .Z(n1282) );
  AND U1123 ( .A(n1283), .B(n1284), .Z(n1281) );
  NAND U1124 ( .A(n1285), .B(n1286), .Z(n1284) );
  NANDN U1125 ( .A(A[191]), .B(B[191]), .Z(n1286) );
  AND U1126 ( .A(n1287), .B(n1288), .Z(n1285) );
  NANDN U1127 ( .A(A[190]), .B(B[190]), .Z(n1288) );
  NAND U1128 ( .A(n1289), .B(n1290), .Z(n1287) );
  NANDN U1129 ( .A(B[190]), .B(A[190]), .Z(n1290) );
  AND U1130 ( .A(n1291), .B(n1292), .Z(n1289) );
  NAND U1131 ( .A(n1293), .B(n1294), .Z(n1292) );
  NANDN U1132 ( .A(A[189]), .B(B[189]), .Z(n1294) );
  AND U1133 ( .A(n1295), .B(n1296), .Z(n1293) );
  NANDN U1134 ( .A(A[188]), .B(B[188]), .Z(n1296) );
  NAND U1135 ( .A(n1297), .B(n1298), .Z(n1295) );
  NANDN U1136 ( .A(B[188]), .B(A[188]), .Z(n1298) );
  AND U1137 ( .A(n1299), .B(n1300), .Z(n1297) );
  NAND U1138 ( .A(n1301), .B(n1302), .Z(n1300) );
  NANDN U1139 ( .A(A[187]), .B(B[187]), .Z(n1302) );
  AND U1140 ( .A(n1303), .B(n1304), .Z(n1301) );
  NANDN U1141 ( .A(A[186]), .B(B[186]), .Z(n1304) );
  NAND U1142 ( .A(n1305), .B(n1306), .Z(n1303) );
  NANDN U1143 ( .A(B[186]), .B(A[186]), .Z(n1306) );
  AND U1144 ( .A(n1307), .B(n1308), .Z(n1305) );
  NAND U1145 ( .A(n1309), .B(n1310), .Z(n1308) );
  NANDN U1146 ( .A(A[185]), .B(B[185]), .Z(n1310) );
  AND U1147 ( .A(n1311), .B(n1312), .Z(n1309) );
  NANDN U1148 ( .A(A[184]), .B(B[184]), .Z(n1312) );
  NAND U1149 ( .A(n1313), .B(n1314), .Z(n1311) );
  NANDN U1150 ( .A(B[184]), .B(A[184]), .Z(n1314) );
  AND U1151 ( .A(n1315), .B(n1316), .Z(n1313) );
  NAND U1152 ( .A(n1317), .B(n1318), .Z(n1316) );
  NANDN U1153 ( .A(A[183]), .B(B[183]), .Z(n1318) );
  AND U1154 ( .A(n1319), .B(n1320), .Z(n1317) );
  NANDN U1155 ( .A(A[182]), .B(B[182]), .Z(n1320) );
  NAND U1156 ( .A(n1321), .B(n1322), .Z(n1319) );
  NANDN U1157 ( .A(B[182]), .B(A[182]), .Z(n1322) );
  AND U1158 ( .A(n1323), .B(n1324), .Z(n1321) );
  NAND U1159 ( .A(n1325), .B(n1326), .Z(n1324) );
  NANDN U1160 ( .A(A[181]), .B(B[181]), .Z(n1326) );
  AND U1161 ( .A(n1327), .B(n1328), .Z(n1325) );
  NANDN U1162 ( .A(A[180]), .B(B[180]), .Z(n1328) );
  NAND U1163 ( .A(n1329), .B(n1330), .Z(n1327) );
  NANDN U1164 ( .A(B[180]), .B(A[180]), .Z(n1330) );
  AND U1165 ( .A(n1331), .B(n1332), .Z(n1329) );
  NAND U1166 ( .A(n1333), .B(n1334), .Z(n1332) );
  NANDN U1167 ( .A(A[179]), .B(B[179]), .Z(n1334) );
  AND U1168 ( .A(n1335), .B(n1336), .Z(n1333) );
  NANDN U1169 ( .A(A[178]), .B(B[178]), .Z(n1336) );
  NAND U1170 ( .A(n1337), .B(n1338), .Z(n1335) );
  NANDN U1171 ( .A(B[178]), .B(A[178]), .Z(n1338) );
  AND U1172 ( .A(n1339), .B(n1340), .Z(n1337) );
  NAND U1173 ( .A(n1341), .B(n1342), .Z(n1340) );
  NANDN U1174 ( .A(A[177]), .B(B[177]), .Z(n1342) );
  AND U1175 ( .A(n1343), .B(n1344), .Z(n1341) );
  NANDN U1176 ( .A(A[176]), .B(B[176]), .Z(n1344) );
  NAND U1177 ( .A(n1345), .B(n1346), .Z(n1343) );
  NANDN U1178 ( .A(B[176]), .B(A[176]), .Z(n1346) );
  AND U1179 ( .A(n1347), .B(n1348), .Z(n1345) );
  NAND U1180 ( .A(n1349), .B(n1350), .Z(n1348) );
  NANDN U1181 ( .A(A[175]), .B(B[175]), .Z(n1350) );
  AND U1182 ( .A(n1351), .B(n1352), .Z(n1349) );
  NANDN U1183 ( .A(A[174]), .B(B[174]), .Z(n1352) );
  NAND U1184 ( .A(n1353), .B(n1354), .Z(n1351) );
  NANDN U1185 ( .A(B[174]), .B(A[174]), .Z(n1354) );
  AND U1186 ( .A(n1355), .B(n1356), .Z(n1353) );
  NAND U1187 ( .A(n1357), .B(n1358), .Z(n1356) );
  NANDN U1188 ( .A(A[173]), .B(B[173]), .Z(n1358) );
  AND U1189 ( .A(n1359), .B(n1360), .Z(n1357) );
  NANDN U1190 ( .A(A[172]), .B(B[172]), .Z(n1360) );
  NAND U1191 ( .A(n1361), .B(n1362), .Z(n1359) );
  NANDN U1192 ( .A(B[172]), .B(A[172]), .Z(n1362) );
  AND U1193 ( .A(n1363), .B(n1364), .Z(n1361) );
  NAND U1194 ( .A(n1365), .B(n1366), .Z(n1364) );
  NANDN U1195 ( .A(A[171]), .B(B[171]), .Z(n1366) );
  AND U1196 ( .A(n1367), .B(n1368), .Z(n1365) );
  NANDN U1197 ( .A(A[170]), .B(B[170]), .Z(n1368) );
  NAND U1198 ( .A(n1369), .B(n1370), .Z(n1367) );
  NANDN U1199 ( .A(B[170]), .B(A[170]), .Z(n1370) );
  AND U1200 ( .A(n1371), .B(n1372), .Z(n1369) );
  NAND U1201 ( .A(n1373), .B(n1374), .Z(n1372) );
  NANDN U1202 ( .A(A[169]), .B(B[169]), .Z(n1374) );
  AND U1203 ( .A(n1375), .B(n1376), .Z(n1373) );
  NANDN U1204 ( .A(A[168]), .B(B[168]), .Z(n1376) );
  NAND U1205 ( .A(n1377), .B(n1378), .Z(n1375) );
  NANDN U1206 ( .A(B[168]), .B(A[168]), .Z(n1378) );
  AND U1207 ( .A(n1379), .B(n1380), .Z(n1377) );
  NAND U1208 ( .A(n1381), .B(n1382), .Z(n1380) );
  NANDN U1209 ( .A(A[167]), .B(B[167]), .Z(n1382) );
  AND U1210 ( .A(n1383), .B(n1384), .Z(n1381) );
  NANDN U1211 ( .A(A[166]), .B(B[166]), .Z(n1384) );
  NAND U1212 ( .A(n1385), .B(n1386), .Z(n1383) );
  NANDN U1213 ( .A(B[166]), .B(A[166]), .Z(n1386) );
  AND U1214 ( .A(n1387), .B(n1388), .Z(n1385) );
  NAND U1215 ( .A(n1389), .B(n1390), .Z(n1388) );
  NANDN U1216 ( .A(A[165]), .B(B[165]), .Z(n1390) );
  AND U1217 ( .A(n1391), .B(n1392), .Z(n1389) );
  NANDN U1218 ( .A(A[164]), .B(B[164]), .Z(n1392) );
  NAND U1219 ( .A(n1393), .B(n1394), .Z(n1391) );
  NANDN U1220 ( .A(B[164]), .B(A[164]), .Z(n1394) );
  AND U1221 ( .A(n1395), .B(n1396), .Z(n1393) );
  NAND U1222 ( .A(n1397), .B(n1398), .Z(n1396) );
  NANDN U1223 ( .A(A[163]), .B(B[163]), .Z(n1398) );
  AND U1224 ( .A(n1399), .B(n1400), .Z(n1397) );
  NANDN U1225 ( .A(A[162]), .B(B[162]), .Z(n1400) );
  NAND U1226 ( .A(n1401), .B(n1402), .Z(n1399) );
  NANDN U1227 ( .A(B[162]), .B(A[162]), .Z(n1402) );
  AND U1228 ( .A(n1403), .B(n1404), .Z(n1401) );
  NAND U1229 ( .A(n1405), .B(n1406), .Z(n1404) );
  NANDN U1230 ( .A(A[161]), .B(B[161]), .Z(n1406) );
  AND U1231 ( .A(n1407), .B(n1408), .Z(n1405) );
  NANDN U1232 ( .A(A[160]), .B(B[160]), .Z(n1408) );
  NAND U1233 ( .A(n1409), .B(n1410), .Z(n1407) );
  NANDN U1234 ( .A(B[160]), .B(A[160]), .Z(n1410) );
  AND U1235 ( .A(n1411), .B(n1412), .Z(n1409) );
  NAND U1236 ( .A(n1413), .B(n1414), .Z(n1412) );
  NANDN U1237 ( .A(A[159]), .B(B[159]), .Z(n1414) );
  AND U1238 ( .A(n1415), .B(n1416), .Z(n1413) );
  NANDN U1239 ( .A(A[158]), .B(B[158]), .Z(n1416) );
  NAND U1240 ( .A(n1417), .B(n1418), .Z(n1415) );
  NANDN U1241 ( .A(B[158]), .B(A[158]), .Z(n1418) );
  AND U1242 ( .A(n1419), .B(n1420), .Z(n1417) );
  NAND U1243 ( .A(n1421), .B(n1422), .Z(n1420) );
  NANDN U1244 ( .A(A[157]), .B(B[157]), .Z(n1422) );
  AND U1245 ( .A(n1423), .B(n1424), .Z(n1421) );
  NANDN U1246 ( .A(A[156]), .B(B[156]), .Z(n1424) );
  NAND U1247 ( .A(n1425), .B(n1426), .Z(n1423) );
  NANDN U1248 ( .A(B[156]), .B(A[156]), .Z(n1426) );
  AND U1249 ( .A(n1427), .B(n1428), .Z(n1425) );
  NAND U1250 ( .A(n1429), .B(n1430), .Z(n1428) );
  NANDN U1251 ( .A(A[155]), .B(B[155]), .Z(n1430) );
  AND U1252 ( .A(n1431), .B(n1432), .Z(n1429) );
  NANDN U1253 ( .A(A[154]), .B(B[154]), .Z(n1432) );
  NAND U1254 ( .A(n1433), .B(n1434), .Z(n1431) );
  NANDN U1255 ( .A(B[154]), .B(A[154]), .Z(n1434) );
  AND U1256 ( .A(n1435), .B(n1436), .Z(n1433) );
  NAND U1257 ( .A(n1437), .B(n1438), .Z(n1436) );
  NANDN U1258 ( .A(A[153]), .B(B[153]), .Z(n1438) );
  AND U1259 ( .A(n1439), .B(n1440), .Z(n1437) );
  NANDN U1260 ( .A(A[152]), .B(B[152]), .Z(n1440) );
  NAND U1261 ( .A(n1441), .B(n1442), .Z(n1439) );
  NANDN U1262 ( .A(B[152]), .B(A[152]), .Z(n1442) );
  AND U1263 ( .A(n1443), .B(n1444), .Z(n1441) );
  NAND U1264 ( .A(n1445), .B(n1446), .Z(n1444) );
  NANDN U1265 ( .A(A[151]), .B(B[151]), .Z(n1446) );
  AND U1266 ( .A(n1447), .B(n1448), .Z(n1445) );
  NANDN U1267 ( .A(A[150]), .B(B[150]), .Z(n1448) );
  NAND U1268 ( .A(n1449), .B(n1450), .Z(n1447) );
  NANDN U1269 ( .A(B[150]), .B(A[150]), .Z(n1450) );
  AND U1270 ( .A(n1451), .B(n1452), .Z(n1449) );
  NAND U1271 ( .A(n1453), .B(n1454), .Z(n1452) );
  NANDN U1272 ( .A(A[149]), .B(B[149]), .Z(n1454) );
  AND U1273 ( .A(n1455), .B(n1456), .Z(n1453) );
  NANDN U1274 ( .A(A[148]), .B(B[148]), .Z(n1456) );
  NAND U1275 ( .A(n1457), .B(n1458), .Z(n1455) );
  NANDN U1276 ( .A(B[148]), .B(A[148]), .Z(n1458) );
  AND U1277 ( .A(n1459), .B(n1460), .Z(n1457) );
  NAND U1278 ( .A(n1461), .B(n1462), .Z(n1460) );
  NANDN U1279 ( .A(A[147]), .B(B[147]), .Z(n1462) );
  AND U1280 ( .A(n1463), .B(n1464), .Z(n1461) );
  NANDN U1281 ( .A(A[146]), .B(B[146]), .Z(n1464) );
  NAND U1282 ( .A(n1465), .B(n1466), .Z(n1463) );
  NANDN U1283 ( .A(B[146]), .B(A[146]), .Z(n1466) );
  AND U1284 ( .A(n1467), .B(n1468), .Z(n1465) );
  NAND U1285 ( .A(n1469), .B(n1470), .Z(n1468) );
  NANDN U1286 ( .A(A[145]), .B(B[145]), .Z(n1470) );
  AND U1287 ( .A(n1471), .B(n1472), .Z(n1469) );
  NANDN U1288 ( .A(A[144]), .B(B[144]), .Z(n1472) );
  NAND U1289 ( .A(n1473), .B(n1474), .Z(n1471) );
  NANDN U1290 ( .A(B[144]), .B(A[144]), .Z(n1474) );
  AND U1291 ( .A(n1475), .B(n1476), .Z(n1473) );
  NAND U1292 ( .A(n1477), .B(n1478), .Z(n1476) );
  NANDN U1293 ( .A(A[143]), .B(B[143]), .Z(n1478) );
  AND U1294 ( .A(n1479), .B(n1480), .Z(n1477) );
  NANDN U1295 ( .A(A[142]), .B(B[142]), .Z(n1480) );
  NAND U1296 ( .A(n1481), .B(n1482), .Z(n1479) );
  NANDN U1297 ( .A(B[142]), .B(A[142]), .Z(n1482) );
  AND U1298 ( .A(n1483), .B(n1484), .Z(n1481) );
  NAND U1299 ( .A(n1485), .B(n1486), .Z(n1484) );
  NANDN U1300 ( .A(A[141]), .B(B[141]), .Z(n1486) );
  AND U1301 ( .A(n1487), .B(n1488), .Z(n1485) );
  NANDN U1302 ( .A(A[140]), .B(B[140]), .Z(n1488) );
  NAND U1303 ( .A(n1489), .B(n1490), .Z(n1487) );
  NANDN U1304 ( .A(B[140]), .B(A[140]), .Z(n1490) );
  AND U1305 ( .A(n1491), .B(n1492), .Z(n1489) );
  NAND U1306 ( .A(n1493), .B(n1494), .Z(n1492) );
  NANDN U1307 ( .A(A[139]), .B(B[139]), .Z(n1494) );
  AND U1308 ( .A(n1495), .B(n1496), .Z(n1493) );
  NANDN U1309 ( .A(A[138]), .B(B[138]), .Z(n1496) );
  NAND U1310 ( .A(n1497), .B(n1498), .Z(n1495) );
  NANDN U1311 ( .A(B[138]), .B(A[138]), .Z(n1498) );
  AND U1312 ( .A(n1499), .B(n1500), .Z(n1497) );
  NAND U1313 ( .A(n1501), .B(n1502), .Z(n1500) );
  NANDN U1314 ( .A(A[137]), .B(B[137]), .Z(n1502) );
  AND U1315 ( .A(n1503), .B(n1504), .Z(n1501) );
  NANDN U1316 ( .A(A[136]), .B(B[136]), .Z(n1504) );
  NAND U1317 ( .A(n1505), .B(n1506), .Z(n1503) );
  NANDN U1318 ( .A(B[136]), .B(A[136]), .Z(n1506) );
  AND U1319 ( .A(n1507), .B(n1508), .Z(n1505) );
  NAND U1320 ( .A(n1509), .B(n1510), .Z(n1508) );
  NANDN U1321 ( .A(A[135]), .B(B[135]), .Z(n1510) );
  AND U1322 ( .A(n1511), .B(n1512), .Z(n1509) );
  NANDN U1323 ( .A(A[134]), .B(B[134]), .Z(n1512) );
  NAND U1324 ( .A(n1513), .B(n1514), .Z(n1511) );
  NANDN U1325 ( .A(B[134]), .B(A[134]), .Z(n1514) );
  AND U1326 ( .A(n1515), .B(n1516), .Z(n1513) );
  NAND U1327 ( .A(n1517), .B(n1518), .Z(n1516) );
  NANDN U1328 ( .A(A[133]), .B(B[133]), .Z(n1518) );
  AND U1329 ( .A(n1519), .B(n1520), .Z(n1517) );
  NANDN U1330 ( .A(A[132]), .B(B[132]), .Z(n1520) );
  NAND U1331 ( .A(n1521), .B(n1522), .Z(n1519) );
  NANDN U1332 ( .A(B[132]), .B(A[132]), .Z(n1522) );
  AND U1333 ( .A(n1523), .B(n1524), .Z(n1521) );
  NAND U1334 ( .A(n1525), .B(n1526), .Z(n1524) );
  NANDN U1335 ( .A(A[131]), .B(B[131]), .Z(n1526) );
  AND U1336 ( .A(n1527), .B(n1528), .Z(n1525) );
  NANDN U1337 ( .A(A[130]), .B(B[130]), .Z(n1528) );
  NAND U1338 ( .A(n1529), .B(n1530), .Z(n1527) );
  NANDN U1339 ( .A(B[130]), .B(A[130]), .Z(n1530) );
  AND U1340 ( .A(n1531), .B(n1532), .Z(n1529) );
  NAND U1341 ( .A(n1533), .B(n1534), .Z(n1532) );
  NANDN U1342 ( .A(A[129]), .B(B[129]), .Z(n1534) );
  AND U1343 ( .A(n1535), .B(n1536), .Z(n1533) );
  NANDN U1344 ( .A(A[128]), .B(B[128]), .Z(n1536) );
  NAND U1345 ( .A(n1537), .B(n1538), .Z(n1535) );
  NANDN U1346 ( .A(B[128]), .B(A[128]), .Z(n1538) );
  AND U1347 ( .A(n1539), .B(n1540), .Z(n1537) );
  NAND U1348 ( .A(n1541), .B(n1542), .Z(n1540) );
  NANDN U1349 ( .A(A[127]), .B(B[127]), .Z(n1542) );
  AND U1350 ( .A(n1543), .B(n1544), .Z(n1541) );
  NANDN U1351 ( .A(A[126]), .B(B[126]), .Z(n1544) );
  NAND U1352 ( .A(n1545), .B(n1546), .Z(n1543) );
  NANDN U1353 ( .A(B[126]), .B(A[126]), .Z(n1546) );
  AND U1354 ( .A(n1547), .B(n1548), .Z(n1545) );
  NAND U1355 ( .A(n1549), .B(n1550), .Z(n1548) );
  NANDN U1356 ( .A(A[125]), .B(B[125]), .Z(n1550) );
  AND U1357 ( .A(n1551), .B(n1552), .Z(n1549) );
  NANDN U1358 ( .A(A[124]), .B(B[124]), .Z(n1552) );
  NAND U1359 ( .A(n1553), .B(n1554), .Z(n1551) );
  NANDN U1360 ( .A(B[124]), .B(A[124]), .Z(n1554) );
  AND U1361 ( .A(n1555), .B(n1556), .Z(n1553) );
  NAND U1362 ( .A(n1557), .B(n1558), .Z(n1556) );
  NANDN U1363 ( .A(A[123]), .B(B[123]), .Z(n1558) );
  AND U1364 ( .A(n1559), .B(n1560), .Z(n1557) );
  NANDN U1365 ( .A(A[122]), .B(B[122]), .Z(n1560) );
  NAND U1366 ( .A(n1561), .B(n1562), .Z(n1559) );
  NANDN U1367 ( .A(B[122]), .B(A[122]), .Z(n1562) );
  AND U1368 ( .A(n1563), .B(n1564), .Z(n1561) );
  NAND U1369 ( .A(n1565), .B(n1566), .Z(n1564) );
  NANDN U1370 ( .A(A[121]), .B(B[121]), .Z(n1566) );
  AND U1371 ( .A(n1567), .B(n1568), .Z(n1565) );
  NANDN U1372 ( .A(A[120]), .B(B[120]), .Z(n1568) );
  NAND U1373 ( .A(n1569), .B(n1570), .Z(n1567) );
  NANDN U1374 ( .A(B[120]), .B(A[120]), .Z(n1570) );
  AND U1375 ( .A(n1571), .B(n1572), .Z(n1569) );
  NAND U1376 ( .A(n1573), .B(n1574), .Z(n1572) );
  NANDN U1377 ( .A(A[119]), .B(B[119]), .Z(n1574) );
  AND U1378 ( .A(n1575), .B(n1576), .Z(n1573) );
  NANDN U1379 ( .A(A[118]), .B(B[118]), .Z(n1576) );
  NAND U1380 ( .A(n1577), .B(n1578), .Z(n1575) );
  NANDN U1381 ( .A(B[118]), .B(A[118]), .Z(n1578) );
  AND U1382 ( .A(n1579), .B(n1580), .Z(n1577) );
  NAND U1383 ( .A(n1581), .B(n1582), .Z(n1580) );
  NANDN U1384 ( .A(A[117]), .B(B[117]), .Z(n1582) );
  AND U1385 ( .A(n1583), .B(n1584), .Z(n1581) );
  NANDN U1386 ( .A(A[116]), .B(B[116]), .Z(n1584) );
  NAND U1387 ( .A(n1585), .B(n1586), .Z(n1583) );
  NANDN U1388 ( .A(B[116]), .B(A[116]), .Z(n1586) );
  AND U1389 ( .A(n1587), .B(n1588), .Z(n1585) );
  NAND U1390 ( .A(n1589), .B(n1590), .Z(n1588) );
  NANDN U1391 ( .A(A[115]), .B(B[115]), .Z(n1590) );
  AND U1392 ( .A(n1591), .B(n1592), .Z(n1589) );
  NANDN U1393 ( .A(A[114]), .B(B[114]), .Z(n1592) );
  NAND U1394 ( .A(n1593), .B(n1594), .Z(n1591) );
  NANDN U1395 ( .A(B[114]), .B(A[114]), .Z(n1594) );
  AND U1396 ( .A(n1595), .B(n1596), .Z(n1593) );
  NAND U1397 ( .A(n1597), .B(n1598), .Z(n1596) );
  NANDN U1398 ( .A(A[113]), .B(B[113]), .Z(n1598) );
  AND U1399 ( .A(n1599), .B(n1600), .Z(n1597) );
  NANDN U1400 ( .A(A[112]), .B(B[112]), .Z(n1600) );
  NAND U1401 ( .A(n1601), .B(n1602), .Z(n1599) );
  NANDN U1402 ( .A(B[112]), .B(A[112]), .Z(n1602) );
  AND U1403 ( .A(n1603), .B(n1604), .Z(n1601) );
  NAND U1404 ( .A(n1605), .B(n1606), .Z(n1604) );
  NANDN U1405 ( .A(A[111]), .B(B[111]), .Z(n1606) );
  AND U1406 ( .A(n1607), .B(n1608), .Z(n1605) );
  NANDN U1407 ( .A(A[110]), .B(B[110]), .Z(n1608) );
  NAND U1408 ( .A(n1609), .B(n1610), .Z(n1607) );
  NANDN U1409 ( .A(B[110]), .B(A[110]), .Z(n1610) );
  AND U1410 ( .A(n1611), .B(n1612), .Z(n1609) );
  NAND U1411 ( .A(n1613), .B(n1614), .Z(n1612) );
  NANDN U1412 ( .A(A[109]), .B(B[109]), .Z(n1614) );
  AND U1413 ( .A(n1615), .B(n1616), .Z(n1613) );
  NANDN U1414 ( .A(A[108]), .B(B[108]), .Z(n1616) );
  NAND U1415 ( .A(n1617), .B(n1618), .Z(n1615) );
  NANDN U1416 ( .A(B[108]), .B(A[108]), .Z(n1618) );
  AND U1417 ( .A(n1619), .B(n1620), .Z(n1617) );
  NAND U1418 ( .A(n1621), .B(n1622), .Z(n1620) );
  NANDN U1419 ( .A(A[107]), .B(B[107]), .Z(n1622) );
  AND U1420 ( .A(n1623), .B(n1624), .Z(n1621) );
  NANDN U1421 ( .A(A[106]), .B(B[106]), .Z(n1624) );
  NAND U1422 ( .A(n1625), .B(n1626), .Z(n1623) );
  NANDN U1423 ( .A(B[106]), .B(A[106]), .Z(n1626) );
  AND U1424 ( .A(n1627), .B(n1628), .Z(n1625) );
  NAND U1425 ( .A(n1629), .B(n1630), .Z(n1628) );
  NANDN U1426 ( .A(A[105]), .B(B[105]), .Z(n1630) );
  AND U1427 ( .A(n1631), .B(n1632), .Z(n1629) );
  NANDN U1428 ( .A(A[104]), .B(B[104]), .Z(n1632) );
  NAND U1429 ( .A(n1633), .B(n1634), .Z(n1631) );
  NANDN U1430 ( .A(B[104]), .B(A[104]), .Z(n1634) );
  AND U1431 ( .A(n1635), .B(n1636), .Z(n1633) );
  NAND U1432 ( .A(n1637), .B(n1638), .Z(n1636) );
  NANDN U1433 ( .A(A[103]), .B(B[103]), .Z(n1638) );
  AND U1434 ( .A(n1639), .B(n1640), .Z(n1637) );
  NANDN U1435 ( .A(A[102]), .B(B[102]), .Z(n1640) );
  NAND U1436 ( .A(n1641), .B(n1642), .Z(n1639) );
  NANDN U1437 ( .A(B[102]), .B(A[102]), .Z(n1642) );
  AND U1438 ( .A(n1643), .B(n1644), .Z(n1641) );
  NAND U1439 ( .A(n1645), .B(n1646), .Z(n1644) );
  NANDN U1440 ( .A(A[101]), .B(B[101]), .Z(n1646) );
  AND U1441 ( .A(n1647), .B(n1648), .Z(n1645) );
  NANDN U1442 ( .A(A[100]), .B(B[100]), .Z(n1648) );
  NAND U1443 ( .A(n1649), .B(n1650), .Z(n1647) );
  NANDN U1444 ( .A(B[99]), .B(A[99]), .Z(n1650) );
  AND U1445 ( .A(n1651), .B(n1652), .Z(n1649) );
  NAND U1446 ( .A(n1653), .B(n1654), .Z(n1652) );
  NANDN U1447 ( .A(A[99]), .B(B[99]), .Z(n1654) );
  AND U1448 ( .A(n1655), .B(n1656), .Z(n1653) );
  NANDN U1449 ( .A(A[98]), .B(B[98]), .Z(n1656) );
  NAND U1450 ( .A(n1657), .B(n1658), .Z(n1655) );
  NANDN U1451 ( .A(B[98]), .B(A[98]), .Z(n1658) );
  AND U1452 ( .A(n1659), .B(n1660), .Z(n1657) );
  NAND U1453 ( .A(n1661), .B(n1662), .Z(n1660) );
  NANDN U1454 ( .A(A[97]), .B(B[97]), .Z(n1662) );
  AND U1455 ( .A(n1663), .B(n1664), .Z(n1661) );
  NANDN U1456 ( .A(A[96]), .B(B[96]), .Z(n1664) );
  NAND U1457 ( .A(n1665), .B(n1666), .Z(n1663) );
  NANDN U1458 ( .A(B[96]), .B(A[96]), .Z(n1666) );
  AND U1459 ( .A(n1667), .B(n1668), .Z(n1665) );
  NAND U1460 ( .A(n1669), .B(n1670), .Z(n1668) );
  NANDN U1461 ( .A(A[95]), .B(B[95]), .Z(n1670) );
  AND U1462 ( .A(n1671), .B(n1672), .Z(n1669) );
  NANDN U1463 ( .A(A[94]), .B(B[94]), .Z(n1672) );
  NAND U1464 ( .A(n1673), .B(n1674), .Z(n1671) );
  NANDN U1465 ( .A(B[94]), .B(A[94]), .Z(n1674) );
  AND U1466 ( .A(n1675), .B(n1676), .Z(n1673) );
  NAND U1467 ( .A(n1677), .B(n1678), .Z(n1676) );
  NANDN U1468 ( .A(A[93]), .B(B[93]), .Z(n1678) );
  AND U1469 ( .A(n1679), .B(n1680), .Z(n1677) );
  NANDN U1470 ( .A(A[92]), .B(B[92]), .Z(n1680) );
  NAND U1471 ( .A(n1681), .B(n1682), .Z(n1679) );
  NANDN U1472 ( .A(B[92]), .B(A[92]), .Z(n1682) );
  AND U1473 ( .A(n1683), .B(n1684), .Z(n1681) );
  NAND U1474 ( .A(n1685), .B(n1686), .Z(n1684) );
  NANDN U1475 ( .A(A[91]), .B(B[91]), .Z(n1686) );
  AND U1476 ( .A(n1687), .B(n1688), .Z(n1685) );
  NANDN U1477 ( .A(A[90]), .B(B[90]), .Z(n1688) );
  NAND U1478 ( .A(n1689), .B(n1690), .Z(n1687) );
  NANDN U1479 ( .A(B[90]), .B(A[90]), .Z(n1690) );
  AND U1480 ( .A(n1691), .B(n1692), .Z(n1689) );
  NAND U1481 ( .A(n1693), .B(n1694), .Z(n1692) );
  NANDN U1482 ( .A(A[89]), .B(B[89]), .Z(n1694) );
  AND U1483 ( .A(n1695), .B(n1696), .Z(n1693) );
  NANDN U1484 ( .A(A[88]), .B(B[88]), .Z(n1696) );
  NAND U1485 ( .A(n1697), .B(n1698), .Z(n1695) );
  NANDN U1486 ( .A(B[88]), .B(A[88]), .Z(n1698) );
  AND U1487 ( .A(n1699), .B(n1700), .Z(n1697) );
  NAND U1488 ( .A(n1701), .B(n1702), .Z(n1700) );
  NANDN U1489 ( .A(A[87]), .B(B[87]), .Z(n1702) );
  AND U1490 ( .A(n1703), .B(n1704), .Z(n1701) );
  NANDN U1491 ( .A(A[86]), .B(B[86]), .Z(n1704) );
  NAND U1492 ( .A(n1705), .B(n1706), .Z(n1703) );
  NANDN U1493 ( .A(B[86]), .B(A[86]), .Z(n1706) );
  AND U1494 ( .A(n1707), .B(n1708), .Z(n1705) );
  NAND U1495 ( .A(n1709), .B(n1710), .Z(n1708) );
  NANDN U1496 ( .A(A[85]), .B(B[85]), .Z(n1710) );
  AND U1497 ( .A(n1711), .B(n1712), .Z(n1709) );
  NANDN U1498 ( .A(A[84]), .B(B[84]), .Z(n1712) );
  NAND U1499 ( .A(n1713), .B(n1714), .Z(n1711) );
  NANDN U1500 ( .A(B[84]), .B(A[84]), .Z(n1714) );
  AND U1501 ( .A(n1715), .B(n1716), .Z(n1713) );
  NAND U1502 ( .A(n1717), .B(n1718), .Z(n1716) );
  NANDN U1503 ( .A(A[83]), .B(B[83]), .Z(n1718) );
  AND U1504 ( .A(n1719), .B(n1720), .Z(n1717) );
  NANDN U1505 ( .A(A[82]), .B(B[82]), .Z(n1720) );
  NAND U1506 ( .A(n1721), .B(n1722), .Z(n1719) );
  NANDN U1507 ( .A(B[82]), .B(A[82]), .Z(n1722) );
  AND U1508 ( .A(n1723), .B(n1724), .Z(n1721) );
  NAND U1509 ( .A(n1725), .B(n1726), .Z(n1724) );
  NANDN U1510 ( .A(A[81]), .B(B[81]), .Z(n1726) );
  AND U1511 ( .A(n1727), .B(n1728), .Z(n1725) );
  NANDN U1512 ( .A(A[80]), .B(B[80]), .Z(n1728) );
  NAND U1513 ( .A(n1729), .B(n1730), .Z(n1727) );
  NANDN U1514 ( .A(B[80]), .B(A[80]), .Z(n1730) );
  AND U1515 ( .A(n1731), .B(n1732), .Z(n1729) );
  NAND U1516 ( .A(n1733), .B(n1734), .Z(n1732) );
  NANDN U1517 ( .A(A[79]), .B(B[79]), .Z(n1734) );
  AND U1518 ( .A(n1735), .B(n1736), .Z(n1733) );
  NANDN U1519 ( .A(A[78]), .B(B[78]), .Z(n1736) );
  NAND U1520 ( .A(n1737), .B(n1738), .Z(n1735) );
  NANDN U1521 ( .A(B[78]), .B(A[78]), .Z(n1738) );
  AND U1522 ( .A(n1739), .B(n1740), .Z(n1737) );
  NAND U1523 ( .A(n1741), .B(n1742), .Z(n1740) );
  NANDN U1524 ( .A(A[77]), .B(B[77]), .Z(n1742) );
  AND U1525 ( .A(n1743), .B(n1744), .Z(n1741) );
  NANDN U1526 ( .A(A[76]), .B(B[76]), .Z(n1744) );
  NAND U1527 ( .A(n1745), .B(n1746), .Z(n1743) );
  NANDN U1528 ( .A(B[76]), .B(A[76]), .Z(n1746) );
  AND U1529 ( .A(n1747), .B(n1748), .Z(n1745) );
  NAND U1530 ( .A(n1749), .B(n1750), .Z(n1748) );
  NANDN U1531 ( .A(A[75]), .B(B[75]), .Z(n1750) );
  AND U1532 ( .A(n1751), .B(n1752), .Z(n1749) );
  NANDN U1533 ( .A(A[74]), .B(B[74]), .Z(n1752) );
  NAND U1534 ( .A(n1753), .B(n1754), .Z(n1751) );
  NANDN U1535 ( .A(B[74]), .B(A[74]), .Z(n1754) );
  AND U1536 ( .A(n1755), .B(n1756), .Z(n1753) );
  NAND U1537 ( .A(n1757), .B(n1758), .Z(n1756) );
  NANDN U1538 ( .A(A[73]), .B(B[73]), .Z(n1758) );
  AND U1539 ( .A(n1759), .B(n1760), .Z(n1757) );
  NANDN U1540 ( .A(A[72]), .B(B[72]), .Z(n1760) );
  NAND U1541 ( .A(n1761), .B(n1762), .Z(n1759) );
  NANDN U1542 ( .A(B[72]), .B(A[72]), .Z(n1762) );
  AND U1543 ( .A(n1763), .B(n1764), .Z(n1761) );
  NAND U1544 ( .A(n1765), .B(n1766), .Z(n1764) );
  NANDN U1545 ( .A(A[71]), .B(B[71]), .Z(n1766) );
  AND U1546 ( .A(n1767), .B(n1768), .Z(n1765) );
  NANDN U1547 ( .A(A[70]), .B(B[70]), .Z(n1768) );
  NAND U1548 ( .A(n1769), .B(n1770), .Z(n1767) );
  NANDN U1549 ( .A(B[70]), .B(A[70]), .Z(n1770) );
  AND U1550 ( .A(n1771), .B(n1772), .Z(n1769) );
  NAND U1551 ( .A(n1773), .B(n1774), .Z(n1772) );
  NANDN U1552 ( .A(A[69]), .B(B[69]), .Z(n1774) );
  AND U1553 ( .A(n1775), .B(n1776), .Z(n1773) );
  NANDN U1554 ( .A(A[68]), .B(B[68]), .Z(n1776) );
  NAND U1555 ( .A(n1777), .B(n1778), .Z(n1775) );
  NANDN U1556 ( .A(B[68]), .B(A[68]), .Z(n1778) );
  AND U1557 ( .A(n1779), .B(n1780), .Z(n1777) );
  NAND U1558 ( .A(n1781), .B(n1782), .Z(n1780) );
  NANDN U1559 ( .A(A[67]), .B(B[67]), .Z(n1782) );
  AND U1560 ( .A(n1783), .B(n1784), .Z(n1781) );
  NANDN U1561 ( .A(A[66]), .B(B[66]), .Z(n1784) );
  NAND U1562 ( .A(n1785), .B(n1786), .Z(n1783) );
  NANDN U1563 ( .A(B[66]), .B(A[66]), .Z(n1786) );
  AND U1564 ( .A(n1787), .B(n1788), .Z(n1785) );
  NAND U1565 ( .A(n1789), .B(n1790), .Z(n1788) );
  NANDN U1566 ( .A(A[65]), .B(B[65]), .Z(n1790) );
  AND U1567 ( .A(n1791), .B(n1792), .Z(n1789) );
  NANDN U1568 ( .A(A[64]), .B(B[64]), .Z(n1792) );
  NAND U1569 ( .A(n1793), .B(n1794), .Z(n1791) );
  NANDN U1570 ( .A(B[64]), .B(A[64]), .Z(n1794) );
  AND U1571 ( .A(n1795), .B(n1796), .Z(n1793) );
  NAND U1572 ( .A(n1797), .B(n1798), .Z(n1796) );
  NANDN U1573 ( .A(A[63]), .B(B[63]), .Z(n1798) );
  AND U1574 ( .A(n1799), .B(n1800), .Z(n1797) );
  NANDN U1575 ( .A(A[62]), .B(B[62]), .Z(n1800) );
  NAND U1576 ( .A(n1801), .B(n1802), .Z(n1799) );
  NANDN U1577 ( .A(B[62]), .B(A[62]), .Z(n1802) );
  AND U1578 ( .A(n1803), .B(n1804), .Z(n1801) );
  NAND U1579 ( .A(n1805), .B(n1806), .Z(n1804) );
  NANDN U1580 ( .A(A[61]), .B(B[61]), .Z(n1806) );
  AND U1581 ( .A(n1807), .B(n1808), .Z(n1805) );
  NANDN U1582 ( .A(A[60]), .B(B[60]), .Z(n1808) );
  NAND U1583 ( .A(n1809), .B(n1810), .Z(n1807) );
  NANDN U1584 ( .A(B[60]), .B(A[60]), .Z(n1810) );
  AND U1585 ( .A(n1811), .B(n1812), .Z(n1809) );
  NAND U1586 ( .A(n1813), .B(n1814), .Z(n1812) );
  NANDN U1587 ( .A(A[59]), .B(B[59]), .Z(n1814) );
  AND U1588 ( .A(n1815), .B(n1816), .Z(n1813) );
  NANDN U1589 ( .A(A[58]), .B(B[58]), .Z(n1816) );
  NAND U1590 ( .A(n1817), .B(n1818), .Z(n1815) );
  NANDN U1591 ( .A(B[58]), .B(A[58]), .Z(n1818) );
  AND U1592 ( .A(n1819), .B(n1820), .Z(n1817) );
  NAND U1593 ( .A(n1821), .B(n1822), .Z(n1820) );
  NANDN U1594 ( .A(A[57]), .B(B[57]), .Z(n1822) );
  AND U1595 ( .A(n1823), .B(n1824), .Z(n1821) );
  NANDN U1596 ( .A(A[56]), .B(B[56]), .Z(n1824) );
  NAND U1597 ( .A(n1825), .B(n1826), .Z(n1823) );
  NANDN U1598 ( .A(B[56]), .B(A[56]), .Z(n1826) );
  AND U1599 ( .A(n1827), .B(n1828), .Z(n1825) );
  NAND U1600 ( .A(n1829), .B(n1830), .Z(n1828) );
  NANDN U1601 ( .A(A[55]), .B(B[55]), .Z(n1830) );
  AND U1602 ( .A(n1831), .B(n1832), .Z(n1829) );
  NANDN U1603 ( .A(A[54]), .B(B[54]), .Z(n1832) );
  NAND U1604 ( .A(n1833), .B(n1834), .Z(n1831) );
  NANDN U1605 ( .A(B[54]), .B(A[54]), .Z(n1834) );
  AND U1606 ( .A(n1835), .B(n1836), .Z(n1833) );
  NAND U1607 ( .A(n1837), .B(n1838), .Z(n1836) );
  NANDN U1608 ( .A(A[53]), .B(B[53]), .Z(n1838) );
  AND U1609 ( .A(n1839), .B(n1840), .Z(n1837) );
  NANDN U1610 ( .A(A[52]), .B(B[52]), .Z(n1840) );
  NAND U1611 ( .A(n1841), .B(n1842), .Z(n1839) );
  NANDN U1612 ( .A(B[52]), .B(A[52]), .Z(n1842) );
  AND U1613 ( .A(n1843), .B(n1844), .Z(n1841) );
  NAND U1614 ( .A(n1845), .B(n1846), .Z(n1844) );
  NANDN U1615 ( .A(A[51]), .B(B[51]), .Z(n1846) );
  AND U1616 ( .A(n1847), .B(n1848), .Z(n1845) );
  NANDN U1617 ( .A(A[50]), .B(B[50]), .Z(n1848) );
  NAND U1618 ( .A(n1849), .B(n1850), .Z(n1847) );
  NANDN U1619 ( .A(B[50]), .B(A[50]), .Z(n1850) );
  AND U1620 ( .A(n1851), .B(n1852), .Z(n1849) );
  NAND U1621 ( .A(n1853), .B(n1854), .Z(n1852) );
  NANDN U1622 ( .A(A[49]), .B(B[49]), .Z(n1854) );
  AND U1623 ( .A(n1855), .B(n1856), .Z(n1853) );
  NANDN U1624 ( .A(A[48]), .B(B[48]), .Z(n1856) );
  NAND U1625 ( .A(n1857), .B(n1858), .Z(n1855) );
  NANDN U1626 ( .A(B[48]), .B(A[48]), .Z(n1858) );
  AND U1627 ( .A(n1859), .B(n1860), .Z(n1857) );
  NAND U1628 ( .A(n1861), .B(n1862), .Z(n1860) );
  NANDN U1629 ( .A(A[47]), .B(B[47]), .Z(n1862) );
  AND U1630 ( .A(n1863), .B(n1864), .Z(n1861) );
  NANDN U1631 ( .A(A[46]), .B(B[46]), .Z(n1864) );
  NAND U1632 ( .A(n1865), .B(n1866), .Z(n1863) );
  NANDN U1633 ( .A(B[46]), .B(A[46]), .Z(n1866) );
  AND U1634 ( .A(n1867), .B(n1868), .Z(n1865) );
  NAND U1635 ( .A(n1869), .B(n1870), .Z(n1868) );
  NANDN U1636 ( .A(A[45]), .B(B[45]), .Z(n1870) );
  AND U1637 ( .A(n1871), .B(n1872), .Z(n1869) );
  NANDN U1638 ( .A(A[44]), .B(B[44]), .Z(n1872) );
  NAND U1639 ( .A(n1873), .B(n1874), .Z(n1871) );
  NANDN U1640 ( .A(B[44]), .B(A[44]), .Z(n1874) );
  AND U1641 ( .A(n1875), .B(n1876), .Z(n1873) );
  NAND U1642 ( .A(n1877), .B(n1878), .Z(n1876) );
  NANDN U1643 ( .A(A[43]), .B(B[43]), .Z(n1878) );
  AND U1644 ( .A(n1879), .B(n1880), .Z(n1877) );
  NANDN U1645 ( .A(A[42]), .B(B[42]), .Z(n1880) );
  NAND U1646 ( .A(n1881), .B(n1882), .Z(n1879) );
  NANDN U1647 ( .A(B[42]), .B(A[42]), .Z(n1882) );
  AND U1648 ( .A(n1883), .B(n1884), .Z(n1881) );
  NAND U1649 ( .A(n1885), .B(n1886), .Z(n1884) );
  NANDN U1650 ( .A(A[41]), .B(B[41]), .Z(n1886) );
  AND U1651 ( .A(n1887), .B(n1888), .Z(n1885) );
  NANDN U1652 ( .A(A[40]), .B(B[40]), .Z(n1888) );
  NAND U1653 ( .A(n1889), .B(n1890), .Z(n1887) );
  NANDN U1654 ( .A(B[40]), .B(A[40]), .Z(n1890) );
  AND U1655 ( .A(n1891), .B(n1892), .Z(n1889) );
  NAND U1656 ( .A(n1893), .B(n1894), .Z(n1892) );
  NANDN U1657 ( .A(A[39]), .B(B[39]), .Z(n1894) );
  AND U1658 ( .A(n1895), .B(n1896), .Z(n1893) );
  NANDN U1659 ( .A(A[38]), .B(B[38]), .Z(n1896) );
  NAND U1660 ( .A(n1897), .B(n1898), .Z(n1895) );
  NANDN U1661 ( .A(B[38]), .B(A[38]), .Z(n1898) );
  AND U1662 ( .A(n1899), .B(n1900), .Z(n1897) );
  NAND U1663 ( .A(n1901), .B(n1902), .Z(n1900) );
  NANDN U1664 ( .A(A[37]), .B(B[37]), .Z(n1902) );
  AND U1665 ( .A(n1903), .B(n1904), .Z(n1901) );
  NANDN U1666 ( .A(A[36]), .B(B[36]), .Z(n1904) );
  NAND U1667 ( .A(n1905), .B(n1906), .Z(n1903) );
  NANDN U1668 ( .A(B[36]), .B(A[36]), .Z(n1906) );
  AND U1669 ( .A(n1907), .B(n1908), .Z(n1905) );
  NAND U1670 ( .A(n1909), .B(n1910), .Z(n1908) );
  NANDN U1671 ( .A(A[35]), .B(B[35]), .Z(n1910) );
  AND U1672 ( .A(n1911), .B(n1912), .Z(n1909) );
  NANDN U1673 ( .A(A[34]), .B(B[34]), .Z(n1912) );
  NAND U1674 ( .A(n1913), .B(n1914), .Z(n1911) );
  NANDN U1675 ( .A(B[34]), .B(A[34]), .Z(n1914) );
  AND U1676 ( .A(n1915), .B(n1916), .Z(n1913) );
  NAND U1677 ( .A(n1917), .B(n1918), .Z(n1916) );
  NANDN U1678 ( .A(A[33]), .B(B[33]), .Z(n1918) );
  AND U1679 ( .A(n1919), .B(n1920), .Z(n1917) );
  NANDN U1680 ( .A(A[32]), .B(B[32]), .Z(n1920) );
  NAND U1681 ( .A(n1921), .B(n1922), .Z(n1919) );
  NANDN U1682 ( .A(B[32]), .B(A[32]), .Z(n1922) );
  AND U1683 ( .A(n1923), .B(n1924), .Z(n1921) );
  NAND U1684 ( .A(n1925), .B(n1926), .Z(n1924) );
  NANDN U1685 ( .A(A[31]), .B(B[31]), .Z(n1926) );
  AND U1686 ( .A(n1927), .B(n1928), .Z(n1925) );
  NANDN U1687 ( .A(A[30]), .B(B[30]), .Z(n1928) );
  NAND U1688 ( .A(n1929), .B(n1930), .Z(n1927) );
  NANDN U1689 ( .A(B[30]), .B(A[30]), .Z(n1930) );
  AND U1690 ( .A(n1931), .B(n1932), .Z(n1929) );
  NAND U1691 ( .A(n1933), .B(n1934), .Z(n1932) );
  NANDN U1692 ( .A(A[29]), .B(B[29]), .Z(n1934) );
  AND U1693 ( .A(n1935), .B(n1936), .Z(n1933) );
  NANDN U1694 ( .A(A[28]), .B(B[28]), .Z(n1936) );
  NAND U1695 ( .A(n1937), .B(n1938), .Z(n1935) );
  NANDN U1696 ( .A(B[28]), .B(A[28]), .Z(n1938) );
  AND U1697 ( .A(n1939), .B(n1940), .Z(n1937) );
  NAND U1698 ( .A(n1941), .B(n1942), .Z(n1940) );
  NANDN U1699 ( .A(A[27]), .B(B[27]), .Z(n1942) );
  AND U1700 ( .A(n1943), .B(n1944), .Z(n1941) );
  NANDN U1701 ( .A(A[26]), .B(B[26]), .Z(n1944) );
  NAND U1702 ( .A(n1945), .B(n1946), .Z(n1943) );
  NANDN U1703 ( .A(B[26]), .B(A[26]), .Z(n1946) );
  AND U1704 ( .A(n1947), .B(n1948), .Z(n1945) );
  NAND U1705 ( .A(n1949), .B(n1950), .Z(n1948) );
  NANDN U1706 ( .A(A[25]), .B(B[25]), .Z(n1950) );
  AND U1707 ( .A(n1951), .B(n1952), .Z(n1949) );
  NANDN U1708 ( .A(A[24]), .B(B[24]), .Z(n1952) );
  NAND U1709 ( .A(n1953), .B(n1954), .Z(n1951) );
  NANDN U1710 ( .A(B[24]), .B(A[24]), .Z(n1954) );
  AND U1711 ( .A(n1955), .B(n1956), .Z(n1953) );
  NAND U1712 ( .A(n1957), .B(n1958), .Z(n1956) );
  NANDN U1713 ( .A(A[23]), .B(B[23]), .Z(n1958) );
  AND U1714 ( .A(n1959), .B(n1960), .Z(n1957) );
  NANDN U1715 ( .A(A[22]), .B(B[22]), .Z(n1960) );
  NAND U1716 ( .A(n1961), .B(n1962), .Z(n1959) );
  NANDN U1717 ( .A(B[22]), .B(A[22]), .Z(n1962) );
  AND U1718 ( .A(n1963), .B(n1964), .Z(n1961) );
  NAND U1719 ( .A(n1965), .B(n1966), .Z(n1964) );
  NANDN U1720 ( .A(A[21]), .B(B[21]), .Z(n1966) );
  AND U1721 ( .A(n1967), .B(n1968), .Z(n1965) );
  NANDN U1722 ( .A(A[20]), .B(B[20]), .Z(n1968) );
  NAND U1723 ( .A(n1969), .B(n1970), .Z(n1967) );
  NANDN U1724 ( .A(B[20]), .B(A[20]), .Z(n1970) );
  AND U1725 ( .A(n1971), .B(n1972), .Z(n1969) );
  NAND U1726 ( .A(n1973), .B(n1974), .Z(n1972) );
  NANDN U1727 ( .A(A[19]), .B(B[19]), .Z(n1974) );
  AND U1728 ( .A(n1975), .B(n1976), .Z(n1973) );
  NANDN U1729 ( .A(A[18]), .B(B[18]), .Z(n1976) );
  NAND U1730 ( .A(n1977), .B(n1978), .Z(n1975) );
  NANDN U1731 ( .A(B[18]), .B(A[18]), .Z(n1978) );
  AND U1732 ( .A(n1979), .B(n1980), .Z(n1977) );
  NAND U1733 ( .A(n1981), .B(n1982), .Z(n1980) );
  NANDN U1734 ( .A(A[17]), .B(B[17]), .Z(n1982) );
  AND U1735 ( .A(n1983), .B(n1984), .Z(n1981) );
  NANDN U1736 ( .A(A[16]), .B(B[16]), .Z(n1984) );
  NAND U1737 ( .A(n1985), .B(n1986), .Z(n1983) );
  NANDN U1738 ( .A(B[16]), .B(A[16]), .Z(n1986) );
  AND U1739 ( .A(n1987), .B(n1988), .Z(n1985) );
  NAND U1740 ( .A(n1989), .B(n1990), .Z(n1988) );
  NANDN U1741 ( .A(A[15]), .B(B[15]), .Z(n1990) );
  AND U1742 ( .A(n1991), .B(n1992), .Z(n1989) );
  NANDN U1743 ( .A(A[14]), .B(B[14]), .Z(n1992) );
  NAND U1744 ( .A(n1993), .B(n1994), .Z(n1991) );
  NANDN U1745 ( .A(B[14]), .B(A[14]), .Z(n1994) );
  AND U1746 ( .A(n1995), .B(n1996), .Z(n1993) );
  NAND U1747 ( .A(n1997), .B(n1998), .Z(n1996) );
  NANDN U1748 ( .A(A[13]), .B(B[13]), .Z(n1998) );
  AND U1749 ( .A(n1999), .B(n2000), .Z(n1997) );
  NANDN U1750 ( .A(A[12]), .B(B[12]), .Z(n2000) );
  NAND U1751 ( .A(n2001), .B(n2002), .Z(n1999) );
  NANDN U1752 ( .A(B[12]), .B(A[12]), .Z(n2002) );
  AND U1753 ( .A(n2003), .B(n2004), .Z(n2001) );
  NAND U1754 ( .A(n2005), .B(n2006), .Z(n2004) );
  NANDN U1755 ( .A(A[11]), .B(B[11]), .Z(n2006) );
  AND U1756 ( .A(n2007), .B(n2008), .Z(n2005) );
  NANDN U1757 ( .A(A[10]), .B(B[10]), .Z(n2008) );
  NAND U1758 ( .A(n2009), .B(n2010), .Z(n2007) );
  NANDN U1759 ( .A(B[9]), .B(A[9]), .Z(n2010) );
  AND U1760 ( .A(n2011), .B(n2012), .Z(n2009) );
  NAND U1761 ( .A(n2013), .B(n2014), .Z(n2012) );
  NANDN U1762 ( .A(A[9]), .B(B[9]), .Z(n2014) );
  AND U1763 ( .A(n2015), .B(n2016), .Z(n2013) );
  NANDN U1764 ( .A(A[8]), .B(B[8]), .Z(n2016) );
  NAND U1765 ( .A(n2017), .B(n2018), .Z(n2015) );
  NANDN U1766 ( .A(B[8]), .B(A[8]), .Z(n2018) );
  AND U1767 ( .A(n2019), .B(n2020), .Z(n2017) );
  NAND U1768 ( .A(n2021), .B(n2022), .Z(n2020) );
  NANDN U1769 ( .A(A[7]), .B(B[7]), .Z(n2022) );
  AND U1770 ( .A(n2023), .B(n2024), .Z(n2021) );
  NANDN U1771 ( .A(A[6]), .B(B[6]), .Z(n2024) );
  NAND U1772 ( .A(n2025), .B(n2026), .Z(n2023) );
  NANDN U1773 ( .A(B[6]), .B(A[6]), .Z(n2026) );
  AND U1774 ( .A(n2027), .B(n2028), .Z(n2025) );
  NAND U1775 ( .A(n2029), .B(n2030), .Z(n2028) );
  NANDN U1776 ( .A(A[5]), .B(B[5]), .Z(n2030) );
  AND U1777 ( .A(n2031), .B(n2032), .Z(n2029) );
  NANDN U1778 ( .A(A[4]), .B(B[4]), .Z(n2032) );
  NAND U1779 ( .A(n2033), .B(n2034), .Z(n2031) );
  NANDN U1780 ( .A(B[4]), .B(A[4]), .Z(n2034) );
  AND U1781 ( .A(n2035), .B(n2036), .Z(n2033) );
  NAND U1782 ( .A(n2037), .B(n2038), .Z(n2036) );
  NANDN U1783 ( .A(A[3]), .B(B[3]), .Z(n2038) );
  AND U1784 ( .A(n2039), .B(n2040), .Z(n2037) );
  NANDN U1785 ( .A(A[2]), .B(B[2]), .Z(n2040) );
  NAND U1786 ( .A(n2041), .B(n2042), .Z(n2039) );
  NANDN U1787 ( .A(B[2]), .B(A[2]), .Z(n2042) );
  AND U1788 ( .A(n2043), .B(n2044), .Z(n2041) );
  NANDN U1789 ( .A(B[1]), .B(n2045), .Z(n2044) );
  NANDN U1790 ( .A(A[1]), .B(n2046), .Z(n2045) );
  NANDN U1791 ( .A(n2046), .B(A[1]), .Z(n2043) );
  ANDN U1792 ( .B(B[0]), .A(A[0]), .Z(n2046) );
  NANDN U1793 ( .A(B[3]), .B(A[3]), .Z(n2035) );
  NANDN U1794 ( .A(B[5]), .B(A[5]), .Z(n2027) );
  NANDN U1795 ( .A(B[7]), .B(A[7]), .Z(n2019) );
  NANDN U1796 ( .A(B[10]), .B(A[10]), .Z(n2011) );
  NANDN U1797 ( .A(B[11]), .B(A[11]), .Z(n2003) );
  NANDN U1798 ( .A(B[13]), .B(A[13]), .Z(n1995) );
  NANDN U1799 ( .A(B[15]), .B(A[15]), .Z(n1987) );
  NANDN U1800 ( .A(B[17]), .B(A[17]), .Z(n1979) );
  NANDN U1801 ( .A(B[19]), .B(A[19]), .Z(n1971) );
  NANDN U1802 ( .A(B[21]), .B(A[21]), .Z(n1963) );
  NANDN U1803 ( .A(B[23]), .B(A[23]), .Z(n1955) );
  NANDN U1804 ( .A(B[25]), .B(A[25]), .Z(n1947) );
  NANDN U1805 ( .A(B[27]), .B(A[27]), .Z(n1939) );
  NANDN U1806 ( .A(B[29]), .B(A[29]), .Z(n1931) );
  NANDN U1807 ( .A(B[31]), .B(A[31]), .Z(n1923) );
  NANDN U1808 ( .A(B[33]), .B(A[33]), .Z(n1915) );
  NANDN U1809 ( .A(B[35]), .B(A[35]), .Z(n1907) );
  NANDN U1810 ( .A(B[37]), .B(A[37]), .Z(n1899) );
  NANDN U1811 ( .A(B[39]), .B(A[39]), .Z(n1891) );
  NANDN U1812 ( .A(B[41]), .B(A[41]), .Z(n1883) );
  NANDN U1813 ( .A(B[43]), .B(A[43]), .Z(n1875) );
  NANDN U1814 ( .A(B[45]), .B(A[45]), .Z(n1867) );
  NANDN U1815 ( .A(B[47]), .B(A[47]), .Z(n1859) );
  NANDN U1816 ( .A(B[49]), .B(A[49]), .Z(n1851) );
  NANDN U1817 ( .A(B[51]), .B(A[51]), .Z(n1843) );
  NANDN U1818 ( .A(B[53]), .B(A[53]), .Z(n1835) );
  NANDN U1819 ( .A(B[55]), .B(A[55]), .Z(n1827) );
  NANDN U1820 ( .A(B[57]), .B(A[57]), .Z(n1819) );
  NANDN U1821 ( .A(B[59]), .B(A[59]), .Z(n1811) );
  NANDN U1822 ( .A(B[61]), .B(A[61]), .Z(n1803) );
  NANDN U1823 ( .A(B[63]), .B(A[63]), .Z(n1795) );
  NANDN U1824 ( .A(B[65]), .B(A[65]), .Z(n1787) );
  NANDN U1825 ( .A(B[67]), .B(A[67]), .Z(n1779) );
  NANDN U1826 ( .A(B[69]), .B(A[69]), .Z(n1771) );
  NANDN U1827 ( .A(B[71]), .B(A[71]), .Z(n1763) );
  NANDN U1828 ( .A(B[73]), .B(A[73]), .Z(n1755) );
  NANDN U1829 ( .A(B[75]), .B(A[75]), .Z(n1747) );
  NANDN U1830 ( .A(B[77]), .B(A[77]), .Z(n1739) );
  NANDN U1831 ( .A(B[79]), .B(A[79]), .Z(n1731) );
  NANDN U1832 ( .A(B[81]), .B(A[81]), .Z(n1723) );
  NANDN U1833 ( .A(B[83]), .B(A[83]), .Z(n1715) );
  NANDN U1834 ( .A(B[85]), .B(A[85]), .Z(n1707) );
  NANDN U1835 ( .A(B[87]), .B(A[87]), .Z(n1699) );
  NANDN U1836 ( .A(B[89]), .B(A[89]), .Z(n1691) );
  NANDN U1837 ( .A(B[91]), .B(A[91]), .Z(n1683) );
  NANDN U1838 ( .A(B[93]), .B(A[93]), .Z(n1675) );
  NANDN U1839 ( .A(B[95]), .B(A[95]), .Z(n1667) );
  NANDN U1840 ( .A(B[97]), .B(A[97]), .Z(n1659) );
  NANDN U1841 ( .A(B[100]), .B(A[100]), .Z(n1651) );
  NANDN U1842 ( .A(B[101]), .B(A[101]), .Z(n1643) );
  NANDN U1843 ( .A(B[103]), .B(A[103]), .Z(n1635) );
  NANDN U1844 ( .A(B[105]), .B(A[105]), .Z(n1627) );
  NANDN U1845 ( .A(B[107]), .B(A[107]), .Z(n1619) );
  NANDN U1846 ( .A(B[109]), .B(A[109]), .Z(n1611) );
  NANDN U1847 ( .A(B[111]), .B(A[111]), .Z(n1603) );
  NANDN U1848 ( .A(B[113]), .B(A[113]), .Z(n1595) );
  NANDN U1849 ( .A(B[115]), .B(A[115]), .Z(n1587) );
  NANDN U1850 ( .A(B[117]), .B(A[117]), .Z(n1579) );
  NANDN U1851 ( .A(B[119]), .B(A[119]), .Z(n1571) );
  NANDN U1852 ( .A(B[121]), .B(A[121]), .Z(n1563) );
  NANDN U1853 ( .A(B[123]), .B(A[123]), .Z(n1555) );
  NANDN U1854 ( .A(B[125]), .B(A[125]), .Z(n1547) );
  NANDN U1855 ( .A(B[127]), .B(A[127]), .Z(n1539) );
  NANDN U1856 ( .A(B[129]), .B(A[129]), .Z(n1531) );
  NANDN U1857 ( .A(B[131]), .B(A[131]), .Z(n1523) );
  NANDN U1858 ( .A(B[133]), .B(A[133]), .Z(n1515) );
  NANDN U1859 ( .A(B[135]), .B(A[135]), .Z(n1507) );
  NANDN U1860 ( .A(B[137]), .B(A[137]), .Z(n1499) );
  NANDN U1861 ( .A(B[139]), .B(A[139]), .Z(n1491) );
  NANDN U1862 ( .A(B[141]), .B(A[141]), .Z(n1483) );
  NANDN U1863 ( .A(B[143]), .B(A[143]), .Z(n1475) );
  NANDN U1864 ( .A(B[145]), .B(A[145]), .Z(n1467) );
  NANDN U1865 ( .A(B[147]), .B(A[147]), .Z(n1459) );
  NANDN U1866 ( .A(B[149]), .B(A[149]), .Z(n1451) );
  NANDN U1867 ( .A(B[151]), .B(A[151]), .Z(n1443) );
  NANDN U1868 ( .A(B[153]), .B(A[153]), .Z(n1435) );
  NANDN U1869 ( .A(B[155]), .B(A[155]), .Z(n1427) );
  NANDN U1870 ( .A(B[157]), .B(A[157]), .Z(n1419) );
  NANDN U1871 ( .A(B[159]), .B(A[159]), .Z(n1411) );
  NANDN U1872 ( .A(B[161]), .B(A[161]), .Z(n1403) );
  NANDN U1873 ( .A(B[163]), .B(A[163]), .Z(n1395) );
  NANDN U1874 ( .A(B[165]), .B(A[165]), .Z(n1387) );
  NANDN U1875 ( .A(B[167]), .B(A[167]), .Z(n1379) );
  NANDN U1876 ( .A(B[169]), .B(A[169]), .Z(n1371) );
  NANDN U1877 ( .A(B[171]), .B(A[171]), .Z(n1363) );
  NANDN U1878 ( .A(B[173]), .B(A[173]), .Z(n1355) );
  NANDN U1879 ( .A(B[175]), .B(A[175]), .Z(n1347) );
  NANDN U1880 ( .A(B[177]), .B(A[177]), .Z(n1339) );
  NANDN U1881 ( .A(B[179]), .B(A[179]), .Z(n1331) );
  NANDN U1882 ( .A(B[181]), .B(A[181]), .Z(n1323) );
  NANDN U1883 ( .A(B[183]), .B(A[183]), .Z(n1315) );
  NANDN U1884 ( .A(B[185]), .B(A[185]), .Z(n1307) );
  NANDN U1885 ( .A(B[187]), .B(A[187]), .Z(n1299) );
  NANDN U1886 ( .A(B[189]), .B(A[189]), .Z(n1291) );
  NANDN U1887 ( .A(B[191]), .B(A[191]), .Z(n1283) );
  NANDN U1888 ( .A(B[193]), .B(A[193]), .Z(n1275) );
  NANDN U1889 ( .A(B[195]), .B(A[195]), .Z(n1267) );
  NANDN U1890 ( .A(B[197]), .B(A[197]), .Z(n1259) );
  NANDN U1891 ( .A(B[199]), .B(A[199]), .Z(n1251) );
  NANDN U1892 ( .A(B[201]), .B(A[201]), .Z(n1243) );
  NANDN U1893 ( .A(B[203]), .B(A[203]), .Z(n1235) );
  NANDN U1894 ( .A(B[205]), .B(A[205]), .Z(n1227) );
  NANDN U1895 ( .A(B[207]), .B(A[207]), .Z(n1219) );
  NANDN U1896 ( .A(B[209]), .B(A[209]), .Z(n1211) );
  NANDN U1897 ( .A(B[211]), .B(A[211]), .Z(n1203) );
  NANDN U1898 ( .A(B[213]), .B(A[213]), .Z(n1195) );
  NANDN U1899 ( .A(B[215]), .B(A[215]), .Z(n1187) );
  NANDN U1900 ( .A(B[217]), .B(A[217]), .Z(n1179) );
  NANDN U1901 ( .A(B[219]), .B(A[219]), .Z(n1171) );
  NANDN U1902 ( .A(B[221]), .B(A[221]), .Z(n1163) );
  NANDN U1903 ( .A(B[223]), .B(A[223]), .Z(n1155) );
  NANDN U1904 ( .A(B[225]), .B(A[225]), .Z(n1147) );
  NANDN U1905 ( .A(B[227]), .B(A[227]), .Z(n1139) );
  NANDN U1906 ( .A(B[229]), .B(A[229]), .Z(n1131) );
  NANDN U1907 ( .A(B[231]), .B(A[231]), .Z(n1123) );
  NANDN U1908 ( .A(B[233]), .B(A[233]), .Z(n1115) );
  NANDN U1909 ( .A(B[235]), .B(A[235]), .Z(n1107) );
  NANDN U1910 ( .A(B[237]), .B(A[237]), .Z(n1099) );
  NANDN U1911 ( .A(B[239]), .B(A[239]), .Z(n1091) );
  NANDN U1912 ( .A(B[241]), .B(A[241]), .Z(n1083) );
  NANDN U1913 ( .A(B[243]), .B(A[243]), .Z(n1075) );
  NANDN U1914 ( .A(B[245]), .B(A[245]), .Z(n1067) );
  NANDN U1915 ( .A(B[247]), .B(A[247]), .Z(n1059) );
  NANDN U1916 ( .A(B[249]), .B(A[249]), .Z(n1051) );
  NANDN U1917 ( .A(B[251]), .B(A[251]), .Z(n1043) );
  NANDN U1918 ( .A(B[253]), .B(A[253]), .Z(n1035) );
  NANDN U1919 ( .A(B[255]), .B(A[255]), .Z(n1027) );
  NANDN U1920 ( .A(B[257]), .B(A[257]), .Z(n1019) );
  NANDN U1921 ( .A(B[259]), .B(A[259]), .Z(n1011) );
  NANDN U1922 ( .A(B[261]), .B(A[261]), .Z(n1003) );
  NANDN U1923 ( .A(B[263]), .B(A[263]), .Z(n995) );
  NANDN U1924 ( .A(B[265]), .B(A[265]), .Z(n987) );
  NANDN U1925 ( .A(B[267]), .B(A[267]), .Z(n979) );
  NANDN U1926 ( .A(B[269]), .B(A[269]), .Z(n971) );
  NANDN U1927 ( .A(B[271]), .B(A[271]), .Z(n963) );
  NANDN U1928 ( .A(B[273]), .B(A[273]), .Z(n955) );
  NANDN U1929 ( .A(B[275]), .B(A[275]), .Z(n947) );
  NANDN U1930 ( .A(B[277]), .B(A[277]), .Z(n939) );
  NANDN U1931 ( .A(B[279]), .B(A[279]), .Z(n931) );
  NANDN U1932 ( .A(B[281]), .B(A[281]), .Z(n923) );
  NANDN U1933 ( .A(B[283]), .B(A[283]), .Z(n915) );
  NANDN U1934 ( .A(B[285]), .B(A[285]), .Z(n907) );
  NANDN U1935 ( .A(B[287]), .B(A[287]), .Z(n899) );
  NANDN U1936 ( .A(B[289]), .B(A[289]), .Z(n891) );
  NANDN U1937 ( .A(B[291]), .B(A[291]), .Z(n883) );
  NANDN U1938 ( .A(B[293]), .B(A[293]), .Z(n875) );
  NANDN U1939 ( .A(B[295]), .B(A[295]), .Z(n867) );
  NANDN U1940 ( .A(B[297]), .B(A[297]), .Z(n859) );
  NANDN U1941 ( .A(B[299]), .B(A[299]), .Z(n851) );
  NANDN U1942 ( .A(B[301]), .B(A[301]), .Z(n843) );
  NANDN U1943 ( .A(B[303]), .B(A[303]), .Z(n835) );
  NANDN U1944 ( .A(B[305]), .B(A[305]), .Z(n827) );
  NANDN U1945 ( .A(B[307]), .B(A[307]), .Z(n819) );
  NANDN U1946 ( .A(B[309]), .B(A[309]), .Z(n811) );
  NANDN U1947 ( .A(B[311]), .B(A[311]), .Z(n803) );
  NANDN U1948 ( .A(B[313]), .B(A[313]), .Z(n795) );
  NANDN U1949 ( .A(B[315]), .B(A[315]), .Z(n787) );
  NANDN U1950 ( .A(B[317]), .B(A[317]), .Z(n779) );
  NANDN U1951 ( .A(B[319]), .B(A[319]), .Z(n771) );
  NANDN U1952 ( .A(B[321]), .B(A[321]), .Z(n763) );
  NANDN U1953 ( .A(B[323]), .B(A[323]), .Z(n755) );
  NANDN U1954 ( .A(B[325]), .B(A[325]), .Z(n747) );
  NANDN U1955 ( .A(B[327]), .B(A[327]), .Z(n739) );
  NANDN U1956 ( .A(B[329]), .B(A[329]), .Z(n731) );
  NANDN U1957 ( .A(B[331]), .B(A[331]), .Z(n723) );
  NANDN U1958 ( .A(B[333]), .B(A[333]), .Z(n715) );
  NANDN U1959 ( .A(B[335]), .B(A[335]), .Z(n707) );
  NANDN U1960 ( .A(B[337]), .B(A[337]), .Z(n699) );
  NANDN U1961 ( .A(B[339]), .B(A[339]), .Z(n691) );
  NANDN U1962 ( .A(B[341]), .B(A[341]), .Z(n683) );
  NANDN U1963 ( .A(B[343]), .B(A[343]), .Z(n675) );
  NANDN U1964 ( .A(B[345]), .B(A[345]), .Z(n667) );
  NANDN U1965 ( .A(B[347]), .B(A[347]), .Z(n659) );
  NANDN U1966 ( .A(B[349]), .B(A[349]), .Z(n651) );
  NANDN U1967 ( .A(B[351]), .B(A[351]), .Z(n643) );
  NANDN U1968 ( .A(B[353]), .B(A[353]), .Z(n635) );
  NANDN U1969 ( .A(B[355]), .B(A[355]), .Z(n627) );
  NANDN U1970 ( .A(B[357]), .B(A[357]), .Z(n619) );
  NANDN U1971 ( .A(B[359]), .B(A[359]), .Z(n611) );
  NANDN U1972 ( .A(B[361]), .B(A[361]), .Z(n603) );
  NANDN U1973 ( .A(B[363]), .B(A[363]), .Z(n595) );
  NANDN U1974 ( .A(B[365]), .B(A[365]), .Z(n587) );
  NANDN U1975 ( .A(B[367]), .B(A[367]), .Z(n579) );
  NANDN U1976 ( .A(B[369]), .B(A[369]), .Z(n571) );
  NANDN U1977 ( .A(B[371]), .B(A[371]), .Z(n563) );
  NANDN U1978 ( .A(B[373]), .B(A[373]), .Z(n555) );
  NANDN U1979 ( .A(B[375]), .B(A[375]), .Z(n547) );
  NANDN U1980 ( .A(B[377]), .B(A[377]), .Z(n539) );
  NANDN U1981 ( .A(B[379]), .B(A[379]), .Z(n531) );
  NANDN U1982 ( .A(B[381]), .B(A[381]), .Z(n523) );
  NANDN U1983 ( .A(B[383]), .B(A[383]), .Z(n515) );
  NANDN U1984 ( .A(B[385]), .B(A[385]), .Z(n507) );
  NANDN U1985 ( .A(B[387]), .B(A[387]), .Z(n499) );
  NANDN U1986 ( .A(B[389]), .B(A[389]), .Z(n491) );
  NANDN U1987 ( .A(B[391]), .B(A[391]), .Z(n483) );
  NANDN U1988 ( .A(B[393]), .B(A[393]), .Z(n475) );
  NANDN U1989 ( .A(B[395]), .B(A[395]), .Z(n467) );
  NANDN U1990 ( .A(B[397]), .B(A[397]), .Z(n459) );
  NANDN U1991 ( .A(B[399]), .B(A[399]), .Z(n451) );
  NANDN U1992 ( .A(B[401]), .B(A[401]), .Z(n443) );
  NANDN U1993 ( .A(B[403]), .B(A[403]), .Z(n435) );
  NANDN U1994 ( .A(B[405]), .B(A[405]), .Z(n427) );
  NANDN U1995 ( .A(B[407]), .B(A[407]), .Z(n419) );
  NANDN U1996 ( .A(B[409]), .B(A[409]), .Z(n411) );
  NANDN U1997 ( .A(B[411]), .B(A[411]), .Z(n403) );
  NANDN U1998 ( .A(B[413]), .B(A[413]), .Z(n395) );
  NANDN U1999 ( .A(B[415]), .B(A[415]), .Z(n387) );
  NANDN U2000 ( .A(B[417]), .B(A[417]), .Z(n379) );
  NANDN U2001 ( .A(B[419]), .B(A[419]), .Z(n371) );
  NANDN U2002 ( .A(B[421]), .B(A[421]), .Z(n363) );
  NANDN U2003 ( .A(B[423]), .B(A[423]), .Z(n355) );
  NANDN U2004 ( .A(B[425]), .B(A[425]), .Z(n347) );
  NANDN U2005 ( .A(B[427]), .B(A[427]), .Z(n339) );
  NANDN U2006 ( .A(B[429]), .B(A[429]), .Z(n331) );
  NANDN U2007 ( .A(B[431]), .B(A[431]), .Z(n323) );
  NANDN U2008 ( .A(B[433]), .B(A[433]), .Z(n315) );
  NANDN U2009 ( .A(B[435]), .B(A[435]), .Z(n307) );
  NANDN U2010 ( .A(B[437]), .B(A[437]), .Z(n299) );
  NANDN U2011 ( .A(B[439]), .B(A[439]), .Z(n291) );
  NANDN U2012 ( .A(B[441]), .B(A[441]), .Z(n283) );
  NANDN U2013 ( .A(B[443]), .B(A[443]), .Z(n275) );
  NANDN U2014 ( .A(B[445]), .B(A[445]), .Z(n267) );
  NANDN U2015 ( .A(B[447]), .B(A[447]), .Z(n259) );
  NANDN U2016 ( .A(B[449]), .B(A[449]), .Z(n251) );
  NANDN U2017 ( .A(B[451]), .B(A[451]), .Z(n243) );
  NANDN U2018 ( .A(B[453]), .B(A[453]), .Z(n235) );
  NANDN U2019 ( .A(B[455]), .B(A[455]), .Z(n227) );
  NANDN U2020 ( .A(B[457]), .B(A[457]), .Z(n219) );
  NANDN U2021 ( .A(B[459]), .B(A[459]), .Z(n211) );
  NANDN U2022 ( .A(B[461]), .B(A[461]), .Z(n203) );
  NANDN U2023 ( .A(B[463]), .B(A[463]), .Z(n195) );
  NANDN U2024 ( .A(B[465]), .B(A[465]), .Z(n187) );
  NANDN U2025 ( .A(B[467]), .B(A[467]), .Z(n179) );
  NANDN U2026 ( .A(B[469]), .B(A[469]), .Z(n171) );
  NANDN U2027 ( .A(B[471]), .B(A[471]), .Z(n163) );
  NANDN U2028 ( .A(B[473]), .B(A[473]), .Z(n155) );
  NANDN U2029 ( .A(B[475]), .B(A[475]), .Z(n147) );
  NANDN U2030 ( .A(B[477]), .B(A[477]), .Z(n139) );
  NANDN U2031 ( .A(B[479]), .B(A[479]), .Z(n131) );
  NANDN U2032 ( .A(B[481]), .B(A[481]), .Z(n123) );
  NANDN U2033 ( .A(B[483]), .B(A[483]), .Z(n115) );
  NANDN U2034 ( .A(B[485]), .B(A[485]), .Z(n107) );
  NANDN U2035 ( .A(B[487]), .B(A[487]), .Z(n99) );
  NANDN U2036 ( .A(B[489]), .B(A[489]), .Z(n91) );
  NANDN U2037 ( .A(B[491]), .B(A[491]), .Z(n83) );
  NANDN U2038 ( .A(B[493]), .B(A[493]), .Z(n75) );
  NANDN U2039 ( .A(B[495]), .B(A[495]), .Z(n67) );
  NANDN U2040 ( .A(B[497]), .B(A[497]), .Z(n59) );
  NANDN U2041 ( .A(B[499]), .B(A[499]), .Z(n51) );
  NANDN U2042 ( .A(B[501]), .B(A[501]), .Z(n43) );
  NANDN U2043 ( .A(B[503]), .B(A[503]), .Z(n35) );
  NANDN U2044 ( .A(B[505]), .B(A[505]), .Z(n27) );
  NANDN U2045 ( .A(B[507]), .B(A[507]), .Z(n19) );
  NANDN U2046 ( .A(B[509]), .B(A[509]), .Z(n11) );
  NANDN U2047 ( .A(A[511]), .B(B[511]), .Z(n3) );
endmodule


module modmult_step_N512_DW01_add_0 ( A, B, CI, SUM, CO );
  input [513:0] A;
  input [513:0] B;
  output [513:0] SUM;
  input CI;
  output CO;
  wire   \B[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
         n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
         n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
         n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
         n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
         n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
         n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
         n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
         n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
         n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
         n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
         n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
         n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
         n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
         n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
         n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
         n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
         n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
         n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
         n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
         n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
         n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
         n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711,
         n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
         n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
         n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
         n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
         n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
         n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
         n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
         n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791,
         n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
         n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
         n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
         n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831,
         n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
         n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
         n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
         n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
         n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
         n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
         n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
         n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
         n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
         n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931,
         n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
         n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
         n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
         n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971,
         n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981,
         n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
         n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
         n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011,
         n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021,
         n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
         n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
         n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
         n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
         n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
         n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
         n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
         n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
         n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
         n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
         n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
         n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
         n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
         n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
         n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
         n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
         n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
         n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
         n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
         n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
         n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
         n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
         n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
         n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
         n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
         n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
         n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
         n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
         n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
         n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
         n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
         n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
         n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
         n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
         n2552;
  assign SUM[0] = \B[0] ;
  assign \B[0]  = B[0];

  XNOR U1 ( .A(n1), .B(n2), .Z(SUM[9]) );
  XNOR U2 ( .A(B[9]), .B(A[9]), .Z(n2) );
  XNOR U3 ( .A(n3), .B(n4), .Z(SUM[99]) );
  XNOR U4 ( .A(B[99]), .B(A[99]), .Z(n4) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[98]) );
  XNOR U6 ( .A(B[98]), .B(A[98]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(SUM[97]) );
  XNOR U8 ( .A(B[97]), .B(A[97]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(SUM[96]) );
  XNOR U10 ( .A(B[96]), .B(A[96]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(SUM[95]) );
  XNOR U12 ( .A(B[95]), .B(A[95]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(SUM[94]) );
  XNOR U14 ( .A(B[94]), .B(A[94]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(SUM[93]) );
  XNOR U16 ( .A(B[93]), .B(A[93]), .Z(n16) );
  XOR U17 ( .A(n17), .B(n18), .Z(SUM[92]) );
  XNOR U18 ( .A(B[92]), .B(A[92]), .Z(n18) );
  XOR U19 ( .A(n19), .B(n20), .Z(SUM[91]) );
  XNOR U20 ( .A(B[91]), .B(A[91]), .Z(n20) );
  XOR U21 ( .A(n21), .B(n22), .Z(SUM[90]) );
  XNOR U22 ( .A(B[90]), .B(A[90]), .Z(n22) );
  XOR U23 ( .A(n23), .B(n24), .Z(SUM[8]) );
  XNOR U24 ( .A(B[8]), .B(A[8]), .Z(n24) );
  XOR U25 ( .A(n25), .B(n26), .Z(SUM[89]) );
  XNOR U26 ( .A(B[89]), .B(A[89]), .Z(n26) );
  XOR U27 ( .A(n27), .B(n28), .Z(SUM[88]) );
  XNOR U28 ( .A(B[88]), .B(A[88]), .Z(n28) );
  XOR U29 ( .A(n29), .B(n30), .Z(SUM[87]) );
  XNOR U30 ( .A(B[87]), .B(A[87]), .Z(n30) );
  XOR U31 ( .A(n31), .B(n32), .Z(SUM[86]) );
  XNOR U32 ( .A(B[86]), .B(A[86]), .Z(n32) );
  XOR U33 ( .A(n33), .B(n34), .Z(SUM[85]) );
  XNOR U34 ( .A(B[85]), .B(A[85]), .Z(n34) );
  XOR U35 ( .A(n35), .B(n36), .Z(SUM[84]) );
  XNOR U36 ( .A(B[84]), .B(A[84]), .Z(n36) );
  XOR U37 ( .A(n37), .B(n38), .Z(SUM[83]) );
  XNOR U38 ( .A(B[83]), .B(A[83]), .Z(n38) );
  XOR U39 ( .A(n39), .B(n40), .Z(SUM[82]) );
  XNOR U40 ( .A(B[82]), .B(A[82]), .Z(n40) );
  XOR U41 ( .A(n41), .B(n42), .Z(SUM[81]) );
  XNOR U42 ( .A(B[81]), .B(A[81]), .Z(n42) );
  XOR U43 ( .A(n43), .B(n44), .Z(SUM[80]) );
  XNOR U44 ( .A(B[80]), .B(A[80]), .Z(n44) );
  XOR U45 ( .A(n45), .B(n46), .Z(SUM[7]) );
  XNOR U46 ( .A(B[7]), .B(A[7]), .Z(n46) );
  XOR U47 ( .A(n47), .B(n48), .Z(SUM[79]) );
  XNOR U48 ( .A(B[79]), .B(A[79]), .Z(n48) );
  XOR U49 ( .A(n49), .B(n50), .Z(SUM[78]) );
  XNOR U50 ( .A(B[78]), .B(A[78]), .Z(n50) );
  XOR U51 ( .A(n51), .B(n52), .Z(SUM[77]) );
  XNOR U52 ( .A(B[77]), .B(A[77]), .Z(n52) );
  XOR U53 ( .A(n53), .B(n54), .Z(SUM[76]) );
  XNOR U54 ( .A(B[76]), .B(A[76]), .Z(n54) );
  XOR U55 ( .A(n55), .B(n56), .Z(SUM[75]) );
  XNOR U56 ( .A(B[75]), .B(A[75]), .Z(n56) );
  XOR U57 ( .A(n57), .B(n58), .Z(SUM[74]) );
  XNOR U58 ( .A(B[74]), .B(A[74]), .Z(n58) );
  XOR U59 ( .A(n59), .B(n60), .Z(SUM[73]) );
  XNOR U60 ( .A(B[73]), .B(A[73]), .Z(n60) );
  XOR U61 ( .A(n61), .B(n62), .Z(SUM[72]) );
  XNOR U62 ( .A(B[72]), .B(A[72]), .Z(n62) );
  XOR U63 ( .A(n63), .B(n64), .Z(SUM[71]) );
  XNOR U64 ( .A(B[71]), .B(A[71]), .Z(n64) );
  XOR U65 ( .A(n65), .B(n66), .Z(SUM[70]) );
  XNOR U66 ( .A(B[70]), .B(A[70]), .Z(n66) );
  XOR U67 ( .A(n67), .B(n68), .Z(SUM[6]) );
  XNOR U68 ( .A(B[6]), .B(A[6]), .Z(n68) );
  XOR U69 ( .A(n69), .B(n70), .Z(SUM[69]) );
  XNOR U70 ( .A(B[69]), .B(A[69]), .Z(n70) );
  XOR U71 ( .A(n71), .B(n72), .Z(SUM[68]) );
  XNOR U72 ( .A(B[68]), .B(A[68]), .Z(n72) );
  XOR U73 ( .A(n73), .B(n74), .Z(SUM[67]) );
  XNOR U74 ( .A(B[67]), .B(A[67]), .Z(n74) );
  XOR U75 ( .A(n75), .B(n76), .Z(SUM[66]) );
  XNOR U76 ( .A(B[66]), .B(A[66]), .Z(n76) );
  XOR U77 ( .A(n77), .B(n78), .Z(SUM[65]) );
  XNOR U78 ( .A(B[65]), .B(A[65]), .Z(n78) );
  XOR U79 ( .A(n79), .B(n80), .Z(SUM[64]) );
  XNOR U80 ( .A(B[64]), .B(A[64]), .Z(n80) );
  XOR U81 ( .A(n81), .B(n82), .Z(SUM[63]) );
  XNOR U82 ( .A(B[63]), .B(A[63]), .Z(n82) );
  XOR U83 ( .A(n83), .B(n84), .Z(SUM[62]) );
  XNOR U84 ( .A(B[62]), .B(A[62]), .Z(n84) );
  XOR U85 ( .A(n85), .B(n86), .Z(SUM[61]) );
  XNOR U86 ( .A(B[61]), .B(A[61]), .Z(n86) );
  XOR U87 ( .A(n87), .B(n88), .Z(SUM[60]) );
  XNOR U88 ( .A(B[60]), .B(A[60]), .Z(n88) );
  XOR U89 ( .A(n89), .B(n90), .Z(SUM[5]) );
  XNOR U90 ( .A(B[5]), .B(A[5]), .Z(n90) );
  XOR U91 ( .A(n91), .B(n92), .Z(SUM[59]) );
  XNOR U92 ( .A(B[59]), .B(A[59]), .Z(n92) );
  XOR U93 ( .A(n93), .B(n94), .Z(SUM[58]) );
  XNOR U94 ( .A(B[58]), .B(A[58]), .Z(n94) );
  XOR U95 ( .A(n95), .B(n96), .Z(SUM[57]) );
  XNOR U96 ( .A(B[57]), .B(A[57]), .Z(n96) );
  XOR U97 ( .A(n97), .B(n98), .Z(SUM[56]) );
  XNOR U98 ( .A(B[56]), .B(A[56]), .Z(n98) );
  XOR U99 ( .A(n99), .B(n100), .Z(SUM[55]) );
  XNOR U100 ( .A(B[55]), .B(A[55]), .Z(n100) );
  XOR U101 ( .A(n101), .B(n102), .Z(SUM[54]) );
  XNOR U102 ( .A(B[54]), .B(A[54]), .Z(n102) );
  XOR U103 ( .A(n103), .B(n104), .Z(SUM[53]) );
  XNOR U104 ( .A(B[53]), .B(A[53]), .Z(n104) );
  XOR U105 ( .A(n105), .B(n106), .Z(SUM[52]) );
  XNOR U106 ( .A(B[52]), .B(A[52]), .Z(n106) );
  XOR U107 ( .A(n107), .B(n108), .Z(SUM[51]) );
  XNOR U108 ( .A(B[51]), .B(A[51]), .Z(n108) );
  XOR U109 ( .A(A[513]), .B(n109), .Z(SUM[513]) );
  AND U110 ( .A(A[512]), .B(n110), .Z(n109) );
  XOR U111 ( .A(A[512]), .B(n110), .Z(SUM[512]) );
  NAND U112 ( .A(n111), .B(n112), .Z(n110) );
  NAND U113 ( .A(B[511]), .B(n113), .Z(n112) );
  NANDN U114 ( .A(A[511]), .B(n114), .Z(n113) );
  NANDN U115 ( .A(n114), .B(A[511]), .Z(n111) );
  XOR U116 ( .A(n114), .B(n115), .Z(SUM[511]) );
  XNOR U117 ( .A(B[511]), .B(A[511]), .Z(n115) );
  AND U118 ( .A(n116), .B(n117), .Z(n114) );
  NAND U119 ( .A(B[510]), .B(n118), .Z(n117) );
  NANDN U120 ( .A(A[510]), .B(n119), .Z(n118) );
  NANDN U121 ( .A(n119), .B(A[510]), .Z(n116) );
  XOR U122 ( .A(n119), .B(n120), .Z(SUM[510]) );
  XNOR U123 ( .A(B[510]), .B(A[510]), .Z(n120) );
  AND U124 ( .A(n121), .B(n122), .Z(n119) );
  NAND U125 ( .A(B[509]), .B(n123), .Z(n122) );
  NANDN U126 ( .A(A[509]), .B(n124), .Z(n123) );
  NANDN U127 ( .A(n124), .B(A[509]), .Z(n121) );
  XOR U128 ( .A(n125), .B(n126), .Z(SUM[50]) );
  XNOR U129 ( .A(B[50]), .B(A[50]), .Z(n126) );
  XOR U130 ( .A(n124), .B(n127), .Z(SUM[509]) );
  XNOR U131 ( .A(B[509]), .B(A[509]), .Z(n127) );
  AND U132 ( .A(n128), .B(n129), .Z(n124) );
  NAND U133 ( .A(B[508]), .B(n130), .Z(n129) );
  NANDN U134 ( .A(A[508]), .B(n131), .Z(n130) );
  NANDN U135 ( .A(n131), .B(A[508]), .Z(n128) );
  XOR U136 ( .A(n131), .B(n132), .Z(SUM[508]) );
  XNOR U137 ( .A(B[508]), .B(A[508]), .Z(n132) );
  AND U138 ( .A(n133), .B(n134), .Z(n131) );
  NAND U139 ( .A(B[507]), .B(n135), .Z(n134) );
  NANDN U140 ( .A(A[507]), .B(n136), .Z(n135) );
  NANDN U141 ( .A(n136), .B(A[507]), .Z(n133) );
  XOR U142 ( .A(n136), .B(n137), .Z(SUM[507]) );
  XNOR U143 ( .A(B[507]), .B(A[507]), .Z(n137) );
  AND U144 ( .A(n138), .B(n139), .Z(n136) );
  NAND U145 ( .A(B[506]), .B(n140), .Z(n139) );
  NANDN U146 ( .A(A[506]), .B(n141), .Z(n140) );
  NANDN U147 ( .A(n141), .B(A[506]), .Z(n138) );
  XOR U148 ( .A(n141), .B(n142), .Z(SUM[506]) );
  XNOR U149 ( .A(B[506]), .B(A[506]), .Z(n142) );
  AND U150 ( .A(n143), .B(n144), .Z(n141) );
  NAND U151 ( .A(B[505]), .B(n145), .Z(n144) );
  NANDN U152 ( .A(A[505]), .B(n146), .Z(n145) );
  NANDN U153 ( .A(n146), .B(A[505]), .Z(n143) );
  XOR U154 ( .A(n146), .B(n147), .Z(SUM[505]) );
  XNOR U155 ( .A(B[505]), .B(A[505]), .Z(n147) );
  AND U156 ( .A(n148), .B(n149), .Z(n146) );
  NAND U157 ( .A(B[504]), .B(n150), .Z(n149) );
  NANDN U158 ( .A(A[504]), .B(n151), .Z(n150) );
  NANDN U159 ( .A(n151), .B(A[504]), .Z(n148) );
  XOR U160 ( .A(n151), .B(n152), .Z(SUM[504]) );
  XNOR U161 ( .A(B[504]), .B(A[504]), .Z(n152) );
  AND U162 ( .A(n153), .B(n154), .Z(n151) );
  NAND U163 ( .A(B[503]), .B(n155), .Z(n154) );
  NANDN U164 ( .A(A[503]), .B(n156), .Z(n155) );
  NANDN U165 ( .A(n156), .B(A[503]), .Z(n153) );
  XOR U166 ( .A(n156), .B(n157), .Z(SUM[503]) );
  XNOR U167 ( .A(B[503]), .B(A[503]), .Z(n157) );
  AND U168 ( .A(n158), .B(n159), .Z(n156) );
  NAND U169 ( .A(B[502]), .B(n160), .Z(n159) );
  NANDN U170 ( .A(A[502]), .B(n161), .Z(n160) );
  NANDN U171 ( .A(n161), .B(A[502]), .Z(n158) );
  XOR U172 ( .A(n161), .B(n162), .Z(SUM[502]) );
  XNOR U173 ( .A(B[502]), .B(A[502]), .Z(n162) );
  AND U174 ( .A(n163), .B(n164), .Z(n161) );
  NAND U175 ( .A(B[501]), .B(n165), .Z(n164) );
  NANDN U176 ( .A(A[501]), .B(n166), .Z(n165) );
  NANDN U177 ( .A(n166), .B(A[501]), .Z(n163) );
  XOR U178 ( .A(n166), .B(n167), .Z(SUM[501]) );
  XNOR U179 ( .A(B[501]), .B(A[501]), .Z(n167) );
  AND U180 ( .A(n168), .B(n169), .Z(n166) );
  NAND U181 ( .A(B[500]), .B(n170), .Z(n169) );
  NANDN U182 ( .A(A[500]), .B(n171), .Z(n170) );
  NANDN U183 ( .A(n171), .B(A[500]), .Z(n168) );
  XOR U184 ( .A(n171), .B(n172), .Z(SUM[500]) );
  XNOR U185 ( .A(B[500]), .B(A[500]), .Z(n172) );
  AND U186 ( .A(n173), .B(n174), .Z(n171) );
  NAND U187 ( .A(B[499]), .B(n175), .Z(n174) );
  NANDN U188 ( .A(A[499]), .B(n176), .Z(n175) );
  NANDN U189 ( .A(n176), .B(A[499]), .Z(n173) );
  XOR U190 ( .A(n177), .B(n178), .Z(SUM[4]) );
  XNOR U191 ( .A(B[4]), .B(A[4]), .Z(n178) );
  XOR U192 ( .A(n179), .B(n180), .Z(SUM[49]) );
  XNOR U193 ( .A(B[49]), .B(A[49]), .Z(n180) );
  XOR U194 ( .A(n176), .B(n181), .Z(SUM[499]) );
  XNOR U195 ( .A(B[499]), .B(A[499]), .Z(n181) );
  AND U196 ( .A(n182), .B(n183), .Z(n176) );
  NAND U197 ( .A(B[498]), .B(n184), .Z(n183) );
  NANDN U198 ( .A(A[498]), .B(n185), .Z(n184) );
  NANDN U199 ( .A(n185), .B(A[498]), .Z(n182) );
  XOR U200 ( .A(n185), .B(n186), .Z(SUM[498]) );
  XNOR U201 ( .A(B[498]), .B(A[498]), .Z(n186) );
  AND U202 ( .A(n187), .B(n188), .Z(n185) );
  NAND U203 ( .A(B[497]), .B(n189), .Z(n188) );
  NANDN U204 ( .A(A[497]), .B(n190), .Z(n189) );
  NANDN U205 ( .A(n190), .B(A[497]), .Z(n187) );
  XOR U206 ( .A(n190), .B(n191), .Z(SUM[497]) );
  XNOR U207 ( .A(B[497]), .B(A[497]), .Z(n191) );
  AND U208 ( .A(n192), .B(n193), .Z(n190) );
  NAND U209 ( .A(B[496]), .B(n194), .Z(n193) );
  NANDN U210 ( .A(A[496]), .B(n195), .Z(n194) );
  NANDN U211 ( .A(n195), .B(A[496]), .Z(n192) );
  XOR U212 ( .A(n195), .B(n196), .Z(SUM[496]) );
  XNOR U213 ( .A(B[496]), .B(A[496]), .Z(n196) );
  AND U214 ( .A(n197), .B(n198), .Z(n195) );
  NAND U215 ( .A(B[495]), .B(n199), .Z(n198) );
  NANDN U216 ( .A(A[495]), .B(n200), .Z(n199) );
  NANDN U217 ( .A(n200), .B(A[495]), .Z(n197) );
  XOR U218 ( .A(n200), .B(n201), .Z(SUM[495]) );
  XNOR U219 ( .A(B[495]), .B(A[495]), .Z(n201) );
  AND U220 ( .A(n202), .B(n203), .Z(n200) );
  NAND U221 ( .A(B[494]), .B(n204), .Z(n203) );
  NANDN U222 ( .A(A[494]), .B(n205), .Z(n204) );
  NANDN U223 ( .A(n205), .B(A[494]), .Z(n202) );
  XOR U224 ( .A(n205), .B(n206), .Z(SUM[494]) );
  XNOR U225 ( .A(B[494]), .B(A[494]), .Z(n206) );
  AND U226 ( .A(n207), .B(n208), .Z(n205) );
  NAND U227 ( .A(B[493]), .B(n209), .Z(n208) );
  NANDN U228 ( .A(A[493]), .B(n210), .Z(n209) );
  NANDN U229 ( .A(n210), .B(A[493]), .Z(n207) );
  XOR U230 ( .A(n210), .B(n211), .Z(SUM[493]) );
  XNOR U231 ( .A(B[493]), .B(A[493]), .Z(n211) );
  AND U232 ( .A(n212), .B(n213), .Z(n210) );
  NAND U233 ( .A(B[492]), .B(n214), .Z(n213) );
  NANDN U234 ( .A(A[492]), .B(n215), .Z(n214) );
  NANDN U235 ( .A(n215), .B(A[492]), .Z(n212) );
  XOR U236 ( .A(n215), .B(n216), .Z(SUM[492]) );
  XNOR U237 ( .A(B[492]), .B(A[492]), .Z(n216) );
  AND U238 ( .A(n217), .B(n218), .Z(n215) );
  NAND U239 ( .A(B[491]), .B(n219), .Z(n218) );
  NANDN U240 ( .A(A[491]), .B(n220), .Z(n219) );
  NANDN U241 ( .A(n220), .B(A[491]), .Z(n217) );
  XOR U242 ( .A(n220), .B(n221), .Z(SUM[491]) );
  XNOR U243 ( .A(B[491]), .B(A[491]), .Z(n221) );
  AND U244 ( .A(n222), .B(n223), .Z(n220) );
  NAND U245 ( .A(B[490]), .B(n224), .Z(n223) );
  NANDN U246 ( .A(A[490]), .B(n225), .Z(n224) );
  NANDN U247 ( .A(n225), .B(A[490]), .Z(n222) );
  XOR U248 ( .A(n225), .B(n226), .Z(SUM[490]) );
  XNOR U249 ( .A(B[490]), .B(A[490]), .Z(n226) );
  AND U250 ( .A(n227), .B(n228), .Z(n225) );
  NAND U251 ( .A(B[489]), .B(n229), .Z(n228) );
  NANDN U252 ( .A(A[489]), .B(n230), .Z(n229) );
  NANDN U253 ( .A(n230), .B(A[489]), .Z(n227) );
  XOR U254 ( .A(n231), .B(n232), .Z(SUM[48]) );
  XNOR U255 ( .A(B[48]), .B(A[48]), .Z(n232) );
  XOR U256 ( .A(n230), .B(n233), .Z(SUM[489]) );
  XNOR U257 ( .A(B[489]), .B(A[489]), .Z(n233) );
  AND U258 ( .A(n234), .B(n235), .Z(n230) );
  NAND U259 ( .A(B[488]), .B(n236), .Z(n235) );
  NANDN U260 ( .A(A[488]), .B(n237), .Z(n236) );
  NANDN U261 ( .A(n237), .B(A[488]), .Z(n234) );
  XOR U262 ( .A(n237), .B(n238), .Z(SUM[488]) );
  XNOR U263 ( .A(B[488]), .B(A[488]), .Z(n238) );
  AND U264 ( .A(n239), .B(n240), .Z(n237) );
  NAND U265 ( .A(B[487]), .B(n241), .Z(n240) );
  NANDN U266 ( .A(A[487]), .B(n242), .Z(n241) );
  NANDN U267 ( .A(n242), .B(A[487]), .Z(n239) );
  XOR U268 ( .A(n242), .B(n243), .Z(SUM[487]) );
  XNOR U269 ( .A(B[487]), .B(A[487]), .Z(n243) );
  AND U270 ( .A(n244), .B(n245), .Z(n242) );
  NAND U271 ( .A(B[486]), .B(n246), .Z(n245) );
  NANDN U272 ( .A(A[486]), .B(n247), .Z(n246) );
  NANDN U273 ( .A(n247), .B(A[486]), .Z(n244) );
  XOR U274 ( .A(n247), .B(n248), .Z(SUM[486]) );
  XNOR U275 ( .A(B[486]), .B(A[486]), .Z(n248) );
  AND U276 ( .A(n249), .B(n250), .Z(n247) );
  NAND U277 ( .A(B[485]), .B(n251), .Z(n250) );
  NANDN U278 ( .A(A[485]), .B(n252), .Z(n251) );
  NANDN U279 ( .A(n252), .B(A[485]), .Z(n249) );
  XOR U280 ( .A(n252), .B(n253), .Z(SUM[485]) );
  XNOR U281 ( .A(B[485]), .B(A[485]), .Z(n253) );
  AND U282 ( .A(n254), .B(n255), .Z(n252) );
  NAND U283 ( .A(B[484]), .B(n256), .Z(n255) );
  NANDN U284 ( .A(A[484]), .B(n257), .Z(n256) );
  NANDN U285 ( .A(n257), .B(A[484]), .Z(n254) );
  XOR U286 ( .A(n257), .B(n258), .Z(SUM[484]) );
  XNOR U287 ( .A(B[484]), .B(A[484]), .Z(n258) );
  AND U288 ( .A(n259), .B(n260), .Z(n257) );
  NAND U289 ( .A(B[483]), .B(n261), .Z(n260) );
  NANDN U290 ( .A(A[483]), .B(n262), .Z(n261) );
  NANDN U291 ( .A(n262), .B(A[483]), .Z(n259) );
  XOR U292 ( .A(n262), .B(n263), .Z(SUM[483]) );
  XNOR U293 ( .A(B[483]), .B(A[483]), .Z(n263) );
  AND U294 ( .A(n264), .B(n265), .Z(n262) );
  NAND U295 ( .A(B[482]), .B(n266), .Z(n265) );
  NANDN U296 ( .A(A[482]), .B(n267), .Z(n266) );
  NANDN U297 ( .A(n267), .B(A[482]), .Z(n264) );
  XOR U298 ( .A(n267), .B(n268), .Z(SUM[482]) );
  XNOR U299 ( .A(B[482]), .B(A[482]), .Z(n268) );
  AND U300 ( .A(n269), .B(n270), .Z(n267) );
  NAND U301 ( .A(B[481]), .B(n271), .Z(n270) );
  NANDN U302 ( .A(A[481]), .B(n272), .Z(n271) );
  NANDN U303 ( .A(n272), .B(A[481]), .Z(n269) );
  XOR U304 ( .A(n272), .B(n273), .Z(SUM[481]) );
  XNOR U305 ( .A(B[481]), .B(A[481]), .Z(n273) );
  AND U306 ( .A(n274), .B(n275), .Z(n272) );
  NAND U307 ( .A(B[480]), .B(n276), .Z(n275) );
  NANDN U308 ( .A(A[480]), .B(n277), .Z(n276) );
  NANDN U309 ( .A(n277), .B(A[480]), .Z(n274) );
  XOR U310 ( .A(n277), .B(n278), .Z(SUM[480]) );
  XNOR U311 ( .A(B[480]), .B(A[480]), .Z(n278) );
  AND U312 ( .A(n279), .B(n280), .Z(n277) );
  NAND U313 ( .A(B[479]), .B(n281), .Z(n280) );
  NANDN U314 ( .A(A[479]), .B(n282), .Z(n281) );
  NANDN U315 ( .A(n282), .B(A[479]), .Z(n279) );
  XOR U316 ( .A(n283), .B(n284), .Z(SUM[47]) );
  XNOR U317 ( .A(B[47]), .B(A[47]), .Z(n284) );
  XOR U318 ( .A(n282), .B(n285), .Z(SUM[479]) );
  XNOR U319 ( .A(B[479]), .B(A[479]), .Z(n285) );
  AND U320 ( .A(n286), .B(n287), .Z(n282) );
  NAND U321 ( .A(B[478]), .B(n288), .Z(n287) );
  NANDN U322 ( .A(A[478]), .B(n289), .Z(n288) );
  NANDN U323 ( .A(n289), .B(A[478]), .Z(n286) );
  XOR U324 ( .A(n289), .B(n290), .Z(SUM[478]) );
  XNOR U325 ( .A(B[478]), .B(A[478]), .Z(n290) );
  AND U326 ( .A(n291), .B(n292), .Z(n289) );
  NAND U327 ( .A(B[477]), .B(n293), .Z(n292) );
  NANDN U328 ( .A(A[477]), .B(n294), .Z(n293) );
  NANDN U329 ( .A(n294), .B(A[477]), .Z(n291) );
  XOR U330 ( .A(n294), .B(n295), .Z(SUM[477]) );
  XNOR U331 ( .A(B[477]), .B(A[477]), .Z(n295) );
  AND U332 ( .A(n296), .B(n297), .Z(n294) );
  NAND U333 ( .A(B[476]), .B(n298), .Z(n297) );
  NANDN U334 ( .A(A[476]), .B(n299), .Z(n298) );
  NANDN U335 ( .A(n299), .B(A[476]), .Z(n296) );
  XOR U336 ( .A(n299), .B(n300), .Z(SUM[476]) );
  XNOR U337 ( .A(B[476]), .B(A[476]), .Z(n300) );
  AND U338 ( .A(n301), .B(n302), .Z(n299) );
  NAND U339 ( .A(B[475]), .B(n303), .Z(n302) );
  NANDN U340 ( .A(A[475]), .B(n304), .Z(n303) );
  NANDN U341 ( .A(n304), .B(A[475]), .Z(n301) );
  XOR U342 ( .A(n304), .B(n305), .Z(SUM[475]) );
  XNOR U343 ( .A(B[475]), .B(A[475]), .Z(n305) );
  AND U344 ( .A(n306), .B(n307), .Z(n304) );
  NAND U345 ( .A(B[474]), .B(n308), .Z(n307) );
  NANDN U346 ( .A(A[474]), .B(n309), .Z(n308) );
  NANDN U347 ( .A(n309), .B(A[474]), .Z(n306) );
  XOR U348 ( .A(n309), .B(n310), .Z(SUM[474]) );
  XNOR U349 ( .A(B[474]), .B(A[474]), .Z(n310) );
  AND U350 ( .A(n311), .B(n312), .Z(n309) );
  NAND U351 ( .A(B[473]), .B(n313), .Z(n312) );
  NANDN U352 ( .A(A[473]), .B(n314), .Z(n313) );
  NANDN U353 ( .A(n314), .B(A[473]), .Z(n311) );
  XOR U354 ( .A(n314), .B(n315), .Z(SUM[473]) );
  XNOR U355 ( .A(B[473]), .B(A[473]), .Z(n315) );
  AND U356 ( .A(n316), .B(n317), .Z(n314) );
  NAND U357 ( .A(B[472]), .B(n318), .Z(n317) );
  NANDN U358 ( .A(A[472]), .B(n319), .Z(n318) );
  NANDN U359 ( .A(n319), .B(A[472]), .Z(n316) );
  XOR U360 ( .A(n319), .B(n320), .Z(SUM[472]) );
  XNOR U361 ( .A(B[472]), .B(A[472]), .Z(n320) );
  AND U362 ( .A(n321), .B(n322), .Z(n319) );
  NAND U363 ( .A(B[471]), .B(n323), .Z(n322) );
  NANDN U364 ( .A(A[471]), .B(n324), .Z(n323) );
  NANDN U365 ( .A(n324), .B(A[471]), .Z(n321) );
  XOR U366 ( .A(n324), .B(n325), .Z(SUM[471]) );
  XNOR U367 ( .A(B[471]), .B(A[471]), .Z(n325) );
  AND U368 ( .A(n326), .B(n327), .Z(n324) );
  NAND U369 ( .A(B[470]), .B(n328), .Z(n327) );
  NANDN U370 ( .A(A[470]), .B(n329), .Z(n328) );
  NANDN U371 ( .A(n329), .B(A[470]), .Z(n326) );
  XOR U372 ( .A(n329), .B(n330), .Z(SUM[470]) );
  XNOR U373 ( .A(B[470]), .B(A[470]), .Z(n330) );
  AND U374 ( .A(n331), .B(n332), .Z(n329) );
  NAND U375 ( .A(B[469]), .B(n333), .Z(n332) );
  NANDN U376 ( .A(A[469]), .B(n334), .Z(n333) );
  NANDN U377 ( .A(n334), .B(A[469]), .Z(n331) );
  XOR U378 ( .A(n335), .B(n336), .Z(SUM[46]) );
  XNOR U379 ( .A(B[46]), .B(A[46]), .Z(n336) );
  XOR U380 ( .A(n334), .B(n337), .Z(SUM[469]) );
  XNOR U381 ( .A(B[469]), .B(A[469]), .Z(n337) );
  AND U382 ( .A(n338), .B(n339), .Z(n334) );
  NAND U383 ( .A(B[468]), .B(n340), .Z(n339) );
  NANDN U384 ( .A(A[468]), .B(n341), .Z(n340) );
  NANDN U385 ( .A(n341), .B(A[468]), .Z(n338) );
  XOR U386 ( .A(n341), .B(n342), .Z(SUM[468]) );
  XNOR U387 ( .A(B[468]), .B(A[468]), .Z(n342) );
  AND U388 ( .A(n343), .B(n344), .Z(n341) );
  NAND U389 ( .A(B[467]), .B(n345), .Z(n344) );
  NANDN U390 ( .A(A[467]), .B(n346), .Z(n345) );
  NANDN U391 ( .A(n346), .B(A[467]), .Z(n343) );
  XOR U392 ( .A(n346), .B(n347), .Z(SUM[467]) );
  XNOR U393 ( .A(B[467]), .B(A[467]), .Z(n347) );
  AND U394 ( .A(n348), .B(n349), .Z(n346) );
  NAND U395 ( .A(B[466]), .B(n350), .Z(n349) );
  NANDN U396 ( .A(A[466]), .B(n351), .Z(n350) );
  NANDN U397 ( .A(n351), .B(A[466]), .Z(n348) );
  XOR U398 ( .A(n351), .B(n352), .Z(SUM[466]) );
  XNOR U399 ( .A(B[466]), .B(A[466]), .Z(n352) );
  AND U400 ( .A(n353), .B(n354), .Z(n351) );
  NAND U401 ( .A(B[465]), .B(n355), .Z(n354) );
  NANDN U402 ( .A(A[465]), .B(n356), .Z(n355) );
  NANDN U403 ( .A(n356), .B(A[465]), .Z(n353) );
  XOR U404 ( .A(n356), .B(n357), .Z(SUM[465]) );
  XNOR U405 ( .A(B[465]), .B(A[465]), .Z(n357) );
  AND U406 ( .A(n358), .B(n359), .Z(n356) );
  NAND U407 ( .A(B[464]), .B(n360), .Z(n359) );
  NANDN U408 ( .A(A[464]), .B(n361), .Z(n360) );
  NANDN U409 ( .A(n361), .B(A[464]), .Z(n358) );
  XOR U410 ( .A(n361), .B(n362), .Z(SUM[464]) );
  XNOR U411 ( .A(B[464]), .B(A[464]), .Z(n362) );
  AND U412 ( .A(n363), .B(n364), .Z(n361) );
  NAND U413 ( .A(B[463]), .B(n365), .Z(n364) );
  NANDN U414 ( .A(A[463]), .B(n366), .Z(n365) );
  NANDN U415 ( .A(n366), .B(A[463]), .Z(n363) );
  XOR U416 ( .A(n366), .B(n367), .Z(SUM[463]) );
  XNOR U417 ( .A(B[463]), .B(A[463]), .Z(n367) );
  AND U418 ( .A(n368), .B(n369), .Z(n366) );
  NAND U419 ( .A(B[462]), .B(n370), .Z(n369) );
  NANDN U420 ( .A(A[462]), .B(n371), .Z(n370) );
  NANDN U421 ( .A(n371), .B(A[462]), .Z(n368) );
  XOR U422 ( .A(n371), .B(n372), .Z(SUM[462]) );
  XNOR U423 ( .A(B[462]), .B(A[462]), .Z(n372) );
  AND U424 ( .A(n373), .B(n374), .Z(n371) );
  NAND U425 ( .A(B[461]), .B(n375), .Z(n374) );
  NANDN U426 ( .A(A[461]), .B(n376), .Z(n375) );
  NANDN U427 ( .A(n376), .B(A[461]), .Z(n373) );
  XOR U428 ( .A(n376), .B(n377), .Z(SUM[461]) );
  XNOR U429 ( .A(B[461]), .B(A[461]), .Z(n377) );
  AND U430 ( .A(n378), .B(n379), .Z(n376) );
  NAND U431 ( .A(B[460]), .B(n380), .Z(n379) );
  NANDN U432 ( .A(A[460]), .B(n381), .Z(n380) );
  NANDN U433 ( .A(n381), .B(A[460]), .Z(n378) );
  XOR U434 ( .A(n381), .B(n382), .Z(SUM[460]) );
  XNOR U435 ( .A(B[460]), .B(A[460]), .Z(n382) );
  AND U436 ( .A(n383), .B(n384), .Z(n381) );
  NAND U437 ( .A(B[459]), .B(n385), .Z(n384) );
  NANDN U438 ( .A(A[459]), .B(n386), .Z(n385) );
  NANDN U439 ( .A(n386), .B(A[459]), .Z(n383) );
  XOR U440 ( .A(n387), .B(n388), .Z(SUM[45]) );
  XNOR U441 ( .A(B[45]), .B(A[45]), .Z(n388) );
  XOR U442 ( .A(n386), .B(n389), .Z(SUM[459]) );
  XNOR U443 ( .A(B[459]), .B(A[459]), .Z(n389) );
  AND U444 ( .A(n390), .B(n391), .Z(n386) );
  NAND U445 ( .A(B[458]), .B(n392), .Z(n391) );
  NANDN U446 ( .A(A[458]), .B(n393), .Z(n392) );
  NANDN U447 ( .A(n393), .B(A[458]), .Z(n390) );
  XOR U448 ( .A(n393), .B(n394), .Z(SUM[458]) );
  XNOR U449 ( .A(B[458]), .B(A[458]), .Z(n394) );
  AND U450 ( .A(n395), .B(n396), .Z(n393) );
  NAND U451 ( .A(B[457]), .B(n397), .Z(n396) );
  NANDN U452 ( .A(A[457]), .B(n398), .Z(n397) );
  NANDN U453 ( .A(n398), .B(A[457]), .Z(n395) );
  XOR U454 ( .A(n398), .B(n399), .Z(SUM[457]) );
  XNOR U455 ( .A(B[457]), .B(A[457]), .Z(n399) );
  AND U456 ( .A(n400), .B(n401), .Z(n398) );
  NAND U457 ( .A(B[456]), .B(n402), .Z(n401) );
  NANDN U458 ( .A(A[456]), .B(n403), .Z(n402) );
  NANDN U459 ( .A(n403), .B(A[456]), .Z(n400) );
  XOR U460 ( .A(n403), .B(n404), .Z(SUM[456]) );
  XNOR U461 ( .A(B[456]), .B(A[456]), .Z(n404) );
  AND U462 ( .A(n405), .B(n406), .Z(n403) );
  NAND U463 ( .A(B[455]), .B(n407), .Z(n406) );
  NANDN U464 ( .A(A[455]), .B(n408), .Z(n407) );
  NANDN U465 ( .A(n408), .B(A[455]), .Z(n405) );
  XOR U466 ( .A(n408), .B(n409), .Z(SUM[455]) );
  XNOR U467 ( .A(B[455]), .B(A[455]), .Z(n409) );
  AND U468 ( .A(n410), .B(n411), .Z(n408) );
  NAND U469 ( .A(B[454]), .B(n412), .Z(n411) );
  NANDN U470 ( .A(A[454]), .B(n413), .Z(n412) );
  NANDN U471 ( .A(n413), .B(A[454]), .Z(n410) );
  XOR U472 ( .A(n413), .B(n414), .Z(SUM[454]) );
  XNOR U473 ( .A(B[454]), .B(A[454]), .Z(n414) );
  AND U474 ( .A(n415), .B(n416), .Z(n413) );
  NAND U475 ( .A(B[453]), .B(n417), .Z(n416) );
  NANDN U476 ( .A(A[453]), .B(n418), .Z(n417) );
  NANDN U477 ( .A(n418), .B(A[453]), .Z(n415) );
  XOR U478 ( .A(n418), .B(n419), .Z(SUM[453]) );
  XNOR U479 ( .A(B[453]), .B(A[453]), .Z(n419) );
  AND U480 ( .A(n420), .B(n421), .Z(n418) );
  NAND U481 ( .A(B[452]), .B(n422), .Z(n421) );
  NANDN U482 ( .A(A[452]), .B(n423), .Z(n422) );
  NANDN U483 ( .A(n423), .B(A[452]), .Z(n420) );
  XOR U484 ( .A(n423), .B(n424), .Z(SUM[452]) );
  XNOR U485 ( .A(B[452]), .B(A[452]), .Z(n424) );
  AND U486 ( .A(n425), .B(n426), .Z(n423) );
  NAND U487 ( .A(B[451]), .B(n427), .Z(n426) );
  NANDN U488 ( .A(A[451]), .B(n428), .Z(n427) );
  NANDN U489 ( .A(n428), .B(A[451]), .Z(n425) );
  XOR U490 ( .A(n428), .B(n429), .Z(SUM[451]) );
  XNOR U491 ( .A(B[451]), .B(A[451]), .Z(n429) );
  AND U492 ( .A(n430), .B(n431), .Z(n428) );
  NAND U493 ( .A(B[450]), .B(n432), .Z(n431) );
  NANDN U494 ( .A(A[450]), .B(n433), .Z(n432) );
  NANDN U495 ( .A(n433), .B(A[450]), .Z(n430) );
  XOR U496 ( .A(n433), .B(n434), .Z(SUM[450]) );
  XNOR U497 ( .A(B[450]), .B(A[450]), .Z(n434) );
  AND U498 ( .A(n435), .B(n436), .Z(n433) );
  NAND U499 ( .A(B[449]), .B(n437), .Z(n436) );
  NANDN U500 ( .A(A[449]), .B(n438), .Z(n437) );
  NANDN U501 ( .A(n438), .B(A[449]), .Z(n435) );
  XOR U502 ( .A(n439), .B(n440), .Z(SUM[44]) );
  XNOR U503 ( .A(B[44]), .B(A[44]), .Z(n440) );
  XOR U504 ( .A(n438), .B(n441), .Z(SUM[449]) );
  XNOR U505 ( .A(B[449]), .B(A[449]), .Z(n441) );
  AND U506 ( .A(n442), .B(n443), .Z(n438) );
  NAND U507 ( .A(B[448]), .B(n444), .Z(n443) );
  NANDN U508 ( .A(A[448]), .B(n445), .Z(n444) );
  NANDN U509 ( .A(n445), .B(A[448]), .Z(n442) );
  XOR U510 ( .A(n445), .B(n446), .Z(SUM[448]) );
  XNOR U511 ( .A(B[448]), .B(A[448]), .Z(n446) );
  AND U512 ( .A(n447), .B(n448), .Z(n445) );
  NAND U513 ( .A(B[447]), .B(n449), .Z(n448) );
  NANDN U514 ( .A(A[447]), .B(n450), .Z(n449) );
  NANDN U515 ( .A(n450), .B(A[447]), .Z(n447) );
  XOR U516 ( .A(n450), .B(n451), .Z(SUM[447]) );
  XNOR U517 ( .A(B[447]), .B(A[447]), .Z(n451) );
  AND U518 ( .A(n452), .B(n453), .Z(n450) );
  NAND U519 ( .A(B[446]), .B(n454), .Z(n453) );
  NANDN U520 ( .A(A[446]), .B(n455), .Z(n454) );
  NANDN U521 ( .A(n455), .B(A[446]), .Z(n452) );
  XOR U522 ( .A(n455), .B(n456), .Z(SUM[446]) );
  XNOR U523 ( .A(B[446]), .B(A[446]), .Z(n456) );
  AND U524 ( .A(n457), .B(n458), .Z(n455) );
  NAND U525 ( .A(B[445]), .B(n459), .Z(n458) );
  NANDN U526 ( .A(A[445]), .B(n460), .Z(n459) );
  NANDN U527 ( .A(n460), .B(A[445]), .Z(n457) );
  XOR U528 ( .A(n460), .B(n461), .Z(SUM[445]) );
  XNOR U529 ( .A(B[445]), .B(A[445]), .Z(n461) );
  AND U530 ( .A(n462), .B(n463), .Z(n460) );
  NAND U531 ( .A(B[444]), .B(n464), .Z(n463) );
  NANDN U532 ( .A(A[444]), .B(n465), .Z(n464) );
  NANDN U533 ( .A(n465), .B(A[444]), .Z(n462) );
  XOR U534 ( .A(n465), .B(n466), .Z(SUM[444]) );
  XNOR U535 ( .A(B[444]), .B(A[444]), .Z(n466) );
  AND U536 ( .A(n467), .B(n468), .Z(n465) );
  NAND U537 ( .A(B[443]), .B(n469), .Z(n468) );
  NANDN U538 ( .A(A[443]), .B(n470), .Z(n469) );
  NANDN U539 ( .A(n470), .B(A[443]), .Z(n467) );
  XOR U540 ( .A(n470), .B(n471), .Z(SUM[443]) );
  XNOR U541 ( .A(B[443]), .B(A[443]), .Z(n471) );
  AND U542 ( .A(n472), .B(n473), .Z(n470) );
  NAND U543 ( .A(B[442]), .B(n474), .Z(n473) );
  NANDN U544 ( .A(A[442]), .B(n475), .Z(n474) );
  NANDN U545 ( .A(n475), .B(A[442]), .Z(n472) );
  XOR U546 ( .A(n475), .B(n476), .Z(SUM[442]) );
  XNOR U547 ( .A(B[442]), .B(A[442]), .Z(n476) );
  AND U548 ( .A(n477), .B(n478), .Z(n475) );
  NAND U549 ( .A(B[441]), .B(n479), .Z(n478) );
  NANDN U550 ( .A(A[441]), .B(n480), .Z(n479) );
  NANDN U551 ( .A(n480), .B(A[441]), .Z(n477) );
  XOR U552 ( .A(n480), .B(n481), .Z(SUM[441]) );
  XNOR U553 ( .A(B[441]), .B(A[441]), .Z(n481) );
  AND U554 ( .A(n482), .B(n483), .Z(n480) );
  NAND U555 ( .A(B[440]), .B(n484), .Z(n483) );
  NANDN U556 ( .A(A[440]), .B(n485), .Z(n484) );
  NANDN U557 ( .A(n485), .B(A[440]), .Z(n482) );
  XOR U558 ( .A(n485), .B(n486), .Z(SUM[440]) );
  XNOR U559 ( .A(B[440]), .B(A[440]), .Z(n486) );
  AND U560 ( .A(n487), .B(n488), .Z(n485) );
  NAND U561 ( .A(B[439]), .B(n489), .Z(n488) );
  NANDN U562 ( .A(A[439]), .B(n490), .Z(n489) );
  NANDN U563 ( .A(n490), .B(A[439]), .Z(n487) );
  XOR U564 ( .A(n491), .B(n492), .Z(SUM[43]) );
  XNOR U565 ( .A(B[43]), .B(A[43]), .Z(n492) );
  XOR U566 ( .A(n490), .B(n493), .Z(SUM[439]) );
  XNOR U567 ( .A(B[439]), .B(A[439]), .Z(n493) );
  AND U568 ( .A(n494), .B(n495), .Z(n490) );
  NAND U569 ( .A(B[438]), .B(n496), .Z(n495) );
  NANDN U570 ( .A(A[438]), .B(n497), .Z(n496) );
  NANDN U571 ( .A(n497), .B(A[438]), .Z(n494) );
  XOR U572 ( .A(n497), .B(n498), .Z(SUM[438]) );
  XNOR U573 ( .A(B[438]), .B(A[438]), .Z(n498) );
  AND U574 ( .A(n499), .B(n500), .Z(n497) );
  NAND U575 ( .A(B[437]), .B(n501), .Z(n500) );
  NANDN U576 ( .A(A[437]), .B(n502), .Z(n501) );
  NANDN U577 ( .A(n502), .B(A[437]), .Z(n499) );
  XOR U578 ( .A(n502), .B(n503), .Z(SUM[437]) );
  XNOR U579 ( .A(B[437]), .B(A[437]), .Z(n503) );
  AND U580 ( .A(n504), .B(n505), .Z(n502) );
  NAND U581 ( .A(B[436]), .B(n506), .Z(n505) );
  NANDN U582 ( .A(A[436]), .B(n507), .Z(n506) );
  NANDN U583 ( .A(n507), .B(A[436]), .Z(n504) );
  XOR U584 ( .A(n507), .B(n508), .Z(SUM[436]) );
  XNOR U585 ( .A(B[436]), .B(A[436]), .Z(n508) );
  AND U586 ( .A(n509), .B(n510), .Z(n507) );
  NAND U587 ( .A(B[435]), .B(n511), .Z(n510) );
  NANDN U588 ( .A(A[435]), .B(n512), .Z(n511) );
  NANDN U589 ( .A(n512), .B(A[435]), .Z(n509) );
  XOR U590 ( .A(n512), .B(n513), .Z(SUM[435]) );
  XNOR U591 ( .A(B[435]), .B(A[435]), .Z(n513) );
  AND U592 ( .A(n514), .B(n515), .Z(n512) );
  NAND U593 ( .A(B[434]), .B(n516), .Z(n515) );
  NANDN U594 ( .A(A[434]), .B(n517), .Z(n516) );
  NANDN U595 ( .A(n517), .B(A[434]), .Z(n514) );
  XOR U596 ( .A(n517), .B(n518), .Z(SUM[434]) );
  XNOR U597 ( .A(B[434]), .B(A[434]), .Z(n518) );
  AND U598 ( .A(n519), .B(n520), .Z(n517) );
  NAND U599 ( .A(B[433]), .B(n521), .Z(n520) );
  NANDN U600 ( .A(A[433]), .B(n522), .Z(n521) );
  NANDN U601 ( .A(n522), .B(A[433]), .Z(n519) );
  XOR U602 ( .A(n522), .B(n523), .Z(SUM[433]) );
  XNOR U603 ( .A(B[433]), .B(A[433]), .Z(n523) );
  AND U604 ( .A(n524), .B(n525), .Z(n522) );
  NAND U605 ( .A(B[432]), .B(n526), .Z(n525) );
  NANDN U606 ( .A(A[432]), .B(n527), .Z(n526) );
  NANDN U607 ( .A(n527), .B(A[432]), .Z(n524) );
  XOR U608 ( .A(n527), .B(n528), .Z(SUM[432]) );
  XNOR U609 ( .A(B[432]), .B(A[432]), .Z(n528) );
  AND U610 ( .A(n529), .B(n530), .Z(n527) );
  NAND U611 ( .A(B[431]), .B(n531), .Z(n530) );
  NANDN U612 ( .A(A[431]), .B(n532), .Z(n531) );
  NANDN U613 ( .A(n532), .B(A[431]), .Z(n529) );
  XOR U614 ( .A(n532), .B(n533), .Z(SUM[431]) );
  XNOR U615 ( .A(B[431]), .B(A[431]), .Z(n533) );
  AND U616 ( .A(n534), .B(n535), .Z(n532) );
  NAND U617 ( .A(B[430]), .B(n536), .Z(n535) );
  NANDN U618 ( .A(A[430]), .B(n537), .Z(n536) );
  NANDN U619 ( .A(n537), .B(A[430]), .Z(n534) );
  XOR U620 ( .A(n537), .B(n538), .Z(SUM[430]) );
  XNOR U621 ( .A(B[430]), .B(A[430]), .Z(n538) );
  AND U622 ( .A(n539), .B(n540), .Z(n537) );
  NAND U623 ( .A(B[429]), .B(n541), .Z(n540) );
  NANDN U624 ( .A(A[429]), .B(n542), .Z(n541) );
  NANDN U625 ( .A(n542), .B(A[429]), .Z(n539) );
  XOR U626 ( .A(n543), .B(n544), .Z(SUM[42]) );
  XNOR U627 ( .A(B[42]), .B(A[42]), .Z(n544) );
  XOR U628 ( .A(n542), .B(n545), .Z(SUM[429]) );
  XNOR U629 ( .A(B[429]), .B(A[429]), .Z(n545) );
  AND U630 ( .A(n546), .B(n547), .Z(n542) );
  NAND U631 ( .A(B[428]), .B(n548), .Z(n547) );
  NANDN U632 ( .A(A[428]), .B(n549), .Z(n548) );
  NANDN U633 ( .A(n549), .B(A[428]), .Z(n546) );
  XOR U634 ( .A(n549), .B(n550), .Z(SUM[428]) );
  XNOR U635 ( .A(B[428]), .B(A[428]), .Z(n550) );
  AND U636 ( .A(n551), .B(n552), .Z(n549) );
  NAND U637 ( .A(B[427]), .B(n553), .Z(n552) );
  NANDN U638 ( .A(A[427]), .B(n554), .Z(n553) );
  NANDN U639 ( .A(n554), .B(A[427]), .Z(n551) );
  XOR U640 ( .A(n554), .B(n555), .Z(SUM[427]) );
  XNOR U641 ( .A(B[427]), .B(A[427]), .Z(n555) );
  AND U642 ( .A(n556), .B(n557), .Z(n554) );
  NAND U643 ( .A(B[426]), .B(n558), .Z(n557) );
  NANDN U644 ( .A(A[426]), .B(n559), .Z(n558) );
  NANDN U645 ( .A(n559), .B(A[426]), .Z(n556) );
  XOR U646 ( .A(n559), .B(n560), .Z(SUM[426]) );
  XNOR U647 ( .A(B[426]), .B(A[426]), .Z(n560) );
  AND U648 ( .A(n561), .B(n562), .Z(n559) );
  NAND U649 ( .A(B[425]), .B(n563), .Z(n562) );
  NANDN U650 ( .A(A[425]), .B(n564), .Z(n563) );
  NANDN U651 ( .A(n564), .B(A[425]), .Z(n561) );
  XOR U652 ( .A(n564), .B(n565), .Z(SUM[425]) );
  XNOR U653 ( .A(B[425]), .B(A[425]), .Z(n565) );
  AND U654 ( .A(n566), .B(n567), .Z(n564) );
  NAND U655 ( .A(B[424]), .B(n568), .Z(n567) );
  NANDN U656 ( .A(A[424]), .B(n569), .Z(n568) );
  NANDN U657 ( .A(n569), .B(A[424]), .Z(n566) );
  XOR U658 ( .A(n569), .B(n570), .Z(SUM[424]) );
  XNOR U659 ( .A(B[424]), .B(A[424]), .Z(n570) );
  AND U660 ( .A(n571), .B(n572), .Z(n569) );
  NAND U661 ( .A(B[423]), .B(n573), .Z(n572) );
  NANDN U662 ( .A(A[423]), .B(n574), .Z(n573) );
  NANDN U663 ( .A(n574), .B(A[423]), .Z(n571) );
  XOR U664 ( .A(n574), .B(n575), .Z(SUM[423]) );
  XNOR U665 ( .A(B[423]), .B(A[423]), .Z(n575) );
  AND U666 ( .A(n576), .B(n577), .Z(n574) );
  NAND U667 ( .A(B[422]), .B(n578), .Z(n577) );
  NANDN U668 ( .A(A[422]), .B(n579), .Z(n578) );
  NANDN U669 ( .A(n579), .B(A[422]), .Z(n576) );
  XOR U670 ( .A(n579), .B(n580), .Z(SUM[422]) );
  XNOR U671 ( .A(B[422]), .B(A[422]), .Z(n580) );
  AND U672 ( .A(n581), .B(n582), .Z(n579) );
  NAND U673 ( .A(B[421]), .B(n583), .Z(n582) );
  NANDN U674 ( .A(A[421]), .B(n584), .Z(n583) );
  NANDN U675 ( .A(n584), .B(A[421]), .Z(n581) );
  XOR U676 ( .A(n584), .B(n585), .Z(SUM[421]) );
  XNOR U677 ( .A(B[421]), .B(A[421]), .Z(n585) );
  AND U678 ( .A(n586), .B(n587), .Z(n584) );
  NAND U679 ( .A(B[420]), .B(n588), .Z(n587) );
  NANDN U680 ( .A(A[420]), .B(n589), .Z(n588) );
  NANDN U681 ( .A(n589), .B(A[420]), .Z(n586) );
  XOR U682 ( .A(n589), .B(n590), .Z(SUM[420]) );
  XNOR U683 ( .A(B[420]), .B(A[420]), .Z(n590) );
  AND U684 ( .A(n591), .B(n592), .Z(n589) );
  NAND U685 ( .A(B[419]), .B(n593), .Z(n592) );
  NANDN U686 ( .A(A[419]), .B(n594), .Z(n593) );
  NANDN U687 ( .A(n594), .B(A[419]), .Z(n591) );
  XOR U688 ( .A(n595), .B(n596), .Z(SUM[41]) );
  XNOR U689 ( .A(B[41]), .B(A[41]), .Z(n596) );
  XOR U690 ( .A(n594), .B(n597), .Z(SUM[419]) );
  XNOR U691 ( .A(B[419]), .B(A[419]), .Z(n597) );
  AND U692 ( .A(n598), .B(n599), .Z(n594) );
  NAND U693 ( .A(B[418]), .B(n600), .Z(n599) );
  NANDN U694 ( .A(A[418]), .B(n601), .Z(n600) );
  NANDN U695 ( .A(n601), .B(A[418]), .Z(n598) );
  XOR U696 ( .A(n601), .B(n602), .Z(SUM[418]) );
  XNOR U697 ( .A(B[418]), .B(A[418]), .Z(n602) );
  AND U698 ( .A(n603), .B(n604), .Z(n601) );
  NAND U699 ( .A(B[417]), .B(n605), .Z(n604) );
  NANDN U700 ( .A(A[417]), .B(n606), .Z(n605) );
  NANDN U701 ( .A(n606), .B(A[417]), .Z(n603) );
  XOR U702 ( .A(n606), .B(n607), .Z(SUM[417]) );
  XNOR U703 ( .A(B[417]), .B(A[417]), .Z(n607) );
  AND U704 ( .A(n608), .B(n609), .Z(n606) );
  NAND U705 ( .A(B[416]), .B(n610), .Z(n609) );
  NANDN U706 ( .A(A[416]), .B(n611), .Z(n610) );
  NANDN U707 ( .A(n611), .B(A[416]), .Z(n608) );
  XOR U708 ( .A(n611), .B(n612), .Z(SUM[416]) );
  XNOR U709 ( .A(B[416]), .B(A[416]), .Z(n612) );
  AND U710 ( .A(n613), .B(n614), .Z(n611) );
  NAND U711 ( .A(B[415]), .B(n615), .Z(n614) );
  NANDN U712 ( .A(A[415]), .B(n616), .Z(n615) );
  NANDN U713 ( .A(n616), .B(A[415]), .Z(n613) );
  XOR U714 ( .A(n616), .B(n617), .Z(SUM[415]) );
  XNOR U715 ( .A(B[415]), .B(A[415]), .Z(n617) );
  AND U716 ( .A(n618), .B(n619), .Z(n616) );
  NAND U717 ( .A(B[414]), .B(n620), .Z(n619) );
  NANDN U718 ( .A(A[414]), .B(n621), .Z(n620) );
  NANDN U719 ( .A(n621), .B(A[414]), .Z(n618) );
  XOR U720 ( .A(n621), .B(n622), .Z(SUM[414]) );
  XNOR U721 ( .A(B[414]), .B(A[414]), .Z(n622) );
  AND U722 ( .A(n623), .B(n624), .Z(n621) );
  NAND U723 ( .A(B[413]), .B(n625), .Z(n624) );
  NANDN U724 ( .A(A[413]), .B(n626), .Z(n625) );
  NANDN U725 ( .A(n626), .B(A[413]), .Z(n623) );
  XOR U726 ( .A(n626), .B(n627), .Z(SUM[413]) );
  XNOR U727 ( .A(B[413]), .B(A[413]), .Z(n627) );
  AND U728 ( .A(n628), .B(n629), .Z(n626) );
  NAND U729 ( .A(B[412]), .B(n630), .Z(n629) );
  NANDN U730 ( .A(A[412]), .B(n631), .Z(n630) );
  NANDN U731 ( .A(n631), .B(A[412]), .Z(n628) );
  XOR U732 ( .A(n631), .B(n632), .Z(SUM[412]) );
  XNOR U733 ( .A(B[412]), .B(A[412]), .Z(n632) );
  AND U734 ( .A(n633), .B(n634), .Z(n631) );
  NAND U735 ( .A(B[411]), .B(n635), .Z(n634) );
  NANDN U736 ( .A(A[411]), .B(n636), .Z(n635) );
  NANDN U737 ( .A(n636), .B(A[411]), .Z(n633) );
  XOR U738 ( .A(n636), .B(n637), .Z(SUM[411]) );
  XNOR U739 ( .A(B[411]), .B(A[411]), .Z(n637) );
  AND U740 ( .A(n638), .B(n639), .Z(n636) );
  NAND U741 ( .A(B[410]), .B(n640), .Z(n639) );
  NANDN U742 ( .A(A[410]), .B(n641), .Z(n640) );
  NANDN U743 ( .A(n641), .B(A[410]), .Z(n638) );
  XOR U744 ( .A(n641), .B(n642), .Z(SUM[410]) );
  XNOR U745 ( .A(B[410]), .B(A[410]), .Z(n642) );
  AND U746 ( .A(n643), .B(n644), .Z(n641) );
  NAND U747 ( .A(B[409]), .B(n645), .Z(n644) );
  NANDN U748 ( .A(A[409]), .B(n646), .Z(n645) );
  NANDN U749 ( .A(n646), .B(A[409]), .Z(n643) );
  XOR U750 ( .A(n647), .B(n648), .Z(SUM[40]) );
  XNOR U751 ( .A(B[40]), .B(A[40]), .Z(n648) );
  XOR U752 ( .A(n646), .B(n649), .Z(SUM[409]) );
  XNOR U753 ( .A(B[409]), .B(A[409]), .Z(n649) );
  AND U754 ( .A(n650), .B(n651), .Z(n646) );
  NAND U755 ( .A(B[408]), .B(n652), .Z(n651) );
  NANDN U756 ( .A(A[408]), .B(n653), .Z(n652) );
  NANDN U757 ( .A(n653), .B(A[408]), .Z(n650) );
  XOR U758 ( .A(n653), .B(n654), .Z(SUM[408]) );
  XNOR U759 ( .A(B[408]), .B(A[408]), .Z(n654) );
  AND U760 ( .A(n655), .B(n656), .Z(n653) );
  NAND U761 ( .A(B[407]), .B(n657), .Z(n656) );
  NANDN U762 ( .A(A[407]), .B(n658), .Z(n657) );
  NANDN U763 ( .A(n658), .B(A[407]), .Z(n655) );
  XOR U764 ( .A(n658), .B(n659), .Z(SUM[407]) );
  XNOR U765 ( .A(B[407]), .B(A[407]), .Z(n659) );
  AND U766 ( .A(n660), .B(n661), .Z(n658) );
  NAND U767 ( .A(B[406]), .B(n662), .Z(n661) );
  NANDN U768 ( .A(A[406]), .B(n663), .Z(n662) );
  NANDN U769 ( .A(n663), .B(A[406]), .Z(n660) );
  XOR U770 ( .A(n663), .B(n664), .Z(SUM[406]) );
  XNOR U771 ( .A(B[406]), .B(A[406]), .Z(n664) );
  AND U772 ( .A(n665), .B(n666), .Z(n663) );
  NAND U773 ( .A(B[405]), .B(n667), .Z(n666) );
  NANDN U774 ( .A(A[405]), .B(n668), .Z(n667) );
  NANDN U775 ( .A(n668), .B(A[405]), .Z(n665) );
  XOR U776 ( .A(n668), .B(n669), .Z(SUM[405]) );
  XNOR U777 ( .A(B[405]), .B(A[405]), .Z(n669) );
  AND U778 ( .A(n670), .B(n671), .Z(n668) );
  NAND U779 ( .A(B[404]), .B(n672), .Z(n671) );
  NANDN U780 ( .A(A[404]), .B(n673), .Z(n672) );
  NANDN U781 ( .A(n673), .B(A[404]), .Z(n670) );
  XOR U782 ( .A(n673), .B(n674), .Z(SUM[404]) );
  XNOR U783 ( .A(B[404]), .B(A[404]), .Z(n674) );
  AND U784 ( .A(n675), .B(n676), .Z(n673) );
  NAND U785 ( .A(B[403]), .B(n677), .Z(n676) );
  NANDN U786 ( .A(A[403]), .B(n678), .Z(n677) );
  NANDN U787 ( .A(n678), .B(A[403]), .Z(n675) );
  XOR U788 ( .A(n678), .B(n679), .Z(SUM[403]) );
  XNOR U789 ( .A(B[403]), .B(A[403]), .Z(n679) );
  AND U790 ( .A(n680), .B(n681), .Z(n678) );
  NAND U791 ( .A(B[402]), .B(n682), .Z(n681) );
  NANDN U792 ( .A(A[402]), .B(n683), .Z(n682) );
  NANDN U793 ( .A(n683), .B(A[402]), .Z(n680) );
  XOR U794 ( .A(n683), .B(n684), .Z(SUM[402]) );
  XNOR U795 ( .A(B[402]), .B(A[402]), .Z(n684) );
  AND U796 ( .A(n685), .B(n686), .Z(n683) );
  NAND U797 ( .A(B[401]), .B(n687), .Z(n686) );
  NANDN U798 ( .A(A[401]), .B(n688), .Z(n687) );
  NANDN U799 ( .A(n688), .B(A[401]), .Z(n685) );
  XOR U800 ( .A(n688), .B(n689), .Z(SUM[401]) );
  XNOR U801 ( .A(B[401]), .B(A[401]), .Z(n689) );
  AND U802 ( .A(n690), .B(n691), .Z(n688) );
  NAND U803 ( .A(B[400]), .B(n692), .Z(n691) );
  NANDN U804 ( .A(A[400]), .B(n693), .Z(n692) );
  NANDN U805 ( .A(n693), .B(A[400]), .Z(n690) );
  XOR U806 ( .A(n693), .B(n694), .Z(SUM[400]) );
  XNOR U807 ( .A(B[400]), .B(A[400]), .Z(n694) );
  AND U808 ( .A(n695), .B(n696), .Z(n693) );
  NAND U809 ( .A(B[399]), .B(n697), .Z(n696) );
  NANDN U810 ( .A(A[399]), .B(n698), .Z(n697) );
  NANDN U811 ( .A(n698), .B(A[399]), .Z(n695) );
  XOR U812 ( .A(n699), .B(n700), .Z(SUM[3]) );
  XNOR U813 ( .A(B[3]), .B(A[3]), .Z(n700) );
  XOR U814 ( .A(n701), .B(n702), .Z(SUM[39]) );
  XNOR U815 ( .A(B[39]), .B(A[39]), .Z(n702) );
  XOR U816 ( .A(n698), .B(n703), .Z(SUM[399]) );
  XNOR U817 ( .A(B[399]), .B(A[399]), .Z(n703) );
  AND U818 ( .A(n704), .B(n705), .Z(n698) );
  NAND U819 ( .A(B[398]), .B(n706), .Z(n705) );
  NANDN U820 ( .A(A[398]), .B(n707), .Z(n706) );
  NANDN U821 ( .A(n707), .B(A[398]), .Z(n704) );
  XOR U822 ( .A(n707), .B(n708), .Z(SUM[398]) );
  XNOR U823 ( .A(B[398]), .B(A[398]), .Z(n708) );
  AND U824 ( .A(n709), .B(n710), .Z(n707) );
  NAND U825 ( .A(B[397]), .B(n711), .Z(n710) );
  NANDN U826 ( .A(A[397]), .B(n712), .Z(n711) );
  NANDN U827 ( .A(n712), .B(A[397]), .Z(n709) );
  XOR U828 ( .A(n712), .B(n713), .Z(SUM[397]) );
  XNOR U829 ( .A(B[397]), .B(A[397]), .Z(n713) );
  AND U830 ( .A(n714), .B(n715), .Z(n712) );
  NAND U831 ( .A(B[396]), .B(n716), .Z(n715) );
  NANDN U832 ( .A(A[396]), .B(n717), .Z(n716) );
  NANDN U833 ( .A(n717), .B(A[396]), .Z(n714) );
  XOR U834 ( .A(n717), .B(n718), .Z(SUM[396]) );
  XNOR U835 ( .A(B[396]), .B(A[396]), .Z(n718) );
  AND U836 ( .A(n719), .B(n720), .Z(n717) );
  NAND U837 ( .A(B[395]), .B(n721), .Z(n720) );
  NANDN U838 ( .A(A[395]), .B(n722), .Z(n721) );
  NANDN U839 ( .A(n722), .B(A[395]), .Z(n719) );
  XOR U840 ( .A(n722), .B(n723), .Z(SUM[395]) );
  XNOR U841 ( .A(B[395]), .B(A[395]), .Z(n723) );
  AND U842 ( .A(n724), .B(n725), .Z(n722) );
  NAND U843 ( .A(B[394]), .B(n726), .Z(n725) );
  NANDN U844 ( .A(A[394]), .B(n727), .Z(n726) );
  NANDN U845 ( .A(n727), .B(A[394]), .Z(n724) );
  XOR U846 ( .A(n727), .B(n728), .Z(SUM[394]) );
  XNOR U847 ( .A(B[394]), .B(A[394]), .Z(n728) );
  AND U848 ( .A(n729), .B(n730), .Z(n727) );
  NAND U849 ( .A(B[393]), .B(n731), .Z(n730) );
  NANDN U850 ( .A(A[393]), .B(n732), .Z(n731) );
  NANDN U851 ( .A(n732), .B(A[393]), .Z(n729) );
  XOR U852 ( .A(n732), .B(n733), .Z(SUM[393]) );
  XNOR U853 ( .A(B[393]), .B(A[393]), .Z(n733) );
  AND U854 ( .A(n734), .B(n735), .Z(n732) );
  NAND U855 ( .A(B[392]), .B(n736), .Z(n735) );
  NANDN U856 ( .A(A[392]), .B(n737), .Z(n736) );
  NANDN U857 ( .A(n737), .B(A[392]), .Z(n734) );
  XOR U858 ( .A(n737), .B(n738), .Z(SUM[392]) );
  XNOR U859 ( .A(B[392]), .B(A[392]), .Z(n738) );
  AND U860 ( .A(n739), .B(n740), .Z(n737) );
  NAND U861 ( .A(B[391]), .B(n741), .Z(n740) );
  NANDN U862 ( .A(A[391]), .B(n742), .Z(n741) );
  NANDN U863 ( .A(n742), .B(A[391]), .Z(n739) );
  XOR U864 ( .A(n742), .B(n743), .Z(SUM[391]) );
  XNOR U865 ( .A(B[391]), .B(A[391]), .Z(n743) );
  AND U866 ( .A(n744), .B(n745), .Z(n742) );
  NAND U867 ( .A(B[390]), .B(n746), .Z(n745) );
  NANDN U868 ( .A(A[390]), .B(n747), .Z(n746) );
  NANDN U869 ( .A(n747), .B(A[390]), .Z(n744) );
  XOR U870 ( .A(n747), .B(n748), .Z(SUM[390]) );
  XNOR U871 ( .A(B[390]), .B(A[390]), .Z(n748) );
  AND U872 ( .A(n749), .B(n750), .Z(n747) );
  NAND U873 ( .A(B[389]), .B(n751), .Z(n750) );
  NANDN U874 ( .A(A[389]), .B(n752), .Z(n751) );
  NANDN U875 ( .A(n752), .B(A[389]), .Z(n749) );
  XOR U876 ( .A(n753), .B(n754), .Z(SUM[38]) );
  XNOR U877 ( .A(B[38]), .B(A[38]), .Z(n754) );
  XOR U878 ( .A(n752), .B(n755), .Z(SUM[389]) );
  XNOR U879 ( .A(B[389]), .B(A[389]), .Z(n755) );
  AND U880 ( .A(n756), .B(n757), .Z(n752) );
  NAND U881 ( .A(B[388]), .B(n758), .Z(n757) );
  NANDN U882 ( .A(A[388]), .B(n759), .Z(n758) );
  NANDN U883 ( .A(n759), .B(A[388]), .Z(n756) );
  XOR U884 ( .A(n759), .B(n760), .Z(SUM[388]) );
  XNOR U885 ( .A(B[388]), .B(A[388]), .Z(n760) );
  AND U886 ( .A(n761), .B(n762), .Z(n759) );
  NAND U887 ( .A(B[387]), .B(n763), .Z(n762) );
  NANDN U888 ( .A(A[387]), .B(n764), .Z(n763) );
  NANDN U889 ( .A(n764), .B(A[387]), .Z(n761) );
  XOR U890 ( .A(n764), .B(n765), .Z(SUM[387]) );
  XNOR U891 ( .A(B[387]), .B(A[387]), .Z(n765) );
  AND U892 ( .A(n766), .B(n767), .Z(n764) );
  NAND U893 ( .A(B[386]), .B(n768), .Z(n767) );
  NANDN U894 ( .A(A[386]), .B(n769), .Z(n768) );
  NANDN U895 ( .A(n769), .B(A[386]), .Z(n766) );
  XOR U896 ( .A(n769), .B(n770), .Z(SUM[386]) );
  XNOR U897 ( .A(B[386]), .B(A[386]), .Z(n770) );
  AND U898 ( .A(n771), .B(n772), .Z(n769) );
  NAND U899 ( .A(B[385]), .B(n773), .Z(n772) );
  NANDN U900 ( .A(A[385]), .B(n774), .Z(n773) );
  NANDN U901 ( .A(n774), .B(A[385]), .Z(n771) );
  XOR U902 ( .A(n774), .B(n775), .Z(SUM[385]) );
  XNOR U903 ( .A(B[385]), .B(A[385]), .Z(n775) );
  AND U904 ( .A(n776), .B(n777), .Z(n774) );
  NAND U905 ( .A(B[384]), .B(n778), .Z(n777) );
  NANDN U906 ( .A(A[384]), .B(n779), .Z(n778) );
  NANDN U907 ( .A(n779), .B(A[384]), .Z(n776) );
  XOR U908 ( .A(n779), .B(n780), .Z(SUM[384]) );
  XNOR U909 ( .A(B[384]), .B(A[384]), .Z(n780) );
  AND U910 ( .A(n781), .B(n782), .Z(n779) );
  NAND U911 ( .A(B[383]), .B(n783), .Z(n782) );
  NANDN U912 ( .A(A[383]), .B(n784), .Z(n783) );
  NANDN U913 ( .A(n784), .B(A[383]), .Z(n781) );
  XOR U914 ( .A(n784), .B(n785), .Z(SUM[383]) );
  XNOR U915 ( .A(B[383]), .B(A[383]), .Z(n785) );
  AND U916 ( .A(n786), .B(n787), .Z(n784) );
  NAND U917 ( .A(B[382]), .B(n788), .Z(n787) );
  NANDN U918 ( .A(A[382]), .B(n789), .Z(n788) );
  NANDN U919 ( .A(n789), .B(A[382]), .Z(n786) );
  XOR U920 ( .A(n789), .B(n790), .Z(SUM[382]) );
  XNOR U921 ( .A(B[382]), .B(A[382]), .Z(n790) );
  AND U922 ( .A(n791), .B(n792), .Z(n789) );
  NAND U923 ( .A(B[381]), .B(n793), .Z(n792) );
  NANDN U924 ( .A(A[381]), .B(n794), .Z(n793) );
  NANDN U925 ( .A(n794), .B(A[381]), .Z(n791) );
  XOR U926 ( .A(n794), .B(n795), .Z(SUM[381]) );
  XNOR U927 ( .A(B[381]), .B(A[381]), .Z(n795) );
  AND U928 ( .A(n796), .B(n797), .Z(n794) );
  NAND U929 ( .A(B[380]), .B(n798), .Z(n797) );
  NANDN U930 ( .A(A[380]), .B(n799), .Z(n798) );
  NANDN U931 ( .A(n799), .B(A[380]), .Z(n796) );
  XOR U932 ( .A(n799), .B(n800), .Z(SUM[380]) );
  XNOR U933 ( .A(B[380]), .B(A[380]), .Z(n800) );
  AND U934 ( .A(n801), .B(n802), .Z(n799) );
  NAND U935 ( .A(B[379]), .B(n803), .Z(n802) );
  NANDN U936 ( .A(A[379]), .B(n804), .Z(n803) );
  NANDN U937 ( .A(n804), .B(A[379]), .Z(n801) );
  XOR U938 ( .A(n805), .B(n806), .Z(SUM[37]) );
  XNOR U939 ( .A(B[37]), .B(A[37]), .Z(n806) );
  XOR U940 ( .A(n804), .B(n807), .Z(SUM[379]) );
  XNOR U941 ( .A(B[379]), .B(A[379]), .Z(n807) );
  AND U942 ( .A(n808), .B(n809), .Z(n804) );
  NAND U943 ( .A(B[378]), .B(n810), .Z(n809) );
  NANDN U944 ( .A(A[378]), .B(n811), .Z(n810) );
  NANDN U945 ( .A(n811), .B(A[378]), .Z(n808) );
  XOR U946 ( .A(n811), .B(n812), .Z(SUM[378]) );
  XNOR U947 ( .A(B[378]), .B(A[378]), .Z(n812) );
  AND U948 ( .A(n813), .B(n814), .Z(n811) );
  NAND U949 ( .A(B[377]), .B(n815), .Z(n814) );
  NANDN U950 ( .A(A[377]), .B(n816), .Z(n815) );
  NANDN U951 ( .A(n816), .B(A[377]), .Z(n813) );
  XOR U952 ( .A(n816), .B(n817), .Z(SUM[377]) );
  XNOR U953 ( .A(B[377]), .B(A[377]), .Z(n817) );
  AND U954 ( .A(n818), .B(n819), .Z(n816) );
  NAND U955 ( .A(B[376]), .B(n820), .Z(n819) );
  NANDN U956 ( .A(A[376]), .B(n821), .Z(n820) );
  NANDN U957 ( .A(n821), .B(A[376]), .Z(n818) );
  XOR U958 ( .A(n821), .B(n822), .Z(SUM[376]) );
  XNOR U959 ( .A(B[376]), .B(A[376]), .Z(n822) );
  AND U960 ( .A(n823), .B(n824), .Z(n821) );
  NAND U961 ( .A(B[375]), .B(n825), .Z(n824) );
  NANDN U962 ( .A(A[375]), .B(n826), .Z(n825) );
  NANDN U963 ( .A(n826), .B(A[375]), .Z(n823) );
  XOR U964 ( .A(n826), .B(n827), .Z(SUM[375]) );
  XNOR U965 ( .A(B[375]), .B(A[375]), .Z(n827) );
  AND U966 ( .A(n828), .B(n829), .Z(n826) );
  NAND U967 ( .A(B[374]), .B(n830), .Z(n829) );
  NANDN U968 ( .A(A[374]), .B(n831), .Z(n830) );
  NANDN U969 ( .A(n831), .B(A[374]), .Z(n828) );
  XOR U970 ( .A(n831), .B(n832), .Z(SUM[374]) );
  XNOR U971 ( .A(B[374]), .B(A[374]), .Z(n832) );
  AND U972 ( .A(n833), .B(n834), .Z(n831) );
  NAND U973 ( .A(B[373]), .B(n835), .Z(n834) );
  NANDN U974 ( .A(A[373]), .B(n836), .Z(n835) );
  NANDN U975 ( .A(n836), .B(A[373]), .Z(n833) );
  XOR U976 ( .A(n836), .B(n837), .Z(SUM[373]) );
  XNOR U977 ( .A(B[373]), .B(A[373]), .Z(n837) );
  AND U978 ( .A(n838), .B(n839), .Z(n836) );
  NAND U979 ( .A(B[372]), .B(n840), .Z(n839) );
  NANDN U980 ( .A(A[372]), .B(n841), .Z(n840) );
  NANDN U981 ( .A(n841), .B(A[372]), .Z(n838) );
  XOR U982 ( .A(n841), .B(n842), .Z(SUM[372]) );
  XNOR U983 ( .A(B[372]), .B(A[372]), .Z(n842) );
  AND U984 ( .A(n843), .B(n844), .Z(n841) );
  NAND U985 ( .A(B[371]), .B(n845), .Z(n844) );
  NANDN U986 ( .A(A[371]), .B(n846), .Z(n845) );
  NANDN U987 ( .A(n846), .B(A[371]), .Z(n843) );
  XOR U988 ( .A(n846), .B(n847), .Z(SUM[371]) );
  XNOR U989 ( .A(B[371]), .B(A[371]), .Z(n847) );
  AND U990 ( .A(n848), .B(n849), .Z(n846) );
  NAND U991 ( .A(B[370]), .B(n850), .Z(n849) );
  NANDN U992 ( .A(A[370]), .B(n851), .Z(n850) );
  NANDN U993 ( .A(n851), .B(A[370]), .Z(n848) );
  XOR U994 ( .A(n851), .B(n852), .Z(SUM[370]) );
  XNOR U995 ( .A(B[370]), .B(A[370]), .Z(n852) );
  AND U996 ( .A(n853), .B(n854), .Z(n851) );
  NAND U997 ( .A(B[369]), .B(n855), .Z(n854) );
  NANDN U998 ( .A(A[369]), .B(n856), .Z(n855) );
  NANDN U999 ( .A(n856), .B(A[369]), .Z(n853) );
  XOR U1000 ( .A(n857), .B(n858), .Z(SUM[36]) );
  XNOR U1001 ( .A(B[36]), .B(A[36]), .Z(n858) );
  XOR U1002 ( .A(n856), .B(n859), .Z(SUM[369]) );
  XNOR U1003 ( .A(B[369]), .B(A[369]), .Z(n859) );
  AND U1004 ( .A(n860), .B(n861), .Z(n856) );
  NAND U1005 ( .A(B[368]), .B(n862), .Z(n861) );
  NANDN U1006 ( .A(A[368]), .B(n863), .Z(n862) );
  NANDN U1007 ( .A(n863), .B(A[368]), .Z(n860) );
  XOR U1008 ( .A(n863), .B(n864), .Z(SUM[368]) );
  XNOR U1009 ( .A(B[368]), .B(A[368]), .Z(n864) );
  AND U1010 ( .A(n865), .B(n866), .Z(n863) );
  NAND U1011 ( .A(B[367]), .B(n867), .Z(n866) );
  NANDN U1012 ( .A(A[367]), .B(n868), .Z(n867) );
  NANDN U1013 ( .A(n868), .B(A[367]), .Z(n865) );
  XOR U1014 ( .A(n868), .B(n869), .Z(SUM[367]) );
  XNOR U1015 ( .A(B[367]), .B(A[367]), .Z(n869) );
  AND U1016 ( .A(n870), .B(n871), .Z(n868) );
  NAND U1017 ( .A(B[366]), .B(n872), .Z(n871) );
  NANDN U1018 ( .A(A[366]), .B(n873), .Z(n872) );
  NANDN U1019 ( .A(n873), .B(A[366]), .Z(n870) );
  XOR U1020 ( .A(n873), .B(n874), .Z(SUM[366]) );
  XNOR U1021 ( .A(B[366]), .B(A[366]), .Z(n874) );
  AND U1022 ( .A(n875), .B(n876), .Z(n873) );
  NAND U1023 ( .A(B[365]), .B(n877), .Z(n876) );
  NANDN U1024 ( .A(A[365]), .B(n878), .Z(n877) );
  NANDN U1025 ( .A(n878), .B(A[365]), .Z(n875) );
  XOR U1026 ( .A(n878), .B(n879), .Z(SUM[365]) );
  XNOR U1027 ( .A(B[365]), .B(A[365]), .Z(n879) );
  AND U1028 ( .A(n880), .B(n881), .Z(n878) );
  NAND U1029 ( .A(B[364]), .B(n882), .Z(n881) );
  NANDN U1030 ( .A(A[364]), .B(n883), .Z(n882) );
  NANDN U1031 ( .A(n883), .B(A[364]), .Z(n880) );
  XOR U1032 ( .A(n883), .B(n884), .Z(SUM[364]) );
  XNOR U1033 ( .A(B[364]), .B(A[364]), .Z(n884) );
  AND U1034 ( .A(n885), .B(n886), .Z(n883) );
  NAND U1035 ( .A(B[363]), .B(n887), .Z(n886) );
  NANDN U1036 ( .A(A[363]), .B(n888), .Z(n887) );
  NANDN U1037 ( .A(n888), .B(A[363]), .Z(n885) );
  XOR U1038 ( .A(n888), .B(n889), .Z(SUM[363]) );
  XNOR U1039 ( .A(B[363]), .B(A[363]), .Z(n889) );
  AND U1040 ( .A(n890), .B(n891), .Z(n888) );
  NAND U1041 ( .A(B[362]), .B(n892), .Z(n891) );
  NANDN U1042 ( .A(A[362]), .B(n893), .Z(n892) );
  NANDN U1043 ( .A(n893), .B(A[362]), .Z(n890) );
  XOR U1044 ( .A(n893), .B(n894), .Z(SUM[362]) );
  XNOR U1045 ( .A(B[362]), .B(A[362]), .Z(n894) );
  AND U1046 ( .A(n895), .B(n896), .Z(n893) );
  NAND U1047 ( .A(B[361]), .B(n897), .Z(n896) );
  NANDN U1048 ( .A(A[361]), .B(n898), .Z(n897) );
  NANDN U1049 ( .A(n898), .B(A[361]), .Z(n895) );
  XOR U1050 ( .A(n898), .B(n899), .Z(SUM[361]) );
  XNOR U1051 ( .A(B[361]), .B(A[361]), .Z(n899) );
  AND U1052 ( .A(n900), .B(n901), .Z(n898) );
  NAND U1053 ( .A(B[360]), .B(n902), .Z(n901) );
  NANDN U1054 ( .A(A[360]), .B(n903), .Z(n902) );
  NANDN U1055 ( .A(n903), .B(A[360]), .Z(n900) );
  XOR U1056 ( .A(n903), .B(n904), .Z(SUM[360]) );
  XNOR U1057 ( .A(B[360]), .B(A[360]), .Z(n904) );
  AND U1058 ( .A(n905), .B(n906), .Z(n903) );
  NAND U1059 ( .A(B[359]), .B(n907), .Z(n906) );
  NANDN U1060 ( .A(A[359]), .B(n908), .Z(n907) );
  NANDN U1061 ( .A(n908), .B(A[359]), .Z(n905) );
  XOR U1062 ( .A(n909), .B(n910), .Z(SUM[35]) );
  XNOR U1063 ( .A(B[35]), .B(A[35]), .Z(n910) );
  XOR U1064 ( .A(n908), .B(n911), .Z(SUM[359]) );
  XNOR U1065 ( .A(B[359]), .B(A[359]), .Z(n911) );
  AND U1066 ( .A(n912), .B(n913), .Z(n908) );
  NAND U1067 ( .A(B[358]), .B(n914), .Z(n913) );
  NANDN U1068 ( .A(A[358]), .B(n915), .Z(n914) );
  NANDN U1069 ( .A(n915), .B(A[358]), .Z(n912) );
  XOR U1070 ( .A(n915), .B(n916), .Z(SUM[358]) );
  XNOR U1071 ( .A(B[358]), .B(A[358]), .Z(n916) );
  AND U1072 ( .A(n917), .B(n918), .Z(n915) );
  NAND U1073 ( .A(B[357]), .B(n919), .Z(n918) );
  NANDN U1074 ( .A(A[357]), .B(n920), .Z(n919) );
  NANDN U1075 ( .A(n920), .B(A[357]), .Z(n917) );
  XOR U1076 ( .A(n920), .B(n921), .Z(SUM[357]) );
  XNOR U1077 ( .A(B[357]), .B(A[357]), .Z(n921) );
  AND U1078 ( .A(n922), .B(n923), .Z(n920) );
  NAND U1079 ( .A(B[356]), .B(n924), .Z(n923) );
  NANDN U1080 ( .A(A[356]), .B(n925), .Z(n924) );
  NANDN U1081 ( .A(n925), .B(A[356]), .Z(n922) );
  XOR U1082 ( .A(n925), .B(n926), .Z(SUM[356]) );
  XNOR U1083 ( .A(B[356]), .B(A[356]), .Z(n926) );
  AND U1084 ( .A(n927), .B(n928), .Z(n925) );
  NAND U1085 ( .A(B[355]), .B(n929), .Z(n928) );
  NANDN U1086 ( .A(A[355]), .B(n930), .Z(n929) );
  NANDN U1087 ( .A(n930), .B(A[355]), .Z(n927) );
  XOR U1088 ( .A(n930), .B(n931), .Z(SUM[355]) );
  XNOR U1089 ( .A(B[355]), .B(A[355]), .Z(n931) );
  AND U1090 ( .A(n932), .B(n933), .Z(n930) );
  NAND U1091 ( .A(B[354]), .B(n934), .Z(n933) );
  NANDN U1092 ( .A(A[354]), .B(n935), .Z(n934) );
  NANDN U1093 ( .A(n935), .B(A[354]), .Z(n932) );
  XOR U1094 ( .A(n935), .B(n936), .Z(SUM[354]) );
  XNOR U1095 ( .A(B[354]), .B(A[354]), .Z(n936) );
  AND U1096 ( .A(n937), .B(n938), .Z(n935) );
  NAND U1097 ( .A(B[353]), .B(n939), .Z(n938) );
  NANDN U1098 ( .A(A[353]), .B(n940), .Z(n939) );
  NANDN U1099 ( .A(n940), .B(A[353]), .Z(n937) );
  XOR U1100 ( .A(n940), .B(n941), .Z(SUM[353]) );
  XNOR U1101 ( .A(B[353]), .B(A[353]), .Z(n941) );
  AND U1102 ( .A(n942), .B(n943), .Z(n940) );
  NAND U1103 ( .A(B[352]), .B(n944), .Z(n943) );
  NANDN U1104 ( .A(A[352]), .B(n945), .Z(n944) );
  NANDN U1105 ( .A(n945), .B(A[352]), .Z(n942) );
  XOR U1106 ( .A(n945), .B(n946), .Z(SUM[352]) );
  XNOR U1107 ( .A(B[352]), .B(A[352]), .Z(n946) );
  AND U1108 ( .A(n947), .B(n948), .Z(n945) );
  NAND U1109 ( .A(B[351]), .B(n949), .Z(n948) );
  NANDN U1110 ( .A(A[351]), .B(n950), .Z(n949) );
  NANDN U1111 ( .A(n950), .B(A[351]), .Z(n947) );
  XOR U1112 ( .A(n950), .B(n951), .Z(SUM[351]) );
  XNOR U1113 ( .A(B[351]), .B(A[351]), .Z(n951) );
  AND U1114 ( .A(n952), .B(n953), .Z(n950) );
  NAND U1115 ( .A(B[350]), .B(n954), .Z(n953) );
  NANDN U1116 ( .A(A[350]), .B(n955), .Z(n954) );
  NANDN U1117 ( .A(n955), .B(A[350]), .Z(n952) );
  XOR U1118 ( .A(n955), .B(n956), .Z(SUM[350]) );
  XNOR U1119 ( .A(B[350]), .B(A[350]), .Z(n956) );
  AND U1120 ( .A(n957), .B(n958), .Z(n955) );
  NAND U1121 ( .A(B[349]), .B(n959), .Z(n958) );
  NANDN U1122 ( .A(A[349]), .B(n960), .Z(n959) );
  NANDN U1123 ( .A(n960), .B(A[349]), .Z(n957) );
  XOR U1124 ( .A(n961), .B(n962), .Z(SUM[34]) );
  XNOR U1125 ( .A(B[34]), .B(A[34]), .Z(n962) );
  XOR U1126 ( .A(n960), .B(n963), .Z(SUM[349]) );
  XNOR U1127 ( .A(B[349]), .B(A[349]), .Z(n963) );
  AND U1128 ( .A(n964), .B(n965), .Z(n960) );
  NAND U1129 ( .A(B[348]), .B(n966), .Z(n965) );
  NANDN U1130 ( .A(A[348]), .B(n967), .Z(n966) );
  NANDN U1131 ( .A(n967), .B(A[348]), .Z(n964) );
  XOR U1132 ( .A(n967), .B(n968), .Z(SUM[348]) );
  XNOR U1133 ( .A(B[348]), .B(A[348]), .Z(n968) );
  AND U1134 ( .A(n969), .B(n970), .Z(n967) );
  NAND U1135 ( .A(B[347]), .B(n971), .Z(n970) );
  NANDN U1136 ( .A(A[347]), .B(n972), .Z(n971) );
  NANDN U1137 ( .A(n972), .B(A[347]), .Z(n969) );
  XOR U1138 ( .A(n972), .B(n973), .Z(SUM[347]) );
  XNOR U1139 ( .A(B[347]), .B(A[347]), .Z(n973) );
  AND U1140 ( .A(n974), .B(n975), .Z(n972) );
  NAND U1141 ( .A(B[346]), .B(n976), .Z(n975) );
  NANDN U1142 ( .A(A[346]), .B(n977), .Z(n976) );
  NANDN U1143 ( .A(n977), .B(A[346]), .Z(n974) );
  XOR U1144 ( .A(n977), .B(n978), .Z(SUM[346]) );
  XNOR U1145 ( .A(B[346]), .B(A[346]), .Z(n978) );
  AND U1146 ( .A(n979), .B(n980), .Z(n977) );
  NAND U1147 ( .A(B[345]), .B(n981), .Z(n980) );
  NANDN U1148 ( .A(A[345]), .B(n982), .Z(n981) );
  NANDN U1149 ( .A(n982), .B(A[345]), .Z(n979) );
  XOR U1150 ( .A(n982), .B(n983), .Z(SUM[345]) );
  XNOR U1151 ( .A(B[345]), .B(A[345]), .Z(n983) );
  AND U1152 ( .A(n984), .B(n985), .Z(n982) );
  NAND U1153 ( .A(B[344]), .B(n986), .Z(n985) );
  NANDN U1154 ( .A(A[344]), .B(n987), .Z(n986) );
  NANDN U1155 ( .A(n987), .B(A[344]), .Z(n984) );
  XOR U1156 ( .A(n987), .B(n988), .Z(SUM[344]) );
  XNOR U1157 ( .A(B[344]), .B(A[344]), .Z(n988) );
  AND U1158 ( .A(n989), .B(n990), .Z(n987) );
  NAND U1159 ( .A(B[343]), .B(n991), .Z(n990) );
  NANDN U1160 ( .A(A[343]), .B(n992), .Z(n991) );
  NANDN U1161 ( .A(n992), .B(A[343]), .Z(n989) );
  XOR U1162 ( .A(n992), .B(n993), .Z(SUM[343]) );
  XNOR U1163 ( .A(B[343]), .B(A[343]), .Z(n993) );
  AND U1164 ( .A(n994), .B(n995), .Z(n992) );
  NAND U1165 ( .A(B[342]), .B(n996), .Z(n995) );
  NANDN U1166 ( .A(A[342]), .B(n997), .Z(n996) );
  NANDN U1167 ( .A(n997), .B(A[342]), .Z(n994) );
  XOR U1168 ( .A(n997), .B(n998), .Z(SUM[342]) );
  XNOR U1169 ( .A(B[342]), .B(A[342]), .Z(n998) );
  AND U1170 ( .A(n999), .B(n1000), .Z(n997) );
  NAND U1171 ( .A(B[341]), .B(n1001), .Z(n1000) );
  NANDN U1172 ( .A(A[341]), .B(n1002), .Z(n1001) );
  NANDN U1173 ( .A(n1002), .B(A[341]), .Z(n999) );
  XOR U1174 ( .A(n1002), .B(n1003), .Z(SUM[341]) );
  XNOR U1175 ( .A(B[341]), .B(A[341]), .Z(n1003) );
  AND U1176 ( .A(n1004), .B(n1005), .Z(n1002) );
  NAND U1177 ( .A(B[340]), .B(n1006), .Z(n1005) );
  NANDN U1178 ( .A(A[340]), .B(n1007), .Z(n1006) );
  NANDN U1179 ( .A(n1007), .B(A[340]), .Z(n1004) );
  XOR U1180 ( .A(n1007), .B(n1008), .Z(SUM[340]) );
  XNOR U1181 ( .A(B[340]), .B(A[340]), .Z(n1008) );
  AND U1182 ( .A(n1009), .B(n1010), .Z(n1007) );
  NAND U1183 ( .A(B[339]), .B(n1011), .Z(n1010) );
  NANDN U1184 ( .A(A[339]), .B(n1012), .Z(n1011) );
  NANDN U1185 ( .A(n1012), .B(A[339]), .Z(n1009) );
  XOR U1186 ( .A(n1013), .B(n1014), .Z(SUM[33]) );
  XNOR U1187 ( .A(B[33]), .B(A[33]), .Z(n1014) );
  XOR U1188 ( .A(n1012), .B(n1015), .Z(SUM[339]) );
  XNOR U1189 ( .A(B[339]), .B(A[339]), .Z(n1015) );
  AND U1190 ( .A(n1016), .B(n1017), .Z(n1012) );
  NAND U1191 ( .A(B[338]), .B(n1018), .Z(n1017) );
  NANDN U1192 ( .A(A[338]), .B(n1019), .Z(n1018) );
  NANDN U1193 ( .A(n1019), .B(A[338]), .Z(n1016) );
  XOR U1194 ( .A(n1019), .B(n1020), .Z(SUM[338]) );
  XNOR U1195 ( .A(B[338]), .B(A[338]), .Z(n1020) );
  AND U1196 ( .A(n1021), .B(n1022), .Z(n1019) );
  NAND U1197 ( .A(B[337]), .B(n1023), .Z(n1022) );
  NANDN U1198 ( .A(A[337]), .B(n1024), .Z(n1023) );
  NANDN U1199 ( .A(n1024), .B(A[337]), .Z(n1021) );
  XOR U1200 ( .A(n1024), .B(n1025), .Z(SUM[337]) );
  XNOR U1201 ( .A(B[337]), .B(A[337]), .Z(n1025) );
  AND U1202 ( .A(n1026), .B(n1027), .Z(n1024) );
  NAND U1203 ( .A(B[336]), .B(n1028), .Z(n1027) );
  NANDN U1204 ( .A(A[336]), .B(n1029), .Z(n1028) );
  NANDN U1205 ( .A(n1029), .B(A[336]), .Z(n1026) );
  XOR U1206 ( .A(n1029), .B(n1030), .Z(SUM[336]) );
  XNOR U1207 ( .A(B[336]), .B(A[336]), .Z(n1030) );
  AND U1208 ( .A(n1031), .B(n1032), .Z(n1029) );
  NAND U1209 ( .A(B[335]), .B(n1033), .Z(n1032) );
  NANDN U1210 ( .A(A[335]), .B(n1034), .Z(n1033) );
  NANDN U1211 ( .A(n1034), .B(A[335]), .Z(n1031) );
  XOR U1212 ( .A(n1034), .B(n1035), .Z(SUM[335]) );
  XNOR U1213 ( .A(B[335]), .B(A[335]), .Z(n1035) );
  AND U1214 ( .A(n1036), .B(n1037), .Z(n1034) );
  NAND U1215 ( .A(B[334]), .B(n1038), .Z(n1037) );
  NANDN U1216 ( .A(A[334]), .B(n1039), .Z(n1038) );
  NANDN U1217 ( .A(n1039), .B(A[334]), .Z(n1036) );
  XOR U1218 ( .A(n1039), .B(n1040), .Z(SUM[334]) );
  XNOR U1219 ( .A(B[334]), .B(A[334]), .Z(n1040) );
  AND U1220 ( .A(n1041), .B(n1042), .Z(n1039) );
  NAND U1221 ( .A(B[333]), .B(n1043), .Z(n1042) );
  NANDN U1222 ( .A(A[333]), .B(n1044), .Z(n1043) );
  NANDN U1223 ( .A(n1044), .B(A[333]), .Z(n1041) );
  XOR U1224 ( .A(n1044), .B(n1045), .Z(SUM[333]) );
  XNOR U1225 ( .A(B[333]), .B(A[333]), .Z(n1045) );
  AND U1226 ( .A(n1046), .B(n1047), .Z(n1044) );
  NAND U1227 ( .A(B[332]), .B(n1048), .Z(n1047) );
  NANDN U1228 ( .A(A[332]), .B(n1049), .Z(n1048) );
  NANDN U1229 ( .A(n1049), .B(A[332]), .Z(n1046) );
  XOR U1230 ( .A(n1049), .B(n1050), .Z(SUM[332]) );
  XNOR U1231 ( .A(B[332]), .B(A[332]), .Z(n1050) );
  AND U1232 ( .A(n1051), .B(n1052), .Z(n1049) );
  NAND U1233 ( .A(B[331]), .B(n1053), .Z(n1052) );
  NANDN U1234 ( .A(A[331]), .B(n1054), .Z(n1053) );
  NANDN U1235 ( .A(n1054), .B(A[331]), .Z(n1051) );
  XOR U1236 ( .A(n1054), .B(n1055), .Z(SUM[331]) );
  XNOR U1237 ( .A(B[331]), .B(A[331]), .Z(n1055) );
  AND U1238 ( .A(n1056), .B(n1057), .Z(n1054) );
  NAND U1239 ( .A(B[330]), .B(n1058), .Z(n1057) );
  NANDN U1240 ( .A(A[330]), .B(n1059), .Z(n1058) );
  NANDN U1241 ( .A(n1059), .B(A[330]), .Z(n1056) );
  XOR U1242 ( .A(n1059), .B(n1060), .Z(SUM[330]) );
  XNOR U1243 ( .A(B[330]), .B(A[330]), .Z(n1060) );
  AND U1244 ( .A(n1061), .B(n1062), .Z(n1059) );
  NAND U1245 ( .A(B[329]), .B(n1063), .Z(n1062) );
  NANDN U1246 ( .A(A[329]), .B(n1064), .Z(n1063) );
  NANDN U1247 ( .A(n1064), .B(A[329]), .Z(n1061) );
  XOR U1248 ( .A(n1065), .B(n1066), .Z(SUM[32]) );
  XNOR U1249 ( .A(B[32]), .B(A[32]), .Z(n1066) );
  XOR U1250 ( .A(n1064), .B(n1067), .Z(SUM[329]) );
  XNOR U1251 ( .A(B[329]), .B(A[329]), .Z(n1067) );
  AND U1252 ( .A(n1068), .B(n1069), .Z(n1064) );
  NAND U1253 ( .A(B[328]), .B(n1070), .Z(n1069) );
  NANDN U1254 ( .A(A[328]), .B(n1071), .Z(n1070) );
  NANDN U1255 ( .A(n1071), .B(A[328]), .Z(n1068) );
  XOR U1256 ( .A(n1071), .B(n1072), .Z(SUM[328]) );
  XNOR U1257 ( .A(B[328]), .B(A[328]), .Z(n1072) );
  AND U1258 ( .A(n1073), .B(n1074), .Z(n1071) );
  NAND U1259 ( .A(B[327]), .B(n1075), .Z(n1074) );
  NANDN U1260 ( .A(A[327]), .B(n1076), .Z(n1075) );
  NANDN U1261 ( .A(n1076), .B(A[327]), .Z(n1073) );
  XOR U1262 ( .A(n1076), .B(n1077), .Z(SUM[327]) );
  XNOR U1263 ( .A(B[327]), .B(A[327]), .Z(n1077) );
  AND U1264 ( .A(n1078), .B(n1079), .Z(n1076) );
  NAND U1265 ( .A(B[326]), .B(n1080), .Z(n1079) );
  NANDN U1266 ( .A(A[326]), .B(n1081), .Z(n1080) );
  NANDN U1267 ( .A(n1081), .B(A[326]), .Z(n1078) );
  XOR U1268 ( .A(n1081), .B(n1082), .Z(SUM[326]) );
  XNOR U1269 ( .A(B[326]), .B(A[326]), .Z(n1082) );
  AND U1270 ( .A(n1083), .B(n1084), .Z(n1081) );
  NAND U1271 ( .A(B[325]), .B(n1085), .Z(n1084) );
  NANDN U1272 ( .A(A[325]), .B(n1086), .Z(n1085) );
  NANDN U1273 ( .A(n1086), .B(A[325]), .Z(n1083) );
  XOR U1274 ( .A(n1086), .B(n1087), .Z(SUM[325]) );
  XNOR U1275 ( .A(B[325]), .B(A[325]), .Z(n1087) );
  AND U1276 ( .A(n1088), .B(n1089), .Z(n1086) );
  NAND U1277 ( .A(B[324]), .B(n1090), .Z(n1089) );
  NANDN U1278 ( .A(A[324]), .B(n1091), .Z(n1090) );
  NANDN U1279 ( .A(n1091), .B(A[324]), .Z(n1088) );
  XOR U1280 ( .A(n1091), .B(n1092), .Z(SUM[324]) );
  XNOR U1281 ( .A(B[324]), .B(A[324]), .Z(n1092) );
  AND U1282 ( .A(n1093), .B(n1094), .Z(n1091) );
  NAND U1283 ( .A(B[323]), .B(n1095), .Z(n1094) );
  NANDN U1284 ( .A(A[323]), .B(n1096), .Z(n1095) );
  NANDN U1285 ( .A(n1096), .B(A[323]), .Z(n1093) );
  XOR U1286 ( .A(n1096), .B(n1097), .Z(SUM[323]) );
  XNOR U1287 ( .A(B[323]), .B(A[323]), .Z(n1097) );
  AND U1288 ( .A(n1098), .B(n1099), .Z(n1096) );
  NAND U1289 ( .A(B[322]), .B(n1100), .Z(n1099) );
  NANDN U1290 ( .A(A[322]), .B(n1101), .Z(n1100) );
  NANDN U1291 ( .A(n1101), .B(A[322]), .Z(n1098) );
  XOR U1292 ( .A(n1101), .B(n1102), .Z(SUM[322]) );
  XNOR U1293 ( .A(B[322]), .B(A[322]), .Z(n1102) );
  AND U1294 ( .A(n1103), .B(n1104), .Z(n1101) );
  NAND U1295 ( .A(B[321]), .B(n1105), .Z(n1104) );
  NANDN U1296 ( .A(A[321]), .B(n1106), .Z(n1105) );
  NANDN U1297 ( .A(n1106), .B(A[321]), .Z(n1103) );
  XOR U1298 ( .A(n1106), .B(n1107), .Z(SUM[321]) );
  XNOR U1299 ( .A(B[321]), .B(A[321]), .Z(n1107) );
  AND U1300 ( .A(n1108), .B(n1109), .Z(n1106) );
  NAND U1301 ( .A(B[320]), .B(n1110), .Z(n1109) );
  NANDN U1302 ( .A(A[320]), .B(n1111), .Z(n1110) );
  NANDN U1303 ( .A(n1111), .B(A[320]), .Z(n1108) );
  XOR U1304 ( .A(n1111), .B(n1112), .Z(SUM[320]) );
  XNOR U1305 ( .A(B[320]), .B(A[320]), .Z(n1112) );
  AND U1306 ( .A(n1113), .B(n1114), .Z(n1111) );
  NAND U1307 ( .A(B[319]), .B(n1115), .Z(n1114) );
  NANDN U1308 ( .A(A[319]), .B(n1116), .Z(n1115) );
  NANDN U1309 ( .A(n1116), .B(A[319]), .Z(n1113) );
  XOR U1310 ( .A(n1117), .B(n1118), .Z(SUM[31]) );
  XNOR U1311 ( .A(B[31]), .B(A[31]), .Z(n1118) );
  XOR U1312 ( .A(n1116), .B(n1119), .Z(SUM[319]) );
  XNOR U1313 ( .A(B[319]), .B(A[319]), .Z(n1119) );
  AND U1314 ( .A(n1120), .B(n1121), .Z(n1116) );
  NAND U1315 ( .A(B[318]), .B(n1122), .Z(n1121) );
  NANDN U1316 ( .A(A[318]), .B(n1123), .Z(n1122) );
  NANDN U1317 ( .A(n1123), .B(A[318]), .Z(n1120) );
  XOR U1318 ( .A(n1123), .B(n1124), .Z(SUM[318]) );
  XNOR U1319 ( .A(B[318]), .B(A[318]), .Z(n1124) );
  AND U1320 ( .A(n1125), .B(n1126), .Z(n1123) );
  NAND U1321 ( .A(B[317]), .B(n1127), .Z(n1126) );
  NANDN U1322 ( .A(A[317]), .B(n1128), .Z(n1127) );
  NANDN U1323 ( .A(n1128), .B(A[317]), .Z(n1125) );
  XOR U1324 ( .A(n1128), .B(n1129), .Z(SUM[317]) );
  XNOR U1325 ( .A(B[317]), .B(A[317]), .Z(n1129) );
  AND U1326 ( .A(n1130), .B(n1131), .Z(n1128) );
  NAND U1327 ( .A(B[316]), .B(n1132), .Z(n1131) );
  NANDN U1328 ( .A(A[316]), .B(n1133), .Z(n1132) );
  NANDN U1329 ( .A(n1133), .B(A[316]), .Z(n1130) );
  XOR U1330 ( .A(n1133), .B(n1134), .Z(SUM[316]) );
  XNOR U1331 ( .A(B[316]), .B(A[316]), .Z(n1134) );
  AND U1332 ( .A(n1135), .B(n1136), .Z(n1133) );
  NAND U1333 ( .A(B[315]), .B(n1137), .Z(n1136) );
  NANDN U1334 ( .A(A[315]), .B(n1138), .Z(n1137) );
  NANDN U1335 ( .A(n1138), .B(A[315]), .Z(n1135) );
  XOR U1336 ( .A(n1138), .B(n1139), .Z(SUM[315]) );
  XNOR U1337 ( .A(B[315]), .B(A[315]), .Z(n1139) );
  AND U1338 ( .A(n1140), .B(n1141), .Z(n1138) );
  NAND U1339 ( .A(B[314]), .B(n1142), .Z(n1141) );
  NANDN U1340 ( .A(A[314]), .B(n1143), .Z(n1142) );
  NANDN U1341 ( .A(n1143), .B(A[314]), .Z(n1140) );
  XOR U1342 ( .A(n1143), .B(n1144), .Z(SUM[314]) );
  XNOR U1343 ( .A(B[314]), .B(A[314]), .Z(n1144) );
  AND U1344 ( .A(n1145), .B(n1146), .Z(n1143) );
  NAND U1345 ( .A(B[313]), .B(n1147), .Z(n1146) );
  NANDN U1346 ( .A(A[313]), .B(n1148), .Z(n1147) );
  NANDN U1347 ( .A(n1148), .B(A[313]), .Z(n1145) );
  XOR U1348 ( .A(n1148), .B(n1149), .Z(SUM[313]) );
  XNOR U1349 ( .A(B[313]), .B(A[313]), .Z(n1149) );
  AND U1350 ( .A(n1150), .B(n1151), .Z(n1148) );
  NAND U1351 ( .A(B[312]), .B(n1152), .Z(n1151) );
  NANDN U1352 ( .A(A[312]), .B(n1153), .Z(n1152) );
  NANDN U1353 ( .A(n1153), .B(A[312]), .Z(n1150) );
  XOR U1354 ( .A(n1153), .B(n1154), .Z(SUM[312]) );
  XNOR U1355 ( .A(B[312]), .B(A[312]), .Z(n1154) );
  AND U1356 ( .A(n1155), .B(n1156), .Z(n1153) );
  NAND U1357 ( .A(B[311]), .B(n1157), .Z(n1156) );
  NANDN U1358 ( .A(A[311]), .B(n1158), .Z(n1157) );
  NANDN U1359 ( .A(n1158), .B(A[311]), .Z(n1155) );
  XOR U1360 ( .A(n1158), .B(n1159), .Z(SUM[311]) );
  XNOR U1361 ( .A(B[311]), .B(A[311]), .Z(n1159) );
  AND U1362 ( .A(n1160), .B(n1161), .Z(n1158) );
  NAND U1363 ( .A(B[310]), .B(n1162), .Z(n1161) );
  NANDN U1364 ( .A(A[310]), .B(n1163), .Z(n1162) );
  NANDN U1365 ( .A(n1163), .B(A[310]), .Z(n1160) );
  XOR U1366 ( .A(n1163), .B(n1164), .Z(SUM[310]) );
  XNOR U1367 ( .A(B[310]), .B(A[310]), .Z(n1164) );
  AND U1368 ( .A(n1165), .B(n1166), .Z(n1163) );
  NAND U1369 ( .A(B[309]), .B(n1167), .Z(n1166) );
  NANDN U1370 ( .A(A[309]), .B(n1168), .Z(n1167) );
  NANDN U1371 ( .A(n1168), .B(A[309]), .Z(n1165) );
  XOR U1372 ( .A(n1169), .B(n1170), .Z(SUM[30]) );
  XNOR U1373 ( .A(B[30]), .B(A[30]), .Z(n1170) );
  XOR U1374 ( .A(n1168), .B(n1171), .Z(SUM[309]) );
  XNOR U1375 ( .A(B[309]), .B(A[309]), .Z(n1171) );
  AND U1376 ( .A(n1172), .B(n1173), .Z(n1168) );
  NAND U1377 ( .A(B[308]), .B(n1174), .Z(n1173) );
  NANDN U1378 ( .A(A[308]), .B(n1175), .Z(n1174) );
  NANDN U1379 ( .A(n1175), .B(A[308]), .Z(n1172) );
  XOR U1380 ( .A(n1175), .B(n1176), .Z(SUM[308]) );
  XNOR U1381 ( .A(B[308]), .B(A[308]), .Z(n1176) );
  AND U1382 ( .A(n1177), .B(n1178), .Z(n1175) );
  NAND U1383 ( .A(B[307]), .B(n1179), .Z(n1178) );
  NANDN U1384 ( .A(A[307]), .B(n1180), .Z(n1179) );
  NANDN U1385 ( .A(n1180), .B(A[307]), .Z(n1177) );
  XOR U1386 ( .A(n1180), .B(n1181), .Z(SUM[307]) );
  XNOR U1387 ( .A(B[307]), .B(A[307]), .Z(n1181) );
  AND U1388 ( .A(n1182), .B(n1183), .Z(n1180) );
  NAND U1389 ( .A(B[306]), .B(n1184), .Z(n1183) );
  NANDN U1390 ( .A(A[306]), .B(n1185), .Z(n1184) );
  NANDN U1391 ( .A(n1185), .B(A[306]), .Z(n1182) );
  XOR U1392 ( .A(n1185), .B(n1186), .Z(SUM[306]) );
  XNOR U1393 ( .A(B[306]), .B(A[306]), .Z(n1186) );
  AND U1394 ( .A(n1187), .B(n1188), .Z(n1185) );
  NAND U1395 ( .A(B[305]), .B(n1189), .Z(n1188) );
  NANDN U1396 ( .A(A[305]), .B(n1190), .Z(n1189) );
  NANDN U1397 ( .A(n1190), .B(A[305]), .Z(n1187) );
  XOR U1398 ( .A(n1190), .B(n1191), .Z(SUM[305]) );
  XNOR U1399 ( .A(B[305]), .B(A[305]), .Z(n1191) );
  AND U1400 ( .A(n1192), .B(n1193), .Z(n1190) );
  NAND U1401 ( .A(B[304]), .B(n1194), .Z(n1193) );
  NANDN U1402 ( .A(A[304]), .B(n1195), .Z(n1194) );
  NANDN U1403 ( .A(n1195), .B(A[304]), .Z(n1192) );
  XOR U1404 ( .A(n1195), .B(n1196), .Z(SUM[304]) );
  XNOR U1405 ( .A(B[304]), .B(A[304]), .Z(n1196) );
  AND U1406 ( .A(n1197), .B(n1198), .Z(n1195) );
  NAND U1407 ( .A(B[303]), .B(n1199), .Z(n1198) );
  NANDN U1408 ( .A(A[303]), .B(n1200), .Z(n1199) );
  NANDN U1409 ( .A(n1200), .B(A[303]), .Z(n1197) );
  XOR U1410 ( .A(n1200), .B(n1201), .Z(SUM[303]) );
  XNOR U1411 ( .A(B[303]), .B(A[303]), .Z(n1201) );
  AND U1412 ( .A(n1202), .B(n1203), .Z(n1200) );
  NAND U1413 ( .A(B[302]), .B(n1204), .Z(n1203) );
  NANDN U1414 ( .A(A[302]), .B(n1205), .Z(n1204) );
  NANDN U1415 ( .A(n1205), .B(A[302]), .Z(n1202) );
  XOR U1416 ( .A(n1205), .B(n1206), .Z(SUM[302]) );
  XNOR U1417 ( .A(B[302]), .B(A[302]), .Z(n1206) );
  AND U1418 ( .A(n1207), .B(n1208), .Z(n1205) );
  NAND U1419 ( .A(B[301]), .B(n1209), .Z(n1208) );
  NANDN U1420 ( .A(A[301]), .B(n1210), .Z(n1209) );
  NANDN U1421 ( .A(n1210), .B(A[301]), .Z(n1207) );
  XOR U1422 ( .A(n1210), .B(n1211), .Z(SUM[301]) );
  XNOR U1423 ( .A(B[301]), .B(A[301]), .Z(n1211) );
  AND U1424 ( .A(n1212), .B(n1213), .Z(n1210) );
  NAND U1425 ( .A(B[300]), .B(n1214), .Z(n1213) );
  NANDN U1426 ( .A(A[300]), .B(n1215), .Z(n1214) );
  NANDN U1427 ( .A(n1215), .B(A[300]), .Z(n1212) );
  XOR U1428 ( .A(n1215), .B(n1216), .Z(SUM[300]) );
  XNOR U1429 ( .A(B[300]), .B(A[300]), .Z(n1216) );
  AND U1430 ( .A(n1217), .B(n1218), .Z(n1215) );
  NAND U1431 ( .A(B[299]), .B(n1219), .Z(n1218) );
  NANDN U1432 ( .A(A[299]), .B(n1220), .Z(n1219) );
  NANDN U1433 ( .A(n1220), .B(A[299]), .Z(n1217) );
  XOR U1434 ( .A(n1221), .B(n1222), .Z(SUM[2]) );
  XOR U1435 ( .A(B[2]), .B(A[2]), .Z(n1222) );
  XOR U1436 ( .A(n1223), .B(n1224), .Z(SUM[29]) );
  XNOR U1437 ( .A(B[29]), .B(A[29]), .Z(n1224) );
  XOR U1438 ( .A(n1220), .B(n1225), .Z(SUM[299]) );
  XNOR U1439 ( .A(B[299]), .B(A[299]), .Z(n1225) );
  AND U1440 ( .A(n1226), .B(n1227), .Z(n1220) );
  NAND U1441 ( .A(B[298]), .B(n1228), .Z(n1227) );
  NANDN U1442 ( .A(A[298]), .B(n1229), .Z(n1228) );
  NANDN U1443 ( .A(n1229), .B(A[298]), .Z(n1226) );
  XOR U1444 ( .A(n1229), .B(n1230), .Z(SUM[298]) );
  XNOR U1445 ( .A(B[298]), .B(A[298]), .Z(n1230) );
  AND U1446 ( .A(n1231), .B(n1232), .Z(n1229) );
  NAND U1447 ( .A(B[297]), .B(n1233), .Z(n1232) );
  NANDN U1448 ( .A(A[297]), .B(n1234), .Z(n1233) );
  NANDN U1449 ( .A(n1234), .B(A[297]), .Z(n1231) );
  XOR U1450 ( .A(n1234), .B(n1235), .Z(SUM[297]) );
  XNOR U1451 ( .A(B[297]), .B(A[297]), .Z(n1235) );
  AND U1452 ( .A(n1236), .B(n1237), .Z(n1234) );
  NAND U1453 ( .A(B[296]), .B(n1238), .Z(n1237) );
  NANDN U1454 ( .A(A[296]), .B(n1239), .Z(n1238) );
  NANDN U1455 ( .A(n1239), .B(A[296]), .Z(n1236) );
  XOR U1456 ( .A(n1239), .B(n1240), .Z(SUM[296]) );
  XNOR U1457 ( .A(B[296]), .B(A[296]), .Z(n1240) );
  AND U1458 ( .A(n1241), .B(n1242), .Z(n1239) );
  NAND U1459 ( .A(B[295]), .B(n1243), .Z(n1242) );
  NANDN U1460 ( .A(A[295]), .B(n1244), .Z(n1243) );
  NANDN U1461 ( .A(n1244), .B(A[295]), .Z(n1241) );
  XOR U1462 ( .A(n1244), .B(n1245), .Z(SUM[295]) );
  XNOR U1463 ( .A(B[295]), .B(A[295]), .Z(n1245) );
  AND U1464 ( .A(n1246), .B(n1247), .Z(n1244) );
  NAND U1465 ( .A(B[294]), .B(n1248), .Z(n1247) );
  NANDN U1466 ( .A(A[294]), .B(n1249), .Z(n1248) );
  NANDN U1467 ( .A(n1249), .B(A[294]), .Z(n1246) );
  XOR U1468 ( .A(n1249), .B(n1250), .Z(SUM[294]) );
  XNOR U1469 ( .A(B[294]), .B(A[294]), .Z(n1250) );
  AND U1470 ( .A(n1251), .B(n1252), .Z(n1249) );
  NAND U1471 ( .A(B[293]), .B(n1253), .Z(n1252) );
  NANDN U1472 ( .A(A[293]), .B(n1254), .Z(n1253) );
  NANDN U1473 ( .A(n1254), .B(A[293]), .Z(n1251) );
  XOR U1474 ( .A(n1254), .B(n1255), .Z(SUM[293]) );
  XNOR U1475 ( .A(B[293]), .B(A[293]), .Z(n1255) );
  AND U1476 ( .A(n1256), .B(n1257), .Z(n1254) );
  NAND U1477 ( .A(B[292]), .B(n1258), .Z(n1257) );
  NANDN U1478 ( .A(A[292]), .B(n1259), .Z(n1258) );
  NANDN U1479 ( .A(n1259), .B(A[292]), .Z(n1256) );
  XOR U1480 ( .A(n1259), .B(n1260), .Z(SUM[292]) );
  XNOR U1481 ( .A(B[292]), .B(A[292]), .Z(n1260) );
  AND U1482 ( .A(n1261), .B(n1262), .Z(n1259) );
  NAND U1483 ( .A(B[291]), .B(n1263), .Z(n1262) );
  NANDN U1484 ( .A(A[291]), .B(n1264), .Z(n1263) );
  NANDN U1485 ( .A(n1264), .B(A[291]), .Z(n1261) );
  XOR U1486 ( .A(n1264), .B(n1265), .Z(SUM[291]) );
  XNOR U1487 ( .A(B[291]), .B(A[291]), .Z(n1265) );
  AND U1488 ( .A(n1266), .B(n1267), .Z(n1264) );
  NAND U1489 ( .A(B[290]), .B(n1268), .Z(n1267) );
  NANDN U1490 ( .A(A[290]), .B(n1269), .Z(n1268) );
  NANDN U1491 ( .A(n1269), .B(A[290]), .Z(n1266) );
  XOR U1492 ( .A(n1269), .B(n1270), .Z(SUM[290]) );
  XNOR U1493 ( .A(B[290]), .B(A[290]), .Z(n1270) );
  AND U1494 ( .A(n1271), .B(n1272), .Z(n1269) );
  NAND U1495 ( .A(B[289]), .B(n1273), .Z(n1272) );
  NANDN U1496 ( .A(A[289]), .B(n1274), .Z(n1273) );
  NANDN U1497 ( .A(n1274), .B(A[289]), .Z(n1271) );
  XOR U1498 ( .A(n1275), .B(n1276), .Z(SUM[28]) );
  XNOR U1499 ( .A(B[28]), .B(A[28]), .Z(n1276) );
  XOR U1500 ( .A(n1274), .B(n1277), .Z(SUM[289]) );
  XNOR U1501 ( .A(B[289]), .B(A[289]), .Z(n1277) );
  AND U1502 ( .A(n1278), .B(n1279), .Z(n1274) );
  NAND U1503 ( .A(B[288]), .B(n1280), .Z(n1279) );
  NANDN U1504 ( .A(A[288]), .B(n1281), .Z(n1280) );
  NANDN U1505 ( .A(n1281), .B(A[288]), .Z(n1278) );
  XOR U1506 ( .A(n1281), .B(n1282), .Z(SUM[288]) );
  XNOR U1507 ( .A(B[288]), .B(A[288]), .Z(n1282) );
  AND U1508 ( .A(n1283), .B(n1284), .Z(n1281) );
  NAND U1509 ( .A(B[287]), .B(n1285), .Z(n1284) );
  NANDN U1510 ( .A(A[287]), .B(n1286), .Z(n1285) );
  NANDN U1511 ( .A(n1286), .B(A[287]), .Z(n1283) );
  XOR U1512 ( .A(n1286), .B(n1287), .Z(SUM[287]) );
  XNOR U1513 ( .A(B[287]), .B(A[287]), .Z(n1287) );
  AND U1514 ( .A(n1288), .B(n1289), .Z(n1286) );
  NAND U1515 ( .A(B[286]), .B(n1290), .Z(n1289) );
  NANDN U1516 ( .A(A[286]), .B(n1291), .Z(n1290) );
  NANDN U1517 ( .A(n1291), .B(A[286]), .Z(n1288) );
  XOR U1518 ( .A(n1291), .B(n1292), .Z(SUM[286]) );
  XNOR U1519 ( .A(B[286]), .B(A[286]), .Z(n1292) );
  AND U1520 ( .A(n1293), .B(n1294), .Z(n1291) );
  NAND U1521 ( .A(B[285]), .B(n1295), .Z(n1294) );
  NANDN U1522 ( .A(A[285]), .B(n1296), .Z(n1295) );
  NANDN U1523 ( .A(n1296), .B(A[285]), .Z(n1293) );
  XOR U1524 ( .A(n1296), .B(n1297), .Z(SUM[285]) );
  XNOR U1525 ( .A(B[285]), .B(A[285]), .Z(n1297) );
  AND U1526 ( .A(n1298), .B(n1299), .Z(n1296) );
  NAND U1527 ( .A(B[284]), .B(n1300), .Z(n1299) );
  NANDN U1528 ( .A(A[284]), .B(n1301), .Z(n1300) );
  NANDN U1529 ( .A(n1301), .B(A[284]), .Z(n1298) );
  XOR U1530 ( .A(n1301), .B(n1302), .Z(SUM[284]) );
  XNOR U1531 ( .A(B[284]), .B(A[284]), .Z(n1302) );
  AND U1532 ( .A(n1303), .B(n1304), .Z(n1301) );
  NAND U1533 ( .A(B[283]), .B(n1305), .Z(n1304) );
  NANDN U1534 ( .A(A[283]), .B(n1306), .Z(n1305) );
  NANDN U1535 ( .A(n1306), .B(A[283]), .Z(n1303) );
  XOR U1536 ( .A(n1306), .B(n1307), .Z(SUM[283]) );
  XNOR U1537 ( .A(B[283]), .B(A[283]), .Z(n1307) );
  AND U1538 ( .A(n1308), .B(n1309), .Z(n1306) );
  NAND U1539 ( .A(B[282]), .B(n1310), .Z(n1309) );
  NANDN U1540 ( .A(A[282]), .B(n1311), .Z(n1310) );
  NANDN U1541 ( .A(n1311), .B(A[282]), .Z(n1308) );
  XOR U1542 ( .A(n1311), .B(n1312), .Z(SUM[282]) );
  XNOR U1543 ( .A(B[282]), .B(A[282]), .Z(n1312) );
  AND U1544 ( .A(n1313), .B(n1314), .Z(n1311) );
  NAND U1545 ( .A(B[281]), .B(n1315), .Z(n1314) );
  NANDN U1546 ( .A(A[281]), .B(n1316), .Z(n1315) );
  NANDN U1547 ( .A(n1316), .B(A[281]), .Z(n1313) );
  XOR U1548 ( .A(n1316), .B(n1317), .Z(SUM[281]) );
  XNOR U1549 ( .A(B[281]), .B(A[281]), .Z(n1317) );
  AND U1550 ( .A(n1318), .B(n1319), .Z(n1316) );
  NAND U1551 ( .A(B[280]), .B(n1320), .Z(n1319) );
  NANDN U1552 ( .A(A[280]), .B(n1321), .Z(n1320) );
  NANDN U1553 ( .A(n1321), .B(A[280]), .Z(n1318) );
  XOR U1554 ( .A(n1321), .B(n1322), .Z(SUM[280]) );
  XNOR U1555 ( .A(B[280]), .B(A[280]), .Z(n1322) );
  AND U1556 ( .A(n1323), .B(n1324), .Z(n1321) );
  NAND U1557 ( .A(B[279]), .B(n1325), .Z(n1324) );
  NANDN U1558 ( .A(A[279]), .B(n1326), .Z(n1325) );
  NANDN U1559 ( .A(n1326), .B(A[279]), .Z(n1323) );
  XOR U1560 ( .A(n1327), .B(n1328), .Z(SUM[27]) );
  XNOR U1561 ( .A(B[27]), .B(A[27]), .Z(n1328) );
  XOR U1562 ( .A(n1326), .B(n1329), .Z(SUM[279]) );
  XNOR U1563 ( .A(B[279]), .B(A[279]), .Z(n1329) );
  AND U1564 ( .A(n1330), .B(n1331), .Z(n1326) );
  NAND U1565 ( .A(B[278]), .B(n1332), .Z(n1331) );
  NANDN U1566 ( .A(A[278]), .B(n1333), .Z(n1332) );
  NANDN U1567 ( .A(n1333), .B(A[278]), .Z(n1330) );
  XOR U1568 ( .A(n1333), .B(n1334), .Z(SUM[278]) );
  XNOR U1569 ( .A(B[278]), .B(A[278]), .Z(n1334) );
  AND U1570 ( .A(n1335), .B(n1336), .Z(n1333) );
  NAND U1571 ( .A(B[277]), .B(n1337), .Z(n1336) );
  NANDN U1572 ( .A(A[277]), .B(n1338), .Z(n1337) );
  NANDN U1573 ( .A(n1338), .B(A[277]), .Z(n1335) );
  XOR U1574 ( .A(n1338), .B(n1339), .Z(SUM[277]) );
  XNOR U1575 ( .A(B[277]), .B(A[277]), .Z(n1339) );
  AND U1576 ( .A(n1340), .B(n1341), .Z(n1338) );
  NAND U1577 ( .A(B[276]), .B(n1342), .Z(n1341) );
  NANDN U1578 ( .A(A[276]), .B(n1343), .Z(n1342) );
  NANDN U1579 ( .A(n1343), .B(A[276]), .Z(n1340) );
  XOR U1580 ( .A(n1343), .B(n1344), .Z(SUM[276]) );
  XNOR U1581 ( .A(B[276]), .B(A[276]), .Z(n1344) );
  AND U1582 ( .A(n1345), .B(n1346), .Z(n1343) );
  NAND U1583 ( .A(B[275]), .B(n1347), .Z(n1346) );
  NANDN U1584 ( .A(A[275]), .B(n1348), .Z(n1347) );
  NANDN U1585 ( .A(n1348), .B(A[275]), .Z(n1345) );
  XOR U1586 ( .A(n1348), .B(n1349), .Z(SUM[275]) );
  XNOR U1587 ( .A(B[275]), .B(A[275]), .Z(n1349) );
  AND U1588 ( .A(n1350), .B(n1351), .Z(n1348) );
  NAND U1589 ( .A(B[274]), .B(n1352), .Z(n1351) );
  NANDN U1590 ( .A(A[274]), .B(n1353), .Z(n1352) );
  NANDN U1591 ( .A(n1353), .B(A[274]), .Z(n1350) );
  XOR U1592 ( .A(n1353), .B(n1354), .Z(SUM[274]) );
  XNOR U1593 ( .A(B[274]), .B(A[274]), .Z(n1354) );
  AND U1594 ( .A(n1355), .B(n1356), .Z(n1353) );
  NAND U1595 ( .A(B[273]), .B(n1357), .Z(n1356) );
  NANDN U1596 ( .A(A[273]), .B(n1358), .Z(n1357) );
  NANDN U1597 ( .A(n1358), .B(A[273]), .Z(n1355) );
  XOR U1598 ( .A(n1358), .B(n1359), .Z(SUM[273]) );
  XNOR U1599 ( .A(B[273]), .B(A[273]), .Z(n1359) );
  AND U1600 ( .A(n1360), .B(n1361), .Z(n1358) );
  NAND U1601 ( .A(B[272]), .B(n1362), .Z(n1361) );
  NANDN U1602 ( .A(A[272]), .B(n1363), .Z(n1362) );
  NANDN U1603 ( .A(n1363), .B(A[272]), .Z(n1360) );
  XOR U1604 ( .A(n1363), .B(n1364), .Z(SUM[272]) );
  XNOR U1605 ( .A(B[272]), .B(A[272]), .Z(n1364) );
  AND U1606 ( .A(n1365), .B(n1366), .Z(n1363) );
  NAND U1607 ( .A(B[271]), .B(n1367), .Z(n1366) );
  NANDN U1608 ( .A(A[271]), .B(n1368), .Z(n1367) );
  NANDN U1609 ( .A(n1368), .B(A[271]), .Z(n1365) );
  XOR U1610 ( .A(n1368), .B(n1369), .Z(SUM[271]) );
  XNOR U1611 ( .A(B[271]), .B(A[271]), .Z(n1369) );
  AND U1612 ( .A(n1370), .B(n1371), .Z(n1368) );
  NAND U1613 ( .A(B[270]), .B(n1372), .Z(n1371) );
  NANDN U1614 ( .A(A[270]), .B(n1373), .Z(n1372) );
  NANDN U1615 ( .A(n1373), .B(A[270]), .Z(n1370) );
  XOR U1616 ( .A(n1373), .B(n1374), .Z(SUM[270]) );
  XNOR U1617 ( .A(B[270]), .B(A[270]), .Z(n1374) );
  AND U1618 ( .A(n1375), .B(n1376), .Z(n1373) );
  NAND U1619 ( .A(B[269]), .B(n1377), .Z(n1376) );
  NANDN U1620 ( .A(A[269]), .B(n1378), .Z(n1377) );
  NANDN U1621 ( .A(n1378), .B(A[269]), .Z(n1375) );
  XOR U1622 ( .A(n1379), .B(n1380), .Z(SUM[26]) );
  XNOR U1623 ( .A(B[26]), .B(A[26]), .Z(n1380) );
  XOR U1624 ( .A(n1378), .B(n1381), .Z(SUM[269]) );
  XNOR U1625 ( .A(B[269]), .B(A[269]), .Z(n1381) );
  AND U1626 ( .A(n1382), .B(n1383), .Z(n1378) );
  NAND U1627 ( .A(B[268]), .B(n1384), .Z(n1383) );
  NANDN U1628 ( .A(A[268]), .B(n1385), .Z(n1384) );
  NANDN U1629 ( .A(n1385), .B(A[268]), .Z(n1382) );
  XOR U1630 ( .A(n1385), .B(n1386), .Z(SUM[268]) );
  XNOR U1631 ( .A(B[268]), .B(A[268]), .Z(n1386) );
  AND U1632 ( .A(n1387), .B(n1388), .Z(n1385) );
  NAND U1633 ( .A(B[267]), .B(n1389), .Z(n1388) );
  NANDN U1634 ( .A(A[267]), .B(n1390), .Z(n1389) );
  NANDN U1635 ( .A(n1390), .B(A[267]), .Z(n1387) );
  XOR U1636 ( .A(n1390), .B(n1391), .Z(SUM[267]) );
  XNOR U1637 ( .A(B[267]), .B(A[267]), .Z(n1391) );
  AND U1638 ( .A(n1392), .B(n1393), .Z(n1390) );
  NAND U1639 ( .A(B[266]), .B(n1394), .Z(n1393) );
  NANDN U1640 ( .A(A[266]), .B(n1395), .Z(n1394) );
  NANDN U1641 ( .A(n1395), .B(A[266]), .Z(n1392) );
  XOR U1642 ( .A(n1395), .B(n1396), .Z(SUM[266]) );
  XNOR U1643 ( .A(B[266]), .B(A[266]), .Z(n1396) );
  AND U1644 ( .A(n1397), .B(n1398), .Z(n1395) );
  NAND U1645 ( .A(B[265]), .B(n1399), .Z(n1398) );
  NANDN U1646 ( .A(A[265]), .B(n1400), .Z(n1399) );
  NANDN U1647 ( .A(n1400), .B(A[265]), .Z(n1397) );
  XOR U1648 ( .A(n1400), .B(n1401), .Z(SUM[265]) );
  XNOR U1649 ( .A(B[265]), .B(A[265]), .Z(n1401) );
  AND U1650 ( .A(n1402), .B(n1403), .Z(n1400) );
  NAND U1651 ( .A(B[264]), .B(n1404), .Z(n1403) );
  NANDN U1652 ( .A(A[264]), .B(n1405), .Z(n1404) );
  NANDN U1653 ( .A(n1405), .B(A[264]), .Z(n1402) );
  XOR U1654 ( .A(n1405), .B(n1406), .Z(SUM[264]) );
  XNOR U1655 ( .A(B[264]), .B(A[264]), .Z(n1406) );
  AND U1656 ( .A(n1407), .B(n1408), .Z(n1405) );
  NAND U1657 ( .A(B[263]), .B(n1409), .Z(n1408) );
  NANDN U1658 ( .A(A[263]), .B(n1410), .Z(n1409) );
  NANDN U1659 ( .A(n1410), .B(A[263]), .Z(n1407) );
  XOR U1660 ( .A(n1410), .B(n1411), .Z(SUM[263]) );
  XNOR U1661 ( .A(B[263]), .B(A[263]), .Z(n1411) );
  AND U1662 ( .A(n1412), .B(n1413), .Z(n1410) );
  NAND U1663 ( .A(B[262]), .B(n1414), .Z(n1413) );
  NANDN U1664 ( .A(A[262]), .B(n1415), .Z(n1414) );
  NANDN U1665 ( .A(n1415), .B(A[262]), .Z(n1412) );
  XOR U1666 ( .A(n1415), .B(n1416), .Z(SUM[262]) );
  XNOR U1667 ( .A(B[262]), .B(A[262]), .Z(n1416) );
  AND U1668 ( .A(n1417), .B(n1418), .Z(n1415) );
  NAND U1669 ( .A(B[261]), .B(n1419), .Z(n1418) );
  NANDN U1670 ( .A(A[261]), .B(n1420), .Z(n1419) );
  NANDN U1671 ( .A(n1420), .B(A[261]), .Z(n1417) );
  XOR U1672 ( .A(n1420), .B(n1421), .Z(SUM[261]) );
  XNOR U1673 ( .A(B[261]), .B(A[261]), .Z(n1421) );
  AND U1674 ( .A(n1422), .B(n1423), .Z(n1420) );
  NAND U1675 ( .A(B[260]), .B(n1424), .Z(n1423) );
  NANDN U1676 ( .A(A[260]), .B(n1425), .Z(n1424) );
  NANDN U1677 ( .A(n1425), .B(A[260]), .Z(n1422) );
  XOR U1678 ( .A(n1425), .B(n1426), .Z(SUM[260]) );
  XNOR U1679 ( .A(B[260]), .B(A[260]), .Z(n1426) );
  AND U1680 ( .A(n1427), .B(n1428), .Z(n1425) );
  NAND U1681 ( .A(B[259]), .B(n1429), .Z(n1428) );
  NANDN U1682 ( .A(A[259]), .B(n1430), .Z(n1429) );
  NANDN U1683 ( .A(n1430), .B(A[259]), .Z(n1427) );
  XOR U1684 ( .A(n1431), .B(n1432), .Z(SUM[25]) );
  XNOR U1685 ( .A(B[25]), .B(A[25]), .Z(n1432) );
  XOR U1686 ( .A(n1430), .B(n1433), .Z(SUM[259]) );
  XNOR U1687 ( .A(B[259]), .B(A[259]), .Z(n1433) );
  AND U1688 ( .A(n1434), .B(n1435), .Z(n1430) );
  NAND U1689 ( .A(B[258]), .B(n1436), .Z(n1435) );
  NANDN U1690 ( .A(A[258]), .B(n1437), .Z(n1436) );
  NANDN U1691 ( .A(n1437), .B(A[258]), .Z(n1434) );
  XOR U1692 ( .A(n1437), .B(n1438), .Z(SUM[258]) );
  XNOR U1693 ( .A(B[258]), .B(A[258]), .Z(n1438) );
  AND U1694 ( .A(n1439), .B(n1440), .Z(n1437) );
  NAND U1695 ( .A(B[257]), .B(n1441), .Z(n1440) );
  NANDN U1696 ( .A(A[257]), .B(n1442), .Z(n1441) );
  NANDN U1697 ( .A(n1442), .B(A[257]), .Z(n1439) );
  XOR U1698 ( .A(n1442), .B(n1443), .Z(SUM[257]) );
  XNOR U1699 ( .A(B[257]), .B(A[257]), .Z(n1443) );
  AND U1700 ( .A(n1444), .B(n1445), .Z(n1442) );
  NAND U1701 ( .A(B[256]), .B(n1446), .Z(n1445) );
  NANDN U1702 ( .A(A[256]), .B(n1447), .Z(n1446) );
  NANDN U1703 ( .A(n1447), .B(A[256]), .Z(n1444) );
  XOR U1704 ( .A(n1447), .B(n1448), .Z(SUM[256]) );
  XNOR U1705 ( .A(B[256]), .B(A[256]), .Z(n1448) );
  AND U1706 ( .A(n1449), .B(n1450), .Z(n1447) );
  NAND U1707 ( .A(B[255]), .B(n1451), .Z(n1450) );
  NANDN U1708 ( .A(A[255]), .B(n1452), .Z(n1451) );
  NANDN U1709 ( .A(n1452), .B(A[255]), .Z(n1449) );
  XOR U1710 ( .A(n1452), .B(n1453), .Z(SUM[255]) );
  XNOR U1711 ( .A(B[255]), .B(A[255]), .Z(n1453) );
  AND U1712 ( .A(n1454), .B(n1455), .Z(n1452) );
  NAND U1713 ( .A(B[254]), .B(n1456), .Z(n1455) );
  NANDN U1714 ( .A(A[254]), .B(n1457), .Z(n1456) );
  NANDN U1715 ( .A(n1457), .B(A[254]), .Z(n1454) );
  XOR U1716 ( .A(n1457), .B(n1458), .Z(SUM[254]) );
  XNOR U1717 ( .A(B[254]), .B(A[254]), .Z(n1458) );
  AND U1718 ( .A(n1459), .B(n1460), .Z(n1457) );
  NAND U1719 ( .A(B[253]), .B(n1461), .Z(n1460) );
  NANDN U1720 ( .A(A[253]), .B(n1462), .Z(n1461) );
  NANDN U1721 ( .A(n1462), .B(A[253]), .Z(n1459) );
  XOR U1722 ( .A(n1462), .B(n1463), .Z(SUM[253]) );
  XNOR U1723 ( .A(B[253]), .B(A[253]), .Z(n1463) );
  AND U1724 ( .A(n1464), .B(n1465), .Z(n1462) );
  NAND U1725 ( .A(B[252]), .B(n1466), .Z(n1465) );
  NANDN U1726 ( .A(A[252]), .B(n1467), .Z(n1466) );
  NANDN U1727 ( .A(n1467), .B(A[252]), .Z(n1464) );
  XOR U1728 ( .A(n1467), .B(n1468), .Z(SUM[252]) );
  XNOR U1729 ( .A(B[252]), .B(A[252]), .Z(n1468) );
  AND U1730 ( .A(n1469), .B(n1470), .Z(n1467) );
  NAND U1731 ( .A(B[251]), .B(n1471), .Z(n1470) );
  NANDN U1732 ( .A(A[251]), .B(n1472), .Z(n1471) );
  NANDN U1733 ( .A(n1472), .B(A[251]), .Z(n1469) );
  XOR U1734 ( .A(n1472), .B(n1473), .Z(SUM[251]) );
  XNOR U1735 ( .A(B[251]), .B(A[251]), .Z(n1473) );
  AND U1736 ( .A(n1474), .B(n1475), .Z(n1472) );
  NAND U1737 ( .A(B[250]), .B(n1476), .Z(n1475) );
  NANDN U1738 ( .A(A[250]), .B(n1477), .Z(n1476) );
  NANDN U1739 ( .A(n1477), .B(A[250]), .Z(n1474) );
  XOR U1740 ( .A(n1477), .B(n1478), .Z(SUM[250]) );
  XNOR U1741 ( .A(B[250]), .B(A[250]), .Z(n1478) );
  AND U1742 ( .A(n1479), .B(n1480), .Z(n1477) );
  NAND U1743 ( .A(B[249]), .B(n1481), .Z(n1480) );
  NANDN U1744 ( .A(A[249]), .B(n1482), .Z(n1481) );
  NANDN U1745 ( .A(n1482), .B(A[249]), .Z(n1479) );
  XOR U1746 ( .A(n1483), .B(n1484), .Z(SUM[24]) );
  XNOR U1747 ( .A(B[24]), .B(A[24]), .Z(n1484) );
  XOR U1748 ( .A(n1482), .B(n1485), .Z(SUM[249]) );
  XNOR U1749 ( .A(B[249]), .B(A[249]), .Z(n1485) );
  AND U1750 ( .A(n1486), .B(n1487), .Z(n1482) );
  NAND U1751 ( .A(B[248]), .B(n1488), .Z(n1487) );
  NANDN U1752 ( .A(A[248]), .B(n1489), .Z(n1488) );
  NANDN U1753 ( .A(n1489), .B(A[248]), .Z(n1486) );
  XOR U1754 ( .A(n1489), .B(n1490), .Z(SUM[248]) );
  XNOR U1755 ( .A(B[248]), .B(A[248]), .Z(n1490) );
  AND U1756 ( .A(n1491), .B(n1492), .Z(n1489) );
  NAND U1757 ( .A(B[247]), .B(n1493), .Z(n1492) );
  NANDN U1758 ( .A(A[247]), .B(n1494), .Z(n1493) );
  NANDN U1759 ( .A(n1494), .B(A[247]), .Z(n1491) );
  XOR U1760 ( .A(n1494), .B(n1495), .Z(SUM[247]) );
  XNOR U1761 ( .A(B[247]), .B(A[247]), .Z(n1495) );
  AND U1762 ( .A(n1496), .B(n1497), .Z(n1494) );
  NAND U1763 ( .A(B[246]), .B(n1498), .Z(n1497) );
  NANDN U1764 ( .A(A[246]), .B(n1499), .Z(n1498) );
  NANDN U1765 ( .A(n1499), .B(A[246]), .Z(n1496) );
  XOR U1766 ( .A(n1499), .B(n1500), .Z(SUM[246]) );
  XNOR U1767 ( .A(B[246]), .B(A[246]), .Z(n1500) );
  AND U1768 ( .A(n1501), .B(n1502), .Z(n1499) );
  NAND U1769 ( .A(B[245]), .B(n1503), .Z(n1502) );
  NANDN U1770 ( .A(A[245]), .B(n1504), .Z(n1503) );
  NANDN U1771 ( .A(n1504), .B(A[245]), .Z(n1501) );
  XOR U1772 ( .A(n1504), .B(n1505), .Z(SUM[245]) );
  XNOR U1773 ( .A(B[245]), .B(A[245]), .Z(n1505) );
  AND U1774 ( .A(n1506), .B(n1507), .Z(n1504) );
  NAND U1775 ( .A(B[244]), .B(n1508), .Z(n1507) );
  NANDN U1776 ( .A(A[244]), .B(n1509), .Z(n1508) );
  NANDN U1777 ( .A(n1509), .B(A[244]), .Z(n1506) );
  XOR U1778 ( .A(n1509), .B(n1510), .Z(SUM[244]) );
  XNOR U1779 ( .A(B[244]), .B(A[244]), .Z(n1510) );
  AND U1780 ( .A(n1511), .B(n1512), .Z(n1509) );
  NAND U1781 ( .A(B[243]), .B(n1513), .Z(n1512) );
  NANDN U1782 ( .A(A[243]), .B(n1514), .Z(n1513) );
  NANDN U1783 ( .A(n1514), .B(A[243]), .Z(n1511) );
  XOR U1784 ( .A(n1514), .B(n1515), .Z(SUM[243]) );
  XNOR U1785 ( .A(B[243]), .B(A[243]), .Z(n1515) );
  AND U1786 ( .A(n1516), .B(n1517), .Z(n1514) );
  NAND U1787 ( .A(B[242]), .B(n1518), .Z(n1517) );
  NANDN U1788 ( .A(A[242]), .B(n1519), .Z(n1518) );
  NANDN U1789 ( .A(n1519), .B(A[242]), .Z(n1516) );
  XOR U1790 ( .A(n1519), .B(n1520), .Z(SUM[242]) );
  XNOR U1791 ( .A(B[242]), .B(A[242]), .Z(n1520) );
  AND U1792 ( .A(n1521), .B(n1522), .Z(n1519) );
  NAND U1793 ( .A(B[241]), .B(n1523), .Z(n1522) );
  NANDN U1794 ( .A(A[241]), .B(n1524), .Z(n1523) );
  NANDN U1795 ( .A(n1524), .B(A[241]), .Z(n1521) );
  XOR U1796 ( .A(n1524), .B(n1525), .Z(SUM[241]) );
  XNOR U1797 ( .A(B[241]), .B(A[241]), .Z(n1525) );
  AND U1798 ( .A(n1526), .B(n1527), .Z(n1524) );
  NAND U1799 ( .A(B[240]), .B(n1528), .Z(n1527) );
  NANDN U1800 ( .A(A[240]), .B(n1529), .Z(n1528) );
  NANDN U1801 ( .A(n1529), .B(A[240]), .Z(n1526) );
  XOR U1802 ( .A(n1529), .B(n1530), .Z(SUM[240]) );
  XNOR U1803 ( .A(B[240]), .B(A[240]), .Z(n1530) );
  AND U1804 ( .A(n1531), .B(n1532), .Z(n1529) );
  NAND U1805 ( .A(B[239]), .B(n1533), .Z(n1532) );
  NANDN U1806 ( .A(A[239]), .B(n1534), .Z(n1533) );
  NANDN U1807 ( .A(n1534), .B(A[239]), .Z(n1531) );
  XOR U1808 ( .A(n1535), .B(n1536), .Z(SUM[23]) );
  XNOR U1809 ( .A(B[23]), .B(A[23]), .Z(n1536) );
  XOR U1810 ( .A(n1534), .B(n1537), .Z(SUM[239]) );
  XNOR U1811 ( .A(B[239]), .B(A[239]), .Z(n1537) );
  AND U1812 ( .A(n1538), .B(n1539), .Z(n1534) );
  NAND U1813 ( .A(B[238]), .B(n1540), .Z(n1539) );
  NANDN U1814 ( .A(A[238]), .B(n1541), .Z(n1540) );
  NANDN U1815 ( .A(n1541), .B(A[238]), .Z(n1538) );
  XOR U1816 ( .A(n1541), .B(n1542), .Z(SUM[238]) );
  XNOR U1817 ( .A(B[238]), .B(A[238]), .Z(n1542) );
  AND U1818 ( .A(n1543), .B(n1544), .Z(n1541) );
  NAND U1819 ( .A(B[237]), .B(n1545), .Z(n1544) );
  NANDN U1820 ( .A(A[237]), .B(n1546), .Z(n1545) );
  NANDN U1821 ( .A(n1546), .B(A[237]), .Z(n1543) );
  XOR U1822 ( .A(n1546), .B(n1547), .Z(SUM[237]) );
  XNOR U1823 ( .A(B[237]), .B(A[237]), .Z(n1547) );
  AND U1824 ( .A(n1548), .B(n1549), .Z(n1546) );
  NAND U1825 ( .A(B[236]), .B(n1550), .Z(n1549) );
  NANDN U1826 ( .A(A[236]), .B(n1551), .Z(n1550) );
  NANDN U1827 ( .A(n1551), .B(A[236]), .Z(n1548) );
  XOR U1828 ( .A(n1551), .B(n1552), .Z(SUM[236]) );
  XNOR U1829 ( .A(B[236]), .B(A[236]), .Z(n1552) );
  AND U1830 ( .A(n1553), .B(n1554), .Z(n1551) );
  NAND U1831 ( .A(B[235]), .B(n1555), .Z(n1554) );
  NANDN U1832 ( .A(A[235]), .B(n1556), .Z(n1555) );
  NANDN U1833 ( .A(n1556), .B(A[235]), .Z(n1553) );
  XOR U1834 ( .A(n1556), .B(n1557), .Z(SUM[235]) );
  XNOR U1835 ( .A(B[235]), .B(A[235]), .Z(n1557) );
  AND U1836 ( .A(n1558), .B(n1559), .Z(n1556) );
  NAND U1837 ( .A(B[234]), .B(n1560), .Z(n1559) );
  NANDN U1838 ( .A(A[234]), .B(n1561), .Z(n1560) );
  NANDN U1839 ( .A(n1561), .B(A[234]), .Z(n1558) );
  XOR U1840 ( .A(n1561), .B(n1562), .Z(SUM[234]) );
  XNOR U1841 ( .A(B[234]), .B(A[234]), .Z(n1562) );
  AND U1842 ( .A(n1563), .B(n1564), .Z(n1561) );
  NAND U1843 ( .A(B[233]), .B(n1565), .Z(n1564) );
  NANDN U1844 ( .A(A[233]), .B(n1566), .Z(n1565) );
  NANDN U1845 ( .A(n1566), .B(A[233]), .Z(n1563) );
  XOR U1846 ( .A(n1566), .B(n1567), .Z(SUM[233]) );
  XNOR U1847 ( .A(B[233]), .B(A[233]), .Z(n1567) );
  AND U1848 ( .A(n1568), .B(n1569), .Z(n1566) );
  NAND U1849 ( .A(B[232]), .B(n1570), .Z(n1569) );
  NANDN U1850 ( .A(A[232]), .B(n1571), .Z(n1570) );
  NANDN U1851 ( .A(n1571), .B(A[232]), .Z(n1568) );
  XOR U1852 ( .A(n1571), .B(n1572), .Z(SUM[232]) );
  XNOR U1853 ( .A(B[232]), .B(A[232]), .Z(n1572) );
  AND U1854 ( .A(n1573), .B(n1574), .Z(n1571) );
  NAND U1855 ( .A(B[231]), .B(n1575), .Z(n1574) );
  NANDN U1856 ( .A(A[231]), .B(n1576), .Z(n1575) );
  NANDN U1857 ( .A(n1576), .B(A[231]), .Z(n1573) );
  XOR U1858 ( .A(n1576), .B(n1577), .Z(SUM[231]) );
  XNOR U1859 ( .A(B[231]), .B(A[231]), .Z(n1577) );
  AND U1860 ( .A(n1578), .B(n1579), .Z(n1576) );
  NAND U1861 ( .A(B[230]), .B(n1580), .Z(n1579) );
  NANDN U1862 ( .A(A[230]), .B(n1581), .Z(n1580) );
  NANDN U1863 ( .A(n1581), .B(A[230]), .Z(n1578) );
  XOR U1864 ( .A(n1581), .B(n1582), .Z(SUM[230]) );
  XNOR U1865 ( .A(B[230]), .B(A[230]), .Z(n1582) );
  AND U1866 ( .A(n1583), .B(n1584), .Z(n1581) );
  NAND U1867 ( .A(B[229]), .B(n1585), .Z(n1584) );
  NANDN U1868 ( .A(A[229]), .B(n1586), .Z(n1585) );
  NANDN U1869 ( .A(n1586), .B(A[229]), .Z(n1583) );
  XOR U1870 ( .A(n1587), .B(n1588), .Z(SUM[22]) );
  XNOR U1871 ( .A(B[22]), .B(A[22]), .Z(n1588) );
  XOR U1872 ( .A(n1586), .B(n1589), .Z(SUM[229]) );
  XNOR U1873 ( .A(B[229]), .B(A[229]), .Z(n1589) );
  AND U1874 ( .A(n1590), .B(n1591), .Z(n1586) );
  NAND U1875 ( .A(B[228]), .B(n1592), .Z(n1591) );
  NANDN U1876 ( .A(A[228]), .B(n1593), .Z(n1592) );
  NANDN U1877 ( .A(n1593), .B(A[228]), .Z(n1590) );
  XOR U1878 ( .A(n1593), .B(n1594), .Z(SUM[228]) );
  XNOR U1879 ( .A(B[228]), .B(A[228]), .Z(n1594) );
  AND U1880 ( .A(n1595), .B(n1596), .Z(n1593) );
  NAND U1881 ( .A(B[227]), .B(n1597), .Z(n1596) );
  NANDN U1882 ( .A(A[227]), .B(n1598), .Z(n1597) );
  NANDN U1883 ( .A(n1598), .B(A[227]), .Z(n1595) );
  XOR U1884 ( .A(n1598), .B(n1599), .Z(SUM[227]) );
  XNOR U1885 ( .A(B[227]), .B(A[227]), .Z(n1599) );
  AND U1886 ( .A(n1600), .B(n1601), .Z(n1598) );
  NAND U1887 ( .A(B[226]), .B(n1602), .Z(n1601) );
  NANDN U1888 ( .A(A[226]), .B(n1603), .Z(n1602) );
  NANDN U1889 ( .A(n1603), .B(A[226]), .Z(n1600) );
  XOR U1890 ( .A(n1603), .B(n1604), .Z(SUM[226]) );
  XNOR U1891 ( .A(B[226]), .B(A[226]), .Z(n1604) );
  AND U1892 ( .A(n1605), .B(n1606), .Z(n1603) );
  NAND U1893 ( .A(B[225]), .B(n1607), .Z(n1606) );
  NANDN U1894 ( .A(A[225]), .B(n1608), .Z(n1607) );
  NANDN U1895 ( .A(n1608), .B(A[225]), .Z(n1605) );
  XOR U1896 ( .A(n1608), .B(n1609), .Z(SUM[225]) );
  XNOR U1897 ( .A(B[225]), .B(A[225]), .Z(n1609) );
  AND U1898 ( .A(n1610), .B(n1611), .Z(n1608) );
  NAND U1899 ( .A(B[224]), .B(n1612), .Z(n1611) );
  NANDN U1900 ( .A(A[224]), .B(n1613), .Z(n1612) );
  NANDN U1901 ( .A(n1613), .B(A[224]), .Z(n1610) );
  XOR U1902 ( .A(n1613), .B(n1614), .Z(SUM[224]) );
  XNOR U1903 ( .A(B[224]), .B(A[224]), .Z(n1614) );
  AND U1904 ( .A(n1615), .B(n1616), .Z(n1613) );
  NAND U1905 ( .A(B[223]), .B(n1617), .Z(n1616) );
  NANDN U1906 ( .A(A[223]), .B(n1618), .Z(n1617) );
  NANDN U1907 ( .A(n1618), .B(A[223]), .Z(n1615) );
  XOR U1908 ( .A(n1618), .B(n1619), .Z(SUM[223]) );
  XNOR U1909 ( .A(B[223]), .B(A[223]), .Z(n1619) );
  AND U1910 ( .A(n1620), .B(n1621), .Z(n1618) );
  NAND U1911 ( .A(B[222]), .B(n1622), .Z(n1621) );
  NANDN U1912 ( .A(A[222]), .B(n1623), .Z(n1622) );
  NANDN U1913 ( .A(n1623), .B(A[222]), .Z(n1620) );
  XOR U1914 ( .A(n1623), .B(n1624), .Z(SUM[222]) );
  XNOR U1915 ( .A(B[222]), .B(A[222]), .Z(n1624) );
  AND U1916 ( .A(n1625), .B(n1626), .Z(n1623) );
  NAND U1917 ( .A(B[221]), .B(n1627), .Z(n1626) );
  NANDN U1918 ( .A(A[221]), .B(n1628), .Z(n1627) );
  NANDN U1919 ( .A(n1628), .B(A[221]), .Z(n1625) );
  XOR U1920 ( .A(n1628), .B(n1629), .Z(SUM[221]) );
  XNOR U1921 ( .A(B[221]), .B(A[221]), .Z(n1629) );
  AND U1922 ( .A(n1630), .B(n1631), .Z(n1628) );
  NAND U1923 ( .A(B[220]), .B(n1632), .Z(n1631) );
  NANDN U1924 ( .A(A[220]), .B(n1633), .Z(n1632) );
  NANDN U1925 ( .A(n1633), .B(A[220]), .Z(n1630) );
  XOR U1926 ( .A(n1633), .B(n1634), .Z(SUM[220]) );
  XNOR U1927 ( .A(B[220]), .B(A[220]), .Z(n1634) );
  AND U1928 ( .A(n1635), .B(n1636), .Z(n1633) );
  NAND U1929 ( .A(B[219]), .B(n1637), .Z(n1636) );
  NANDN U1930 ( .A(A[219]), .B(n1638), .Z(n1637) );
  NANDN U1931 ( .A(n1638), .B(A[219]), .Z(n1635) );
  XOR U1932 ( .A(n1639), .B(n1640), .Z(SUM[21]) );
  XNOR U1933 ( .A(B[21]), .B(A[21]), .Z(n1640) );
  XOR U1934 ( .A(n1638), .B(n1641), .Z(SUM[219]) );
  XNOR U1935 ( .A(B[219]), .B(A[219]), .Z(n1641) );
  AND U1936 ( .A(n1642), .B(n1643), .Z(n1638) );
  NAND U1937 ( .A(B[218]), .B(n1644), .Z(n1643) );
  NANDN U1938 ( .A(A[218]), .B(n1645), .Z(n1644) );
  NANDN U1939 ( .A(n1645), .B(A[218]), .Z(n1642) );
  XOR U1940 ( .A(n1645), .B(n1646), .Z(SUM[218]) );
  XNOR U1941 ( .A(B[218]), .B(A[218]), .Z(n1646) );
  AND U1942 ( .A(n1647), .B(n1648), .Z(n1645) );
  NAND U1943 ( .A(B[217]), .B(n1649), .Z(n1648) );
  NANDN U1944 ( .A(A[217]), .B(n1650), .Z(n1649) );
  NANDN U1945 ( .A(n1650), .B(A[217]), .Z(n1647) );
  XOR U1946 ( .A(n1650), .B(n1651), .Z(SUM[217]) );
  XNOR U1947 ( .A(B[217]), .B(A[217]), .Z(n1651) );
  AND U1948 ( .A(n1652), .B(n1653), .Z(n1650) );
  NAND U1949 ( .A(B[216]), .B(n1654), .Z(n1653) );
  NANDN U1950 ( .A(A[216]), .B(n1655), .Z(n1654) );
  NANDN U1951 ( .A(n1655), .B(A[216]), .Z(n1652) );
  XOR U1952 ( .A(n1655), .B(n1656), .Z(SUM[216]) );
  XNOR U1953 ( .A(B[216]), .B(A[216]), .Z(n1656) );
  AND U1954 ( .A(n1657), .B(n1658), .Z(n1655) );
  NAND U1955 ( .A(B[215]), .B(n1659), .Z(n1658) );
  NANDN U1956 ( .A(A[215]), .B(n1660), .Z(n1659) );
  NANDN U1957 ( .A(n1660), .B(A[215]), .Z(n1657) );
  XOR U1958 ( .A(n1660), .B(n1661), .Z(SUM[215]) );
  XNOR U1959 ( .A(B[215]), .B(A[215]), .Z(n1661) );
  AND U1960 ( .A(n1662), .B(n1663), .Z(n1660) );
  NAND U1961 ( .A(B[214]), .B(n1664), .Z(n1663) );
  NANDN U1962 ( .A(A[214]), .B(n1665), .Z(n1664) );
  NANDN U1963 ( .A(n1665), .B(A[214]), .Z(n1662) );
  XOR U1964 ( .A(n1665), .B(n1666), .Z(SUM[214]) );
  XNOR U1965 ( .A(B[214]), .B(A[214]), .Z(n1666) );
  AND U1966 ( .A(n1667), .B(n1668), .Z(n1665) );
  NAND U1967 ( .A(B[213]), .B(n1669), .Z(n1668) );
  NANDN U1968 ( .A(A[213]), .B(n1670), .Z(n1669) );
  NANDN U1969 ( .A(n1670), .B(A[213]), .Z(n1667) );
  XOR U1970 ( .A(n1670), .B(n1671), .Z(SUM[213]) );
  XNOR U1971 ( .A(B[213]), .B(A[213]), .Z(n1671) );
  AND U1972 ( .A(n1672), .B(n1673), .Z(n1670) );
  NAND U1973 ( .A(B[212]), .B(n1674), .Z(n1673) );
  NANDN U1974 ( .A(A[212]), .B(n1675), .Z(n1674) );
  NANDN U1975 ( .A(n1675), .B(A[212]), .Z(n1672) );
  XOR U1976 ( .A(n1675), .B(n1676), .Z(SUM[212]) );
  XNOR U1977 ( .A(B[212]), .B(A[212]), .Z(n1676) );
  AND U1978 ( .A(n1677), .B(n1678), .Z(n1675) );
  NAND U1979 ( .A(B[211]), .B(n1679), .Z(n1678) );
  NANDN U1980 ( .A(A[211]), .B(n1680), .Z(n1679) );
  NANDN U1981 ( .A(n1680), .B(A[211]), .Z(n1677) );
  XOR U1982 ( .A(n1680), .B(n1681), .Z(SUM[211]) );
  XNOR U1983 ( .A(B[211]), .B(A[211]), .Z(n1681) );
  AND U1984 ( .A(n1682), .B(n1683), .Z(n1680) );
  NAND U1985 ( .A(B[210]), .B(n1684), .Z(n1683) );
  NANDN U1986 ( .A(A[210]), .B(n1685), .Z(n1684) );
  NANDN U1987 ( .A(n1685), .B(A[210]), .Z(n1682) );
  XOR U1988 ( .A(n1685), .B(n1686), .Z(SUM[210]) );
  XNOR U1989 ( .A(B[210]), .B(A[210]), .Z(n1686) );
  AND U1990 ( .A(n1687), .B(n1688), .Z(n1685) );
  NAND U1991 ( .A(B[209]), .B(n1689), .Z(n1688) );
  NANDN U1992 ( .A(A[209]), .B(n1690), .Z(n1689) );
  NANDN U1993 ( .A(n1690), .B(A[209]), .Z(n1687) );
  XOR U1994 ( .A(n1691), .B(n1692), .Z(SUM[20]) );
  XNOR U1995 ( .A(B[20]), .B(A[20]), .Z(n1692) );
  XOR U1996 ( .A(n1690), .B(n1693), .Z(SUM[209]) );
  XNOR U1997 ( .A(B[209]), .B(A[209]), .Z(n1693) );
  AND U1998 ( .A(n1694), .B(n1695), .Z(n1690) );
  NAND U1999 ( .A(B[208]), .B(n1696), .Z(n1695) );
  NANDN U2000 ( .A(A[208]), .B(n1697), .Z(n1696) );
  NANDN U2001 ( .A(n1697), .B(A[208]), .Z(n1694) );
  XOR U2002 ( .A(n1697), .B(n1698), .Z(SUM[208]) );
  XNOR U2003 ( .A(B[208]), .B(A[208]), .Z(n1698) );
  AND U2004 ( .A(n1699), .B(n1700), .Z(n1697) );
  NAND U2005 ( .A(B[207]), .B(n1701), .Z(n1700) );
  NANDN U2006 ( .A(A[207]), .B(n1702), .Z(n1701) );
  NANDN U2007 ( .A(n1702), .B(A[207]), .Z(n1699) );
  XOR U2008 ( .A(n1702), .B(n1703), .Z(SUM[207]) );
  XNOR U2009 ( .A(B[207]), .B(A[207]), .Z(n1703) );
  AND U2010 ( .A(n1704), .B(n1705), .Z(n1702) );
  NAND U2011 ( .A(B[206]), .B(n1706), .Z(n1705) );
  NANDN U2012 ( .A(A[206]), .B(n1707), .Z(n1706) );
  NANDN U2013 ( .A(n1707), .B(A[206]), .Z(n1704) );
  XOR U2014 ( .A(n1707), .B(n1708), .Z(SUM[206]) );
  XNOR U2015 ( .A(B[206]), .B(A[206]), .Z(n1708) );
  AND U2016 ( .A(n1709), .B(n1710), .Z(n1707) );
  NAND U2017 ( .A(B[205]), .B(n1711), .Z(n1710) );
  NANDN U2018 ( .A(A[205]), .B(n1712), .Z(n1711) );
  NANDN U2019 ( .A(n1712), .B(A[205]), .Z(n1709) );
  XOR U2020 ( .A(n1712), .B(n1713), .Z(SUM[205]) );
  XNOR U2021 ( .A(B[205]), .B(A[205]), .Z(n1713) );
  AND U2022 ( .A(n1714), .B(n1715), .Z(n1712) );
  NAND U2023 ( .A(B[204]), .B(n1716), .Z(n1715) );
  NANDN U2024 ( .A(A[204]), .B(n1717), .Z(n1716) );
  NANDN U2025 ( .A(n1717), .B(A[204]), .Z(n1714) );
  XOR U2026 ( .A(n1717), .B(n1718), .Z(SUM[204]) );
  XNOR U2027 ( .A(B[204]), .B(A[204]), .Z(n1718) );
  AND U2028 ( .A(n1719), .B(n1720), .Z(n1717) );
  NAND U2029 ( .A(B[203]), .B(n1721), .Z(n1720) );
  NANDN U2030 ( .A(A[203]), .B(n1722), .Z(n1721) );
  NANDN U2031 ( .A(n1722), .B(A[203]), .Z(n1719) );
  XOR U2032 ( .A(n1722), .B(n1723), .Z(SUM[203]) );
  XNOR U2033 ( .A(B[203]), .B(A[203]), .Z(n1723) );
  AND U2034 ( .A(n1724), .B(n1725), .Z(n1722) );
  NAND U2035 ( .A(B[202]), .B(n1726), .Z(n1725) );
  NANDN U2036 ( .A(A[202]), .B(n1727), .Z(n1726) );
  NANDN U2037 ( .A(n1727), .B(A[202]), .Z(n1724) );
  XOR U2038 ( .A(n1727), .B(n1728), .Z(SUM[202]) );
  XNOR U2039 ( .A(B[202]), .B(A[202]), .Z(n1728) );
  AND U2040 ( .A(n1729), .B(n1730), .Z(n1727) );
  NAND U2041 ( .A(B[201]), .B(n1731), .Z(n1730) );
  NANDN U2042 ( .A(A[201]), .B(n1732), .Z(n1731) );
  NANDN U2043 ( .A(n1732), .B(A[201]), .Z(n1729) );
  XOR U2044 ( .A(n1732), .B(n1733), .Z(SUM[201]) );
  XNOR U2045 ( .A(B[201]), .B(A[201]), .Z(n1733) );
  AND U2046 ( .A(n1734), .B(n1735), .Z(n1732) );
  NAND U2047 ( .A(B[200]), .B(n1736), .Z(n1735) );
  NANDN U2048 ( .A(A[200]), .B(n1737), .Z(n1736) );
  NANDN U2049 ( .A(n1737), .B(A[200]), .Z(n1734) );
  XOR U2050 ( .A(n1737), .B(n1738), .Z(SUM[200]) );
  XNOR U2051 ( .A(B[200]), .B(A[200]), .Z(n1738) );
  AND U2052 ( .A(n1739), .B(n1740), .Z(n1737) );
  NAND U2053 ( .A(B[199]), .B(n1741), .Z(n1740) );
  NANDN U2054 ( .A(A[199]), .B(n1742), .Z(n1741) );
  NANDN U2055 ( .A(n1742), .B(A[199]), .Z(n1739) );
  XOR U2056 ( .A(B[1]), .B(A[1]), .Z(SUM[1]) );
  XOR U2057 ( .A(n1743), .B(n1744), .Z(SUM[19]) );
  XNOR U2058 ( .A(B[19]), .B(A[19]), .Z(n1744) );
  XOR U2059 ( .A(n1742), .B(n1745), .Z(SUM[199]) );
  XNOR U2060 ( .A(B[199]), .B(A[199]), .Z(n1745) );
  AND U2061 ( .A(n1746), .B(n1747), .Z(n1742) );
  NAND U2062 ( .A(B[198]), .B(n1748), .Z(n1747) );
  NANDN U2063 ( .A(A[198]), .B(n1749), .Z(n1748) );
  NANDN U2064 ( .A(n1749), .B(A[198]), .Z(n1746) );
  XOR U2065 ( .A(n1749), .B(n1750), .Z(SUM[198]) );
  XNOR U2066 ( .A(B[198]), .B(A[198]), .Z(n1750) );
  AND U2067 ( .A(n1751), .B(n1752), .Z(n1749) );
  NAND U2068 ( .A(B[197]), .B(n1753), .Z(n1752) );
  NANDN U2069 ( .A(A[197]), .B(n1754), .Z(n1753) );
  NANDN U2070 ( .A(n1754), .B(A[197]), .Z(n1751) );
  XOR U2071 ( .A(n1754), .B(n1755), .Z(SUM[197]) );
  XNOR U2072 ( .A(B[197]), .B(A[197]), .Z(n1755) );
  AND U2073 ( .A(n1756), .B(n1757), .Z(n1754) );
  NAND U2074 ( .A(B[196]), .B(n1758), .Z(n1757) );
  NANDN U2075 ( .A(A[196]), .B(n1759), .Z(n1758) );
  NANDN U2076 ( .A(n1759), .B(A[196]), .Z(n1756) );
  XOR U2077 ( .A(n1759), .B(n1760), .Z(SUM[196]) );
  XNOR U2078 ( .A(B[196]), .B(A[196]), .Z(n1760) );
  AND U2079 ( .A(n1761), .B(n1762), .Z(n1759) );
  NAND U2080 ( .A(B[195]), .B(n1763), .Z(n1762) );
  NANDN U2081 ( .A(A[195]), .B(n1764), .Z(n1763) );
  NANDN U2082 ( .A(n1764), .B(A[195]), .Z(n1761) );
  XOR U2083 ( .A(n1764), .B(n1765), .Z(SUM[195]) );
  XNOR U2084 ( .A(B[195]), .B(A[195]), .Z(n1765) );
  AND U2085 ( .A(n1766), .B(n1767), .Z(n1764) );
  NAND U2086 ( .A(B[194]), .B(n1768), .Z(n1767) );
  NANDN U2087 ( .A(A[194]), .B(n1769), .Z(n1768) );
  NANDN U2088 ( .A(n1769), .B(A[194]), .Z(n1766) );
  XOR U2089 ( .A(n1769), .B(n1770), .Z(SUM[194]) );
  XNOR U2090 ( .A(B[194]), .B(A[194]), .Z(n1770) );
  AND U2091 ( .A(n1771), .B(n1772), .Z(n1769) );
  NAND U2092 ( .A(B[193]), .B(n1773), .Z(n1772) );
  NANDN U2093 ( .A(A[193]), .B(n1774), .Z(n1773) );
  NANDN U2094 ( .A(n1774), .B(A[193]), .Z(n1771) );
  XOR U2095 ( .A(n1774), .B(n1775), .Z(SUM[193]) );
  XNOR U2096 ( .A(B[193]), .B(A[193]), .Z(n1775) );
  AND U2097 ( .A(n1776), .B(n1777), .Z(n1774) );
  NAND U2098 ( .A(B[192]), .B(n1778), .Z(n1777) );
  NANDN U2099 ( .A(A[192]), .B(n1779), .Z(n1778) );
  NANDN U2100 ( .A(n1779), .B(A[192]), .Z(n1776) );
  XOR U2101 ( .A(n1779), .B(n1780), .Z(SUM[192]) );
  XNOR U2102 ( .A(B[192]), .B(A[192]), .Z(n1780) );
  AND U2103 ( .A(n1781), .B(n1782), .Z(n1779) );
  NAND U2104 ( .A(B[191]), .B(n1783), .Z(n1782) );
  NANDN U2105 ( .A(A[191]), .B(n1784), .Z(n1783) );
  NANDN U2106 ( .A(n1784), .B(A[191]), .Z(n1781) );
  XOR U2107 ( .A(n1784), .B(n1785), .Z(SUM[191]) );
  XNOR U2108 ( .A(B[191]), .B(A[191]), .Z(n1785) );
  AND U2109 ( .A(n1786), .B(n1787), .Z(n1784) );
  NAND U2110 ( .A(B[190]), .B(n1788), .Z(n1787) );
  NANDN U2111 ( .A(A[190]), .B(n1789), .Z(n1788) );
  NANDN U2112 ( .A(n1789), .B(A[190]), .Z(n1786) );
  XOR U2113 ( .A(n1789), .B(n1790), .Z(SUM[190]) );
  XNOR U2114 ( .A(B[190]), .B(A[190]), .Z(n1790) );
  AND U2115 ( .A(n1791), .B(n1792), .Z(n1789) );
  NAND U2116 ( .A(B[189]), .B(n1793), .Z(n1792) );
  NANDN U2117 ( .A(A[189]), .B(n1794), .Z(n1793) );
  NANDN U2118 ( .A(n1794), .B(A[189]), .Z(n1791) );
  XOR U2119 ( .A(n1795), .B(n1796), .Z(SUM[18]) );
  XNOR U2120 ( .A(B[18]), .B(A[18]), .Z(n1796) );
  XOR U2121 ( .A(n1794), .B(n1797), .Z(SUM[189]) );
  XNOR U2122 ( .A(B[189]), .B(A[189]), .Z(n1797) );
  AND U2123 ( .A(n1798), .B(n1799), .Z(n1794) );
  NAND U2124 ( .A(B[188]), .B(n1800), .Z(n1799) );
  NANDN U2125 ( .A(A[188]), .B(n1801), .Z(n1800) );
  NANDN U2126 ( .A(n1801), .B(A[188]), .Z(n1798) );
  XOR U2127 ( .A(n1801), .B(n1802), .Z(SUM[188]) );
  XNOR U2128 ( .A(B[188]), .B(A[188]), .Z(n1802) );
  AND U2129 ( .A(n1803), .B(n1804), .Z(n1801) );
  NAND U2130 ( .A(B[187]), .B(n1805), .Z(n1804) );
  NANDN U2131 ( .A(A[187]), .B(n1806), .Z(n1805) );
  NANDN U2132 ( .A(n1806), .B(A[187]), .Z(n1803) );
  XOR U2133 ( .A(n1806), .B(n1807), .Z(SUM[187]) );
  XNOR U2134 ( .A(B[187]), .B(A[187]), .Z(n1807) );
  AND U2135 ( .A(n1808), .B(n1809), .Z(n1806) );
  NAND U2136 ( .A(B[186]), .B(n1810), .Z(n1809) );
  NANDN U2137 ( .A(A[186]), .B(n1811), .Z(n1810) );
  NANDN U2138 ( .A(n1811), .B(A[186]), .Z(n1808) );
  XOR U2139 ( .A(n1811), .B(n1812), .Z(SUM[186]) );
  XNOR U2140 ( .A(B[186]), .B(A[186]), .Z(n1812) );
  AND U2141 ( .A(n1813), .B(n1814), .Z(n1811) );
  NAND U2142 ( .A(B[185]), .B(n1815), .Z(n1814) );
  NANDN U2143 ( .A(A[185]), .B(n1816), .Z(n1815) );
  NANDN U2144 ( .A(n1816), .B(A[185]), .Z(n1813) );
  XOR U2145 ( .A(n1816), .B(n1817), .Z(SUM[185]) );
  XNOR U2146 ( .A(B[185]), .B(A[185]), .Z(n1817) );
  AND U2147 ( .A(n1818), .B(n1819), .Z(n1816) );
  NAND U2148 ( .A(B[184]), .B(n1820), .Z(n1819) );
  NANDN U2149 ( .A(A[184]), .B(n1821), .Z(n1820) );
  NANDN U2150 ( .A(n1821), .B(A[184]), .Z(n1818) );
  XOR U2151 ( .A(n1821), .B(n1822), .Z(SUM[184]) );
  XNOR U2152 ( .A(B[184]), .B(A[184]), .Z(n1822) );
  AND U2153 ( .A(n1823), .B(n1824), .Z(n1821) );
  NAND U2154 ( .A(B[183]), .B(n1825), .Z(n1824) );
  NANDN U2155 ( .A(A[183]), .B(n1826), .Z(n1825) );
  NANDN U2156 ( .A(n1826), .B(A[183]), .Z(n1823) );
  XOR U2157 ( .A(n1826), .B(n1827), .Z(SUM[183]) );
  XNOR U2158 ( .A(B[183]), .B(A[183]), .Z(n1827) );
  AND U2159 ( .A(n1828), .B(n1829), .Z(n1826) );
  NAND U2160 ( .A(B[182]), .B(n1830), .Z(n1829) );
  NANDN U2161 ( .A(A[182]), .B(n1831), .Z(n1830) );
  NANDN U2162 ( .A(n1831), .B(A[182]), .Z(n1828) );
  XOR U2163 ( .A(n1831), .B(n1832), .Z(SUM[182]) );
  XNOR U2164 ( .A(B[182]), .B(A[182]), .Z(n1832) );
  AND U2165 ( .A(n1833), .B(n1834), .Z(n1831) );
  NAND U2166 ( .A(B[181]), .B(n1835), .Z(n1834) );
  NANDN U2167 ( .A(A[181]), .B(n1836), .Z(n1835) );
  NANDN U2168 ( .A(n1836), .B(A[181]), .Z(n1833) );
  XOR U2169 ( .A(n1836), .B(n1837), .Z(SUM[181]) );
  XNOR U2170 ( .A(B[181]), .B(A[181]), .Z(n1837) );
  AND U2171 ( .A(n1838), .B(n1839), .Z(n1836) );
  NAND U2172 ( .A(B[180]), .B(n1840), .Z(n1839) );
  NANDN U2173 ( .A(A[180]), .B(n1841), .Z(n1840) );
  NANDN U2174 ( .A(n1841), .B(A[180]), .Z(n1838) );
  XOR U2175 ( .A(n1841), .B(n1842), .Z(SUM[180]) );
  XNOR U2176 ( .A(B[180]), .B(A[180]), .Z(n1842) );
  AND U2177 ( .A(n1843), .B(n1844), .Z(n1841) );
  NAND U2178 ( .A(B[179]), .B(n1845), .Z(n1844) );
  NANDN U2179 ( .A(A[179]), .B(n1846), .Z(n1845) );
  NANDN U2180 ( .A(n1846), .B(A[179]), .Z(n1843) );
  XOR U2181 ( .A(n1847), .B(n1848), .Z(SUM[17]) );
  XNOR U2182 ( .A(B[17]), .B(A[17]), .Z(n1848) );
  XOR U2183 ( .A(n1846), .B(n1849), .Z(SUM[179]) );
  XNOR U2184 ( .A(B[179]), .B(A[179]), .Z(n1849) );
  AND U2185 ( .A(n1850), .B(n1851), .Z(n1846) );
  NAND U2186 ( .A(B[178]), .B(n1852), .Z(n1851) );
  NANDN U2187 ( .A(A[178]), .B(n1853), .Z(n1852) );
  NANDN U2188 ( .A(n1853), .B(A[178]), .Z(n1850) );
  XOR U2189 ( .A(n1853), .B(n1854), .Z(SUM[178]) );
  XNOR U2190 ( .A(B[178]), .B(A[178]), .Z(n1854) );
  AND U2191 ( .A(n1855), .B(n1856), .Z(n1853) );
  NAND U2192 ( .A(B[177]), .B(n1857), .Z(n1856) );
  NANDN U2193 ( .A(A[177]), .B(n1858), .Z(n1857) );
  NANDN U2194 ( .A(n1858), .B(A[177]), .Z(n1855) );
  XOR U2195 ( .A(n1858), .B(n1859), .Z(SUM[177]) );
  XNOR U2196 ( .A(B[177]), .B(A[177]), .Z(n1859) );
  AND U2197 ( .A(n1860), .B(n1861), .Z(n1858) );
  NAND U2198 ( .A(B[176]), .B(n1862), .Z(n1861) );
  NANDN U2199 ( .A(A[176]), .B(n1863), .Z(n1862) );
  NANDN U2200 ( .A(n1863), .B(A[176]), .Z(n1860) );
  XOR U2201 ( .A(n1863), .B(n1864), .Z(SUM[176]) );
  XNOR U2202 ( .A(B[176]), .B(A[176]), .Z(n1864) );
  AND U2203 ( .A(n1865), .B(n1866), .Z(n1863) );
  NAND U2204 ( .A(B[175]), .B(n1867), .Z(n1866) );
  NANDN U2205 ( .A(A[175]), .B(n1868), .Z(n1867) );
  NANDN U2206 ( .A(n1868), .B(A[175]), .Z(n1865) );
  XOR U2207 ( .A(n1868), .B(n1869), .Z(SUM[175]) );
  XNOR U2208 ( .A(B[175]), .B(A[175]), .Z(n1869) );
  AND U2209 ( .A(n1870), .B(n1871), .Z(n1868) );
  NAND U2210 ( .A(B[174]), .B(n1872), .Z(n1871) );
  NANDN U2211 ( .A(A[174]), .B(n1873), .Z(n1872) );
  NANDN U2212 ( .A(n1873), .B(A[174]), .Z(n1870) );
  XOR U2213 ( .A(n1873), .B(n1874), .Z(SUM[174]) );
  XNOR U2214 ( .A(B[174]), .B(A[174]), .Z(n1874) );
  AND U2215 ( .A(n1875), .B(n1876), .Z(n1873) );
  NAND U2216 ( .A(B[173]), .B(n1877), .Z(n1876) );
  NANDN U2217 ( .A(A[173]), .B(n1878), .Z(n1877) );
  NANDN U2218 ( .A(n1878), .B(A[173]), .Z(n1875) );
  XOR U2219 ( .A(n1878), .B(n1879), .Z(SUM[173]) );
  XNOR U2220 ( .A(B[173]), .B(A[173]), .Z(n1879) );
  AND U2221 ( .A(n1880), .B(n1881), .Z(n1878) );
  NAND U2222 ( .A(B[172]), .B(n1882), .Z(n1881) );
  NANDN U2223 ( .A(A[172]), .B(n1883), .Z(n1882) );
  NANDN U2224 ( .A(n1883), .B(A[172]), .Z(n1880) );
  XOR U2225 ( .A(n1883), .B(n1884), .Z(SUM[172]) );
  XNOR U2226 ( .A(B[172]), .B(A[172]), .Z(n1884) );
  AND U2227 ( .A(n1885), .B(n1886), .Z(n1883) );
  NAND U2228 ( .A(B[171]), .B(n1887), .Z(n1886) );
  NANDN U2229 ( .A(A[171]), .B(n1888), .Z(n1887) );
  NANDN U2230 ( .A(n1888), .B(A[171]), .Z(n1885) );
  XOR U2231 ( .A(n1888), .B(n1889), .Z(SUM[171]) );
  XNOR U2232 ( .A(B[171]), .B(A[171]), .Z(n1889) );
  AND U2233 ( .A(n1890), .B(n1891), .Z(n1888) );
  NAND U2234 ( .A(B[170]), .B(n1892), .Z(n1891) );
  NANDN U2235 ( .A(A[170]), .B(n1893), .Z(n1892) );
  NANDN U2236 ( .A(n1893), .B(A[170]), .Z(n1890) );
  XOR U2237 ( .A(n1893), .B(n1894), .Z(SUM[170]) );
  XNOR U2238 ( .A(B[170]), .B(A[170]), .Z(n1894) );
  AND U2239 ( .A(n1895), .B(n1896), .Z(n1893) );
  NAND U2240 ( .A(B[169]), .B(n1897), .Z(n1896) );
  NANDN U2241 ( .A(A[169]), .B(n1898), .Z(n1897) );
  NANDN U2242 ( .A(n1898), .B(A[169]), .Z(n1895) );
  XOR U2243 ( .A(n1899), .B(n1900), .Z(SUM[16]) );
  XNOR U2244 ( .A(B[16]), .B(A[16]), .Z(n1900) );
  XOR U2245 ( .A(n1898), .B(n1901), .Z(SUM[169]) );
  XNOR U2246 ( .A(B[169]), .B(A[169]), .Z(n1901) );
  AND U2247 ( .A(n1902), .B(n1903), .Z(n1898) );
  NAND U2248 ( .A(B[168]), .B(n1904), .Z(n1903) );
  NANDN U2249 ( .A(A[168]), .B(n1905), .Z(n1904) );
  NANDN U2250 ( .A(n1905), .B(A[168]), .Z(n1902) );
  XOR U2251 ( .A(n1905), .B(n1906), .Z(SUM[168]) );
  XNOR U2252 ( .A(B[168]), .B(A[168]), .Z(n1906) );
  AND U2253 ( .A(n1907), .B(n1908), .Z(n1905) );
  NAND U2254 ( .A(B[167]), .B(n1909), .Z(n1908) );
  NANDN U2255 ( .A(A[167]), .B(n1910), .Z(n1909) );
  NANDN U2256 ( .A(n1910), .B(A[167]), .Z(n1907) );
  XOR U2257 ( .A(n1910), .B(n1911), .Z(SUM[167]) );
  XNOR U2258 ( .A(B[167]), .B(A[167]), .Z(n1911) );
  AND U2259 ( .A(n1912), .B(n1913), .Z(n1910) );
  NAND U2260 ( .A(B[166]), .B(n1914), .Z(n1913) );
  NANDN U2261 ( .A(A[166]), .B(n1915), .Z(n1914) );
  NANDN U2262 ( .A(n1915), .B(A[166]), .Z(n1912) );
  XOR U2263 ( .A(n1915), .B(n1916), .Z(SUM[166]) );
  XNOR U2264 ( .A(B[166]), .B(A[166]), .Z(n1916) );
  AND U2265 ( .A(n1917), .B(n1918), .Z(n1915) );
  NAND U2266 ( .A(B[165]), .B(n1919), .Z(n1918) );
  NANDN U2267 ( .A(A[165]), .B(n1920), .Z(n1919) );
  NANDN U2268 ( .A(n1920), .B(A[165]), .Z(n1917) );
  XOR U2269 ( .A(n1920), .B(n1921), .Z(SUM[165]) );
  XNOR U2270 ( .A(B[165]), .B(A[165]), .Z(n1921) );
  AND U2271 ( .A(n1922), .B(n1923), .Z(n1920) );
  NAND U2272 ( .A(B[164]), .B(n1924), .Z(n1923) );
  NANDN U2273 ( .A(A[164]), .B(n1925), .Z(n1924) );
  NANDN U2274 ( .A(n1925), .B(A[164]), .Z(n1922) );
  XOR U2275 ( .A(n1925), .B(n1926), .Z(SUM[164]) );
  XNOR U2276 ( .A(B[164]), .B(A[164]), .Z(n1926) );
  AND U2277 ( .A(n1927), .B(n1928), .Z(n1925) );
  NAND U2278 ( .A(B[163]), .B(n1929), .Z(n1928) );
  NANDN U2279 ( .A(A[163]), .B(n1930), .Z(n1929) );
  NANDN U2280 ( .A(n1930), .B(A[163]), .Z(n1927) );
  XOR U2281 ( .A(n1930), .B(n1931), .Z(SUM[163]) );
  XNOR U2282 ( .A(B[163]), .B(A[163]), .Z(n1931) );
  AND U2283 ( .A(n1932), .B(n1933), .Z(n1930) );
  NAND U2284 ( .A(B[162]), .B(n1934), .Z(n1933) );
  NANDN U2285 ( .A(A[162]), .B(n1935), .Z(n1934) );
  NANDN U2286 ( .A(n1935), .B(A[162]), .Z(n1932) );
  XOR U2287 ( .A(n1935), .B(n1936), .Z(SUM[162]) );
  XNOR U2288 ( .A(B[162]), .B(A[162]), .Z(n1936) );
  AND U2289 ( .A(n1937), .B(n1938), .Z(n1935) );
  NAND U2290 ( .A(B[161]), .B(n1939), .Z(n1938) );
  NANDN U2291 ( .A(A[161]), .B(n1940), .Z(n1939) );
  NANDN U2292 ( .A(n1940), .B(A[161]), .Z(n1937) );
  XOR U2293 ( .A(n1940), .B(n1941), .Z(SUM[161]) );
  XNOR U2294 ( .A(B[161]), .B(A[161]), .Z(n1941) );
  AND U2295 ( .A(n1942), .B(n1943), .Z(n1940) );
  NAND U2296 ( .A(B[160]), .B(n1944), .Z(n1943) );
  NANDN U2297 ( .A(A[160]), .B(n1945), .Z(n1944) );
  NANDN U2298 ( .A(n1945), .B(A[160]), .Z(n1942) );
  XOR U2299 ( .A(n1945), .B(n1946), .Z(SUM[160]) );
  XNOR U2300 ( .A(B[160]), .B(A[160]), .Z(n1946) );
  AND U2301 ( .A(n1947), .B(n1948), .Z(n1945) );
  NAND U2302 ( .A(B[159]), .B(n1949), .Z(n1948) );
  NANDN U2303 ( .A(A[159]), .B(n1950), .Z(n1949) );
  NANDN U2304 ( .A(n1950), .B(A[159]), .Z(n1947) );
  XOR U2305 ( .A(n1951), .B(n1952), .Z(SUM[15]) );
  XNOR U2306 ( .A(B[15]), .B(A[15]), .Z(n1952) );
  XOR U2307 ( .A(n1950), .B(n1953), .Z(SUM[159]) );
  XNOR U2308 ( .A(B[159]), .B(A[159]), .Z(n1953) );
  AND U2309 ( .A(n1954), .B(n1955), .Z(n1950) );
  NAND U2310 ( .A(B[158]), .B(n1956), .Z(n1955) );
  NANDN U2311 ( .A(A[158]), .B(n1957), .Z(n1956) );
  NANDN U2312 ( .A(n1957), .B(A[158]), .Z(n1954) );
  XOR U2313 ( .A(n1957), .B(n1958), .Z(SUM[158]) );
  XNOR U2314 ( .A(B[158]), .B(A[158]), .Z(n1958) );
  AND U2315 ( .A(n1959), .B(n1960), .Z(n1957) );
  NAND U2316 ( .A(B[157]), .B(n1961), .Z(n1960) );
  NANDN U2317 ( .A(A[157]), .B(n1962), .Z(n1961) );
  NANDN U2318 ( .A(n1962), .B(A[157]), .Z(n1959) );
  XOR U2319 ( .A(n1962), .B(n1963), .Z(SUM[157]) );
  XNOR U2320 ( .A(B[157]), .B(A[157]), .Z(n1963) );
  AND U2321 ( .A(n1964), .B(n1965), .Z(n1962) );
  NAND U2322 ( .A(B[156]), .B(n1966), .Z(n1965) );
  NANDN U2323 ( .A(A[156]), .B(n1967), .Z(n1966) );
  NANDN U2324 ( .A(n1967), .B(A[156]), .Z(n1964) );
  XOR U2325 ( .A(n1967), .B(n1968), .Z(SUM[156]) );
  XNOR U2326 ( .A(B[156]), .B(A[156]), .Z(n1968) );
  AND U2327 ( .A(n1969), .B(n1970), .Z(n1967) );
  NAND U2328 ( .A(B[155]), .B(n1971), .Z(n1970) );
  NANDN U2329 ( .A(A[155]), .B(n1972), .Z(n1971) );
  NANDN U2330 ( .A(n1972), .B(A[155]), .Z(n1969) );
  XOR U2331 ( .A(n1972), .B(n1973), .Z(SUM[155]) );
  XNOR U2332 ( .A(B[155]), .B(A[155]), .Z(n1973) );
  AND U2333 ( .A(n1974), .B(n1975), .Z(n1972) );
  NAND U2334 ( .A(B[154]), .B(n1976), .Z(n1975) );
  NANDN U2335 ( .A(A[154]), .B(n1977), .Z(n1976) );
  NANDN U2336 ( .A(n1977), .B(A[154]), .Z(n1974) );
  XOR U2337 ( .A(n1977), .B(n1978), .Z(SUM[154]) );
  XNOR U2338 ( .A(B[154]), .B(A[154]), .Z(n1978) );
  AND U2339 ( .A(n1979), .B(n1980), .Z(n1977) );
  NAND U2340 ( .A(B[153]), .B(n1981), .Z(n1980) );
  NANDN U2341 ( .A(A[153]), .B(n1982), .Z(n1981) );
  NANDN U2342 ( .A(n1982), .B(A[153]), .Z(n1979) );
  XOR U2343 ( .A(n1982), .B(n1983), .Z(SUM[153]) );
  XNOR U2344 ( .A(B[153]), .B(A[153]), .Z(n1983) );
  AND U2345 ( .A(n1984), .B(n1985), .Z(n1982) );
  NAND U2346 ( .A(B[152]), .B(n1986), .Z(n1985) );
  NANDN U2347 ( .A(A[152]), .B(n1987), .Z(n1986) );
  NANDN U2348 ( .A(n1987), .B(A[152]), .Z(n1984) );
  XOR U2349 ( .A(n1987), .B(n1988), .Z(SUM[152]) );
  XNOR U2350 ( .A(B[152]), .B(A[152]), .Z(n1988) );
  AND U2351 ( .A(n1989), .B(n1990), .Z(n1987) );
  NAND U2352 ( .A(B[151]), .B(n1991), .Z(n1990) );
  NANDN U2353 ( .A(A[151]), .B(n1992), .Z(n1991) );
  NANDN U2354 ( .A(n1992), .B(A[151]), .Z(n1989) );
  XOR U2355 ( .A(n1992), .B(n1993), .Z(SUM[151]) );
  XNOR U2356 ( .A(B[151]), .B(A[151]), .Z(n1993) );
  AND U2357 ( .A(n1994), .B(n1995), .Z(n1992) );
  NAND U2358 ( .A(B[150]), .B(n1996), .Z(n1995) );
  NANDN U2359 ( .A(A[150]), .B(n1997), .Z(n1996) );
  NANDN U2360 ( .A(n1997), .B(A[150]), .Z(n1994) );
  XOR U2361 ( .A(n1997), .B(n1998), .Z(SUM[150]) );
  XNOR U2362 ( .A(B[150]), .B(A[150]), .Z(n1998) );
  AND U2363 ( .A(n1999), .B(n2000), .Z(n1997) );
  NAND U2364 ( .A(B[149]), .B(n2001), .Z(n2000) );
  NANDN U2365 ( .A(A[149]), .B(n2002), .Z(n2001) );
  NANDN U2366 ( .A(n2002), .B(A[149]), .Z(n1999) );
  XOR U2367 ( .A(n2003), .B(n2004), .Z(SUM[14]) );
  XNOR U2368 ( .A(B[14]), .B(A[14]), .Z(n2004) );
  XOR U2369 ( .A(n2002), .B(n2005), .Z(SUM[149]) );
  XNOR U2370 ( .A(B[149]), .B(A[149]), .Z(n2005) );
  AND U2371 ( .A(n2006), .B(n2007), .Z(n2002) );
  NAND U2372 ( .A(B[148]), .B(n2008), .Z(n2007) );
  NANDN U2373 ( .A(A[148]), .B(n2009), .Z(n2008) );
  NANDN U2374 ( .A(n2009), .B(A[148]), .Z(n2006) );
  XOR U2375 ( .A(n2009), .B(n2010), .Z(SUM[148]) );
  XNOR U2376 ( .A(B[148]), .B(A[148]), .Z(n2010) );
  AND U2377 ( .A(n2011), .B(n2012), .Z(n2009) );
  NAND U2378 ( .A(B[147]), .B(n2013), .Z(n2012) );
  NANDN U2379 ( .A(A[147]), .B(n2014), .Z(n2013) );
  NANDN U2380 ( .A(n2014), .B(A[147]), .Z(n2011) );
  XOR U2381 ( .A(n2014), .B(n2015), .Z(SUM[147]) );
  XNOR U2382 ( .A(B[147]), .B(A[147]), .Z(n2015) );
  AND U2383 ( .A(n2016), .B(n2017), .Z(n2014) );
  NAND U2384 ( .A(B[146]), .B(n2018), .Z(n2017) );
  NANDN U2385 ( .A(A[146]), .B(n2019), .Z(n2018) );
  NANDN U2386 ( .A(n2019), .B(A[146]), .Z(n2016) );
  XOR U2387 ( .A(n2019), .B(n2020), .Z(SUM[146]) );
  XNOR U2388 ( .A(B[146]), .B(A[146]), .Z(n2020) );
  AND U2389 ( .A(n2021), .B(n2022), .Z(n2019) );
  NAND U2390 ( .A(B[145]), .B(n2023), .Z(n2022) );
  NANDN U2391 ( .A(A[145]), .B(n2024), .Z(n2023) );
  NANDN U2392 ( .A(n2024), .B(A[145]), .Z(n2021) );
  XOR U2393 ( .A(n2024), .B(n2025), .Z(SUM[145]) );
  XNOR U2394 ( .A(B[145]), .B(A[145]), .Z(n2025) );
  AND U2395 ( .A(n2026), .B(n2027), .Z(n2024) );
  NAND U2396 ( .A(B[144]), .B(n2028), .Z(n2027) );
  NANDN U2397 ( .A(A[144]), .B(n2029), .Z(n2028) );
  NANDN U2398 ( .A(n2029), .B(A[144]), .Z(n2026) );
  XOR U2399 ( .A(n2029), .B(n2030), .Z(SUM[144]) );
  XNOR U2400 ( .A(B[144]), .B(A[144]), .Z(n2030) );
  AND U2401 ( .A(n2031), .B(n2032), .Z(n2029) );
  NAND U2402 ( .A(B[143]), .B(n2033), .Z(n2032) );
  NANDN U2403 ( .A(A[143]), .B(n2034), .Z(n2033) );
  NANDN U2404 ( .A(n2034), .B(A[143]), .Z(n2031) );
  XOR U2405 ( .A(n2034), .B(n2035), .Z(SUM[143]) );
  XNOR U2406 ( .A(B[143]), .B(A[143]), .Z(n2035) );
  AND U2407 ( .A(n2036), .B(n2037), .Z(n2034) );
  NAND U2408 ( .A(B[142]), .B(n2038), .Z(n2037) );
  NANDN U2409 ( .A(A[142]), .B(n2039), .Z(n2038) );
  NANDN U2410 ( .A(n2039), .B(A[142]), .Z(n2036) );
  XOR U2411 ( .A(n2039), .B(n2040), .Z(SUM[142]) );
  XNOR U2412 ( .A(B[142]), .B(A[142]), .Z(n2040) );
  AND U2413 ( .A(n2041), .B(n2042), .Z(n2039) );
  NAND U2414 ( .A(B[141]), .B(n2043), .Z(n2042) );
  NANDN U2415 ( .A(A[141]), .B(n2044), .Z(n2043) );
  NANDN U2416 ( .A(n2044), .B(A[141]), .Z(n2041) );
  XOR U2417 ( .A(n2044), .B(n2045), .Z(SUM[141]) );
  XNOR U2418 ( .A(B[141]), .B(A[141]), .Z(n2045) );
  AND U2419 ( .A(n2046), .B(n2047), .Z(n2044) );
  NAND U2420 ( .A(B[140]), .B(n2048), .Z(n2047) );
  NANDN U2421 ( .A(A[140]), .B(n2049), .Z(n2048) );
  NANDN U2422 ( .A(n2049), .B(A[140]), .Z(n2046) );
  XOR U2423 ( .A(n2049), .B(n2050), .Z(SUM[140]) );
  XNOR U2424 ( .A(B[140]), .B(A[140]), .Z(n2050) );
  AND U2425 ( .A(n2051), .B(n2052), .Z(n2049) );
  NAND U2426 ( .A(B[139]), .B(n2053), .Z(n2052) );
  NANDN U2427 ( .A(A[139]), .B(n2054), .Z(n2053) );
  NANDN U2428 ( .A(n2054), .B(A[139]), .Z(n2051) );
  XOR U2429 ( .A(n2055), .B(n2056), .Z(SUM[13]) );
  XNOR U2430 ( .A(B[13]), .B(A[13]), .Z(n2056) );
  XOR U2431 ( .A(n2054), .B(n2057), .Z(SUM[139]) );
  XNOR U2432 ( .A(B[139]), .B(A[139]), .Z(n2057) );
  AND U2433 ( .A(n2058), .B(n2059), .Z(n2054) );
  NAND U2434 ( .A(B[138]), .B(n2060), .Z(n2059) );
  NANDN U2435 ( .A(A[138]), .B(n2061), .Z(n2060) );
  NANDN U2436 ( .A(n2061), .B(A[138]), .Z(n2058) );
  XOR U2437 ( .A(n2061), .B(n2062), .Z(SUM[138]) );
  XNOR U2438 ( .A(B[138]), .B(A[138]), .Z(n2062) );
  AND U2439 ( .A(n2063), .B(n2064), .Z(n2061) );
  NAND U2440 ( .A(B[137]), .B(n2065), .Z(n2064) );
  NANDN U2441 ( .A(A[137]), .B(n2066), .Z(n2065) );
  NANDN U2442 ( .A(n2066), .B(A[137]), .Z(n2063) );
  XOR U2443 ( .A(n2066), .B(n2067), .Z(SUM[137]) );
  XNOR U2444 ( .A(B[137]), .B(A[137]), .Z(n2067) );
  AND U2445 ( .A(n2068), .B(n2069), .Z(n2066) );
  NAND U2446 ( .A(B[136]), .B(n2070), .Z(n2069) );
  NANDN U2447 ( .A(A[136]), .B(n2071), .Z(n2070) );
  NANDN U2448 ( .A(n2071), .B(A[136]), .Z(n2068) );
  XOR U2449 ( .A(n2071), .B(n2072), .Z(SUM[136]) );
  XNOR U2450 ( .A(B[136]), .B(A[136]), .Z(n2072) );
  AND U2451 ( .A(n2073), .B(n2074), .Z(n2071) );
  NAND U2452 ( .A(B[135]), .B(n2075), .Z(n2074) );
  NANDN U2453 ( .A(A[135]), .B(n2076), .Z(n2075) );
  NANDN U2454 ( .A(n2076), .B(A[135]), .Z(n2073) );
  XOR U2455 ( .A(n2076), .B(n2077), .Z(SUM[135]) );
  XNOR U2456 ( .A(B[135]), .B(A[135]), .Z(n2077) );
  AND U2457 ( .A(n2078), .B(n2079), .Z(n2076) );
  NAND U2458 ( .A(B[134]), .B(n2080), .Z(n2079) );
  NANDN U2459 ( .A(A[134]), .B(n2081), .Z(n2080) );
  NANDN U2460 ( .A(n2081), .B(A[134]), .Z(n2078) );
  XOR U2461 ( .A(n2081), .B(n2082), .Z(SUM[134]) );
  XNOR U2462 ( .A(B[134]), .B(A[134]), .Z(n2082) );
  AND U2463 ( .A(n2083), .B(n2084), .Z(n2081) );
  NAND U2464 ( .A(B[133]), .B(n2085), .Z(n2084) );
  NANDN U2465 ( .A(A[133]), .B(n2086), .Z(n2085) );
  NANDN U2466 ( .A(n2086), .B(A[133]), .Z(n2083) );
  XOR U2467 ( .A(n2086), .B(n2087), .Z(SUM[133]) );
  XNOR U2468 ( .A(B[133]), .B(A[133]), .Z(n2087) );
  AND U2469 ( .A(n2088), .B(n2089), .Z(n2086) );
  NAND U2470 ( .A(B[132]), .B(n2090), .Z(n2089) );
  NANDN U2471 ( .A(A[132]), .B(n2091), .Z(n2090) );
  NANDN U2472 ( .A(n2091), .B(A[132]), .Z(n2088) );
  XOR U2473 ( .A(n2091), .B(n2092), .Z(SUM[132]) );
  XNOR U2474 ( .A(B[132]), .B(A[132]), .Z(n2092) );
  AND U2475 ( .A(n2093), .B(n2094), .Z(n2091) );
  NAND U2476 ( .A(B[131]), .B(n2095), .Z(n2094) );
  NANDN U2477 ( .A(A[131]), .B(n2096), .Z(n2095) );
  NANDN U2478 ( .A(n2096), .B(A[131]), .Z(n2093) );
  XOR U2479 ( .A(n2096), .B(n2097), .Z(SUM[131]) );
  XNOR U2480 ( .A(B[131]), .B(A[131]), .Z(n2097) );
  AND U2481 ( .A(n2098), .B(n2099), .Z(n2096) );
  NAND U2482 ( .A(B[130]), .B(n2100), .Z(n2099) );
  NANDN U2483 ( .A(A[130]), .B(n2101), .Z(n2100) );
  NANDN U2484 ( .A(n2101), .B(A[130]), .Z(n2098) );
  XOR U2485 ( .A(n2101), .B(n2102), .Z(SUM[130]) );
  XNOR U2486 ( .A(B[130]), .B(A[130]), .Z(n2102) );
  AND U2487 ( .A(n2103), .B(n2104), .Z(n2101) );
  NAND U2488 ( .A(B[129]), .B(n2105), .Z(n2104) );
  NANDN U2489 ( .A(A[129]), .B(n2106), .Z(n2105) );
  NANDN U2490 ( .A(n2106), .B(A[129]), .Z(n2103) );
  XOR U2491 ( .A(n2107), .B(n2108), .Z(SUM[12]) );
  XNOR U2492 ( .A(B[12]), .B(A[12]), .Z(n2108) );
  XOR U2493 ( .A(n2106), .B(n2109), .Z(SUM[129]) );
  XNOR U2494 ( .A(B[129]), .B(A[129]), .Z(n2109) );
  AND U2495 ( .A(n2110), .B(n2111), .Z(n2106) );
  NAND U2496 ( .A(B[128]), .B(n2112), .Z(n2111) );
  NANDN U2497 ( .A(A[128]), .B(n2113), .Z(n2112) );
  NANDN U2498 ( .A(n2113), .B(A[128]), .Z(n2110) );
  XOR U2499 ( .A(n2113), .B(n2114), .Z(SUM[128]) );
  XNOR U2500 ( .A(B[128]), .B(A[128]), .Z(n2114) );
  AND U2501 ( .A(n2115), .B(n2116), .Z(n2113) );
  NAND U2502 ( .A(B[127]), .B(n2117), .Z(n2116) );
  NANDN U2503 ( .A(A[127]), .B(n2118), .Z(n2117) );
  NANDN U2504 ( .A(n2118), .B(A[127]), .Z(n2115) );
  XOR U2505 ( .A(n2118), .B(n2119), .Z(SUM[127]) );
  XNOR U2506 ( .A(B[127]), .B(A[127]), .Z(n2119) );
  AND U2507 ( .A(n2120), .B(n2121), .Z(n2118) );
  NAND U2508 ( .A(B[126]), .B(n2122), .Z(n2121) );
  NANDN U2509 ( .A(A[126]), .B(n2123), .Z(n2122) );
  NANDN U2510 ( .A(n2123), .B(A[126]), .Z(n2120) );
  XOR U2511 ( .A(n2123), .B(n2124), .Z(SUM[126]) );
  XNOR U2512 ( .A(B[126]), .B(A[126]), .Z(n2124) );
  AND U2513 ( .A(n2125), .B(n2126), .Z(n2123) );
  NAND U2514 ( .A(B[125]), .B(n2127), .Z(n2126) );
  NANDN U2515 ( .A(A[125]), .B(n2128), .Z(n2127) );
  NANDN U2516 ( .A(n2128), .B(A[125]), .Z(n2125) );
  XOR U2517 ( .A(n2128), .B(n2129), .Z(SUM[125]) );
  XNOR U2518 ( .A(B[125]), .B(A[125]), .Z(n2129) );
  AND U2519 ( .A(n2130), .B(n2131), .Z(n2128) );
  NAND U2520 ( .A(B[124]), .B(n2132), .Z(n2131) );
  NANDN U2521 ( .A(A[124]), .B(n2133), .Z(n2132) );
  NANDN U2522 ( .A(n2133), .B(A[124]), .Z(n2130) );
  XOR U2523 ( .A(n2133), .B(n2134), .Z(SUM[124]) );
  XNOR U2524 ( .A(B[124]), .B(A[124]), .Z(n2134) );
  AND U2525 ( .A(n2135), .B(n2136), .Z(n2133) );
  NAND U2526 ( .A(B[123]), .B(n2137), .Z(n2136) );
  NANDN U2527 ( .A(A[123]), .B(n2138), .Z(n2137) );
  NANDN U2528 ( .A(n2138), .B(A[123]), .Z(n2135) );
  XOR U2529 ( .A(n2138), .B(n2139), .Z(SUM[123]) );
  XNOR U2530 ( .A(B[123]), .B(A[123]), .Z(n2139) );
  AND U2531 ( .A(n2140), .B(n2141), .Z(n2138) );
  NAND U2532 ( .A(B[122]), .B(n2142), .Z(n2141) );
  NANDN U2533 ( .A(A[122]), .B(n2143), .Z(n2142) );
  NANDN U2534 ( .A(n2143), .B(A[122]), .Z(n2140) );
  XOR U2535 ( .A(n2143), .B(n2144), .Z(SUM[122]) );
  XNOR U2536 ( .A(B[122]), .B(A[122]), .Z(n2144) );
  AND U2537 ( .A(n2145), .B(n2146), .Z(n2143) );
  NAND U2538 ( .A(B[121]), .B(n2147), .Z(n2146) );
  NANDN U2539 ( .A(A[121]), .B(n2148), .Z(n2147) );
  NANDN U2540 ( .A(n2148), .B(A[121]), .Z(n2145) );
  XOR U2541 ( .A(n2148), .B(n2149), .Z(SUM[121]) );
  XNOR U2542 ( .A(B[121]), .B(A[121]), .Z(n2149) );
  AND U2543 ( .A(n2150), .B(n2151), .Z(n2148) );
  NAND U2544 ( .A(B[120]), .B(n2152), .Z(n2151) );
  NANDN U2545 ( .A(A[120]), .B(n2153), .Z(n2152) );
  NANDN U2546 ( .A(n2153), .B(A[120]), .Z(n2150) );
  XOR U2547 ( .A(n2153), .B(n2154), .Z(SUM[120]) );
  XNOR U2548 ( .A(B[120]), .B(A[120]), .Z(n2154) );
  AND U2549 ( .A(n2155), .B(n2156), .Z(n2153) );
  NAND U2550 ( .A(B[119]), .B(n2157), .Z(n2156) );
  NANDN U2551 ( .A(A[119]), .B(n2158), .Z(n2157) );
  NANDN U2552 ( .A(n2158), .B(A[119]), .Z(n2155) );
  XOR U2553 ( .A(n2159), .B(n2160), .Z(SUM[11]) );
  XNOR U2554 ( .A(B[11]), .B(A[11]), .Z(n2160) );
  XOR U2555 ( .A(n2158), .B(n2161), .Z(SUM[119]) );
  XNOR U2556 ( .A(B[119]), .B(A[119]), .Z(n2161) );
  AND U2557 ( .A(n2162), .B(n2163), .Z(n2158) );
  NAND U2558 ( .A(B[118]), .B(n2164), .Z(n2163) );
  NANDN U2559 ( .A(A[118]), .B(n2165), .Z(n2164) );
  NANDN U2560 ( .A(n2165), .B(A[118]), .Z(n2162) );
  XOR U2561 ( .A(n2165), .B(n2166), .Z(SUM[118]) );
  XNOR U2562 ( .A(B[118]), .B(A[118]), .Z(n2166) );
  AND U2563 ( .A(n2167), .B(n2168), .Z(n2165) );
  NAND U2564 ( .A(B[117]), .B(n2169), .Z(n2168) );
  NANDN U2565 ( .A(A[117]), .B(n2170), .Z(n2169) );
  NANDN U2566 ( .A(n2170), .B(A[117]), .Z(n2167) );
  XOR U2567 ( .A(n2170), .B(n2171), .Z(SUM[117]) );
  XNOR U2568 ( .A(B[117]), .B(A[117]), .Z(n2171) );
  AND U2569 ( .A(n2172), .B(n2173), .Z(n2170) );
  NAND U2570 ( .A(B[116]), .B(n2174), .Z(n2173) );
  NANDN U2571 ( .A(A[116]), .B(n2175), .Z(n2174) );
  NANDN U2572 ( .A(n2175), .B(A[116]), .Z(n2172) );
  XOR U2573 ( .A(n2175), .B(n2176), .Z(SUM[116]) );
  XNOR U2574 ( .A(B[116]), .B(A[116]), .Z(n2176) );
  AND U2575 ( .A(n2177), .B(n2178), .Z(n2175) );
  NAND U2576 ( .A(B[115]), .B(n2179), .Z(n2178) );
  NANDN U2577 ( .A(A[115]), .B(n2180), .Z(n2179) );
  NANDN U2578 ( .A(n2180), .B(A[115]), .Z(n2177) );
  XOR U2579 ( .A(n2180), .B(n2181), .Z(SUM[115]) );
  XNOR U2580 ( .A(B[115]), .B(A[115]), .Z(n2181) );
  AND U2581 ( .A(n2182), .B(n2183), .Z(n2180) );
  NAND U2582 ( .A(B[114]), .B(n2184), .Z(n2183) );
  NANDN U2583 ( .A(A[114]), .B(n2185), .Z(n2184) );
  NANDN U2584 ( .A(n2185), .B(A[114]), .Z(n2182) );
  XOR U2585 ( .A(n2185), .B(n2186), .Z(SUM[114]) );
  XNOR U2586 ( .A(B[114]), .B(A[114]), .Z(n2186) );
  AND U2587 ( .A(n2187), .B(n2188), .Z(n2185) );
  NAND U2588 ( .A(B[113]), .B(n2189), .Z(n2188) );
  NANDN U2589 ( .A(A[113]), .B(n2190), .Z(n2189) );
  NANDN U2590 ( .A(n2190), .B(A[113]), .Z(n2187) );
  XOR U2591 ( .A(n2190), .B(n2191), .Z(SUM[113]) );
  XNOR U2592 ( .A(B[113]), .B(A[113]), .Z(n2191) );
  AND U2593 ( .A(n2192), .B(n2193), .Z(n2190) );
  NAND U2594 ( .A(B[112]), .B(n2194), .Z(n2193) );
  NANDN U2595 ( .A(A[112]), .B(n2195), .Z(n2194) );
  NANDN U2596 ( .A(n2195), .B(A[112]), .Z(n2192) );
  XOR U2597 ( .A(n2195), .B(n2196), .Z(SUM[112]) );
  XNOR U2598 ( .A(B[112]), .B(A[112]), .Z(n2196) );
  AND U2599 ( .A(n2197), .B(n2198), .Z(n2195) );
  NAND U2600 ( .A(B[111]), .B(n2199), .Z(n2198) );
  NANDN U2601 ( .A(A[111]), .B(n2200), .Z(n2199) );
  NANDN U2602 ( .A(n2200), .B(A[111]), .Z(n2197) );
  XOR U2603 ( .A(n2200), .B(n2201), .Z(SUM[111]) );
  XNOR U2604 ( .A(B[111]), .B(A[111]), .Z(n2201) );
  AND U2605 ( .A(n2202), .B(n2203), .Z(n2200) );
  NAND U2606 ( .A(B[110]), .B(n2204), .Z(n2203) );
  NANDN U2607 ( .A(A[110]), .B(n2205), .Z(n2204) );
  NANDN U2608 ( .A(n2205), .B(A[110]), .Z(n2202) );
  XOR U2609 ( .A(n2205), .B(n2206), .Z(SUM[110]) );
  XNOR U2610 ( .A(B[110]), .B(A[110]), .Z(n2206) );
  AND U2611 ( .A(n2207), .B(n2208), .Z(n2205) );
  NAND U2612 ( .A(B[109]), .B(n2209), .Z(n2208) );
  NANDN U2613 ( .A(A[109]), .B(n2210), .Z(n2209) );
  NANDN U2614 ( .A(n2210), .B(A[109]), .Z(n2207) );
  XOR U2615 ( .A(n2211), .B(n2212), .Z(SUM[10]) );
  XNOR U2616 ( .A(B[10]), .B(A[10]), .Z(n2212) );
  XOR U2617 ( .A(n2210), .B(n2213), .Z(SUM[109]) );
  XNOR U2618 ( .A(B[109]), .B(A[109]), .Z(n2213) );
  AND U2619 ( .A(n2214), .B(n2215), .Z(n2210) );
  NAND U2620 ( .A(B[108]), .B(n2216), .Z(n2215) );
  NANDN U2621 ( .A(A[108]), .B(n2217), .Z(n2216) );
  NANDN U2622 ( .A(n2217), .B(A[108]), .Z(n2214) );
  XOR U2623 ( .A(n2217), .B(n2218), .Z(SUM[108]) );
  XNOR U2624 ( .A(B[108]), .B(A[108]), .Z(n2218) );
  AND U2625 ( .A(n2219), .B(n2220), .Z(n2217) );
  NAND U2626 ( .A(B[107]), .B(n2221), .Z(n2220) );
  NANDN U2627 ( .A(A[107]), .B(n2222), .Z(n2221) );
  NANDN U2628 ( .A(n2222), .B(A[107]), .Z(n2219) );
  XOR U2629 ( .A(n2222), .B(n2223), .Z(SUM[107]) );
  XNOR U2630 ( .A(B[107]), .B(A[107]), .Z(n2223) );
  AND U2631 ( .A(n2224), .B(n2225), .Z(n2222) );
  NAND U2632 ( .A(B[106]), .B(n2226), .Z(n2225) );
  NANDN U2633 ( .A(A[106]), .B(n2227), .Z(n2226) );
  NANDN U2634 ( .A(n2227), .B(A[106]), .Z(n2224) );
  XOR U2635 ( .A(n2227), .B(n2228), .Z(SUM[106]) );
  XNOR U2636 ( .A(B[106]), .B(A[106]), .Z(n2228) );
  AND U2637 ( .A(n2229), .B(n2230), .Z(n2227) );
  NAND U2638 ( .A(B[105]), .B(n2231), .Z(n2230) );
  NANDN U2639 ( .A(A[105]), .B(n2232), .Z(n2231) );
  NANDN U2640 ( .A(n2232), .B(A[105]), .Z(n2229) );
  XOR U2641 ( .A(n2232), .B(n2233), .Z(SUM[105]) );
  XNOR U2642 ( .A(B[105]), .B(A[105]), .Z(n2233) );
  AND U2643 ( .A(n2234), .B(n2235), .Z(n2232) );
  NAND U2644 ( .A(B[104]), .B(n2236), .Z(n2235) );
  NANDN U2645 ( .A(A[104]), .B(n2237), .Z(n2236) );
  NANDN U2646 ( .A(n2237), .B(A[104]), .Z(n2234) );
  XOR U2647 ( .A(n2237), .B(n2238), .Z(SUM[104]) );
  XNOR U2648 ( .A(B[104]), .B(A[104]), .Z(n2238) );
  AND U2649 ( .A(n2239), .B(n2240), .Z(n2237) );
  NAND U2650 ( .A(B[103]), .B(n2241), .Z(n2240) );
  NANDN U2651 ( .A(A[103]), .B(n2242), .Z(n2241) );
  NANDN U2652 ( .A(n2242), .B(A[103]), .Z(n2239) );
  XOR U2653 ( .A(n2242), .B(n2243), .Z(SUM[103]) );
  XNOR U2654 ( .A(B[103]), .B(A[103]), .Z(n2243) );
  AND U2655 ( .A(n2244), .B(n2245), .Z(n2242) );
  NAND U2656 ( .A(B[102]), .B(n2246), .Z(n2245) );
  NANDN U2657 ( .A(A[102]), .B(n2247), .Z(n2246) );
  NANDN U2658 ( .A(n2247), .B(A[102]), .Z(n2244) );
  XOR U2659 ( .A(n2247), .B(n2248), .Z(SUM[102]) );
  XNOR U2660 ( .A(B[102]), .B(A[102]), .Z(n2248) );
  AND U2661 ( .A(n2249), .B(n2250), .Z(n2247) );
  NAND U2662 ( .A(B[101]), .B(n2251), .Z(n2250) );
  NANDN U2663 ( .A(A[101]), .B(n2252), .Z(n2251) );
  NANDN U2664 ( .A(n2252), .B(A[101]), .Z(n2249) );
  XOR U2665 ( .A(n2252), .B(n2253), .Z(SUM[101]) );
  XNOR U2666 ( .A(B[101]), .B(A[101]), .Z(n2253) );
  AND U2667 ( .A(n2254), .B(n2255), .Z(n2252) );
  NAND U2668 ( .A(B[100]), .B(n2256), .Z(n2255) );
  NANDN U2669 ( .A(A[100]), .B(n2257), .Z(n2256) );
  NANDN U2670 ( .A(n2257), .B(A[100]), .Z(n2254) );
  XOR U2671 ( .A(n2257), .B(n2258), .Z(SUM[100]) );
  XNOR U2672 ( .A(B[100]), .B(A[100]), .Z(n2258) );
  AND U2673 ( .A(n2259), .B(n2260), .Z(n2257) );
  NAND U2674 ( .A(B[99]), .B(n2261), .Z(n2260) );
  OR U2675 ( .A(n3), .B(A[99]), .Z(n2261) );
  NAND U2676 ( .A(A[99]), .B(n3), .Z(n2259) );
  NAND U2677 ( .A(n2262), .B(n2263), .Z(n3) );
  NAND U2678 ( .A(B[98]), .B(n2264), .Z(n2263) );
  NANDN U2679 ( .A(A[98]), .B(n5), .Z(n2264) );
  NANDN U2680 ( .A(n5), .B(A[98]), .Z(n2262) );
  AND U2681 ( .A(n2265), .B(n2266), .Z(n5) );
  NAND U2682 ( .A(B[97]), .B(n2267), .Z(n2266) );
  NANDN U2683 ( .A(A[97]), .B(n7), .Z(n2267) );
  NANDN U2684 ( .A(n7), .B(A[97]), .Z(n2265) );
  AND U2685 ( .A(n2268), .B(n2269), .Z(n7) );
  NAND U2686 ( .A(B[96]), .B(n2270), .Z(n2269) );
  NANDN U2687 ( .A(A[96]), .B(n9), .Z(n2270) );
  NANDN U2688 ( .A(n9), .B(A[96]), .Z(n2268) );
  AND U2689 ( .A(n2271), .B(n2272), .Z(n9) );
  NAND U2690 ( .A(B[95]), .B(n2273), .Z(n2272) );
  NANDN U2691 ( .A(A[95]), .B(n11), .Z(n2273) );
  NANDN U2692 ( .A(n11), .B(A[95]), .Z(n2271) );
  AND U2693 ( .A(n2274), .B(n2275), .Z(n11) );
  NAND U2694 ( .A(B[94]), .B(n2276), .Z(n2275) );
  NANDN U2695 ( .A(A[94]), .B(n13), .Z(n2276) );
  NANDN U2696 ( .A(n13), .B(A[94]), .Z(n2274) );
  AND U2697 ( .A(n2277), .B(n2278), .Z(n13) );
  NAND U2698 ( .A(B[93]), .B(n2279), .Z(n2278) );
  NANDN U2699 ( .A(A[93]), .B(n15), .Z(n2279) );
  NANDN U2700 ( .A(n15), .B(A[93]), .Z(n2277) );
  AND U2701 ( .A(n2280), .B(n2281), .Z(n15) );
  NAND U2702 ( .A(B[92]), .B(n2282), .Z(n2281) );
  NANDN U2703 ( .A(A[92]), .B(n17), .Z(n2282) );
  NANDN U2704 ( .A(n17), .B(A[92]), .Z(n2280) );
  AND U2705 ( .A(n2283), .B(n2284), .Z(n17) );
  NAND U2706 ( .A(B[91]), .B(n2285), .Z(n2284) );
  NANDN U2707 ( .A(A[91]), .B(n19), .Z(n2285) );
  NANDN U2708 ( .A(n19), .B(A[91]), .Z(n2283) );
  AND U2709 ( .A(n2286), .B(n2287), .Z(n19) );
  NAND U2710 ( .A(B[90]), .B(n2288), .Z(n2287) );
  NANDN U2711 ( .A(A[90]), .B(n21), .Z(n2288) );
  NANDN U2712 ( .A(n21), .B(A[90]), .Z(n2286) );
  AND U2713 ( .A(n2289), .B(n2290), .Z(n21) );
  NAND U2714 ( .A(B[89]), .B(n2291), .Z(n2290) );
  NANDN U2715 ( .A(A[89]), .B(n25), .Z(n2291) );
  NANDN U2716 ( .A(n25), .B(A[89]), .Z(n2289) );
  AND U2717 ( .A(n2292), .B(n2293), .Z(n25) );
  NAND U2718 ( .A(B[88]), .B(n2294), .Z(n2293) );
  NANDN U2719 ( .A(A[88]), .B(n27), .Z(n2294) );
  NANDN U2720 ( .A(n27), .B(A[88]), .Z(n2292) );
  AND U2721 ( .A(n2295), .B(n2296), .Z(n27) );
  NAND U2722 ( .A(B[87]), .B(n2297), .Z(n2296) );
  NANDN U2723 ( .A(A[87]), .B(n29), .Z(n2297) );
  NANDN U2724 ( .A(n29), .B(A[87]), .Z(n2295) );
  AND U2725 ( .A(n2298), .B(n2299), .Z(n29) );
  NAND U2726 ( .A(B[86]), .B(n2300), .Z(n2299) );
  NANDN U2727 ( .A(A[86]), .B(n31), .Z(n2300) );
  NANDN U2728 ( .A(n31), .B(A[86]), .Z(n2298) );
  AND U2729 ( .A(n2301), .B(n2302), .Z(n31) );
  NAND U2730 ( .A(B[85]), .B(n2303), .Z(n2302) );
  NANDN U2731 ( .A(A[85]), .B(n33), .Z(n2303) );
  NANDN U2732 ( .A(n33), .B(A[85]), .Z(n2301) );
  AND U2733 ( .A(n2304), .B(n2305), .Z(n33) );
  NAND U2734 ( .A(B[84]), .B(n2306), .Z(n2305) );
  NANDN U2735 ( .A(A[84]), .B(n35), .Z(n2306) );
  NANDN U2736 ( .A(n35), .B(A[84]), .Z(n2304) );
  AND U2737 ( .A(n2307), .B(n2308), .Z(n35) );
  NAND U2738 ( .A(B[83]), .B(n2309), .Z(n2308) );
  NANDN U2739 ( .A(A[83]), .B(n37), .Z(n2309) );
  NANDN U2740 ( .A(n37), .B(A[83]), .Z(n2307) );
  AND U2741 ( .A(n2310), .B(n2311), .Z(n37) );
  NAND U2742 ( .A(B[82]), .B(n2312), .Z(n2311) );
  NANDN U2743 ( .A(A[82]), .B(n39), .Z(n2312) );
  NANDN U2744 ( .A(n39), .B(A[82]), .Z(n2310) );
  AND U2745 ( .A(n2313), .B(n2314), .Z(n39) );
  NAND U2746 ( .A(B[81]), .B(n2315), .Z(n2314) );
  NANDN U2747 ( .A(A[81]), .B(n41), .Z(n2315) );
  NANDN U2748 ( .A(n41), .B(A[81]), .Z(n2313) );
  AND U2749 ( .A(n2316), .B(n2317), .Z(n41) );
  NAND U2750 ( .A(B[80]), .B(n2318), .Z(n2317) );
  NANDN U2751 ( .A(A[80]), .B(n43), .Z(n2318) );
  NANDN U2752 ( .A(n43), .B(A[80]), .Z(n2316) );
  AND U2753 ( .A(n2319), .B(n2320), .Z(n43) );
  NAND U2754 ( .A(B[79]), .B(n2321), .Z(n2320) );
  NANDN U2755 ( .A(A[79]), .B(n47), .Z(n2321) );
  NANDN U2756 ( .A(n47), .B(A[79]), .Z(n2319) );
  AND U2757 ( .A(n2322), .B(n2323), .Z(n47) );
  NAND U2758 ( .A(B[78]), .B(n2324), .Z(n2323) );
  NANDN U2759 ( .A(A[78]), .B(n49), .Z(n2324) );
  NANDN U2760 ( .A(n49), .B(A[78]), .Z(n2322) );
  AND U2761 ( .A(n2325), .B(n2326), .Z(n49) );
  NAND U2762 ( .A(B[77]), .B(n2327), .Z(n2326) );
  NANDN U2763 ( .A(A[77]), .B(n51), .Z(n2327) );
  NANDN U2764 ( .A(n51), .B(A[77]), .Z(n2325) );
  AND U2765 ( .A(n2328), .B(n2329), .Z(n51) );
  NAND U2766 ( .A(B[76]), .B(n2330), .Z(n2329) );
  NANDN U2767 ( .A(A[76]), .B(n53), .Z(n2330) );
  NANDN U2768 ( .A(n53), .B(A[76]), .Z(n2328) );
  AND U2769 ( .A(n2331), .B(n2332), .Z(n53) );
  NAND U2770 ( .A(B[75]), .B(n2333), .Z(n2332) );
  NANDN U2771 ( .A(A[75]), .B(n55), .Z(n2333) );
  NANDN U2772 ( .A(n55), .B(A[75]), .Z(n2331) );
  AND U2773 ( .A(n2334), .B(n2335), .Z(n55) );
  NAND U2774 ( .A(B[74]), .B(n2336), .Z(n2335) );
  NANDN U2775 ( .A(A[74]), .B(n57), .Z(n2336) );
  NANDN U2776 ( .A(n57), .B(A[74]), .Z(n2334) );
  AND U2777 ( .A(n2337), .B(n2338), .Z(n57) );
  NAND U2778 ( .A(B[73]), .B(n2339), .Z(n2338) );
  NANDN U2779 ( .A(A[73]), .B(n59), .Z(n2339) );
  NANDN U2780 ( .A(n59), .B(A[73]), .Z(n2337) );
  AND U2781 ( .A(n2340), .B(n2341), .Z(n59) );
  NAND U2782 ( .A(B[72]), .B(n2342), .Z(n2341) );
  NANDN U2783 ( .A(A[72]), .B(n61), .Z(n2342) );
  NANDN U2784 ( .A(n61), .B(A[72]), .Z(n2340) );
  AND U2785 ( .A(n2343), .B(n2344), .Z(n61) );
  NAND U2786 ( .A(B[71]), .B(n2345), .Z(n2344) );
  NANDN U2787 ( .A(A[71]), .B(n63), .Z(n2345) );
  NANDN U2788 ( .A(n63), .B(A[71]), .Z(n2343) );
  AND U2789 ( .A(n2346), .B(n2347), .Z(n63) );
  NAND U2790 ( .A(B[70]), .B(n2348), .Z(n2347) );
  NANDN U2791 ( .A(A[70]), .B(n65), .Z(n2348) );
  NANDN U2792 ( .A(n65), .B(A[70]), .Z(n2346) );
  AND U2793 ( .A(n2349), .B(n2350), .Z(n65) );
  NAND U2794 ( .A(B[69]), .B(n2351), .Z(n2350) );
  NANDN U2795 ( .A(A[69]), .B(n69), .Z(n2351) );
  NANDN U2796 ( .A(n69), .B(A[69]), .Z(n2349) );
  AND U2797 ( .A(n2352), .B(n2353), .Z(n69) );
  NAND U2798 ( .A(B[68]), .B(n2354), .Z(n2353) );
  NANDN U2799 ( .A(A[68]), .B(n71), .Z(n2354) );
  NANDN U2800 ( .A(n71), .B(A[68]), .Z(n2352) );
  AND U2801 ( .A(n2355), .B(n2356), .Z(n71) );
  NAND U2802 ( .A(B[67]), .B(n2357), .Z(n2356) );
  NANDN U2803 ( .A(A[67]), .B(n73), .Z(n2357) );
  NANDN U2804 ( .A(n73), .B(A[67]), .Z(n2355) );
  AND U2805 ( .A(n2358), .B(n2359), .Z(n73) );
  NAND U2806 ( .A(B[66]), .B(n2360), .Z(n2359) );
  NANDN U2807 ( .A(A[66]), .B(n75), .Z(n2360) );
  NANDN U2808 ( .A(n75), .B(A[66]), .Z(n2358) );
  AND U2809 ( .A(n2361), .B(n2362), .Z(n75) );
  NAND U2810 ( .A(B[65]), .B(n2363), .Z(n2362) );
  NANDN U2811 ( .A(A[65]), .B(n77), .Z(n2363) );
  NANDN U2812 ( .A(n77), .B(A[65]), .Z(n2361) );
  AND U2813 ( .A(n2364), .B(n2365), .Z(n77) );
  NAND U2814 ( .A(B[64]), .B(n2366), .Z(n2365) );
  NANDN U2815 ( .A(A[64]), .B(n79), .Z(n2366) );
  NANDN U2816 ( .A(n79), .B(A[64]), .Z(n2364) );
  AND U2817 ( .A(n2367), .B(n2368), .Z(n79) );
  NAND U2818 ( .A(B[63]), .B(n2369), .Z(n2368) );
  NANDN U2819 ( .A(A[63]), .B(n81), .Z(n2369) );
  NANDN U2820 ( .A(n81), .B(A[63]), .Z(n2367) );
  AND U2821 ( .A(n2370), .B(n2371), .Z(n81) );
  NAND U2822 ( .A(B[62]), .B(n2372), .Z(n2371) );
  NANDN U2823 ( .A(A[62]), .B(n83), .Z(n2372) );
  NANDN U2824 ( .A(n83), .B(A[62]), .Z(n2370) );
  AND U2825 ( .A(n2373), .B(n2374), .Z(n83) );
  NAND U2826 ( .A(B[61]), .B(n2375), .Z(n2374) );
  NANDN U2827 ( .A(A[61]), .B(n85), .Z(n2375) );
  NANDN U2828 ( .A(n85), .B(A[61]), .Z(n2373) );
  AND U2829 ( .A(n2376), .B(n2377), .Z(n85) );
  NAND U2830 ( .A(B[60]), .B(n2378), .Z(n2377) );
  NANDN U2831 ( .A(A[60]), .B(n87), .Z(n2378) );
  NANDN U2832 ( .A(n87), .B(A[60]), .Z(n2376) );
  AND U2833 ( .A(n2379), .B(n2380), .Z(n87) );
  NAND U2834 ( .A(B[59]), .B(n2381), .Z(n2380) );
  NANDN U2835 ( .A(A[59]), .B(n91), .Z(n2381) );
  NANDN U2836 ( .A(n91), .B(A[59]), .Z(n2379) );
  AND U2837 ( .A(n2382), .B(n2383), .Z(n91) );
  NAND U2838 ( .A(B[58]), .B(n2384), .Z(n2383) );
  NANDN U2839 ( .A(A[58]), .B(n93), .Z(n2384) );
  NANDN U2840 ( .A(n93), .B(A[58]), .Z(n2382) );
  AND U2841 ( .A(n2385), .B(n2386), .Z(n93) );
  NAND U2842 ( .A(B[57]), .B(n2387), .Z(n2386) );
  NANDN U2843 ( .A(A[57]), .B(n95), .Z(n2387) );
  NANDN U2844 ( .A(n95), .B(A[57]), .Z(n2385) );
  AND U2845 ( .A(n2388), .B(n2389), .Z(n95) );
  NAND U2846 ( .A(B[56]), .B(n2390), .Z(n2389) );
  NANDN U2847 ( .A(A[56]), .B(n97), .Z(n2390) );
  NANDN U2848 ( .A(n97), .B(A[56]), .Z(n2388) );
  AND U2849 ( .A(n2391), .B(n2392), .Z(n97) );
  NAND U2850 ( .A(B[55]), .B(n2393), .Z(n2392) );
  NANDN U2851 ( .A(A[55]), .B(n99), .Z(n2393) );
  NANDN U2852 ( .A(n99), .B(A[55]), .Z(n2391) );
  AND U2853 ( .A(n2394), .B(n2395), .Z(n99) );
  NAND U2854 ( .A(B[54]), .B(n2396), .Z(n2395) );
  NANDN U2855 ( .A(A[54]), .B(n101), .Z(n2396) );
  NANDN U2856 ( .A(n101), .B(A[54]), .Z(n2394) );
  AND U2857 ( .A(n2397), .B(n2398), .Z(n101) );
  NAND U2858 ( .A(B[53]), .B(n2399), .Z(n2398) );
  NANDN U2859 ( .A(A[53]), .B(n103), .Z(n2399) );
  NANDN U2860 ( .A(n103), .B(A[53]), .Z(n2397) );
  AND U2861 ( .A(n2400), .B(n2401), .Z(n103) );
  NAND U2862 ( .A(B[52]), .B(n2402), .Z(n2401) );
  NANDN U2863 ( .A(A[52]), .B(n105), .Z(n2402) );
  NANDN U2864 ( .A(n105), .B(A[52]), .Z(n2400) );
  AND U2865 ( .A(n2403), .B(n2404), .Z(n105) );
  NAND U2866 ( .A(B[51]), .B(n2405), .Z(n2404) );
  NANDN U2867 ( .A(A[51]), .B(n107), .Z(n2405) );
  NANDN U2868 ( .A(n107), .B(A[51]), .Z(n2403) );
  AND U2869 ( .A(n2406), .B(n2407), .Z(n107) );
  NAND U2870 ( .A(B[50]), .B(n2408), .Z(n2407) );
  NANDN U2871 ( .A(A[50]), .B(n125), .Z(n2408) );
  NANDN U2872 ( .A(n125), .B(A[50]), .Z(n2406) );
  AND U2873 ( .A(n2409), .B(n2410), .Z(n125) );
  NAND U2874 ( .A(B[49]), .B(n2411), .Z(n2410) );
  NANDN U2875 ( .A(A[49]), .B(n179), .Z(n2411) );
  NANDN U2876 ( .A(n179), .B(A[49]), .Z(n2409) );
  AND U2877 ( .A(n2412), .B(n2413), .Z(n179) );
  NAND U2878 ( .A(B[48]), .B(n2414), .Z(n2413) );
  NANDN U2879 ( .A(A[48]), .B(n231), .Z(n2414) );
  NANDN U2880 ( .A(n231), .B(A[48]), .Z(n2412) );
  AND U2881 ( .A(n2415), .B(n2416), .Z(n231) );
  NAND U2882 ( .A(B[47]), .B(n2417), .Z(n2416) );
  NANDN U2883 ( .A(A[47]), .B(n283), .Z(n2417) );
  NANDN U2884 ( .A(n283), .B(A[47]), .Z(n2415) );
  AND U2885 ( .A(n2418), .B(n2419), .Z(n283) );
  NAND U2886 ( .A(B[46]), .B(n2420), .Z(n2419) );
  NANDN U2887 ( .A(A[46]), .B(n335), .Z(n2420) );
  NANDN U2888 ( .A(n335), .B(A[46]), .Z(n2418) );
  AND U2889 ( .A(n2421), .B(n2422), .Z(n335) );
  NAND U2890 ( .A(B[45]), .B(n2423), .Z(n2422) );
  NANDN U2891 ( .A(A[45]), .B(n387), .Z(n2423) );
  NANDN U2892 ( .A(n387), .B(A[45]), .Z(n2421) );
  AND U2893 ( .A(n2424), .B(n2425), .Z(n387) );
  NAND U2894 ( .A(B[44]), .B(n2426), .Z(n2425) );
  NANDN U2895 ( .A(A[44]), .B(n439), .Z(n2426) );
  NANDN U2896 ( .A(n439), .B(A[44]), .Z(n2424) );
  AND U2897 ( .A(n2427), .B(n2428), .Z(n439) );
  NAND U2898 ( .A(B[43]), .B(n2429), .Z(n2428) );
  NANDN U2899 ( .A(A[43]), .B(n491), .Z(n2429) );
  NANDN U2900 ( .A(n491), .B(A[43]), .Z(n2427) );
  AND U2901 ( .A(n2430), .B(n2431), .Z(n491) );
  NAND U2902 ( .A(B[42]), .B(n2432), .Z(n2431) );
  NANDN U2903 ( .A(A[42]), .B(n543), .Z(n2432) );
  NANDN U2904 ( .A(n543), .B(A[42]), .Z(n2430) );
  AND U2905 ( .A(n2433), .B(n2434), .Z(n543) );
  NAND U2906 ( .A(B[41]), .B(n2435), .Z(n2434) );
  NANDN U2907 ( .A(A[41]), .B(n595), .Z(n2435) );
  NANDN U2908 ( .A(n595), .B(A[41]), .Z(n2433) );
  AND U2909 ( .A(n2436), .B(n2437), .Z(n595) );
  NAND U2910 ( .A(B[40]), .B(n2438), .Z(n2437) );
  NANDN U2911 ( .A(A[40]), .B(n647), .Z(n2438) );
  NANDN U2912 ( .A(n647), .B(A[40]), .Z(n2436) );
  AND U2913 ( .A(n2439), .B(n2440), .Z(n647) );
  NAND U2914 ( .A(B[39]), .B(n2441), .Z(n2440) );
  NANDN U2915 ( .A(A[39]), .B(n701), .Z(n2441) );
  NANDN U2916 ( .A(n701), .B(A[39]), .Z(n2439) );
  AND U2917 ( .A(n2442), .B(n2443), .Z(n701) );
  NAND U2918 ( .A(B[38]), .B(n2444), .Z(n2443) );
  NANDN U2919 ( .A(A[38]), .B(n753), .Z(n2444) );
  NANDN U2920 ( .A(n753), .B(A[38]), .Z(n2442) );
  AND U2921 ( .A(n2445), .B(n2446), .Z(n753) );
  NAND U2922 ( .A(B[37]), .B(n2447), .Z(n2446) );
  NANDN U2923 ( .A(A[37]), .B(n805), .Z(n2447) );
  NANDN U2924 ( .A(n805), .B(A[37]), .Z(n2445) );
  AND U2925 ( .A(n2448), .B(n2449), .Z(n805) );
  NAND U2926 ( .A(B[36]), .B(n2450), .Z(n2449) );
  NANDN U2927 ( .A(A[36]), .B(n857), .Z(n2450) );
  NANDN U2928 ( .A(n857), .B(A[36]), .Z(n2448) );
  AND U2929 ( .A(n2451), .B(n2452), .Z(n857) );
  NAND U2930 ( .A(B[35]), .B(n2453), .Z(n2452) );
  NANDN U2931 ( .A(A[35]), .B(n909), .Z(n2453) );
  NANDN U2932 ( .A(n909), .B(A[35]), .Z(n2451) );
  AND U2933 ( .A(n2454), .B(n2455), .Z(n909) );
  NAND U2934 ( .A(B[34]), .B(n2456), .Z(n2455) );
  NANDN U2935 ( .A(A[34]), .B(n961), .Z(n2456) );
  NANDN U2936 ( .A(n961), .B(A[34]), .Z(n2454) );
  AND U2937 ( .A(n2457), .B(n2458), .Z(n961) );
  NAND U2938 ( .A(B[33]), .B(n2459), .Z(n2458) );
  NANDN U2939 ( .A(A[33]), .B(n1013), .Z(n2459) );
  NANDN U2940 ( .A(n1013), .B(A[33]), .Z(n2457) );
  AND U2941 ( .A(n2460), .B(n2461), .Z(n1013) );
  NAND U2942 ( .A(B[32]), .B(n2462), .Z(n2461) );
  NANDN U2943 ( .A(A[32]), .B(n1065), .Z(n2462) );
  NANDN U2944 ( .A(n1065), .B(A[32]), .Z(n2460) );
  AND U2945 ( .A(n2463), .B(n2464), .Z(n1065) );
  NAND U2946 ( .A(B[31]), .B(n2465), .Z(n2464) );
  NANDN U2947 ( .A(A[31]), .B(n1117), .Z(n2465) );
  NANDN U2948 ( .A(n1117), .B(A[31]), .Z(n2463) );
  AND U2949 ( .A(n2466), .B(n2467), .Z(n1117) );
  NAND U2950 ( .A(B[30]), .B(n2468), .Z(n2467) );
  NANDN U2951 ( .A(A[30]), .B(n1169), .Z(n2468) );
  NANDN U2952 ( .A(n1169), .B(A[30]), .Z(n2466) );
  AND U2953 ( .A(n2469), .B(n2470), .Z(n1169) );
  NAND U2954 ( .A(B[29]), .B(n2471), .Z(n2470) );
  NANDN U2955 ( .A(A[29]), .B(n1223), .Z(n2471) );
  NANDN U2956 ( .A(n1223), .B(A[29]), .Z(n2469) );
  AND U2957 ( .A(n2472), .B(n2473), .Z(n1223) );
  NAND U2958 ( .A(B[28]), .B(n2474), .Z(n2473) );
  NANDN U2959 ( .A(A[28]), .B(n1275), .Z(n2474) );
  NANDN U2960 ( .A(n1275), .B(A[28]), .Z(n2472) );
  AND U2961 ( .A(n2475), .B(n2476), .Z(n1275) );
  NAND U2962 ( .A(B[27]), .B(n2477), .Z(n2476) );
  NANDN U2963 ( .A(A[27]), .B(n1327), .Z(n2477) );
  NANDN U2964 ( .A(n1327), .B(A[27]), .Z(n2475) );
  AND U2965 ( .A(n2478), .B(n2479), .Z(n1327) );
  NAND U2966 ( .A(B[26]), .B(n2480), .Z(n2479) );
  NANDN U2967 ( .A(A[26]), .B(n1379), .Z(n2480) );
  NANDN U2968 ( .A(n1379), .B(A[26]), .Z(n2478) );
  AND U2969 ( .A(n2481), .B(n2482), .Z(n1379) );
  NAND U2970 ( .A(B[25]), .B(n2483), .Z(n2482) );
  NANDN U2971 ( .A(A[25]), .B(n1431), .Z(n2483) );
  NANDN U2972 ( .A(n1431), .B(A[25]), .Z(n2481) );
  AND U2973 ( .A(n2484), .B(n2485), .Z(n1431) );
  NAND U2974 ( .A(B[24]), .B(n2486), .Z(n2485) );
  NANDN U2975 ( .A(A[24]), .B(n1483), .Z(n2486) );
  NANDN U2976 ( .A(n1483), .B(A[24]), .Z(n2484) );
  AND U2977 ( .A(n2487), .B(n2488), .Z(n1483) );
  NAND U2978 ( .A(B[23]), .B(n2489), .Z(n2488) );
  NANDN U2979 ( .A(A[23]), .B(n1535), .Z(n2489) );
  NANDN U2980 ( .A(n1535), .B(A[23]), .Z(n2487) );
  AND U2981 ( .A(n2490), .B(n2491), .Z(n1535) );
  NAND U2982 ( .A(B[22]), .B(n2492), .Z(n2491) );
  NANDN U2983 ( .A(A[22]), .B(n1587), .Z(n2492) );
  NANDN U2984 ( .A(n1587), .B(A[22]), .Z(n2490) );
  AND U2985 ( .A(n2493), .B(n2494), .Z(n1587) );
  NAND U2986 ( .A(B[21]), .B(n2495), .Z(n2494) );
  NANDN U2987 ( .A(A[21]), .B(n1639), .Z(n2495) );
  NANDN U2988 ( .A(n1639), .B(A[21]), .Z(n2493) );
  AND U2989 ( .A(n2496), .B(n2497), .Z(n1639) );
  NAND U2990 ( .A(B[20]), .B(n2498), .Z(n2497) );
  NANDN U2991 ( .A(A[20]), .B(n1691), .Z(n2498) );
  NANDN U2992 ( .A(n1691), .B(A[20]), .Z(n2496) );
  AND U2993 ( .A(n2499), .B(n2500), .Z(n1691) );
  NAND U2994 ( .A(B[19]), .B(n2501), .Z(n2500) );
  NANDN U2995 ( .A(A[19]), .B(n1743), .Z(n2501) );
  NANDN U2996 ( .A(n1743), .B(A[19]), .Z(n2499) );
  AND U2997 ( .A(n2502), .B(n2503), .Z(n1743) );
  NAND U2998 ( .A(B[18]), .B(n2504), .Z(n2503) );
  NANDN U2999 ( .A(A[18]), .B(n1795), .Z(n2504) );
  NANDN U3000 ( .A(n1795), .B(A[18]), .Z(n2502) );
  AND U3001 ( .A(n2505), .B(n2506), .Z(n1795) );
  NAND U3002 ( .A(B[17]), .B(n2507), .Z(n2506) );
  NANDN U3003 ( .A(A[17]), .B(n1847), .Z(n2507) );
  NANDN U3004 ( .A(n1847), .B(A[17]), .Z(n2505) );
  AND U3005 ( .A(n2508), .B(n2509), .Z(n1847) );
  NAND U3006 ( .A(B[16]), .B(n2510), .Z(n2509) );
  NANDN U3007 ( .A(A[16]), .B(n1899), .Z(n2510) );
  NANDN U3008 ( .A(n1899), .B(A[16]), .Z(n2508) );
  AND U3009 ( .A(n2511), .B(n2512), .Z(n1899) );
  NAND U3010 ( .A(B[15]), .B(n2513), .Z(n2512) );
  NANDN U3011 ( .A(A[15]), .B(n1951), .Z(n2513) );
  NANDN U3012 ( .A(n1951), .B(A[15]), .Z(n2511) );
  AND U3013 ( .A(n2514), .B(n2515), .Z(n1951) );
  NAND U3014 ( .A(B[14]), .B(n2516), .Z(n2515) );
  NANDN U3015 ( .A(A[14]), .B(n2003), .Z(n2516) );
  NANDN U3016 ( .A(n2003), .B(A[14]), .Z(n2514) );
  AND U3017 ( .A(n2517), .B(n2518), .Z(n2003) );
  NAND U3018 ( .A(B[13]), .B(n2519), .Z(n2518) );
  NANDN U3019 ( .A(A[13]), .B(n2055), .Z(n2519) );
  NANDN U3020 ( .A(n2055), .B(A[13]), .Z(n2517) );
  AND U3021 ( .A(n2520), .B(n2521), .Z(n2055) );
  NAND U3022 ( .A(B[12]), .B(n2522), .Z(n2521) );
  NANDN U3023 ( .A(A[12]), .B(n2107), .Z(n2522) );
  NANDN U3024 ( .A(n2107), .B(A[12]), .Z(n2520) );
  AND U3025 ( .A(n2523), .B(n2524), .Z(n2107) );
  NAND U3026 ( .A(B[11]), .B(n2525), .Z(n2524) );
  NANDN U3027 ( .A(A[11]), .B(n2159), .Z(n2525) );
  NANDN U3028 ( .A(n2159), .B(A[11]), .Z(n2523) );
  AND U3029 ( .A(n2526), .B(n2527), .Z(n2159) );
  NAND U3030 ( .A(B[10]), .B(n2528), .Z(n2527) );
  NANDN U3031 ( .A(A[10]), .B(n2211), .Z(n2528) );
  NANDN U3032 ( .A(n2211), .B(A[10]), .Z(n2526) );
  AND U3033 ( .A(n2529), .B(n2530), .Z(n2211) );
  NAND U3034 ( .A(B[9]), .B(n2531), .Z(n2530) );
  OR U3035 ( .A(n1), .B(A[9]), .Z(n2531) );
  NAND U3036 ( .A(A[9]), .B(n1), .Z(n2529) );
  NAND U3037 ( .A(n2532), .B(n2533), .Z(n1) );
  NAND U3038 ( .A(B[8]), .B(n2534), .Z(n2533) );
  NANDN U3039 ( .A(A[8]), .B(n23), .Z(n2534) );
  NANDN U3040 ( .A(n23), .B(A[8]), .Z(n2532) );
  AND U3041 ( .A(n2535), .B(n2536), .Z(n23) );
  NAND U3042 ( .A(B[7]), .B(n2537), .Z(n2536) );
  NANDN U3043 ( .A(A[7]), .B(n45), .Z(n2537) );
  NANDN U3044 ( .A(n45), .B(A[7]), .Z(n2535) );
  AND U3045 ( .A(n2538), .B(n2539), .Z(n45) );
  NAND U3046 ( .A(B[6]), .B(n2540), .Z(n2539) );
  NANDN U3047 ( .A(A[6]), .B(n67), .Z(n2540) );
  NANDN U3048 ( .A(n67), .B(A[6]), .Z(n2538) );
  AND U3049 ( .A(n2541), .B(n2542), .Z(n67) );
  NAND U3050 ( .A(B[5]), .B(n2543), .Z(n2542) );
  NANDN U3051 ( .A(A[5]), .B(n89), .Z(n2543) );
  NANDN U3052 ( .A(n89), .B(A[5]), .Z(n2541) );
  AND U3053 ( .A(n2544), .B(n2545), .Z(n89) );
  NAND U3054 ( .A(B[4]), .B(n2546), .Z(n2545) );
  NANDN U3055 ( .A(A[4]), .B(n177), .Z(n2546) );
  NANDN U3056 ( .A(n177), .B(A[4]), .Z(n2544) );
  AND U3057 ( .A(n2547), .B(n2548), .Z(n177) );
  NAND U3058 ( .A(B[3]), .B(n2549), .Z(n2548) );
  NANDN U3059 ( .A(A[3]), .B(n699), .Z(n2549) );
  NANDN U3060 ( .A(n699), .B(A[3]), .Z(n2547) );
  AND U3061 ( .A(n2550), .B(n2551), .Z(n699) );
  NAND U3062 ( .A(B[2]), .B(n2552), .Z(n2551) );
  OR U3063 ( .A(n1221), .B(A[2]), .Z(n2552) );
  NAND U3064 ( .A(A[2]), .B(n1221), .Z(n2550) );
  AND U3065 ( .A(B[1]), .B(A[1]), .Z(n1221) );
endmodule


module modmult_step_N512 ( xregN_1, y, n, zin, zout );
  input [511:0] y;
  input [511:0] n;
  input [513:0] zin;
  output [513:0] zout;
  input xregN_1;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18,
         N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N74,
         N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88,
         N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101,
         N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, N112,
         N113, N114, N115, N116, N117, N118, N119, N120, N121, N122, N123,
         N124, N125, N126, N127, N128, N129, N130, N131, N132, N133, N134,
         N135, N136, N137, N138, N139, N140, N141, N142, N143, N144, N145,
         N146, N147, N148, N149, N150, N151, N152, N153, N154, N155, N156,
         N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167,
         N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178,
         N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189,
         N190, N191, N192, N193, N194, N195, N196, N197, N198, N199, N200,
         N201, N202, N203, N204, N205, N206, N207, N208, N209, N210, N211,
         N212, N213, N214, N215, N216, N217, N218, N219, N220, N221, N222,
         N223, N224, N225, N226, N227, N228, N229, N230, N231, N232, N233,
         N234, N235, N236, N237, N238, N239, N240, N241, N242, N243, N244,
         N245, N246, N247, N248, N249, N250, N251, N252, N253, N254, N255,
         N256, N257, N258, N259, N260, N261, N262, N263, N264, N265, N266,
         N267, N268, N269, N270, N271, N272, N273, N274, N275, N276, N277,
         N278, N279, N280, N281, N282, N283, N284, N285, N286, N287, N288,
         N289, N290, N291, N292, N293, N294, N295, N296, N297, N298, N299,
         N300, N301, N302, N303, N304, N305, N306, N307, N308, N309, N310,
         N311, N312, N313, N314, N315, N316, N317, N318, N319, N320, N321,
         N322, N323, N324, N325, N326, N327, N328, N329, N330, N331, N332,
         N333, N334, N335, N336, N337, N338, N339, N340, N341, N342, N343,
         N344, N345, N346, N347, N348, N349, N350, N351, N352, N353, N354,
         N355, N356, N357, N358, N359, N360, N361, N362, N363, N364, N365,
         N366, N367, N368, N369, N370, N371, N372, N373, N374, N375, N376,
         N377, N378, N379, N380, N381, N382, N383, N384, N385, N386, N387,
         N388, N389, N390, N391, N392, N393, N394, N395, N396, N397, N398,
         N399, N400, N401, N402, N403, N404, N405, N406, N407, N408, N409,
         N410, N411, N412, N413, N414, N415, N416, N417, N418, N419, N420,
         N421, N422, N423, N424, N425, N426, N427, N428, N429, N430, N431,
         N432, N433, N434, N435, N436, N437, N438, N439, N440, N441, N442,
         N443, N444, N445, N446, N447, N448, N449, N450, N451, N452, N453,
         N454, N455, N456, N457, N458, N459, N460, N461, N462, N463, N464,
         N465, N466, N467, N468, N469, N470, N471, N472, N473, N474, N475,
         N476, N477, N478, N479, N480, N481, N482, N483, N484, N485, N486,
         N487, N488, N489, N490, N491, N492, N493, N494, N495, N496, N497,
         N498, N499, N500, N501, N502, N503, N504, N505, N506, N507, N508,
         N509, N510, N511, N512, N513, N514, N515, N516, N517, N518, N520,
         N521, N522, N523, N524, N525, N526, N527, N528, N529, N530, N531,
         N532, N533, N534, N535, N536, N537, N538, N539, N540, N541, N542,
         N543, N544, N545, N546, N547, N548, N549, N550, N551, N552, N553,
         N554, N555, N556, N557, N558, N559, N560, N561, N562, N563, N564,
         N565, N566, N567, N568, N569, N570, N571, N572, N573, N574, N575,
         N576, N577, N578, N579, N580, N581, N582, N583, N584, N585, N586,
         N587, N588, N589, N590, N591, N592, N593, N594, N595, N596, N597,
         N598, N599, N600, N601, N602, N603, N604, N605, N606, N607, N608,
         N609, N610, N611, N612, N613, N614, N615, N616, N617, N618, N619,
         N620, N621, N622, N623, N624, N625, N626, N627, N628, N629, N630,
         N631, N632, N633, N634, N635, N636, N637, N638, N639, N640, N641,
         N642, N643, N644, N645, N646, N647, N648, N649, N650, N651, N652,
         N653, N654, N655, N656, N657, N658, N659, N660, N661, N662, N663,
         N664, N665, N666, N667, N668, N669, N670, N671, N672, N673, N674,
         N675, N676, N677, N678, N679, N680, N681, N682, N683, N684, N685,
         N686, N687, N688, N689, N690, N691, N692, N693, N694, N695, N696,
         N697, N698, N699, N700, N701, N702, N703, N704, N705, N706, N707,
         N708, N709, N710, N711, N712, N713, N714, N715, N716, N717, N718,
         N719, N720, N721, N722, N723, N724, N725, N726, N727, N728, N729,
         N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740,
         N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751,
         N752, N753, N754, N755, N756, N757, N758, N759, N760, N761, N762,
         N763, N764, N765, N766, N767, N768, N769, N770, N771, N772, N773,
         N774, N775, N776, N777, N778, N779, N780, N781, N782, N783, N784,
         N785, N786, N787, N788, N789, N790, N791, N792, N793, N794, N795,
         N796, N797, N798, N799, N800, N801, N802, N803, N804, N805, N806,
         N807, N808, N809, N810, N811, N812, N813, N814, N815, N816, N817,
         N818, N819, N820, N821, N822, N823, N824, N825, N826, N827, N828,
         N829, N830, N831, N832, N833, N834, N835, N836, N837, N838, N839,
         N840, N841, N842, N843, N844, N845, N846, N847, N848, N849, N850,
         N851, N852, N853, N854, N855, N856, N857, N858, N859, N860, N861,
         N862, N863, N864, N865, N866, N867, N868, N869, N870, N871, N872,
         N873, N874, N875, N876, N877, N878, N879, N880, N881, N882, N883,
         N884, N885, N886, N887, N888, N889, N890, N891, N892, N893, N894,
         N895, N896, N897, N898, N899, N900, N901, N902, N903, N904, N905,
         N906, N907, N908, N909, N910, N911, N912, N913, N914, N915, N916,
         N917, N918, N919, N920, N921, N922, N923, N924, N925, N926, N927,
         N928, N929, N930, N931, N932, N933, N934, N935, N936, N937, N938,
         N939, N940, N941, N942, N943, N944, N945, N946, N947, N948, N949,
         N950, N951, N952, N953, N954, N955, N956, N957, N958, N959, N960,
         N961, N962, N963, N964, N965, N966, N967, N968, N969, N970, N971,
         N972, N973, N974, N975, N976, N977, N978, N979, N980, N981, N982,
         N983, N984, N985, N986, N987, N988, N989, N990, N991, N992, N993,
         N994, N995, N996, N997, N998, N999, N1000, N1001, N1002, N1003, N1004,
         N1005, N1006, N1007, N1008, N1009, N1010, N1011, N1012, N1013, N1014,
         N1015, N1016, N1017, N1018, N1019, N1020, N1021, N1022, N1023, N1024,
         N1025, N1026, N1027, N1028, N1029, N1030, N1031, N1032, N1033, N1548,
         N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538,
         N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528,
         N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518,
         N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508,
         N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498,
         N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488,
         N1487, N1486, N1485, N1484, N1483, N1482, N1481, N1480, N1479, N1478,
         N1477, N1476, N1475, N1474, N1473, N1472, N1471, N1470, N1469, N1468,
         N1467, N1466, N1465, N1464, N1463, N1462, N1461, N1460, N1459, N1458,
         N1457, N1456, N1455, N1454, N1453, N1452, N1451, N1450, N1449, N1448,
         N1447, N1446, N1445, N1444, N1443, N1442, N1441, N1440, N1439, N1438,
         N1437, N1436, N1435, N1434, N1433, N1432, N1431, N1430, N1429, N1428,
         N1427, N1426, N1425, N1424, N1423, N1422, N1421, N1420, N1419, N1418,
         N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408,
         N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398,
         N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388,
         N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378,
         N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368,
         N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358,
         N1357, N1356, N1355, N1354, N1353, N1352, N1351, N1350, N1349, N1348,
         N1347, N1346, N1345, N1344, N1343, N1342, N1341, N1340, N1339, N1338,
         N1337, N1336, N1335, N1334, N1333, N1332, N1331, N1330, N1329, N1328,
         N1327, N1326, N1325, N1324, N1323, N1322, N1321, N1320, N1319, N1318,
         N1317, N1316, N1315, N1314, N1313, N1312, N1311, N1310, N1309, N1308,
         N1307, N1306, N1305, N1304, N1303, N1302, N1301, N1300, N1299, N1298,
         N1297, N1296, N1295, N1294, N1293, N1292, N1291, N1290, N1289, N1288,
         N1287, N1286, N1285, N1284, N1283, N1282, N1281, N1280, N1279, N1278,
         N1277, N1276, N1275, N1274, N1273, N1272, N1271, N1270, N1269, N1268,
         N1267, N1266, N1265, N1264, N1263, N1262, N1261, N1260, N1259, N1258,
         N1257, N1256, N1255, N1254, N1253, N1252, N1251, N1250, N1249, N1248,
         N1247, N1246, N1245, N1244, N1243, N1242, N1241, N1240, N1239, N1238,
         N1237, N1236, N1235, N1234, N1233, N1232, N1231, N1230, N1229, N1228,
         N1227, N1226, N1225, N1224, N1223, N1222, N1221, N1220, N1219, N1218,
         N1217, N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208,
         N1207, N1206, N1205, N1204, N1203, N1202, N1201, N1200, N1199, N1198,
         N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190, N1189, N1188,
         N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178,
         N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1169, N1168,
         N1167, N1166, N1165, N1164, N1163, N1162, N1161, N1160, N1159, N1158,
         N1157, N1156, N1155, N1154, N1153, N1152, N1151, N1150, N1149, N1148,
         N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138,
         N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128,
         N1127, N1126, N1125, N1124, N1123, N1122, N1121, N1120, N1119, N1118,
         N1117, N1116, N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108,
         N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099, N1098,
         N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088,
         N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078,
         N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069, N1068,
         N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058,
         N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049, N1048,
         N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038,
         N1037, N1034, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
         n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
         n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
         n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
         n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
         n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
         n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
         n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
         n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
         n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
         n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
         n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
         n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
         n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
         n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
         n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
         n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
         n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
         n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
         n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
         n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
         n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
         n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
         n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
         n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
         n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
         n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
         n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
         n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
         n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
         n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
         n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895,
         n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
         n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
         n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
         n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
         n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
         n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
         n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
         n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
         n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
         n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
         n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
         n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
         n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
         n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
         n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
         n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
         n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063;
  wire   [513:0] z2;
  wire   [513:0] z3;
  wire   SYNOPSYS_UNCONNECTED__0;

  modmult_step_N512_DW01_sub_0 sub_129_aco ( .A(z3), .B({1'b0, 1'b0, N1548, 
        N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, 
        N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, 
        N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, 
        N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, 
        N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, 
        N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, 
        N1487, N1486, N1485, N1484, N1483, N1482, N1481, N1480, N1479, N1478, 
        N1477, N1476, N1475, N1474, N1473, N1472, N1471, N1470, N1469, N1468, 
        N1467, N1466, N1465, N1464, N1463, N1462, N1461, N1460, N1459, N1458, 
        N1457, N1456, N1455, N1454, N1453, N1452, N1451, N1450, N1449, N1448, 
        N1447, N1446, N1445, N1444, N1443, N1442, N1441, N1440, N1439, N1438, 
        N1437, N1436, N1435, N1434, N1433, N1432, N1431, N1430, N1429, N1428, 
        N1427, N1426, N1425, N1424, N1423, N1422, N1421, N1420, N1419, N1418, 
        N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, 
        N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, 
        N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, 
        N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, 
        N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, 
        N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, 
        N1357, N1356, N1355, N1354, N1353, N1352, N1351, N1350, N1349, N1348, 
        N1347, N1346, N1345, N1344, N1343, N1342, N1341, N1340, N1339, N1338, 
        N1337, N1336, N1335, N1334, N1333, N1332, N1331, N1330, N1329, N1328, 
        N1327, N1326, N1325, N1324, N1323, N1322, N1321, N1320, N1319, N1318, 
        N1317, N1316, N1315, N1314, N1313, N1312, N1311, N1310, N1309, N1308, 
        N1307, N1306, N1305, N1304, N1303, N1302, N1301, N1300, N1299, N1298, 
        N1297, N1296, N1295, N1294, N1293, N1292, N1291, N1290, N1289, N1288, 
        N1287, N1286, N1285, N1284, N1283, N1282, N1281, N1280, N1279, N1278, 
        N1277, N1276, N1275, N1274, N1273, N1272, N1271, N1270, N1269, N1268, 
        N1267, N1266, N1265, N1264, N1263, N1262, N1261, N1260, N1259, N1258, 
        N1257, N1256, N1255, N1254, N1253, N1252, N1251, N1250, N1249, N1248, 
        N1247, N1246, N1245, N1244, N1243, N1242, N1241, N1240, N1239, N1238, 
        N1237, N1236, N1235, N1234, N1233, N1232, N1231, N1230, N1229, N1228, 
        N1227, N1226, N1225, N1224, N1223, N1222, N1221, N1220, N1219, N1218, 
        N1217, N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208, 
        N1207, N1206, N1205, N1204, N1203, N1202, N1201, N1200, N1199, N1198, 
        N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190, N1189, N1188, 
        N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178, 
        N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1169, N1168, 
        N1167, N1166, N1165, N1164, N1163, N1162, N1161, N1160, N1159, N1158, 
        N1157, N1156, N1155, N1154, N1153, N1152, N1151, N1150, N1149, N1148, 
        N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, 
        N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, 
        N1127, N1126, N1125, N1124, N1123, N1122, N1121, N1120, N1119, N1118, 
        N1117, N1116, N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, 
        N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099, N1098, 
        N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, 
        N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, 
        N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069, N1068, 
        N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058, 
        N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049, N1048, 
        N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, 
        N1037}), .CI(1'b0), .DIFF(zout) );
  modmult_step_N512_DW02_mult_0 mult_sub_129_aco ( .A(n), .B(N1034), .TC(1'b0), 
        .PRODUCT({SYNOPSYS_UNCONNECTED__0, N1548, N1547, N1546, N1545, N1544, 
        N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, 
        N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, 
        N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, 
        N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, 
        N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, 
        N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486, N1485, N1484, 
        N1483, N1482, N1481, N1480, N1479, N1478, N1477, N1476, N1475, N1474, 
        N1473, N1472, N1471, N1470, N1469, N1468, N1467, N1466, N1465, N1464, 
        N1463, N1462, N1461, N1460, N1459, N1458, N1457, N1456, N1455, N1454, 
        N1453, N1452, N1451, N1450, N1449, N1448, N1447, N1446, N1445, N1444, 
        N1443, N1442, N1441, N1440, N1439, N1438, N1437, N1436, N1435, N1434, 
        N1433, N1432, N1431, N1430, N1429, N1428, N1427, N1426, N1425, N1424, 
        N1423, N1422, N1421, N1420, N1419, N1418, N1417, N1416, N1415, N1414, 
        N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, 
        N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, 
        N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, 
        N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, 
        N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, 
        N1363, N1362, N1361, N1360, N1359, N1358, N1357, N1356, N1355, N1354, 
        N1353, N1352, N1351, N1350, N1349, N1348, N1347, N1346, N1345, N1344, 
        N1343, N1342, N1341, N1340, N1339, N1338, N1337, N1336, N1335, N1334, 
        N1333, N1332, N1331, N1330, N1329, N1328, N1327, N1326, N1325, N1324, 
        N1323, N1322, N1321, N1320, N1319, N1318, N1317, N1316, N1315, N1314, 
        N1313, N1312, N1311, N1310, N1309, N1308, N1307, N1306, N1305, N1304, 
        N1303, N1302, N1301, N1300, N1299, N1298, N1297, N1296, N1295, N1294, 
        N1293, N1292, N1291, N1290, N1289, N1288, N1287, N1286, N1285, N1284, 
        N1283, N1282, N1281, N1280, N1279, N1278, N1277, N1276, N1275, N1274, 
        N1273, N1272, N1271, N1270, N1269, N1268, N1267, N1266, N1265, N1264, 
        N1263, N1262, N1261, N1260, N1259, N1258, N1257, N1256, N1255, N1254, 
        N1253, N1252, N1251, N1250, N1249, N1248, N1247, N1246, N1245, N1244, 
        N1243, N1242, N1241, N1240, N1239, N1238, N1237, N1236, N1235, N1234, 
        N1233, N1232, N1231, N1230, N1229, N1228, N1227, N1226, N1225, N1224, 
        N1223, N1222, N1221, N1220, N1219, N1218, N1217, N1216, N1215, N1214, 
        N1213, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N1205, N1204, 
        N1203, N1202, N1201, N1200, N1199, N1198, N1197, N1196, N1195, N1194, 
        N1193, N1192, N1191, N1190, N1189, N1188, N1187, N1186, N1185, N1184, 
        N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, 
        N1173, N1172, N1171, N1170, N1169, N1168, N1167, N1166, N1165, N1164, 
        N1163, N1162, N1161, N1160, N1159, N1158, N1157, N1156, N1155, N1154, 
        N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, 
        N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, 
        N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126, N1125, N1124, 
        N1123, N1122, N1121, N1120, N1119, N1118, N1117, N1116, N1115, N1114, 
        N1113, N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1105, N1104, 
        N1103, N1102, N1101, N1100, N1099, N1098, N1097, N1096, N1095, N1094, 
        N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, 
        N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, N1075, N1074, 
        N1073, N1072, N1071, N1070, N1069, N1068, N1067, N1066, N1065, N1064, 
        N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, N1054, 
        N1053, N1052, N1051, N1050, N1049, N1048, N1047, N1046, N1045, N1044, 
        N1043, N1042, N1041, N1040, N1039, N1038, N1037}) );
  modmult_step_N512_DW01_cmp2_0 gte_128 ( .A({1'b0, 1'b0, n}), .B(z3), .LEQ(
        1'b1), .TC(1'b0), .LT_LE(N1034) );
  modmult_step_N512_DW01_sub_1 sub_124 ( .A(z2), .B({1'b0, 1'b0, n}), .CI(1'b0), .DIFF({N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, 
        N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, 
        N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, 
        N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, 
        N992, N991, N990, N989, N988, N987, N986, N985, N984, N983, N982, N981, 
        N980, N979, N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, 
        N968, N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, 
        N956, N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, 
        N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, 
        N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922, N921, 
        N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, N909, 
        N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897, 
        N896, N895, N894, N893, N892, N891, N890, N889, N888, N887, N886, N885, 
        N884, N883, N882, N881, N880, N879, N878, N877, N876, N875, N874, N873, 
        N872, N871, N870, N869, N868, N867, N866, N865, N864, N863, N862, N861, 
        N860, N859, N858, N857, N856, N855, N854, N853, N852, N851, N850, N849, 
        N848, N847, N846, N845, N844, N843, N842, N841, N840, N839, N838, N837, 
        N836, N835, N834, N833, N832, N831, N830, N829, N828, N827, N826, N825, 
        N824, N823, N822, N821, N820, N819, N818, N817, N816, N815, N814, N813, 
        N812, N811, N810, N809, N808, N807, N806, N805, N804, N803, N802, N801, 
        N800, N799, N798, N797, N796, N795, N794, N793, N792, N791, N790, N789, 
        N788, N787, N786, N785, N784, N783, N782, N781, N780, N779, N778, N777, 
        N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, 
        N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, 
        N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, 
        N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, 
        N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, 
        N716, N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705, 
        N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694, N693, 
        N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, 
        N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, 
        N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, 
        N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, 
        N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, 
        N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, 
        N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, 
        N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, 
        N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, 
        N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, 
        N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, 
        N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, 
        N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, 
        N536, N535, N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, 
        N524, N523, N522, N521, N520}) );
  modmult_step_N512_DW01_cmp2_1 gt_123 ( .A({1'b0, 1'b0, n}), .B(z2), .LEQ(
        1'b0), .TC(1'b0), .LT_LE(N518) );
  modmult_step_N512_DW01_add_0 add_119 ( .A({zin[512:0], 1'b0}), .B({1'b0, 
        1'b0, y}), .CI(1'b0), .SUM({N517, N516, N515, N514, N513, N512, N511, 
        N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, 
        N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, 
        N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, 
        N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, 
        N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, 
        N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, 
        N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, 
        N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, 
        N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, 
        N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, 
        N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, 
        N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, 
        N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, 
        N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, 
        N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, 
        N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, 
        N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, 
        N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, 
        N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, 
        N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, 
        N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, 
        N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, 
        N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, 
        N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, 
        N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, 
        N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, 
        N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, 
        N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, 
        N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, 
        N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, 
        N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, 
        N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, 
        N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, 
        N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, 
        N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, 
        N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, 
        N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, 
        N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, 
        N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, 
        N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, 
        N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, 
        N4}) );
  NAND U5 ( .A(n1), .B(n2), .Z(z3[9]) );
  NANDN U6 ( .A(N518), .B(z2[9]), .Z(n2) );
  NANDN U7 ( .A(n3), .B(N529), .Z(n1) );
  NAND U8 ( .A(n4), .B(n5), .Z(z3[99]) );
  NANDN U9 ( .A(N518), .B(z2[99]), .Z(n5) );
  NANDN U10 ( .A(n3), .B(N619), .Z(n4) );
  NAND U11 ( .A(n6), .B(n7), .Z(z3[98]) );
  NANDN U17 ( .A(N518), .B(z2[98]), .Z(n7) );
  NANDN U18 ( .A(n3), .B(N618), .Z(n6) );
  NAND U19 ( .A(n8), .B(n9), .Z(z3[97]) );
  NANDN U20 ( .A(N518), .B(z2[97]), .Z(n9) );
  NANDN U21 ( .A(n3), .B(N617), .Z(n8) );
  NAND U22 ( .A(n10), .B(n11), .Z(z3[96]) );
  NANDN U23 ( .A(N518), .B(z2[96]), .Z(n11) );
  NANDN U24 ( .A(n3), .B(N616), .Z(n10) );
  NAND U25 ( .A(n12), .B(n13), .Z(z3[95]) );
  NANDN U26 ( .A(N518), .B(z2[95]), .Z(n13) );
  NANDN U27 ( .A(n3), .B(N615), .Z(n12) );
  NAND U28 ( .A(n14), .B(n23), .Z(z3[94]) );
  NANDN U29 ( .A(N518), .B(z2[94]), .Z(n23) );
  NANDN U30 ( .A(n3), .B(N614), .Z(n14) );
  NAND U31 ( .A(n24), .B(n25), .Z(z3[93]) );
  NANDN U32 ( .A(N518), .B(z2[93]), .Z(n25) );
  NANDN U33 ( .A(n3), .B(N613), .Z(n24) );
  NAND U34 ( .A(n26), .B(n27), .Z(z3[92]) );
  NANDN U35 ( .A(N518), .B(z2[92]), .Z(n27) );
  NANDN U36 ( .A(n3), .B(N612), .Z(n26) );
  NAND U37 ( .A(n28), .B(n29), .Z(z3[91]) );
  NANDN U38 ( .A(N518), .B(z2[91]), .Z(n29) );
  NANDN U39 ( .A(n3), .B(N611), .Z(n28) );
  NAND U40 ( .A(n30), .B(n31), .Z(z3[90]) );
  NANDN U41 ( .A(N518), .B(z2[90]), .Z(n31) );
  NANDN U42 ( .A(n3), .B(N610), .Z(n30) );
  NAND U43 ( .A(n32), .B(n33), .Z(z3[8]) );
  NANDN U44 ( .A(N518), .B(z2[8]), .Z(n33) );
  NANDN U45 ( .A(n3), .B(N528), .Z(n32) );
  NAND U46 ( .A(n34), .B(n35), .Z(z3[89]) );
  NANDN U47 ( .A(N518), .B(z2[89]), .Z(n35) );
  NANDN U48 ( .A(n3), .B(N609), .Z(n34) );
  NAND U49 ( .A(n36), .B(n37), .Z(z3[88]) );
  NANDN U50 ( .A(N518), .B(z2[88]), .Z(n37) );
  NANDN U51 ( .A(n3), .B(N608), .Z(n36) );
  NAND U52 ( .A(n38), .B(n39), .Z(z3[87]) );
  NANDN U53 ( .A(N518), .B(z2[87]), .Z(n39) );
  NANDN U54 ( .A(n3), .B(N607), .Z(n38) );
  NAND U55 ( .A(n40), .B(n41), .Z(z3[86]) );
  NANDN U56 ( .A(N518), .B(z2[86]), .Z(n41) );
  NANDN U57 ( .A(n3), .B(N606), .Z(n40) );
  NAND U58 ( .A(n42), .B(n43), .Z(z3[85]) );
  NANDN U59 ( .A(N518), .B(z2[85]), .Z(n43) );
  NANDN U60 ( .A(n3), .B(N605), .Z(n42) );
  NAND U61 ( .A(n44), .B(n45), .Z(z3[84]) );
  NANDN U62 ( .A(N518), .B(z2[84]), .Z(n45) );
  NANDN U63 ( .A(n3), .B(N604), .Z(n44) );
  NAND U64 ( .A(n46), .B(n47), .Z(z3[83]) );
  NANDN U65 ( .A(N518), .B(z2[83]), .Z(n47) );
  NANDN U66 ( .A(n3), .B(N603), .Z(n46) );
  NAND U67 ( .A(n48), .B(n49), .Z(z3[82]) );
  NANDN U68 ( .A(N518), .B(z2[82]), .Z(n49) );
  NANDN U69 ( .A(n3), .B(N602), .Z(n48) );
  NAND U70 ( .A(n50), .B(n51), .Z(z3[81]) );
  NANDN U71 ( .A(N518), .B(z2[81]), .Z(n51) );
  NANDN U72 ( .A(n3), .B(N601), .Z(n50) );
  NAND U73 ( .A(n52), .B(n53), .Z(z3[80]) );
  NANDN U74 ( .A(N518), .B(z2[80]), .Z(n53) );
  NANDN U75 ( .A(n3), .B(N600), .Z(n52) );
  NAND U76 ( .A(n54), .B(n55), .Z(z3[7]) );
  NANDN U77 ( .A(N518), .B(z2[7]), .Z(n55) );
  NANDN U78 ( .A(n3), .B(N527), .Z(n54) );
  NAND U79 ( .A(n56), .B(n57), .Z(z3[79]) );
  NANDN U80 ( .A(N518), .B(z2[79]), .Z(n57) );
  NANDN U81 ( .A(n3), .B(N599), .Z(n56) );
  NAND U82 ( .A(n58), .B(n59), .Z(z3[78]) );
  NANDN U83 ( .A(N518), .B(z2[78]), .Z(n59) );
  NANDN U84 ( .A(n3), .B(N598), .Z(n58) );
  NAND U85 ( .A(n60), .B(n61), .Z(z3[77]) );
  NANDN U86 ( .A(N518), .B(z2[77]), .Z(n61) );
  NANDN U87 ( .A(n3), .B(N597), .Z(n60) );
  NAND U88 ( .A(n62), .B(n63), .Z(z3[76]) );
  NANDN U89 ( .A(N518), .B(z2[76]), .Z(n63) );
  NANDN U90 ( .A(n3), .B(N596), .Z(n62) );
  NAND U91 ( .A(n64), .B(n65), .Z(z3[75]) );
  NANDN U92 ( .A(N518), .B(z2[75]), .Z(n65) );
  NANDN U93 ( .A(n3), .B(N595), .Z(n64) );
  NAND U94 ( .A(n66), .B(n67), .Z(z3[74]) );
  NANDN U95 ( .A(N518), .B(z2[74]), .Z(n67) );
  NANDN U96 ( .A(n3), .B(N594), .Z(n66) );
  NAND U97 ( .A(n68), .B(n69), .Z(z3[73]) );
  NANDN U98 ( .A(N518), .B(z2[73]), .Z(n69) );
  NANDN U99 ( .A(n3), .B(N593), .Z(n68) );
  NAND U100 ( .A(n70), .B(n71), .Z(z3[72]) );
  NANDN U101 ( .A(N518), .B(z2[72]), .Z(n71) );
  NANDN U102 ( .A(n3), .B(N592), .Z(n70) );
  NAND U103 ( .A(n72), .B(n73), .Z(z3[71]) );
  NANDN U104 ( .A(N518), .B(z2[71]), .Z(n73) );
  NANDN U105 ( .A(n3), .B(N591), .Z(n72) );
  NAND U106 ( .A(n74), .B(n75), .Z(z3[70]) );
  NANDN U107 ( .A(N518), .B(z2[70]), .Z(n75) );
  NANDN U108 ( .A(n3), .B(N590), .Z(n74) );
  NAND U109 ( .A(n76), .B(n77), .Z(z3[6]) );
  NANDN U110 ( .A(N518), .B(z2[6]), .Z(n77) );
  NANDN U111 ( .A(n3), .B(N526), .Z(n76) );
  NAND U112 ( .A(n78), .B(n79), .Z(z3[69]) );
  NANDN U113 ( .A(N518), .B(z2[69]), .Z(n79) );
  NANDN U114 ( .A(n3), .B(N589), .Z(n78) );
  NAND U115 ( .A(n80), .B(n81), .Z(z3[68]) );
  NANDN U116 ( .A(N518), .B(z2[68]), .Z(n81) );
  NANDN U117 ( .A(n3), .B(N588), .Z(n80) );
  NAND U118 ( .A(n82), .B(n83), .Z(z3[67]) );
  NANDN U119 ( .A(N518), .B(z2[67]), .Z(n83) );
  NANDN U120 ( .A(n3), .B(N587), .Z(n82) );
  NAND U121 ( .A(n84), .B(n85), .Z(z3[66]) );
  NANDN U122 ( .A(N518), .B(z2[66]), .Z(n85) );
  NANDN U123 ( .A(n3), .B(N586), .Z(n84) );
  NAND U124 ( .A(n86), .B(n87), .Z(z3[65]) );
  NANDN U125 ( .A(N518), .B(z2[65]), .Z(n87) );
  NANDN U126 ( .A(n3), .B(N585), .Z(n86) );
  NAND U127 ( .A(n88), .B(n89), .Z(z3[64]) );
  NANDN U128 ( .A(N518), .B(z2[64]), .Z(n89) );
  NANDN U129 ( .A(n3), .B(N584), .Z(n88) );
  NAND U130 ( .A(n90), .B(n91), .Z(z3[63]) );
  NANDN U131 ( .A(N518), .B(z2[63]), .Z(n91) );
  NANDN U132 ( .A(n3), .B(N583), .Z(n90) );
  NAND U133 ( .A(n92), .B(n93), .Z(z3[62]) );
  NANDN U134 ( .A(N518), .B(z2[62]), .Z(n93) );
  NANDN U135 ( .A(n3), .B(N582), .Z(n92) );
  NAND U136 ( .A(n94), .B(n95), .Z(z3[61]) );
  NANDN U137 ( .A(N518), .B(z2[61]), .Z(n95) );
  NANDN U138 ( .A(n3), .B(N581), .Z(n94) );
  NAND U139 ( .A(n96), .B(n97), .Z(z3[60]) );
  NANDN U140 ( .A(N518), .B(z2[60]), .Z(n97) );
  NANDN U141 ( .A(n3), .B(N580), .Z(n96) );
  NAND U142 ( .A(n98), .B(n99), .Z(z3[5]) );
  NANDN U143 ( .A(N518), .B(z2[5]), .Z(n99) );
  NANDN U144 ( .A(n3), .B(N525), .Z(n98) );
  NAND U145 ( .A(n100), .B(n101), .Z(z3[59]) );
  NANDN U146 ( .A(N518), .B(z2[59]), .Z(n101) );
  NANDN U147 ( .A(n3), .B(N579), .Z(n100) );
  NAND U148 ( .A(n102), .B(n103), .Z(z3[58]) );
  NANDN U149 ( .A(N518), .B(z2[58]), .Z(n103) );
  NANDN U150 ( .A(n3), .B(N578), .Z(n102) );
  NAND U151 ( .A(n104), .B(n105), .Z(z3[57]) );
  NANDN U152 ( .A(N518), .B(z2[57]), .Z(n105) );
  NANDN U153 ( .A(n3), .B(N577), .Z(n104) );
  NAND U154 ( .A(n106), .B(n107), .Z(z3[56]) );
  NANDN U155 ( .A(N518), .B(z2[56]), .Z(n107) );
  NANDN U156 ( .A(n3), .B(N576), .Z(n106) );
  NAND U157 ( .A(n108), .B(n109), .Z(z3[55]) );
  NANDN U158 ( .A(N518), .B(z2[55]), .Z(n109) );
  NANDN U159 ( .A(n3), .B(N575), .Z(n108) );
  NAND U160 ( .A(n110), .B(n111), .Z(z3[54]) );
  NANDN U161 ( .A(N518), .B(z2[54]), .Z(n111) );
  NANDN U162 ( .A(n3), .B(N574), .Z(n110) );
  NAND U163 ( .A(n112), .B(n113), .Z(z3[53]) );
  NANDN U164 ( .A(N518), .B(z2[53]), .Z(n113) );
  NANDN U165 ( .A(n3), .B(N573), .Z(n112) );
  NAND U166 ( .A(n114), .B(n115), .Z(z3[52]) );
  NANDN U167 ( .A(N518), .B(z2[52]), .Z(n115) );
  NANDN U168 ( .A(n3), .B(N572), .Z(n114) );
  NAND U169 ( .A(n116), .B(n117), .Z(z3[51]) );
  NANDN U170 ( .A(N518), .B(z2[51]), .Z(n117) );
  NANDN U171 ( .A(n3), .B(N571), .Z(n116) );
  NAND U172 ( .A(n118), .B(n119), .Z(z3[513]) );
  NANDN U173 ( .A(N518), .B(z2[513]), .Z(n119) );
  NANDN U174 ( .A(n3), .B(N1033), .Z(n118) );
  NAND U175 ( .A(n120), .B(n121), .Z(z3[512]) );
  NANDN U176 ( .A(N518), .B(z2[512]), .Z(n121) );
  NANDN U177 ( .A(n3), .B(N1032), .Z(n120) );
  NAND U178 ( .A(n122), .B(n123), .Z(z3[511]) );
  NANDN U179 ( .A(N518), .B(z2[511]), .Z(n123) );
  NANDN U180 ( .A(n3), .B(N1031), .Z(n122) );
  NAND U181 ( .A(n124), .B(n125), .Z(z3[510]) );
  NANDN U182 ( .A(N518), .B(z2[510]), .Z(n125) );
  NANDN U183 ( .A(n3), .B(N1030), .Z(n124) );
  NAND U184 ( .A(n126), .B(n127), .Z(z3[50]) );
  NANDN U185 ( .A(N518), .B(z2[50]), .Z(n127) );
  NANDN U186 ( .A(n3), .B(N570), .Z(n126) );
  NAND U187 ( .A(n128), .B(n129), .Z(z3[509]) );
  NANDN U188 ( .A(N518), .B(z2[509]), .Z(n129) );
  NANDN U189 ( .A(n3), .B(N1029), .Z(n128) );
  NAND U190 ( .A(n130), .B(n131), .Z(z3[508]) );
  NANDN U191 ( .A(N518), .B(z2[508]), .Z(n131) );
  NANDN U192 ( .A(n3), .B(N1028), .Z(n130) );
  NAND U193 ( .A(n132), .B(n133), .Z(z3[507]) );
  NANDN U194 ( .A(N518), .B(z2[507]), .Z(n133) );
  NANDN U195 ( .A(n3), .B(N1027), .Z(n132) );
  NAND U196 ( .A(n134), .B(n135), .Z(z3[506]) );
  NANDN U197 ( .A(N518), .B(z2[506]), .Z(n135) );
  NANDN U198 ( .A(n3), .B(N1026), .Z(n134) );
  NAND U199 ( .A(n136), .B(n137), .Z(z3[505]) );
  NANDN U200 ( .A(N518), .B(z2[505]), .Z(n137) );
  NANDN U201 ( .A(n3), .B(N1025), .Z(n136) );
  NAND U202 ( .A(n138), .B(n139), .Z(z3[504]) );
  NANDN U203 ( .A(N518), .B(z2[504]), .Z(n139) );
  NANDN U204 ( .A(n3), .B(N1024), .Z(n138) );
  NAND U205 ( .A(n140), .B(n141), .Z(z3[503]) );
  NANDN U206 ( .A(N518), .B(z2[503]), .Z(n141) );
  NANDN U207 ( .A(n3), .B(N1023), .Z(n140) );
  NAND U208 ( .A(n142), .B(n143), .Z(z3[502]) );
  NANDN U209 ( .A(N518), .B(z2[502]), .Z(n143) );
  NANDN U210 ( .A(n3), .B(N1022), .Z(n142) );
  NAND U211 ( .A(n144), .B(n145), .Z(z3[501]) );
  NANDN U212 ( .A(N518), .B(z2[501]), .Z(n145) );
  NANDN U213 ( .A(n3), .B(N1021), .Z(n144) );
  NAND U214 ( .A(n146), .B(n147), .Z(z3[500]) );
  NANDN U215 ( .A(N518), .B(z2[500]), .Z(n147) );
  NANDN U216 ( .A(n3), .B(N1020), .Z(n146) );
  NAND U217 ( .A(n148), .B(n149), .Z(z3[4]) );
  NANDN U218 ( .A(N518), .B(z2[4]), .Z(n149) );
  NANDN U219 ( .A(n3), .B(N524), .Z(n148) );
  NAND U220 ( .A(n150), .B(n151), .Z(z3[49]) );
  NANDN U221 ( .A(N518), .B(z2[49]), .Z(n151) );
  NANDN U222 ( .A(n3), .B(N569), .Z(n150) );
  NAND U223 ( .A(n152), .B(n153), .Z(z3[499]) );
  NANDN U224 ( .A(N518), .B(z2[499]), .Z(n153) );
  NANDN U225 ( .A(n3), .B(N1019), .Z(n152) );
  NAND U226 ( .A(n154), .B(n155), .Z(z3[498]) );
  NANDN U227 ( .A(N518), .B(z2[498]), .Z(n155) );
  NANDN U228 ( .A(n3), .B(N1018), .Z(n154) );
  NAND U229 ( .A(n156), .B(n157), .Z(z3[497]) );
  NANDN U230 ( .A(N518), .B(z2[497]), .Z(n157) );
  NANDN U231 ( .A(n3), .B(N1017), .Z(n156) );
  NAND U232 ( .A(n158), .B(n159), .Z(z3[496]) );
  NANDN U233 ( .A(N518), .B(z2[496]), .Z(n159) );
  NANDN U234 ( .A(n3), .B(N1016), .Z(n158) );
  NAND U235 ( .A(n160), .B(n161), .Z(z3[495]) );
  NANDN U236 ( .A(N518), .B(z2[495]), .Z(n161) );
  NANDN U237 ( .A(n3), .B(N1015), .Z(n160) );
  NAND U238 ( .A(n162), .B(n163), .Z(z3[494]) );
  NANDN U239 ( .A(N518), .B(z2[494]), .Z(n163) );
  NANDN U240 ( .A(n3), .B(N1014), .Z(n162) );
  NAND U241 ( .A(n164), .B(n165), .Z(z3[493]) );
  NANDN U242 ( .A(N518), .B(z2[493]), .Z(n165) );
  NANDN U243 ( .A(n3), .B(N1013), .Z(n164) );
  NAND U244 ( .A(n166), .B(n167), .Z(z3[492]) );
  NANDN U245 ( .A(N518), .B(z2[492]), .Z(n167) );
  NANDN U246 ( .A(n3), .B(N1012), .Z(n166) );
  NAND U247 ( .A(n168), .B(n169), .Z(z3[491]) );
  NANDN U248 ( .A(N518), .B(z2[491]), .Z(n169) );
  NANDN U249 ( .A(n3), .B(N1011), .Z(n168) );
  NAND U250 ( .A(n170), .B(n171), .Z(z3[490]) );
  NANDN U251 ( .A(N518), .B(z2[490]), .Z(n171) );
  NANDN U252 ( .A(n3), .B(N1010), .Z(n170) );
  NAND U253 ( .A(n172), .B(n173), .Z(z3[48]) );
  NANDN U254 ( .A(N518), .B(z2[48]), .Z(n173) );
  NANDN U255 ( .A(n3), .B(N568), .Z(n172) );
  NAND U256 ( .A(n174), .B(n175), .Z(z3[489]) );
  NANDN U257 ( .A(N518), .B(z2[489]), .Z(n175) );
  NANDN U258 ( .A(n3), .B(N1009), .Z(n174) );
  NAND U259 ( .A(n176), .B(n177), .Z(z3[488]) );
  NANDN U260 ( .A(N518), .B(z2[488]), .Z(n177) );
  NANDN U261 ( .A(n3), .B(N1008), .Z(n176) );
  NAND U262 ( .A(n178), .B(n179), .Z(z3[487]) );
  NANDN U263 ( .A(N518), .B(z2[487]), .Z(n179) );
  NANDN U264 ( .A(n3), .B(N1007), .Z(n178) );
  NAND U265 ( .A(n180), .B(n181), .Z(z3[486]) );
  NANDN U266 ( .A(N518), .B(z2[486]), .Z(n181) );
  NANDN U267 ( .A(n3), .B(N1006), .Z(n180) );
  NAND U268 ( .A(n182), .B(n183), .Z(z3[485]) );
  NANDN U269 ( .A(N518), .B(z2[485]), .Z(n183) );
  NANDN U270 ( .A(n3), .B(N1005), .Z(n182) );
  NAND U271 ( .A(n184), .B(n185), .Z(z3[484]) );
  NANDN U272 ( .A(N518), .B(z2[484]), .Z(n185) );
  NANDN U273 ( .A(n3), .B(N1004), .Z(n184) );
  NAND U274 ( .A(n186), .B(n187), .Z(z3[483]) );
  NANDN U275 ( .A(N518), .B(z2[483]), .Z(n187) );
  NANDN U276 ( .A(n3), .B(N1003), .Z(n186) );
  NAND U277 ( .A(n188), .B(n189), .Z(z3[482]) );
  NANDN U278 ( .A(N518), .B(z2[482]), .Z(n189) );
  NANDN U279 ( .A(n3), .B(N1002), .Z(n188) );
  NAND U280 ( .A(n190), .B(n191), .Z(z3[481]) );
  NANDN U281 ( .A(N518), .B(z2[481]), .Z(n191) );
  NANDN U282 ( .A(n3), .B(N1001), .Z(n190) );
  NAND U283 ( .A(n192), .B(n193), .Z(z3[480]) );
  NANDN U284 ( .A(N518), .B(z2[480]), .Z(n193) );
  NANDN U285 ( .A(n3), .B(N1000), .Z(n192) );
  NAND U286 ( .A(n194), .B(n195), .Z(z3[47]) );
  NANDN U287 ( .A(N518), .B(z2[47]), .Z(n195) );
  NANDN U288 ( .A(n3), .B(N567), .Z(n194) );
  NAND U289 ( .A(n196), .B(n197), .Z(z3[479]) );
  NANDN U290 ( .A(N518), .B(z2[479]), .Z(n197) );
  NANDN U291 ( .A(n3), .B(N999), .Z(n196) );
  NAND U292 ( .A(n198), .B(n199), .Z(z3[478]) );
  NANDN U293 ( .A(N518), .B(z2[478]), .Z(n199) );
  NANDN U294 ( .A(n3), .B(N998), .Z(n198) );
  NAND U295 ( .A(n200), .B(n201), .Z(z3[477]) );
  NANDN U296 ( .A(N518), .B(z2[477]), .Z(n201) );
  NANDN U297 ( .A(n3), .B(N997), .Z(n200) );
  NAND U298 ( .A(n202), .B(n203), .Z(z3[476]) );
  NANDN U299 ( .A(N518), .B(z2[476]), .Z(n203) );
  NANDN U300 ( .A(n3), .B(N996), .Z(n202) );
  NAND U301 ( .A(n204), .B(n205), .Z(z3[475]) );
  NANDN U302 ( .A(N518), .B(z2[475]), .Z(n205) );
  NANDN U303 ( .A(n3), .B(N995), .Z(n204) );
  NAND U304 ( .A(n206), .B(n207), .Z(z3[474]) );
  NANDN U305 ( .A(N518), .B(z2[474]), .Z(n207) );
  NANDN U306 ( .A(n3), .B(N994), .Z(n206) );
  NAND U307 ( .A(n208), .B(n209), .Z(z3[473]) );
  NANDN U308 ( .A(N518), .B(z2[473]), .Z(n209) );
  NANDN U309 ( .A(n3), .B(N993), .Z(n208) );
  NAND U310 ( .A(n210), .B(n211), .Z(z3[472]) );
  NANDN U311 ( .A(N518), .B(z2[472]), .Z(n211) );
  NANDN U312 ( .A(n3), .B(N992), .Z(n210) );
  NAND U313 ( .A(n212), .B(n213), .Z(z3[471]) );
  NANDN U314 ( .A(N518), .B(z2[471]), .Z(n213) );
  NANDN U315 ( .A(n3), .B(N991), .Z(n212) );
  NAND U316 ( .A(n214), .B(n215), .Z(z3[470]) );
  NANDN U317 ( .A(N518), .B(z2[470]), .Z(n215) );
  NANDN U318 ( .A(n3), .B(N990), .Z(n214) );
  NAND U319 ( .A(n216), .B(n217), .Z(z3[46]) );
  NANDN U320 ( .A(N518), .B(z2[46]), .Z(n217) );
  NANDN U321 ( .A(n3), .B(N566), .Z(n216) );
  NAND U322 ( .A(n218), .B(n219), .Z(z3[469]) );
  NANDN U323 ( .A(N518), .B(z2[469]), .Z(n219) );
  NANDN U324 ( .A(n3), .B(N989), .Z(n218) );
  NAND U325 ( .A(n220), .B(n221), .Z(z3[468]) );
  NANDN U326 ( .A(N518), .B(z2[468]), .Z(n221) );
  NANDN U327 ( .A(n3), .B(N988), .Z(n220) );
  NAND U328 ( .A(n222), .B(n223), .Z(z3[467]) );
  NANDN U329 ( .A(N518), .B(z2[467]), .Z(n223) );
  NANDN U330 ( .A(n3), .B(N987), .Z(n222) );
  NAND U331 ( .A(n224), .B(n225), .Z(z3[466]) );
  NANDN U332 ( .A(N518), .B(z2[466]), .Z(n225) );
  NANDN U333 ( .A(n3), .B(N986), .Z(n224) );
  NAND U334 ( .A(n226), .B(n227), .Z(z3[465]) );
  NANDN U335 ( .A(N518), .B(z2[465]), .Z(n227) );
  NANDN U336 ( .A(n3), .B(N985), .Z(n226) );
  NAND U337 ( .A(n228), .B(n229), .Z(z3[464]) );
  NANDN U338 ( .A(N518), .B(z2[464]), .Z(n229) );
  NANDN U339 ( .A(n3), .B(N984), .Z(n228) );
  NAND U340 ( .A(n230), .B(n231), .Z(z3[463]) );
  NANDN U341 ( .A(N518), .B(z2[463]), .Z(n231) );
  NANDN U342 ( .A(n3), .B(N983), .Z(n230) );
  NAND U343 ( .A(n232), .B(n233), .Z(z3[462]) );
  NANDN U344 ( .A(N518), .B(z2[462]), .Z(n233) );
  NANDN U345 ( .A(n3), .B(N982), .Z(n232) );
  NAND U346 ( .A(n234), .B(n235), .Z(z3[461]) );
  NANDN U347 ( .A(N518), .B(z2[461]), .Z(n235) );
  NANDN U348 ( .A(n3), .B(N981), .Z(n234) );
  NAND U349 ( .A(n236), .B(n237), .Z(z3[460]) );
  NANDN U350 ( .A(N518), .B(z2[460]), .Z(n237) );
  NANDN U351 ( .A(n3), .B(N980), .Z(n236) );
  NAND U352 ( .A(n238), .B(n239), .Z(z3[45]) );
  NANDN U353 ( .A(N518), .B(z2[45]), .Z(n239) );
  NANDN U354 ( .A(n3), .B(N565), .Z(n238) );
  NAND U355 ( .A(n240), .B(n241), .Z(z3[459]) );
  NANDN U356 ( .A(N518), .B(z2[459]), .Z(n241) );
  NANDN U357 ( .A(n3), .B(N979), .Z(n240) );
  NAND U358 ( .A(n242), .B(n243), .Z(z3[458]) );
  NANDN U359 ( .A(N518), .B(z2[458]), .Z(n243) );
  NANDN U360 ( .A(n3), .B(N978), .Z(n242) );
  NAND U361 ( .A(n244), .B(n245), .Z(z3[457]) );
  NANDN U362 ( .A(N518), .B(z2[457]), .Z(n245) );
  NANDN U363 ( .A(n3), .B(N977), .Z(n244) );
  NAND U364 ( .A(n246), .B(n247), .Z(z3[456]) );
  NANDN U365 ( .A(N518), .B(z2[456]), .Z(n247) );
  NANDN U366 ( .A(n3), .B(N976), .Z(n246) );
  NAND U367 ( .A(n248), .B(n249), .Z(z3[455]) );
  NANDN U368 ( .A(N518), .B(z2[455]), .Z(n249) );
  NANDN U369 ( .A(n3), .B(N975), .Z(n248) );
  NAND U370 ( .A(n250), .B(n251), .Z(z3[454]) );
  NANDN U371 ( .A(N518), .B(z2[454]), .Z(n251) );
  NANDN U372 ( .A(n3), .B(N974), .Z(n250) );
  NAND U373 ( .A(n252), .B(n253), .Z(z3[453]) );
  NANDN U374 ( .A(N518), .B(z2[453]), .Z(n253) );
  NANDN U375 ( .A(n3), .B(N973), .Z(n252) );
  NAND U376 ( .A(n254), .B(n255), .Z(z3[452]) );
  NANDN U377 ( .A(N518), .B(z2[452]), .Z(n255) );
  NANDN U378 ( .A(n3), .B(N972), .Z(n254) );
  NAND U379 ( .A(n256), .B(n257), .Z(z3[451]) );
  NANDN U380 ( .A(N518), .B(z2[451]), .Z(n257) );
  NANDN U381 ( .A(n3), .B(N971), .Z(n256) );
  NAND U382 ( .A(n258), .B(n259), .Z(z3[450]) );
  NANDN U383 ( .A(N518), .B(z2[450]), .Z(n259) );
  NANDN U384 ( .A(n3), .B(N970), .Z(n258) );
  NAND U385 ( .A(n260), .B(n261), .Z(z3[44]) );
  NANDN U386 ( .A(N518), .B(z2[44]), .Z(n261) );
  NANDN U387 ( .A(n3), .B(N564), .Z(n260) );
  NAND U388 ( .A(n262), .B(n263), .Z(z3[449]) );
  NANDN U389 ( .A(N518), .B(z2[449]), .Z(n263) );
  NANDN U390 ( .A(n3), .B(N969), .Z(n262) );
  NAND U391 ( .A(n264), .B(n265), .Z(z3[448]) );
  NANDN U392 ( .A(N518), .B(z2[448]), .Z(n265) );
  NANDN U393 ( .A(n3), .B(N968), .Z(n264) );
  NAND U394 ( .A(n266), .B(n267), .Z(z3[447]) );
  NANDN U395 ( .A(N518), .B(z2[447]), .Z(n267) );
  NANDN U396 ( .A(n3), .B(N967), .Z(n266) );
  NAND U397 ( .A(n268), .B(n269), .Z(z3[446]) );
  NANDN U398 ( .A(N518), .B(z2[446]), .Z(n269) );
  NANDN U399 ( .A(n3), .B(N966), .Z(n268) );
  NAND U400 ( .A(n270), .B(n271), .Z(z3[445]) );
  NANDN U401 ( .A(N518), .B(z2[445]), .Z(n271) );
  NANDN U402 ( .A(n3), .B(N965), .Z(n270) );
  NAND U403 ( .A(n272), .B(n273), .Z(z3[444]) );
  NANDN U404 ( .A(N518), .B(z2[444]), .Z(n273) );
  NANDN U405 ( .A(n3), .B(N964), .Z(n272) );
  NAND U406 ( .A(n274), .B(n275), .Z(z3[443]) );
  NANDN U407 ( .A(N518), .B(z2[443]), .Z(n275) );
  NANDN U408 ( .A(n3), .B(N963), .Z(n274) );
  NAND U409 ( .A(n276), .B(n277), .Z(z3[442]) );
  NANDN U410 ( .A(N518), .B(z2[442]), .Z(n277) );
  NANDN U411 ( .A(n3), .B(N962), .Z(n276) );
  NAND U412 ( .A(n278), .B(n279), .Z(z3[441]) );
  NANDN U413 ( .A(N518), .B(z2[441]), .Z(n279) );
  NANDN U414 ( .A(n3), .B(N961), .Z(n278) );
  NAND U415 ( .A(n280), .B(n281), .Z(z3[440]) );
  NANDN U416 ( .A(N518), .B(z2[440]), .Z(n281) );
  NANDN U417 ( .A(n3), .B(N960), .Z(n280) );
  NAND U418 ( .A(n282), .B(n283), .Z(z3[43]) );
  NANDN U419 ( .A(N518), .B(z2[43]), .Z(n283) );
  NANDN U420 ( .A(n3), .B(N563), .Z(n282) );
  NAND U421 ( .A(n284), .B(n285), .Z(z3[439]) );
  NANDN U422 ( .A(N518), .B(z2[439]), .Z(n285) );
  NANDN U423 ( .A(n3), .B(N959), .Z(n284) );
  NAND U424 ( .A(n286), .B(n287), .Z(z3[438]) );
  NANDN U425 ( .A(N518), .B(z2[438]), .Z(n287) );
  NANDN U426 ( .A(n3), .B(N958), .Z(n286) );
  NAND U427 ( .A(n288), .B(n289), .Z(z3[437]) );
  NANDN U428 ( .A(N518), .B(z2[437]), .Z(n289) );
  NANDN U429 ( .A(n3), .B(N957), .Z(n288) );
  NAND U430 ( .A(n290), .B(n291), .Z(z3[436]) );
  NANDN U431 ( .A(N518), .B(z2[436]), .Z(n291) );
  NANDN U432 ( .A(n3), .B(N956), .Z(n290) );
  NAND U433 ( .A(n292), .B(n293), .Z(z3[435]) );
  NANDN U434 ( .A(N518), .B(z2[435]), .Z(n293) );
  NANDN U435 ( .A(n3), .B(N955), .Z(n292) );
  NAND U436 ( .A(n294), .B(n295), .Z(z3[434]) );
  NANDN U437 ( .A(N518), .B(z2[434]), .Z(n295) );
  NANDN U438 ( .A(n3), .B(N954), .Z(n294) );
  NAND U439 ( .A(n296), .B(n297), .Z(z3[433]) );
  NANDN U440 ( .A(N518), .B(z2[433]), .Z(n297) );
  NANDN U441 ( .A(n3), .B(N953), .Z(n296) );
  NAND U442 ( .A(n298), .B(n299), .Z(z3[432]) );
  NANDN U443 ( .A(N518), .B(z2[432]), .Z(n299) );
  NANDN U444 ( .A(n3), .B(N952), .Z(n298) );
  NAND U445 ( .A(n300), .B(n301), .Z(z3[431]) );
  NANDN U446 ( .A(N518), .B(z2[431]), .Z(n301) );
  NANDN U447 ( .A(n3), .B(N951), .Z(n300) );
  NAND U448 ( .A(n302), .B(n303), .Z(z3[430]) );
  NANDN U449 ( .A(N518), .B(z2[430]), .Z(n303) );
  NANDN U450 ( .A(n3), .B(N950), .Z(n302) );
  NAND U451 ( .A(n304), .B(n305), .Z(z3[42]) );
  NANDN U452 ( .A(N518), .B(z2[42]), .Z(n305) );
  NANDN U453 ( .A(n3), .B(N562), .Z(n304) );
  NAND U454 ( .A(n306), .B(n307), .Z(z3[429]) );
  NANDN U455 ( .A(N518), .B(z2[429]), .Z(n307) );
  NANDN U456 ( .A(n3), .B(N949), .Z(n306) );
  NAND U457 ( .A(n308), .B(n309), .Z(z3[428]) );
  NANDN U458 ( .A(N518), .B(z2[428]), .Z(n309) );
  NANDN U459 ( .A(n3), .B(N948), .Z(n308) );
  NAND U460 ( .A(n310), .B(n311), .Z(z3[427]) );
  NANDN U461 ( .A(N518), .B(z2[427]), .Z(n311) );
  NANDN U462 ( .A(n3), .B(N947), .Z(n310) );
  NAND U463 ( .A(n312), .B(n313), .Z(z3[426]) );
  NANDN U464 ( .A(N518), .B(z2[426]), .Z(n313) );
  NANDN U465 ( .A(n3), .B(N946), .Z(n312) );
  NAND U466 ( .A(n314), .B(n315), .Z(z3[425]) );
  NANDN U467 ( .A(N518), .B(z2[425]), .Z(n315) );
  NANDN U468 ( .A(n3), .B(N945), .Z(n314) );
  NAND U469 ( .A(n316), .B(n317), .Z(z3[424]) );
  NANDN U470 ( .A(N518), .B(z2[424]), .Z(n317) );
  NANDN U471 ( .A(n3), .B(N944), .Z(n316) );
  NAND U472 ( .A(n318), .B(n319), .Z(z3[423]) );
  NANDN U473 ( .A(N518), .B(z2[423]), .Z(n319) );
  NANDN U474 ( .A(n3), .B(N943), .Z(n318) );
  NAND U475 ( .A(n320), .B(n321), .Z(z3[422]) );
  NANDN U476 ( .A(N518), .B(z2[422]), .Z(n321) );
  NANDN U477 ( .A(n3), .B(N942), .Z(n320) );
  NAND U478 ( .A(n322), .B(n323), .Z(z3[421]) );
  NANDN U479 ( .A(N518), .B(z2[421]), .Z(n323) );
  NANDN U480 ( .A(n3), .B(N941), .Z(n322) );
  NAND U481 ( .A(n324), .B(n325), .Z(z3[420]) );
  NANDN U482 ( .A(N518), .B(z2[420]), .Z(n325) );
  NANDN U483 ( .A(n3), .B(N940), .Z(n324) );
  NAND U484 ( .A(n326), .B(n327), .Z(z3[41]) );
  NANDN U485 ( .A(N518), .B(z2[41]), .Z(n327) );
  NANDN U486 ( .A(n3), .B(N561), .Z(n326) );
  NAND U487 ( .A(n328), .B(n329), .Z(z3[419]) );
  NANDN U488 ( .A(N518), .B(z2[419]), .Z(n329) );
  NANDN U489 ( .A(n3), .B(N939), .Z(n328) );
  NAND U490 ( .A(n330), .B(n331), .Z(z3[418]) );
  NANDN U491 ( .A(N518), .B(z2[418]), .Z(n331) );
  NANDN U492 ( .A(n3), .B(N938), .Z(n330) );
  NAND U493 ( .A(n332), .B(n333), .Z(z3[417]) );
  NANDN U494 ( .A(N518), .B(z2[417]), .Z(n333) );
  NANDN U495 ( .A(n3), .B(N937), .Z(n332) );
  NAND U496 ( .A(n334), .B(n335), .Z(z3[416]) );
  NANDN U497 ( .A(N518), .B(z2[416]), .Z(n335) );
  NANDN U498 ( .A(n3), .B(N936), .Z(n334) );
  NAND U499 ( .A(n336), .B(n337), .Z(z3[415]) );
  NANDN U500 ( .A(N518), .B(z2[415]), .Z(n337) );
  NANDN U501 ( .A(n3), .B(N935), .Z(n336) );
  NAND U502 ( .A(n338), .B(n339), .Z(z3[414]) );
  NANDN U503 ( .A(N518), .B(z2[414]), .Z(n339) );
  NANDN U504 ( .A(n3), .B(N934), .Z(n338) );
  NAND U505 ( .A(n340), .B(n341), .Z(z3[413]) );
  NANDN U506 ( .A(N518), .B(z2[413]), .Z(n341) );
  NANDN U507 ( .A(n3), .B(N933), .Z(n340) );
  NAND U508 ( .A(n342), .B(n343), .Z(z3[412]) );
  NANDN U509 ( .A(N518), .B(z2[412]), .Z(n343) );
  NANDN U510 ( .A(n3), .B(N932), .Z(n342) );
  NAND U511 ( .A(n344), .B(n345), .Z(z3[411]) );
  NANDN U512 ( .A(N518), .B(z2[411]), .Z(n345) );
  NANDN U513 ( .A(n3), .B(N931), .Z(n344) );
  NAND U514 ( .A(n346), .B(n347), .Z(z3[410]) );
  NANDN U515 ( .A(N518), .B(z2[410]), .Z(n347) );
  NANDN U516 ( .A(n3), .B(N930), .Z(n346) );
  NAND U517 ( .A(n348), .B(n349), .Z(z3[40]) );
  NANDN U518 ( .A(N518), .B(z2[40]), .Z(n349) );
  NANDN U519 ( .A(n3), .B(N560), .Z(n348) );
  NAND U520 ( .A(n350), .B(n351), .Z(z3[409]) );
  NANDN U521 ( .A(N518), .B(z2[409]), .Z(n351) );
  NANDN U522 ( .A(n3), .B(N929), .Z(n350) );
  NAND U523 ( .A(n352), .B(n353), .Z(z3[408]) );
  NANDN U524 ( .A(N518), .B(z2[408]), .Z(n353) );
  NANDN U525 ( .A(n3), .B(N928), .Z(n352) );
  NAND U526 ( .A(n354), .B(n355), .Z(z3[407]) );
  NANDN U527 ( .A(N518), .B(z2[407]), .Z(n355) );
  NANDN U528 ( .A(n3), .B(N927), .Z(n354) );
  NAND U529 ( .A(n356), .B(n357), .Z(z3[406]) );
  NANDN U530 ( .A(N518), .B(z2[406]), .Z(n357) );
  NANDN U531 ( .A(n3), .B(N926), .Z(n356) );
  NAND U532 ( .A(n358), .B(n359), .Z(z3[405]) );
  NANDN U533 ( .A(N518), .B(z2[405]), .Z(n359) );
  NANDN U534 ( .A(n3), .B(N925), .Z(n358) );
  NAND U535 ( .A(n360), .B(n361), .Z(z3[404]) );
  NANDN U536 ( .A(N518), .B(z2[404]), .Z(n361) );
  NANDN U537 ( .A(n3), .B(N924), .Z(n360) );
  NAND U538 ( .A(n362), .B(n363), .Z(z3[403]) );
  NANDN U539 ( .A(N518), .B(z2[403]), .Z(n363) );
  NANDN U540 ( .A(n3), .B(N923), .Z(n362) );
  NAND U541 ( .A(n364), .B(n365), .Z(z3[402]) );
  NANDN U542 ( .A(N518), .B(z2[402]), .Z(n365) );
  NANDN U543 ( .A(n3), .B(N922), .Z(n364) );
  NAND U544 ( .A(n366), .B(n367), .Z(z3[401]) );
  NANDN U545 ( .A(N518), .B(z2[401]), .Z(n367) );
  NANDN U546 ( .A(n3), .B(N921), .Z(n366) );
  NAND U547 ( .A(n368), .B(n369), .Z(z3[400]) );
  NANDN U548 ( .A(N518), .B(z2[400]), .Z(n369) );
  NANDN U549 ( .A(n3), .B(N920), .Z(n368) );
  NAND U550 ( .A(n370), .B(n371), .Z(z3[3]) );
  NANDN U551 ( .A(N518), .B(z2[3]), .Z(n371) );
  NANDN U552 ( .A(n3), .B(N523), .Z(n370) );
  NAND U553 ( .A(n372), .B(n373), .Z(z3[39]) );
  NANDN U554 ( .A(N518), .B(z2[39]), .Z(n373) );
  NANDN U555 ( .A(n3), .B(N559), .Z(n372) );
  NAND U556 ( .A(n374), .B(n375), .Z(z3[399]) );
  NANDN U557 ( .A(N518), .B(z2[399]), .Z(n375) );
  NANDN U558 ( .A(n3), .B(N919), .Z(n374) );
  NAND U559 ( .A(n376), .B(n377), .Z(z3[398]) );
  NANDN U560 ( .A(N518), .B(z2[398]), .Z(n377) );
  NANDN U561 ( .A(n3), .B(N918), .Z(n376) );
  NAND U562 ( .A(n378), .B(n379), .Z(z3[397]) );
  NANDN U563 ( .A(N518), .B(z2[397]), .Z(n379) );
  NANDN U564 ( .A(n3), .B(N917), .Z(n378) );
  NAND U565 ( .A(n380), .B(n381), .Z(z3[396]) );
  NANDN U566 ( .A(N518), .B(z2[396]), .Z(n381) );
  NANDN U567 ( .A(n3), .B(N916), .Z(n380) );
  NAND U568 ( .A(n382), .B(n383), .Z(z3[395]) );
  NANDN U569 ( .A(N518), .B(z2[395]), .Z(n383) );
  NANDN U570 ( .A(n3), .B(N915), .Z(n382) );
  NAND U571 ( .A(n384), .B(n385), .Z(z3[394]) );
  NANDN U572 ( .A(N518), .B(z2[394]), .Z(n385) );
  NANDN U573 ( .A(n3), .B(N914), .Z(n384) );
  NAND U574 ( .A(n386), .B(n387), .Z(z3[393]) );
  NANDN U575 ( .A(N518), .B(z2[393]), .Z(n387) );
  NANDN U576 ( .A(n3), .B(N913), .Z(n386) );
  NAND U577 ( .A(n388), .B(n389), .Z(z3[392]) );
  NANDN U578 ( .A(N518), .B(z2[392]), .Z(n389) );
  NANDN U579 ( .A(n3), .B(N912), .Z(n388) );
  NAND U580 ( .A(n390), .B(n391), .Z(z3[391]) );
  NANDN U581 ( .A(N518), .B(z2[391]), .Z(n391) );
  NANDN U582 ( .A(n3), .B(N911), .Z(n390) );
  NAND U583 ( .A(n392), .B(n393), .Z(z3[390]) );
  NANDN U584 ( .A(N518), .B(z2[390]), .Z(n393) );
  NANDN U585 ( .A(n3), .B(N910), .Z(n392) );
  NAND U586 ( .A(n394), .B(n395), .Z(z3[38]) );
  NANDN U587 ( .A(N518), .B(z2[38]), .Z(n395) );
  NANDN U588 ( .A(n3), .B(N558), .Z(n394) );
  NAND U589 ( .A(n396), .B(n397), .Z(z3[389]) );
  NANDN U590 ( .A(N518), .B(z2[389]), .Z(n397) );
  NANDN U591 ( .A(n3), .B(N909), .Z(n396) );
  NAND U592 ( .A(n398), .B(n399), .Z(z3[388]) );
  NANDN U593 ( .A(N518), .B(z2[388]), .Z(n399) );
  NANDN U594 ( .A(n3), .B(N908), .Z(n398) );
  NAND U595 ( .A(n400), .B(n401), .Z(z3[387]) );
  NANDN U596 ( .A(N518), .B(z2[387]), .Z(n401) );
  NANDN U597 ( .A(n3), .B(N907), .Z(n400) );
  NAND U598 ( .A(n402), .B(n403), .Z(z3[386]) );
  NANDN U599 ( .A(N518), .B(z2[386]), .Z(n403) );
  NANDN U600 ( .A(n3), .B(N906), .Z(n402) );
  NAND U601 ( .A(n404), .B(n405), .Z(z3[385]) );
  NANDN U602 ( .A(N518), .B(z2[385]), .Z(n405) );
  NANDN U603 ( .A(n3), .B(N905), .Z(n404) );
  NAND U604 ( .A(n406), .B(n407), .Z(z3[384]) );
  NANDN U605 ( .A(N518), .B(z2[384]), .Z(n407) );
  NANDN U606 ( .A(n3), .B(N904), .Z(n406) );
  NAND U607 ( .A(n408), .B(n409), .Z(z3[383]) );
  NANDN U608 ( .A(N518), .B(z2[383]), .Z(n409) );
  NANDN U609 ( .A(n3), .B(N903), .Z(n408) );
  NAND U610 ( .A(n410), .B(n411), .Z(z3[382]) );
  NANDN U611 ( .A(N518), .B(z2[382]), .Z(n411) );
  NANDN U612 ( .A(n3), .B(N902), .Z(n410) );
  NAND U613 ( .A(n412), .B(n413), .Z(z3[381]) );
  NANDN U614 ( .A(N518), .B(z2[381]), .Z(n413) );
  NANDN U615 ( .A(n3), .B(N901), .Z(n412) );
  NAND U616 ( .A(n414), .B(n415), .Z(z3[380]) );
  NANDN U617 ( .A(N518), .B(z2[380]), .Z(n415) );
  NANDN U618 ( .A(n3), .B(N900), .Z(n414) );
  NAND U619 ( .A(n416), .B(n417), .Z(z3[37]) );
  NANDN U620 ( .A(N518), .B(z2[37]), .Z(n417) );
  NANDN U621 ( .A(n3), .B(N557), .Z(n416) );
  NAND U622 ( .A(n418), .B(n419), .Z(z3[379]) );
  NANDN U623 ( .A(N518), .B(z2[379]), .Z(n419) );
  NANDN U624 ( .A(n3), .B(N899), .Z(n418) );
  NAND U625 ( .A(n420), .B(n421), .Z(z3[378]) );
  NANDN U626 ( .A(N518), .B(z2[378]), .Z(n421) );
  NANDN U627 ( .A(n3), .B(N898), .Z(n420) );
  NAND U628 ( .A(n422), .B(n423), .Z(z3[377]) );
  NANDN U629 ( .A(N518), .B(z2[377]), .Z(n423) );
  NANDN U630 ( .A(n3), .B(N897), .Z(n422) );
  NAND U631 ( .A(n424), .B(n425), .Z(z3[376]) );
  NANDN U632 ( .A(N518), .B(z2[376]), .Z(n425) );
  NANDN U633 ( .A(n3), .B(N896), .Z(n424) );
  NAND U634 ( .A(n426), .B(n427), .Z(z3[375]) );
  NANDN U635 ( .A(N518), .B(z2[375]), .Z(n427) );
  NANDN U636 ( .A(n3), .B(N895), .Z(n426) );
  NAND U637 ( .A(n428), .B(n429), .Z(z3[374]) );
  NANDN U638 ( .A(N518), .B(z2[374]), .Z(n429) );
  NANDN U639 ( .A(n3), .B(N894), .Z(n428) );
  NAND U640 ( .A(n430), .B(n431), .Z(z3[373]) );
  NANDN U641 ( .A(N518), .B(z2[373]), .Z(n431) );
  NANDN U642 ( .A(n3), .B(N893), .Z(n430) );
  NAND U643 ( .A(n432), .B(n433), .Z(z3[372]) );
  NANDN U644 ( .A(N518), .B(z2[372]), .Z(n433) );
  NANDN U645 ( .A(n3), .B(N892), .Z(n432) );
  NAND U646 ( .A(n434), .B(n435), .Z(z3[371]) );
  NANDN U647 ( .A(N518), .B(z2[371]), .Z(n435) );
  NANDN U648 ( .A(n3), .B(N891), .Z(n434) );
  NAND U649 ( .A(n436), .B(n437), .Z(z3[370]) );
  NANDN U650 ( .A(N518), .B(z2[370]), .Z(n437) );
  NANDN U651 ( .A(n3), .B(N890), .Z(n436) );
  NAND U652 ( .A(n438), .B(n439), .Z(z3[36]) );
  NANDN U653 ( .A(N518), .B(z2[36]), .Z(n439) );
  NANDN U654 ( .A(n3), .B(N556), .Z(n438) );
  NAND U655 ( .A(n440), .B(n441), .Z(z3[369]) );
  NANDN U656 ( .A(N518), .B(z2[369]), .Z(n441) );
  NANDN U657 ( .A(n3), .B(N889), .Z(n440) );
  NAND U658 ( .A(n442), .B(n443), .Z(z3[368]) );
  NANDN U659 ( .A(N518), .B(z2[368]), .Z(n443) );
  NANDN U660 ( .A(n3), .B(N888), .Z(n442) );
  NAND U661 ( .A(n444), .B(n445), .Z(z3[367]) );
  NANDN U662 ( .A(N518), .B(z2[367]), .Z(n445) );
  NANDN U663 ( .A(n3), .B(N887), .Z(n444) );
  NAND U664 ( .A(n446), .B(n447), .Z(z3[366]) );
  NANDN U665 ( .A(N518), .B(z2[366]), .Z(n447) );
  NANDN U666 ( .A(n3), .B(N886), .Z(n446) );
  NAND U667 ( .A(n448), .B(n449), .Z(z3[365]) );
  NANDN U668 ( .A(N518), .B(z2[365]), .Z(n449) );
  NANDN U669 ( .A(n3), .B(N885), .Z(n448) );
  NAND U670 ( .A(n450), .B(n451), .Z(z3[364]) );
  NANDN U671 ( .A(N518), .B(z2[364]), .Z(n451) );
  NANDN U672 ( .A(n3), .B(N884), .Z(n450) );
  NAND U673 ( .A(n452), .B(n453), .Z(z3[363]) );
  NANDN U674 ( .A(N518), .B(z2[363]), .Z(n453) );
  NANDN U675 ( .A(n3), .B(N883), .Z(n452) );
  NAND U676 ( .A(n454), .B(n455), .Z(z3[362]) );
  NANDN U677 ( .A(N518), .B(z2[362]), .Z(n455) );
  NANDN U678 ( .A(n3), .B(N882), .Z(n454) );
  NAND U679 ( .A(n456), .B(n457), .Z(z3[361]) );
  NANDN U680 ( .A(N518), .B(z2[361]), .Z(n457) );
  NANDN U681 ( .A(n3), .B(N881), .Z(n456) );
  NAND U682 ( .A(n458), .B(n459), .Z(z3[360]) );
  NANDN U683 ( .A(N518), .B(z2[360]), .Z(n459) );
  NANDN U684 ( .A(n3), .B(N880), .Z(n458) );
  NAND U685 ( .A(n460), .B(n461), .Z(z3[35]) );
  NANDN U686 ( .A(N518), .B(z2[35]), .Z(n461) );
  NANDN U687 ( .A(n3), .B(N555), .Z(n460) );
  NAND U688 ( .A(n462), .B(n463), .Z(z3[359]) );
  NANDN U689 ( .A(N518), .B(z2[359]), .Z(n463) );
  NANDN U690 ( .A(n3), .B(N879), .Z(n462) );
  NAND U691 ( .A(n464), .B(n465), .Z(z3[358]) );
  NANDN U692 ( .A(N518), .B(z2[358]), .Z(n465) );
  NANDN U693 ( .A(n3), .B(N878), .Z(n464) );
  NAND U694 ( .A(n466), .B(n467), .Z(z3[357]) );
  NANDN U695 ( .A(N518), .B(z2[357]), .Z(n467) );
  NANDN U696 ( .A(n3), .B(N877), .Z(n466) );
  NAND U697 ( .A(n468), .B(n469), .Z(z3[356]) );
  NANDN U698 ( .A(N518), .B(z2[356]), .Z(n469) );
  NANDN U699 ( .A(n3), .B(N876), .Z(n468) );
  NAND U700 ( .A(n470), .B(n471), .Z(z3[355]) );
  NANDN U701 ( .A(N518), .B(z2[355]), .Z(n471) );
  NANDN U702 ( .A(n3), .B(N875), .Z(n470) );
  NAND U703 ( .A(n472), .B(n473), .Z(z3[354]) );
  NANDN U704 ( .A(N518), .B(z2[354]), .Z(n473) );
  NANDN U705 ( .A(n3), .B(N874), .Z(n472) );
  NAND U706 ( .A(n474), .B(n475), .Z(z3[353]) );
  NANDN U707 ( .A(N518), .B(z2[353]), .Z(n475) );
  NANDN U708 ( .A(n3), .B(N873), .Z(n474) );
  NAND U709 ( .A(n476), .B(n477), .Z(z3[352]) );
  NANDN U710 ( .A(N518), .B(z2[352]), .Z(n477) );
  NANDN U711 ( .A(n3), .B(N872), .Z(n476) );
  NAND U712 ( .A(n478), .B(n479), .Z(z3[351]) );
  NANDN U713 ( .A(N518), .B(z2[351]), .Z(n479) );
  NANDN U714 ( .A(n3), .B(N871), .Z(n478) );
  NAND U715 ( .A(n480), .B(n481), .Z(z3[350]) );
  NANDN U716 ( .A(N518), .B(z2[350]), .Z(n481) );
  NANDN U717 ( .A(n3), .B(N870), .Z(n480) );
  NAND U718 ( .A(n482), .B(n483), .Z(z3[34]) );
  NANDN U719 ( .A(N518), .B(z2[34]), .Z(n483) );
  NANDN U720 ( .A(n3), .B(N554), .Z(n482) );
  NAND U721 ( .A(n484), .B(n485), .Z(z3[349]) );
  NANDN U722 ( .A(N518), .B(z2[349]), .Z(n485) );
  NANDN U723 ( .A(n3), .B(N869), .Z(n484) );
  NAND U724 ( .A(n486), .B(n487), .Z(z3[348]) );
  NANDN U725 ( .A(N518), .B(z2[348]), .Z(n487) );
  NANDN U726 ( .A(n3), .B(N868), .Z(n486) );
  NAND U727 ( .A(n488), .B(n489), .Z(z3[347]) );
  NANDN U728 ( .A(N518), .B(z2[347]), .Z(n489) );
  NANDN U729 ( .A(n3), .B(N867), .Z(n488) );
  NAND U730 ( .A(n490), .B(n491), .Z(z3[346]) );
  NANDN U731 ( .A(N518), .B(z2[346]), .Z(n491) );
  NANDN U732 ( .A(n3), .B(N866), .Z(n490) );
  NAND U733 ( .A(n492), .B(n493), .Z(z3[345]) );
  NANDN U734 ( .A(N518), .B(z2[345]), .Z(n493) );
  NANDN U735 ( .A(n3), .B(N865), .Z(n492) );
  NAND U736 ( .A(n494), .B(n495), .Z(z3[344]) );
  NANDN U737 ( .A(N518), .B(z2[344]), .Z(n495) );
  NANDN U738 ( .A(n3), .B(N864), .Z(n494) );
  NAND U739 ( .A(n496), .B(n497), .Z(z3[343]) );
  NANDN U740 ( .A(N518), .B(z2[343]), .Z(n497) );
  NANDN U741 ( .A(n3), .B(N863), .Z(n496) );
  NAND U742 ( .A(n498), .B(n499), .Z(z3[342]) );
  NANDN U743 ( .A(N518), .B(z2[342]), .Z(n499) );
  NANDN U744 ( .A(n3), .B(N862), .Z(n498) );
  NAND U745 ( .A(n500), .B(n501), .Z(z3[341]) );
  NANDN U746 ( .A(N518), .B(z2[341]), .Z(n501) );
  NANDN U747 ( .A(n3), .B(N861), .Z(n500) );
  NAND U748 ( .A(n502), .B(n503), .Z(z3[340]) );
  NANDN U749 ( .A(N518), .B(z2[340]), .Z(n503) );
  NANDN U750 ( .A(n3), .B(N860), .Z(n502) );
  NAND U751 ( .A(n504), .B(n505), .Z(z3[33]) );
  NANDN U752 ( .A(N518), .B(z2[33]), .Z(n505) );
  NANDN U753 ( .A(n3), .B(N553), .Z(n504) );
  NAND U754 ( .A(n506), .B(n507), .Z(z3[339]) );
  NANDN U755 ( .A(N518), .B(z2[339]), .Z(n507) );
  NANDN U756 ( .A(n3), .B(N859), .Z(n506) );
  NAND U757 ( .A(n508), .B(n509), .Z(z3[338]) );
  NANDN U758 ( .A(N518), .B(z2[338]), .Z(n509) );
  NANDN U759 ( .A(n3), .B(N858), .Z(n508) );
  NAND U760 ( .A(n510), .B(n511), .Z(z3[337]) );
  NANDN U761 ( .A(N518), .B(z2[337]), .Z(n511) );
  NANDN U762 ( .A(n3), .B(N857), .Z(n510) );
  NAND U763 ( .A(n512), .B(n513), .Z(z3[336]) );
  NANDN U764 ( .A(N518), .B(z2[336]), .Z(n513) );
  NANDN U765 ( .A(n3), .B(N856), .Z(n512) );
  NAND U766 ( .A(n514), .B(n515), .Z(z3[335]) );
  NANDN U767 ( .A(N518), .B(z2[335]), .Z(n515) );
  NANDN U768 ( .A(n3), .B(N855), .Z(n514) );
  NAND U769 ( .A(n516), .B(n517), .Z(z3[334]) );
  NANDN U770 ( .A(N518), .B(z2[334]), .Z(n517) );
  NANDN U771 ( .A(n3), .B(N854), .Z(n516) );
  NAND U772 ( .A(n518), .B(n519), .Z(z3[333]) );
  NANDN U773 ( .A(N518), .B(z2[333]), .Z(n519) );
  NANDN U774 ( .A(n3), .B(N853), .Z(n518) );
  NAND U775 ( .A(n520), .B(n521), .Z(z3[332]) );
  NANDN U776 ( .A(N518), .B(z2[332]), .Z(n521) );
  NANDN U777 ( .A(n3), .B(N852), .Z(n520) );
  NAND U778 ( .A(n522), .B(n523), .Z(z3[331]) );
  NANDN U779 ( .A(N518), .B(z2[331]), .Z(n523) );
  NANDN U780 ( .A(n3), .B(N851), .Z(n522) );
  NAND U781 ( .A(n524), .B(n525), .Z(z3[330]) );
  NANDN U782 ( .A(N518), .B(z2[330]), .Z(n525) );
  NANDN U783 ( .A(n3), .B(N850), .Z(n524) );
  NAND U784 ( .A(n526), .B(n527), .Z(z3[32]) );
  NANDN U785 ( .A(N518), .B(z2[32]), .Z(n527) );
  NANDN U786 ( .A(n3), .B(N552), .Z(n526) );
  NAND U787 ( .A(n528), .B(n529), .Z(z3[329]) );
  NANDN U788 ( .A(N518), .B(z2[329]), .Z(n529) );
  NANDN U789 ( .A(n3), .B(N849), .Z(n528) );
  NAND U790 ( .A(n530), .B(n531), .Z(z3[328]) );
  NANDN U791 ( .A(N518), .B(z2[328]), .Z(n531) );
  NANDN U792 ( .A(n3), .B(N848), .Z(n530) );
  NAND U793 ( .A(n532), .B(n533), .Z(z3[327]) );
  NANDN U794 ( .A(N518), .B(z2[327]), .Z(n533) );
  NANDN U795 ( .A(n3), .B(N847), .Z(n532) );
  NAND U796 ( .A(n534), .B(n535), .Z(z3[326]) );
  NANDN U797 ( .A(N518), .B(z2[326]), .Z(n535) );
  NANDN U798 ( .A(n3), .B(N846), .Z(n534) );
  NAND U799 ( .A(n536), .B(n537), .Z(z3[325]) );
  NANDN U800 ( .A(N518), .B(z2[325]), .Z(n537) );
  NANDN U801 ( .A(n3), .B(N845), .Z(n536) );
  NAND U802 ( .A(n538), .B(n539), .Z(z3[324]) );
  NANDN U803 ( .A(N518), .B(z2[324]), .Z(n539) );
  NANDN U804 ( .A(n3), .B(N844), .Z(n538) );
  NAND U805 ( .A(n540), .B(n541), .Z(z3[323]) );
  NANDN U806 ( .A(N518), .B(z2[323]), .Z(n541) );
  NANDN U807 ( .A(n3), .B(N843), .Z(n540) );
  NAND U808 ( .A(n542), .B(n543), .Z(z3[322]) );
  NANDN U809 ( .A(N518), .B(z2[322]), .Z(n543) );
  NANDN U810 ( .A(n3), .B(N842), .Z(n542) );
  NAND U811 ( .A(n544), .B(n545), .Z(z3[321]) );
  NANDN U812 ( .A(N518), .B(z2[321]), .Z(n545) );
  NANDN U813 ( .A(n3), .B(N841), .Z(n544) );
  NAND U814 ( .A(n546), .B(n547), .Z(z3[320]) );
  NANDN U815 ( .A(N518), .B(z2[320]), .Z(n547) );
  NANDN U816 ( .A(n3), .B(N840), .Z(n546) );
  NAND U817 ( .A(n548), .B(n549), .Z(z3[31]) );
  NANDN U818 ( .A(N518), .B(z2[31]), .Z(n549) );
  NANDN U819 ( .A(n3), .B(N551), .Z(n548) );
  NAND U820 ( .A(n550), .B(n551), .Z(z3[319]) );
  NANDN U821 ( .A(N518), .B(z2[319]), .Z(n551) );
  NANDN U822 ( .A(n3), .B(N839), .Z(n550) );
  NAND U823 ( .A(n552), .B(n553), .Z(z3[318]) );
  NANDN U824 ( .A(N518), .B(z2[318]), .Z(n553) );
  NANDN U825 ( .A(n3), .B(N838), .Z(n552) );
  NAND U826 ( .A(n554), .B(n555), .Z(z3[317]) );
  NANDN U827 ( .A(N518), .B(z2[317]), .Z(n555) );
  NANDN U828 ( .A(n3), .B(N837), .Z(n554) );
  NAND U829 ( .A(n556), .B(n557), .Z(z3[316]) );
  NANDN U830 ( .A(N518), .B(z2[316]), .Z(n557) );
  NANDN U831 ( .A(n3), .B(N836), .Z(n556) );
  NAND U832 ( .A(n558), .B(n559), .Z(z3[315]) );
  NANDN U833 ( .A(N518), .B(z2[315]), .Z(n559) );
  NANDN U834 ( .A(n3), .B(N835), .Z(n558) );
  NAND U835 ( .A(n560), .B(n561), .Z(z3[314]) );
  NANDN U836 ( .A(N518), .B(z2[314]), .Z(n561) );
  NANDN U837 ( .A(n3), .B(N834), .Z(n560) );
  NAND U838 ( .A(n562), .B(n563), .Z(z3[313]) );
  NANDN U839 ( .A(N518), .B(z2[313]), .Z(n563) );
  NANDN U840 ( .A(n3), .B(N833), .Z(n562) );
  NAND U841 ( .A(n564), .B(n565), .Z(z3[312]) );
  NANDN U842 ( .A(N518), .B(z2[312]), .Z(n565) );
  NANDN U843 ( .A(n3), .B(N832), .Z(n564) );
  NAND U844 ( .A(n566), .B(n567), .Z(z3[311]) );
  NANDN U845 ( .A(N518), .B(z2[311]), .Z(n567) );
  NANDN U846 ( .A(n3), .B(N831), .Z(n566) );
  NAND U847 ( .A(n568), .B(n569), .Z(z3[310]) );
  NANDN U848 ( .A(N518), .B(z2[310]), .Z(n569) );
  NANDN U849 ( .A(n3), .B(N830), .Z(n568) );
  NAND U850 ( .A(n570), .B(n571), .Z(z3[30]) );
  NANDN U851 ( .A(N518), .B(z2[30]), .Z(n571) );
  NANDN U852 ( .A(n3), .B(N550), .Z(n570) );
  NAND U853 ( .A(n572), .B(n573), .Z(z3[309]) );
  NANDN U854 ( .A(N518), .B(z2[309]), .Z(n573) );
  NANDN U855 ( .A(n3), .B(N829), .Z(n572) );
  NAND U856 ( .A(n574), .B(n575), .Z(z3[308]) );
  NANDN U857 ( .A(N518), .B(z2[308]), .Z(n575) );
  NANDN U858 ( .A(n3), .B(N828), .Z(n574) );
  NAND U859 ( .A(n576), .B(n577), .Z(z3[307]) );
  NANDN U860 ( .A(N518), .B(z2[307]), .Z(n577) );
  NANDN U861 ( .A(n3), .B(N827), .Z(n576) );
  NAND U862 ( .A(n578), .B(n579), .Z(z3[306]) );
  NANDN U863 ( .A(N518), .B(z2[306]), .Z(n579) );
  NANDN U864 ( .A(n3), .B(N826), .Z(n578) );
  NAND U865 ( .A(n580), .B(n581), .Z(z3[305]) );
  NANDN U866 ( .A(N518), .B(z2[305]), .Z(n581) );
  NANDN U867 ( .A(n3), .B(N825), .Z(n580) );
  NAND U868 ( .A(n582), .B(n583), .Z(z3[304]) );
  NANDN U869 ( .A(N518), .B(z2[304]), .Z(n583) );
  NANDN U870 ( .A(n3), .B(N824), .Z(n582) );
  NAND U871 ( .A(n584), .B(n585), .Z(z3[303]) );
  NANDN U872 ( .A(N518), .B(z2[303]), .Z(n585) );
  NANDN U873 ( .A(n3), .B(N823), .Z(n584) );
  NAND U874 ( .A(n586), .B(n587), .Z(z3[302]) );
  NANDN U875 ( .A(N518), .B(z2[302]), .Z(n587) );
  NANDN U876 ( .A(n3), .B(N822), .Z(n586) );
  NAND U877 ( .A(n588), .B(n589), .Z(z3[301]) );
  NANDN U878 ( .A(N518), .B(z2[301]), .Z(n589) );
  NANDN U879 ( .A(n3), .B(N821), .Z(n588) );
  NAND U880 ( .A(n590), .B(n591), .Z(z3[300]) );
  NANDN U881 ( .A(N518), .B(z2[300]), .Z(n591) );
  NANDN U882 ( .A(n3), .B(N820), .Z(n590) );
  NAND U883 ( .A(n592), .B(n593), .Z(z3[2]) );
  NANDN U884 ( .A(N518), .B(z2[2]), .Z(n593) );
  NANDN U885 ( .A(n3), .B(N522), .Z(n592) );
  NAND U886 ( .A(n594), .B(n595), .Z(z3[29]) );
  NANDN U887 ( .A(N518), .B(z2[29]), .Z(n595) );
  NANDN U888 ( .A(n3), .B(N549), .Z(n594) );
  NAND U889 ( .A(n596), .B(n597), .Z(z3[299]) );
  NANDN U890 ( .A(N518), .B(z2[299]), .Z(n597) );
  NANDN U891 ( .A(n3), .B(N819), .Z(n596) );
  NAND U892 ( .A(n598), .B(n599), .Z(z3[298]) );
  NANDN U893 ( .A(N518), .B(z2[298]), .Z(n599) );
  NANDN U894 ( .A(n3), .B(N818), .Z(n598) );
  NAND U895 ( .A(n600), .B(n601), .Z(z3[297]) );
  NANDN U896 ( .A(N518), .B(z2[297]), .Z(n601) );
  NANDN U897 ( .A(n3), .B(N817), .Z(n600) );
  NAND U898 ( .A(n602), .B(n603), .Z(z3[296]) );
  NANDN U899 ( .A(N518), .B(z2[296]), .Z(n603) );
  NANDN U900 ( .A(n3), .B(N816), .Z(n602) );
  NAND U901 ( .A(n604), .B(n605), .Z(z3[295]) );
  NANDN U902 ( .A(N518), .B(z2[295]), .Z(n605) );
  NANDN U903 ( .A(n3), .B(N815), .Z(n604) );
  NAND U904 ( .A(n606), .B(n607), .Z(z3[294]) );
  NANDN U905 ( .A(N518), .B(z2[294]), .Z(n607) );
  NANDN U906 ( .A(n3), .B(N814), .Z(n606) );
  NAND U907 ( .A(n608), .B(n609), .Z(z3[293]) );
  NANDN U908 ( .A(N518), .B(z2[293]), .Z(n609) );
  NANDN U909 ( .A(n3), .B(N813), .Z(n608) );
  NAND U910 ( .A(n610), .B(n611), .Z(z3[292]) );
  NANDN U911 ( .A(N518), .B(z2[292]), .Z(n611) );
  NANDN U912 ( .A(n3), .B(N812), .Z(n610) );
  NAND U913 ( .A(n612), .B(n613), .Z(z3[291]) );
  NANDN U914 ( .A(N518), .B(z2[291]), .Z(n613) );
  NANDN U915 ( .A(n3), .B(N811), .Z(n612) );
  NAND U916 ( .A(n614), .B(n615), .Z(z3[290]) );
  NANDN U917 ( .A(N518), .B(z2[290]), .Z(n615) );
  NANDN U918 ( .A(n3), .B(N810), .Z(n614) );
  NAND U919 ( .A(n616), .B(n617), .Z(z3[28]) );
  NANDN U920 ( .A(N518), .B(z2[28]), .Z(n617) );
  NANDN U921 ( .A(n3), .B(N548), .Z(n616) );
  NAND U922 ( .A(n618), .B(n619), .Z(z3[289]) );
  NANDN U923 ( .A(N518), .B(z2[289]), .Z(n619) );
  NANDN U924 ( .A(n3), .B(N809), .Z(n618) );
  NAND U925 ( .A(n620), .B(n621), .Z(z3[288]) );
  NANDN U926 ( .A(N518), .B(z2[288]), .Z(n621) );
  NANDN U927 ( .A(n3), .B(N808), .Z(n620) );
  NAND U928 ( .A(n622), .B(n623), .Z(z3[287]) );
  NANDN U929 ( .A(N518), .B(z2[287]), .Z(n623) );
  NANDN U930 ( .A(n3), .B(N807), .Z(n622) );
  NAND U931 ( .A(n624), .B(n625), .Z(z3[286]) );
  NANDN U932 ( .A(N518), .B(z2[286]), .Z(n625) );
  NANDN U933 ( .A(n3), .B(N806), .Z(n624) );
  NAND U934 ( .A(n626), .B(n627), .Z(z3[285]) );
  NANDN U935 ( .A(N518), .B(z2[285]), .Z(n627) );
  NANDN U936 ( .A(n3), .B(N805), .Z(n626) );
  NAND U937 ( .A(n628), .B(n629), .Z(z3[284]) );
  NANDN U938 ( .A(N518), .B(z2[284]), .Z(n629) );
  NANDN U939 ( .A(n3), .B(N804), .Z(n628) );
  NAND U940 ( .A(n630), .B(n631), .Z(z3[283]) );
  NANDN U941 ( .A(N518), .B(z2[283]), .Z(n631) );
  NANDN U942 ( .A(n3), .B(N803), .Z(n630) );
  NAND U943 ( .A(n632), .B(n633), .Z(z3[282]) );
  NANDN U944 ( .A(N518), .B(z2[282]), .Z(n633) );
  NANDN U945 ( .A(n3), .B(N802), .Z(n632) );
  NAND U946 ( .A(n634), .B(n635), .Z(z3[281]) );
  NANDN U947 ( .A(N518), .B(z2[281]), .Z(n635) );
  NANDN U948 ( .A(n3), .B(N801), .Z(n634) );
  NAND U949 ( .A(n636), .B(n637), .Z(z3[280]) );
  NANDN U950 ( .A(N518), .B(z2[280]), .Z(n637) );
  NANDN U951 ( .A(n3), .B(N800), .Z(n636) );
  NAND U952 ( .A(n638), .B(n639), .Z(z3[27]) );
  NANDN U953 ( .A(N518), .B(z2[27]), .Z(n639) );
  NANDN U954 ( .A(n3), .B(N547), .Z(n638) );
  NAND U955 ( .A(n640), .B(n641), .Z(z3[279]) );
  NANDN U956 ( .A(N518), .B(z2[279]), .Z(n641) );
  NANDN U957 ( .A(n3), .B(N799), .Z(n640) );
  NAND U958 ( .A(n642), .B(n643), .Z(z3[278]) );
  NANDN U959 ( .A(N518), .B(z2[278]), .Z(n643) );
  NANDN U960 ( .A(n3), .B(N798), .Z(n642) );
  NAND U961 ( .A(n644), .B(n645), .Z(z3[277]) );
  NANDN U962 ( .A(N518), .B(z2[277]), .Z(n645) );
  NANDN U963 ( .A(n3), .B(N797), .Z(n644) );
  NAND U964 ( .A(n646), .B(n647), .Z(z3[276]) );
  NANDN U965 ( .A(N518), .B(z2[276]), .Z(n647) );
  NANDN U966 ( .A(n3), .B(N796), .Z(n646) );
  NAND U967 ( .A(n648), .B(n649), .Z(z3[275]) );
  NANDN U968 ( .A(N518), .B(z2[275]), .Z(n649) );
  NANDN U969 ( .A(n3), .B(N795), .Z(n648) );
  NAND U970 ( .A(n650), .B(n651), .Z(z3[274]) );
  NANDN U971 ( .A(N518), .B(z2[274]), .Z(n651) );
  NANDN U972 ( .A(n3), .B(N794), .Z(n650) );
  NAND U973 ( .A(n652), .B(n653), .Z(z3[273]) );
  NANDN U974 ( .A(N518), .B(z2[273]), .Z(n653) );
  NANDN U975 ( .A(n3), .B(N793), .Z(n652) );
  NAND U976 ( .A(n654), .B(n655), .Z(z3[272]) );
  NANDN U977 ( .A(N518), .B(z2[272]), .Z(n655) );
  NANDN U978 ( .A(n3), .B(N792), .Z(n654) );
  NAND U979 ( .A(n656), .B(n657), .Z(z3[271]) );
  NANDN U980 ( .A(N518), .B(z2[271]), .Z(n657) );
  NANDN U981 ( .A(n3), .B(N791), .Z(n656) );
  NAND U982 ( .A(n658), .B(n659), .Z(z3[270]) );
  NANDN U983 ( .A(N518), .B(z2[270]), .Z(n659) );
  NANDN U984 ( .A(n3), .B(N790), .Z(n658) );
  NAND U985 ( .A(n660), .B(n661), .Z(z3[26]) );
  NANDN U986 ( .A(N518), .B(z2[26]), .Z(n661) );
  NANDN U987 ( .A(n3), .B(N546), .Z(n660) );
  NAND U988 ( .A(n662), .B(n663), .Z(z3[269]) );
  NANDN U989 ( .A(N518), .B(z2[269]), .Z(n663) );
  NANDN U990 ( .A(n3), .B(N789), .Z(n662) );
  NAND U991 ( .A(n664), .B(n665), .Z(z3[268]) );
  NANDN U992 ( .A(N518), .B(z2[268]), .Z(n665) );
  NANDN U993 ( .A(n3), .B(N788), .Z(n664) );
  NAND U994 ( .A(n666), .B(n667), .Z(z3[267]) );
  NANDN U995 ( .A(N518), .B(z2[267]), .Z(n667) );
  NANDN U996 ( .A(n3), .B(N787), .Z(n666) );
  NAND U997 ( .A(n668), .B(n669), .Z(z3[266]) );
  NANDN U998 ( .A(N518), .B(z2[266]), .Z(n669) );
  NANDN U999 ( .A(n3), .B(N786), .Z(n668) );
  NAND U1000 ( .A(n670), .B(n671), .Z(z3[265]) );
  NANDN U1001 ( .A(N518), .B(z2[265]), .Z(n671) );
  NANDN U1002 ( .A(n3), .B(N785), .Z(n670) );
  NAND U1003 ( .A(n672), .B(n673), .Z(z3[264]) );
  NANDN U1004 ( .A(N518), .B(z2[264]), .Z(n673) );
  NANDN U1005 ( .A(n3), .B(N784), .Z(n672) );
  NAND U1006 ( .A(n674), .B(n675), .Z(z3[263]) );
  NANDN U1007 ( .A(N518), .B(z2[263]), .Z(n675) );
  NANDN U1008 ( .A(n3), .B(N783), .Z(n674) );
  NAND U1009 ( .A(n676), .B(n677), .Z(z3[262]) );
  NANDN U1010 ( .A(N518), .B(z2[262]), .Z(n677) );
  NANDN U1011 ( .A(n3), .B(N782), .Z(n676) );
  NAND U1012 ( .A(n678), .B(n679), .Z(z3[261]) );
  NANDN U1013 ( .A(N518), .B(z2[261]), .Z(n679) );
  NANDN U1014 ( .A(n3), .B(N781), .Z(n678) );
  NAND U1015 ( .A(n680), .B(n681), .Z(z3[260]) );
  NANDN U1016 ( .A(N518), .B(z2[260]), .Z(n681) );
  NANDN U1017 ( .A(n3), .B(N780), .Z(n680) );
  NAND U1018 ( .A(n682), .B(n683), .Z(z3[25]) );
  NANDN U1019 ( .A(N518), .B(z2[25]), .Z(n683) );
  NANDN U1020 ( .A(n3), .B(N545), .Z(n682) );
  NAND U1021 ( .A(n684), .B(n685), .Z(z3[259]) );
  NANDN U1022 ( .A(N518), .B(z2[259]), .Z(n685) );
  NANDN U1023 ( .A(n3), .B(N779), .Z(n684) );
  NAND U1024 ( .A(n686), .B(n687), .Z(z3[258]) );
  NANDN U1025 ( .A(N518), .B(z2[258]), .Z(n687) );
  NANDN U1026 ( .A(n3), .B(N778), .Z(n686) );
  NAND U1027 ( .A(n688), .B(n689), .Z(z3[257]) );
  NANDN U1028 ( .A(N518), .B(z2[257]), .Z(n689) );
  NANDN U1029 ( .A(n3), .B(N777), .Z(n688) );
  NAND U1030 ( .A(n690), .B(n691), .Z(z3[256]) );
  NANDN U1031 ( .A(N518), .B(z2[256]), .Z(n691) );
  NANDN U1032 ( .A(n3), .B(N776), .Z(n690) );
  NAND U1033 ( .A(n692), .B(n693), .Z(z3[255]) );
  NANDN U1034 ( .A(N518), .B(z2[255]), .Z(n693) );
  NANDN U1035 ( .A(n3), .B(N775), .Z(n692) );
  NAND U1036 ( .A(n694), .B(n695), .Z(z3[254]) );
  NANDN U1037 ( .A(N518), .B(z2[254]), .Z(n695) );
  NANDN U1038 ( .A(n3), .B(N774), .Z(n694) );
  NAND U1039 ( .A(n696), .B(n697), .Z(z3[253]) );
  NANDN U1040 ( .A(N518), .B(z2[253]), .Z(n697) );
  NANDN U1041 ( .A(n3), .B(N773), .Z(n696) );
  NAND U1042 ( .A(n698), .B(n699), .Z(z3[252]) );
  NANDN U1043 ( .A(N518), .B(z2[252]), .Z(n699) );
  NANDN U1044 ( .A(n3), .B(N772), .Z(n698) );
  NAND U1045 ( .A(n700), .B(n701), .Z(z3[251]) );
  NANDN U1046 ( .A(N518), .B(z2[251]), .Z(n701) );
  NANDN U1047 ( .A(n3), .B(N771), .Z(n700) );
  NAND U1048 ( .A(n702), .B(n703), .Z(z3[250]) );
  NANDN U1049 ( .A(N518), .B(z2[250]), .Z(n703) );
  NANDN U1050 ( .A(n3), .B(N770), .Z(n702) );
  NAND U1051 ( .A(n704), .B(n705), .Z(z3[24]) );
  NANDN U1052 ( .A(N518), .B(z2[24]), .Z(n705) );
  NANDN U1053 ( .A(n3), .B(N544), .Z(n704) );
  NAND U1054 ( .A(n706), .B(n707), .Z(z3[249]) );
  NANDN U1055 ( .A(N518), .B(z2[249]), .Z(n707) );
  NANDN U1056 ( .A(n3), .B(N769), .Z(n706) );
  NAND U1057 ( .A(n708), .B(n709), .Z(z3[248]) );
  NANDN U1058 ( .A(N518), .B(z2[248]), .Z(n709) );
  NANDN U1059 ( .A(n3), .B(N768), .Z(n708) );
  NAND U1060 ( .A(n710), .B(n711), .Z(z3[247]) );
  NANDN U1061 ( .A(N518), .B(z2[247]), .Z(n711) );
  NANDN U1062 ( .A(n3), .B(N767), .Z(n710) );
  NAND U1063 ( .A(n712), .B(n713), .Z(z3[246]) );
  NANDN U1064 ( .A(N518), .B(z2[246]), .Z(n713) );
  NANDN U1065 ( .A(n3), .B(N766), .Z(n712) );
  NAND U1066 ( .A(n714), .B(n715), .Z(z3[245]) );
  NANDN U1067 ( .A(N518), .B(z2[245]), .Z(n715) );
  NANDN U1068 ( .A(n3), .B(N765), .Z(n714) );
  NAND U1069 ( .A(n716), .B(n717), .Z(z3[244]) );
  NANDN U1070 ( .A(N518), .B(z2[244]), .Z(n717) );
  NANDN U1071 ( .A(n3), .B(N764), .Z(n716) );
  NAND U1072 ( .A(n718), .B(n719), .Z(z3[243]) );
  NANDN U1073 ( .A(N518), .B(z2[243]), .Z(n719) );
  NANDN U1074 ( .A(n3), .B(N763), .Z(n718) );
  NAND U1075 ( .A(n720), .B(n721), .Z(z3[242]) );
  NANDN U1076 ( .A(N518), .B(z2[242]), .Z(n721) );
  NANDN U1077 ( .A(n3), .B(N762), .Z(n720) );
  NAND U1078 ( .A(n722), .B(n723), .Z(z3[241]) );
  NANDN U1079 ( .A(N518), .B(z2[241]), .Z(n723) );
  NANDN U1080 ( .A(n3), .B(N761), .Z(n722) );
  NAND U1081 ( .A(n724), .B(n725), .Z(z3[240]) );
  NANDN U1082 ( .A(N518), .B(z2[240]), .Z(n725) );
  NANDN U1083 ( .A(n3), .B(N760), .Z(n724) );
  NAND U1084 ( .A(n726), .B(n727), .Z(z3[23]) );
  NANDN U1085 ( .A(N518), .B(z2[23]), .Z(n727) );
  NANDN U1086 ( .A(n3), .B(N543), .Z(n726) );
  NAND U1087 ( .A(n728), .B(n729), .Z(z3[239]) );
  NANDN U1088 ( .A(N518), .B(z2[239]), .Z(n729) );
  NANDN U1089 ( .A(n3), .B(N759), .Z(n728) );
  NAND U1090 ( .A(n730), .B(n731), .Z(z3[238]) );
  NANDN U1091 ( .A(N518), .B(z2[238]), .Z(n731) );
  NANDN U1092 ( .A(n3), .B(N758), .Z(n730) );
  NAND U1093 ( .A(n732), .B(n733), .Z(z3[237]) );
  NANDN U1094 ( .A(N518), .B(z2[237]), .Z(n733) );
  NANDN U1095 ( .A(n3), .B(N757), .Z(n732) );
  NAND U1096 ( .A(n734), .B(n735), .Z(z3[236]) );
  NANDN U1097 ( .A(N518), .B(z2[236]), .Z(n735) );
  NANDN U1098 ( .A(n3), .B(N756), .Z(n734) );
  NAND U1099 ( .A(n736), .B(n737), .Z(z3[235]) );
  NANDN U1100 ( .A(N518), .B(z2[235]), .Z(n737) );
  NANDN U1101 ( .A(n3), .B(N755), .Z(n736) );
  NAND U1102 ( .A(n738), .B(n739), .Z(z3[234]) );
  NANDN U1103 ( .A(N518), .B(z2[234]), .Z(n739) );
  NANDN U1104 ( .A(n3), .B(N754), .Z(n738) );
  NAND U1105 ( .A(n740), .B(n741), .Z(z3[233]) );
  NANDN U1106 ( .A(N518), .B(z2[233]), .Z(n741) );
  NANDN U1107 ( .A(n3), .B(N753), .Z(n740) );
  NAND U1108 ( .A(n742), .B(n743), .Z(z3[232]) );
  NANDN U1109 ( .A(N518), .B(z2[232]), .Z(n743) );
  NANDN U1110 ( .A(n3), .B(N752), .Z(n742) );
  NAND U1111 ( .A(n744), .B(n745), .Z(z3[231]) );
  NANDN U1112 ( .A(N518), .B(z2[231]), .Z(n745) );
  NANDN U1113 ( .A(n3), .B(N751), .Z(n744) );
  NAND U1114 ( .A(n746), .B(n747), .Z(z3[230]) );
  NANDN U1115 ( .A(N518), .B(z2[230]), .Z(n747) );
  NANDN U1116 ( .A(n3), .B(N750), .Z(n746) );
  NAND U1117 ( .A(n748), .B(n749), .Z(z3[22]) );
  NANDN U1118 ( .A(N518), .B(z2[22]), .Z(n749) );
  NANDN U1119 ( .A(n3), .B(N542), .Z(n748) );
  NAND U1120 ( .A(n750), .B(n751), .Z(z3[229]) );
  NANDN U1121 ( .A(N518), .B(z2[229]), .Z(n751) );
  NANDN U1122 ( .A(n3), .B(N749), .Z(n750) );
  NAND U1123 ( .A(n752), .B(n753), .Z(z3[228]) );
  NANDN U1124 ( .A(N518), .B(z2[228]), .Z(n753) );
  NANDN U1125 ( .A(n3), .B(N748), .Z(n752) );
  NAND U1126 ( .A(n754), .B(n755), .Z(z3[227]) );
  NANDN U1127 ( .A(N518), .B(z2[227]), .Z(n755) );
  NANDN U1128 ( .A(n3), .B(N747), .Z(n754) );
  NAND U1129 ( .A(n756), .B(n757), .Z(z3[226]) );
  NANDN U1130 ( .A(N518), .B(z2[226]), .Z(n757) );
  NANDN U1131 ( .A(n3), .B(N746), .Z(n756) );
  NAND U1132 ( .A(n758), .B(n759), .Z(z3[225]) );
  NANDN U1133 ( .A(N518), .B(z2[225]), .Z(n759) );
  NANDN U1134 ( .A(n3), .B(N745), .Z(n758) );
  NAND U1135 ( .A(n760), .B(n761), .Z(z3[224]) );
  NANDN U1136 ( .A(N518), .B(z2[224]), .Z(n761) );
  NANDN U1137 ( .A(n3), .B(N744), .Z(n760) );
  NAND U1138 ( .A(n762), .B(n763), .Z(z3[223]) );
  NANDN U1139 ( .A(N518), .B(z2[223]), .Z(n763) );
  NANDN U1140 ( .A(n3), .B(N743), .Z(n762) );
  NAND U1141 ( .A(n764), .B(n765), .Z(z3[222]) );
  NANDN U1142 ( .A(N518), .B(z2[222]), .Z(n765) );
  NANDN U1143 ( .A(n3), .B(N742), .Z(n764) );
  NAND U1144 ( .A(n766), .B(n767), .Z(z3[221]) );
  NANDN U1145 ( .A(N518), .B(z2[221]), .Z(n767) );
  NANDN U1146 ( .A(n3), .B(N741), .Z(n766) );
  NAND U1147 ( .A(n768), .B(n769), .Z(z3[220]) );
  NANDN U1148 ( .A(N518), .B(z2[220]), .Z(n769) );
  NANDN U1149 ( .A(n3), .B(N740), .Z(n768) );
  NAND U1150 ( .A(n770), .B(n771), .Z(z3[21]) );
  NANDN U1151 ( .A(N518), .B(z2[21]), .Z(n771) );
  NANDN U1152 ( .A(n3), .B(N541), .Z(n770) );
  NAND U1153 ( .A(n772), .B(n773), .Z(z3[219]) );
  NANDN U1154 ( .A(N518), .B(z2[219]), .Z(n773) );
  NANDN U1155 ( .A(n3), .B(N739), .Z(n772) );
  NAND U1156 ( .A(n774), .B(n775), .Z(z3[218]) );
  NANDN U1157 ( .A(N518), .B(z2[218]), .Z(n775) );
  NANDN U1158 ( .A(n3), .B(N738), .Z(n774) );
  NAND U1159 ( .A(n776), .B(n777), .Z(z3[217]) );
  NANDN U1160 ( .A(N518), .B(z2[217]), .Z(n777) );
  NANDN U1161 ( .A(n3), .B(N737), .Z(n776) );
  NAND U1162 ( .A(n778), .B(n779), .Z(z3[216]) );
  NANDN U1163 ( .A(N518), .B(z2[216]), .Z(n779) );
  NANDN U1164 ( .A(n3), .B(N736), .Z(n778) );
  NAND U1165 ( .A(n780), .B(n781), .Z(z3[215]) );
  NANDN U1166 ( .A(N518), .B(z2[215]), .Z(n781) );
  NANDN U1167 ( .A(n3), .B(N735), .Z(n780) );
  NAND U1168 ( .A(n782), .B(n783), .Z(z3[214]) );
  NANDN U1169 ( .A(N518), .B(z2[214]), .Z(n783) );
  NANDN U1170 ( .A(n3), .B(N734), .Z(n782) );
  NAND U1171 ( .A(n784), .B(n785), .Z(z3[213]) );
  NANDN U1172 ( .A(N518), .B(z2[213]), .Z(n785) );
  NANDN U1173 ( .A(n3), .B(N733), .Z(n784) );
  NAND U1174 ( .A(n786), .B(n787), .Z(z3[212]) );
  NANDN U1175 ( .A(N518), .B(z2[212]), .Z(n787) );
  NANDN U1176 ( .A(n3), .B(N732), .Z(n786) );
  NAND U1177 ( .A(n788), .B(n789), .Z(z3[211]) );
  NANDN U1178 ( .A(N518), .B(z2[211]), .Z(n789) );
  NANDN U1179 ( .A(n3), .B(N731), .Z(n788) );
  NAND U1180 ( .A(n790), .B(n791), .Z(z3[210]) );
  NANDN U1181 ( .A(N518), .B(z2[210]), .Z(n791) );
  NANDN U1182 ( .A(n3), .B(N730), .Z(n790) );
  NAND U1183 ( .A(n792), .B(n793), .Z(z3[20]) );
  NANDN U1184 ( .A(N518), .B(z2[20]), .Z(n793) );
  NANDN U1185 ( .A(n3), .B(N540), .Z(n792) );
  NAND U1186 ( .A(n794), .B(n795), .Z(z3[209]) );
  NANDN U1187 ( .A(N518), .B(z2[209]), .Z(n795) );
  NANDN U1188 ( .A(n3), .B(N729), .Z(n794) );
  NAND U1189 ( .A(n796), .B(n797), .Z(z3[208]) );
  NANDN U1190 ( .A(N518), .B(z2[208]), .Z(n797) );
  NANDN U1191 ( .A(n3), .B(N728), .Z(n796) );
  NAND U1192 ( .A(n798), .B(n799), .Z(z3[207]) );
  NANDN U1193 ( .A(N518), .B(z2[207]), .Z(n799) );
  NANDN U1194 ( .A(n3), .B(N727), .Z(n798) );
  NAND U1195 ( .A(n800), .B(n801), .Z(z3[206]) );
  NANDN U1196 ( .A(N518), .B(z2[206]), .Z(n801) );
  NANDN U1197 ( .A(n3), .B(N726), .Z(n800) );
  NAND U1198 ( .A(n802), .B(n803), .Z(z3[205]) );
  NANDN U1199 ( .A(N518), .B(z2[205]), .Z(n803) );
  NANDN U1200 ( .A(n3), .B(N725), .Z(n802) );
  NAND U1201 ( .A(n804), .B(n805), .Z(z3[204]) );
  NANDN U1202 ( .A(N518), .B(z2[204]), .Z(n805) );
  NANDN U1203 ( .A(n3), .B(N724), .Z(n804) );
  NAND U1204 ( .A(n806), .B(n807), .Z(z3[203]) );
  NANDN U1205 ( .A(N518), .B(z2[203]), .Z(n807) );
  NANDN U1206 ( .A(n3), .B(N723), .Z(n806) );
  NAND U1207 ( .A(n808), .B(n809), .Z(z3[202]) );
  NANDN U1208 ( .A(N518), .B(z2[202]), .Z(n809) );
  NANDN U1209 ( .A(n3), .B(N722), .Z(n808) );
  NAND U1210 ( .A(n810), .B(n811), .Z(z3[201]) );
  NANDN U1211 ( .A(N518), .B(z2[201]), .Z(n811) );
  NANDN U1212 ( .A(n3), .B(N721), .Z(n810) );
  NAND U1213 ( .A(n812), .B(n813), .Z(z3[200]) );
  NANDN U1214 ( .A(N518), .B(z2[200]), .Z(n813) );
  NANDN U1215 ( .A(n3), .B(N720), .Z(n812) );
  NAND U1216 ( .A(n814), .B(n815), .Z(z3[1]) );
  NANDN U1217 ( .A(N518), .B(z2[1]), .Z(n815) );
  NANDN U1218 ( .A(n3), .B(N521), .Z(n814) );
  NAND U1219 ( .A(n816), .B(n817), .Z(z3[19]) );
  NANDN U1220 ( .A(N518), .B(z2[19]), .Z(n817) );
  NANDN U1221 ( .A(n3), .B(N539), .Z(n816) );
  NAND U1222 ( .A(n818), .B(n819), .Z(z3[199]) );
  NANDN U1223 ( .A(N518), .B(z2[199]), .Z(n819) );
  NANDN U1224 ( .A(n3), .B(N719), .Z(n818) );
  NAND U1225 ( .A(n820), .B(n821), .Z(z3[198]) );
  NANDN U1226 ( .A(N518), .B(z2[198]), .Z(n821) );
  NANDN U1227 ( .A(n3), .B(N718), .Z(n820) );
  NAND U1228 ( .A(n822), .B(n823), .Z(z3[197]) );
  NANDN U1229 ( .A(N518), .B(z2[197]), .Z(n823) );
  NANDN U1230 ( .A(n3), .B(N717), .Z(n822) );
  NAND U1231 ( .A(n824), .B(n825), .Z(z3[196]) );
  NANDN U1232 ( .A(N518), .B(z2[196]), .Z(n825) );
  NANDN U1233 ( .A(n3), .B(N716), .Z(n824) );
  NAND U1234 ( .A(n826), .B(n827), .Z(z3[195]) );
  NANDN U1235 ( .A(N518), .B(z2[195]), .Z(n827) );
  NANDN U1236 ( .A(n3), .B(N715), .Z(n826) );
  NAND U1237 ( .A(n828), .B(n829), .Z(z3[194]) );
  NANDN U1238 ( .A(N518), .B(z2[194]), .Z(n829) );
  NANDN U1239 ( .A(n3), .B(N714), .Z(n828) );
  NAND U1240 ( .A(n830), .B(n831), .Z(z3[193]) );
  NANDN U1241 ( .A(N518), .B(z2[193]), .Z(n831) );
  NANDN U1242 ( .A(n3), .B(N713), .Z(n830) );
  NAND U1243 ( .A(n832), .B(n833), .Z(z3[192]) );
  NANDN U1244 ( .A(N518), .B(z2[192]), .Z(n833) );
  NANDN U1245 ( .A(n3), .B(N712), .Z(n832) );
  NAND U1246 ( .A(n834), .B(n835), .Z(z3[191]) );
  NANDN U1247 ( .A(N518), .B(z2[191]), .Z(n835) );
  NANDN U1248 ( .A(n3), .B(N711), .Z(n834) );
  NAND U1249 ( .A(n836), .B(n837), .Z(z3[190]) );
  NANDN U1250 ( .A(N518), .B(z2[190]), .Z(n837) );
  NANDN U1251 ( .A(n3), .B(N710), .Z(n836) );
  NAND U1252 ( .A(n838), .B(n839), .Z(z3[18]) );
  NANDN U1253 ( .A(N518), .B(z2[18]), .Z(n839) );
  NANDN U1254 ( .A(n3), .B(N538), .Z(n838) );
  NAND U1255 ( .A(n840), .B(n841), .Z(z3[189]) );
  NANDN U1256 ( .A(N518), .B(z2[189]), .Z(n841) );
  NANDN U1257 ( .A(n3), .B(N709), .Z(n840) );
  NAND U1258 ( .A(n842), .B(n843), .Z(z3[188]) );
  NANDN U1259 ( .A(N518), .B(z2[188]), .Z(n843) );
  NANDN U1260 ( .A(n3), .B(N708), .Z(n842) );
  NAND U1261 ( .A(n844), .B(n845), .Z(z3[187]) );
  NANDN U1262 ( .A(N518), .B(z2[187]), .Z(n845) );
  NANDN U1263 ( .A(n3), .B(N707), .Z(n844) );
  NAND U1264 ( .A(n846), .B(n847), .Z(z3[186]) );
  NANDN U1265 ( .A(N518), .B(z2[186]), .Z(n847) );
  NANDN U1266 ( .A(n3), .B(N706), .Z(n846) );
  NAND U1267 ( .A(n848), .B(n849), .Z(z3[185]) );
  NANDN U1268 ( .A(N518), .B(z2[185]), .Z(n849) );
  NANDN U1269 ( .A(n3), .B(N705), .Z(n848) );
  NAND U1270 ( .A(n850), .B(n851), .Z(z3[184]) );
  NANDN U1271 ( .A(N518), .B(z2[184]), .Z(n851) );
  NANDN U1272 ( .A(n3), .B(N704), .Z(n850) );
  NAND U1273 ( .A(n852), .B(n853), .Z(z3[183]) );
  NANDN U1274 ( .A(N518), .B(z2[183]), .Z(n853) );
  NANDN U1275 ( .A(n3), .B(N703), .Z(n852) );
  NAND U1276 ( .A(n854), .B(n855), .Z(z3[182]) );
  NANDN U1277 ( .A(N518), .B(z2[182]), .Z(n855) );
  NANDN U1278 ( .A(n3), .B(N702), .Z(n854) );
  NAND U1279 ( .A(n856), .B(n857), .Z(z3[181]) );
  NANDN U1280 ( .A(N518), .B(z2[181]), .Z(n857) );
  NANDN U1281 ( .A(n3), .B(N701), .Z(n856) );
  NAND U1282 ( .A(n858), .B(n859), .Z(z3[180]) );
  NANDN U1283 ( .A(N518), .B(z2[180]), .Z(n859) );
  NANDN U1284 ( .A(n3), .B(N700), .Z(n858) );
  NAND U1285 ( .A(n860), .B(n861), .Z(z3[17]) );
  NANDN U1286 ( .A(N518), .B(z2[17]), .Z(n861) );
  NANDN U1287 ( .A(n3), .B(N537), .Z(n860) );
  NAND U1288 ( .A(n862), .B(n863), .Z(z3[179]) );
  NANDN U1289 ( .A(N518), .B(z2[179]), .Z(n863) );
  NANDN U1290 ( .A(n3), .B(N699), .Z(n862) );
  NAND U1291 ( .A(n864), .B(n865), .Z(z3[178]) );
  NANDN U1292 ( .A(N518), .B(z2[178]), .Z(n865) );
  NANDN U1293 ( .A(n3), .B(N698), .Z(n864) );
  NAND U1294 ( .A(n866), .B(n867), .Z(z3[177]) );
  NANDN U1295 ( .A(N518), .B(z2[177]), .Z(n867) );
  NANDN U1296 ( .A(n3), .B(N697), .Z(n866) );
  NAND U1297 ( .A(n868), .B(n869), .Z(z3[176]) );
  NANDN U1298 ( .A(N518), .B(z2[176]), .Z(n869) );
  NANDN U1299 ( .A(n3), .B(N696), .Z(n868) );
  NAND U1300 ( .A(n870), .B(n871), .Z(z3[175]) );
  NANDN U1301 ( .A(N518), .B(z2[175]), .Z(n871) );
  NANDN U1302 ( .A(n3), .B(N695), .Z(n870) );
  NAND U1303 ( .A(n872), .B(n873), .Z(z3[174]) );
  NANDN U1304 ( .A(N518), .B(z2[174]), .Z(n873) );
  NANDN U1305 ( .A(n3), .B(N694), .Z(n872) );
  NAND U1306 ( .A(n874), .B(n875), .Z(z3[173]) );
  NANDN U1307 ( .A(N518), .B(z2[173]), .Z(n875) );
  NANDN U1308 ( .A(n3), .B(N693), .Z(n874) );
  NAND U1309 ( .A(n876), .B(n877), .Z(z3[172]) );
  NANDN U1310 ( .A(N518), .B(z2[172]), .Z(n877) );
  NANDN U1311 ( .A(n3), .B(N692), .Z(n876) );
  NAND U1312 ( .A(n878), .B(n879), .Z(z3[171]) );
  NANDN U1313 ( .A(N518), .B(z2[171]), .Z(n879) );
  NANDN U1314 ( .A(n3), .B(N691), .Z(n878) );
  NAND U1315 ( .A(n880), .B(n881), .Z(z3[170]) );
  NANDN U1316 ( .A(N518), .B(z2[170]), .Z(n881) );
  NANDN U1317 ( .A(n3), .B(N690), .Z(n880) );
  NAND U1318 ( .A(n882), .B(n883), .Z(z3[16]) );
  NANDN U1319 ( .A(N518), .B(z2[16]), .Z(n883) );
  NANDN U1320 ( .A(n3), .B(N536), .Z(n882) );
  NAND U1321 ( .A(n884), .B(n885), .Z(z3[169]) );
  NANDN U1322 ( .A(N518), .B(z2[169]), .Z(n885) );
  NANDN U1323 ( .A(n3), .B(N689), .Z(n884) );
  NAND U1324 ( .A(n886), .B(n887), .Z(z3[168]) );
  NANDN U1325 ( .A(N518), .B(z2[168]), .Z(n887) );
  NANDN U1326 ( .A(n3), .B(N688), .Z(n886) );
  NAND U1327 ( .A(n888), .B(n889), .Z(z3[167]) );
  NANDN U1328 ( .A(N518), .B(z2[167]), .Z(n889) );
  NANDN U1329 ( .A(n3), .B(N687), .Z(n888) );
  NAND U1330 ( .A(n890), .B(n891), .Z(z3[166]) );
  NANDN U1331 ( .A(N518), .B(z2[166]), .Z(n891) );
  NANDN U1332 ( .A(n3), .B(N686), .Z(n890) );
  NAND U1333 ( .A(n892), .B(n893), .Z(z3[165]) );
  NANDN U1334 ( .A(N518), .B(z2[165]), .Z(n893) );
  NANDN U1335 ( .A(n3), .B(N685), .Z(n892) );
  NAND U1336 ( .A(n894), .B(n895), .Z(z3[164]) );
  NANDN U1337 ( .A(N518), .B(z2[164]), .Z(n895) );
  NANDN U1338 ( .A(n3), .B(N684), .Z(n894) );
  NAND U1339 ( .A(n896), .B(n897), .Z(z3[163]) );
  NANDN U1340 ( .A(N518), .B(z2[163]), .Z(n897) );
  NANDN U1341 ( .A(n3), .B(N683), .Z(n896) );
  NAND U1342 ( .A(n898), .B(n899), .Z(z3[162]) );
  NANDN U1343 ( .A(N518), .B(z2[162]), .Z(n899) );
  NANDN U1344 ( .A(n3), .B(N682), .Z(n898) );
  NAND U1345 ( .A(n900), .B(n901), .Z(z3[161]) );
  NANDN U1346 ( .A(N518), .B(z2[161]), .Z(n901) );
  NANDN U1347 ( .A(n3), .B(N681), .Z(n900) );
  NAND U1348 ( .A(n902), .B(n903), .Z(z3[160]) );
  NANDN U1349 ( .A(N518), .B(z2[160]), .Z(n903) );
  NANDN U1350 ( .A(n3), .B(N680), .Z(n902) );
  NAND U1351 ( .A(n904), .B(n905), .Z(z3[15]) );
  NANDN U1352 ( .A(N518), .B(z2[15]), .Z(n905) );
  NANDN U1353 ( .A(n3), .B(N535), .Z(n904) );
  NAND U1354 ( .A(n906), .B(n907), .Z(z3[159]) );
  NANDN U1355 ( .A(N518), .B(z2[159]), .Z(n907) );
  NANDN U1356 ( .A(n3), .B(N679), .Z(n906) );
  NAND U1357 ( .A(n908), .B(n909), .Z(z3[158]) );
  NANDN U1358 ( .A(N518), .B(z2[158]), .Z(n909) );
  NANDN U1359 ( .A(n3), .B(N678), .Z(n908) );
  NAND U1360 ( .A(n910), .B(n911), .Z(z3[157]) );
  NANDN U1361 ( .A(N518), .B(z2[157]), .Z(n911) );
  NANDN U1362 ( .A(n3), .B(N677), .Z(n910) );
  NAND U1363 ( .A(n912), .B(n913), .Z(z3[156]) );
  NANDN U1364 ( .A(N518), .B(z2[156]), .Z(n913) );
  NANDN U1365 ( .A(n3), .B(N676), .Z(n912) );
  NAND U1366 ( .A(n914), .B(n915), .Z(z3[155]) );
  NANDN U1367 ( .A(N518), .B(z2[155]), .Z(n915) );
  NANDN U1368 ( .A(n3), .B(N675), .Z(n914) );
  NAND U1369 ( .A(n916), .B(n917), .Z(z3[154]) );
  NANDN U1370 ( .A(N518), .B(z2[154]), .Z(n917) );
  NANDN U1371 ( .A(n3), .B(N674), .Z(n916) );
  NAND U1372 ( .A(n918), .B(n919), .Z(z3[153]) );
  NANDN U1373 ( .A(N518), .B(z2[153]), .Z(n919) );
  NANDN U1374 ( .A(n3), .B(N673), .Z(n918) );
  NAND U1375 ( .A(n920), .B(n921), .Z(z3[152]) );
  NANDN U1376 ( .A(N518), .B(z2[152]), .Z(n921) );
  NANDN U1377 ( .A(n3), .B(N672), .Z(n920) );
  NAND U1378 ( .A(n922), .B(n923), .Z(z3[151]) );
  NANDN U1379 ( .A(N518), .B(z2[151]), .Z(n923) );
  NANDN U1380 ( .A(n3), .B(N671), .Z(n922) );
  NAND U1381 ( .A(n924), .B(n925), .Z(z3[150]) );
  NANDN U1382 ( .A(N518), .B(z2[150]), .Z(n925) );
  NANDN U1383 ( .A(n3), .B(N670), .Z(n924) );
  NAND U1384 ( .A(n926), .B(n927), .Z(z3[14]) );
  NANDN U1385 ( .A(N518), .B(z2[14]), .Z(n927) );
  NANDN U1386 ( .A(n3), .B(N534), .Z(n926) );
  NAND U1387 ( .A(n928), .B(n929), .Z(z3[149]) );
  NANDN U1388 ( .A(N518), .B(z2[149]), .Z(n929) );
  NANDN U1389 ( .A(n3), .B(N669), .Z(n928) );
  NAND U1390 ( .A(n930), .B(n931), .Z(z3[148]) );
  NANDN U1391 ( .A(N518), .B(z2[148]), .Z(n931) );
  NANDN U1392 ( .A(n3), .B(N668), .Z(n930) );
  NAND U1393 ( .A(n932), .B(n933), .Z(z3[147]) );
  NANDN U1394 ( .A(N518), .B(z2[147]), .Z(n933) );
  NANDN U1395 ( .A(n3), .B(N667), .Z(n932) );
  NAND U1396 ( .A(n934), .B(n935), .Z(z3[146]) );
  NANDN U1397 ( .A(N518), .B(z2[146]), .Z(n935) );
  NANDN U1398 ( .A(n3), .B(N666), .Z(n934) );
  NAND U1399 ( .A(n936), .B(n937), .Z(z3[145]) );
  NANDN U1400 ( .A(N518), .B(z2[145]), .Z(n937) );
  NANDN U1401 ( .A(n3), .B(N665), .Z(n936) );
  NAND U1402 ( .A(n938), .B(n939), .Z(z3[144]) );
  NANDN U1403 ( .A(N518), .B(z2[144]), .Z(n939) );
  NANDN U1404 ( .A(n3), .B(N664), .Z(n938) );
  NAND U1405 ( .A(n940), .B(n941), .Z(z3[143]) );
  NANDN U1406 ( .A(N518), .B(z2[143]), .Z(n941) );
  NANDN U1407 ( .A(n3), .B(N663), .Z(n940) );
  NAND U1408 ( .A(n942), .B(n943), .Z(z3[142]) );
  NANDN U1409 ( .A(N518), .B(z2[142]), .Z(n943) );
  NANDN U1410 ( .A(n3), .B(N662), .Z(n942) );
  NAND U1411 ( .A(n944), .B(n945), .Z(z3[141]) );
  NANDN U1412 ( .A(N518), .B(z2[141]), .Z(n945) );
  NANDN U1413 ( .A(n3), .B(N661), .Z(n944) );
  NAND U1414 ( .A(n946), .B(n947), .Z(z3[140]) );
  NANDN U1415 ( .A(N518), .B(z2[140]), .Z(n947) );
  NANDN U1416 ( .A(n3), .B(N660), .Z(n946) );
  NAND U1417 ( .A(n948), .B(n949), .Z(z3[13]) );
  NANDN U1418 ( .A(N518), .B(z2[13]), .Z(n949) );
  NANDN U1419 ( .A(n3), .B(N533), .Z(n948) );
  NAND U1420 ( .A(n950), .B(n951), .Z(z3[139]) );
  NANDN U1421 ( .A(N518), .B(z2[139]), .Z(n951) );
  NANDN U1422 ( .A(n3), .B(N659), .Z(n950) );
  NAND U1423 ( .A(n952), .B(n953), .Z(z3[138]) );
  NANDN U1424 ( .A(N518), .B(z2[138]), .Z(n953) );
  NANDN U1425 ( .A(n3), .B(N658), .Z(n952) );
  NAND U1426 ( .A(n954), .B(n955), .Z(z3[137]) );
  NANDN U1427 ( .A(N518), .B(z2[137]), .Z(n955) );
  NANDN U1428 ( .A(n3), .B(N657), .Z(n954) );
  NAND U1429 ( .A(n956), .B(n957), .Z(z3[136]) );
  NANDN U1430 ( .A(N518), .B(z2[136]), .Z(n957) );
  NANDN U1431 ( .A(n3), .B(N656), .Z(n956) );
  NAND U1432 ( .A(n958), .B(n959), .Z(z3[135]) );
  NANDN U1433 ( .A(N518), .B(z2[135]), .Z(n959) );
  NANDN U1434 ( .A(n3), .B(N655), .Z(n958) );
  NAND U1435 ( .A(n960), .B(n961), .Z(z3[134]) );
  NANDN U1436 ( .A(N518), .B(z2[134]), .Z(n961) );
  NANDN U1437 ( .A(n3), .B(N654), .Z(n960) );
  NAND U1438 ( .A(n962), .B(n963), .Z(z3[133]) );
  NANDN U1439 ( .A(N518), .B(z2[133]), .Z(n963) );
  NANDN U1440 ( .A(n3), .B(N653), .Z(n962) );
  NAND U1441 ( .A(n964), .B(n965), .Z(z3[132]) );
  NANDN U1442 ( .A(N518), .B(z2[132]), .Z(n965) );
  NANDN U1443 ( .A(n3), .B(N652), .Z(n964) );
  NAND U1444 ( .A(n966), .B(n967), .Z(z3[131]) );
  NANDN U1445 ( .A(N518), .B(z2[131]), .Z(n967) );
  NANDN U1446 ( .A(n3), .B(N651), .Z(n966) );
  NAND U1447 ( .A(n968), .B(n969), .Z(z3[130]) );
  NANDN U1448 ( .A(N518), .B(z2[130]), .Z(n969) );
  NANDN U1449 ( .A(n3), .B(N650), .Z(n968) );
  NAND U1450 ( .A(n970), .B(n971), .Z(z3[12]) );
  NANDN U1451 ( .A(N518), .B(z2[12]), .Z(n971) );
  NANDN U1452 ( .A(n3), .B(N532), .Z(n970) );
  NAND U1453 ( .A(n972), .B(n973), .Z(z3[129]) );
  NANDN U1454 ( .A(N518), .B(z2[129]), .Z(n973) );
  NANDN U1455 ( .A(n3), .B(N649), .Z(n972) );
  NAND U1456 ( .A(n974), .B(n975), .Z(z3[128]) );
  NANDN U1457 ( .A(N518), .B(z2[128]), .Z(n975) );
  NANDN U1458 ( .A(n3), .B(N648), .Z(n974) );
  NAND U1459 ( .A(n976), .B(n977), .Z(z3[127]) );
  NANDN U1460 ( .A(N518), .B(z2[127]), .Z(n977) );
  NANDN U1461 ( .A(n3), .B(N647), .Z(n976) );
  NAND U1462 ( .A(n978), .B(n979), .Z(z3[126]) );
  NANDN U1463 ( .A(N518), .B(z2[126]), .Z(n979) );
  NANDN U1464 ( .A(n3), .B(N646), .Z(n978) );
  NAND U1465 ( .A(n980), .B(n981), .Z(z3[125]) );
  NANDN U1466 ( .A(N518), .B(z2[125]), .Z(n981) );
  NANDN U1467 ( .A(n3), .B(N645), .Z(n980) );
  NAND U1468 ( .A(n982), .B(n983), .Z(z3[124]) );
  NANDN U1469 ( .A(N518), .B(z2[124]), .Z(n983) );
  NANDN U1470 ( .A(n3), .B(N644), .Z(n982) );
  NAND U1471 ( .A(n984), .B(n985), .Z(z3[123]) );
  NANDN U1472 ( .A(N518), .B(z2[123]), .Z(n985) );
  NANDN U1473 ( .A(n3), .B(N643), .Z(n984) );
  NAND U1474 ( .A(n986), .B(n987), .Z(z3[122]) );
  NANDN U1475 ( .A(N518), .B(z2[122]), .Z(n987) );
  NANDN U1476 ( .A(n3), .B(N642), .Z(n986) );
  NAND U1477 ( .A(n988), .B(n989), .Z(z3[121]) );
  NANDN U1478 ( .A(N518), .B(z2[121]), .Z(n989) );
  NANDN U1479 ( .A(n3), .B(N641), .Z(n988) );
  NAND U1480 ( .A(n990), .B(n991), .Z(z3[120]) );
  NANDN U1481 ( .A(N518), .B(z2[120]), .Z(n991) );
  NANDN U1482 ( .A(n3), .B(N640), .Z(n990) );
  NAND U1483 ( .A(n992), .B(n993), .Z(z3[11]) );
  NANDN U1484 ( .A(N518), .B(z2[11]), .Z(n993) );
  NANDN U1485 ( .A(n3), .B(N531), .Z(n992) );
  NAND U1486 ( .A(n994), .B(n995), .Z(z3[119]) );
  NANDN U1487 ( .A(N518), .B(z2[119]), .Z(n995) );
  NANDN U1488 ( .A(n3), .B(N639), .Z(n994) );
  NAND U1489 ( .A(n996), .B(n997), .Z(z3[118]) );
  NANDN U1490 ( .A(N518), .B(z2[118]), .Z(n997) );
  NANDN U1491 ( .A(n3), .B(N638), .Z(n996) );
  NAND U1492 ( .A(n998), .B(n999), .Z(z3[117]) );
  NANDN U1493 ( .A(N518), .B(z2[117]), .Z(n999) );
  NANDN U1494 ( .A(n3), .B(N637), .Z(n998) );
  NAND U1495 ( .A(n1000), .B(n1001), .Z(z3[116]) );
  NANDN U1496 ( .A(N518), .B(z2[116]), .Z(n1001) );
  NANDN U1497 ( .A(n3), .B(N636), .Z(n1000) );
  NAND U1498 ( .A(n1002), .B(n1003), .Z(z3[115]) );
  NANDN U1499 ( .A(N518), .B(z2[115]), .Z(n1003) );
  NANDN U1500 ( .A(n3), .B(N635), .Z(n1002) );
  NAND U1501 ( .A(n1004), .B(n1005), .Z(z3[114]) );
  NANDN U1502 ( .A(N518), .B(z2[114]), .Z(n1005) );
  NANDN U1503 ( .A(n3), .B(N634), .Z(n1004) );
  NAND U1504 ( .A(n1006), .B(n1007), .Z(z3[113]) );
  NANDN U1505 ( .A(N518), .B(z2[113]), .Z(n1007) );
  NANDN U1506 ( .A(n3), .B(N633), .Z(n1006) );
  NAND U1507 ( .A(n1008), .B(n1009), .Z(z3[112]) );
  NANDN U1508 ( .A(N518), .B(z2[112]), .Z(n1009) );
  NANDN U1509 ( .A(n3), .B(N632), .Z(n1008) );
  NAND U1510 ( .A(n1010), .B(n1011), .Z(z3[111]) );
  NANDN U1511 ( .A(N518), .B(z2[111]), .Z(n1011) );
  NANDN U1512 ( .A(n3), .B(N631), .Z(n1010) );
  NAND U1513 ( .A(n1012), .B(n1013), .Z(z3[110]) );
  NANDN U1514 ( .A(N518), .B(z2[110]), .Z(n1013) );
  NANDN U1515 ( .A(n3), .B(N630), .Z(n1012) );
  NAND U1516 ( .A(n1014), .B(n1015), .Z(z3[10]) );
  NANDN U1517 ( .A(N518), .B(z2[10]), .Z(n1015) );
  NANDN U1518 ( .A(n3), .B(N530), .Z(n1014) );
  NAND U1519 ( .A(n1016), .B(n1017), .Z(z3[109]) );
  NANDN U1520 ( .A(N518), .B(z2[109]), .Z(n1017) );
  NANDN U1521 ( .A(n3), .B(N629), .Z(n1016) );
  NAND U1522 ( .A(n1018), .B(n1019), .Z(z3[108]) );
  NANDN U1523 ( .A(N518), .B(z2[108]), .Z(n1019) );
  NANDN U1524 ( .A(n3), .B(N628), .Z(n1018) );
  NAND U1525 ( .A(n1020), .B(n1021), .Z(z3[107]) );
  NANDN U1526 ( .A(N518), .B(z2[107]), .Z(n1021) );
  NANDN U1527 ( .A(n3), .B(N627), .Z(n1020) );
  NAND U1528 ( .A(n1022), .B(n1023), .Z(z3[106]) );
  NANDN U1529 ( .A(N518), .B(z2[106]), .Z(n1023) );
  NANDN U1530 ( .A(n3), .B(N626), .Z(n1022) );
  NAND U1531 ( .A(n1024), .B(n1025), .Z(z3[105]) );
  NANDN U1532 ( .A(N518), .B(z2[105]), .Z(n1025) );
  NANDN U1533 ( .A(n3), .B(N625), .Z(n1024) );
  NAND U1534 ( .A(n1026), .B(n1027), .Z(z3[104]) );
  NANDN U1535 ( .A(N518), .B(z2[104]), .Z(n1027) );
  NANDN U1536 ( .A(n3), .B(N624), .Z(n1026) );
  NAND U1537 ( .A(n1028), .B(n1029), .Z(z3[103]) );
  NANDN U1538 ( .A(N518), .B(z2[103]), .Z(n1029) );
  NANDN U1539 ( .A(n3), .B(N623), .Z(n1028) );
  NAND U1540 ( .A(n1030), .B(n1031), .Z(z3[102]) );
  NANDN U1541 ( .A(N518), .B(z2[102]), .Z(n1031) );
  NANDN U1542 ( .A(n3), .B(N622), .Z(n1030) );
  NAND U1543 ( .A(n1032), .B(n1033), .Z(z3[101]) );
  NANDN U1544 ( .A(N518), .B(z2[101]), .Z(n1033) );
  NANDN U1545 ( .A(n3), .B(N621), .Z(n1032) );
  NAND U1546 ( .A(n1034), .B(n1035), .Z(z3[100]) );
  NANDN U1547 ( .A(N518), .B(z2[100]), .Z(n1035) );
  NANDN U1548 ( .A(n3), .B(N620), .Z(n1034) );
  NAND U1549 ( .A(n1036), .B(n1037), .Z(z3[0]) );
  NANDN U1550 ( .A(N518), .B(z2[0]), .Z(n1037) );
  NANDN U1551 ( .A(n3), .B(N520), .Z(n1036) );
  IV U1552 ( .A(N518), .Z(n3) );
  NAND U1553 ( .A(n1038), .B(n1039), .Z(z2[9]) );
  NANDN U1554 ( .A(xregN_1), .B(zin[8]), .Z(n1039) );
  NAND U1555 ( .A(N13), .B(xregN_1), .Z(n1038) );
  NAND U1556 ( .A(n1040), .B(n1041), .Z(z2[99]) );
  NANDN U1557 ( .A(xregN_1), .B(zin[98]), .Z(n1041) );
  NAND U1558 ( .A(N103), .B(xregN_1), .Z(n1040) );
  NAND U1559 ( .A(n1042), .B(n1043), .Z(z2[98]) );
  NANDN U1560 ( .A(xregN_1), .B(zin[97]), .Z(n1043) );
  NAND U1561 ( .A(N102), .B(xregN_1), .Z(n1042) );
  NAND U1562 ( .A(n1044), .B(n1045), .Z(z2[97]) );
  NANDN U1563 ( .A(xregN_1), .B(zin[96]), .Z(n1045) );
  NAND U1564 ( .A(N101), .B(xregN_1), .Z(n1044) );
  NAND U1565 ( .A(n1046), .B(n1047), .Z(z2[96]) );
  NANDN U1566 ( .A(xregN_1), .B(zin[95]), .Z(n1047) );
  NAND U1567 ( .A(N100), .B(xregN_1), .Z(n1046) );
  NAND U1568 ( .A(n1048), .B(n1049), .Z(z2[95]) );
  NANDN U1569 ( .A(xregN_1), .B(zin[94]), .Z(n1049) );
  NAND U1570 ( .A(N99), .B(xregN_1), .Z(n1048) );
  NAND U1571 ( .A(n1050), .B(n1051), .Z(z2[94]) );
  NANDN U1572 ( .A(xregN_1), .B(zin[93]), .Z(n1051) );
  NAND U1573 ( .A(N98), .B(xregN_1), .Z(n1050) );
  NAND U1574 ( .A(n1052), .B(n1053), .Z(z2[93]) );
  NANDN U1575 ( .A(xregN_1), .B(zin[92]), .Z(n1053) );
  NAND U1576 ( .A(N97), .B(xregN_1), .Z(n1052) );
  NAND U1577 ( .A(n1054), .B(n1055), .Z(z2[92]) );
  NANDN U1578 ( .A(xregN_1), .B(zin[91]), .Z(n1055) );
  NAND U1579 ( .A(N96), .B(xregN_1), .Z(n1054) );
  NAND U1580 ( .A(n1056), .B(n1057), .Z(z2[91]) );
  NANDN U1581 ( .A(xregN_1), .B(zin[90]), .Z(n1057) );
  NAND U1582 ( .A(N95), .B(xregN_1), .Z(n1056) );
  NAND U1583 ( .A(n1058), .B(n1059), .Z(z2[90]) );
  NANDN U1584 ( .A(xregN_1), .B(zin[89]), .Z(n1059) );
  NAND U1585 ( .A(N94), .B(xregN_1), .Z(n1058) );
  NAND U1586 ( .A(n1060), .B(n1061), .Z(z2[8]) );
  NANDN U1587 ( .A(xregN_1), .B(zin[7]), .Z(n1061) );
  NAND U1588 ( .A(N12), .B(xregN_1), .Z(n1060) );
  NAND U1589 ( .A(n1062), .B(n1063), .Z(z2[89]) );
  NANDN U1590 ( .A(xregN_1), .B(zin[88]), .Z(n1063) );
  NAND U1591 ( .A(N93), .B(xregN_1), .Z(n1062) );
  NAND U1592 ( .A(n1064), .B(n1065), .Z(z2[88]) );
  NANDN U1593 ( .A(xregN_1), .B(zin[87]), .Z(n1065) );
  NAND U1594 ( .A(N92), .B(xregN_1), .Z(n1064) );
  NAND U1595 ( .A(n1066), .B(n1067), .Z(z2[87]) );
  NANDN U1596 ( .A(xregN_1), .B(zin[86]), .Z(n1067) );
  NAND U1597 ( .A(N91), .B(xregN_1), .Z(n1066) );
  NAND U1598 ( .A(n1068), .B(n1069), .Z(z2[86]) );
  NANDN U1599 ( .A(xregN_1), .B(zin[85]), .Z(n1069) );
  NAND U1600 ( .A(N90), .B(xregN_1), .Z(n1068) );
  NAND U1601 ( .A(n1070), .B(n1071), .Z(z2[85]) );
  NANDN U1602 ( .A(xregN_1), .B(zin[84]), .Z(n1071) );
  NAND U1603 ( .A(N89), .B(xregN_1), .Z(n1070) );
  NAND U1604 ( .A(n1072), .B(n1073), .Z(z2[84]) );
  NANDN U1605 ( .A(xregN_1), .B(zin[83]), .Z(n1073) );
  NAND U1606 ( .A(N88), .B(xregN_1), .Z(n1072) );
  NAND U1607 ( .A(n1074), .B(n1075), .Z(z2[83]) );
  NANDN U1608 ( .A(xregN_1), .B(zin[82]), .Z(n1075) );
  NAND U1609 ( .A(N87), .B(xregN_1), .Z(n1074) );
  NAND U1610 ( .A(n1076), .B(n1077), .Z(z2[82]) );
  NANDN U1611 ( .A(xregN_1), .B(zin[81]), .Z(n1077) );
  NAND U1612 ( .A(N86), .B(xregN_1), .Z(n1076) );
  NAND U1613 ( .A(n1078), .B(n1079), .Z(z2[81]) );
  NANDN U1614 ( .A(xregN_1), .B(zin[80]), .Z(n1079) );
  NAND U1615 ( .A(N85), .B(xregN_1), .Z(n1078) );
  NAND U1616 ( .A(n1080), .B(n1081), .Z(z2[80]) );
  NANDN U1617 ( .A(xregN_1), .B(zin[79]), .Z(n1081) );
  NAND U1618 ( .A(N84), .B(xregN_1), .Z(n1080) );
  NAND U1619 ( .A(n1082), .B(n1083), .Z(z2[7]) );
  NANDN U1620 ( .A(xregN_1), .B(zin[6]), .Z(n1083) );
  NAND U1621 ( .A(N11), .B(xregN_1), .Z(n1082) );
  NAND U1622 ( .A(n1084), .B(n1085), .Z(z2[79]) );
  NANDN U1623 ( .A(xregN_1), .B(zin[78]), .Z(n1085) );
  NAND U1624 ( .A(N83), .B(xregN_1), .Z(n1084) );
  NAND U1625 ( .A(n1086), .B(n1087), .Z(z2[78]) );
  NANDN U1626 ( .A(xregN_1), .B(zin[77]), .Z(n1087) );
  NAND U1627 ( .A(N82), .B(xregN_1), .Z(n1086) );
  NAND U1628 ( .A(n1088), .B(n1089), .Z(z2[77]) );
  NANDN U1629 ( .A(xregN_1), .B(zin[76]), .Z(n1089) );
  NAND U1630 ( .A(N81), .B(xregN_1), .Z(n1088) );
  NAND U1631 ( .A(n1090), .B(n1091), .Z(z2[76]) );
  NANDN U1632 ( .A(xregN_1), .B(zin[75]), .Z(n1091) );
  NAND U1633 ( .A(N80), .B(xregN_1), .Z(n1090) );
  NAND U1634 ( .A(n1092), .B(n1093), .Z(z2[75]) );
  NANDN U1635 ( .A(xregN_1), .B(zin[74]), .Z(n1093) );
  NAND U1636 ( .A(N79), .B(xregN_1), .Z(n1092) );
  NAND U1637 ( .A(n1094), .B(n1095), .Z(z2[74]) );
  NANDN U1638 ( .A(xregN_1), .B(zin[73]), .Z(n1095) );
  NAND U1639 ( .A(N78), .B(xregN_1), .Z(n1094) );
  NAND U1640 ( .A(n1096), .B(n1097), .Z(z2[73]) );
  NANDN U1641 ( .A(xregN_1), .B(zin[72]), .Z(n1097) );
  NAND U1642 ( .A(N77), .B(xregN_1), .Z(n1096) );
  NAND U1643 ( .A(n1098), .B(n1099), .Z(z2[72]) );
  NANDN U1644 ( .A(xregN_1), .B(zin[71]), .Z(n1099) );
  NAND U1645 ( .A(N76), .B(xregN_1), .Z(n1098) );
  NAND U1646 ( .A(n1100), .B(n1101), .Z(z2[71]) );
  NANDN U1647 ( .A(xregN_1), .B(zin[70]), .Z(n1101) );
  NAND U1648 ( .A(N75), .B(xregN_1), .Z(n1100) );
  NAND U1649 ( .A(n1102), .B(n1103), .Z(z2[70]) );
  NANDN U1650 ( .A(xregN_1), .B(zin[69]), .Z(n1103) );
  NAND U1651 ( .A(N74), .B(xregN_1), .Z(n1102) );
  NAND U1652 ( .A(n1104), .B(n1105), .Z(z2[6]) );
  NANDN U1653 ( .A(xregN_1), .B(zin[5]), .Z(n1105) );
  NAND U1654 ( .A(N10), .B(xregN_1), .Z(n1104) );
  NAND U1655 ( .A(n1106), .B(n1107), .Z(z2[69]) );
  NANDN U1656 ( .A(xregN_1), .B(zin[68]), .Z(n1107) );
  NAND U1657 ( .A(N73), .B(xregN_1), .Z(n1106) );
  NAND U1658 ( .A(n1108), .B(n1109), .Z(z2[68]) );
  NANDN U1659 ( .A(xregN_1), .B(zin[67]), .Z(n1109) );
  NAND U1660 ( .A(N72), .B(xregN_1), .Z(n1108) );
  NAND U1661 ( .A(n1110), .B(n1111), .Z(z2[67]) );
  NANDN U1662 ( .A(xregN_1), .B(zin[66]), .Z(n1111) );
  NAND U1663 ( .A(N71), .B(xregN_1), .Z(n1110) );
  NAND U1664 ( .A(n1112), .B(n1113), .Z(z2[66]) );
  NANDN U1665 ( .A(xregN_1), .B(zin[65]), .Z(n1113) );
  NAND U1666 ( .A(N70), .B(xregN_1), .Z(n1112) );
  NAND U1667 ( .A(n1114), .B(n1115), .Z(z2[65]) );
  NANDN U1668 ( .A(xregN_1), .B(zin[64]), .Z(n1115) );
  NAND U1669 ( .A(N69), .B(xregN_1), .Z(n1114) );
  NAND U1670 ( .A(n1116), .B(n1117), .Z(z2[64]) );
  NANDN U1671 ( .A(xregN_1), .B(zin[63]), .Z(n1117) );
  NAND U1672 ( .A(N68), .B(xregN_1), .Z(n1116) );
  NAND U1673 ( .A(n1118), .B(n1119), .Z(z2[63]) );
  NANDN U1674 ( .A(xregN_1), .B(zin[62]), .Z(n1119) );
  NAND U1675 ( .A(N67), .B(xregN_1), .Z(n1118) );
  NAND U1676 ( .A(n1120), .B(n1121), .Z(z2[62]) );
  NANDN U1677 ( .A(xregN_1), .B(zin[61]), .Z(n1121) );
  NAND U1678 ( .A(N66), .B(xregN_1), .Z(n1120) );
  NAND U1679 ( .A(n1122), .B(n1123), .Z(z2[61]) );
  NANDN U1680 ( .A(xregN_1), .B(zin[60]), .Z(n1123) );
  NAND U1681 ( .A(N65), .B(xregN_1), .Z(n1122) );
  NAND U1682 ( .A(n1124), .B(n1125), .Z(z2[60]) );
  NANDN U1683 ( .A(xregN_1), .B(zin[59]), .Z(n1125) );
  NAND U1684 ( .A(N64), .B(xregN_1), .Z(n1124) );
  NAND U1685 ( .A(n1126), .B(n1127), .Z(z2[5]) );
  NANDN U1686 ( .A(xregN_1), .B(zin[4]), .Z(n1127) );
  NAND U1687 ( .A(N9), .B(xregN_1), .Z(n1126) );
  NAND U1688 ( .A(n1128), .B(n1129), .Z(z2[59]) );
  NANDN U1689 ( .A(xregN_1), .B(zin[58]), .Z(n1129) );
  NAND U1690 ( .A(N63), .B(xregN_1), .Z(n1128) );
  NAND U1691 ( .A(n1130), .B(n1131), .Z(z2[58]) );
  NANDN U1692 ( .A(xregN_1), .B(zin[57]), .Z(n1131) );
  NAND U1693 ( .A(N62), .B(xregN_1), .Z(n1130) );
  NAND U1694 ( .A(n1132), .B(n1133), .Z(z2[57]) );
  NANDN U1695 ( .A(xregN_1), .B(zin[56]), .Z(n1133) );
  NAND U1696 ( .A(N61), .B(xregN_1), .Z(n1132) );
  NAND U1697 ( .A(n1134), .B(n1135), .Z(z2[56]) );
  NANDN U1698 ( .A(xregN_1), .B(zin[55]), .Z(n1135) );
  NAND U1699 ( .A(N60), .B(xregN_1), .Z(n1134) );
  NAND U1700 ( .A(n1136), .B(n1137), .Z(z2[55]) );
  NANDN U1701 ( .A(xregN_1), .B(zin[54]), .Z(n1137) );
  NAND U1702 ( .A(N59), .B(xregN_1), .Z(n1136) );
  NAND U1703 ( .A(n1138), .B(n1139), .Z(z2[54]) );
  NANDN U1704 ( .A(xregN_1), .B(zin[53]), .Z(n1139) );
  NAND U1705 ( .A(N58), .B(xregN_1), .Z(n1138) );
  NAND U1706 ( .A(n1140), .B(n1141), .Z(z2[53]) );
  NANDN U1707 ( .A(xregN_1), .B(zin[52]), .Z(n1141) );
  NAND U1708 ( .A(N57), .B(xregN_1), .Z(n1140) );
  NAND U1709 ( .A(n1142), .B(n1143), .Z(z2[52]) );
  NANDN U1710 ( .A(xregN_1), .B(zin[51]), .Z(n1143) );
  NAND U1711 ( .A(N56), .B(xregN_1), .Z(n1142) );
  NAND U1712 ( .A(n1144), .B(n1145), .Z(z2[51]) );
  NANDN U1713 ( .A(xregN_1), .B(zin[50]), .Z(n1145) );
  NAND U1714 ( .A(N55), .B(xregN_1), .Z(n1144) );
  NAND U1715 ( .A(n1146), .B(n1147), .Z(z2[513]) );
  NANDN U1716 ( .A(xregN_1), .B(zin[512]), .Z(n1147) );
  NAND U1717 ( .A(N517), .B(xregN_1), .Z(n1146) );
  NAND U1718 ( .A(n1148), .B(n1149), .Z(z2[512]) );
  NANDN U1719 ( .A(xregN_1), .B(zin[511]), .Z(n1149) );
  NAND U1720 ( .A(N516), .B(xregN_1), .Z(n1148) );
  NAND U1721 ( .A(n1150), .B(n1151), .Z(z2[511]) );
  NANDN U1722 ( .A(xregN_1), .B(zin[510]), .Z(n1151) );
  NAND U1723 ( .A(N515), .B(xregN_1), .Z(n1150) );
  NAND U1724 ( .A(n1152), .B(n1153), .Z(z2[510]) );
  NANDN U1725 ( .A(xregN_1), .B(zin[509]), .Z(n1153) );
  NAND U1726 ( .A(N514), .B(xregN_1), .Z(n1152) );
  NAND U1727 ( .A(n1154), .B(n1155), .Z(z2[50]) );
  NANDN U1728 ( .A(xregN_1), .B(zin[49]), .Z(n1155) );
  NAND U1729 ( .A(N54), .B(xregN_1), .Z(n1154) );
  NAND U1730 ( .A(n1156), .B(n1157), .Z(z2[509]) );
  NANDN U1731 ( .A(xregN_1), .B(zin[508]), .Z(n1157) );
  NAND U1732 ( .A(N513), .B(xregN_1), .Z(n1156) );
  NAND U1733 ( .A(n1158), .B(n1159), .Z(z2[508]) );
  NANDN U1734 ( .A(xregN_1), .B(zin[507]), .Z(n1159) );
  NAND U1735 ( .A(N512), .B(xregN_1), .Z(n1158) );
  NAND U1736 ( .A(n1160), .B(n1161), .Z(z2[507]) );
  NANDN U1737 ( .A(xregN_1), .B(zin[506]), .Z(n1161) );
  NAND U1738 ( .A(N511), .B(xregN_1), .Z(n1160) );
  NAND U1739 ( .A(n1162), .B(n1163), .Z(z2[506]) );
  NANDN U1740 ( .A(xregN_1), .B(zin[505]), .Z(n1163) );
  NAND U1741 ( .A(N510), .B(xregN_1), .Z(n1162) );
  NAND U1742 ( .A(n1164), .B(n1165), .Z(z2[505]) );
  NANDN U1743 ( .A(xregN_1), .B(zin[504]), .Z(n1165) );
  NAND U1744 ( .A(N509), .B(xregN_1), .Z(n1164) );
  NAND U1745 ( .A(n1166), .B(n1167), .Z(z2[504]) );
  NANDN U1746 ( .A(xregN_1), .B(zin[503]), .Z(n1167) );
  NAND U1747 ( .A(N508), .B(xregN_1), .Z(n1166) );
  NAND U1748 ( .A(n1168), .B(n1169), .Z(z2[503]) );
  NANDN U1749 ( .A(xregN_1), .B(zin[502]), .Z(n1169) );
  NAND U1750 ( .A(N507), .B(xregN_1), .Z(n1168) );
  NAND U1751 ( .A(n1170), .B(n1171), .Z(z2[502]) );
  NANDN U1752 ( .A(xregN_1), .B(zin[501]), .Z(n1171) );
  NAND U1753 ( .A(N506), .B(xregN_1), .Z(n1170) );
  NAND U1754 ( .A(n1172), .B(n1173), .Z(z2[501]) );
  NANDN U1755 ( .A(xregN_1), .B(zin[500]), .Z(n1173) );
  NAND U1756 ( .A(N505), .B(xregN_1), .Z(n1172) );
  NAND U1757 ( .A(n1174), .B(n1175), .Z(z2[500]) );
  NANDN U1758 ( .A(xregN_1), .B(zin[499]), .Z(n1175) );
  NAND U1759 ( .A(N504), .B(xregN_1), .Z(n1174) );
  NAND U1760 ( .A(n1176), .B(n1177), .Z(z2[4]) );
  NANDN U1761 ( .A(xregN_1), .B(zin[3]), .Z(n1177) );
  NAND U1762 ( .A(N8), .B(xregN_1), .Z(n1176) );
  NAND U1763 ( .A(n1178), .B(n1179), .Z(z2[49]) );
  NANDN U1764 ( .A(xregN_1), .B(zin[48]), .Z(n1179) );
  NAND U1765 ( .A(N53), .B(xregN_1), .Z(n1178) );
  NAND U1766 ( .A(n1180), .B(n1181), .Z(z2[499]) );
  NANDN U1767 ( .A(xregN_1), .B(zin[498]), .Z(n1181) );
  NAND U1768 ( .A(N503), .B(xregN_1), .Z(n1180) );
  NAND U1769 ( .A(n1182), .B(n1183), .Z(z2[498]) );
  NANDN U1770 ( .A(xregN_1), .B(zin[497]), .Z(n1183) );
  NAND U1771 ( .A(N502), .B(xregN_1), .Z(n1182) );
  NAND U1772 ( .A(n1184), .B(n1185), .Z(z2[497]) );
  NANDN U1773 ( .A(xregN_1), .B(zin[496]), .Z(n1185) );
  NAND U1774 ( .A(N501), .B(xregN_1), .Z(n1184) );
  NAND U1775 ( .A(n1186), .B(n1187), .Z(z2[496]) );
  NANDN U1776 ( .A(xregN_1), .B(zin[495]), .Z(n1187) );
  NAND U1777 ( .A(N500), .B(xregN_1), .Z(n1186) );
  NAND U1778 ( .A(n1188), .B(n1189), .Z(z2[495]) );
  NANDN U1779 ( .A(xregN_1), .B(zin[494]), .Z(n1189) );
  NAND U1780 ( .A(N499), .B(xregN_1), .Z(n1188) );
  NAND U1781 ( .A(n1190), .B(n1191), .Z(z2[494]) );
  NANDN U1782 ( .A(xregN_1), .B(zin[493]), .Z(n1191) );
  NAND U1783 ( .A(N498), .B(xregN_1), .Z(n1190) );
  NAND U1784 ( .A(n1192), .B(n1193), .Z(z2[493]) );
  NANDN U1785 ( .A(xregN_1), .B(zin[492]), .Z(n1193) );
  NAND U1786 ( .A(N497), .B(xregN_1), .Z(n1192) );
  NAND U1787 ( .A(n1194), .B(n1195), .Z(z2[492]) );
  NANDN U1788 ( .A(xregN_1), .B(zin[491]), .Z(n1195) );
  NAND U1789 ( .A(N496), .B(xregN_1), .Z(n1194) );
  NAND U1790 ( .A(n1196), .B(n1197), .Z(z2[491]) );
  NANDN U1791 ( .A(xregN_1), .B(zin[490]), .Z(n1197) );
  NAND U1792 ( .A(N495), .B(xregN_1), .Z(n1196) );
  NAND U1793 ( .A(n1198), .B(n1199), .Z(z2[490]) );
  NANDN U1794 ( .A(xregN_1), .B(zin[489]), .Z(n1199) );
  NAND U1795 ( .A(N494), .B(xregN_1), .Z(n1198) );
  NAND U1796 ( .A(n1200), .B(n1201), .Z(z2[48]) );
  NANDN U1797 ( .A(xregN_1), .B(zin[47]), .Z(n1201) );
  NAND U1798 ( .A(N52), .B(xregN_1), .Z(n1200) );
  NAND U1799 ( .A(n1202), .B(n1203), .Z(z2[489]) );
  NANDN U1800 ( .A(xregN_1), .B(zin[488]), .Z(n1203) );
  NAND U1801 ( .A(N493), .B(xregN_1), .Z(n1202) );
  NAND U1802 ( .A(n1204), .B(n1205), .Z(z2[488]) );
  NANDN U1803 ( .A(xregN_1), .B(zin[487]), .Z(n1205) );
  NAND U1804 ( .A(N492), .B(xregN_1), .Z(n1204) );
  NAND U1805 ( .A(n1206), .B(n1207), .Z(z2[487]) );
  NANDN U1806 ( .A(xregN_1), .B(zin[486]), .Z(n1207) );
  NAND U1807 ( .A(N491), .B(xregN_1), .Z(n1206) );
  NAND U1808 ( .A(n1208), .B(n1209), .Z(z2[486]) );
  NANDN U1809 ( .A(xregN_1), .B(zin[485]), .Z(n1209) );
  NAND U1810 ( .A(N490), .B(xregN_1), .Z(n1208) );
  NAND U1811 ( .A(n1210), .B(n1211), .Z(z2[485]) );
  NANDN U1812 ( .A(xregN_1), .B(zin[484]), .Z(n1211) );
  NAND U1813 ( .A(N489), .B(xregN_1), .Z(n1210) );
  NAND U1814 ( .A(n1212), .B(n1213), .Z(z2[484]) );
  NANDN U1815 ( .A(xregN_1), .B(zin[483]), .Z(n1213) );
  NAND U1816 ( .A(N488), .B(xregN_1), .Z(n1212) );
  NAND U1817 ( .A(n1214), .B(n1215), .Z(z2[483]) );
  NANDN U1818 ( .A(xregN_1), .B(zin[482]), .Z(n1215) );
  NAND U1819 ( .A(N487), .B(xregN_1), .Z(n1214) );
  NAND U1820 ( .A(n1216), .B(n1217), .Z(z2[482]) );
  NANDN U1821 ( .A(xregN_1), .B(zin[481]), .Z(n1217) );
  NAND U1822 ( .A(N486), .B(xregN_1), .Z(n1216) );
  NAND U1823 ( .A(n1218), .B(n1219), .Z(z2[481]) );
  NANDN U1824 ( .A(xregN_1), .B(zin[480]), .Z(n1219) );
  NAND U1825 ( .A(N485), .B(xregN_1), .Z(n1218) );
  NAND U1826 ( .A(n1220), .B(n1221), .Z(z2[480]) );
  NANDN U1827 ( .A(xregN_1), .B(zin[479]), .Z(n1221) );
  NAND U1828 ( .A(N484), .B(xregN_1), .Z(n1220) );
  NAND U1829 ( .A(n1222), .B(n1223), .Z(z2[47]) );
  NANDN U1830 ( .A(xregN_1), .B(zin[46]), .Z(n1223) );
  NAND U1831 ( .A(N51), .B(xregN_1), .Z(n1222) );
  NAND U1832 ( .A(n1224), .B(n1225), .Z(z2[479]) );
  NANDN U1833 ( .A(xregN_1), .B(zin[478]), .Z(n1225) );
  NAND U1834 ( .A(N483), .B(xregN_1), .Z(n1224) );
  NAND U1835 ( .A(n1226), .B(n1227), .Z(z2[478]) );
  NANDN U1836 ( .A(xregN_1), .B(zin[477]), .Z(n1227) );
  NAND U1837 ( .A(N482), .B(xregN_1), .Z(n1226) );
  NAND U1838 ( .A(n1228), .B(n1229), .Z(z2[477]) );
  NANDN U1839 ( .A(xregN_1), .B(zin[476]), .Z(n1229) );
  NAND U1840 ( .A(N481), .B(xregN_1), .Z(n1228) );
  NAND U1841 ( .A(n1230), .B(n1231), .Z(z2[476]) );
  NANDN U1842 ( .A(xregN_1), .B(zin[475]), .Z(n1231) );
  NAND U1843 ( .A(N480), .B(xregN_1), .Z(n1230) );
  NAND U1844 ( .A(n1232), .B(n1233), .Z(z2[475]) );
  NANDN U1845 ( .A(xregN_1), .B(zin[474]), .Z(n1233) );
  NAND U1846 ( .A(N479), .B(xregN_1), .Z(n1232) );
  NAND U1847 ( .A(n1234), .B(n1235), .Z(z2[474]) );
  NANDN U1848 ( .A(xregN_1), .B(zin[473]), .Z(n1235) );
  NAND U1849 ( .A(N478), .B(xregN_1), .Z(n1234) );
  NAND U1850 ( .A(n1236), .B(n1237), .Z(z2[473]) );
  NANDN U1851 ( .A(xregN_1), .B(zin[472]), .Z(n1237) );
  NAND U1852 ( .A(N477), .B(xregN_1), .Z(n1236) );
  NAND U1853 ( .A(n1238), .B(n1239), .Z(z2[472]) );
  NANDN U1854 ( .A(xregN_1), .B(zin[471]), .Z(n1239) );
  NAND U1855 ( .A(N476), .B(xregN_1), .Z(n1238) );
  NAND U1856 ( .A(n1240), .B(n1241), .Z(z2[471]) );
  NANDN U1857 ( .A(xregN_1), .B(zin[470]), .Z(n1241) );
  NAND U1858 ( .A(N475), .B(xregN_1), .Z(n1240) );
  NAND U1859 ( .A(n1242), .B(n1243), .Z(z2[470]) );
  NANDN U1860 ( .A(xregN_1), .B(zin[469]), .Z(n1243) );
  NAND U1861 ( .A(N474), .B(xregN_1), .Z(n1242) );
  NAND U1862 ( .A(n1244), .B(n1245), .Z(z2[46]) );
  NANDN U1863 ( .A(xregN_1), .B(zin[45]), .Z(n1245) );
  NAND U1864 ( .A(N50), .B(xregN_1), .Z(n1244) );
  NAND U1865 ( .A(n1246), .B(n1247), .Z(z2[469]) );
  NANDN U1866 ( .A(xregN_1), .B(zin[468]), .Z(n1247) );
  NAND U1867 ( .A(N473), .B(xregN_1), .Z(n1246) );
  NAND U1868 ( .A(n1248), .B(n1249), .Z(z2[468]) );
  NANDN U1869 ( .A(xregN_1), .B(zin[467]), .Z(n1249) );
  NAND U1870 ( .A(N472), .B(xregN_1), .Z(n1248) );
  NAND U1871 ( .A(n1250), .B(n1251), .Z(z2[467]) );
  NANDN U1872 ( .A(xregN_1), .B(zin[466]), .Z(n1251) );
  NAND U1873 ( .A(N471), .B(xregN_1), .Z(n1250) );
  NAND U1874 ( .A(n1252), .B(n1253), .Z(z2[466]) );
  NANDN U1875 ( .A(xregN_1), .B(zin[465]), .Z(n1253) );
  NAND U1876 ( .A(N470), .B(xregN_1), .Z(n1252) );
  NAND U1877 ( .A(n1254), .B(n1255), .Z(z2[465]) );
  NANDN U1878 ( .A(xregN_1), .B(zin[464]), .Z(n1255) );
  NAND U1879 ( .A(N469), .B(xregN_1), .Z(n1254) );
  NAND U1880 ( .A(n1256), .B(n1257), .Z(z2[464]) );
  NANDN U1881 ( .A(xregN_1), .B(zin[463]), .Z(n1257) );
  NAND U1882 ( .A(N468), .B(xregN_1), .Z(n1256) );
  NAND U1883 ( .A(n1258), .B(n1259), .Z(z2[463]) );
  NANDN U1884 ( .A(xregN_1), .B(zin[462]), .Z(n1259) );
  NAND U1885 ( .A(N467), .B(xregN_1), .Z(n1258) );
  NAND U1886 ( .A(n1260), .B(n1261), .Z(z2[462]) );
  NANDN U1887 ( .A(xregN_1), .B(zin[461]), .Z(n1261) );
  NAND U1888 ( .A(N466), .B(xregN_1), .Z(n1260) );
  NAND U1889 ( .A(n1262), .B(n1263), .Z(z2[461]) );
  NANDN U1890 ( .A(xregN_1), .B(zin[460]), .Z(n1263) );
  NAND U1891 ( .A(N465), .B(xregN_1), .Z(n1262) );
  NAND U1892 ( .A(n1264), .B(n1265), .Z(z2[460]) );
  NANDN U1893 ( .A(xregN_1), .B(zin[459]), .Z(n1265) );
  NAND U1894 ( .A(N464), .B(xregN_1), .Z(n1264) );
  NAND U1895 ( .A(n1266), .B(n1267), .Z(z2[45]) );
  NANDN U1896 ( .A(xregN_1), .B(zin[44]), .Z(n1267) );
  NAND U1897 ( .A(N49), .B(xregN_1), .Z(n1266) );
  NAND U1898 ( .A(n1268), .B(n1269), .Z(z2[459]) );
  NANDN U1899 ( .A(xregN_1), .B(zin[458]), .Z(n1269) );
  NAND U1900 ( .A(N463), .B(xregN_1), .Z(n1268) );
  NAND U1901 ( .A(n1270), .B(n1271), .Z(z2[458]) );
  NANDN U1902 ( .A(xregN_1), .B(zin[457]), .Z(n1271) );
  NAND U1903 ( .A(N462), .B(xregN_1), .Z(n1270) );
  NAND U1904 ( .A(n1272), .B(n1273), .Z(z2[457]) );
  NANDN U1905 ( .A(xregN_1), .B(zin[456]), .Z(n1273) );
  NAND U1906 ( .A(N461), .B(xregN_1), .Z(n1272) );
  NAND U1907 ( .A(n1274), .B(n1275), .Z(z2[456]) );
  NANDN U1908 ( .A(xregN_1), .B(zin[455]), .Z(n1275) );
  NAND U1909 ( .A(N460), .B(xregN_1), .Z(n1274) );
  NAND U1910 ( .A(n1276), .B(n1277), .Z(z2[455]) );
  NANDN U1911 ( .A(xregN_1), .B(zin[454]), .Z(n1277) );
  NAND U1912 ( .A(N459), .B(xregN_1), .Z(n1276) );
  NAND U1913 ( .A(n1278), .B(n1279), .Z(z2[454]) );
  NANDN U1914 ( .A(xregN_1), .B(zin[453]), .Z(n1279) );
  NAND U1915 ( .A(N458), .B(xregN_1), .Z(n1278) );
  NAND U1916 ( .A(n1280), .B(n1281), .Z(z2[453]) );
  NANDN U1917 ( .A(xregN_1), .B(zin[452]), .Z(n1281) );
  NAND U1918 ( .A(N457), .B(xregN_1), .Z(n1280) );
  NAND U1919 ( .A(n1282), .B(n1283), .Z(z2[452]) );
  NANDN U1920 ( .A(xregN_1), .B(zin[451]), .Z(n1283) );
  NAND U1921 ( .A(N456), .B(xregN_1), .Z(n1282) );
  NAND U1922 ( .A(n1284), .B(n1285), .Z(z2[451]) );
  NANDN U1923 ( .A(xregN_1), .B(zin[450]), .Z(n1285) );
  NAND U1924 ( .A(N455), .B(xregN_1), .Z(n1284) );
  NAND U1925 ( .A(n1286), .B(n1287), .Z(z2[450]) );
  NANDN U1926 ( .A(xregN_1), .B(zin[449]), .Z(n1287) );
  NAND U1927 ( .A(N454), .B(xregN_1), .Z(n1286) );
  NAND U1928 ( .A(n1288), .B(n1289), .Z(z2[44]) );
  NANDN U1929 ( .A(xregN_1), .B(zin[43]), .Z(n1289) );
  NAND U1930 ( .A(N48), .B(xregN_1), .Z(n1288) );
  NAND U1931 ( .A(n1290), .B(n1291), .Z(z2[449]) );
  NANDN U1932 ( .A(xregN_1), .B(zin[448]), .Z(n1291) );
  NAND U1933 ( .A(N453), .B(xregN_1), .Z(n1290) );
  NAND U1934 ( .A(n1292), .B(n1293), .Z(z2[448]) );
  NANDN U1935 ( .A(xregN_1), .B(zin[447]), .Z(n1293) );
  NAND U1936 ( .A(N452), .B(xregN_1), .Z(n1292) );
  NAND U1937 ( .A(n1294), .B(n1295), .Z(z2[447]) );
  NANDN U1938 ( .A(xregN_1), .B(zin[446]), .Z(n1295) );
  NAND U1939 ( .A(N451), .B(xregN_1), .Z(n1294) );
  NAND U1940 ( .A(n1296), .B(n1297), .Z(z2[446]) );
  NANDN U1941 ( .A(xregN_1), .B(zin[445]), .Z(n1297) );
  NAND U1942 ( .A(N450), .B(xregN_1), .Z(n1296) );
  NAND U1943 ( .A(n1298), .B(n1299), .Z(z2[445]) );
  NANDN U1944 ( .A(xregN_1), .B(zin[444]), .Z(n1299) );
  NAND U1945 ( .A(N449), .B(xregN_1), .Z(n1298) );
  NAND U1946 ( .A(n1300), .B(n1301), .Z(z2[444]) );
  NANDN U1947 ( .A(xregN_1), .B(zin[443]), .Z(n1301) );
  NAND U1948 ( .A(N448), .B(xregN_1), .Z(n1300) );
  NAND U1949 ( .A(n1302), .B(n1303), .Z(z2[443]) );
  NANDN U1950 ( .A(xregN_1), .B(zin[442]), .Z(n1303) );
  NAND U1951 ( .A(N447), .B(xregN_1), .Z(n1302) );
  NAND U1952 ( .A(n1304), .B(n1305), .Z(z2[442]) );
  NANDN U1953 ( .A(xregN_1), .B(zin[441]), .Z(n1305) );
  NAND U1954 ( .A(N446), .B(xregN_1), .Z(n1304) );
  NAND U1955 ( .A(n1306), .B(n1307), .Z(z2[441]) );
  NANDN U1956 ( .A(xregN_1), .B(zin[440]), .Z(n1307) );
  NAND U1957 ( .A(N445), .B(xregN_1), .Z(n1306) );
  NAND U1958 ( .A(n1308), .B(n1309), .Z(z2[440]) );
  NANDN U1959 ( .A(xregN_1), .B(zin[439]), .Z(n1309) );
  NAND U1960 ( .A(N444), .B(xregN_1), .Z(n1308) );
  NAND U1961 ( .A(n1310), .B(n1311), .Z(z2[43]) );
  NANDN U1962 ( .A(xregN_1), .B(zin[42]), .Z(n1311) );
  NAND U1963 ( .A(N47), .B(xregN_1), .Z(n1310) );
  NAND U1964 ( .A(n1312), .B(n1313), .Z(z2[439]) );
  NANDN U1965 ( .A(xregN_1), .B(zin[438]), .Z(n1313) );
  NAND U1966 ( .A(N443), .B(xregN_1), .Z(n1312) );
  NAND U1967 ( .A(n1314), .B(n1315), .Z(z2[438]) );
  NANDN U1968 ( .A(xregN_1), .B(zin[437]), .Z(n1315) );
  NAND U1969 ( .A(N442), .B(xregN_1), .Z(n1314) );
  NAND U1970 ( .A(n1316), .B(n1317), .Z(z2[437]) );
  NANDN U1971 ( .A(xregN_1), .B(zin[436]), .Z(n1317) );
  NAND U1972 ( .A(N441), .B(xregN_1), .Z(n1316) );
  NAND U1973 ( .A(n1318), .B(n1319), .Z(z2[436]) );
  NANDN U1974 ( .A(xregN_1), .B(zin[435]), .Z(n1319) );
  NAND U1975 ( .A(N440), .B(xregN_1), .Z(n1318) );
  NAND U1976 ( .A(n1320), .B(n1321), .Z(z2[435]) );
  NANDN U1977 ( .A(xregN_1), .B(zin[434]), .Z(n1321) );
  NAND U1978 ( .A(N439), .B(xregN_1), .Z(n1320) );
  NAND U1979 ( .A(n1322), .B(n1323), .Z(z2[434]) );
  NANDN U1980 ( .A(xregN_1), .B(zin[433]), .Z(n1323) );
  NAND U1981 ( .A(N438), .B(xregN_1), .Z(n1322) );
  NAND U1982 ( .A(n1324), .B(n1325), .Z(z2[433]) );
  NANDN U1983 ( .A(xregN_1), .B(zin[432]), .Z(n1325) );
  NAND U1984 ( .A(N437), .B(xregN_1), .Z(n1324) );
  NAND U1985 ( .A(n1326), .B(n1327), .Z(z2[432]) );
  NANDN U1986 ( .A(xregN_1), .B(zin[431]), .Z(n1327) );
  NAND U1987 ( .A(N436), .B(xregN_1), .Z(n1326) );
  NAND U1988 ( .A(n1328), .B(n1329), .Z(z2[431]) );
  NANDN U1989 ( .A(xregN_1), .B(zin[430]), .Z(n1329) );
  NAND U1990 ( .A(N435), .B(xregN_1), .Z(n1328) );
  NAND U1991 ( .A(n1330), .B(n1331), .Z(z2[430]) );
  NANDN U1992 ( .A(xregN_1), .B(zin[429]), .Z(n1331) );
  NAND U1993 ( .A(N434), .B(xregN_1), .Z(n1330) );
  NAND U1994 ( .A(n1332), .B(n1333), .Z(z2[42]) );
  NANDN U1995 ( .A(xregN_1), .B(zin[41]), .Z(n1333) );
  NAND U1996 ( .A(N46), .B(xregN_1), .Z(n1332) );
  NAND U1997 ( .A(n1334), .B(n1335), .Z(z2[429]) );
  NANDN U1998 ( .A(xregN_1), .B(zin[428]), .Z(n1335) );
  NAND U1999 ( .A(N433), .B(xregN_1), .Z(n1334) );
  NAND U2000 ( .A(n1336), .B(n1337), .Z(z2[428]) );
  NANDN U2001 ( .A(xregN_1), .B(zin[427]), .Z(n1337) );
  NAND U2002 ( .A(N432), .B(xregN_1), .Z(n1336) );
  NAND U2003 ( .A(n1338), .B(n1339), .Z(z2[427]) );
  NANDN U2004 ( .A(xregN_1), .B(zin[426]), .Z(n1339) );
  NAND U2005 ( .A(N431), .B(xregN_1), .Z(n1338) );
  NAND U2006 ( .A(n1340), .B(n1341), .Z(z2[426]) );
  NANDN U2007 ( .A(xregN_1), .B(zin[425]), .Z(n1341) );
  NAND U2008 ( .A(N430), .B(xregN_1), .Z(n1340) );
  NAND U2009 ( .A(n1342), .B(n1343), .Z(z2[425]) );
  NANDN U2010 ( .A(xregN_1), .B(zin[424]), .Z(n1343) );
  NAND U2011 ( .A(N429), .B(xregN_1), .Z(n1342) );
  NAND U2012 ( .A(n1344), .B(n1345), .Z(z2[424]) );
  NANDN U2013 ( .A(xregN_1), .B(zin[423]), .Z(n1345) );
  NAND U2014 ( .A(N428), .B(xregN_1), .Z(n1344) );
  NAND U2015 ( .A(n1346), .B(n1347), .Z(z2[423]) );
  NANDN U2016 ( .A(xregN_1), .B(zin[422]), .Z(n1347) );
  NAND U2017 ( .A(N427), .B(xregN_1), .Z(n1346) );
  NAND U2018 ( .A(n1348), .B(n1349), .Z(z2[422]) );
  NANDN U2019 ( .A(xregN_1), .B(zin[421]), .Z(n1349) );
  NAND U2020 ( .A(N426), .B(xregN_1), .Z(n1348) );
  NAND U2021 ( .A(n1350), .B(n1351), .Z(z2[421]) );
  NANDN U2022 ( .A(xregN_1), .B(zin[420]), .Z(n1351) );
  NAND U2023 ( .A(N425), .B(xregN_1), .Z(n1350) );
  NAND U2024 ( .A(n1352), .B(n1353), .Z(z2[420]) );
  NANDN U2025 ( .A(xregN_1), .B(zin[419]), .Z(n1353) );
  NAND U2026 ( .A(N424), .B(xregN_1), .Z(n1352) );
  NAND U2027 ( .A(n1354), .B(n1355), .Z(z2[41]) );
  NANDN U2028 ( .A(xregN_1), .B(zin[40]), .Z(n1355) );
  NAND U2029 ( .A(N45), .B(xregN_1), .Z(n1354) );
  NAND U2030 ( .A(n1356), .B(n1357), .Z(z2[419]) );
  NANDN U2031 ( .A(xregN_1), .B(zin[418]), .Z(n1357) );
  NAND U2032 ( .A(N423), .B(xregN_1), .Z(n1356) );
  NAND U2033 ( .A(n1358), .B(n1359), .Z(z2[418]) );
  NANDN U2034 ( .A(xregN_1), .B(zin[417]), .Z(n1359) );
  NAND U2035 ( .A(N422), .B(xregN_1), .Z(n1358) );
  NAND U2036 ( .A(n1360), .B(n1361), .Z(z2[417]) );
  NANDN U2037 ( .A(xregN_1), .B(zin[416]), .Z(n1361) );
  NAND U2038 ( .A(N421), .B(xregN_1), .Z(n1360) );
  NAND U2039 ( .A(n1362), .B(n1363), .Z(z2[416]) );
  NANDN U2040 ( .A(xregN_1), .B(zin[415]), .Z(n1363) );
  NAND U2041 ( .A(N420), .B(xregN_1), .Z(n1362) );
  NAND U2042 ( .A(n1364), .B(n1365), .Z(z2[415]) );
  NANDN U2043 ( .A(xregN_1), .B(zin[414]), .Z(n1365) );
  NAND U2044 ( .A(N419), .B(xregN_1), .Z(n1364) );
  NAND U2045 ( .A(n1366), .B(n1367), .Z(z2[414]) );
  NANDN U2046 ( .A(xregN_1), .B(zin[413]), .Z(n1367) );
  NAND U2047 ( .A(N418), .B(xregN_1), .Z(n1366) );
  NAND U2048 ( .A(n1368), .B(n1369), .Z(z2[413]) );
  NANDN U2049 ( .A(xregN_1), .B(zin[412]), .Z(n1369) );
  NAND U2050 ( .A(N417), .B(xregN_1), .Z(n1368) );
  NAND U2051 ( .A(n1370), .B(n1371), .Z(z2[412]) );
  NANDN U2052 ( .A(xregN_1), .B(zin[411]), .Z(n1371) );
  NAND U2053 ( .A(N416), .B(xregN_1), .Z(n1370) );
  NAND U2054 ( .A(n1372), .B(n1373), .Z(z2[411]) );
  NANDN U2055 ( .A(xregN_1), .B(zin[410]), .Z(n1373) );
  NAND U2056 ( .A(N415), .B(xregN_1), .Z(n1372) );
  NAND U2057 ( .A(n1374), .B(n1375), .Z(z2[410]) );
  NANDN U2058 ( .A(xregN_1), .B(zin[409]), .Z(n1375) );
  NAND U2059 ( .A(N414), .B(xregN_1), .Z(n1374) );
  NAND U2060 ( .A(n1376), .B(n1377), .Z(z2[40]) );
  NANDN U2061 ( .A(xregN_1), .B(zin[39]), .Z(n1377) );
  NAND U2062 ( .A(N44), .B(xregN_1), .Z(n1376) );
  NAND U2063 ( .A(n1378), .B(n1379), .Z(z2[409]) );
  NANDN U2064 ( .A(xregN_1), .B(zin[408]), .Z(n1379) );
  NAND U2065 ( .A(N413), .B(xregN_1), .Z(n1378) );
  NAND U2066 ( .A(n1380), .B(n1381), .Z(z2[408]) );
  NANDN U2067 ( .A(xregN_1), .B(zin[407]), .Z(n1381) );
  NAND U2068 ( .A(N412), .B(xregN_1), .Z(n1380) );
  NAND U2069 ( .A(n1382), .B(n1383), .Z(z2[407]) );
  NANDN U2070 ( .A(xregN_1), .B(zin[406]), .Z(n1383) );
  NAND U2071 ( .A(N411), .B(xregN_1), .Z(n1382) );
  NAND U2072 ( .A(n1384), .B(n1385), .Z(z2[406]) );
  NANDN U2073 ( .A(xregN_1), .B(zin[405]), .Z(n1385) );
  NAND U2074 ( .A(N410), .B(xregN_1), .Z(n1384) );
  NAND U2075 ( .A(n1386), .B(n1387), .Z(z2[405]) );
  NANDN U2076 ( .A(xregN_1), .B(zin[404]), .Z(n1387) );
  NAND U2077 ( .A(N409), .B(xregN_1), .Z(n1386) );
  NAND U2078 ( .A(n1388), .B(n1389), .Z(z2[404]) );
  NANDN U2079 ( .A(xregN_1), .B(zin[403]), .Z(n1389) );
  NAND U2080 ( .A(N408), .B(xregN_1), .Z(n1388) );
  NAND U2081 ( .A(n1390), .B(n1391), .Z(z2[403]) );
  NANDN U2082 ( .A(xregN_1), .B(zin[402]), .Z(n1391) );
  NAND U2083 ( .A(N407), .B(xregN_1), .Z(n1390) );
  NAND U2084 ( .A(n1392), .B(n1393), .Z(z2[402]) );
  NANDN U2085 ( .A(xregN_1), .B(zin[401]), .Z(n1393) );
  NAND U2086 ( .A(N406), .B(xregN_1), .Z(n1392) );
  NAND U2087 ( .A(n1394), .B(n1395), .Z(z2[401]) );
  NANDN U2088 ( .A(xregN_1), .B(zin[400]), .Z(n1395) );
  NAND U2089 ( .A(N405), .B(xregN_1), .Z(n1394) );
  NAND U2090 ( .A(n1396), .B(n1397), .Z(z2[400]) );
  NANDN U2091 ( .A(xregN_1), .B(zin[399]), .Z(n1397) );
  NAND U2092 ( .A(N404), .B(xregN_1), .Z(n1396) );
  NAND U2093 ( .A(n1398), .B(n1399), .Z(z2[3]) );
  NANDN U2094 ( .A(xregN_1), .B(zin[2]), .Z(n1399) );
  NAND U2095 ( .A(N7), .B(xregN_1), .Z(n1398) );
  NAND U2096 ( .A(n1400), .B(n1401), .Z(z2[39]) );
  NANDN U2097 ( .A(xregN_1), .B(zin[38]), .Z(n1401) );
  NAND U2098 ( .A(N43), .B(xregN_1), .Z(n1400) );
  NAND U2099 ( .A(n1402), .B(n1403), .Z(z2[399]) );
  NANDN U2100 ( .A(xregN_1), .B(zin[398]), .Z(n1403) );
  NAND U2101 ( .A(N403), .B(xregN_1), .Z(n1402) );
  NAND U2102 ( .A(n1404), .B(n1405), .Z(z2[398]) );
  NANDN U2103 ( .A(xregN_1), .B(zin[397]), .Z(n1405) );
  NAND U2104 ( .A(N402), .B(xregN_1), .Z(n1404) );
  NAND U2105 ( .A(n1406), .B(n1407), .Z(z2[397]) );
  NANDN U2106 ( .A(xregN_1), .B(zin[396]), .Z(n1407) );
  NAND U2107 ( .A(N401), .B(xregN_1), .Z(n1406) );
  NAND U2108 ( .A(n1408), .B(n1409), .Z(z2[396]) );
  NANDN U2109 ( .A(xregN_1), .B(zin[395]), .Z(n1409) );
  NAND U2110 ( .A(N400), .B(xregN_1), .Z(n1408) );
  NAND U2111 ( .A(n1410), .B(n1411), .Z(z2[395]) );
  NANDN U2112 ( .A(xregN_1), .B(zin[394]), .Z(n1411) );
  NAND U2113 ( .A(N399), .B(xregN_1), .Z(n1410) );
  NAND U2114 ( .A(n1412), .B(n1413), .Z(z2[394]) );
  NANDN U2115 ( .A(xregN_1), .B(zin[393]), .Z(n1413) );
  NAND U2116 ( .A(N398), .B(xregN_1), .Z(n1412) );
  NAND U2117 ( .A(n1414), .B(n1415), .Z(z2[393]) );
  NANDN U2118 ( .A(xregN_1), .B(zin[392]), .Z(n1415) );
  NAND U2119 ( .A(N397), .B(xregN_1), .Z(n1414) );
  NAND U2120 ( .A(n1416), .B(n1417), .Z(z2[392]) );
  NANDN U2121 ( .A(xregN_1), .B(zin[391]), .Z(n1417) );
  NAND U2122 ( .A(N396), .B(xregN_1), .Z(n1416) );
  NAND U2123 ( .A(n1418), .B(n1419), .Z(z2[391]) );
  NANDN U2124 ( .A(xregN_1), .B(zin[390]), .Z(n1419) );
  NAND U2125 ( .A(N395), .B(xregN_1), .Z(n1418) );
  NAND U2126 ( .A(n1420), .B(n1421), .Z(z2[390]) );
  NANDN U2127 ( .A(xregN_1), .B(zin[389]), .Z(n1421) );
  NAND U2128 ( .A(N394), .B(xregN_1), .Z(n1420) );
  NAND U2129 ( .A(n1422), .B(n1423), .Z(z2[38]) );
  NANDN U2130 ( .A(xregN_1), .B(zin[37]), .Z(n1423) );
  NAND U2131 ( .A(N42), .B(xregN_1), .Z(n1422) );
  NAND U2132 ( .A(n1424), .B(n1425), .Z(z2[389]) );
  NANDN U2133 ( .A(xregN_1), .B(zin[388]), .Z(n1425) );
  NAND U2134 ( .A(N393), .B(xregN_1), .Z(n1424) );
  NAND U2135 ( .A(n1426), .B(n1427), .Z(z2[388]) );
  NANDN U2136 ( .A(xregN_1), .B(zin[387]), .Z(n1427) );
  NAND U2137 ( .A(N392), .B(xregN_1), .Z(n1426) );
  NAND U2138 ( .A(n1428), .B(n1429), .Z(z2[387]) );
  NANDN U2139 ( .A(xregN_1), .B(zin[386]), .Z(n1429) );
  NAND U2140 ( .A(N391), .B(xregN_1), .Z(n1428) );
  NAND U2141 ( .A(n1430), .B(n1431), .Z(z2[386]) );
  NANDN U2142 ( .A(xregN_1), .B(zin[385]), .Z(n1431) );
  NAND U2143 ( .A(N390), .B(xregN_1), .Z(n1430) );
  NAND U2144 ( .A(n1432), .B(n1433), .Z(z2[385]) );
  NANDN U2145 ( .A(xregN_1), .B(zin[384]), .Z(n1433) );
  NAND U2146 ( .A(N389), .B(xregN_1), .Z(n1432) );
  NAND U2147 ( .A(n1434), .B(n1435), .Z(z2[384]) );
  NANDN U2148 ( .A(xregN_1), .B(zin[383]), .Z(n1435) );
  NAND U2149 ( .A(N388), .B(xregN_1), .Z(n1434) );
  NAND U2150 ( .A(n1436), .B(n1437), .Z(z2[383]) );
  NANDN U2151 ( .A(xregN_1), .B(zin[382]), .Z(n1437) );
  NAND U2152 ( .A(N387), .B(xregN_1), .Z(n1436) );
  NAND U2153 ( .A(n1438), .B(n1439), .Z(z2[382]) );
  NANDN U2154 ( .A(xregN_1), .B(zin[381]), .Z(n1439) );
  NAND U2155 ( .A(N386), .B(xregN_1), .Z(n1438) );
  NAND U2156 ( .A(n1440), .B(n1441), .Z(z2[381]) );
  NANDN U2157 ( .A(xregN_1), .B(zin[380]), .Z(n1441) );
  NAND U2158 ( .A(N385), .B(xregN_1), .Z(n1440) );
  NAND U2159 ( .A(n1442), .B(n1443), .Z(z2[380]) );
  NANDN U2160 ( .A(xregN_1), .B(zin[379]), .Z(n1443) );
  NAND U2161 ( .A(N384), .B(xregN_1), .Z(n1442) );
  NAND U2162 ( .A(n1444), .B(n1445), .Z(z2[37]) );
  NANDN U2163 ( .A(xregN_1), .B(zin[36]), .Z(n1445) );
  NAND U2164 ( .A(N41), .B(xregN_1), .Z(n1444) );
  NAND U2165 ( .A(n1446), .B(n1447), .Z(z2[379]) );
  NANDN U2166 ( .A(xregN_1), .B(zin[378]), .Z(n1447) );
  NAND U2167 ( .A(N383), .B(xregN_1), .Z(n1446) );
  NAND U2168 ( .A(n1448), .B(n1449), .Z(z2[378]) );
  NANDN U2169 ( .A(xregN_1), .B(zin[377]), .Z(n1449) );
  NAND U2170 ( .A(N382), .B(xregN_1), .Z(n1448) );
  NAND U2171 ( .A(n1450), .B(n1451), .Z(z2[377]) );
  NANDN U2172 ( .A(xregN_1), .B(zin[376]), .Z(n1451) );
  NAND U2173 ( .A(N381), .B(xregN_1), .Z(n1450) );
  NAND U2174 ( .A(n1452), .B(n1453), .Z(z2[376]) );
  NANDN U2175 ( .A(xregN_1), .B(zin[375]), .Z(n1453) );
  NAND U2176 ( .A(N380), .B(xregN_1), .Z(n1452) );
  NAND U2177 ( .A(n1454), .B(n1455), .Z(z2[375]) );
  NANDN U2178 ( .A(xregN_1), .B(zin[374]), .Z(n1455) );
  NAND U2179 ( .A(N379), .B(xregN_1), .Z(n1454) );
  NAND U2180 ( .A(n1456), .B(n1457), .Z(z2[374]) );
  NANDN U2181 ( .A(xregN_1), .B(zin[373]), .Z(n1457) );
  NAND U2182 ( .A(N378), .B(xregN_1), .Z(n1456) );
  NAND U2183 ( .A(n1458), .B(n1459), .Z(z2[373]) );
  NANDN U2184 ( .A(xregN_1), .B(zin[372]), .Z(n1459) );
  NAND U2185 ( .A(N377), .B(xregN_1), .Z(n1458) );
  NAND U2186 ( .A(n1460), .B(n1461), .Z(z2[372]) );
  NANDN U2187 ( .A(xregN_1), .B(zin[371]), .Z(n1461) );
  NAND U2188 ( .A(N376), .B(xregN_1), .Z(n1460) );
  NAND U2189 ( .A(n1462), .B(n1463), .Z(z2[371]) );
  NANDN U2190 ( .A(xregN_1), .B(zin[370]), .Z(n1463) );
  NAND U2191 ( .A(N375), .B(xregN_1), .Z(n1462) );
  NAND U2192 ( .A(n1464), .B(n1465), .Z(z2[370]) );
  NANDN U2193 ( .A(xregN_1), .B(zin[369]), .Z(n1465) );
  NAND U2194 ( .A(N374), .B(xregN_1), .Z(n1464) );
  NAND U2195 ( .A(n1466), .B(n1467), .Z(z2[36]) );
  NANDN U2196 ( .A(xregN_1), .B(zin[35]), .Z(n1467) );
  NAND U2197 ( .A(N40), .B(xregN_1), .Z(n1466) );
  NAND U2198 ( .A(n1468), .B(n1469), .Z(z2[369]) );
  NANDN U2199 ( .A(xregN_1), .B(zin[368]), .Z(n1469) );
  NAND U2200 ( .A(N373), .B(xregN_1), .Z(n1468) );
  NAND U2201 ( .A(n1470), .B(n1471), .Z(z2[368]) );
  NANDN U2202 ( .A(xregN_1), .B(zin[367]), .Z(n1471) );
  NAND U2203 ( .A(N372), .B(xregN_1), .Z(n1470) );
  NAND U2204 ( .A(n1472), .B(n1473), .Z(z2[367]) );
  NANDN U2205 ( .A(xregN_1), .B(zin[366]), .Z(n1473) );
  NAND U2206 ( .A(N371), .B(xregN_1), .Z(n1472) );
  NAND U2207 ( .A(n1474), .B(n1475), .Z(z2[366]) );
  NANDN U2208 ( .A(xregN_1), .B(zin[365]), .Z(n1475) );
  NAND U2209 ( .A(N370), .B(xregN_1), .Z(n1474) );
  NAND U2210 ( .A(n1476), .B(n1477), .Z(z2[365]) );
  NANDN U2211 ( .A(xregN_1), .B(zin[364]), .Z(n1477) );
  NAND U2212 ( .A(N369), .B(xregN_1), .Z(n1476) );
  NAND U2213 ( .A(n1478), .B(n1479), .Z(z2[364]) );
  NANDN U2214 ( .A(xregN_1), .B(zin[363]), .Z(n1479) );
  NAND U2215 ( .A(N368), .B(xregN_1), .Z(n1478) );
  NAND U2216 ( .A(n1480), .B(n1481), .Z(z2[363]) );
  NANDN U2217 ( .A(xregN_1), .B(zin[362]), .Z(n1481) );
  NAND U2218 ( .A(N367), .B(xregN_1), .Z(n1480) );
  NAND U2219 ( .A(n1482), .B(n1483), .Z(z2[362]) );
  NANDN U2220 ( .A(xregN_1), .B(zin[361]), .Z(n1483) );
  NAND U2221 ( .A(N366), .B(xregN_1), .Z(n1482) );
  NAND U2222 ( .A(n1484), .B(n1485), .Z(z2[361]) );
  NANDN U2223 ( .A(xregN_1), .B(zin[360]), .Z(n1485) );
  NAND U2224 ( .A(N365), .B(xregN_1), .Z(n1484) );
  NAND U2225 ( .A(n1486), .B(n1487), .Z(z2[360]) );
  NANDN U2226 ( .A(xregN_1), .B(zin[359]), .Z(n1487) );
  NAND U2227 ( .A(N364), .B(xregN_1), .Z(n1486) );
  NAND U2228 ( .A(n1488), .B(n1489), .Z(z2[35]) );
  NANDN U2229 ( .A(xregN_1), .B(zin[34]), .Z(n1489) );
  NAND U2230 ( .A(N39), .B(xregN_1), .Z(n1488) );
  NAND U2231 ( .A(n1490), .B(n1491), .Z(z2[359]) );
  NANDN U2232 ( .A(xregN_1), .B(zin[358]), .Z(n1491) );
  NAND U2233 ( .A(N363), .B(xregN_1), .Z(n1490) );
  NAND U2234 ( .A(n1492), .B(n1493), .Z(z2[358]) );
  NANDN U2235 ( .A(xregN_1), .B(zin[357]), .Z(n1493) );
  NAND U2236 ( .A(N362), .B(xregN_1), .Z(n1492) );
  NAND U2237 ( .A(n1494), .B(n1495), .Z(z2[357]) );
  NANDN U2238 ( .A(xregN_1), .B(zin[356]), .Z(n1495) );
  NAND U2239 ( .A(N361), .B(xregN_1), .Z(n1494) );
  NAND U2240 ( .A(n1496), .B(n1497), .Z(z2[356]) );
  NANDN U2241 ( .A(xregN_1), .B(zin[355]), .Z(n1497) );
  NAND U2242 ( .A(N360), .B(xregN_1), .Z(n1496) );
  NAND U2243 ( .A(n1498), .B(n1499), .Z(z2[355]) );
  NANDN U2244 ( .A(xregN_1), .B(zin[354]), .Z(n1499) );
  NAND U2245 ( .A(N359), .B(xregN_1), .Z(n1498) );
  NAND U2246 ( .A(n1500), .B(n1501), .Z(z2[354]) );
  NANDN U2247 ( .A(xregN_1), .B(zin[353]), .Z(n1501) );
  NAND U2248 ( .A(N358), .B(xregN_1), .Z(n1500) );
  NAND U2249 ( .A(n1502), .B(n1503), .Z(z2[353]) );
  NANDN U2250 ( .A(xregN_1), .B(zin[352]), .Z(n1503) );
  NAND U2251 ( .A(N357), .B(xregN_1), .Z(n1502) );
  NAND U2252 ( .A(n1504), .B(n1505), .Z(z2[352]) );
  NANDN U2253 ( .A(xregN_1), .B(zin[351]), .Z(n1505) );
  NAND U2254 ( .A(N356), .B(xregN_1), .Z(n1504) );
  NAND U2255 ( .A(n1506), .B(n1507), .Z(z2[351]) );
  NANDN U2256 ( .A(xregN_1), .B(zin[350]), .Z(n1507) );
  NAND U2257 ( .A(N355), .B(xregN_1), .Z(n1506) );
  NAND U2258 ( .A(n1508), .B(n1509), .Z(z2[350]) );
  NANDN U2259 ( .A(xregN_1), .B(zin[349]), .Z(n1509) );
  NAND U2260 ( .A(N354), .B(xregN_1), .Z(n1508) );
  NAND U2261 ( .A(n1510), .B(n1511), .Z(z2[34]) );
  NANDN U2262 ( .A(xregN_1), .B(zin[33]), .Z(n1511) );
  NAND U2263 ( .A(N38), .B(xregN_1), .Z(n1510) );
  NAND U2264 ( .A(n1512), .B(n1513), .Z(z2[349]) );
  NANDN U2265 ( .A(xregN_1), .B(zin[348]), .Z(n1513) );
  NAND U2266 ( .A(N353), .B(xregN_1), .Z(n1512) );
  NAND U2267 ( .A(n1514), .B(n1515), .Z(z2[348]) );
  NANDN U2268 ( .A(xregN_1), .B(zin[347]), .Z(n1515) );
  NAND U2269 ( .A(N352), .B(xregN_1), .Z(n1514) );
  NAND U2270 ( .A(n1516), .B(n1517), .Z(z2[347]) );
  NANDN U2271 ( .A(xregN_1), .B(zin[346]), .Z(n1517) );
  NAND U2272 ( .A(N351), .B(xregN_1), .Z(n1516) );
  NAND U2273 ( .A(n1518), .B(n1519), .Z(z2[346]) );
  NANDN U2274 ( .A(xregN_1), .B(zin[345]), .Z(n1519) );
  NAND U2275 ( .A(N350), .B(xregN_1), .Z(n1518) );
  NAND U2276 ( .A(n1520), .B(n1521), .Z(z2[345]) );
  NANDN U2277 ( .A(xregN_1), .B(zin[344]), .Z(n1521) );
  NAND U2278 ( .A(N349), .B(xregN_1), .Z(n1520) );
  NAND U2279 ( .A(n1522), .B(n1523), .Z(z2[344]) );
  NANDN U2280 ( .A(xregN_1), .B(zin[343]), .Z(n1523) );
  NAND U2281 ( .A(N348), .B(xregN_1), .Z(n1522) );
  NAND U2282 ( .A(n1524), .B(n1525), .Z(z2[343]) );
  NANDN U2283 ( .A(xregN_1), .B(zin[342]), .Z(n1525) );
  NAND U2284 ( .A(N347), .B(xregN_1), .Z(n1524) );
  NAND U2285 ( .A(n1526), .B(n1527), .Z(z2[342]) );
  NANDN U2286 ( .A(xregN_1), .B(zin[341]), .Z(n1527) );
  NAND U2287 ( .A(N346), .B(xregN_1), .Z(n1526) );
  NAND U2288 ( .A(n1528), .B(n1529), .Z(z2[341]) );
  NANDN U2289 ( .A(xregN_1), .B(zin[340]), .Z(n1529) );
  NAND U2290 ( .A(N345), .B(xregN_1), .Z(n1528) );
  NAND U2291 ( .A(n1530), .B(n1531), .Z(z2[340]) );
  NANDN U2292 ( .A(xregN_1), .B(zin[339]), .Z(n1531) );
  NAND U2293 ( .A(N344), .B(xregN_1), .Z(n1530) );
  NAND U2294 ( .A(n1532), .B(n1533), .Z(z2[33]) );
  NANDN U2295 ( .A(xregN_1), .B(zin[32]), .Z(n1533) );
  NAND U2296 ( .A(N37), .B(xregN_1), .Z(n1532) );
  NAND U2297 ( .A(n1534), .B(n1535), .Z(z2[339]) );
  NANDN U2298 ( .A(xregN_1), .B(zin[338]), .Z(n1535) );
  NAND U2299 ( .A(N343), .B(xregN_1), .Z(n1534) );
  NAND U2300 ( .A(n1536), .B(n1537), .Z(z2[338]) );
  NANDN U2301 ( .A(xregN_1), .B(zin[337]), .Z(n1537) );
  NAND U2302 ( .A(N342), .B(xregN_1), .Z(n1536) );
  NAND U2303 ( .A(n1538), .B(n1539), .Z(z2[337]) );
  NANDN U2304 ( .A(xregN_1), .B(zin[336]), .Z(n1539) );
  NAND U2305 ( .A(N341), .B(xregN_1), .Z(n1538) );
  NAND U2306 ( .A(n1540), .B(n1541), .Z(z2[336]) );
  NANDN U2307 ( .A(xregN_1), .B(zin[335]), .Z(n1541) );
  NAND U2308 ( .A(N340), .B(xregN_1), .Z(n1540) );
  NAND U2309 ( .A(n1542), .B(n1543), .Z(z2[335]) );
  NANDN U2310 ( .A(xregN_1), .B(zin[334]), .Z(n1543) );
  NAND U2311 ( .A(N339), .B(xregN_1), .Z(n1542) );
  NAND U2312 ( .A(n1544), .B(n1545), .Z(z2[334]) );
  NANDN U2313 ( .A(xregN_1), .B(zin[333]), .Z(n1545) );
  NAND U2314 ( .A(N338), .B(xregN_1), .Z(n1544) );
  NAND U2315 ( .A(n1546), .B(n1547), .Z(z2[333]) );
  NANDN U2316 ( .A(xregN_1), .B(zin[332]), .Z(n1547) );
  NAND U2317 ( .A(N337), .B(xregN_1), .Z(n1546) );
  NAND U2318 ( .A(n1548), .B(n1549), .Z(z2[332]) );
  NANDN U2319 ( .A(xregN_1), .B(zin[331]), .Z(n1549) );
  NAND U2320 ( .A(N336), .B(xregN_1), .Z(n1548) );
  NAND U2321 ( .A(n1550), .B(n1551), .Z(z2[331]) );
  NANDN U2322 ( .A(xregN_1), .B(zin[330]), .Z(n1551) );
  NAND U2323 ( .A(N335), .B(xregN_1), .Z(n1550) );
  NAND U2324 ( .A(n1552), .B(n1553), .Z(z2[330]) );
  NANDN U2325 ( .A(xregN_1), .B(zin[329]), .Z(n1553) );
  NAND U2326 ( .A(N334), .B(xregN_1), .Z(n1552) );
  NAND U2327 ( .A(n1554), .B(n1555), .Z(z2[32]) );
  NANDN U2328 ( .A(xregN_1), .B(zin[31]), .Z(n1555) );
  NAND U2329 ( .A(N36), .B(xregN_1), .Z(n1554) );
  NAND U2330 ( .A(n1556), .B(n1557), .Z(z2[329]) );
  NANDN U2331 ( .A(xregN_1), .B(zin[328]), .Z(n1557) );
  NAND U2332 ( .A(N333), .B(xregN_1), .Z(n1556) );
  NAND U2333 ( .A(n1558), .B(n1559), .Z(z2[328]) );
  NANDN U2334 ( .A(xregN_1), .B(zin[327]), .Z(n1559) );
  NAND U2335 ( .A(N332), .B(xregN_1), .Z(n1558) );
  NAND U2336 ( .A(n1560), .B(n1561), .Z(z2[327]) );
  NANDN U2337 ( .A(xregN_1), .B(zin[326]), .Z(n1561) );
  NAND U2338 ( .A(N331), .B(xregN_1), .Z(n1560) );
  NAND U2339 ( .A(n1562), .B(n1563), .Z(z2[326]) );
  NANDN U2340 ( .A(xregN_1), .B(zin[325]), .Z(n1563) );
  NAND U2341 ( .A(N330), .B(xregN_1), .Z(n1562) );
  NAND U2342 ( .A(n1564), .B(n1565), .Z(z2[325]) );
  NANDN U2343 ( .A(xregN_1), .B(zin[324]), .Z(n1565) );
  NAND U2344 ( .A(N329), .B(xregN_1), .Z(n1564) );
  NAND U2345 ( .A(n1566), .B(n1567), .Z(z2[324]) );
  NANDN U2346 ( .A(xregN_1), .B(zin[323]), .Z(n1567) );
  NAND U2347 ( .A(N328), .B(xregN_1), .Z(n1566) );
  NAND U2348 ( .A(n1568), .B(n1569), .Z(z2[323]) );
  NANDN U2349 ( .A(xregN_1), .B(zin[322]), .Z(n1569) );
  NAND U2350 ( .A(N327), .B(xregN_1), .Z(n1568) );
  NAND U2351 ( .A(n1570), .B(n1571), .Z(z2[322]) );
  NANDN U2352 ( .A(xregN_1), .B(zin[321]), .Z(n1571) );
  NAND U2353 ( .A(N326), .B(xregN_1), .Z(n1570) );
  NAND U2354 ( .A(n1572), .B(n1573), .Z(z2[321]) );
  NANDN U2355 ( .A(xregN_1), .B(zin[320]), .Z(n1573) );
  NAND U2356 ( .A(N325), .B(xregN_1), .Z(n1572) );
  NAND U2357 ( .A(n1574), .B(n1575), .Z(z2[320]) );
  NANDN U2358 ( .A(xregN_1), .B(zin[319]), .Z(n1575) );
  NAND U2359 ( .A(N324), .B(xregN_1), .Z(n1574) );
  NAND U2360 ( .A(n1576), .B(n1577), .Z(z2[31]) );
  NANDN U2361 ( .A(xregN_1), .B(zin[30]), .Z(n1577) );
  NAND U2362 ( .A(N35), .B(xregN_1), .Z(n1576) );
  NAND U2363 ( .A(n1578), .B(n1579), .Z(z2[319]) );
  NANDN U2364 ( .A(xregN_1), .B(zin[318]), .Z(n1579) );
  NAND U2365 ( .A(N323), .B(xregN_1), .Z(n1578) );
  NAND U2366 ( .A(n1580), .B(n1581), .Z(z2[318]) );
  NANDN U2367 ( .A(xregN_1), .B(zin[317]), .Z(n1581) );
  NAND U2368 ( .A(N322), .B(xregN_1), .Z(n1580) );
  NAND U2369 ( .A(n1582), .B(n1583), .Z(z2[317]) );
  NANDN U2370 ( .A(xregN_1), .B(zin[316]), .Z(n1583) );
  NAND U2371 ( .A(N321), .B(xregN_1), .Z(n1582) );
  NAND U2372 ( .A(n1584), .B(n1585), .Z(z2[316]) );
  NANDN U2373 ( .A(xregN_1), .B(zin[315]), .Z(n1585) );
  NAND U2374 ( .A(N320), .B(xregN_1), .Z(n1584) );
  NAND U2375 ( .A(n1586), .B(n1587), .Z(z2[315]) );
  NANDN U2376 ( .A(xregN_1), .B(zin[314]), .Z(n1587) );
  NAND U2377 ( .A(N319), .B(xregN_1), .Z(n1586) );
  NAND U2378 ( .A(n1588), .B(n1589), .Z(z2[314]) );
  NANDN U2379 ( .A(xregN_1), .B(zin[313]), .Z(n1589) );
  NAND U2380 ( .A(N318), .B(xregN_1), .Z(n1588) );
  NAND U2381 ( .A(n1590), .B(n1591), .Z(z2[313]) );
  NANDN U2382 ( .A(xregN_1), .B(zin[312]), .Z(n1591) );
  NAND U2383 ( .A(N317), .B(xregN_1), .Z(n1590) );
  NAND U2384 ( .A(n1592), .B(n1593), .Z(z2[312]) );
  NANDN U2385 ( .A(xregN_1), .B(zin[311]), .Z(n1593) );
  NAND U2386 ( .A(N316), .B(xregN_1), .Z(n1592) );
  NAND U2387 ( .A(n1594), .B(n1595), .Z(z2[311]) );
  NANDN U2388 ( .A(xregN_1), .B(zin[310]), .Z(n1595) );
  NAND U2389 ( .A(N315), .B(xregN_1), .Z(n1594) );
  NAND U2390 ( .A(n1596), .B(n1597), .Z(z2[310]) );
  NANDN U2391 ( .A(xregN_1), .B(zin[309]), .Z(n1597) );
  NAND U2392 ( .A(N314), .B(xregN_1), .Z(n1596) );
  NAND U2393 ( .A(n1598), .B(n1599), .Z(z2[30]) );
  NANDN U2394 ( .A(xregN_1), .B(zin[29]), .Z(n1599) );
  NAND U2395 ( .A(N34), .B(xregN_1), .Z(n1598) );
  NAND U2396 ( .A(n1600), .B(n1601), .Z(z2[309]) );
  NANDN U2397 ( .A(xregN_1), .B(zin[308]), .Z(n1601) );
  NAND U2398 ( .A(N313), .B(xregN_1), .Z(n1600) );
  NAND U2399 ( .A(n1602), .B(n1603), .Z(z2[308]) );
  NANDN U2400 ( .A(xregN_1), .B(zin[307]), .Z(n1603) );
  NAND U2401 ( .A(N312), .B(xregN_1), .Z(n1602) );
  NAND U2402 ( .A(n1604), .B(n1605), .Z(z2[307]) );
  NANDN U2403 ( .A(xregN_1), .B(zin[306]), .Z(n1605) );
  NAND U2404 ( .A(N311), .B(xregN_1), .Z(n1604) );
  NAND U2405 ( .A(n1606), .B(n1607), .Z(z2[306]) );
  NANDN U2406 ( .A(xregN_1), .B(zin[305]), .Z(n1607) );
  NAND U2407 ( .A(N310), .B(xregN_1), .Z(n1606) );
  NAND U2408 ( .A(n1608), .B(n1609), .Z(z2[305]) );
  NANDN U2409 ( .A(xregN_1), .B(zin[304]), .Z(n1609) );
  NAND U2410 ( .A(N309), .B(xregN_1), .Z(n1608) );
  NAND U2411 ( .A(n1610), .B(n1611), .Z(z2[304]) );
  NANDN U2412 ( .A(xregN_1), .B(zin[303]), .Z(n1611) );
  NAND U2413 ( .A(N308), .B(xregN_1), .Z(n1610) );
  NAND U2414 ( .A(n1612), .B(n1613), .Z(z2[303]) );
  NANDN U2415 ( .A(xregN_1), .B(zin[302]), .Z(n1613) );
  NAND U2416 ( .A(N307), .B(xregN_1), .Z(n1612) );
  NAND U2417 ( .A(n1614), .B(n1615), .Z(z2[302]) );
  NANDN U2418 ( .A(xregN_1), .B(zin[301]), .Z(n1615) );
  NAND U2419 ( .A(N306), .B(xregN_1), .Z(n1614) );
  NAND U2420 ( .A(n1616), .B(n1617), .Z(z2[301]) );
  NANDN U2421 ( .A(xregN_1), .B(zin[300]), .Z(n1617) );
  NAND U2422 ( .A(N305), .B(xregN_1), .Z(n1616) );
  NAND U2423 ( .A(n1618), .B(n1619), .Z(z2[300]) );
  NANDN U2424 ( .A(xregN_1), .B(zin[299]), .Z(n1619) );
  NAND U2425 ( .A(N304), .B(xregN_1), .Z(n1618) );
  NAND U2426 ( .A(n1620), .B(n1621), .Z(z2[2]) );
  NANDN U2427 ( .A(xregN_1), .B(zin[1]), .Z(n1621) );
  NAND U2428 ( .A(N6), .B(xregN_1), .Z(n1620) );
  NAND U2429 ( .A(n1622), .B(n1623), .Z(z2[29]) );
  NANDN U2430 ( .A(xregN_1), .B(zin[28]), .Z(n1623) );
  NAND U2431 ( .A(N33), .B(xregN_1), .Z(n1622) );
  NAND U2432 ( .A(n1624), .B(n1625), .Z(z2[299]) );
  NANDN U2433 ( .A(xregN_1), .B(zin[298]), .Z(n1625) );
  NAND U2434 ( .A(N303), .B(xregN_1), .Z(n1624) );
  NAND U2435 ( .A(n1626), .B(n1627), .Z(z2[298]) );
  NANDN U2436 ( .A(xregN_1), .B(zin[297]), .Z(n1627) );
  NAND U2437 ( .A(N302), .B(xregN_1), .Z(n1626) );
  NAND U2438 ( .A(n1628), .B(n1629), .Z(z2[297]) );
  NANDN U2439 ( .A(xregN_1), .B(zin[296]), .Z(n1629) );
  NAND U2440 ( .A(N301), .B(xregN_1), .Z(n1628) );
  NAND U2441 ( .A(n1630), .B(n1631), .Z(z2[296]) );
  NANDN U2442 ( .A(xregN_1), .B(zin[295]), .Z(n1631) );
  NAND U2443 ( .A(N300), .B(xregN_1), .Z(n1630) );
  NAND U2444 ( .A(n1632), .B(n1633), .Z(z2[295]) );
  NANDN U2445 ( .A(xregN_1), .B(zin[294]), .Z(n1633) );
  NAND U2446 ( .A(N299), .B(xregN_1), .Z(n1632) );
  NAND U2447 ( .A(n1634), .B(n1635), .Z(z2[294]) );
  NANDN U2448 ( .A(xregN_1), .B(zin[293]), .Z(n1635) );
  NAND U2449 ( .A(N298), .B(xregN_1), .Z(n1634) );
  NAND U2450 ( .A(n1636), .B(n1637), .Z(z2[293]) );
  NANDN U2451 ( .A(xregN_1), .B(zin[292]), .Z(n1637) );
  NAND U2452 ( .A(N297), .B(xregN_1), .Z(n1636) );
  NAND U2453 ( .A(n1638), .B(n1639), .Z(z2[292]) );
  NANDN U2454 ( .A(xregN_1), .B(zin[291]), .Z(n1639) );
  NAND U2455 ( .A(N296), .B(xregN_1), .Z(n1638) );
  NAND U2456 ( .A(n1640), .B(n1641), .Z(z2[291]) );
  NANDN U2457 ( .A(xregN_1), .B(zin[290]), .Z(n1641) );
  NAND U2458 ( .A(N295), .B(xregN_1), .Z(n1640) );
  NAND U2459 ( .A(n1642), .B(n1643), .Z(z2[290]) );
  NANDN U2460 ( .A(xregN_1), .B(zin[289]), .Z(n1643) );
  NAND U2461 ( .A(N294), .B(xregN_1), .Z(n1642) );
  NAND U2462 ( .A(n1644), .B(n1645), .Z(z2[28]) );
  NANDN U2463 ( .A(xregN_1), .B(zin[27]), .Z(n1645) );
  NAND U2464 ( .A(N32), .B(xregN_1), .Z(n1644) );
  NAND U2465 ( .A(n1646), .B(n1647), .Z(z2[289]) );
  NANDN U2466 ( .A(xregN_1), .B(zin[288]), .Z(n1647) );
  NAND U2467 ( .A(N293), .B(xregN_1), .Z(n1646) );
  NAND U2468 ( .A(n1648), .B(n1649), .Z(z2[288]) );
  NANDN U2469 ( .A(xregN_1), .B(zin[287]), .Z(n1649) );
  NAND U2470 ( .A(N292), .B(xregN_1), .Z(n1648) );
  NAND U2471 ( .A(n1650), .B(n1651), .Z(z2[287]) );
  NANDN U2472 ( .A(xregN_1), .B(zin[286]), .Z(n1651) );
  NAND U2473 ( .A(N291), .B(xregN_1), .Z(n1650) );
  NAND U2474 ( .A(n1652), .B(n1653), .Z(z2[286]) );
  NANDN U2475 ( .A(xregN_1), .B(zin[285]), .Z(n1653) );
  NAND U2476 ( .A(N290), .B(xregN_1), .Z(n1652) );
  NAND U2477 ( .A(n1654), .B(n1655), .Z(z2[285]) );
  NANDN U2478 ( .A(xregN_1), .B(zin[284]), .Z(n1655) );
  NAND U2479 ( .A(N289), .B(xregN_1), .Z(n1654) );
  NAND U2480 ( .A(n1656), .B(n1657), .Z(z2[284]) );
  NANDN U2481 ( .A(xregN_1), .B(zin[283]), .Z(n1657) );
  NAND U2482 ( .A(N288), .B(xregN_1), .Z(n1656) );
  NAND U2483 ( .A(n1658), .B(n1659), .Z(z2[283]) );
  NANDN U2484 ( .A(xregN_1), .B(zin[282]), .Z(n1659) );
  NAND U2485 ( .A(N287), .B(xregN_1), .Z(n1658) );
  NAND U2486 ( .A(n1660), .B(n1661), .Z(z2[282]) );
  NANDN U2487 ( .A(xregN_1), .B(zin[281]), .Z(n1661) );
  NAND U2488 ( .A(N286), .B(xregN_1), .Z(n1660) );
  NAND U2489 ( .A(n1662), .B(n1663), .Z(z2[281]) );
  NANDN U2490 ( .A(xregN_1), .B(zin[280]), .Z(n1663) );
  NAND U2491 ( .A(N285), .B(xregN_1), .Z(n1662) );
  NAND U2492 ( .A(n1664), .B(n1665), .Z(z2[280]) );
  NANDN U2493 ( .A(xregN_1), .B(zin[279]), .Z(n1665) );
  NAND U2494 ( .A(N284), .B(xregN_1), .Z(n1664) );
  NAND U2495 ( .A(n1666), .B(n1667), .Z(z2[27]) );
  NANDN U2496 ( .A(xregN_1), .B(zin[26]), .Z(n1667) );
  NAND U2497 ( .A(N31), .B(xregN_1), .Z(n1666) );
  NAND U2498 ( .A(n1668), .B(n1669), .Z(z2[279]) );
  NANDN U2499 ( .A(xregN_1), .B(zin[278]), .Z(n1669) );
  NAND U2500 ( .A(N283), .B(xregN_1), .Z(n1668) );
  NAND U2501 ( .A(n1670), .B(n1671), .Z(z2[278]) );
  NANDN U2502 ( .A(xregN_1), .B(zin[277]), .Z(n1671) );
  NAND U2503 ( .A(N282), .B(xregN_1), .Z(n1670) );
  NAND U2504 ( .A(n1672), .B(n1673), .Z(z2[277]) );
  NANDN U2505 ( .A(xregN_1), .B(zin[276]), .Z(n1673) );
  NAND U2506 ( .A(N281), .B(xregN_1), .Z(n1672) );
  NAND U2507 ( .A(n1674), .B(n1675), .Z(z2[276]) );
  NANDN U2508 ( .A(xregN_1), .B(zin[275]), .Z(n1675) );
  NAND U2509 ( .A(N280), .B(xregN_1), .Z(n1674) );
  NAND U2510 ( .A(n1676), .B(n1677), .Z(z2[275]) );
  NANDN U2511 ( .A(xregN_1), .B(zin[274]), .Z(n1677) );
  NAND U2512 ( .A(N279), .B(xregN_1), .Z(n1676) );
  NAND U2513 ( .A(n1678), .B(n1679), .Z(z2[274]) );
  NANDN U2514 ( .A(xregN_1), .B(zin[273]), .Z(n1679) );
  NAND U2515 ( .A(N278), .B(xregN_1), .Z(n1678) );
  NAND U2516 ( .A(n1680), .B(n1681), .Z(z2[273]) );
  NANDN U2517 ( .A(xregN_1), .B(zin[272]), .Z(n1681) );
  NAND U2518 ( .A(N277), .B(xregN_1), .Z(n1680) );
  NAND U2519 ( .A(n1682), .B(n1683), .Z(z2[272]) );
  NANDN U2520 ( .A(xregN_1), .B(zin[271]), .Z(n1683) );
  NAND U2521 ( .A(N276), .B(xregN_1), .Z(n1682) );
  NAND U2522 ( .A(n1684), .B(n1685), .Z(z2[271]) );
  NANDN U2523 ( .A(xregN_1), .B(zin[270]), .Z(n1685) );
  NAND U2524 ( .A(N275), .B(xregN_1), .Z(n1684) );
  NAND U2525 ( .A(n1686), .B(n1687), .Z(z2[270]) );
  NANDN U2526 ( .A(xregN_1), .B(zin[269]), .Z(n1687) );
  NAND U2527 ( .A(N274), .B(xregN_1), .Z(n1686) );
  NAND U2528 ( .A(n1688), .B(n1689), .Z(z2[26]) );
  NANDN U2529 ( .A(xregN_1), .B(zin[25]), .Z(n1689) );
  NAND U2530 ( .A(N30), .B(xregN_1), .Z(n1688) );
  NAND U2531 ( .A(n1690), .B(n1691), .Z(z2[269]) );
  NANDN U2532 ( .A(xregN_1), .B(zin[268]), .Z(n1691) );
  NAND U2533 ( .A(N273), .B(xregN_1), .Z(n1690) );
  NAND U2534 ( .A(n1692), .B(n1693), .Z(z2[268]) );
  NANDN U2535 ( .A(xregN_1), .B(zin[267]), .Z(n1693) );
  NAND U2536 ( .A(N272), .B(xregN_1), .Z(n1692) );
  NAND U2537 ( .A(n1694), .B(n1695), .Z(z2[267]) );
  NANDN U2538 ( .A(xregN_1), .B(zin[266]), .Z(n1695) );
  NAND U2539 ( .A(N271), .B(xregN_1), .Z(n1694) );
  NAND U2540 ( .A(n1696), .B(n1697), .Z(z2[266]) );
  NANDN U2541 ( .A(xregN_1), .B(zin[265]), .Z(n1697) );
  NAND U2542 ( .A(N270), .B(xregN_1), .Z(n1696) );
  NAND U2543 ( .A(n1698), .B(n1699), .Z(z2[265]) );
  NANDN U2544 ( .A(xregN_1), .B(zin[264]), .Z(n1699) );
  NAND U2545 ( .A(N269), .B(xregN_1), .Z(n1698) );
  NAND U2546 ( .A(n1700), .B(n1701), .Z(z2[264]) );
  NANDN U2547 ( .A(xregN_1), .B(zin[263]), .Z(n1701) );
  NAND U2548 ( .A(N268), .B(xregN_1), .Z(n1700) );
  NAND U2549 ( .A(n1702), .B(n1703), .Z(z2[263]) );
  NANDN U2550 ( .A(xregN_1), .B(zin[262]), .Z(n1703) );
  NAND U2551 ( .A(N267), .B(xregN_1), .Z(n1702) );
  NAND U2552 ( .A(n1704), .B(n1705), .Z(z2[262]) );
  NANDN U2553 ( .A(xregN_1), .B(zin[261]), .Z(n1705) );
  NAND U2554 ( .A(N266), .B(xregN_1), .Z(n1704) );
  NAND U2555 ( .A(n1706), .B(n1707), .Z(z2[261]) );
  NANDN U2556 ( .A(xregN_1), .B(zin[260]), .Z(n1707) );
  NAND U2557 ( .A(N265), .B(xregN_1), .Z(n1706) );
  NAND U2558 ( .A(n1708), .B(n1709), .Z(z2[260]) );
  NANDN U2559 ( .A(xregN_1), .B(zin[259]), .Z(n1709) );
  NAND U2560 ( .A(N264), .B(xregN_1), .Z(n1708) );
  NAND U2561 ( .A(n1710), .B(n1711), .Z(z2[25]) );
  NANDN U2562 ( .A(xregN_1), .B(zin[24]), .Z(n1711) );
  NAND U2563 ( .A(N29), .B(xregN_1), .Z(n1710) );
  NAND U2564 ( .A(n1712), .B(n1713), .Z(z2[259]) );
  NANDN U2565 ( .A(xregN_1), .B(zin[258]), .Z(n1713) );
  NAND U2566 ( .A(N263), .B(xregN_1), .Z(n1712) );
  NAND U2567 ( .A(n1714), .B(n1715), .Z(z2[258]) );
  NANDN U2568 ( .A(xregN_1), .B(zin[257]), .Z(n1715) );
  NAND U2569 ( .A(N262), .B(xregN_1), .Z(n1714) );
  NAND U2570 ( .A(n1716), .B(n1717), .Z(z2[257]) );
  NANDN U2571 ( .A(xregN_1), .B(zin[256]), .Z(n1717) );
  NAND U2572 ( .A(N261), .B(xregN_1), .Z(n1716) );
  NAND U2573 ( .A(n1718), .B(n1719), .Z(z2[256]) );
  NANDN U2574 ( .A(xregN_1), .B(zin[255]), .Z(n1719) );
  NAND U2575 ( .A(N260), .B(xregN_1), .Z(n1718) );
  NAND U2576 ( .A(n1720), .B(n1721), .Z(z2[255]) );
  NANDN U2577 ( .A(xregN_1), .B(zin[254]), .Z(n1721) );
  NAND U2578 ( .A(N259), .B(xregN_1), .Z(n1720) );
  NAND U2579 ( .A(n1722), .B(n1723), .Z(z2[254]) );
  NANDN U2580 ( .A(xregN_1), .B(zin[253]), .Z(n1723) );
  NAND U2581 ( .A(N258), .B(xregN_1), .Z(n1722) );
  NAND U2582 ( .A(n1724), .B(n1725), .Z(z2[253]) );
  NANDN U2583 ( .A(xregN_1), .B(zin[252]), .Z(n1725) );
  NAND U2584 ( .A(N257), .B(xregN_1), .Z(n1724) );
  NAND U2585 ( .A(n1726), .B(n1727), .Z(z2[252]) );
  NANDN U2586 ( .A(xregN_1), .B(zin[251]), .Z(n1727) );
  NAND U2587 ( .A(N256), .B(xregN_1), .Z(n1726) );
  NAND U2588 ( .A(n1728), .B(n1729), .Z(z2[251]) );
  NANDN U2589 ( .A(xregN_1), .B(zin[250]), .Z(n1729) );
  NAND U2590 ( .A(N255), .B(xregN_1), .Z(n1728) );
  NAND U2591 ( .A(n1730), .B(n1731), .Z(z2[250]) );
  NANDN U2592 ( .A(xregN_1), .B(zin[249]), .Z(n1731) );
  NAND U2593 ( .A(N254), .B(xregN_1), .Z(n1730) );
  NAND U2594 ( .A(n1732), .B(n1733), .Z(z2[24]) );
  NANDN U2595 ( .A(xregN_1), .B(zin[23]), .Z(n1733) );
  NAND U2596 ( .A(N28), .B(xregN_1), .Z(n1732) );
  NAND U2597 ( .A(n1734), .B(n1735), .Z(z2[249]) );
  NANDN U2598 ( .A(xregN_1), .B(zin[248]), .Z(n1735) );
  NAND U2599 ( .A(N253), .B(xregN_1), .Z(n1734) );
  NAND U2600 ( .A(n1736), .B(n1737), .Z(z2[248]) );
  NANDN U2601 ( .A(xregN_1), .B(zin[247]), .Z(n1737) );
  NAND U2602 ( .A(N252), .B(xregN_1), .Z(n1736) );
  NAND U2603 ( .A(n1738), .B(n1739), .Z(z2[247]) );
  NANDN U2604 ( .A(xregN_1), .B(zin[246]), .Z(n1739) );
  NAND U2605 ( .A(N251), .B(xregN_1), .Z(n1738) );
  NAND U2606 ( .A(n1740), .B(n1741), .Z(z2[246]) );
  NANDN U2607 ( .A(xregN_1), .B(zin[245]), .Z(n1741) );
  NAND U2608 ( .A(N250), .B(xregN_1), .Z(n1740) );
  NAND U2609 ( .A(n1742), .B(n1743), .Z(z2[245]) );
  NANDN U2610 ( .A(xregN_1), .B(zin[244]), .Z(n1743) );
  NAND U2611 ( .A(N249), .B(xregN_1), .Z(n1742) );
  NAND U2612 ( .A(n1744), .B(n1745), .Z(z2[244]) );
  NANDN U2613 ( .A(xregN_1), .B(zin[243]), .Z(n1745) );
  NAND U2614 ( .A(N248), .B(xregN_1), .Z(n1744) );
  NAND U2615 ( .A(n1746), .B(n1747), .Z(z2[243]) );
  NANDN U2616 ( .A(xregN_1), .B(zin[242]), .Z(n1747) );
  NAND U2617 ( .A(N247), .B(xregN_1), .Z(n1746) );
  NAND U2618 ( .A(n1748), .B(n1749), .Z(z2[242]) );
  NANDN U2619 ( .A(xregN_1), .B(zin[241]), .Z(n1749) );
  NAND U2620 ( .A(N246), .B(xregN_1), .Z(n1748) );
  NAND U2621 ( .A(n1750), .B(n1751), .Z(z2[241]) );
  NANDN U2622 ( .A(xregN_1), .B(zin[240]), .Z(n1751) );
  NAND U2623 ( .A(N245), .B(xregN_1), .Z(n1750) );
  NAND U2624 ( .A(n1752), .B(n1753), .Z(z2[240]) );
  NANDN U2625 ( .A(xregN_1), .B(zin[239]), .Z(n1753) );
  NAND U2626 ( .A(N244), .B(xregN_1), .Z(n1752) );
  NAND U2627 ( .A(n1754), .B(n1755), .Z(z2[23]) );
  NANDN U2628 ( .A(xregN_1), .B(zin[22]), .Z(n1755) );
  NAND U2629 ( .A(N27), .B(xregN_1), .Z(n1754) );
  NAND U2630 ( .A(n1756), .B(n1757), .Z(z2[239]) );
  NANDN U2631 ( .A(xregN_1), .B(zin[238]), .Z(n1757) );
  NAND U2632 ( .A(N243), .B(xregN_1), .Z(n1756) );
  NAND U2633 ( .A(n1758), .B(n1759), .Z(z2[238]) );
  NANDN U2634 ( .A(xregN_1), .B(zin[237]), .Z(n1759) );
  NAND U2635 ( .A(N242), .B(xregN_1), .Z(n1758) );
  NAND U2636 ( .A(n1760), .B(n1761), .Z(z2[237]) );
  NANDN U2637 ( .A(xregN_1), .B(zin[236]), .Z(n1761) );
  NAND U2638 ( .A(N241), .B(xregN_1), .Z(n1760) );
  NAND U2639 ( .A(n1762), .B(n1763), .Z(z2[236]) );
  NANDN U2640 ( .A(xregN_1), .B(zin[235]), .Z(n1763) );
  NAND U2641 ( .A(N240), .B(xregN_1), .Z(n1762) );
  NAND U2642 ( .A(n1764), .B(n1765), .Z(z2[235]) );
  NANDN U2643 ( .A(xregN_1), .B(zin[234]), .Z(n1765) );
  NAND U2644 ( .A(N239), .B(xregN_1), .Z(n1764) );
  NAND U2645 ( .A(n1766), .B(n1767), .Z(z2[234]) );
  NANDN U2646 ( .A(xregN_1), .B(zin[233]), .Z(n1767) );
  NAND U2647 ( .A(N238), .B(xregN_1), .Z(n1766) );
  NAND U2648 ( .A(n1768), .B(n1769), .Z(z2[233]) );
  NANDN U2649 ( .A(xregN_1), .B(zin[232]), .Z(n1769) );
  NAND U2650 ( .A(N237), .B(xregN_1), .Z(n1768) );
  NAND U2651 ( .A(n1770), .B(n1771), .Z(z2[232]) );
  NANDN U2652 ( .A(xregN_1), .B(zin[231]), .Z(n1771) );
  NAND U2653 ( .A(N236), .B(xregN_1), .Z(n1770) );
  NAND U2654 ( .A(n1772), .B(n1773), .Z(z2[231]) );
  NANDN U2655 ( .A(xregN_1), .B(zin[230]), .Z(n1773) );
  NAND U2656 ( .A(N235), .B(xregN_1), .Z(n1772) );
  NAND U2657 ( .A(n1774), .B(n1775), .Z(z2[230]) );
  NANDN U2658 ( .A(xregN_1), .B(zin[229]), .Z(n1775) );
  NAND U2659 ( .A(N234), .B(xregN_1), .Z(n1774) );
  NAND U2660 ( .A(n1776), .B(n1777), .Z(z2[22]) );
  NANDN U2661 ( .A(xregN_1), .B(zin[21]), .Z(n1777) );
  NAND U2662 ( .A(N26), .B(xregN_1), .Z(n1776) );
  NAND U2663 ( .A(n1778), .B(n1779), .Z(z2[229]) );
  NANDN U2664 ( .A(xregN_1), .B(zin[228]), .Z(n1779) );
  NAND U2665 ( .A(N233), .B(xregN_1), .Z(n1778) );
  NAND U2666 ( .A(n1780), .B(n1781), .Z(z2[228]) );
  NANDN U2667 ( .A(xregN_1), .B(zin[227]), .Z(n1781) );
  NAND U2668 ( .A(N232), .B(xregN_1), .Z(n1780) );
  NAND U2669 ( .A(n1782), .B(n1783), .Z(z2[227]) );
  NANDN U2670 ( .A(xregN_1), .B(zin[226]), .Z(n1783) );
  NAND U2671 ( .A(N231), .B(xregN_1), .Z(n1782) );
  NAND U2672 ( .A(n1784), .B(n1785), .Z(z2[226]) );
  NANDN U2673 ( .A(xregN_1), .B(zin[225]), .Z(n1785) );
  NAND U2674 ( .A(N230), .B(xregN_1), .Z(n1784) );
  NAND U2675 ( .A(n1786), .B(n1787), .Z(z2[225]) );
  NANDN U2676 ( .A(xregN_1), .B(zin[224]), .Z(n1787) );
  NAND U2677 ( .A(N229), .B(xregN_1), .Z(n1786) );
  NAND U2678 ( .A(n1788), .B(n1789), .Z(z2[224]) );
  NANDN U2679 ( .A(xregN_1), .B(zin[223]), .Z(n1789) );
  NAND U2680 ( .A(N228), .B(xregN_1), .Z(n1788) );
  NAND U2681 ( .A(n1790), .B(n1791), .Z(z2[223]) );
  NANDN U2682 ( .A(xregN_1), .B(zin[222]), .Z(n1791) );
  NAND U2683 ( .A(N227), .B(xregN_1), .Z(n1790) );
  NAND U2684 ( .A(n1792), .B(n1793), .Z(z2[222]) );
  NANDN U2685 ( .A(xregN_1), .B(zin[221]), .Z(n1793) );
  NAND U2686 ( .A(N226), .B(xregN_1), .Z(n1792) );
  NAND U2687 ( .A(n1794), .B(n1795), .Z(z2[221]) );
  NANDN U2688 ( .A(xregN_1), .B(zin[220]), .Z(n1795) );
  NAND U2689 ( .A(N225), .B(xregN_1), .Z(n1794) );
  NAND U2690 ( .A(n1796), .B(n1797), .Z(z2[220]) );
  NANDN U2691 ( .A(xregN_1), .B(zin[219]), .Z(n1797) );
  NAND U2692 ( .A(N224), .B(xregN_1), .Z(n1796) );
  NAND U2693 ( .A(n1798), .B(n1799), .Z(z2[21]) );
  NANDN U2694 ( .A(xregN_1), .B(zin[20]), .Z(n1799) );
  NAND U2695 ( .A(N25), .B(xregN_1), .Z(n1798) );
  NAND U2696 ( .A(n1800), .B(n1801), .Z(z2[219]) );
  NANDN U2697 ( .A(xregN_1), .B(zin[218]), .Z(n1801) );
  NAND U2698 ( .A(N223), .B(xregN_1), .Z(n1800) );
  NAND U2699 ( .A(n1802), .B(n1803), .Z(z2[218]) );
  NANDN U2700 ( .A(xregN_1), .B(zin[217]), .Z(n1803) );
  NAND U2701 ( .A(N222), .B(xregN_1), .Z(n1802) );
  NAND U2702 ( .A(n1804), .B(n1805), .Z(z2[217]) );
  NANDN U2703 ( .A(xregN_1), .B(zin[216]), .Z(n1805) );
  NAND U2704 ( .A(N221), .B(xregN_1), .Z(n1804) );
  NAND U2705 ( .A(n1806), .B(n1807), .Z(z2[216]) );
  NANDN U2706 ( .A(xregN_1), .B(zin[215]), .Z(n1807) );
  NAND U2707 ( .A(N220), .B(xregN_1), .Z(n1806) );
  NAND U2708 ( .A(n1808), .B(n1809), .Z(z2[215]) );
  NANDN U2709 ( .A(xregN_1), .B(zin[214]), .Z(n1809) );
  NAND U2710 ( .A(N219), .B(xregN_1), .Z(n1808) );
  NAND U2711 ( .A(n1810), .B(n1811), .Z(z2[214]) );
  NANDN U2712 ( .A(xregN_1), .B(zin[213]), .Z(n1811) );
  NAND U2713 ( .A(N218), .B(xregN_1), .Z(n1810) );
  NAND U2714 ( .A(n1812), .B(n1813), .Z(z2[213]) );
  NANDN U2715 ( .A(xregN_1), .B(zin[212]), .Z(n1813) );
  NAND U2716 ( .A(N217), .B(xregN_1), .Z(n1812) );
  NAND U2717 ( .A(n1814), .B(n1815), .Z(z2[212]) );
  NANDN U2718 ( .A(xregN_1), .B(zin[211]), .Z(n1815) );
  NAND U2719 ( .A(N216), .B(xregN_1), .Z(n1814) );
  NAND U2720 ( .A(n1816), .B(n1817), .Z(z2[211]) );
  NANDN U2721 ( .A(xregN_1), .B(zin[210]), .Z(n1817) );
  NAND U2722 ( .A(N215), .B(xregN_1), .Z(n1816) );
  NAND U2723 ( .A(n1818), .B(n1819), .Z(z2[210]) );
  NANDN U2724 ( .A(xregN_1), .B(zin[209]), .Z(n1819) );
  NAND U2725 ( .A(N214), .B(xregN_1), .Z(n1818) );
  NAND U2726 ( .A(n1820), .B(n1821), .Z(z2[20]) );
  NANDN U2727 ( .A(xregN_1), .B(zin[19]), .Z(n1821) );
  NAND U2728 ( .A(N24), .B(xregN_1), .Z(n1820) );
  NAND U2729 ( .A(n1822), .B(n1823), .Z(z2[209]) );
  NANDN U2730 ( .A(xregN_1), .B(zin[208]), .Z(n1823) );
  NAND U2731 ( .A(N213), .B(xregN_1), .Z(n1822) );
  NAND U2732 ( .A(n1824), .B(n1825), .Z(z2[208]) );
  NANDN U2733 ( .A(xregN_1), .B(zin[207]), .Z(n1825) );
  NAND U2734 ( .A(N212), .B(xregN_1), .Z(n1824) );
  NAND U2735 ( .A(n1826), .B(n1827), .Z(z2[207]) );
  NANDN U2736 ( .A(xregN_1), .B(zin[206]), .Z(n1827) );
  NAND U2737 ( .A(N211), .B(xregN_1), .Z(n1826) );
  NAND U2738 ( .A(n1828), .B(n1829), .Z(z2[206]) );
  NANDN U2739 ( .A(xregN_1), .B(zin[205]), .Z(n1829) );
  NAND U2740 ( .A(N210), .B(xregN_1), .Z(n1828) );
  NAND U2741 ( .A(n1830), .B(n1831), .Z(z2[205]) );
  NANDN U2742 ( .A(xregN_1), .B(zin[204]), .Z(n1831) );
  NAND U2743 ( .A(N209), .B(xregN_1), .Z(n1830) );
  NAND U2744 ( .A(n1832), .B(n1833), .Z(z2[204]) );
  NANDN U2745 ( .A(xregN_1), .B(zin[203]), .Z(n1833) );
  NAND U2746 ( .A(N208), .B(xregN_1), .Z(n1832) );
  NAND U2747 ( .A(n1834), .B(n1835), .Z(z2[203]) );
  NANDN U2748 ( .A(xregN_1), .B(zin[202]), .Z(n1835) );
  NAND U2749 ( .A(N207), .B(xregN_1), .Z(n1834) );
  NAND U2750 ( .A(n1836), .B(n1837), .Z(z2[202]) );
  NANDN U2751 ( .A(xregN_1), .B(zin[201]), .Z(n1837) );
  NAND U2752 ( .A(N206), .B(xregN_1), .Z(n1836) );
  NAND U2753 ( .A(n1838), .B(n1839), .Z(z2[201]) );
  NANDN U2754 ( .A(xregN_1), .B(zin[200]), .Z(n1839) );
  NAND U2755 ( .A(N205), .B(xregN_1), .Z(n1838) );
  NAND U2756 ( .A(n1840), .B(n1841), .Z(z2[200]) );
  NANDN U2757 ( .A(xregN_1), .B(zin[199]), .Z(n1841) );
  NAND U2758 ( .A(N204), .B(xregN_1), .Z(n1840) );
  NAND U2759 ( .A(n1842), .B(n1843), .Z(z2[1]) );
  NANDN U2760 ( .A(xregN_1), .B(zin[0]), .Z(n1843) );
  NAND U2761 ( .A(N5), .B(xregN_1), .Z(n1842) );
  NAND U2762 ( .A(n1844), .B(n1845), .Z(z2[19]) );
  NANDN U2763 ( .A(xregN_1), .B(zin[18]), .Z(n1845) );
  NAND U2764 ( .A(N23), .B(xregN_1), .Z(n1844) );
  NAND U2765 ( .A(n1846), .B(n1847), .Z(z2[199]) );
  NANDN U2766 ( .A(xregN_1), .B(zin[198]), .Z(n1847) );
  NAND U2767 ( .A(N203), .B(xregN_1), .Z(n1846) );
  NAND U2768 ( .A(n1848), .B(n1849), .Z(z2[198]) );
  NANDN U2769 ( .A(xregN_1), .B(zin[197]), .Z(n1849) );
  NAND U2770 ( .A(N202), .B(xregN_1), .Z(n1848) );
  NAND U2771 ( .A(n1850), .B(n1851), .Z(z2[197]) );
  NANDN U2772 ( .A(xregN_1), .B(zin[196]), .Z(n1851) );
  NAND U2773 ( .A(N201), .B(xregN_1), .Z(n1850) );
  NAND U2774 ( .A(n1852), .B(n1853), .Z(z2[196]) );
  NANDN U2775 ( .A(xregN_1), .B(zin[195]), .Z(n1853) );
  NAND U2776 ( .A(N200), .B(xregN_1), .Z(n1852) );
  NAND U2777 ( .A(n1854), .B(n1855), .Z(z2[195]) );
  NANDN U2778 ( .A(xregN_1), .B(zin[194]), .Z(n1855) );
  NAND U2779 ( .A(N199), .B(xregN_1), .Z(n1854) );
  NAND U2780 ( .A(n1856), .B(n1857), .Z(z2[194]) );
  NANDN U2781 ( .A(xregN_1), .B(zin[193]), .Z(n1857) );
  NAND U2782 ( .A(N198), .B(xregN_1), .Z(n1856) );
  NAND U2783 ( .A(n1858), .B(n1859), .Z(z2[193]) );
  NANDN U2784 ( .A(xregN_1), .B(zin[192]), .Z(n1859) );
  NAND U2785 ( .A(N197), .B(xregN_1), .Z(n1858) );
  NAND U2786 ( .A(n1860), .B(n1861), .Z(z2[192]) );
  NANDN U2787 ( .A(xregN_1), .B(zin[191]), .Z(n1861) );
  NAND U2788 ( .A(N196), .B(xregN_1), .Z(n1860) );
  NAND U2789 ( .A(n1862), .B(n1863), .Z(z2[191]) );
  NANDN U2790 ( .A(xregN_1), .B(zin[190]), .Z(n1863) );
  NAND U2791 ( .A(N195), .B(xregN_1), .Z(n1862) );
  NAND U2792 ( .A(n1864), .B(n1865), .Z(z2[190]) );
  NANDN U2793 ( .A(xregN_1), .B(zin[189]), .Z(n1865) );
  NAND U2794 ( .A(N194), .B(xregN_1), .Z(n1864) );
  NAND U2795 ( .A(n1866), .B(n1867), .Z(z2[18]) );
  NANDN U2796 ( .A(xregN_1), .B(zin[17]), .Z(n1867) );
  NAND U2797 ( .A(N22), .B(xregN_1), .Z(n1866) );
  NAND U2798 ( .A(n1868), .B(n1869), .Z(z2[189]) );
  NANDN U2799 ( .A(xregN_1), .B(zin[188]), .Z(n1869) );
  NAND U2800 ( .A(N193), .B(xregN_1), .Z(n1868) );
  NAND U2801 ( .A(n1870), .B(n1871), .Z(z2[188]) );
  NANDN U2802 ( .A(xregN_1), .B(zin[187]), .Z(n1871) );
  NAND U2803 ( .A(N192), .B(xregN_1), .Z(n1870) );
  NAND U2804 ( .A(n1872), .B(n1873), .Z(z2[187]) );
  NANDN U2805 ( .A(xregN_1), .B(zin[186]), .Z(n1873) );
  NAND U2806 ( .A(N191), .B(xregN_1), .Z(n1872) );
  NAND U2807 ( .A(n1874), .B(n1875), .Z(z2[186]) );
  NANDN U2808 ( .A(xregN_1), .B(zin[185]), .Z(n1875) );
  NAND U2809 ( .A(N190), .B(xregN_1), .Z(n1874) );
  NAND U2810 ( .A(n1876), .B(n1877), .Z(z2[185]) );
  NANDN U2811 ( .A(xregN_1), .B(zin[184]), .Z(n1877) );
  NAND U2812 ( .A(N189), .B(xregN_1), .Z(n1876) );
  NAND U2813 ( .A(n1878), .B(n1879), .Z(z2[184]) );
  NANDN U2814 ( .A(xregN_1), .B(zin[183]), .Z(n1879) );
  NAND U2815 ( .A(N188), .B(xregN_1), .Z(n1878) );
  NAND U2816 ( .A(n1880), .B(n1881), .Z(z2[183]) );
  NANDN U2817 ( .A(xregN_1), .B(zin[182]), .Z(n1881) );
  NAND U2818 ( .A(N187), .B(xregN_1), .Z(n1880) );
  NAND U2819 ( .A(n1882), .B(n1883), .Z(z2[182]) );
  NANDN U2820 ( .A(xregN_1), .B(zin[181]), .Z(n1883) );
  NAND U2821 ( .A(N186), .B(xregN_1), .Z(n1882) );
  NAND U2822 ( .A(n1884), .B(n1885), .Z(z2[181]) );
  NANDN U2823 ( .A(xregN_1), .B(zin[180]), .Z(n1885) );
  NAND U2824 ( .A(N185), .B(xregN_1), .Z(n1884) );
  NAND U2825 ( .A(n1886), .B(n1887), .Z(z2[180]) );
  NANDN U2826 ( .A(xregN_1), .B(zin[179]), .Z(n1887) );
  NAND U2827 ( .A(N184), .B(xregN_1), .Z(n1886) );
  NAND U2828 ( .A(n1888), .B(n1889), .Z(z2[17]) );
  NANDN U2829 ( .A(xregN_1), .B(zin[16]), .Z(n1889) );
  NAND U2830 ( .A(N21), .B(xregN_1), .Z(n1888) );
  NAND U2831 ( .A(n1890), .B(n1891), .Z(z2[179]) );
  NANDN U2832 ( .A(xregN_1), .B(zin[178]), .Z(n1891) );
  NAND U2833 ( .A(N183), .B(xregN_1), .Z(n1890) );
  NAND U2834 ( .A(n1892), .B(n1893), .Z(z2[178]) );
  NANDN U2835 ( .A(xregN_1), .B(zin[177]), .Z(n1893) );
  NAND U2836 ( .A(N182), .B(xregN_1), .Z(n1892) );
  NAND U2837 ( .A(n1894), .B(n1895), .Z(z2[177]) );
  NANDN U2838 ( .A(xregN_1), .B(zin[176]), .Z(n1895) );
  NAND U2839 ( .A(N181), .B(xregN_1), .Z(n1894) );
  NAND U2840 ( .A(n1896), .B(n1897), .Z(z2[176]) );
  NANDN U2841 ( .A(xregN_1), .B(zin[175]), .Z(n1897) );
  NAND U2842 ( .A(N180), .B(xregN_1), .Z(n1896) );
  NAND U2843 ( .A(n1898), .B(n1899), .Z(z2[175]) );
  NANDN U2844 ( .A(xregN_1), .B(zin[174]), .Z(n1899) );
  NAND U2845 ( .A(N179), .B(xregN_1), .Z(n1898) );
  NAND U2846 ( .A(n1900), .B(n1901), .Z(z2[174]) );
  NANDN U2847 ( .A(xregN_1), .B(zin[173]), .Z(n1901) );
  NAND U2848 ( .A(N178), .B(xregN_1), .Z(n1900) );
  NAND U2849 ( .A(n1902), .B(n1903), .Z(z2[173]) );
  NANDN U2850 ( .A(xregN_1), .B(zin[172]), .Z(n1903) );
  NAND U2851 ( .A(N177), .B(xregN_1), .Z(n1902) );
  NAND U2852 ( .A(n1904), .B(n1905), .Z(z2[172]) );
  NANDN U2853 ( .A(xregN_1), .B(zin[171]), .Z(n1905) );
  NAND U2854 ( .A(N176), .B(xregN_1), .Z(n1904) );
  NAND U2855 ( .A(n1906), .B(n1907), .Z(z2[171]) );
  NANDN U2856 ( .A(xregN_1), .B(zin[170]), .Z(n1907) );
  NAND U2857 ( .A(N175), .B(xregN_1), .Z(n1906) );
  NAND U2858 ( .A(n1908), .B(n1909), .Z(z2[170]) );
  NANDN U2859 ( .A(xregN_1), .B(zin[169]), .Z(n1909) );
  NAND U2860 ( .A(N174), .B(xregN_1), .Z(n1908) );
  NAND U2861 ( .A(n1910), .B(n1911), .Z(z2[16]) );
  NANDN U2862 ( .A(xregN_1), .B(zin[15]), .Z(n1911) );
  NAND U2863 ( .A(N20), .B(xregN_1), .Z(n1910) );
  NAND U2864 ( .A(n1912), .B(n1913), .Z(z2[169]) );
  NANDN U2865 ( .A(xregN_1), .B(zin[168]), .Z(n1913) );
  NAND U2866 ( .A(N173), .B(xregN_1), .Z(n1912) );
  NAND U2867 ( .A(n1914), .B(n1915), .Z(z2[168]) );
  NANDN U2868 ( .A(xregN_1), .B(zin[167]), .Z(n1915) );
  NAND U2869 ( .A(N172), .B(xregN_1), .Z(n1914) );
  NAND U2870 ( .A(n1916), .B(n1917), .Z(z2[167]) );
  NANDN U2871 ( .A(xregN_1), .B(zin[166]), .Z(n1917) );
  NAND U2872 ( .A(N171), .B(xregN_1), .Z(n1916) );
  NAND U2873 ( .A(n1918), .B(n1919), .Z(z2[166]) );
  NANDN U2874 ( .A(xregN_1), .B(zin[165]), .Z(n1919) );
  NAND U2875 ( .A(N170), .B(xregN_1), .Z(n1918) );
  NAND U2876 ( .A(n1920), .B(n1921), .Z(z2[165]) );
  NANDN U2877 ( .A(xregN_1), .B(zin[164]), .Z(n1921) );
  NAND U2878 ( .A(N169), .B(xregN_1), .Z(n1920) );
  NAND U2879 ( .A(n1922), .B(n1923), .Z(z2[164]) );
  NANDN U2880 ( .A(xregN_1), .B(zin[163]), .Z(n1923) );
  NAND U2881 ( .A(N168), .B(xregN_1), .Z(n1922) );
  NAND U2882 ( .A(n1924), .B(n1925), .Z(z2[163]) );
  NANDN U2883 ( .A(xregN_1), .B(zin[162]), .Z(n1925) );
  NAND U2884 ( .A(N167), .B(xregN_1), .Z(n1924) );
  NAND U2885 ( .A(n1926), .B(n1927), .Z(z2[162]) );
  NANDN U2886 ( .A(xregN_1), .B(zin[161]), .Z(n1927) );
  NAND U2887 ( .A(N166), .B(xregN_1), .Z(n1926) );
  NAND U2888 ( .A(n1928), .B(n1929), .Z(z2[161]) );
  NANDN U2889 ( .A(xregN_1), .B(zin[160]), .Z(n1929) );
  NAND U2890 ( .A(N165), .B(xregN_1), .Z(n1928) );
  NAND U2891 ( .A(n1930), .B(n1931), .Z(z2[160]) );
  NANDN U2892 ( .A(xregN_1), .B(zin[159]), .Z(n1931) );
  NAND U2893 ( .A(N164), .B(xregN_1), .Z(n1930) );
  NAND U2894 ( .A(n1932), .B(n1933), .Z(z2[15]) );
  NANDN U2895 ( .A(xregN_1), .B(zin[14]), .Z(n1933) );
  NAND U2896 ( .A(N19), .B(xregN_1), .Z(n1932) );
  NAND U2897 ( .A(n1934), .B(n1935), .Z(z2[159]) );
  NANDN U2898 ( .A(xregN_1), .B(zin[158]), .Z(n1935) );
  NAND U2899 ( .A(N163), .B(xregN_1), .Z(n1934) );
  NAND U2900 ( .A(n1936), .B(n1937), .Z(z2[158]) );
  NANDN U2901 ( .A(xregN_1), .B(zin[157]), .Z(n1937) );
  NAND U2902 ( .A(N162), .B(xregN_1), .Z(n1936) );
  NAND U2903 ( .A(n1938), .B(n1939), .Z(z2[157]) );
  NANDN U2904 ( .A(xregN_1), .B(zin[156]), .Z(n1939) );
  NAND U2905 ( .A(N161), .B(xregN_1), .Z(n1938) );
  NAND U2906 ( .A(n1940), .B(n1941), .Z(z2[156]) );
  NANDN U2907 ( .A(xregN_1), .B(zin[155]), .Z(n1941) );
  NAND U2908 ( .A(N160), .B(xregN_1), .Z(n1940) );
  NAND U2909 ( .A(n1942), .B(n1943), .Z(z2[155]) );
  NANDN U2910 ( .A(xregN_1), .B(zin[154]), .Z(n1943) );
  NAND U2911 ( .A(N159), .B(xregN_1), .Z(n1942) );
  NAND U2912 ( .A(n1944), .B(n1945), .Z(z2[154]) );
  NANDN U2913 ( .A(xregN_1), .B(zin[153]), .Z(n1945) );
  NAND U2914 ( .A(N158), .B(xregN_1), .Z(n1944) );
  NAND U2915 ( .A(n1946), .B(n1947), .Z(z2[153]) );
  NANDN U2916 ( .A(xregN_1), .B(zin[152]), .Z(n1947) );
  NAND U2917 ( .A(N157), .B(xregN_1), .Z(n1946) );
  NAND U2918 ( .A(n1948), .B(n1949), .Z(z2[152]) );
  NANDN U2919 ( .A(xregN_1), .B(zin[151]), .Z(n1949) );
  NAND U2920 ( .A(N156), .B(xregN_1), .Z(n1948) );
  NAND U2921 ( .A(n1950), .B(n1951), .Z(z2[151]) );
  NANDN U2922 ( .A(xregN_1), .B(zin[150]), .Z(n1951) );
  NAND U2923 ( .A(N155), .B(xregN_1), .Z(n1950) );
  NAND U2924 ( .A(n1952), .B(n1953), .Z(z2[150]) );
  NANDN U2925 ( .A(xregN_1), .B(zin[149]), .Z(n1953) );
  NAND U2926 ( .A(N154), .B(xregN_1), .Z(n1952) );
  NAND U2927 ( .A(n1954), .B(n1955), .Z(z2[14]) );
  NANDN U2928 ( .A(xregN_1), .B(zin[13]), .Z(n1955) );
  NAND U2929 ( .A(N18), .B(xregN_1), .Z(n1954) );
  NAND U2930 ( .A(n1956), .B(n1957), .Z(z2[149]) );
  NANDN U2931 ( .A(xregN_1), .B(zin[148]), .Z(n1957) );
  NAND U2932 ( .A(N153), .B(xregN_1), .Z(n1956) );
  NAND U2933 ( .A(n1958), .B(n1959), .Z(z2[148]) );
  NANDN U2934 ( .A(xregN_1), .B(zin[147]), .Z(n1959) );
  NAND U2935 ( .A(N152), .B(xregN_1), .Z(n1958) );
  NAND U2936 ( .A(n1960), .B(n1961), .Z(z2[147]) );
  NANDN U2937 ( .A(xregN_1), .B(zin[146]), .Z(n1961) );
  NAND U2938 ( .A(N151), .B(xregN_1), .Z(n1960) );
  NAND U2939 ( .A(n1962), .B(n1963), .Z(z2[146]) );
  NANDN U2940 ( .A(xregN_1), .B(zin[145]), .Z(n1963) );
  NAND U2941 ( .A(N150), .B(xregN_1), .Z(n1962) );
  NAND U2942 ( .A(n1964), .B(n1965), .Z(z2[145]) );
  NANDN U2943 ( .A(xregN_1), .B(zin[144]), .Z(n1965) );
  NAND U2944 ( .A(N149), .B(xregN_1), .Z(n1964) );
  NAND U2945 ( .A(n1966), .B(n1967), .Z(z2[144]) );
  NANDN U2946 ( .A(xregN_1), .B(zin[143]), .Z(n1967) );
  NAND U2947 ( .A(N148), .B(xregN_1), .Z(n1966) );
  NAND U2948 ( .A(n1968), .B(n1969), .Z(z2[143]) );
  NANDN U2949 ( .A(xregN_1), .B(zin[142]), .Z(n1969) );
  NAND U2950 ( .A(N147), .B(xregN_1), .Z(n1968) );
  NAND U2951 ( .A(n1970), .B(n1971), .Z(z2[142]) );
  NANDN U2952 ( .A(xregN_1), .B(zin[141]), .Z(n1971) );
  NAND U2953 ( .A(N146), .B(xregN_1), .Z(n1970) );
  NAND U2954 ( .A(n1972), .B(n1973), .Z(z2[141]) );
  NANDN U2955 ( .A(xregN_1), .B(zin[140]), .Z(n1973) );
  NAND U2956 ( .A(N145), .B(xregN_1), .Z(n1972) );
  NAND U2957 ( .A(n1974), .B(n1975), .Z(z2[140]) );
  NANDN U2958 ( .A(xregN_1), .B(zin[139]), .Z(n1975) );
  NAND U2959 ( .A(N144), .B(xregN_1), .Z(n1974) );
  NAND U2960 ( .A(n1976), .B(n1977), .Z(z2[13]) );
  NANDN U2961 ( .A(xregN_1), .B(zin[12]), .Z(n1977) );
  NAND U2962 ( .A(N17), .B(xregN_1), .Z(n1976) );
  NAND U2963 ( .A(n1978), .B(n1979), .Z(z2[139]) );
  NANDN U2964 ( .A(xregN_1), .B(zin[138]), .Z(n1979) );
  NAND U2965 ( .A(N143), .B(xregN_1), .Z(n1978) );
  NAND U2966 ( .A(n1980), .B(n1981), .Z(z2[138]) );
  NANDN U2967 ( .A(xregN_1), .B(zin[137]), .Z(n1981) );
  NAND U2968 ( .A(N142), .B(xregN_1), .Z(n1980) );
  NAND U2969 ( .A(n1982), .B(n1983), .Z(z2[137]) );
  NANDN U2970 ( .A(xregN_1), .B(zin[136]), .Z(n1983) );
  NAND U2971 ( .A(N141), .B(xregN_1), .Z(n1982) );
  NAND U2972 ( .A(n1984), .B(n1985), .Z(z2[136]) );
  NANDN U2973 ( .A(xregN_1), .B(zin[135]), .Z(n1985) );
  NAND U2974 ( .A(N140), .B(xregN_1), .Z(n1984) );
  NAND U2975 ( .A(n1986), .B(n1987), .Z(z2[135]) );
  NANDN U2976 ( .A(xregN_1), .B(zin[134]), .Z(n1987) );
  NAND U2977 ( .A(N139), .B(xregN_1), .Z(n1986) );
  NAND U2978 ( .A(n1988), .B(n1989), .Z(z2[134]) );
  NANDN U2979 ( .A(xregN_1), .B(zin[133]), .Z(n1989) );
  NAND U2980 ( .A(N138), .B(xregN_1), .Z(n1988) );
  NAND U2981 ( .A(n1990), .B(n1991), .Z(z2[133]) );
  NANDN U2982 ( .A(xregN_1), .B(zin[132]), .Z(n1991) );
  NAND U2983 ( .A(N137), .B(xregN_1), .Z(n1990) );
  NAND U2984 ( .A(n1992), .B(n1993), .Z(z2[132]) );
  NANDN U2985 ( .A(xregN_1), .B(zin[131]), .Z(n1993) );
  NAND U2986 ( .A(N136), .B(xregN_1), .Z(n1992) );
  NAND U2987 ( .A(n1994), .B(n1995), .Z(z2[131]) );
  NANDN U2988 ( .A(xregN_1), .B(zin[130]), .Z(n1995) );
  NAND U2989 ( .A(N135), .B(xregN_1), .Z(n1994) );
  NAND U2990 ( .A(n1996), .B(n1997), .Z(z2[130]) );
  NANDN U2991 ( .A(xregN_1), .B(zin[129]), .Z(n1997) );
  NAND U2992 ( .A(N134), .B(xregN_1), .Z(n1996) );
  NAND U2993 ( .A(n1998), .B(n1999), .Z(z2[12]) );
  NANDN U2994 ( .A(xregN_1), .B(zin[11]), .Z(n1999) );
  NAND U2995 ( .A(N16), .B(xregN_1), .Z(n1998) );
  NAND U2996 ( .A(n2000), .B(n2001), .Z(z2[129]) );
  NANDN U2997 ( .A(xregN_1), .B(zin[128]), .Z(n2001) );
  NAND U2998 ( .A(N133), .B(xregN_1), .Z(n2000) );
  NAND U2999 ( .A(n2002), .B(n2003), .Z(z2[128]) );
  NANDN U3000 ( .A(xregN_1), .B(zin[127]), .Z(n2003) );
  NAND U3001 ( .A(N132), .B(xregN_1), .Z(n2002) );
  NAND U3002 ( .A(n2004), .B(n2005), .Z(z2[127]) );
  NANDN U3003 ( .A(xregN_1), .B(zin[126]), .Z(n2005) );
  NAND U3004 ( .A(N131), .B(xregN_1), .Z(n2004) );
  NAND U3005 ( .A(n2006), .B(n2007), .Z(z2[126]) );
  NANDN U3006 ( .A(xregN_1), .B(zin[125]), .Z(n2007) );
  NAND U3007 ( .A(N130), .B(xregN_1), .Z(n2006) );
  NAND U3008 ( .A(n2008), .B(n2009), .Z(z2[125]) );
  NANDN U3009 ( .A(xregN_1), .B(zin[124]), .Z(n2009) );
  NAND U3010 ( .A(N129), .B(xregN_1), .Z(n2008) );
  NAND U3011 ( .A(n2010), .B(n2011), .Z(z2[124]) );
  NANDN U3012 ( .A(xregN_1), .B(zin[123]), .Z(n2011) );
  NAND U3013 ( .A(N128), .B(xregN_1), .Z(n2010) );
  NAND U3014 ( .A(n2012), .B(n2013), .Z(z2[123]) );
  NANDN U3015 ( .A(xregN_1), .B(zin[122]), .Z(n2013) );
  NAND U3016 ( .A(N127), .B(xregN_1), .Z(n2012) );
  NAND U3017 ( .A(n2014), .B(n2015), .Z(z2[122]) );
  NANDN U3018 ( .A(xregN_1), .B(zin[121]), .Z(n2015) );
  NAND U3019 ( .A(N126), .B(xregN_1), .Z(n2014) );
  NAND U3020 ( .A(n2016), .B(n2017), .Z(z2[121]) );
  NANDN U3021 ( .A(xregN_1), .B(zin[120]), .Z(n2017) );
  NAND U3022 ( .A(N125), .B(xregN_1), .Z(n2016) );
  NAND U3023 ( .A(n2018), .B(n2019), .Z(z2[120]) );
  NANDN U3024 ( .A(xregN_1), .B(zin[119]), .Z(n2019) );
  NAND U3025 ( .A(N124), .B(xregN_1), .Z(n2018) );
  NAND U3026 ( .A(n2020), .B(n2021), .Z(z2[11]) );
  NANDN U3027 ( .A(xregN_1), .B(zin[10]), .Z(n2021) );
  NAND U3028 ( .A(N15), .B(xregN_1), .Z(n2020) );
  NAND U3029 ( .A(n2022), .B(n2023), .Z(z2[119]) );
  NANDN U3030 ( .A(xregN_1), .B(zin[118]), .Z(n2023) );
  NAND U3031 ( .A(N123), .B(xregN_1), .Z(n2022) );
  NAND U3032 ( .A(n2024), .B(n2025), .Z(z2[118]) );
  NANDN U3033 ( .A(xregN_1), .B(zin[117]), .Z(n2025) );
  NAND U3034 ( .A(N122), .B(xregN_1), .Z(n2024) );
  NAND U3035 ( .A(n2026), .B(n2027), .Z(z2[117]) );
  NANDN U3036 ( .A(xregN_1), .B(zin[116]), .Z(n2027) );
  NAND U3037 ( .A(N121), .B(xregN_1), .Z(n2026) );
  NAND U3038 ( .A(n2028), .B(n2029), .Z(z2[116]) );
  NANDN U3039 ( .A(xregN_1), .B(zin[115]), .Z(n2029) );
  NAND U3040 ( .A(N120), .B(xregN_1), .Z(n2028) );
  NAND U3041 ( .A(n2030), .B(n2031), .Z(z2[115]) );
  NANDN U3042 ( .A(xregN_1), .B(zin[114]), .Z(n2031) );
  NAND U3043 ( .A(N119), .B(xregN_1), .Z(n2030) );
  NAND U3044 ( .A(n2032), .B(n2033), .Z(z2[114]) );
  NANDN U3045 ( .A(xregN_1), .B(zin[113]), .Z(n2033) );
  NAND U3046 ( .A(N118), .B(xregN_1), .Z(n2032) );
  NAND U3047 ( .A(n2034), .B(n2035), .Z(z2[113]) );
  NANDN U3048 ( .A(xregN_1), .B(zin[112]), .Z(n2035) );
  NAND U3049 ( .A(N117), .B(xregN_1), .Z(n2034) );
  NAND U3050 ( .A(n2036), .B(n2037), .Z(z2[112]) );
  NANDN U3051 ( .A(xregN_1), .B(zin[111]), .Z(n2037) );
  NAND U3052 ( .A(N116), .B(xregN_1), .Z(n2036) );
  NAND U3053 ( .A(n2038), .B(n2039), .Z(z2[111]) );
  NANDN U3054 ( .A(xregN_1), .B(zin[110]), .Z(n2039) );
  NAND U3055 ( .A(N115), .B(xregN_1), .Z(n2038) );
  NAND U3056 ( .A(n2040), .B(n2041), .Z(z2[110]) );
  NANDN U3057 ( .A(xregN_1), .B(zin[109]), .Z(n2041) );
  NAND U3058 ( .A(N114), .B(xregN_1), .Z(n2040) );
  NAND U3059 ( .A(n2042), .B(n2043), .Z(z2[10]) );
  NANDN U3060 ( .A(xregN_1), .B(zin[9]), .Z(n2043) );
  NAND U3061 ( .A(N14), .B(xregN_1), .Z(n2042) );
  NAND U3062 ( .A(n2044), .B(n2045), .Z(z2[109]) );
  NANDN U3063 ( .A(xregN_1), .B(zin[108]), .Z(n2045) );
  NAND U3064 ( .A(N113), .B(xregN_1), .Z(n2044) );
  NAND U3065 ( .A(n2046), .B(n2047), .Z(z2[108]) );
  NANDN U3066 ( .A(xregN_1), .B(zin[107]), .Z(n2047) );
  NAND U3067 ( .A(N112), .B(xregN_1), .Z(n2046) );
  NAND U3068 ( .A(n2048), .B(n2049), .Z(z2[107]) );
  NANDN U3069 ( .A(xregN_1), .B(zin[106]), .Z(n2049) );
  NAND U3070 ( .A(N111), .B(xregN_1), .Z(n2048) );
  NAND U3071 ( .A(n2050), .B(n2051), .Z(z2[106]) );
  NANDN U3072 ( .A(xregN_1), .B(zin[105]), .Z(n2051) );
  NAND U3073 ( .A(N110), .B(xregN_1), .Z(n2050) );
  NAND U3074 ( .A(n2052), .B(n2053), .Z(z2[105]) );
  NANDN U3075 ( .A(xregN_1), .B(zin[104]), .Z(n2053) );
  NAND U3076 ( .A(N109), .B(xregN_1), .Z(n2052) );
  NAND U3077 ( .A(n2054), .B(n2055), .Z(z2[104]) );
  NANDN U3078 ( .A(xregN_1), .B(zin[103]), .Z(n2055) );
  NAND U3079 ( .A(N108), .B(xregN_1), .Z(n2054) );
  NAND U3080 ( .A(n2056), .B(n2057), .Z(z2[103]) );
  NANDN U3081 ( .A(xregN_1), .B(zin[102]), .Z(n2057) );
  NAND U3082 ( .A(N107), .B(xregN_1), .Z(n2056) );
  NAND U3083 ( .A(n2058), .B(n2059), .Z(z2[102]) );
  NANDN U3084 ( .A(xregN_1), .B(zin[101]), .Z(n2059) );
  NAND U3085 ( .A(N106), .B(xregN_1), .Z(n2058) );
  NAND U3086 ( .A(n2060), .B(n2061), .Z(z2[101]) );
  NANDN U3087 ( .A(xregN_1), .B(zin[100]), .Z(n2061) );
  NAND U3088 ( .A(N105), .B(xregN_1), .Z(n2060) );
  NAND U3089 ( .A(n2062), .B(n2063), .Z(z2[100]) );
  NANDN U3090 ( .A(xregN_1), .B(zin[99]), .Z(n2063) );
  NAND U3091 ( .A(N104), .B(xregN_1), .Z(n2062) );
  AND U3092 ( .A(N4), .B(xregN_1), .Z(z2[0]) );
endmodule


module modmult_N512_CC512 ( clk, rst, start, x, y, n, o );
  input [511:0] x;
  input [511:0] y;
  input [511:0] n;
  output [511:0] o;
  input clk, rst, start;
  wire   \zout[0][513] , \zout[0][512] , \zin[0][513] , \zin[0][512] ,
         \zin[0][511] , \zin[0][510] , \zin[0][509] , \zin[0][508] ,
         \zin[0][507] , \zin[0][506] , \zin[0][505] , \zin[0][504] ,
         \zin[0][503] , \zin[0][502] , \zin[0][501] , \zin[0][500] ,
         \zin[0][499] , \zin[0][498] , \zin[0][497] , \zin[0][496] ,
         \zin[0][495] , \zin[0][494] , \zin[0][493] , \zin[0][492] ,
         \zin[0][491] , \zin[0][490] , \zin[0][489] , \zin[0][488] ,
         \zin[0][487] , \zin[0][486] , \zin[0][485] , \zin[0][484] ,
         \zin[0][483] , \zin[0][482] , \zin[0][481] , \zin[0][480] ,
         \zin[0][479] , \zin[0][478] , \zin[0][477] , \zin[0][476] ,
         \zin[0][475] , \zin[0][474] , \zin[0][473] , \zin[0][472] ,
         \zin[0][471] , \zin[0][470] , \zin[0][469] , \zin[0][468] ,
         \zin[0][467] , \zin[0][466] , \zin[0][465] , \zin[0][464] ,
         \zin[0][463] , \zin[0][462] , \zin[0][461] , \zin[0][460] ,
         \zin[0][459] , \zin[0][458] , \zin[0][457] , \zin[0][456] ,
         \zin[0][455] , \zin[0][454] , \zin[0][453] , \zin[0][452] ,
         \zin[0][451] , \zin[0][450] , \zin[0][449] , \zin[0][448] ,
         \zin[0][447] , \zin[0][446] , \zin[0][445] , \zin[0][444] ,
         \zin[0][443] , \zin[0][442] , \zin[0][441] , \zin[0][440] ,
         \zin[0][439] , \zin[0][438] , \zin[0][437] , \zin[0][436] ,
         \zin[0][435] , \zin[0][434] , \zin[0][433] , \zin[0][432] ,
         \zin[0][431] , \zin[0][430] , \zin[0][429] , \zin[0][428] ,
         \zin[0][427] , \zin[0][426] , \zin[0][425] , \zin[0][424] ,
         \zin[0][423] , \zin[0][422] , \zin[0][421] , \zin[0][420] ,
         \zin[0][419] , \zin[0][418] , \zin[0][417] , \zin[0][416] ,
         \zin[0][415] , \zin[0][414] , \zin[0][413] , \zin[0][412] ,
         \zin[0][411] , \zin[0][410] , \zin[0][409] , \zin[0][408] ,
         \zin[0][407] , \zin[0][406] , \zin[0][405] , \zin[0][404] ,
         \zin[0][403] , \zin[0][402] , \zin[0][401] , \zin[0][400] ,
         \zin[0][399] , \zin[0][398] , \zin[0][397] , \zin[0][396] ,
         \zin[0][395] , \zin[0][394] , \zin[0][393] , \zin[0][392] ,
         \zin[0][391] , \zin[0][390] , \zin[0][389] , \zin[0][388] ,
         \zin[0][387] , \zin[0][386] , \zin[0][385] , \zin[0][384] ,
         \zin[0][383] , \zin[0][382] , \zin[0][381] , \zin[0][380] ,
         \zin[0][379] , \zin[0][378] , \zin[0][377] , \zin[0][376] ,
         \zin[0][375] , \zin[0][374] , \zin[0][373] , \zin[0][372] ,
         \zin[0][371] , \zin[0][370] , \zin[0][369] , \zin[0][368] ,
         \zin[0][367] , \zin[0][366] , \zin[0][365] , \zin[0][364] ,
         \zin[0][363] , \zin[0][362] , \zin[0][361] , \zin[0][360] ,
         \zin[0][359] , \zin[0][358] , \zin[0][357] , \zin[0][356] ,
         \zin[0][355] , \zin[0][354] , \zin[0][353] , \zin[0][352] ,
         \zin[0][351] , \zin[0][350] , \zin[0][349] , \zin[0][348] ,
         \zin[0][347] , \zin[0][346] , \zin[0][345] , \zin[0][344] ,
         \zin[0][343] , \zin[0][342] , \zin[0][341] , \zin[0][340] ,
         \zin[0][339] , \zin[0][338] , \zin[0][337] , \zin[0][336] ,
         \zin[0][335] , \zin[0][334] , \zin[0][333] , \zin[0][332] ,
         \zin[0][331] , \zin[0][330] , \zin[0][329] , \zin[0][328] ,
         \zin[0][327] , \zin[0][326] , \zin[0][325] , \zin[0][324] ,
         \zin[0][323] , \zin[0][322] , \zin[0][321] , \zin[0][320] ,
         \zin[0][319] , \zin[0][318] , \zin[0][317] , \zin[0][316] ,
         \zin[0][315] , \zin[0][314] , \zin[0][313] , \zin[0][312] ,
         \zin[0][311] , \zin[0][310] , \zin[0][309] , \zin[0][308] ,
         \zin[0][307] , \zin[0][306] , \zin[0][305] , \zin[0][304] ,
         \zin[0][303] , \zin[0][302] , \zin[0][301] , \zin[0][300] ,
         \zin[0][299] , \zin[0][298] , \zin[0][297] , \zin[0][296] ,
         \zin[0][295] , \zin[0][294] , \zin[0][293] , \zin[0][292] ,
         \zin[0][291] , \zin[0][290] , \zin[0][289] , \zin[0][288] ,
         \zin[0][287] , \zin[0][286] , \zin[0][285] , \zin[0][284] ,
         \zin[0][283] , \zin[0][282] , \zin[0][281] , \zin[0][280] ,
         \zin[0][279] , \zin[0][278] , \zin[0][277] , \zin[0][276] ,
         \zin[0][275] , \zin[0][274] , \zin[0][273] , \zin[0][272] ,
         \zin[0][271] , \zin[0][270] , \zin[0][269] , \zin[0][268] ,
         \zin[0][267] , \zin[0][266] , \zin[0][265] , \zin[0][264] ,
         \zin[0][263] , \zin[0][262] , \zin[0][261] , \zin[0][260] ,
         \zin[0][259] , \zin[0][258] , \zin[0][257] , \zin[0][256] ,
         \zin[0][255] , \zin[0][254] , \zin[0][253] , \zin[0][252] ,
         \zin[0][251] , \zin[0][250] , \zin[0][249] , \zin[0][248] ,
         \zin[0][247] , \zin[0][246] , \zin[0][245] , \zin[0][244] ,
         \zin[0][243] , \zin[0][242] , \zin[0][241] , \zin[0][240] ,
         \zin[0][239] , \zin[0][238] , \zin[0][237] , \zin[0][236] ,
         \zin[0][235] , \zin[0][234] , \zin[0][233] , \zin[0][232] ,
         \zin[0][231] , \zin[0][230] , \zin[0][229] , \zin[0][228] ,
         \zin[0][227] , \zin[0][226] , \zin[0][225] , \zin[0][224] ,
         \zin[0][223] , \zin[0][222] , \zin[0][221] , \zin[0][220] ,
         \zin[0][219] , \zin[0][218] , \zin[0][217] , \zin[0][216] ,
         \zin[0][215] , \zin[0][214] , \zin[0][213] , \zin[0][212] ,
         \zin[0][211] , \zin[0][210] , \zin[0][209] , \zin[0][208] ,
         \zin[0][207] , \zin[0][206] , \zin[0][205] , \zin[0][204] ,
         \zin[0][203] , \zin[0][202] , \zin[0][201] , \zin[0][200] ,
         \zin[0][199] , \zin[0][198] , \zin[0][197] , \zin[0][196] ,
         \zin[0][195] , \zin[0][194] , \zin[0][193] , \zin[0][192] ,
         \zin[0][191] , \zin[0][190] , \zin[0][189] , \zin[0][188] ,
         \zin[0][187] , \zin[0][186] , \zin[0][185] , \zin[0][184] ,
         \zin[0][183] , \zin[0][182] , \zin[0][181] , \zin[0][180] ,
         \zin[0][179] , \zin[0][178] , \zin[0][177] , \zin[0][176] ,
         \zin[0][175] , \zin[0][174] , \zin[0][173] , \zin[0][172] ,
         \zin[0][171] , \zin[0][170] , \zin[0][169] , \zin[0][168] ,
         \zin[0][167] , \zin[0][166] , \zin[0][165] , \zin[0][164] ,
         \zin[0][163] , \zin[0][162] , \zin[0][161] , \zin[0][160] ,
         \zin[0][159] , \zin[0][158] , \zin[0][157] , \zin[0][156] ,
         \zin[0][155] , \zin[0][154] , \zin[0][153] , \zin[0][152] ,
         \zin[0][151] , \zin[0][150] , \zin[0][149] , \zin[0][148] ,
         \zin[0][147] , \zin[0][146] , \zin[0][145] , \zin[0][144] ,
         \zin[0][143] , \zin[0][142] , \zin[0][141] , \zin[0][140] ,
         \zin[0][139] , \zin[0][138] , \zin[0][137] , \zin[0][136] ,
         \zin[0][135] , \zin[0][134] , \zin[0][133] , \zin[0][132] ,
         \zin[0][131] , \zin[0][130] , \zin[0][129] , \zin[0][128] ,
         \zin[0][127] , \zin[0][126] , \zin[0][125] , \zin[0][124] ,
         \zin[0][123] , \zin[0][122] , \zin[0][121] , \zin[0][120] ,
         \zin[0][119] , \zin[0][118] , \zin[0][117] , \zin[0][116] ,
         \zin[0][115] , \zin[0][114] , \zin[0][113] , \zin[0][112] ,
         \zin[0][111] , \zin[0][110] , \zin[0][109] , \zin[0][108] ,
         \zin[0][107] , \zin[0][106] , \zin[0][105] , \zin[0][104] ,
         \zin[0][103] , \zin[0][102] , \zin[0][101] , \zin[0][100] ,
         \zin[0][99] , \zin[0][98] , \zin[0][97] , \zin[0][96] , \zin[0][95] ,
         \zin[0][94] , \zin[0][93] , \zin[0][92] , \zin[0][91] , \zin[0][90] ,
         \zin[0][89] , \zin[0][88] , \zin[0][87] , \zin[0][86] , \zin[0][85] ,
         \zin[0][84] , \zin[0][83] , \zin[0][82] , \zin[0][81] , \zin[0][80] ,
         \zin[0][79] , \zin[0][78] , \zin[0][77] , \zin[0][76] , \zin[0][75] ,
         \zin[0][74] , \zin[0][73] , \zin[0][72] , \zin[0][71] , \zin[0][70] ,
         \zin[0][69] , \zin[0][68] , \zin[0][67] , \zin[0][66] , \zin[0][65] ,
         \zin[0][64] , \zin[0][63] , \zin[0][62] , \zin[0][61] , \zin[0][60] ,
         \zin[0][59] , \zin[0][58] , \zin[0][57] , \zin[0][56] , \zin[0][55] ,
         \zin[0][54] , \zin[0][53] , \zin[0][52] , \zin[0][51] , \zin[0][50] ,
         \zin[0][49] , \zin[0][48] , \zin[0][47] , \zin[0][46] , \zin[0][45] ,
         \zin[0][44] , \zin[0][43] , \zin[0][42] , \zin[0][41] , \zin[0][40] ,
         \zin[0][39] , \zin[0][38] , \zin[0][37] , \zin[0][36] , \zin[0][35] ,
         \zin[0][34] , \zin[0][33] , \zin[0][32] , \zin[0][31] , \zin[0][30] ,
         \zin[0][29] , \zin[0][28] , \zin[0][27] , \zin[0][26] , \zin[0][25] ,
         \zin[0][24] , \zin[0][23] , \zin[0][22] , \zin[0][21] , \zin[0][20] ,
         \zin[0][19] , \zin[0][18] , \zin[0][17] , \zin[0][16] , \zin[0][15] ,
         \zin[0][14] , \zin[0][13] , \zin[0][12] , \zin[0][11] , \zin[0][10] ,
         \zin[0][9] , \zin[0][8] , \zin[0][7] , \zin[0][6] , \zin[0][5] ,
         \zin[0][4] , \zin[0][3] , \zin[0][2] , \zin[0][1] , \zin[0][0] , n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023;
  wire   [513:0] zreg;
  wire   [511:0] xin;
  wire   [511:0] xreg;

  DFF \xreg_reg[1]  ( .D(n1023), .CLK(clk), .RST(rst), .Q(xreg[1]) );
  DFF \xreg_reg[2]  ( .D(xin[1]), .CLK(clk), .RST(rst), .Q(xreg[2]) );
  DFF \xreg_reg[3]  ( .D(xin[2]), .CLK(clk), .RST(rst), .Q(xreg[3]) );
  DFF \xreg_reg[4]  ( .D(xin[3]), .CLK(clk), .RST(rst), .Q(xreg[4]) );
  DFF \xreg_reg[5]  ( .D(xin[4]), .CLK(clk), .RST(rst), .Q(xreg[5]) );
  DFF \xreg_reg[6]  ( .D(xin[5]), .CLK(clk), .RST(rst), .Q(xreg[6]) );
  DFF \xreg_reg[7]  ( .D(xin[6]), .CLK(clk), .RST(rst), .Q(xreg[7]) );
  DFF \xreg_reg[8]  ( .D(xin[7]), .CLK(clk), .RST(rst), .Q(xreg[8]) );
  DFF \xreg_reg[9]  ( .D(xin[8]), .CLK(clk), .RST(rst), .Q(xreg[9]) );
  DFF \xreg_reg[10]  ( .D(xin[9]), .CLK(clk), .RST(rst), .Q(xreg[10]) );
  DFF \xreg_reg[11]  ( .D(xin[10]), .CLK(clk), .RST(rst), .Q(xreg[11]) );
  DFF \xreg_reg[12]  ( .D(xin[11]), .CLK(clk), .RST(rst), .Q(xreg[12]) );
  DFF \xreg_reg[13]  ( .D(xin[12]), .CLK(clk), .RST(rst), .Q(xreg[13]) );
  DFF \xreg_reg[14]  ( .D(xin[13]), .CLK(clk), .RST(rst), .Q(xreg[14]) );
  DFF \xreg_reg[15]  ( .D(xin[14]), .CLK(clk), .RST(rst), .Q(xreg[15]) );
  DFF \xreg_reg[16]  ( .D(xin[15]), .CLK(clk), .RST(rst), .Q(xreg[16]) );
  DFF \xreg_reg[17]  ( .D(xin[16]), .CLK(clk), .RST(rst), .Q(xreg[17]) );
  DFF \xreg_reg[18]  ( .D(xin[17]), .CLK(clk), .RST(rst), .Q(xreg[18]) );
  DFF \xreg_reg[19]  ( .D(xin[18]), .CLK(clk), .RST(rst), .Q(xreg[19]) );
  DFF \xreg_reg[20]  ( .D(xin[19]), .CLK(clk), .RST(rst), .Q(xreg[20]) );
  DFF \xreg_reg[21]  ( .D(xin[20]), .CLK(clk), .RST(rst), .Q(xreg[21]) );
  DFF \xreg_reg[22]  ( .D(xin[21]), .CLK(clk), .RST(rst), .Q(xreg[22]) );
  DFF \xreg_reg[23]  ( .D(xin[22]), .CLK(clk), .RST(rst), .Q(xreg[23]) );
  DFF \xreg_reg[24]  ( .D(xin[23]), .CLK(clk), .RST(rst), .Q(xreg[24]) );
  DFF \xreg_reg[25]  ( .D(xin[24]), .CLK(clk), .RST(rst), .Q(xreg[25]) );
  DFF \xreg_reg[26]  ( .D(xin[25]), .CLK(clk), .RST(rst), .Q(xreg[26]) );
  DFF \xreg_reg[27]  ( .D(xin[26]), .CLK(clk), .RST(rst), .Q(xreg[27]) );
  DFF \xreg_reg[28]  ( .D(xin[27]), .CLK(clk), .RST(rst), .Q(xreg[28]) );
  DFF \xreg_reg[29]  ( .D(xin[28]), .CLK(clk), .RST(rst), .Q(xreg[29]) );
  DFF \xreg_reg[30]  ( .D(xin[29]), .CLK(clk), .RST(rst), .Q(xreg[30]) );
  DFF \xreg_reg[31]  ( .D(xin[30]), .CLK(clk), .RST(rst), .Q(xreg[31]) );
  DFF \xreg_reg[32]  ( .D(xin[31]), .CLK(clk), .RST(rst), .Q(xreg[32]) );
  DFF \xreg_reg[33]  ( .D(xin[32]), .CLK(clk), .RST(rst), .Q(xreg[33]) );
  DFF \xreg_reg[34]  ( .D(xin[33]), .CLK(clk), .RST(rst), .Q(xreg[34]) );
  DFF \xreg_reg[35]  ( .D(xin[34]), .CLK(clk), .RST(rst), .Q(xreg[35]) );
  DFF \xreg_reg[36]  ( .D(xin[35]), .CLK(clk), .RST(rst), .Q(xreg[36]) );
  DFF \xreg_reg[37]  ( .D(xin[36]), .CLK(clk), .RST(rst), .Q(xreg[37]) );
  DFF \xreg_reg[38]  ( .D(xin[37]), .CLK(clk), .RST(rst), .Q(xreg[38]) );
  DFF \xreg_reg[39]  ( .D(xin[38]), .CLK(clk), .RST(rst), .Q(xreg[39]) );
  DFF \xreg_reg[40]  ( .D(xin[39]), .CLK(clk), .RST(rst), .Q(xreg[40]) );
  DFF \xreg_reg[41]  ( .D(xin[40]), .CLK(clk), .RST(rst), .Q(xreg[41]) );
  DFF \xreg_reg[42]  ( .D(xin[41]), .CLK(clk), .RST(rst), .Q(xreg[42]) );
  DFF \xreg_reg[43]  ( .D(xin[42]), .CLK(clk), .RST(rst), .Q(xreg[43]) );
  DFF \xreg_reg[44]  ( .D(xin[43]), .CLK(clk), .RST(rst), .Q(xreg[44]) );
  DFF \xreg_reg[45]  ( .D(xin[44]), .CLK(clk), .RST(rst), .Q(xreg[45]) );
  DFF \xreg_reg[46]  ( .D(xin[45]), .CLK(clk), .RST(rst), .Q(xreg[46]) );
  DFF \xreg_reg[47]  ( .D(xin[46]), .CLK(clk), .RST(rst), .Q(xreg[47]) );
  DFF \xreg_reg[48]  ( .D(xin[47]), .CLK(clk), .RST(rst), .Q(xreg[48]) );
  DFF \xreg_reg[49]  ( .D(xin[48]), .CLK(clk), .RST(rst), .Q(xreg[49]) );
  DFF \xreg_reg[50]  ( .D(xin[49]), .CLK(clk), .RST(rst), .Q(xreg[50]) );
  DFF \xreg_reg[51]  ( .D(xin[50]), .CLK(clk), .RST(rst), .Q(xreg[51]) );
  DFF \xreg_reg[52]  ( .D(xin[51]), .CLK(clk), .RST(rst), .Q(xreg[52]) );
  DFF \xreg_reg[53]  ( .D(xin[52]), .CLK(clk), .RST(rst), .Q(xreg[53]) );
  DFF \xreg_reg[54]  ( .D(xin[53]), .CLK(clk), .RST(rst), .Q(xreg[54]) );
  DFF \xreg_reg[55]  ( .D(xin[54]), .CLK(clk), .RST(rst), .Q(xreg[55]) );
  DFF \xreg_reg[56]  ( .D(xin[55]), .CLK(clk), .RST(rst), .Q(xreg[56]) );
  DFF \xreg_reg[57]  ( .D(xin[56]), .CLK(clk), .RST(rst), .Q(xreg[57]) );
  DFF \xreg_reg[58]  ( .D(xin[57]), .CLK(clk), .RST(rst), .Q(xreg[58]) );
  DFF \xreg_reg[59]  ( .D(xin[58]), .CLK(clk), .RST(rst), .Q(xreg[59]) );
  DFF \xreg_reg[60]  ( .D(xin[59]), .CLK(clk), .RST(rst), .Q(xreg[60]) );
  DFF \xreg_reg[61]  ( .D(xin[60]), .CLK(clk), .RST(rst), .Q(xreg[61]) );
  DFF \xreg_reg[62]  ( .D(xin[61]), .CLK(clk), .RST(rst), .Q(xreg[62]) );
  DFF \xreg_reg[63]  ( .D(xin[62]), .CLK(clk), .RST(rst), .Q(xreg[63]) );
  DFF \xreg_reg[64]  ( .D(xin[63]), .CLK(clk), .RST(rst), .Q(xreg[64]) );
  DFF \xreg_reg[65]  ( .D(xin[64]), .CLK(clk), .RST(rst), .Q(xreg[65]) );
  DFF \xreg_reg[66]  ( .D(xin[65]), .CLK(clk), .RST(rst), .Q(xreg[66]) );
  DFF \xreg_reg[67]  ( .D(xin[66]), .CLK(clk), .RST(rst), .Q(xreg[67]) );
  DFF \xreg_reg[68]  ( .D(xin[67]), .CLK(clk), .RST(rst), .Q(xreg[68]) );
  DFF \xreg_reg[69]  ( .D(xin[68]), .CLK(clk), .RST(rst), .Q(xreg[69]) );
  DFF \xreg_reg[70]  ( .D(xin[69]), .CLK(clk), .RST(rst), .Q(xreg[70]) );
  DFF \xreg_reg[71]  ( .D(xin[70]), .CLK(clk), .RST(rst), .Q(xreg[71]) );
  DFF \xreg_reg[72]  ( .D(xin[71]), .CLK(clk), .RST(rst), .Q(xreg[72]) );
  DFF \xreg_reg[73]  ( .D(xin[72]), .CLK(clk), .RST(rst), .Q(xreg[73]) );
  DFF \xreg_reg[74]  ( .D(xin[73]), .CLK(clk), .RST(rst), .Q(xreg[74]) );
  DFF \xreg_reg[75]  ( .D(xin[74]), .CLK(clk), .RST(rst), .Q(xreg[75]) );
  DFF \xreg_reg[76]  ( .D(xin[75]), .CLK(clk), .RST(rst), .Q(xreg[76]) );
  DFF \xreg_reg[77]  ( .D(xin[76]), .CLK(clk), .RST(rst), .Q(xreg[77]) );
  DFF \xreg_reg[78]  ( .D(xin[77]), .CLK(clk), .RST(rst), .Q(xreg[78]) );
  DFF \xreg_reg[79]  ( .D(xin[78]), .CLK(clk), .RST(rst), .Q(xreg[79]) );
  DFF \xreg_reg[80]  ( .D(xin[79]), .CLK(clk), .RST(rst), .Q(xreg[80]) );
  DFF \xreg_reg[81]  ( .D(xin[80]), .CLK(clk), .RST(rst), .Q(xreg[81]) );
  DFF \xreg_reg[82]  ( .D(xin[81]), .CLK(clk), .RST(rst), .Q(xreg[82]) );
  DFF \xreg_reg[83]  ( .D(xin[82]), .CLK(clk), .RST(rst), .Q(xreg[83]) );
  DFF \xreg_reg[84]  ( .D(xin[83]), .CLK(clk), .RST(rst), .Q(xreg[84]) );
  DFF \xreg_reg[85]  ( .D(xin[84]), .CLK(clk), .RST(rst), .Q(xreg[85]) );
  DFF \xreg_reg[86]  ( .D(xin[85]), .CLK(clk), .RST(rst), .Q(xreg[86]) );
  DFF \xreg_reg[87]  ( .D(xin[86]), .CLK(clk), .RST(rst), .Q(xreg[87]) );
  DFF \xreg_reg[88]  ( .D(xin[87]), .CLK(clk), .RST(rst), .Q(xreg[88]) );
  DFF \xreg_reg[89]  ( .D(xin[88]), .CLK(clk), .RST(rst), .Q(xreg[89]) );
  DFF \xreg_reg[90]  ( .D(xin[89]), .CLK(clk), .RST(rst), .Q(xreg[90]) );
  DFF \xreg_reg[91]  ( .D(xin[90]), .CLK(clk), .RST(rst), .Q(xreg[91]) );
  DFF \xreg_reg[92]  ( .D(xin[91]), .CLK(clk), .RST(rst), .Q(xreg[92]) );
  DFF \xreg_reg[93]  ( .D(xin[92]), .CLK(clk), .RST(rst), .Q(xreg[93]) );
  DFF \xreg_reg[94]  ( .D(xin[93]), .CLK(clk), .RST(rst), .Q(xreg[94]) );
  DFF \xreg_reg[95]  ( .D(xin[94]), .CLK(clk), .RST(rst), .Q(xreg[95]) );
  DFF \xreg_reg[96]  ( .D(xin[95]), .CLK(clk), .RST(rst), .Q(xreg[96]) );
  DFF \xreg_reg[97]  ( .D(xin[96]), .CLK(clk), .RST(rst), .Q(xreg[97]) );
  DFF \xreg_reg[98]  ( .D(xin[97]), .CLK(clk), .RST(rst), .Q(xreg[98]) );
  DFF \xreg_reg[99]  ( .D(xin[98]), .CLK(clk), .RST(rst), .Q(xreg[99]) );
  DFF \xreg_reg[100]  ( .D(xin[99]), .CLK(clk), .RST(rst), .Q(xreg[100]) );
  DFF \xreg_reg[101]  ( .D(xin[100]), .CLK(clk), .RST(rst), .Q(xreg[101]) );
  DFF \xreg_reg[102]  ( .D(xin[101]), .CLK(clk), .RST(rst), .Q(xreg[102]) );
  DFF \xreg_reg[103]  ( .D(xin[102]), .CLK(clk), .RST(rst), .Q(xreg[103]) );
  DFF \xreg_reg[104]  ( .D(xin[103]), .CLK(clk), .RST(rst), .Q(xreg[104]) );
  DFF \xreg_reg[105]  ( .D(xin[104]), .CLK(clk), .RST(rst), .Q(xreg[105]) );
  DFF \xreg_reg[106]  ( .D(xin[105]), .CLK(clk), .RST(rst), .Q(xreg[106]) );
  DFF \xreg_reg[107]  ( .D(xin[106]), .CLK(clk), .RST(rst), .Q(xreg[107]) );
  DFF \xreg_reg[108]  ( .D(xin[107]), .CLK(clk), .RST(rst), .Q(xreg[108]) );
  DFF \xreg_reg[109]  ( .D(xin[108]), .CLK(clk), .RST(rst), .Q(xreg[109]) );
  DFF \xreg_reg[110]  ( .D(xin[109]), .CLK(clk), .RST(rst), .Q(xreg[110]) );
  DFF \xreg_reg[111]  ( .D(xin[110]), .CLK(clk), .RST(rst), .Q(xreg[111]) );
  DFF \xreg_reg[112]  ( .D(xin[111]), .CLK(clk), .RST(rst), .Q(xreg[112]) );
  DFF \xreg_reg[113]  ( .D(xin[112]), .CLK(clk), .RST(rst), .Q(xreg[113]) );
  DFF \xreg_reg[114]  ( .D(xin[113]), .CLK(clk), .RST(rst), .Q(xreg[114]) );
  DFF \xreg_reg[115]  ( .D(xin[114]), .CLK(clk), .RST(rst), .Q(xreg[115]) );
  DFF \xreg_reg[116]  ( .D(xin[115]), .CLK(clk), .RST(rst), .Q(xreg[116]) );
  DFF \xreg_reg[117]  ( .D(xin[116]), .CLK(clk), .RST(rst), .Q(xreg[117]) );
  DFF \xreg_reg[118]  ( .D(xin[117]), .CLK(clk), .RST(rst), .Q(xreg[118]) );
  DFF \xreg_reg[119]  ( .D(xin[118]), .CLK(clk), .RST(rst), .Q(xreg[119]) );
  DFF \xreg_reg[120]  ( .D(xin[119]), .CLK(clk), .RST(rst), .Q(xreg[120]) );
  DFF \xreg_reg[121]  ( .D(xin[120]), .CLK(clk), .RST(rst), .Q(xreg[121]) );
  DFF \xreg_reg[122]  ( .D(xin[121]), .CLK(clk), .RST(rst), .Q(xreg[122]) );
  DFF \xreg_reg[123]  ( .D(xin[122]), .CLK(clk), .RST(rst), .Q(xreg[123]) );
  DFF \xreg_reg[124]  ( .D(xin[123]), .CLK(clk), .RST(rst), .Q(xreg[124]) );
  DFF \xreg_reg[125]  ( .D(xin[124]), .CLK(clk), .RST(rst), .Q(xreg[125]) );
  DFF \xreg_reg[126]  ( .D(xin[125]), .CLK(clk), .RST(rst), .Q(xreg[126]) );
  DFF \xreg_reg[127]  ( .D(xin[126]), .CLK(clk), .RST(rst), .Q(xreg[127]) );
  DFF \xreg_reg[128]  ( .D(xin[127]), .CLK(clk), .RST(rst), .Q(xreg[128]) );
  DFF \xreg_reg[129]  ( .D(xin[128]), .CLK(clk), .RST(rst), .Q(xreg[129]) );
  DFF \xreg_reg[130]  ( .D(xin[129]), .CLK(clk), .RST(rst), .Q(xreg[130]) );
  DFF \xreg_reg[131]  ( .D(xin[130]), .CLK(clk), .RST(rst), .Q(xreg[131]) );
  DFF \xreg_reg[132]  ( .D(xin[131]), .CLK(clk), .RST(rst), .Q(xreg[132]) );
  DFF \xreg_reg[133]  ( .D(xin[132]), .CLK(clk), .RST(rst), .Q(xreg[133]) );
  DFF \xreg_reg[134]  ( .D(xin[133]), .CLK(clk), .RST(rst), .Q(xreg[134]) );
  DFF \xreg_reg[135]  ( .D(xin[134]), .CLK(clk), .RST(rst), .Q(xreg[135]) );
  DFF \xreg_reg[136]  ( .D(xin[135]), .CLK(clk), .RST(rst), .Q(xreg[136]) );
  DFF \xreg_reg[137]  ( .D(xin[136]), .CLK(clk), .RST(rst), .Q(xreg[137]) );
  DFF \xreg_reg[138]  ( .D(xin[137]), .CLK(clk), .RST(rst), .Q(xreg[138]) );
  DFF \xreg_reg[139]  ( .D(xin[138]), .CLK(clk), .RST(rst), .Q(xreg[139]) );
  DFF \xreg_reg[140]  ( .D(xin[139]), .CLK(clk), .RST(rst), .Q(xreg[140]) );
  DFF \xreg_reg[141]  ( .D(xin[140]), .CLK(clk), .RST(rst), .Q(xreg[141]) );
  DFF \xreg_reg[142]  ( .D(xin[141]), .CLK(clk), .RST(rst), .Q(xreg[142]) );
  DFF \xreg_reg[143]  ( .D(xin[142]), .CLK(clk), .RST(rst), .Q(xreg[143]) );
  DFF \xreg_reg[144]  ( .D(xin[143]), .CLK(clk), .RST(rst), .Q(xreg[144]) );
  DFF \xreg_reg[145]  ( .D(xin[144]), .CLK(clk), .RST(rst), .Q(xreg[145]) );
  DFF \xreg_reg[146]  ( .D(xin[145]), .CLK(clk), .RST(rst), .Q(xreg[146]) );
  DFF \xreg_reg[147]  ( .D(xin[146]), .CLK(clk), .RST(rst), .Q(xreg[147]) );
  DFF \xreg_reg[148]  ( .D(xin[147]), .CLK(clk), .RST(rst), .Q(xreg[148]) );
  DFF \xreg_reg[149]  ( .D(xin[148]), .CLK(clk), .RST(rst), .Q(xreg[149]) );
  DFF \xreg_reg[150]  ( .D(xin[149]), .CLK(clk), .RST(rst), .Q(xreg[150]) );
  DFF \xreg_reg[151]  ( .D(xin[150]), .CLK(clk), .RST(rst), .Q(xreg[151]) );
  DFF \xreg_reg[152]  ( .D(xin[151]), .CLK(clk), .RST(rst), .Q(xreg[152]) );
  DFF \xreg_reg[153]  ( .D(xin[152]), .CLK(clk), .RST(rst), .Q(xreg[153]) );
  DFF \xreg_reg[154]  ( .D(xin[153]), .CLK(clk), .RST(rst), .Q(xreg[154]) );
  DFF \xreg_reg[155]  ( .D(xin[154]), .CLK(clk), .RST(rst), .Q(xreg[155]) );
  DFF \xreg_reg[156]  ( .D(xin[155]), .CLK(clk), .RST(rst), .Q(xreg[156]) );
  DFF \xreg_reg[157]  ( .D(xin[156]), .CLK(clk), .RST(rst), .Q(xreg[157]) );
  DFF \xreg_reg[158]  ( .D(xin[157]), .CLK(clk), .RST(rst), .Q(xreg[158]) );
  DFF \xreg_reg[159]  ( .D(xin[158]), .CLK(clk), .RST(rst), .Q(xreg[159]) );
  DFF \xreg_reg[160]  ( .D(xin[159]), .CLK(clk), .RST(rst), .Q(xreg[160]) );
  DFF \xreg_reg[161]  ( .D(xin[160]), .CLK(clk), .RST(rst), .Q(xreg[161]) );
  DFF \xreg_reg[162]  ( .D(xin[161]), .CLK(clk), .RST(rst), .Q(xreg[162]) );
  DFF \xreg_reg[163]  ( .D(xin[162]), .CLK(clk), .RST(rst), .Q(xreg[163]) );
  DFF \xreg_reg[164]  ( .D(xin[163]), .CLK(clk), .RST(rst), .Q(xreg[164]) );
  DFF \xreg_reg[165]  ( .D(xin[164]), .CLK(clk), .RST(rst), .Q(xreg[165]) );
  DFF \xreg_reg[166]  ( .D(xin[165]), .CLK(clk), .RST(rst), .Q(xreg[166]) );
  DFF \xreg_reg[167]  ( .D(xin[166]), .CLK(clk), .RST(rst), .Q(xreg[167]) );
  DFF \xreg_reg[168]  ( .D(xin[167]), .CLK(clk), .RST(rst), .Q(xreg[168]) );
  DFF \xreg_reg[169]  ( .D(xin[168]), .CLK(clk), .RST(rst), .Q(xreg[169]) );
  DFF \xreg_reg[170]  ( .D(xin[169]), .CLK(clk), .RST(rst), .Q(xreg[170]) );
  DFF \xreg_reg[171]  ( .D(xin[170]), .CLK(clk), .RST(rst), .Q(xreg[171]) );
  DFF \xreg_reg[172]  ( .D(xin[171]), .CLK(clk), .RST(rst), .Q(xreg[172]) );
  DFF \xreg_reg[173]  ( .D(xin[172]), .CLK(clk), .RST(rst), .Q(xreg[173]) );
  DFF \xreg_reg[174]  ( .D(xin[173]), .CLK(clk), .RST(rst), .Q(xreg[174]) );
  DFF \xreg_reg[175]  ( .D(xin[174]), .CLK(clk), .RST(rst), .Q(xreg[175]) );
  DFF \xreg_reg[176]  ( .D(xin[175]), .CLK(clk), .RST(rst), .Q(xreg[176]) );
  DFF \xreg_reg[177]  ( .D(xin[176]), .CLK(clk), .RST(rst), .Q(xreg[177]) );
  DFF \xreg_reg[178]  ( .D(xin[177]), .CLK(clk), .RST(rst), .Q(xreg[178]) );
  DFF \xreg_reg[179]  ( .D(xin[178]), .CLK(clk), .RST(rst), .Q(xreg[179]) );
  DFF \xreg_reg[180]  ( .D(xin[179]), .CLK(clk), .RST(rst), .Q(xreg[180]) );
  DFF \xreg_reg[181]  ( .D(xin[180]), .CLK(clk), .RST(rst), .Q(xreg[181]) );
  DFF \xreg_reg[182]  ( .D(xin[181]), .CLK(clk), .RST(rst), .Q(xreg[182]) );
  DFF \xreg_reg[183]  ( .D(xin[182]), .CLK(clk), .RST(rst), .Q(xreg[183]) );
  DFF \xreg_reg[184]  ( .D(xin[183]), .CLK(clk), .RST(rst), .Q(xreg[184]) );
  DFF \xreg_reg[185]  ( .D(xin[184]), .CLK(clk), .RST(rst), .Q(xreg[185]) );
  DFF \xreg_reg[186]  ( .D(xin[185]), .CLK(clk), .RST(rst), .Q(xreg[186]) );
  DFF \xreg_reg[187]  ( .D(xin[186]), .CLK(clk), .RST(rst), .Q(xreg[187]) );
  DFF \xreg_reg[188]  ( .D(xin[187]), .CLK(clk), .RST(rst), .Q(xreg[188]) );
  DFF \xreg_reg[189]  ( .D(xin[188]), .CLK(clk), .RST(rst), .Q(xreg[189]) );
  DFF \xreg_reg[190]  ( .D(xin[189]), .CLK(clk), .RST(rst), .Q(xreg[190]) );
  DFF \xreg_reg[191]  ( .D(xin[190]), .CLK(clk), .RST(rst), .Q(xreg[191]) );
  DFF \xreg_reg[192]  ( .D(xin[191]), .CLK(clk), .RST(rst), .Q(xreg[192]) );
  DFF \xreg_reg[193]  ( .D(xin[192]), .CLK(clk), .RST(rst), .Q(xreg[193]) );
  DFF \xreg_reg[194]  ( .D(xin[193]), .CLK(clk), .RST(rst), .Q(xreg[194]) );
  DFF \xreg_reg[195]  ( .D(xin[194]), .CLK(clk), .RST(rst), .Q(xreg[195]) );
  DFF \xreg_reg[196]  ( .D(xin[195]), .CLK(clk), .RST(rst), .Q(xreg[196]) );
  DFF \xreg_reg[197]  ( .D(xin[196]), .CLK(clk), .RST(rst), .Q(xreg[197]) );
  DFF \xreg_reg[198]  ( .D(xin[197]), .CLK(clk), .RST(rst), .Q(xreg[198]) );
  DFF \xreg_reg[199]  ( .D(xin[198]), .CLK(clk), .RST(rst), .Q(xreg[199]) );
  DFF \xreg_reg[200]  ( .D(xin[199]), .CLK(clk), .RST(rst), .Q(xreg[200]) );
  DFF \xreg_reg[201]  ( .D(xin[200]), .CLK(clk), .RST(rst), .Q(xreg[201]) );
  DFF \xreg_reg[202]  ( .D(xin[201]), .CLK(clk), .RST(rst), .Q(xreg[202]) );
  DFF \xreg_reg[203]  ( .D(xin[202]), .CLK(clk), .RST(rst), .Q(xreg[203]) );
  DFF \xreg_reg[204]  ( .D(xin[203]), .CLK(clk), .RST(rst), .Q(xreg[204]) );
  DFF \xreg_reg[205]  ( .D(xin[204]), .CLK(clk), .RST(rst), .Q(xreg[205]) );
  DFF \xreg_reg[206]  ( .D(xin[205]), .CLK(clk), .RST(rst), .Q(xreg[206]) );
  DFF \xreg_reg[207]  ( .D(xin[206]), .CLK(clk), .RST(rst), .Q(xreg[207]) );
  DFF \xreg_reg[208]  ( .D(xin[207]), .CLK(clk), .RST(rst), .Q(xreg[208]) );
  DFF \xreg_reg[209]  ( .D(xin[208]), .CLK(clk), .RST(rst), .Q(xreg[209]) );
  DFF \xreg_reg[210]  ( .D(xin[209]), .CLK(clk), .RST(rst), .Q(xreg[210]) );
  DFF \xreg_reg[211]  ( .D(xin[210]), .CLK(clk), .RST(rst), .Q(xreg[211]) );
  DFF \xreg_reg[212]  ( .D(xin[211]), .CLK(clk), .RST(rst), .Q(xreg[212]) );
  DFF \xreg_reg[213]  ( .D(xin[212]), .CLK(clk), .RST(rst), .Q(xreg[213]) );
  DFF \xreg_reg[214]  ( .D(xin[213]), .CLK(clk), .RST(rst), .Q(xreg[214]) );
  DFF \xreg_reg[215]  ( .D(xin[214]), .CLK(clk), .RST(rst), .Q(xreg[215]) );
  DFF \xreg_reg[216]  ( .D(xin[215]), .CLK(clk), .RST(rst), .Q(xreg[216]) );
  DFF \xreg_reg[217]  ( .D(xin[216]), .CLK(clk), .RST(rst), .Q(xreg[217]) );
  DFF \xreg_reg[218]  ( .D(xin[217]), .CLK(clk), .RST(rst), .Q(xreg[218]) );
  DFF \xreg_reg[219]  ( .D(xin[218]), .CLK(clk), .RST(rst), .Q(xreg[219]) );
  DFF \xreg_reg[220]  ( .D(xin[219]), .CLK(clk), .RST(rst), .Q(xreg[220]) );
  DFF \xreg_reg[221]  ( .D(xin[220]), .CLK(clk), .RST(rst), .Q(xreg[221]) );
  DFF \xreg_reg[222]  ( .D(xin[221]), .CLK(clk), .RST(rst), .Q(xreg[222]) );
  DFF \xreg_reg[223]  ( .D(xin[222]), .CLK(clk), .RST(rst), .Q(xreg[223]) );
  DFF \xreg_reg[224]  ( .D(xin[223]), .CLK(clk), .RST(rst), .Q(xreg[224]) );
  DFF \xreg_reg[225]  ( .D(xin[224]), .CLK(clk), .RST(rst), .Q(xreg[225]) );
  DFF \xreg_reg[226]  ( .D(xin[225]), .CLK(clk), .RST(rst), .Q(xreg[226]) );
  DFF \xreg_reg[227]  ( .D(xin[226]), .CLK(clk), .RST(rst), .Q(xreg[227]) );
  DFF \xreg_reg[228]  ( .D(xin[227]), .CLK(clk), .RST(rst), .Q(xreg[228]) );
  DFF \xreg_reg[229]  ( .D(xin[228]), .CLK(clk), .RST(rst), .Q(xreg[229]) );
  DFF \xreg_reg[230]  ( .D(xin[229]), .CLK(clk), .RST(rst), .Q(xreg[230]) );
  DFF \xreg_reg[231]  ( .D(xin[230]), .CLK(clk), .RST(rst), .Q(xreg[231]) );
  DFF \xreg_reg[232]  ( .D(xin[231]), .CLK(clk), .RST(rst), .Q(xreg[232]) );
  DFF \xreg_reg[233]  ( .D(xin[232]), .CLK(clk), .RST(rst), .Q(xreg[233]) );
  DFF \xreg_reg[234]  ( .D(xin[233]), .CLK(clk), .RST(rst), .Q(xreg[234]) );
  DFF \xreg_reg[235]  ( .D(xin[234]), .CLK(clk), .RST(rst), .Q(xreg[235]) );
  DFF \xreg_reg[236]  ( .D(xin[235]), .CLK(clk), .RST(rst), .Q(xreg[236]) );
  DFF \xreg_reg[237]  ( .D(xin[236]), .CLK(clk), .RST(rst), .Q(xreg[237]) );
  DFF \xreg_reg[238]  ( .D(xin[237]), .CLK(clk), .RST(rst), .Q(xreg[238]) );
  DFF \xreg_reg[239]  ( .D(xin[238]), .CLK(clk), .RST(rst), .Q(xreg[239]) );
  DFF \xreg_reg[240]  ( .D(xin[239]), .CLK(clk), .RST(rst), .Q(xreg[240]) );
  DFF \xreg_reg[241]  ( .D(xin[240]), .CLK(clk), .RST(rst), .Q(xreg[241]) );
  DFF \xreg_reg[242]  ( .D(xin[241]), .CLK(clk), .RST(rst), .Q(xreg[242]) );
  DFF \xreg_reg[243]  ( .D(xin[242]), .CLK(clk), .RST(rst), .Q(xreg[243]) );
  DFF \xreg_reg[244]  ( .D(xin[243]), .CLK(clk), .RST(rst), .Q(xreg[244]) );
  DFF \xreg_reg[245]  ( .D(xin[244]), .CLK(clk), .RST(rst), .Q(xreg[245]) );
  DFF \xreg_reg[246]  ( .D(xin[245]), .CLK(clk), .RST(rst), .Q(xreg[246]) );
  DFF \xreg_reg[247]  ( .D(xin[246]), .CLK(clk), .RST(rst), .Q(xreg[247]) );
  DFF \xreg_reg[248]  ( .D(xin[247]), .CLK(clk), .RST(rst), .Q(xreg[248]) );
  DFF \xreg_reg[249]  ( .D(xin[248]), .CLK(clk), .RST(rst), .Q(xreg[249]) );
  DFF \xreg_reg[250]  ( .D(xin[249]), .CLK(clk), .RST(rst), .Q(xreg[250]) );
  DFF \xreg_reg[251]  ( .D(xin[250]), .CLK(clk), .RST(rst), .Q(xreg[251]) );
  DFF \xreg_reg[252]  ( .D(xin[251]), .CLK(clk), .RST(rst), .Q(xreg[252]) );
  DFF \xreg_reg[253]  ( .D(xin[252]), .CLK(clk), .RST(rst), .Q(xreg[253]) );
  DFF \xreg_reg[254]  ( .D(xin[253]), .CLK(clk), .RST(rst), .Q(xreg[254]) );
  DFF \xreg_reg[255]  ( .D(xin[254]), .CLK(clk), .RST(rst), .Q(xreg[255]) );
  DFF \xreg_reg[256]  ( .D(xin[255]), .CLK(clk), .RST(rst), .Q(xreg[256]) );
  DFF \xreg_reg[257]  ( .D(xin[256]), .CLK(clk), .RST(rst), .Q(xreg[257]) );
  DFF \xreg_reg[258]  ( .D(xin[257]), .CLK(clk), .RST(rst), .Q(xreg[258]) );
  DFF \xreg_reg[259]  ( .D(xin[258]), .CLK(clk), .RST(rst), .Q(xreg[259]) );
  DFF \xreg_reg[260]  ( .D(xin[259]), .CLK(clk), .RST(rst), .Q(xreg[260]) );
  DFF \xreg_reg[261]  ( .D(xin[260]), .CLK(clk), .RST(rst), .Q(xreg[261]) );
  DFF \xreg_reg[262]  ( .D(xin[261]), .CLK(clk), .RST(rst), .Q(xreg[262]) );
  DFF \xreg_reg[263]  ( .D(xin[262]), .CLK(clk), .RST(rst), .Q(xreg[263]) );
  DFF \xreg_reg[264]  ( .D(xin[263]), .CLK(clk), .RST(rst), .Q(xreg[264]) );
  DFF \xreg_reg[265]  ( .D(xin[264]), .CLK(clk), .RST(rst), .Q(xreg[265]) );
  DFF \xreg_reg[266]  ( .D(xin[265]), .CLK(clk), .RST(rst), .Q(xreg[266]) );
  DFF \xreg_reg[267]  ( .D(xin[266]), .CLK(clk), .RST(rst), .Q(xreg[267]) );
  DFF \xreg_reg[268]  ( .D(xin[267]), .CLK(clk), .RST(rst), .Q(xreg[268]) );
  DFF \xreg_reg[269]  ( .D(xin[268]), .CLK(clk), .RST(rst), .Q(xreg[269]) );
  DFF \xreg_reg[270]  ( .D(xin[269]), .CLK(clk), .RST(rst), .Q(xreg[270]) );
  DFF \xreg_reg[271]  ( .D(xin[270]), .CLK(clk), .RST(rst), .Q(xreg[271]) );
  DFF \xreg_reg[272]  ( .D(xin[271]), .CLK(clk), .RST(rst), .Q(xreg[272]) );
  DFF \xreg_reg[273]  ( .D(xin[272]), .CLK(clk), .RST(rst), .Q(xreg[273]) );
  DFF \xreg_reg[274]  ( .D(xin[273]), .CLK(clk), .RST(rst), .Q(xreg[274]) );
  DFF \xreg_reg[275]  ( .D(xin[274]), .CLK(clk), .RST(rst), .Q(xreg[275]) );
  DFF \xreg_reg[276]  ( .D(xin[275]), .CLK(clk), .RST(rst), .Q(xreg[276]) );
  DFF \xreg_reg[277]  ( .D(xin[276]), .CLK(clk), .RST(rst), .Q(xreg[277]) );
  DFF \xreg_reg[278]  ( .D(xin[277]), .CLK(clk), .RST(rst), .Q(xreg[278]) );
  DFF \xreg_reg[279]  ( .D(xin[278]), .CLK(clk), .RST(rst), .Q(xreg[279]) );
  DFF \xreg_reg[280]  ( .D(xin[279]), .CLK(clk), .RST(rst), .Q(xreg[280]) );
  DFF \xreg_reg[281]  ( .D(xin[280]), .CLK(clk), .RST(rst), .Q(xreg[281]) );
  DFF \xreg_reg[282]  ( .D(xin[281]), .CLK(clk), .RST(rst), .Q(xreg[282]) );
  DFF \xreg_reg[283]  ( .D(xin[282]), .CLK(clk), .RST(rst), .Q(xreg[283]) );
  DFF \xreg_reg[284]  ( .D(xin[283]), .CLK(clk), .RST(rst), .Q(xreg[284]) );
  DFF \xreg_reg[285]  ( .D(xin[284]), .CLK(clk), .RST(rst), .Q(xreg[285]) );
  DFF \xreg_reg[286]  ( .D(xin[285]), .CLK(clk), .RST(rst), .Q(xreg[286]) );
  DFF \xreg_reg[287]  ( .D(xin[286]), .CLK(clk), .RST(rst), .Q(xreg[287]) );
  DFF \xreg_reg[288]  ( .D(xin[287]), .CLK(clk), .RST(rst), .Q(xreg[288]) );
  DFF \xreg_reg[289]  ( .D(xin[288]), .CLK(clk), .RST(rst), .Q(xreg[289]) );
  DFF \xreg_reg[290]  ( .D(xin[289]), .CLK(clk), .RST(rst), .Q(xreg[290]) );
  DFF \xreg_reg[291]  ( .D(xin[290]), .CLK(clk), .RST(rst), .Q(xreg[291]) );
  DFF \xreg_reg[292]  ( .D(xin[291]), .CLK(clk), .RST(rst), .Q(xreg[292]) );
  DFF \xreg_reg[293]  ( .D(xin[292]), .CLK(clk), .RST(rst), .Q(xreg[293]) );
  DFF \xreg_reg[294]  ( .D(xin[293]), .CLK(clk), .RST(rst), .Q(xreg[294]) );
  DFF \xreg_reg[295]  ( .D(xin[294]), .CLK(clk), .RST(rst), .Q(xreg[295]) );
  DFF \xreg_reg[296]  ( .D(xin[295]), .CLK(clk), .RST(rst), .Q(xreg[296]) );
  DFF \xreg_reg[297]  ( .D(xin[296]), .CLK(clk), .RST(rst), .Q(xreg[297]) );
  DFF \xreg_reg[298]  ( .D(xin[297]), .CLK(clk), .RST(rst), .Q(xreg[298]) );
  DFF \xreg_reg[299]  ( .D(xin[298]), .CLK(clk), .RST(rst), .Q(xreg[299]) );
  DFF \xreg_reg[300]  ( .D(xin[299]), .CLK(clk), .RST(rst), .Q(xreg[300]) );
  DFF \xreg_reg[301]  ( .D(xin[300]), .CLK(clk), .RST(rst), .Q(xreg[301]) );
  DFF \xreg_reg[302]  ( .D(xin[301]), .CLK(clk), .RST(rst), .Q(xreg[302]) );
  DFF \xreg_reg[303]  ( .D(xin[302]), .CLK(clk), .RST(rst), .Q(xreg[303]) );
  DFF \xreg_reg[304]  ( .D(xin[303]), .CLK(clk), .RST(rst), .Q(xreg[304]) );
  DFF \xreg_reg[305]  ( .D(xin[304]), .CLK(clk), .RST(rst), .Q(xreg[305]) );
  DFF \xreg_reg[306]  ( .D(xin[305]), .CLK(clk), .RST(rst), .Q(xreg[306]) );
  DFF \xreg_reg[307]  ( .D(xin[306]), .CLK(clk), .RST(rst), .Q(xreg[307]) );
  DFF \xreg_reg[308]  ( .D(xin[307]), .CLK(clk), .RST(rst), .Q(xreg[308]) );
  DFF \xreg_reg[309]  ( .D(xin[308]), .CLK(clk), .RST(rst), .Q(xreg[309]) );
  DFF \xreg_reg[310]  ( .D(xin[309]), .CLK(clk), .RST(rst), .Q(xreg[310]) );
  DFF \xreg_reg[311]  ( .D(xin[310]), .CLK(clk), .RST(rst), .Q(xreg[311]) );
  DFF \xreg_reg[312]  ( .D(xin[311]), .CLK(clk), .RST(rst), .Q(xreg[312]) );
  DFF \xreg_reg[313]  ( .D(xin[312]), .CLK(clk), .RST(rst), .Q(xreg[313]) );
  DFF \xreg_reg[314]  ( .D(xin[313]), .CLK(clk), .RST(rst), .Q(xreg[314]) );
  DFF \xreg_reg[315]  ( .D(xin[314]), .CLK(clk), .RST(rst), .Q(xreg[315]) );
  DFF \xreg_reg[316]  ( .D(xin[315]), .CLK(clk), .RST(rst), .Q(xreg[316]) );
  DFF \xreg_reg[317]  ( .D(xin[316]), .CLK(clk), .RST(rst), .Q(xreg[317]) );
  DFF \xreg_reg[318]  ( .D(xin[317]), .CLK(clk), .RST(rst), .Q(xreg[318]) );
  DFF \xreg_reg[319]  ( .D(xin[318]), .CLK(clk), .RST(rst), .Q(xreg[319]) );
  DFF \xreg_reg[320]  ( .D(xin[319]), .CLK(clk), .RST(rst), .Q(xreg[320]) );
  DFF \xreg_reg[321]  ( .D(xin[320]), .CLK(clk), .RST(rst), .Q(xreg[321]) );
  DFF \xreg_reg[322]  ( .D(xin[321]), .CLK(clk), .RST(rst), .Q(xreg[322]) );
  DFF \xreg_reg[323]  ( .D(xin[322]), .CLK(clk), .RST(rst), .Q(xreg[323]) );
  DFF \xreg_reg[324]  ( .D(xin[323]), .CLK(clk), .RST(rst), .Q(xreg[324]) );
  DFF \xreg_reg[325]  ( .D(xin[324]), .CLK(clk), .RST(rst), .Q(xreg[325]) );
  DFF \xreg_reg[326]  ( .D(xin[325]), .CLK(clk), .RST(rst), .Q(xreg[326]) );
  DFF \xreg_reg[327]  ( .D(xin[326]), .CLK(clk), .RST(rst), .Q(xreg[327]) );
  DFF \xreg_reg[328]  ( .D(xin[327]), .CLK(clk), .RST(rst), .Q(xreg[328]) );
  DFF \xreg_reg[329]  ( .D(xin[328]), .CLK(clk), .RST(rst), .Q(xreg[329]) );
  DFF \xreg_reg[330]  ( .D(xin[329]), .CLK(clk), .RST(rst), .Q(xreg[330]) );
  DFF \xreg_reg[331]  ( .D(xin[330]), .CLK(clk), .RST(rst), .Q(xreg[331]) );
  DFF \xreg_reg[332]  ( .D(xin[331]), .CLK(clk), .RST(rst), .Q(xreg[332]) );
  DFF \xreg_reg[333]  ( .D(xin[332]), .CLK(clk), .RST(rst), .Q(xreg[333]) );
  DFF \xreg_reg[334]  ( .D(xin[333]), .CLK(clk), .RST(rst), .Q(xreg[334]) );
  DFF \xreg_reg[335]  ( .D(xin[334]), .CLK(clk), .RST(rst), .Q(xreg[335]) );
  DFF \xreg_reg[336]  ( .D(xin[335]), .CLK(clk), .RST(rst), .Q(xreg[336]) );
  DFF \xreg_reg[337]  ( .D(xin[336]), .CLK(clk), .RST(rst), .Q(xreg[337]) );
  DFF \xreg_reg[338]  ( .D(xin[337]), .CLK(clk), .RST(rst), .Q(xreg[338]) );
  DFF \xreg_reg[339]  ( .D(xin[338]), .CLK(clk), .RST(rst), .Q(xreg[339]) );
  DFF \xreg_reg[340]  ( .D(xin[339]), .CLK(clk), .RST(rst), .Q(xreg[340]) );
  DFF \xreg_reg[341]  ( .D(xin[340]), .CLK(clk), .RST(rst), .Q(xreg[341]) );
  DFF \xreg_reg[342]  ( .D(xin[341]), .CLK(clk), .RST(rst), .Q(xreg[342]) );
  DFF \xreg_reg[343]  ( .D(xin[342]), .CLK(clk), .RST(rst), .Q(xreg[343]) );
  DFF \xreg_reg[344]  ( .D(xin[343]), .CLK(clk), .RST(rst), .Q(xreg[344]) );
  DFF \xreg_reg[345]  ( .D(xin[344]), .CLK(clk), .RST(rst), .Q(xreg[345]) );
  DFF \xreg_reg[346]  ( .D(xin[345]), .CLK(clk), .RST(rst), .Q(xreg[346]) );
  DFF \xreg_reg[347]  ( .D(xin[346]), .CLK(clk), .RST(rst), .Q(xreg[347]) );
  DFF \xreg_reg[348]  ( .D(xin[347]), .CLK(clk), .RST(rst), .Q(xreg[348]) );
  DFF \xreg_reg[349]  ( .D(xin[348]), .CLK(clk), .RST(rst), .Q(xreg[349]) );
  DFF \xreg_reg[350]  ( .D(xin[349]), .CLK(clk), .RST(rst), .Q(xreg[350]) );
  DFF \xreg_reg[351]  ( .D(xin[350]), .CLK(clk), .RST(rst), .Q(xreg[351]) );
  DFF \xreg_reg[352]  ( .D(xin[351]), .CLK(clk), .RST(rst), .Q(xreg[352]) );
  DFF \xreg_reg[353]  ( .D(xin[352]), .CLK(clk), .RST(rst), .Q(xreg[353]) );
  DFF \xreg_reg[354]  ( .D(xin[353]), .CLK(clk), .RST(rst), .Q(xreg[354]) );
  DFF \xreg_reg[355]  ( .D(xin[354]), .CLK(clk), .RST(rst), .Q(xreg[355]) );
  DFF \xreg_reg[356]  ( .D(xin[355]), .CLK(clk), .RST(rst), .Q(xreg[356]) );
  DFF \xreg_reg[357]  ( .D(xin[356]), .CLK(clk), .RST(rst), .Q(xreg[357]) );
  DFF \xreg_reg[358]  ( .D(xin[357]), .CLK(clk), .RST(rst), .Q(xreg[358]) );
  DFF \xreg_reg[359]  ( .D(xin[358]), .CLK(clk), .RST(rst), .Q(xreg[359]) );
  DFF \xreg_reg[360]  ( .D(xin[359]), .CLK(clk), .RST(rst), .Q(xreg[360]) );
  DFF \xreg_reg[361]  ( .D(xin[360]), .CLK(clk), .RST(rst), .Q(xreg[361]) );
  DFF \xreg_reg[362]  ( .D(xin[361]), .CLK(clk), .RST(rst), .Q(xreg[362]) );
  DFF \xreg_reg[363]  ( .D(xin[362]), .CLK(clk), .RST(rst), .Q(xreg[363]) );
  DFF \xreg_reg[364]  ( .D(xin[363]), .CLK(clk), .RST(rst), .Q(xreg[364]) );
  DFF \xreg_reg[365]  ( .D(xin[364]), .CLK(clk), .RST(rst), .Q(xreg[365]) );
  DFF \xreg_reg[366]  ( .D(xin[365]), .CLK(clk), .RST(rst), .Q(xreg[366]) );
  DFF \xreg_reg[367]  ( .D(xin[366]), .CLK(clk), .RST(rst), .Q(xreg[367]) );
  DFF \xreg_reg[368]  ( .D(xin[367]), .CLK(clk), .RST(rst), .Q(xreg[368]) );
  DFF \xreg_reg[369]  ( .D(xin[368]), .CLK(clk), .RST(rst), .Q(xreg[369]) );
  DFF \xreg_reg[370]  ( .D(xin[369]), .CLK(clk), .RST(rst), .Q(xreg[370]) );
  DFF \xreg_reg[371]  ( .D(xin[370]), .CLK(clk), .RST(rst), .Q(xreg[371]) );
  DFF \xreg_reg[372]  ( .D(xin[371]), .CLK(clk), .RST(rst), .Q(xreg[372]) );
  DFF \xreg_reg[373]  ( .D(xin[372]), .CLK(clk), .RST(rst), .Q(xreg[373]) );
  DFF \xreg_reg[374]  ( .D(xin[373]), .CLK(clk), .RST(rst), .Q(xreg[374]) );
  DFF \xreg_reg[375]  ( .D(xin[374]), .CLK(clk), .RST(rst), .Q(xreg[375]) );
  DFF \xreg_reg[376]  ( .D(xin[375]), .CLK(clk), .RST(rst), .Q(xreg[376]) );
  DFF \xreg_reg[377]  ( .D(xin[376]), .CLK(clk), .RST(rst), .Q(xreg[377]) );
  DFF \xreg_reg[378]  ( .D(xin[377]), .CLK(clk), .RST(rst), .Q(xreg[378]) );
  DFF \xreg_reg[379]  ( .D(xin[378]), .CLK(clk), .RST(rst), .Q(xreg[379]) );
  DFF \xreg_reg[380]  ( .D(xin[379]), .CLK(clk), .RST(rst), .Q(xreg[380]) );
  DFF \xreg_reg[381]  ( .D(xin[380]), .CLK(clk), .RST(rst), .Q(xreg[381]) );
  DFF \xreg_reg[382]  ( .D(xin[381]), .CLK(clk), .RST(rst), .Q(xreg[382]) );
  DFF \xreg_reg[383]  ( .D(xin[382]), .CLK(clk), .RST(rst), .Q(xreg[383]) );
  DFF \xreg_reg[384]  ( .D(xin[383]), .CLK(clk), .RST(rst), .Q(xreg[384]) );
  DFF \xreg_reg[385]  ( .D(xin[384]), .CLK(clk), .RST(rst), .Q(xreg[385]) );
  DFF \xreg_reg[386]  ( .D(xin[385]), .CLK(clk), .RST(rst), .Q(xreg[386]) );
  DFF \xreg_reg[387]  ( .D(xin[386]), .CLK(clk), .RST(rst), .Q(xreg[387]) );
  DFF \xreg_reg[388]  ( .D(xin[387]), .CLK(clk), .RST(rst), .Q(xreg[388]) );
  DFF \xreg_reg[389]  ( .D(xin[388]), .CLK(clk), .RST(rst), .Q(xreg[389]) );
  DFF \xreg_reg[390]  ( .D(xin[389]), .CLK(clk), .RST(rst), .Q(xreg[390]) );
  DFF \xreg_reg[391]  ( .D(xin[390]), .CLK(clk), .RST(rst), .Q(xreg[391]) );
  DFF \xreg_reg[392]  ( .D(xin[391]), .CLK(clk), .RST(rst), .Q(xreg[392]) );
  DFF \xreg_reg[393]  ( .D(xin[392]), .CLK(clk), .RST(rst), .Q(xreg[393]) );
  DFF \xreg_reg[394]  ( .D(xin[393]), .CLK(clk), .RST(rst), .Q(xreg[394]) );
  DFF \xreg_reg[395]  ( .D(xin[394]), .CLK(clk), .RST(rst), .Q(xreg[395]) );
  DFF \xreg_reg[396]  ( .D(xin[395]), .CLK(clk), .RST(rst), .Q(xreg[396]) );
  DFF \xreg_reg[397]  ( .D(xin[396]), .CLK(clk), .RST(rst), .Q(xreg[397]) );
  DFF \xreg_reg[398]  ( .D(xin[397]), .CLK(clk), .RST(rst), .Q(xreg[398]) );
  DFF \xreg_reg[399]  ( .D(xin[398]), .CLK(clk), .RST(rst), .Q(xreg[399]) );
  DFF \xreg_reg[400]  ( .D(xin[399]), .CLK(clk), .RST(rst), .Q(xreg[400]) );
  DFF \xreg_reg[401]  ( .D(xin[400]), .CLK(clk), .RST(rst), .Q(xreg[401]) );
  DFF \xreg_reg[402]  ( .D(xin[401]), .CLK(clk), .RST(rst), .Q(xreg[402]) );
  DFF \xreg_reg[403]  ( .D(xin[402]), .CLK(clk), .RST(rst), .Q(xreg[403]) );
  DFF \xreg_reg[404]  ( .D(xin[403]), .CLK(clk), .RST(rst), .Q(xreg[404]) );
  DFF \xreg_reg[405]  ( .D(xin[404]), .CLK(clk), .RST(rst), .Q(xreg[405]) );
  DFF \xreg_reg[406]  ( .D(xin[405]), .CLK(clk), .RST(rst), .Q(xreg[406]) );
  DFF \xreg_reg[407]  ( .D(xin[406]), .CLK(clk), .RST(rst), .Q(xreg[407]) );
  DFF \xreg_reg[408]  ( .D(xin[407]), .CLK(clk), .RST(rst), .Q(xreg[408]) );
  DFF \xreg_reg[409]  ( .D(xin[408]), .CLK(clk), .RST(rst), .Q(xreg[409]) );
  DFF \xreg_reg[410]  ( .D(xin[409]), .CLK(clk), .RST(rst), .Q(xreg[410]) );
  DFF \xreg_reg[411]  ( .D(xin[410]), .CLK(clk), .RST(rst), .Q(xreg[411]) );
  DFF \xreg_reg[412]  ( .D(xin[411]), .CLK(clk), .RST(rst), .Q(xreg[412]) );
  DFF \xreg_reg[413]  ( .D(xin[412]), .CLK(clk), .RST(rst), .Q(xreg[413]) );
  DFF \xreg_reg[414]  ( .D(xin[413]), .CLK(clk), .RST(rst), .Q(xreg[414]) );
  DFF \xreg_reg[415]  ( .D(xin[414]), .CLK(clk), .RST(rst), .Q(xreg[415]) );
  DFF \xreg_reg[416]  ( .D(xin[415]), .CLK(clk), .RST(rst), .Q(xreg[416]) );
  DFF \xreg_reg[417]  ( .D(xin[416]), .CLK(clk), .RST(rst), .Q(xreg[417]) );
  DFF \xreg_reg[418]  ( .D(xin[417]), .CLK(clk), .RST(rst), .Q(xreg[418]) );
  DFF \xreg_reg[419]  ( .D(xin[418]), .CLK(clk), .RST(rst), .Q(xreg[419]) );
  DFF \xreg_reg[420]  ( .D(xin[419]), .CLK(clk), .RST(rst), .Q(xreg[420]) );
  DFF \xreg_reg[421]  ( .D(xin[420]), .CLK(clk), .RST(rst), .Q(xreg[421]) );
  DFF \xreg_reg[422]  ( .D(xin[421]), .CLK(clk), .RST(rst), .Q(xreg[422]) );
  DFF \xreg_reg[423]  ( .D(xin[422]), .CLK(clk), .RST(rst), .Q(xreg[423]) );
  DFF \xreg_reg[424]  ( .D(xin[423]), .CLK(clk), .RST(rst), .Q(xreg[424]) );
  DFF \xreg_reg[425]  ( .D(xin[424]), .CLK(clk), .RST(rst), .Q(xreg[425]) );
  DFF \xreg_reg[426]  ( .D(xin[425]), .CLK(clk), .RST(rst), .Q(xreg[426]) );
  DFF \xreg_reg[427]  ( .D(xin[426]), .CLK(clk), .RST(rst), .Q(xreg[427]) );
  DFF \xreg_reg[428]  ( .D(xin[427]), .CLK(clk), .RST(rst), .Q(xreg[428]) );
  DFF \xreg_reg[429]  ( .D(xin[428]), .CLK(clk), .RST(rst), .Q(xreg[429]) );
  DFF \xreg_reg[430]  ( .D(xin[429]), .CLK(clk), .RST(rst), .Q(xreg[430]) );
  DFF \xreg_reg[431]  ( .D(xin[430]), .CLK(clk), .RST(rst), .Q(xreg[431]) );
  DFF \xreg_reg[432]  ( .D(xin[431]), .CLK(clk), .RST(rst), .Q(xreg[432]) );
  DFF \xreg_reg[433]  ( .D(xin[432]), .CLK(clk), .RST(rst), .Q(xreg[433]) );
  DFF \xreg_reg[434]  ( .D(xin[433]), .CLK(clk), .RST(rst), .Q(xreg[434]) );
  DFF \xreg_reg[435]  ( .D(xin[434]), .CLK(clk), .RST(rst), .Q(xreg[435]) );
  DFF \xreg_reg[436]  ( .D(xin[435]), .CLK(clk), .RST(rst), .Q(xreg[436]) );
  DFF \xreg_reg[437]  ( .D(xin[436]), .CLK(clk), .RST(rst), .Q(xreg[437]) );
  DFF \xreg_reg[438]  ( .D(xin[437]), .CLK(clk), .RST(rst), .Q(xreg[438]) );
  DFF \xreg_reg[439]  ( .D(xin[438]), .CLK(clk), .RST(rst), .Q(xreg[439]) );
  DFF \xreg_reg[440]  ( .D(xin[439]), .CLK(clk), .RST(rst), .Q(xreg[440]) );
  DFF \xreg_reg[441]  ( .D(xin[440]), .CLK(clk), .RST(rst), .Q(xreg[441]) );
  DFF \xreg_reg[442]  ( .D(xin[441]), .CLK(clk), .RST(rst), .Q(xreg[442]) );
  DFF \xreg_reg[443]  ( .D(xin[442]), .CLK(clk), .RST(rst), .Q(xreg[443]) );
  DFF \xreg_reg[444]  ( .D(xin[443]), .CLK(clk), .RST(rst), .Q(xreg[444]) );
  DFF \xreg_reg[445]  ( .D(xin[444]), .CLK(clk), .RST(rst), .Q(xreg[445]) );
  DFF \xreg_reg[446]  ( .D(xin[445]), .CLK(clk), .RST(rst), .Q(xreg[446]) );
  DFF \xreg_reg[447]  ( .D(xin[446]), .CLK(clk), .RST(rst), .Q(xreg[447]) );
  DFF \xreg_reg[448]  ( .D(xin[447]), .CLK(clk), .RST(rst), .Q(xreg[448]) );
  DFF \xreg_reg[449]  ( .D(xin[448]), .CLK(clk), .RST(rst), .Q(xreg[449]) );
  DFF \xreg_reg[450]  ( .D(xin[449]), .CLK(clk), .RST(rst), .Q(xreg[450]) );
  DFF \xreg_reg[451]  ( .D(xin[450]), .CLK(clk), .RST(rst), .Q(xreg[451]) );
  DFF \xreg_reg[452]  ( .D(xin[451]), .CLK(clk), .RST(rst), .Q(xreg[452]) );
  DFF \xreg_reg[453]  ( .D(xin[452]), .CLK(clk), .RST(rst), .Q(xreg[453]) );
  DFF \xreg_reg[454]  ( .D(xin[453]), .CLK(clk), .RST(rst), .Q(xreg[454]) );
  DFF \xreg_reg[455]  ( .D(xin[454]), .CLK(clk), .RST(rst), .Q(xreg[455]) );
  DFF \xreg_reg[456]  ( .D(xin[455]), .CLK(clk), .RST(rst), .Q(xreg[456]) );
  DFF \xreg_reg[457]  ( .D(xin[456]), .CLK(clk), .RST(rst), .Q(xreg[457]) );
  DFF \xreg_reg[458]  ( .D(xin[457]), .CLK(clk), .RST(rst), .Q(xreg[458]) );
  DFF \xreg_reg[459]  ( .D(xin[458]), .CLK(clk), .RST(rst), .Q(xreg[459]) );
  DFF \xreg_reg[460]  ( .D(xin[459]), .CLK(clk), .RST(rst), .Q(xreg[460]) );
  DFF \xreg_reg[461]  ( .D(xin[460]), .CLK(clk), .RST(rst), .Q(xreg[461]) );
  DFF \xreg_reg[462]  ( .D(xin[461]), .CLK(clk), .RST(rst), .Q(xreg[462]) );
  DFF \xreg_reg[463]  ( .D(xin[462]), .CLK(clk), .RST(rst), .Q(xreg[463]) );
  DFF \xreg_reg[464]  ( .D(xin[463]), .CLK(clk), .RST(rst), .Q(xreg[464]) );
  DFF \xreg_reg[465]  ( .D(xin[464]), .CLK(clk), .RST(rst), .Q(xreg[465]) );
  DFF \xreg_reg[466]  ( .D(xin[465]), .CLK(clk), .RST(rst), .Q(xreg[466]) );
  DFF \xreg_reg[467]  ( .D(xin[466]), .CLK(clk), .RST(rst), .Q(xreg[467]) );
  DFF \xreg_reg[468]  ( .D(xin[467]), .CLK(clk), .RST(rst), .Q(xreg[468]) );
  DFF \xreg_reg[469]  ( .D(xin[468]), .CLK(clk), .RST(rst), .Q(xreg[469]) );
  DFF \xreg_reg[470]  ( .D(xin[469]), .CLK(clk), .RST(rst), .Q(xreg[470]) );
  DFF \xreg_reg[471]  ( .D(xin[470]), .CLK(clk), .RST(rst), .Q(xreg[471]) );
  DFF \xreg_reg[472]  ( .D(xin[471]), .CLK(clk), .RST(rst), .Q(xreg[472]) );
  DFF \xreg_reg[473]  ( .D(xin[472]), .CLK(clk), .RST(rst), .Q(xreg[473]) );
  DFF \xreg_reg[474]  ( .D(xin[473]), .CLK(clk), .RST(rst), .Q(xreg[474]) );
  DFF \xreg_reg[475]  ( .D(xin[474]), .CLK(clk), .RST(rst), .Q(xreg[475]) );
  DFF \xreg_reg[476]  ( .D(xin[475]), .CLK(clk), .RST(rst), .Q(xreg[476]) );
  DFF \xreg_reg[477]  ( .D(xin[476]), .CLK(clk), .RST(rst), .Q(xreg[477]) );
  DFF \xreg_reg[478]  ( .D(xin[477]), .CLK(clk), .RST(rst), .Q(xreg[478]) );
  DFF \xreg_reg[479]  ( .D(xin[478]), .CLK(clk), .RST(rst), .Q(xreg[479]) );
  DFF \xreg_reg[480]  ( .D(xin[479]), .CLK(clk), .RST(rst), .Q(xreg[480]) );
  DFF \xreg_reg[481]  ( .D(xin[480]), .CLK(clk), .RST(rst), .Q(xreg[481]) );
  DFF \xreg_reg[482]  ( .D(xin[481]), .CLK(clk), .RST(rst), .Q(xreg[482]) );
  DFF \xreg_reg[483]  ( .D(xin[482]), .CLK(clk), .RST(rst), .Q(xreg[483]) );
  DFF \xreg_reg[484]  ( .D(xin[483]), .CLK(clk), .RST(rst), .Q(xreg[484]) );
  DFF \xreg_reg[485]  ( .D(xin[484]), .CLK(clk), .RST(rst), .Q(xreg[485]) );
  DFF \xreg_reg[486]  ( .D(xin[485]), .CLK(clk), .RST(rst), .Q(xreg[486]) );
  DFF \xreg_reg[487]  ( .D(xin[486]), .CLK(clk), .RST(rst), .Q(xreg[487]) );
  DFF \xreg_reg[488]  ( .D(xin[487]), .CLK(clk), .RST(rst), .Q(xreg[488]) );
  DFF \xreg_reg[489]  ( .D(xin[488]), .CLK(clk), .RST(rst), .Q(xreg[489]) );
  DFF \xreg_reg[490]  ( .D(xin[489]), .CLK(clk), .RST(rst), .Q(xreg[490]) );
  DFF \xreg_reg[491]  ( .D(xin[490]), .CLK(clk), .RST(rst), .Q(xreg[491]) );
  DFF \xreg_reg[492]  ( .D(xin[491]), .CLK(clk), .RST(rst), .Q(xreg[492]) );
  DFF \xreg_reg[493]  ( .D(xin[492]), .CLK(clk), .RST(rst), .Q(xreg[493]) );
  DFF \xreg_reg[494]  ( .D(xin[493]), .CLK(clk), .RST(rst), .Q(xreg[494]) );
  DFF \xreg_reg[495]  ( .D(xin[494]), .CLK(clk), .RST(rst), .Q(xreg[495]) );
  DFF \xreg_reg[496]  ( .D(xin[495]), .CLK(clk), .RST(rst), .Q(xreg[496]) );
  DFF \xreg_reg[497]  ( .D(xin[496]), .CLK(clk), .RST(rst), .Q(xreg[497]) );
  DFF \xreg_reg[498]  ( .D(xin[497]), .CLK(clk), .RST(rst), .Q(xreg[498]) );
  DFF \xreg_reg[499]  ( .D(xin[498]), .CLK(clk), .RST(rst), .Q(xreg[499]) );
  DFF \xreg_reg[500]  ( .D(xin[499]), .CLK(clk), .RST(rst), .Q(xreg[500]) );
  DFF \xreg_reg[501]  ( .D(xin[500]), .CLK(clk), .RST(rst), .Q(xreg[501]) );
  DFF \xreg_reg[502]  ( .D(xin[501]), .CLK(clk), .RST(rst), .Q(xreg[502]) );
  DFF \xreg_reg[503]  ( .D(xin[502]), .CLK(clk), .RST(rst), .Q(xreg[503]) );
  DFF \xreg_reg[504]  ( .D(xin[503]), .CLK(clk), .RST(rst), .Q(xreg[504]) );
  DFF \xreg_reg[505]  ( .D(xin[504]), .CLK(clk), .RST(rst), .Q(xreg[505]) );
  DFF \xreg_reg[506]  ( .D(xin[505]), .CLK(clk), .RST(rst), .Q(xreg[506]) );
  DFF \xreg_reg[507]  ( .D(xin[506]), .CLK(clk), .RST(rst), .Q(xreg[507]) );
  DFF \xreg_reg[508]  ( .D(xin[507]), .CLK(clk), .RST(rst), .Q(xreg[508]) );
  DFF \xreg_reg[509]  ( .D(xin[508]), .CLK(clk), .RST(rst), .Q(xreg[509]) );
  DFF \xreg_reg[510]  ( .D(xin[509]), .CLK(clk), .RST(rst), .Q(xreg[510]) );
  DFF \xreg_reg[511]  ( .D(xin[510]), .CLK(clk), .RST(rst), .Q(xreg[511]) );
  DFF \zreg_reg[0]  ( .D(o[0]), .CLK(clk), .RST(rst), .Q(zreg[0]) );
  DFF \zreg_reg[1]  ( .D(o[1]), .CLK(clk), .RST(rst), .Q(zreg[1]) );
  DFF \zreg_reg[2]  ( .D(o[2]), .CLK(clk), .RST(rst), .Q(zreg[2]) );
  DFF \zreg_reg[3]  ( .D(o[3]), .CLK(clk), .RST(rst), .Q(zreg[3]) );
  DFF \zreg_reg[4]  ( .D(o[4]), .CLK(clk), .RST(rst), .Q(zreg[4]) );
  DFF \zreg_reg[5]  ( .D(o[5]), .CLK(clk), .RST(rst), .Q(zreg[5]) );
  DFF \zreg_reg[6]  ( .D(o[6]), .CLK(clk), .RST(rst), .Q(zreg[6]) );
  DFF \zreg_reg[7]  ( .D(o[7]), .CLK(clk), .RST(rst), .Q(zreg[7]) );
  DFF \zreg_reg[8]  ( .D(o[8]), .CLK(clk), .RST(rst), .Q(zreg[8]) );
  DFF \zreg_reg[9]  ( .D(o[9]), .CLK(clk), .RST(rst), .Q(zreg[9]) );
  DFF \zreg_reg[10]  ( .D(o[10]), .CLK(clk), .RST(rst), .Q(zreg[10]) );
  DFF \zreg_reg[11]  ( .D(o[11]), .CLK(clk), .RST(rst), .Q(zreg[11]) );
  DFF \zreg_reg[12]  ( .D(o[12]), .CLK(clk), .RST(rst), .Q(zreg[12]) );
  DFF \zreg_reg[13]  ( .D(o[13]), .CLK(clk), .RST(rst), .Q(zreg[13]) );
  DFF \zreg_reg[14]  ( .D(o[14]), .CLK(clk), .RST(rst), .Q(zreg[14]) );
  DFF \zreg_reg[15]  ( .D(o[15]), .CLK(clk), .RST(rst), .Q(zreg[15]) );
  DFF \zreg_reg[16]  ( .D(o[16]), .CLK(clk), .RST(rst), .Q(zreg[16]) );
  DFF \zreg_reg[17]  ( .D(o[17]), .CLK(clk), .RST(rst), .Q(zreg[17]) );
  DFF \zreg_reg[18]  ( .D(o[18]), .CLK(clk), .RST(rst), .Q(zreg[18]) );
  DFF \zreg_reg[19]  ( .D(o[19]), .CLK(clk), .RST(rst), .Q(zreg[19]) );
  DFF \zreg_reg[20]  ( .D(o[20]), .CLK(clk), .RST(rst), .Q(zreg[20]) );
  DFF \zreg_reg[21]  ( .D(o[21]), .CLK(clk), .RST(rst), .Q(zreg[21]) );
  DFF \zreg_reg[22]  ( .D(o[22]), .CLK(clk), .RST(rst), .Q(zreg[22]) );
  DFF \zreg_reg[23]  ( .D(o[23]), .CLK(clk), .RST(rst), .Q(zreg[23]) );
  DFF \zreg_reg[24]  ( .D(o[24]), .CLK(clk), .RST(rst), .Q(zreg[24]) );
  DFF \zreg_reg[25]  ( .D(o[25]), .CLK(clk), .RST(rst), .Q(zreg[25]) );
  DFF \zreg_reg[26]  ( .D(o[26]), .CLK(clk), .RST(rst), .Q(zreg[26]) );
  DFF \zreg_reg[27]  ( .D(o[27]), .CLK(clk), .RST(rst), .Q(zreg[27]) );
  DFF \zreg_reg[28]  ( .D(o[28]), .CLK(clk), .RST(rst), .Q(zreg[28]) );
  DFF \zreg_reg[29]  ( .D(o[29]), .CLK(clk), .RST(rst), .Q(zreg[29]) );
  DFF \zreg_reg[30]  ( .D(o[30]), .CLK(clk), .RST(rst), .Q(zreg[30]) );
  DFF \zreg_reg[31]  ( .D(o[31]), .CLK(clk), .RST(rst), .Q(zreg[31]) );
  DFF \zreg_reg[32]  ( .D(o[32]), .CLK(clk), .RST(rst), .Q(zreg[32]) );
  DFF \zreg_reg[33]  ( .D(o[33]), .CLK(clk), .RST(rst), .Q(zreg[33]) );
  DFF \zreg_reg[34]  ( .D(o[34]), .CLK(clk), .RST(rst), .Q(zreg[34]) );
  DFF \zreg_reg[35]  ( .D(o[35]), .CLK(clk), .RST(rst), .Q(zreg[35]) );
  DFF \zreg_reg[36]  ( .D(o[36]), .CLK(clk), .RST(rst), .Q(zreg[36]) );
  DFF \zreg_reg[37]  ( .D(o[37]), .CLK(clk), .RST(rst), .Q(zreg[37]) );
  DFF \zreg_reg[38]  ( .D(o[38]), .CLK(clk), .RST(rst), .Q(zreg[38]) );
  DFF \zreg_reg[39]  ( .D(o[39]), .CLK(clk), .RST(rst), .Q(zreg[39]) );
  DFF \zreg_reg[40]  ( .D(o[40]), .CLK(clk), .RST(rst), .Q(zreg[40]) );
  DFF \zreg_reg[41]  ( .D(o[41]), .CLK(clk), .RST(rst), .Q(zreg[41]) );
  DFF \zreg_reg[42]  ( .D(o[42]), .CLK(clk), .RST(rst), .Q(zreg[42]) );
  DFF \zreg_reg[43]  ( .D(o[43]), .CLK(clk), .RST(rst), .Q(zreg[43]) );
  DFF \zreg_reg[44]  ( .D(o[44]), .CLK(clk), .RST(rst), .Q(zreg[44]) );
  DFF \zreg_reg[45]  ( .D(o[45]), .CLK(clk), .RST(rst), .Q(zreg[45]) );
  DFF \zreg_reg[46]  ( .D(o[46]), .CLK(clk), .RST(rst), .Q(zreg[46]) );
  DFF \zreg_reg[47]  ( .D(o[47]), .CLK(clk), .RST(rst), .Q(zreg[47]) );
  DFF \zreg_reg[48]  ( .D(o[48]), .CLK(clk), .RST(rst), .Q(zreg[48]) );
  DFF \zreg_reg[49]  ( .D(o[49]), .CLK(clk), .RST(rst), .Q(zreg[49]) );
  DFF \zreg_reg[50]  ( .D(o[50]), .CLK(clk), .RST(rst), .Q(zreg[50]) );
  DFF \zreg_reg[51]  ( .D(o[51]), .CLK(clk), .RST(rst), .Q(zreg[51]) );
  DFF \zreg_reg[52]  ( .D(o[52]), .CLK(clk), .RST(rst), .Q(zreg[52]) );
  DFF \zreg_reg[53]  ( .D(o[53]), .CLK(clk), .RST(rst), .Q(zreg[53]) );
  DFF \zreg_reg[54]  ( .D(o[54]), .CLK(clk), .RST(rst), .Q(zreg[54]) );
  DFF \zreg_reg[55]  ( .D(o[55]), .CLK(clk), .RST(rst), .Q(zreg[55]) );
  DFF \zreg_reg[56]  ( .D(o[56]), .CLK(clk), .RST(rst), .Q(zreg[56]) );
  DFF \zreg_reg[57]  ( .D(o[57]), .CLK(clk), .RST(rst), .Q(zreg[57]) );
  DFF \zreg_reg[58]  ( .D(o[58]), .CLK(clk), .RST(rst), .Q(zreg[58]) );
  DFF \zreg_reg[59]  ( .D(o[59]), .CLK(clk), .RST(rst), .Q(zreg[59]) );
  DFF \zreg_reg[60]  ( .D(o[60]), .CLK(clk), .RST(rst), .Q(zreg[60]) );
  DFF \zreg_reg[61]  ( .D(o[61]), .CLK(clk), .RST(rst), .Q(zreg[61]) );
  DFF \zreg_reg[62]  ( .D(o[62]), .CLK(clk), .RST(rst), .Q(zreg[62]) );
  DFF \zreg_reg[63]  ( .D(o[63]), .CLK(clk), .RST(rst), .Q(zreg[63]) );
  DFF \zreg_reg[64]  ( .D(o[64]), .CLK(clk), .RST(rst), .Q(zreg[64]) );
  DFF \zreg_reg[65]  ( .D(o[65]), .CLK(clk), .RST(rst), .Q(zreg[65]) );
  DFF \zreg_reg[66]  ( .D(o[66]), .CLK(clk), .RST(rst), .Q(zreg[66]) );
  DFF \zreg_reg[67]  ( .D(o[67]), .CLK(clk), .RST(rst), .Q(zreg[67]) );
  DFF \zreg_reg[68]  ( .D(o[68]), .CLK(clk), .RST(rst), .Q(zreg[68]) );
  DFF \zreg_reg[69]  ( .D(o[69]), .CLK(clk), .RST(rst), .Q(zreg[69]) );
  DFF \zreg_reg[70]  ( .D(o[70]), .CLK(clk), .RST(rst), .Q(zreg[70]) );
  DFF \zreg_reg[71]  ( .D(o[71]), .CLK(clk), .RST(rst), .Q(zreg[71]) );
  DFF \zreg_reg[72]  ( .D(o[72]), .CLK(clk), .RST(rst), .Q(zreg[72]) );
  DFF \zreg_reg[73]  ( .D(o[73]), .CLK(clk), .RST(rst), .Q(zreg[73]) );
  DFF \zreg_reg[74]  ( .D(o[74]), .CLK(clk), .RST(rst), .Q(zreg[74]) );
  DFF \zreg_reg[75]  ( .D(o[75]), .CLK(clk), .RST(rst), .Q(zreg[75]) );
  DFF \zreg_reg[76]  ( .D(o[76]), .CLK(clk), .RST(rst), .Q(zreg[76]) );
  DFF \zreg_reg[77]  ( .D(o[77]), .CLK(clk), .RST(rst), .Q(zreg[77]) );
  DFF \zreg_reg[78]  ( .D(o[78]), .CLK(clk), .RST(rst), .Q(zreg[78]) );
  DFF \zreg_reg[79]  ( .D(o[79]), .CLK(clk), .RST(rst), .Q(zreg[79]) );
  DFF \zreg_reg[80]  ( .D(o[80]), .CLK(clk), .RST(rst), .Q(zreg[80]) );
  DFF \zreg_reg[81]  ( .D(o[81]), .CLK(clk), .RST(rst), .Q(zreg[81]) );
  DFF \zreg_reg[82]  ( .D(o[82]), .CLK(clk), .RST(rst), .Q(zreg[82]) );
  DFF \zreg_reg[83]  ( .D(o[83]), .CLK(clk), .RST(rst), .Q(zreg[83]) );
  DFF \zreg_reg[84]  ( .D(o[84]), .CLK(clk), .RST(rst), .Q(zreg[84]) );
  DFF \zreg_reg[85]  ( .D(o[85]), .CLK(clk), .RST(rst), .Q(zreg[85]) );
  DFF \zreg_reg[86]  ( .D(o[86]), .CLK(clk), .RST(rst), .Q(zreg[86]) );
  DFF \zreg_reg[87]  ( .D(o[87]), .CLK(clk), .RST(rst), .Q(zreg[87]) );
  DFF \zreg_reg[88]  ( .D(o[88]), .CLK(clk), .RST(rst), .Q(zreg[88]) );
  DFF \zreg_reg[89]  ( .D(o[89]), .CLK(clk), .RST(rst), .Q(zreg[89]) );
  DFF \zreg_reg[90]  ( .D(o[90]), .CLK(clk), .RST(rst), .Q(zreg[90]) );
  DFF \zreg_reg[91]  ( .D(o[91]), .CLK(clk), .RST(rst), .Q(zreg[91]) );
  DFF \zreg_reg[92]  ( .D(o[92]), .CLK(clk), .RST(rst), .Q(zreg[92]) );
  DFF \zreg_reg[93]  ( .D(o[93]), .CLK(clk), .RST(rst), .Q(zreg[93]) );
  DFF \zreg_reg[94]  ( .D(o[94]), .CLK(clk), .RST(rst), .Q(zreg[94]) );
  DFF \zreg_reg[95]  ( .D(o[95]), .CLK(clk), .RST(rst), .Q(zreg[95]) );
  DFF \zreg_reg[96]  ( .D(o[96]), .CLK(clk), .RST(rst), .Q(zreg[96]) );
  DFF \zreg_reg[97]  ( .D(o[97]), .CLK(clk), .RST(rst), .Q(zreg[97]) );
  DFF \zreg_reg[98]  ( .D(o[98]), .CLK(clk), .RST(rst), .Q(zreg[98]) );
  DFF \zreg_reg[99]  ( .D(o[99]), .CLK(clk), .RST(rst), .Q(zreg[99]) );
  DFF \zreg_reg[100]  ( .D(o[100]), .CLK(clk), .RST(rst), .Q(zreg[100]) );
  DFF \zreg_reg[101]  ( .D(o[101]), .CLK(clk), .RST(rst), .Q(zreg[101]) );
  DFF \zreg_reg[102]  ( .D(o[102]), .CLK(clk), .RST(rst), .Q(zreg[102]) );
  DFF \zreg_reg[103]  ( .D(o[103]), .CLK(clk), .RST(rst), .Q(zreg[103]) );
  DFF \zreg_reg[104]  ( .D(o[104]), .CLK(clk), .RST(rst), .Q(zreg[104]) );
  DFF \zreg_reg[105]  ( .D(o[105]), .CLK(clk), .RST(rst), .Q(zreg[105]) );
  DFF \zreg_reg[106]  ( .D(o[106]), .CLK(clk), .RST(rst), .Q(zreg[106]) );
  DFF \zreg_reg[107]  ( .D(o[107]), .CLK(clk), .RST(rst), .Q(zreg[107]) );
  DFF \zreg_reg[108]  ( .D(o[108]), .CLK(clk), .RST(rst), .Q(zreg[108]) );
  DFF \zreg_reg[109]  ( .D(o[109]), .CLK(clk), .RST(rst), .Q(zreg[109]) );
  DFF \zreg_reg[110]  ( .D(o[110]), .CLK(clk), .RST(rst), .Q(zreg[110]) );
  DFF \zreg_reg[111]  ( .D(o[111]), .CLK(clk), .RST(rst), .Q(zreg[111]) );
  DFF \zreg_reg[112]  ( .D(o[112]), .CLK(clk), .RST(rst), .Q(zreg[112]) );
  DFF \zreg_reg[113]  ( .D(o[113]), .CLK(clk), .RST(rst), .Q(zreg[113]) );
  DFF \zreg_reg[114]  ( .D(o[114]), .CLK(clk), .RST(rst), .Q(zreg[114]) );
  DFF \zreg_reg[115]  ( .D(o[115]), .CLK(clk), .RST(rst), .Q(zreg[115]) );
  DFF \zreg_reg[116]  ( .D(o[116]), .CLK(clk), .RST(rst), .Q(zreg[116]) );
  DFF \zreg_reg[117]  ( .D(o[117]), .CLK(clk), .RST(rst), .Q(zreg[117]) );
  DFF \zreg_reg[118]  ( .D(o[118]), .CLK(clk), .RST(rst), .Q(zreg[118]) );
  DFF \zreg_reg[119]  ( .D(o[119]), .CLK(clk), .RST(rst), .Q(zreg[119]) );
  DFF \zreg_reg[120]  ( .D(o[120]), .CLK(clk), .RST(rst), .Q(zreg[120]) );
  DFF \zreg_reg[121]  ( .D(o[121]), .CLK(clk), .RST(rst), .Q(zreg[121]) );
  DFF \zreg_reg[122]  ( .D(o[122]), .CLK(clk), .RST(rst), .Q(zreg[122]) );
  DFF \zreg_reg[123]  ( .D(o[123]), .CLK(clk), .RST(rst), .Q(zreg[123]) );
  DFF \zreg_reg[124]  ( .D(o[124]), .CLK(clk), .RST(rst), .Q(zreg[124]) );
  DFF \zreg_reg[125]  ( .D(o[125]), .CLK(clk), .RST(rst), .Q(zreg[125]) );
  DFF \zreg_reg[126]  ( .D(o[126]), .CLK(clk), .RST(rst), .Q(zreg[126]) );
  DFF \zreg_reg[127]  ( .D(o[127]), .CLK(clk), .RST(rst), .Q(zreg[127]) );
  DFF \zreg_reg[128]  ( .D(o[128]), .CLK(clk), .RST(rst), .Q(zreg[128]) );
  DFF \zreg_reg[129]  ( .D(o[129]), .CLK(clk), .RST(rst), .Q(zreg[129]) );
  DFF \zreg_reg[130]  ( .D(o[130]), .CLK(clk), .RST(rst), .Q(zreg[130]) );
  DFF \zreg_reg[131]  ( .D(o[131]), .CLK(clk), .RST(rst), .Q(zreg[131]) );
  DFF \zreg_reg[132]  ( .D(o[132]), .CLK(clk), .RST(rst), .Q(zreg[132]) );
  DFF \zreg_reg[133]  ( .D(o[133]), .CLK(clk), .RST(rst), .Q(zreg[133]) );
  DFF \zreg_reg[134]  ( .D(o[134]), .CLK(clk), .RST(rst), .Q(zreg[134]) );
  DFF \zreg_reg[135]  ( .D(o[135]), .CLK(clk), .RST(rst), .Q(zreg[135]) );
  DFF \zreg_reg[136]  ( .D(o[136]), .CLK(clk), .RST(rst), .Q(zreg[136]) );
  DFF \zreg_reg[137]  ( .D(o[137]), .CLK(clk), .RST(rst), .Q(zreg[137]) );
  DFF \zreg_reg[138]  ( .D(o[138]), .CLK(clk), .RST(rst), .Q(zreg[138]) );
  DFF \zreg_reg[139]  ( .D(o[139]), .CLK(clk), .RST(rst), .Q(zreg[139]) );
  DFF \zreg_reg[140]  ( .D(o[140]), .CLK(clk), .RST(rst), .Q(zreg[140]) );
  DFF \zreg_reg[141]  ( .D(o[141]), .CLK(clk), .RST(rst), .Q(zreg[141]) );
  DFF \zreg_reg[142]  ( .D(o[142]), .CLK(clk), .RST(rst), .Q(zreg[142]) );
  DFF \zreg_reg[143]  ( .D(o[143]), .CLK(clk), .RST(rst), .Q(zreg[143]) );
  DFF \zreg_reg[144]  ( .D(o[144]), .CLK(clk), .RST(rst), .Q(zreg[144]) );
  DFF \zreg_reg[145]  ( .D(o[145]), .CLK(clk), .RST(rst), .Q(zreg[145]) );
  DFF \zreg_reg[146]  ( .D(o[146]), .CLK(clk), .RST(rst), .Q(zreg[146]) );
  DFF \zreg_reg[147]  ( .D(o[147]), .CLK(clk), .RST(rst), .Q(zreg[147]) );
  DFF \zreg_reg[148]  ( .D(o[148]), .CLK(clk), .RST(rst), .Q(zreg[148]) );
  DFF \zreg_reg[149]  ( .D(o[149]), .CLK(clk), .RST(rst), .Q(zreg[149]) );
  DFF \zreg_reg[150]  ( .D(o[150]), .CLK(clk), .RST(rst), .Q(zreg[150]) );
  DFF \zreg_reg[151]  ( .D(o[151]), .CLK(clk), .RST(rst), .Q(zreg[151]) );
  DFF \zreg_reg[152]  ( .D(o[152]), .CLK(clk), .RST(rst), .Q(zreg[152]) );
  DFF \zreg_reg[153]  ( .D(o[153]), .CLK(clk), .RST(rst), .Q(zreg[153]) );
  DFF \zreg_reg[154]  ( .D(o[154]), .CLK(clk), .RST(rst), .Q(zreg[154]) );
  DFF \zreg_reg[155]  ( .D(o[155]), .CLK(clk), .RST(rst), .Q(zreg[155]) );
  DFF \zreg_reg[156]  ( .D(o[156]), .CLK(clk), .RST(rst), .Q(zreg[156]) );
  DFF \zreg_reg[157]  ( .D(o[157]), .CLK(clk), .RST(rst), .Q(zreg[157]) );
  DFF \zreg_reg[158]  ( .D(o[158]), .CLK(clk), .RST(rst), .Q(zreg[158]) );
  DFF \zreg_reg[159]  ( .D(o[159]), .CLK(clk), .RST(rst), .Q(zreg[159]) );
  DFF \zreg_reg[160]  ( .D(o[160]), .CLK(clk), .RST(rst), .Q(zreg[160]) );
  DFF \zreg_reg[161]  ( .D(o[161]), .CLK(clk), .RST(rst), .Q(zreg[161]) );
  DFF \zreg_reg[162]  ( .D(o[162]), .CLK(clk), .RST(rst), .Q(zreg[162]) );
  DFF \zreg_reg[163]  ( .D(o[163]), .CLK(clk), .RST(rst), .Q(zreg[163]) );
  DFF \zreg_reg[164]  ( .D(o[164]), .CLK(clk), .RST(rst), .Q(zreg[164]) );
  DFF \zreg_reg[165]  ( .D(o[165]), .CLK(clk), .RST(rst), .Q(zreg[165]) );
  DFF \zreg_reg[166]  ( .D(o[166]), .CLK(clk), .RST(rst), .Q(zreg[166]) );
  DFF \zreg_reg[167]  ( .D(o[167]), .CLK(clk), .RST(rst), .Q(zreg[167]) );
  DFF \zreg_reg[168]  ( .D(o[168]), .CLK(clk), .RST(rst), .Q(zreg[168]) );
  DFF \zreg_reg[169]  ( .D(o[169]), .CLK(clk), .RST(rst), .Q(zreg[169]) );
  DFF \zreg_reg[170]  ( .D(o[170]), .CLK(clk), .RST(rst), .Q(zreg[170]) );
  DFF \zreg_reg[171]  ( .D(o[171]), .CLK(clk), .RST(rst), .Q(zreg[171]) );
  DFF \zreg_reg[172]  ( .D(o[172]), .CLK(clk), .RST(rst), .Q(zreg[172]) );
  DFF \zreg_reg[173]  ( .D(o[173]), .CLK(clk), .RST(rst), .Q(zreg[173]) );
  DFF \zreg_reg[174]  ( .D(o[174]), .CLK(clk), .RST(rst), .Q(zreg[174]) );
  DFF \zreg_reg[175]  ( .D(o[175]), .CLK(clk), .RST(rst), .Q(zreg[175]) );
  DFF \zreg_reg[176]  ( .D(o[176]), .CLK(clk), .RST(rst), .Q(zreg[176]) );
  DFF \zreg_reg[177]  ( .D(o[177]), .CLK(clk), .RST(rst), .Q(zreg[177]) );
  DFF \zreg_reg[178]  ( .D(o[178]), .CLK(clk), .RST(rst), .Q(zreg[178]) );
  DFF \zreg_reg[179]  ( .D(o[179]), .CLK(clk), .RST(rst), .Q(zreg[179]) );
  DFF \zreg_reg[180]  ( .D(o[180]), .CLK(clk), .RST(rst), .Q(zreg[180]) );
  DFF \zreg_reg[181]  ( .D(o[181]), .CLK(clk), .RST(rst), .Q(zreg[181]) );
  DFF \zreg_reg[182]  ( .D(o[182]), .CLK(clk), .RST(rst), .Q(zreg[182]) );
  DFF \zreg_reg[183]  ( .D(o[183]), .CLK(clk), .RST(rst), .Q(zreg[183]) );
  DFF \zreg_reg[184]  ( .D(o[184]), .CLK(clk), .RST(rst), .Q(zreg[184]) );
  DFF \zreg_reg[185]  ( .D(o[185]), .CLK(clk), .RST(rst), .Q(zreg[185]) );
  DFF \zreg_reg[186]  ( .D(o[186]), .CLK(clk), .RST(rst), .Q(zreg[186]) );
  DFF \zreg_reg[187]  ( .D(o[187]), .CLK(clk), .RST(rst), .Q(zreg[187]) );
  DFF \zreg_reg[188]  ( .D(o[188]), .CLK(clk), .RST(rst), .Q(zreg[188]) );
  DFF \zreg_reg[189]  ( .D(o[189]), .CLK(clk), .RST(rst), .Q(zreg[189]) );
  DFF \zreg_reg[190]  ( .D(o[190]), .CLK(clk), .RST(rst), .Q(zreg[190]) );
  DFF \zreg_reg[191]  ( .D(o[191]), .CLK(clk), .RST(rst), .Q(zreg[191]) );
  DFF \zreg_reg[192]  ( .D(o[192]), .CLK(clk), .RST(rst), .Q(zreg[192]) );
  DFF \zreg_reg[193]  ( .D(o[193]), .CLK(clk), .RST(rst), .Q(zreg[193]) );
  DFF \zreg_reg[194]  ( .D(o[194]), .CLK(clk), .RST(rst), .Q(zreg[194]) );
  DFF \zreg_reg[195]  ( .D(o[195]), .CLK(clk), .RST(rst), .Q(zreg[195]) );
  DFF \zreg_reg[196]  ( .D(o[196]), .CLK(clk), .RST(rst), .Q(zreg[196]) );
  DFF \zreg_reg[197]  ( .D(o[197]), .CLK(clk), .RST(rst), .Q(zreg[197]) );
  DFF \zreg_reg[198]  ( .D(o[198]), .CLK(clk), .RST(rst), .Q(zreg[198]) );
  DFF \zreg_reg[199]  ( .D(o[199]), .CLK(clk), .RST(rst), .Q(zreg[199]) );
  DFF \zreg_reg[200]  ( .D(o[200]), .CLK(clk), .RST(rst), .Q(zreg[200]) );
  DFF \zreg_reg[201]  ( .D(o[201]), .CLK(clk), .RST(rst), .Q(zreg[201]) );
  DFF \zreg_reg[202]  ( .D(o[202]), .CLK(clk), .RST(rst), .Q(zreg[202]) );
  DFF \zreg_reg[203]  ( .D(o[203]), .CLK(clk), .RST(rst), .Q(zreg[203]) );
  DFF \zreg_reg[204]  ( .D(o[204]), .CLK(clk), .RST(rst), .Q(zreg[204]) );
  DFF \zreg_reg[205]  ( .D(o[205]), .CLK(clk), .RST(rst), .Q(zreg[205]) );
  DFF \zreg_reg[206]  ( .D(o[206]), .CLK(clk), .RST(rst), .Q(zreg[206]) );
  DFF \zreg_reg[207]  ( .D(o[207]), .CLK(clk), .RST(rst), .Q(zreg[207]) );
  DFF \zreg_reg[208]  ( .D(o[208]), .CLK(clk), .RST(rst), .Q(zreg[208]) );
  DFF \zreg_reg[209]  ( .D(o[209]), .CLK(clk), .RST(rst), .Q(zreg[209]) );
  DFF \zreg_reg[210]  ( .D(o[210]), .CLK(clk), .RST(rst), .Q(zreg[210]) );
  DFF \zreg_reg[211]  ( .D(o[211]), .CLK(clk), .RST(rst), .Q(zreg[211]) );
  DFF \zreg_reg[212]  ( .D(o[212]), .CLK(clk), .RST(rst), .Q(zreg[212]) );
  DFF \zreg_reg[213]  ( .D(o[213]), .CLK(clk), .RST(rst), .Q(zreg[213]) );
  DFF \zreg_reg[214]  ( .D(o[214]), .CLK(clk), .RST(rst), .Q(zreg[214]) );
  DFF \zreg_reg[215]  ( .D(o[215]), .CLK(clk), .RST(rst), .Q(zreg[215]) );
  DFF \zreg_reg[216]  ( .D(o[216]), .CLK(clk), .RST(rst), .Q(zreg[216]) );
  DFF \zreg_reg[217]  ( .D(o[217]), .CLK(clk), .RST(rst), .Q(zreg[217]) );
  DFF \zreg_reg[218]  ( .D(o[218]), .CLK(clk), .RST(rst), .Q(zreg[218]) );
  DFF \zreg_reg[219]  ( .D(o[219]), .CLK(clk), .RST(rst), .Q(zreg[219]) );
  DFF \zreg_reg[220]  ( .D(o[220]), .CLK(clk), .RST(rst), .Q(zreg[220]) );
  DFF \zreg_reg[221]  ( .D(o[221]), .CLK(clk), .RST(rst), .Q(zreg[221]) );
  DFF \zreg_reg[222]  ( .D(o[222]), .CLK(clk), .RST(rst), .Q(zreg[222]) );
  DFF \zreg_reg[223]  ( .D(o[223]), .CLK(clk), .RST(rst), .Q(zreg[223]) );
  DFF \zreg_reg[224]  ( .D(o[224]), .CLK(clk), .RST(rst), .Q(zreg[224]) );
  DFF \zreg_reg[225]  ( .D(o[225]), .CLK(clk), .RST(rst), .Q(zreg[225]) );
  DFF \zreg_reg[226]  ( .D(o[226]), .CLK(clk), .RST(rst), .Q(zreg[226]) );
  DFF \zreg_reg[227]  ( .D(o[227]), .CLK(clk), .RST(rst), .Q(zreg[227]) );
  DFF \zreg_reg[228]  ( .D(o[228]), .CLK(clk), .RST(rst), .Q(zreg[228]) );
  DFF \zreg_reg[229]  ( .D(o[229]), .CLK(clk), .RST(rst), .Q(zreg[229]) );
  DFF \zreg_reg[230]  ( .D(o[230]), .CLK(clk), .RST(rst), .Q(zreg[230]) );
  DFF \zreg_reg[231]  ( .D(o[231]), .CLK(clk), .RST(rst), .Q(zreg[231]) );
  DFF \zreg_reg[232]  ( .D(o[232]), .CLK(clk), .RST(rst), .Q(zreg[232]) );
  DFF \zreg_reg[233]  ( .D(o[233]), .CLK(clk), .RST(rst), .Q(zreg[233]) );
  DFF \zreg_reg[234]  ( .D(o[234]), .CLK(clk), .RST(rst), .Q(zreg[234]) );
  DFF \zreg_reg[235]  ( .D(o[235]), .CLK(clk), .RST(rst), .Q(zreg[235]) );
  DFF \zreg_reg[236]  ( .D(o[236]), .CLK(clk), .RST(rst), .Q(zreg[236]) );
  DFF \zreg_reg[237]  ( .D(o[237]), .CLK(clk), .RST(rst), .Q(zreg[237]) );
  DFF \zreg_reg[238]  ( .D(o[238]), .CLK(clk), .RST(rst), .Q(zreg[238]) );
  DFF \zreg_reg[239]  ( .D(o[239]), .CLK(clk), .RST(rst), .Q(zreg[239]) );
  DFF \zreg_reg[240]  ( .D(o[240]), .CLK(clk), .RST(rst), .Q(zreg[240]) );
  DFF \zreg_reg[241]  ( .D(o[241]), .CLK(clk), .RST(rst), .Q(zreg[241]) );
  DFF \zreg_reg[242]  ( .D(o[242]), .CLK(clk), .RST(rst), .Q(zreg[242]) );
  DFF \zreg_reg[243]  ( .D(o[243]), .CLK(clk), .RST(rst), .Q(zreg[243]) );
  DFF \zreg_reg[244]  ( .D(o[244]), .CLK(clk), .RST(rst), .Q(zreg[244]) );
  DFF \zreg_reg[245]  ( .D(o[245]), .CLK(clk), .RST(rst), .Q(zreg[245]) );
  DFF \zreg_reg[246]  ( .D(o[246]), .CLK(clk), .RST(rst), .Q(zreg[246]) );
  DFF \zreg_reg[247]  ( .D(o[247]), .CLK(clk), .RST(rst), .Q(zreg[247]) );
  DFF \zreg_reg[248]  ( .D(o[248]), .CLK(clk), .RST(rst), .Q(zreg[248]) );
  DFF \zreg_reg[249]  ( .D(o[249]), .CLK(clk), .RST(rst), .Q(zreg[249]) );
  DFF \zreg_reg[250]  ( .D(o[250]), .CLK(clk), .RST(rst), .Q(zreg[250]) );
  DFF \zreg_reg[251]  ( .D(o[251]), .CLK(clk), .RST(rst), .Q(zreg[251]) );
  DFF \zreg_reg[252]  ( .D(o[252]), .CLK(clk), .RST(rst), .Q(zreg[252]) );
  DFF \zreg_reg[253]  ( .D(o[253]), .CLK(clk), .RST(rst), .Q(zreg[253]) );
  DFF \zreg_reg[254]  ( .D(o[254]), .CLK(clk), .RST(rst), .Q(zreg[254]) );
  DFF \zreg_reg[255]  ( .D(o[255]), .CLK(clk), .RST(rst), .Q(zreg[255]) );
  DFF \zreg_reg[256]  ( .D(o[256]), .CLK(clk), .RST(rst), .Q(zreg[256]) );
  DFF \zreg_reg[257]  ( .D(o[257]), .CLK(clk), .RST(rst), .Q(zreg[257]) );
  DFF \zreg_reg[258]  ( .D(o[258]), .CLK(clk), .RST(rst), .Q(zreg[258]) );
  DFF \zreg_reg[259]  ( .D(o[259]), .CLK(clk), .RST(rst), .Q(zreg[259]) );
  DFF \zreg_reg[260]  ( .D(o[260]), .CLK(clk), .RST(rst), .Q(zreg[260]) );
  DFF \zreg_reg[261]  ( .D(o[261]), .CLK(clk), .RST(rst), .Q(zreg[261]) );
  DFF \zreg_reg[262]  ( .D(o[262]), .CLK(clk), .RST(rst), .Q(zreg[262]) );
  DFF \zreg_reg[263]  ( .D(o[263]), .CLK(clk), .RST(rst), .Q(zreg[263]) );
  DFF \zreg_reg[264]  ( .D(o[264]), .CLK(clk), .RST(rst), .Q(zreg[264]) );
  DFF \zreg_reg[265]  ( .D(o[265]), .CLK(clk), .RST(rst), .Q(zreg[265]) );
  DFF \zreg_reg[266]  ( .D(o[266]), .CLK(clk), .RST(rst), .Q(zreg[266]) );
  DFF \zreg_reg[267]  ( .D(o[267]), .CLK(clk), .RST(rst), .Q(zreg[267]) );
  DFF \zreg_reg[268]  ( .D(o[268]), .CLK(clk), .RST(rst), .Q(zreg[268]) );
  DFF \zreg_reg[269]  ( .D(o[269]), .CLK(clk), .RST(rst), .Q(zreg[269]) );
  DFF \zreg_reg[270]  ( .D(o[270]), .CLK(clk), .RST(rst), .Q(zreg[270]) );
  DFF \zreg_reg[271]  ( .D(o[271]), .CLK(clk), .RST(rst), .Q(zreg[271]) );
  DFF \zreg_reg[272]  ( .D(o[272]), .CLK(clk), .RST(rst), .Q(zreg[272]) );
  DFF \zreg_reg[273]  ( .D(o[273]), .CLK(clk), .RST(rst), .Q(zreg[273]) );
  DFF \zreg_reg[274]  ( .D(o[274]), .CLK(clk), .RST(rst), .Q(zreg[274]) );
  DFF \zreg_reg[275]  ( .D(o[275]), .CLK(clk), .RST(rst), .Q(zreg[275]) );
  DFF \zreg_reg[276]  ( .D(o[276]), .CLK(clk), .RST(rst), .Q(zreg[276]) );
  DFF \zreg_reg[277]  ( .D(o[277]), .CLK(clk), .RST(rst), .Q(zreg[277]) );
  DFF \zreg_reg[278]  ( .D(o[278]), .CLK(clk), .RST(rst), .Q(zreg[278]) );
  DFF \zreg_reg[279]  ( .D(o[279]), .CLK(clk), .RST(rst), .Q(zreg[279]) );
  DFF \zreg_reg[280]  ( .D(o[280]), .CLK(clk), .RST(rst), .Q(zreg[280]) );
  DFF \zreg_reg[281]  ( .D(o[281]), .CLK(clk), .RST(rst), .Q(zreg[281]) );
  DFF \zreg_reg[282]  ( .D(o[282]), .CLK(clk), .RST(rst), .Q(zreg[282]) );
  DFF \zreg_reg[283]  ( .D(o[283]), .CLK(clk), .RST(rst), .Q(zreg[283]) );
  DFF \zreg_reg[284]  ( .D(o[284]), .CLK(clk), .RST(rst), .Q(zreg[284]) );
  DFF \zreg_reg[285]  ( .D(o[285]), .CLK(clk), .RST(rst), .Q(zreg[285]) );
  DFF \zreg_reg[286]  ( .D(o[286]), .CLK(clk), .RST(rst), .Q(zreg[286]) );
  DFF \zreg_reg[287]  ( .D(o[287]), .CLK(clk), .RST(rst), .Q(zreg[287]) );
  DFF \zreg_reg[288]  ( .D(o[288]), .CLK(clk), .RST(rst), .Q(zreg[288]) );
  DFF \zreg_reg[289]  ( .D(o[289]), .CLK(clk), .RST(rst), .Q(zreg[289]) );
  DFF \zreg_reg[290]  ( .D(o[290]), .CLK(clk), .RST(rst), .Q(zreg[290]) );
  DFF \zreg_reg[291]  ( .D(o[291]), .CLK(clk), .RST(rst), .Q(zreg[291]) );
  DFF \zreg_reg[292]  ( .D(o[292]), .CLK(clk), .RST(rst), .Q(zreg[292]) );
  DFF \zreg_reg[293]  ( .D(o[293]), .CLK(clk), .RST(rst), .Q(zreg[293]) );
  DFF \zreg_reg[294]  ( .D(o[294]), .CLK(clk), .RST(rst), .Q(zreg[294]) );
  DFF \zreg_reg[295]  ( .D(o[295]), .CLK(clk), .RST(rst), .Q(zreg[295]) );
  DFF \zreg_reg[296]  ( .D(o[296]), .CLK(clk), .RST(rst), .Q(zreg[296]) );
  DFF \zreg_reg[297]  ( .D(o[297]), .CLK(clk), .RST(rst), .Q(zreg[297]) );
  DFF \zreg_reg[298]  ( .D(o[298]), .CLK(clk), .RST(rst), .Q(zreg[298]) );
  DFF \zreg_reg[299]  ( .D(o[299]), .CLK(clk), .RST(rst), .Q(zreg[299]) );
  DFF \zreg_reg[300]  ( .D(o[300]), .CLK(clk), .RST(rst), .Q(zreg[300]) );
  DFF \zreg_reg[301]  ( .D(o[301]), .CLK(clk), .RST(rst), .Q(zreg[301]) );
  DFF \zreg_reg[302]  ( .D(o[302]), .CLK(clk), .RST(rst), .Q(zreg[302]) );
  DFF \zreg_reg[303]  ( .D(o[303]), .CLK(clk), .RST(rst), .Q(zreg[303]) );
  DFF \zreg_reg[304]  ( .D(o[304]), .CLK(clk), .RST(rst), .Q(zreg[304]) );
  DFF \zreg_reg[305]  ( .D(o[305]), .CLK(clk), .RST(rst), .Q(zreg[305]) );
  DFF \zreg_reg[306]  ( .D(o[306]), .CLK(clk), .RST(rst), .Q(zreg[306]) );
  DFF \zreg_reg[307]  ( .D(o[307]), .CLK(clk), .RST(rst), .Q(zreg[307]) );
  DFF \zreg_reg[308]  ( .D(o[308]), .CLK(clk), .RST(rst), .Q(zreg[308]) );
  DFF \zreg_reg[309]  ( .D(o[309]), .CLK(clk), .RST(rst), .Q(zreg[309]) );
  DFF \zreg_reg[310]  ( .D(o[310]), .CLK(clk), .RST(rst), .Q(zreg[310]) );
  DFF \zreg_reg[311]  ( .D(o[311]), .CLK(clk), .RST(rst), .Q(zreg[311]) );
  DFF \zreg_reg[312]  ( .D(o[312]), .CLK(clk), .RST(rst), .Q(zreg[312]) );
  DFF \zreg_reg[313]  ( .D(o[313]), .CLK(clk), .RST(rst), .Q(zreg[313]) );
  DFF \zreg_reg[314]  ( .D(o[314]), .CLK(clk), .RST(rst), .Q(zreg[314]) );
  DFF \zreg_reg[315]  ( .D(o[315]), .CLK(clk), .RST(rst), .Q(zreg[315]) );
  DFF \zreg_reg[316]  ( .D(o[316]), .CLK(clk), .RST(rst), .Q(zreg[316]) );
  DFF \zreg_reg[317]  ( .D(o[317]), .CLK(clk), .RST(rst), .Q(zreg[317]) );
  DFF \zreg_reg[318]  ( .D(o[318]), .CLK(clk), .RST(rst), .Q(zreg[318]) );
  DFF \zreg_reg[319]  ( .D(o[319]), .CLK(clk), .RST(rst), .Q(zreg[319]) );
  DFF \zreg_reg[320]  ( .D(o[320]), .CLK(clk), .RST(rst), .Q(zreg[320]) );
  DFF \zreg_reg[321]  ( .D(o[321]), .CLK(clk), .RST(rst), .Q(zreg[321]) );
  DFF \zreg_reg[322]  ( .D(o[322]), .CLK(clk), .RST(rst), .Q(zreg[322]) );
  DFF \zreg_reg[323]  ( .D(o[323]), .CLK(clk), .RST(rst), .Q(zreg[323]) );
  DFF \zreg_reg[324]  ( .D(o[324]), .CLK(clk), .RST(rst), .Q(zreg[324]) );
  DFF \zreg_reg[325]  ( .D(o[325]), .CLK(clk), .RST(rst), .Q(zreg[325]) );
  DFF \zreg_reg[326]  ( .D(o[326]), .CLK(clk), .RST(rst), .Q(zreg[326]) );
  DFF \zreg_reg[327]  ( .D(o[327]), .CLK(clk), .RST(rst), .Q(zreg[327]) );
  DFF \zreg_reg[328]  ( .D(o[328]), .CLK(clk), .RST(rst), .Q(zreg[328]) );
  DFF \zreg_reg[329]  ( .D(o[329]), .CLK(clk), .RST(rst), .Q(zreg[329]) );
  DFF \zreg_reg[330]  ( .D(o[330]), .CLK(clk), .RST(rst), .Q(zreg[330]) );
  DFF \zreg_reg[331]  ( .D(o[331]), .CLK(clk), .RST(rst), .Q(zreg[331]) );
  DFF \zreg_reg[332]  ( .D(o[332]), .CLK(clk), .RST(rst), .Q(zreg[332]) );
  DFF \zreg_reg[333]  ( .D(o[333]), .CLK(clk), .RST(rst), .Q(zreg[333]) );
  DFF \zreg_reg[334]  ( .D(o[334]), .CLK(clk), .RST(rst), .Q(zreg[334]) );
  DFF \zreg_reg[335]  ( .D(o[335]), .CLK(clk), .RST(rst), .Q(zreg[335]) );
  DFF \zreg_reg[336]  ( .D(o[336]), .CLK(clk), .RST(rst), .Q(zreg[336]) );
  DFF \zreg_reg[337]  ( .D(o[337]), .CLK(clk), .RST(rst), .Q(zreg[337]) );
  DFF \zreg_reg[338]  ( .D(o[338]), .CLK(clk), .RST(rst), .Q(zreg[338]) );
  DFF \zreg_reg[339]  ( .D(o[339]), .CLK(clk), .RST(rst), .Q(zreg[339]) );
  DFF \zreg_reg[340]  ( .D(o[340]), .CLK(clk), .RST(rst), .Q(zreg[340]) );
  DFF \zreg_reg[341]  ( .D(o[341]), .CLK(clk), .RST(rst), .Q(zreg[341]) );
  DFF \zreg_reg[342]  ( .D(o[342]), .CLK(clk), .RST(rst), .Q(zreg[342]) );
  DFF \zreg_reg[343]  ( .D(o[343]), .CLK(clk), .RST(rst), .Q(zreg[343]) );
  DFF \zreg_reg[344]  ( .D(o[344]), .CLK(clk), .RST(rst), .Q(zreg[344]) );
  DFF \zreg_reg[345]  ( .D(o[345]), .CLK(clk), .RST(rst), .Q(zreg[345]) );
  DFF \zreg_reg[346]  ( .D(o[346]), .CLK(clk), .RST(rst), .Q(zreg[346]) );
  DFF \zreg_reg[347]  ( .D(o[347]), .CLK(clk), .RST(rst), .Q(zreg[347]) );
  DFF \zreg_reg[348]  ( .D(o[348]), .CLK(clk), .RST(rst), .Q(zreg[348]) );
  DFF \zreg_reg[349]  ( .D(o[349]), .CLK(clk), .RST(rst), .Q(zreg[349]) );
  DFF \zreg_reg[350]  ( .D(o[350]), .CLK(clk), .RST(rst), .Q(zreg[350]) );
  DFF \zreg_reg[351]  ( .D(o[351]), .CLK(clk), .RST(rst), .Q(zreg[351]) );
  DFF \zreg_reg[352]  ( .D(o[352]), .CLK(clk), .RST(rst), .Q(zreg[352]) );
  DFF \zreg_reg[353]  ( .D(o[353]), .CLK(clk), .RST(rst), .Q(zreg[353]) );
  DFF \zreg_reg[354]  ( .D(o[354]), .CLK(clk), .RST(rst), .Q(zreg[354]) );
  DFF \zreg_reg[355]  ( .D(o[355]), .CLK(clk), .RST(rst), .Q(zreg[355]) );
  DFF \zreg_reg[356]  ( .D(o[356]), .CLK(clk), .RST(rst), .Q(zreg[356]) );
  DFF \zreg_reg[357]  ( .D(o[357]), .CLK(clk), .RST(rst), .Q(zreg[357]) );
  DFF \zreg_reg[358]  ( .D(o[358]), .CLK(clk), .RST(rst), .Q(zreg[358]) );
  DFF \zreg_reg[359]  ( .D(o[359]), .CLK(clk), .RST(rst), .Q(zreg[359]) );
  DFF \zreg_reg[360]  ( .D(o[360]), .CLK(clk), .RST(rst), .Q(zreg[360]) );
  DFF \zreg_reg[361]  ( .D(o[361]), .CLK(clk), .RST(rst), .Q(zreg[361]) );
  DFF \zreg_reg[362]  ( .D(o[362]), .CLK(clk), .RST(rst), .Q(zreg[362]) );
  DFF \zreg_reg[363]  ( .D(o[363]), .CLK(clk), .RST(rst), .Q(zreg[363]) );
  DFF \zreg_reg[364]  ( .D(o[364]), .CLK(clk), .RST(rst), .Q(zreg[364]) );
  DFF \zreg_reg[365]  ( .D(o[365]), .CLK(clk), .RST(rst), .Q(zreg[365]) );
  DFF \zreg_reg[366]  ( .D(o[366]), .CLK(clk), .RST(rst), .Q(zreg[366]) );
  DFF \zreg_reg[367]  ( .D(o[367]), .CLK(clk), .RST(rst), .Q(zreg[367]) );
  DFF \zreg_reg[368]  ( .D(o[368]), .CLK(clk), .RST(rst), .Q(zreg[368]) );
  DFF \zreg_reg[369]  ( .D(o[369]), .CLK(clk), .RST(rst), .Q(zreg[369]) );
  DFF \zreg_reg[370]  ( .D(o[370]), .CLK(clk), .RST(rst), .Q(zreg[370]) );
  DFF \zreg_reg[371]  ( .D(o[371]), .CLK(clk), .RST(rst), .Q(zreg[371]) );
  DFF \zreg_reg[372]  ( .D(o[372]), .CLK(clk), .RST(rst), .Q(zreg[372]) );
  DFF \zreg_reg[373]  ( .D(o[373]), .CLK(clk), .RST(rst), .Q(zreg[373]) );
  DFF \zreg_reg[374]  ( .D(o[374]), .CLK(clk), .RST(rst), .Q(zreg[374]) );
  DFF \zreg_reg[375]  ( .D(o[375]), .CLK(clk), .RST(rst), .Q(zreg[375]) );
  DFF \zreg_reg[376]  ( .D(o[376]), .CLK(clk), .RST(rst), .Q(zreg[376]) );
  DFF \zreg_reg[377]  ( .D(o[377]), .CLK(clk), .RST(rst), .Q(zreg[377]) );
  DFF \zreg_reg[378]  ( .D(o[378]), .CLK(clk), .RST(rst), .Q(zreg[378]) );
  DFF \zreg_reg[379]  ( .D(o[379]), .CLK(clk), .RST(rst), .Q(zreg[379]) );
  DFF \zreg_reg[380]  ( .D(o[380]), .CLK(clk), .RST(rst), .Q(zreg[380]) );
  DFF \zreg_reg[381]  ( .D(o[381]), .CLK(clk), .RST(rst), .Q(zreg[381]) );
  DFF \zreg_reg[382]  ( .D(o[382]), .CLK(clk), .RST(rst), .Q(zreg[382]) );
  DFF \zreg_reg[383]  ( .D(o[383]), .CLK(clk), .RST(rst), .Q(zreg[383]) );
  DFF \zreg_reg[384]  ( .D(o[384]), .CLK(clk), .RST(rst), .Q(zreg[384]) );
  DFF \zreg_reg[385]  ( .D(o[385]), .CLK(clk), .RST(rst), .Q(zreg[385]) );
  DFF \zreg_reg[386]  ( .D(o[386]), .CLK(clk), .RST(rst), .Q(zreg[386]) );
  DFF \zreg_reg[387]  ( .D(o[387]), .CLK(clk), .RST(rst), .Q(zreg[387]) );
  DFF \zreg_reg[388]  ( .D(o[388]), .CLK(clk), .RST(rst), .Q(zreg[388]) );
  DFF \zreg_reg[389]  ( .D(o[389]), .CLK(clk), .RST(rst), .Q(zreg[389]) );
  DFF \zreg_reg[390]  ( .D(o[390]), .CLK(clk), .RST(rst), .Q(zreg[390]) );
  DFF \zreg_reg[391]  ( .D(o[391]), .CLK(clk), .RST(rst), .Q(zreg[391]) );
  DFF \zreg_reg[392]  ( .D(o[392]), .CLK(clk), .RST(rst), .Q(zreg[392]) );
  DFF \zreg_reg[393]  ( .D(o[393]), .CLK(clk), .RST(rst), .Q(zreg[393]) );
  DFF \zreg_reg[394]  ( .D(o[394]), .CLK(clk), .RST(rst), .Q(zreg[394]) );
  DFF \zreg_reg[395]  ( .D(o[395]), .CLK(clk), .RST(rst), .Q(zreg[395]) );
  DFF \zreg_reg[396]  ( .D(o[396]), .CLK(clk), .RST(rst), .Q(zreg[396]) );
  DFF \zreg_reg[397]  ( .D(o[397]), .CLK(clk), .RST(rst), .Q(zreg[397]) );
  DFF \zreg_reg[398]  ( .D(o[398]), .CLK(clk), .RST(rst), .Q(zreg[398]) );
  DFF \zreg_reg[399]  ( .D(o[399]), .CLK(clk), .RST(rst), .Q(zreg[399]) );
  DFF \zreg_reg[400]  ( .D(o[400]), .CLK(clk), .RST(rst), .Q(zreg[400]) );
  DFF \zreg_reg[401]  ( .D(o[401]), .CLK(clk), .RST(rst), .Q(zreg[401]) );
  DFF \zreg_reg[402]  ( .D(o[402]), .CLK(clk), .RST(rst), .Q(zreg[402]) );
  DFF \zreg_reg[403]  ( .D(o[403]), .CLK(clk), .RST(rst), .Q(zreg[403]) );
  DFF \zreg_reg[404]  ( .D(o[404]), .CLK(clk), .RST(rst), .Q(zreg[404]) );
  DFF \zreg_reg[405]  ( .D(o[405]), .CLK(clk), .RST(rst), .Q(zreg[405]) );
  DFF \zreg_reg[406]  ( .D(o[406]), .CLK(clk), .RST(rst), .Q(zreg[406]) );
  DFF \zreg_reg[407]  ( .D(o[407]), .CLK(clk), .RST(rst), .Q(zreg[407]) );
  DFF \zreg_reg[408]  ( .D(o[408]), .CLK(clk), .RST(rst), .Q(zreg[408]) );
  DFF \zreg_reg[409]  ( .D(o[409]), .CLK(clk), .RST(rst), .Q(zreg[409]) );
  DFF \zreg_reg[410]  ( .D(o[410]), .CLK(clk), .RST(rst), .Q(zreg[410]) );
  DFF \zreg_reg[411]  ( .D(o[411]), .CLK(clk), .RST(rst), .Q(zreg[411]) );
  DFF \zreg_reg[412]  ( .D(o[412]), .CLK(clk), .RST(rst), .Q(zreg[412]) );
  DFF \zreg_reg[413]  ( .D(o[413]), .CLK(clk), .RST(rst), .Q(zreg[413]) );
  DFF \zreg_reg[414]  ( .D(o[414]), .CLK(clk), .RST(rst), .Q(zreg[414]) );
  DFF \zreg_reg[415]  ( .D(o[415]), .CLK(clk), .RST(rst), .Q(zreg[415]) );
  DFF \zreg_reg[416]  ( .D(o[416]), .CLK(clk), .RST(rst), .Q(zreg[416]) );
  DFF \zreg_reg[417]  ( .D(o[417]), .CLK(clk), .RST(rst), .Q(zreg[417]) );
  DFF \zreg_reg[418]  ( .D(o[418]), .CLK(clk), .RST(rst), .Q(zreg[418]) );
  DFF \zreg_reg[419]  ( .D(o[419]), .CLK(clk), .RST(rst), .Q(zreg[419]) );
  DFF \zreg_reg[420]  ( .D(o[420]), .CLK(clk), .RST(rst), .Q(zreg[420]) );
  DFF \zreg_reg[421]  ( .D(o[421]), .CLK(clk), .RST(rst), .Q(zreg[421]) );
  DFF \zreg_reg[422]  ( .D(o[422]), .CLK(clk), .RST(rst), .Q(zreg[422]) );
  DFF \zreg_reg[423]  ( .D(o[423]), .CLK(clk), .RST(rst), .Q(zreg[423]) );
  DFF \zreg_reg[424]  ( .D(o[424]), .CLK(clk), .RST(rst), .Q(zreg[424]) );
  DFF \zreg_reg[425]  ( .D(o[425]), .CLK(clk), .RST(rst), .Q(zreg[425]) );
  DFF \zreg_reg[426]  ( .D(o[426]), .CLK(clk), .RST(rst), .Q(zreg[426]) );
  DFF \zreg_reg[427]  ( .D(o[427]), .CLK(clk), .RST(rst), .Q(zreg[427]) );
  DFF \zreg_reg[428]  ( .D(o[428]), .CLK(clk), .RST(rst), .Q(zreg[428]) );
  DFF \zreg_reg[429]  ( .D(o[429]), .CLK(clk), .RST(rst), .Q(zreg[429]) );
  DFF \zreg_reg[430]  ( .D(o[430]), .CLK(clk), .RST(rst), .Q(zreg[430]) );
  DFF \zreg_reg[431]  ( .D(o[431]), .CLK(clk), .RST(rst), .Q(zreg[431]) );
  DFF \zreg_reg[432]  ( .D(o[432]), .CLK(clk), .RST(rst), .Q(zreg[432]) );
  DFF \zreg_reg[433]  ( .D(o[433]), .CLK(clk), .RST(rst), .Q(zreg[433]) );
  DFF \zreg_reg[434]  ( .D(o[434]), .CLK(clk), .RST(rst), .Q(zreg[434]) );
  DFF \zreg_reg[435]  ( .D(o[435]), .CLK(clk), .RST(rst), .Q(zreg[435]) );
  DFF \zreg_reg[436]  ( .D(o[436]), .CLK(clk), .RST(rst), .Q(zreg[436]) );
  DFF \zreg_reg[437]  ( .D(o[437]), .CLK(clk), .RST(rst), .Q(zreg[437]) );
  DFF \zreg_reg[438]  ( .D(o[438]), .CLK(clk), .RST(rst), .Q(zreg[438]) );
  DFF \zreg_reg[439]  ( .D(o[439]), .CLK(clk), .RST(rst), .Q(zreg[439]) );
  DFF \zreg_reg[440]  ( .D(o[440]), .CLK(clk), .RST(rst), .Q(zreg[440]) );
  DFF \zreg_reg[441]  ( .D(o[441]), .CLK(clk), .RST(rst), .Q(zreg[441]) );
  DFF \zreg_reg[442]  ( .D(o[442]), .CLK(clk), .RST(rst), .Q(zreg[442]) );
  DFF \zreg_reg[443]  ( .D(o[443]), .CLK(clk), .RST(rst), .Q(zreg[443]) );
  DFF \zreg_reg[444]  ( .D(o[444]), .CLK(clk), .RST(rst), .Q(zreg[444]) );
  DFF \zreg_reg[445]  ( .D(o[445]), .CLK(clk), .RST(rst), .Q(zreg[445]) );
  DFF \zreg_reg[446]  ( .D(o[446]), .CLK(clk), .RST(rst), .Q(zreg[446]) );
  DFF \zreg_reg[447]  ( .D(o[447]), .CLK(clk), .RST(rst), .Q(zreg[447]) );
  DFF \zreg_reg[448]  ( .D(o[448]), .CLK(clk), .RST(rst), .Q(zreg[448]) );
  DFF \zreg_reg[449]  ( .D(o[449]), .CLK(clk), .RST(rst), .Q(zreg[449]) );
  DFF \zreg_reg[450]  ( .D(o[450]), .CLK(clk), .RST(rst), .Q(zreg[450]) );
  DFF \zreg_reg[451]  ( .D(o[451]), .CLK(clk), .RST(rst), .Q(zreg[451]) );
  DFF \zreg_reg[452]  ( .D(o[452]), .CLK(clk), .RST(rst), .Q(zreg[452]) );
  DFF \zreg_reg[453]  ( .D(o[453]), .CLK(clk), .RST(rst), .Q(zreg[453]) );
  DFF \zreg_reg[454]  ( .D(o[454]), .CLK(clk), .RST(rst), .Q(zreg[454]) );
  DFF \zreg_reg[455]  ( .D(o[455]), .CLK(clk), .RST(rst), .Q(zreg[455]) );
  DFF \zreg_reg[456]  ( .D(o[456]), .CLK(clk), .RST(rst), .Q(zreg[456]) );
  DFF \zreg_reg[457]  ( .D(o[457]), .CLK(clk), .RST(rst), .Q(zreg[457]) );
  DFF \zreg_reg[458]  ( .D(o[458]), .CLK(clk), .RST(rst), .Q(zreg[458]) );
  DFF \zreg_reg[459]  ( .D(o[459]), .CLK(clk), .RST(rst), .Q(zreg[459]) );
  DFF \zreg_reg[460]  ( .D(o[460]), .CLK(clk), .RST(rst), .Q(zreg[460]) );
  DFF \zreg_reg[461]  ( .D(o[461]), .CLK(clk), .RST(rst), .Q(zreg[461]) );
  DFF \zreg_reg[462]  ( .D(o[462]), .CLK(clk), .RST(rst), .Q(zreg[462]) );
  DFF \zreg_reg[463]  ( .D(o[463]), .CLK(clk), .RST(rst), .Q(zreg[463]) );
  DFF \zreg_reg[464]  ( .D(o[464]), .CLK(clk), .RST(rst), .Q(zreg[464]) );
  DFF \zreg_reg[465]  ( .D(o[465]), .CLK(clk), .RST(rst), .Q(zreg[465]) );
  DFF \zreg_reg[466]  ( .D(o[466]), .CLK(clk), .RST(rst), .Q(zreg[466]) );
  DFF \zreg_reg[467]  ( .D(o[467]), .CLK(clk), .RST(rst), .Q(zreg[467]) );
  DFF \zreg_reg[468]  ( .D(o[468]), .CLK(clk), .RST(rst), .Q(zreg[468]) );
  DFF \zreg_reg[469]  ( .D(o[469]), .CLK(clk), .RST(rst), .Q(zreg[469]) );
  DFF \zreg_reg[470]  ( .D(o[470]), .CLK(clk), .RST(rst), .Q(zreg[470]) );
  DFF \zreg_reg[471]  ( .D(o[471]), .CLK(clk), .RST(rst), .Q(zreg[471]) );
  DFF \zreg_reg[472]  ( .D(o[472]), .CLK(clk), .RST(rst), .Q(zreg[472]) );
  DFF \zreg_reg[473]  ( .D(o[473]), .CLK(clk), .RST(rst), .Q(zreg[473]) );
  DFF \zreg_reg[474]  ( .D(o[474]), .CLK(clk), .RST(rst), .Q(zreg[474]) );
  DFF \zreg_reg[475]  ( .D(o[475]), .CLK(clk), .RST(rst), .Q(zreg[475]) );
  DFF \zreg_reg[476]  ( .D(o[476]), .CLK(clk), .RST(rst), .Q(zreg[476]) );
  DFF \zreg_reg[477]  ( .D(o[477]), .CLK(clk), .RST(rst), .Q(zreg[477]) );
  DFF \zreg_reg[478]  ( .D(o[478]), .CLK(clk), .RST(rst), .Q(zreg[478]) );
  DFF \zreg_reg[479]  ( .D(o[479]), .CLK(clk), .RST(rst), .Q(zreg[479]) );
  DFF \zreg_reg[480]  ( .D(o[480]), .CLK(clk), .RST(rst), .Q(zreg[480]) );
  DFF \zreg_reg[481]  ( .D(o[481]), .CLK(clk), .RST(rst), .Q(zreg[481]) );
  DFF \zreg_reg[482]  ( .D(o[482]), .CLK(clk), .RST(rst), .Q(zreg[482]) );
  DFF \zreg_reg[483]  ( .D(o[483]), .CLK(clk), .RST(rst), .Q(zreg[483]) );
  DFF \zreg_reg[484]  ( .D(o[484]), .CLK(clk), .RST(rst), .Q(zreg[484]) );
  DFF \zreg_reg[485]  ( .D(o[485]), .CLK(clk), .RST(rst), .Q(zreg[485]) );
  DFF \zreg_reg[486]  ( .D(o[486]), .CLK(clk), .RST(rst), .Q(zreg[486]) );
  DFF \zreg_reg[487]  ( .D(o[487]), .CLK(clk), .RST(rst), .Q(zreg[487]) );
  DFF \zreg_reg[488]  ( .D(o[488]), .CLK(clk), .RST(rst), .Q(zreg[488]) );
  DFF \zreg_reg[489]  ( .D(o[489]), .CLK(clk), .RST(rst), .Q(zreg[489]) );
  DFF \zreg_reg[490]  ( .D(o[490]), .CLK(clk), .RST(rst), .Q(zreg[490]) );
  DFF \zreg_reg[491]  ( .D(o[491]), .CLK(clk), .RST(rst), .Q(zreg[491]) );
  DFF \zreg_reg[492]  ( .D(o[492]), .CLK(clk), .RST(rst), .Q(zreg[492]) );
  DFF \zreg_reg[493]  ( .D(o[493]), .CLK(clk), .RST(rst), .Q(zreg[493]) );
  DFF \zreg_reg[494]  ( .D(o[494]), .CLK(clk), .RST(rst), .Q(zreg[494]) );
  DFF \zreg_reg[495]  ( .D(o[495]), .CLK(clk), .RST(rst), .Q(zreg[495]) );
  DFF \zreg_reg[496]  ( .D(o[496]), .CLK(clk), .RST(rst), .Q(zreg[496]) );
  DFF \zreg_reg[497]  ( .D(o[497]), .CLK(clk), .RST(rst), .Q(zreg[497]) );
  DFF \zreg_reg[498]  ( .D(o[498]), .CLK(clk), .RST(rst), .Q(zreg[498]) );
  DFF \zreg_reg[499]  ( .D(o[499]), .CLK(clk), .RST(rst), .Q(zreg[499]) );
  DFF \zreg_reg[500]  ( .D(o[500]), .CLK(clk), .RST(rst), .Q(zreg[500]) );
  DFF \zreg_reg[501]  ( .D(o[501]), .CLK(clk), .RST(rst), .Q(zreg[501]) );
  DFF \zreg_reg[502]  ( .D(o[502]), .CLK(clk), .RST(rst), .Q(zreg[502]) );
  DFF \zreg_reg[503]  ( .D(o[503]), .CLK(clk), .RST(rst), .Q(zreg[503]) );
  DFF \zreg_reg[504]  ( .D(o[504]), .CLK(clk), .RST(rst), .Q(zreg[504]) );
  DFF \zreg_reg[505]  ( .D(o[505]), .CLK(clk), .RST(rst), .Q(zreg[505]) );
  DFF \zreg_reg[506]  ( .D(o[506]), .CLK(clk), .RST(rst), .Q(zreg[506]) );
  DFF \zreg_reg[507]  ( .D(o[507]), .CLK(clk), .RST(rst), .Q(zreg[507]) );
  DFF \zreg_reg[508]  ( .D(o[508]), .CLK(clk), .RST(rst), .Q(zreg[508]) );
  DFF \zreg_reg[509]  ( .D(o[509]), .CLK(clk), .RST(rst), .Q(zreg[509]) );
  DFF \zreg_reg[510]  ( .D(o[510]), .CLK(clk), .RST(rst), .Q(zreg[510]) );
  DFF \zreg_reg[511]  ( .D(o[511]), .CLK(clk), .RST(rst), .Q(zreg[511]) );
  DFF \zreg_reg[512]  ( .D(\zout[0][512] ), .CLK(clk), .RST(rst), .Q(zreg[512]) );
  DFF \zreg_reg[513]  ( .D(\zout[0][513] ), .CLK(clk), .RST(rst), .Q(zreg[513]) );
  modmult_step_N512 \MODMULT_STEP[0].modmult_step_  ( .xregN_1(xin[511]), .y(y), .n(n), .zin({\zin[0][513] , \zin[0][512] , \zin[0][511] , \zin[0][510] , 
        \zin[0][509] , \zin[0][508] , \zin[0][507] , \zin[0][506] , 
        \zin[0][505] , \zin[0][504] , \zin[0][503] , \zin[0][502] , 
        \zin[0][501] , \zin[0][500] , \zin[0][499] , \zin[0][498] , 
        \zin[0][497] , \zin[0][496] , \zin[0][495] , \zin[0][494] , 
        \zin[0][493] , \zin[0][492] , \zin[0][491] , \zin[0][490] , 
        \zin[0][489] , \zin[0][488] , \zin[0][487] , \zin[0][486] , 
        \zin[0][485] , \zin[0][484] , \zin[0][483] , \zin[0][482] , 
        \zin[0][481] , \zin[0][480] , \zin[0][479] , \zin[0][478] , 
        \zin[0][477] , \zin[0][476] , \zin[0][475] , \zin[0][474] , 
        \zin[0][473] , \zin[0][472] , \zin[0][471] , \zin[0][470] , 
        \zin[0][469] , \zin[0][468] , \zin[0][467] , \zin[0][466] , 
        \zin[0][465] , \zin[0][464] , \zin[0][463] , \zin[0][462] , 
        \zin[0][461] , \zin[0][460] , \zin[0][459] , \zin[0][458] , 
        \zin[0][457] , \zin[0][456] , \zin[0][455] , \zin[0][454] , 
        \zin[0][453] , \zin[0][452] , \zin[0][451] , \zin[0][450] , 
        \zin[0][449] , \zin[0][448] , \zin[0][447] , \zin[0][446] , 
        \zin[0][445] , \zin[0][444] , \zin[0][443] , \zin[0][442] , 
        \zin[0][441] , \zin[0][440] , \zin[0][439] , \zin[0][438] , 
        \zin[0][437] , \zin[0][436] , \zin[0][435] , \zin[0][434] , 
        \zin[0][433] , \zin[0][432] , \zin[0][431] , \zin[0][430] , 
        \zin[0][429] , \zin[0][428] , \zin[0][427] , \zin[0][426] , 
        \zin[0][425] , \zin[0][424] , \zin[0][423] , \zin[0][422] , 
        \zin[0][421] , \zin[0][420] , \zin[0][419] , \zin[0][418] , 
        \zin[0][417] , \zin[0][416] , \zin[0][415] , \zin[0][414] , 
        \zin[0][413] , \zin[0][412] , \zin[0][411] , \zin[0][410] , 
        \zin[0][409] , \zin[0][408] , \zin[0][407] , \zin[0][406] , 
        \zin[0][405] , \zin[0][404] , \zin[0][403] , \zin[0][402] , 
        \zin[0][401] , \zin[0][400] , \zin[0][399] , \zin[0][398] , 
        \zin[0][397] , \zin[0][396] , \zin[0][395] , \zin[0][394] , 
        \zin[0][393] , \zin[0][392] , \zin[0][391] , \zin[0][390] , 
        \zin[0][389] , \zin[0][388] , \zin[0][387] , \zin[0][386] , 
        \zin[0][385] , \zin[0][384] , \zin[0][383] , \zin[0][382] , 
        \zin[0][381] , \zin[0][380] , \zin[0][379] , \zin[0][378] , 
        \zin[0][377] , \zin[0][376] , \zin[0][375] , \zin[0][374] , 
        \zin[0][373] , \zin[0][372] , \zin[0][371] , \zin[0][370] , 
        \zin[0][369] , \zin[0][368] , \zin[0][367] , \zin[0][366] , 
        \zin[0][365] , \zin[0][364] , \zin[0][363] , \zin[0][362] , 
        \zin[0][361] , \zin[0][360] , \zin[0][359] , \zin[0][358] , 
        \zin[0][357] , \zin[0][356] , \zin[0][355] , \zin[0][354] , 
        \zin[0][353] , \zin[0][352] , \zin[0][351] , \zin[0][350] , 
        \zin[0][349] , \zin[0][348] , \zin[0][347] , \zin[0][346] , 
        \zin[0][345] , \zin[0][344] , \zin[0][343] , \zin[0][342] , 
        \zin[0][341] , \zin[0][340] , \zin[0][339] , \zin[0][338] , 
        \zin[0][337] , \zin[0][336] , \zin[0][335] , \zin[0][334] , 
        \zin[0][333] , \zin[0][332] , \zin[0][331] , \zin[0][330] , 
        \zin[0][329] , \zin[0][328] , \zin[0][327] , \zin[0][326] , 
        \zin[0][325] , \zin[0][324] , \zin[0][323] , \zin[0][322] , 
        \zin[0][321] , \zin[0][320] , \zin[0][319] , \zin[0][318] , 
        \zin[0][317] , \zin[0][316] , \zin[0][315] , \zin[0][314] , 
        \zin[0][313] , \zin[0][312] , \zin[0][311] , \zin[0][310] , 
        \zin[0][309] , \zin[0][308] , \zin[0][307] , \zin[0][306] , 
        \zin[0][305] , \zin[0][304] , \zin[0][303] , \zin[0][302] , 
        \zin[0][301] , \zin[0][300] , \zin[0][299] , \zin[0][298] , 
        \zin[0][297] , \zin[0][296] , \zin[0][295] , \zin[0][294] , 
        \zin[0][293] , \zin[0][292] , \zin[0][291] , \zin[0][290] , 
        \zin[0][289] , \zin[0][288] , \zin[0][287] , \zin[0][286] , 
        \zin[0][285] , \zin[0][284] , \zin[0][283] , \zin[0][282] , 
        \zin[0][281] , \zin[0][280] , \zin[0][279] , \zin[0][278] , 
        \zin[0][277] , \zin[0][276] , \zin[0][275] , \zin[0][274] , 
        \zin[0][273] , \zin[0][272] , \zin[0][271] , \zin[0][270] , 
        \zin[0][269] , \zin[0][268] , \zin[0][267] , \zin[0][266] , 
        \zin[0][265] , \zin[0][264] , \zin[0][263] , \zin[0][262] , 
        \zin[0][261] , \zin[0][260] , \zin[0][259] , \zin[0][258] , 
        \zin[0][257] , \zin[0][256] , \zin[0][255] , \zin[0][254] , 
        \zin[0][253] , \zin[0][252] , \zin[0][251] , \zin[0][250] , 
        \zin[0][249] , \zin[0][248] , \zin[0][247] , \zin[0][246] , 
        \zin[0][245] , \zin[0][244] , \zin[0][243] , \zin[0][242] , 
        \zin[0][241] , \zin[0][240] , \zin[0][239] , \zin[0][238] , 
        \zin[0][237] , \zin[0][236] , \zin[0][235] , \zin[0][234] , 
        \zin[0][233] , \zin[0][232] , \zin[0][231] , \zin[0][230] , 
        \zin[0][229] , \zin[0][228] , \zin[0][227] , \zin[0][226] , 
        \zin[0][225] , \zin[0][224] , \zin[0][223] , \zin[0][222] , 
        \zin[0][221] , \zin[0][220] , \zin[0][219] , \zin[0][218] , 
        \zin[0][217] , \zin[0][216] , \zin[0][215] , \zin[0][214] , 
        \zin[0][213] , \zin[0][212] , \zin[0][211] , \zin[0][210] , 
        \zin[0][209] , \zin[0][208] , \zin[0][207] , \zin[0][206] , 
        \zin[0][205] , \zin[0][204] , \zin[0][203] , \zin[0][202] , 
        \zin[0][201] , \zin[0][200] , \zin[0][199] , \zin[0][198] , 
        \zin[0][197] , \zin[0][196] , \zin[0][195] , \zin[0][194] , 
        \zin[0][193] , \zin[0][192] , \zin[0][191] , \zin[0][190] , 
        \zin[0][189] , \zin[0][188] , \zin[0][187] , \zin[0][186] , 
        \zin[0][185] , \zin[0][184] , \zin[0][183] , \zin[0][182] , 
        \zin[0][181] , \zin[0][180] , \zin[0][179] , \zin[0][178] , 
        \zin[0][177] , \zin[0][176] , \zin[0][175] , \zin[0][174] , 
        \zin[0][173] , \zin[0][172] , \zin[0][171] , \zin[0][170] , 
        \zin[0][169] , \zin[0][168] , \zin[0][167] , \zin[0][166] , 
        \zin[0][165] , \zin[0][164] , \zin[0][163] , \zin[0][162] , 
        \zin[0][161] , \zin[0][160] , \zin[0][159] , \zin[0][158] , 
        \zin[0][157] , \zin[0][156] , \zin[0][155] , \zin[0][154] , 
        \zin[0][153] , \zin[0][152] , \zin[0][151] , \zin[0][150] , 
        \zin[0][149] , \zin[0][148] , \zin[0][147] , \zin[0][146] , 
        \zin[0][145] , \zin[0][144] , \zin[0][143] , \zin[0][142] , 
        \zin[0][141] , \zin[0][140] , \zin[0][139] , \zin[0][138] , 
        \zin[0][137] , \zin[0][136] , \zin[0][135] , \zin[0][134] , 
        \zin[0][133] , \zin[0][132] , \zin[0][131] , \zin[0][130] , 
        \zin[0][129] , \zin[0][128] , \zin[0][127] , \zin[0][126] , 
        \zin[0][125] , \zin[0][124] , \zin[0][123] , \zin[0][122] , 
        \zin[0][121] , \zin[0][120] , \zin[0][119] , \zin[0][118] , 
        \zin[0][117] , \zin[0][116] , \zin[0][115] , \zin[0][114] , 
        \zin[0][113] , \zin[0][112] , \zin[0][111] , \zin[0][110] , 
        \zin[0][109] , \zin[0][108] , \zin[0][107] , \zin[0][106] , 
        \zin[0][105] , \zin[0][104] , \zin[0][103] , \zin[0][102] , 
        \zin[0][101] , \zin[0][100] , \zin[0][99] , \zin[0][98] , \zin[0][97] , 
        \zin[0][96] , \zin[0][95] , \zin[0][94] , \zin[0][93] , \zin[0][92] , 
        \zin[0][91] , \zin[0][90] , \zin[0][89] , \zin[0][88] , \zin[0][87] , 
        \zin[0][86] , \zin[0][85] , \zin[0][84] , \zin[0][83] , \zin[0][82] , 
        \zin[0][81] , \zin[0][80] , \zin[0][79] , \zin[0][78] , \zin[0][77] , 
        \zin[0][76] , \zin[0][75] , \zin[0][74] , \zin[0][73] , \zin[0][72] , 
        \zin[0][71] , \zin[0][70] , \zin[0][69] , \zin[0][68] , \zin[0][67] , 
        \zin[0][66] , \zin[0][65] , \zin[0][64] , \zin[0][63] , \zin[0][62] , 
        \zin[0][61] , \zin[0][60] , \zin[0][59] , \zin[0][58] , \zin[0][57] , 
        \zin[0][56] , \zin[0][55] , \zin[0][54] , \zin[0][53] , \zin[0][52] , 
        \zin[0][51] , \zin[0][50] , \zin[0][49] , \zin[0][48] , \zin[0][47] , 
        \zin[0][46] , \zin[0][45] , \zin[0][44] , \zin[0][43] , \zin[0][42] , 
        \zin[0][41] , \zin[0][40] , \zin[0][39] , \zin[0][38] , \zin[0][37] , 
        \zin[0][36] , \zin[0][35] , \zin[0][34] , \zin[0][33] , \zin[0][32] , 
        \zin[0][31] , \zin[0][30] , \zin[0][29] , \zin[0][28] , \zin[0][27] , 
        \zin[0][26] , \zin[0][25] , \zin[0][24] , \zin[0][23] , \zin[0][22] , 
        \zin[0][21] , \zin[0][20] , \zin[0][19] , \zin[0][18] , \zin[0][17] , 
        \zin[0][16] , \zin[0][15] , \zin[0][14] , \zin[0][13] , \zin[0][12] , 
        \zin[0][11] , \zin[0][10] , \zin[0][9] , \zin[0][8] , \zin[0][7] , 
        \zin[0][6] , \zin[0][5] , \zin[0][4] , \zin[0][3] , \zin[0][2] , 
        \zin[0][1] , \zin[0][0] }), .zout({\zout[0][513] , \zout[0][512] , o})
         );
  ANDN U3 ( .B(zreg[9]), .A(start), .Z(\zin[0][9] ) );
  ANDN U4 ( .B(zreg[99]), .A(start), .Z(\zin[0][99] ) );
  ANDN U5 ( .B(zreg[98]), .A(start), .Z(\zin[0][98] ) );
  ANDN U6 ( .B(zreg[97]), .A(start), .Z(\zin[0][97] ) );
  ANDN U7 ( .B(zreg[96]), .A(start), .Z(\zin[0][96] ) );
  ANDN U8 ( .B(zreg[95]), .A(start), .Z(\zin[0][95] ) );
  ANDN U9 ( .B(zreg[94]), .A(start), .Z(\zin[0][94] ) );
  ANDN U10 ( .B(zreg[93]), .A(start), .Z(\zin[0][93] ) );
  ANDN U11 ( .B(zreg[92]), .A(start), .Z(\zin[0][92] ) );
  ANDN U12 ( .B(zreg[91]), .A(start), .Z(\zin[0][91] ) );
  ANDN U13 ( .B(zreg[90]), .A(start), .Z(\zin[0][90] ) );
  ANDN U14 ( .B(zreg[8]), .A(start), .Z(\zin[0][8] ) );
  ANDN U15 ( .B(zreg[89]), .A(start), .Z(\zin[0][89] ) );
  ANDN U16 ( .B(zreg[88]), .A(start), .Z(\zin[0][88] ) );
  ANDN U17 ( .B(zreg[87]), .A(start), .Z(\zin[0][87] ) );
  ANDN U18 ( .B(zreg[86]), .A(start), .Z(\zin[0][86] ) );
  ANDN U19 ( .B(zreg[85]), .A(start), .Z(\zin[0][85] ) );
  ANDN U20 ( .B(zreg[84]), .A(start), .Z(\zin[0][84] ) );
  ANDN U21 ( .B(zreg[83]), .A(start), .Z(\zin[0][83] ) );
  ANDN U22 ( .B(zreg[82]), .A(start), .Z(\zin[0][82] ) );
  ANDN U23 ( .B(zreg[81]), .A(start), .Z(\zin[0][81] ) );
  ANDN U24 ( .B(zreg[80]), .A(start), .Z(\zin[0][80] ) );
  ANDN U25 ( .B(zreg[7]), .A(start), .Z(\zin[0][7] ) );
  ANDN U26 ( .B(zreg[79]), .A(start), .Z(\zin[0][79] ) );
  ANDN U27 ( .B(zreg[78]), .A(start), .Z(\zin[0][78] ) );
  ANDN U28 ( .B(zreg[77]), .A(start), .Z(\zin[0][77] ) );
  ANDN U29 ( .B(zreg[76]), .A(start), .Z(\zin[0][76] ) );
  ANDN U30 ( .B(zreg[75]), .A(start), .Z(\zin[0][75] ) );
  ANDN U31 ( .B(zreg[74]), .A(start), .Z(\zin[0][74] ) );
  ANDN U32 ( .B(zreg[73]), .A(start), .Z(\zin[0][73] ) );
  ANDN U33 ( .B(zreg[72]), .A(start), .Z(\zin[0][72] ) );
  ANDN U34 ( .B(zreg[71]), .A(start), .Z(\zin[0][71] ) );
  ANDN U35 ( .B(zreg[70]), .A(start), .Z(\zin[0][70] ) );
  ANDN U36 ( .B(zreg[6]), .A(start), .Z(\zin[0][6] ) );
  ANDN U37 ( .B(zreg[69]), .A(start), .Z(\zin[0][69] ) );
  ANDN U38 ( .B(zreg[68]), .A(start), .Z(\zin[0][68] ) );
  ANDN U39 ( .B(zreg[67]), .A(start), .Z(\zin[0][67] ) );
  ANDN U40 ( .B(zreg[66]), .A(start), .Z(\zin[0][66] ) );
  ANDN U41 ( .B(zreg[65]), .A(start), .Z(\zin[0][65] ) );
  ANDN U42 ( .B(zreg[64]), .A(start), .Z(\zin[0][64] ) );
  ANDN U43 ( .B(zreg[63]), .A(start), .Z(\zin[0][63] ) );
  ANDN U44 ( .B(zreg[62]), .A(start), .Z(\zin[0][62] ) );
  ANDN U45 ( .B(zreg[61]), .A(start), .Z(\zin[0][61] ) );
  ANDN U46 ( .B(zreg[60]), .A(start), .Z(\zin[0][60] ) );
  ANDN U47 ( .B(zreg[5]), .A(start), .Z(\zin[0][5] ) );
  ANDN U48 ( .B(zreg[59]), .A(start), .Z(\zin[0][59] ) );
  ANDN U49 ( .B(zreg[58]), .A(start), .Z(\zin[0][58] ) );
  ANDN U50 ( .B(zreg[57]), .A(start), .Z(\zin[0][57] ) );
  ANDN U51 ( .B(zreg[56]), .A(start), .Z(\zin[0][56] ) );
  ANDN U52 ( .B(zreg[55]), .A(start), .Z(\zin[0][55] ) );
  ANDN U53 ( .B(zreg[54]), .A(start), .Z(\zin[0][54] ) );
  ANDN U54 ( .B(zreg[53]), .A(start), .Z(\zin[0][53] ) );
  ANDN U55 ( .B(zreg[52]), .A(start), .Z(\zin[0][52] ) );
  ANDN U56 ( .B(zreg[51]), .A(start), .Z(\zin[0][51] ) );
  ANDN U57 ( .B(zreg[513]), .A(start), .Z(\zin[0][513] ) );
  ANDN U58 ( .B(zreg[512]), .A(start), .Z(\zin[0][512] ) );
  ANDN U59 ( .B(zreg[511]), .A(start), .Z(\zin[0][511] ) );
  ANDN U60 ( .B(zreg[510]), .A(start), .Z(\zin[0][510] ) );
  ANDN U61 ( .B(zreg[50]), .A(start), .Z(\zin[0][50] ) );
  ANDN U62 ( .B(zreg[509]), .A(start), .Z(\zin[0][509] ) );
  ANDN U63 ( .B(zreg[508]), .A(start), .Z(\zin[0][508] ) );
  ANDN U64 ( .B(zreg[507]), .A(start), .Z(\zin[0][507] ) );
  ANDN U65 ( .B(zreg[506]), .A(start), .Z(\zin[0][506] ) );
  ANDN U66 ( .B(zreg[505]), .A(start), .Z(\zin[0][505] ) );
  ANDN U67 ( .B(zreg[504]), .A(start), .Z(\zin[0][504] ) );
  ANDN U68 ( .B(zreg[503]), .A(start), .Z(\zin[0][503] ) );
  ANDN U69 ( .B(zreg[502]), .A(start), .Z(\zin[0][502] ) );
  ANDN U70 ( .B(zreg[501]), .A(start), .Z(\zin[0][501] ) );
  ANDN U71 ( .B(zreg[500]), .A(start), .Z(\zin[0][500] ) );
  ANDN U72 ( .B(zreg[4]), .A(start), .Z(\zin[0][4] ) );
  ANDN U73 ( .B(zreg[49]), .A(start), .Z(\zin[0][49] ) );
  ANDN U74 ( .B(zreg[499]), .A(start), .Z(\zin[0][499] ) );
  ANDN U75 ( .B(zreg[498]), .A(start), .Z(\zin[0][498] ) );
  ANDN U76 ( .B(zreg[497]), .A(start), .Z(\zin[0][497] ) );
  ANDN U77 ( .B(zreg[496]), .A(start), .Z(\zin[0][496] ) );
  ANDN U78 ( .B(zreg[495]), .A(start), .Z(\zin[0][495] ) );
  ANDN U79 ( .B(zreg[494]), .A(start), .Z(\zin[0][494] ) );
  ANDN U80 ( .B(zreg[493]), .A(start), .Z(\zin[0][493] ) );
  ANDN U81 ( .B(zreg[492]), .A(start), .Z(\zin[0][492] ) );
  ANDN U82 ( .B(zreg[491]), .A(start), .Z(\zin[0][491] ) );
  ANDN U83 ( .B(zreg[490]), .A(start), .Z(\zin[0][490] ) );
  ANDN U84 ( .B(zreg[48]), .A(start), .Z(\zin[0][48] ) );
  ANDN U85 ( .B(zreg[489]), .A(start), .Z(\zin[0][489] ) );
  ANDN U86 ( .B(zreg[488]), .A(start), .Z(\zin[0][488] ) );
  ANDN U87 ( .B(zreg[487]), .A(start), .Z(\zin[0][487] ) );
  ANDN U88 ( .B(zreg[486]), .A(start), .Z(\zin[0][486] ) );
  ANDN U89 ( .B(zreg[485]), .A(start), .Z(\zin[0][485] ) );
  ANDN U90 ( .B(zreg[484]), .A(start), .Z(\zin[0][484] ) );
  ANDN U91 ( .B(zreg[483]), .A(start), .Z(\zin[0][483] ) );
  ANDN U92 ( .B(zreg[482]), .A(start), .Z(\zin[0][482] ) );
  ANDN U93 ( .B(zreg[481]), .A(start), .Z(\zin[0][481] ) );
  ANDN U94 ( .B(zreg[480]), .A(start), .Z(\zin[0][480] ) );
  ANDN U95 ( .B(zreg[47]), .A(start), .Z(\zin[0][47] ) );
  ANDN U96 ( .B(zreg[479]), .A(start), .Z(\zin[0][479] ) );
  ANDN U97 ( .B(zreg[478]), .A(start), .Z(\zin[0][478] ) );
  ANDN U98 ( .B(zreg[477]), .A(start), .Z(\zin[0][477] ) );
  ANDN U99 ( .B(zreg[476]), .A(start), .Z(\zin[0][476] ) );
  ANDN U100 ( .B(zreg[475]), .A(start), .Z(\zin[0][475] ) );
  ANDN U101 ( .B(zreg[474]), .A(start), .Z(\zin[0][474] ) );
  ANDN U102 ( .B(zreg[473]), .A(start), .Z(\zin[0][473] ) );
  ANDN U103 ( .B(zreg[472]), .A(start), .Z(\zin[0][472] ) );
  ANDN U104 ( .B(zreg[471]), .A(start), .Z(\zin[0][471] ) );
  ANDN U105 ( .B(zreg[470]), .A(start), .Z(\zin[0][470] ) );
  ANDN U106 ( .B(zreg[46]), .A(start), .Z(\zin[0][46] ) );
  ANDN U107 ( .B(zreg[469]), .A(start), .Z(\zin[0][469] ) );
  ANDN U108 ( .B(zreg[468]), .A(start), .Z(\zin[0][468] ) );
  ANDN U109 ( .B(zreg[467]), .A(start), .Z(\zin[0][467] ) );
  ANDN U110 ( .B(zreg[466]), .A(start), .Z(\zin[0][466] ) );
  ANDN U111 ( .B(zreg[465]), .A(start), .Z(\zin[0][465] ) );
  ANDN U112 ( .B(zreg[464]), .A(start), .Z(\zin[0][464] ) );
  ANDN U113 ( .B(zreg[463]), .A(start), .Z(\zin[0][463] ) );
  ANDN U114 ( .B(zreg[462]), .A(start), .Z(\zin[0][462] ) );
  ANDN U115 ( .B(zreg[461]), .A(start), .Z(\zin[0][461] ) );
  ANDN U116 ( .B(zreg[460]), .A(start), .Z(\zin[0][460] ) );
  ANDN U117 ( .B(zreg[45]), .A(start), .Z(\zin[0][45] ) );
  ANDN U118 ( .B(zreg[459]), .A(start), .Z(\zin[0][459] ) );
  ANDN U119 ( .B(zreg[458]), .A(start), .Z(\zin[0][458] ) );
  ANDN U120 ( .B(zreg[457]), .A(start), .Z(\zin[0][457] ) );
  ANDN U121 ( .B(zreg[456]), .A(start), .Z(\zin[0][456] ) );
  ANDN U122 ( .B(zreg[455]), .A(start), .Z(\zin[0][455] ) );
  ANDN U123 ( .B(zreg[454]), .A(start), .Z(\zin[0][454] ) );
  ANDN U124 ( .B(zreg[453]), .A(start), .Z(\zin[0][453] ) );
  ANDN U125 ( .B(zreg[452]), .A(start), .Z(\zin[0][452] ) );
  ANDN U126 ( .B(zreg[451]), .A(start), .Z(\zin[0][451] ) );
  ANDN U127 ( .B(zreg[450]), .A(start), .Z(\zin[0][450] ) );
  ANDN U128 ( .B(zreg[44]), .A(start), .Z(\zin[0][44] ) );
  ANDN U129 ( .B(zreg[449]), .A(start), .Z(\zin[0][449] ) );
  ANDN U130 ( .B(zreg[448]), .A(start), .Z(\zin[0][448] ) );
  ANDN U131 ( .B(zreg[447]), .A(start), .Z(\zin[0][447] ) );
  ANDN U132 ( .B(zreg[446]), .A(start), .Z(\zin[0][446] ) );
  ANDN U133 ( .B(zreg[445]), .A(start), .Z(\zin[0][445] ) );
  ANDN U134 ( .B(zreg[444]), .A(start), .Z(\zin[0][444] ) );
  ANDN U135 ( .B(zreg[443]), .A(start), .Z(\zin[0][443] ) );
  ANDN U136 ( .B(zreg[442]), .A(start), .Z(\zin[0][442] ) );
  ANDN U137 ( .B(zreg[441]), .A(start), .Z(\zin[0][441] ) );
  ANDN U138 ( .B(zreg[440]), .A(start), .Z(\zin[0][440] ) );
  ANDN U139 ( .B(zreg[43]), .A(start), .Z(\zin[0][43] ) );
  ANDN U140 ( .B(zreg[439]), .A(start), .Z(\zin[0][439] ) );
  ANDN U141 ( .B(zreg[438]), .A(start), .Z(\zin[0][438] ) );
  ANDN U142 ( .B(zreg[437]), .A(start), .Z(\zin[0][437] ) );
  ANDN U143 ( .B(zreg[436]), .A(start), .Z(\zin[0][436] ) );
  ANDN U144 ( .B(zreg[435]), .A(start), .Z(\zin[0][435] ) );
  ANDN U145 ( .B(zreg[434]), .A(start), .Z(\zin[0][434] ) );
  ANDN U146 ( .B(zreg[433]), .A(start), .Z(\zin[0][433] ) );
  ANDN U147 ( .B(zreg[432]), .A(start), .Z(\zin[0][432] ) );
  ANDN U148 ( .B(zreg[431]), .A(start), .Z(\zin[0][431] ) );
  ANDN U149 ( .B(zreg[430]), .A(start), .Z(\zin[0][430] ) );
  ANDN U150 ( .B(zreg[42]), .A(start), .Z(\zin[0][42] ) );
  ANDN U151 ( .B(zreg[429]), .A(start), .Z(\zin[0][429] ) );
  ANDN U152 ( .B(zreg[428]), .A(start), .Z(\zin[0][428] ) );
  ANDN U153 ( .B(zreg[427]), .A(start), .Z(\zin[0][427] ) );
  ANDN U154 ( .B(zreg[426]), .A(start), .Z(\zin[0][426] ) );
  ANDN U155 ( .B(zreg[425]), .A(start), .Z(\zin[0][425] ) );
  ANDN U156 ( .B(zreg[424]), .A(start), .Z(\zin[0][424] ) );
  ANDN U157 ( .B(zreg[423]), .A(start), .Z(\zin[0][423] ) );
  ANDN U158 ( .B(zreg[422]), .A(start), .Z(\zin[0][422] ) );
  ANDN U159 ( .B(zreg[421]), .A(start), .Z(\zin[0][421] ) );
  ANDN U160 ( .B(zreg[420]), .A(start), .Z(\zin[0][420] ) );
  ANDN U161 ( .B(zreg[41]), .A(start), .Z(\zin[0][41] ) );
  ANDN U162 ( .B(zreg[419]), .A(start), .Z(\zin[0][419] ) );
  ANDN U163 ( .B(zreg[418]), .A(start), .Z(\zin[0][418] ) );
  ANDN U164 ( .B(zreg[417]), .A(start), .Z(\zin[0][417] ) );
  ANDN U165 ( .B(zreg[416]), .A(start), .Z(\zin[0][416] ) );
  ANDN U166 ( .B(zreg[415]), .A(start), .Z(\zin[0][415] ) );
  ANDN U167 ( .B(zreg[414]), .A(start), .Z(\zin[0][414] ) );
  ANDN U168 ( .B(zreg[413]), .A(start), .Z(\zin[0][413] ) );
  ANDN U169 ( .B(zreg[412]), .A(start), .Z(\zin[0][412] ) );
  ANDN U170 ( .B(zreg[411]), .A(start), .Z(\zin[0][411] ) );
  ANDN U171 ( .B(zreg[410]), .A(start), .Z(\zin[0][410] ) );
  ANDN U172 ( .B(zreg[40]), .A(start), .Z(\zin[0][40] ) );
  ANDN U173 ( .B(zreg[409]), .A(start), .Z(\zin[0][409] ) );
  ANDN U174 ( .B(zreg[408]), .A(start), .Z(\zin[0][408] ) );
  ANDN U175 ( .B(zreg[407]), .A(start), .Z(\zin[0][407] ) );
  ANDN U176 ( .B(zreg[406]), .A(start), .Z(\zin[0][406] ) );
  ANDN U177 ( .B(zreg[405]), .A(start), .Z(\zin[0][405] ) );
  ANDN U178 ( .B(zreg[404]), .A(start), .Z(\zin[0][404] ) );
  ANDN U179 ( .B(zreg[403]), .A(start), .Z(\zin[0][403] ) );
  ANDN U180 ( .B(zreg[402]), .A(start), .Z(\zin[0][402] ) );
  ANDN U181 ( .B(zreg[401]), .A(start), .Z(\zin[0][401] ) );
  ANDN U182 ( .B(zreg[400]), .A(start), .Z(\zin[0][400] ) );
  ANDN U183 ( .B(zreg[3]), .A(start), .Z(\zin[0][3] ) );
  ANDN U184 ( .B(zreg[39]), .A(start), .Z(\zin[0][39] ) );
  ANDN U185 ( .B(zreg[399]), .A(start), .Z(\zin[0][399] ) );
  ANDN U186 ( .B(zreg[398]), .A(start), .Z(\zin[0][398] ) );
  ANDN U187 ( .B(zreg[397]), .A(start), .Z(\zin[0][397] ) );
  ANDN U188 ( .B(zreg[396]), .A(start), .Z(\zin[0][396] ) );
  ANDN U189 ( .B(zreg[395]), .A(start), .Z(\zin[0][395] ) );
  ANDN U190 ( .B(zreg[394]), .A(start), .Z(\zin[0][394] ) );
  ANDN U191 ( .B(zreg[393]), .A(start), .Z(\zin[0][393] ) );
  ANDN U192 ( .B(zreg[392]), .A(start), .Z(\zin[0][392] ) );
  ANDN U193 ( .B(zreg[391]), .A(start), .Z(\zin[0][391] ) );
  ANDN U194 ( .B(zreg[390]), .A(start), .Z(\zin[0][390] ) );
  ANDN U195 ( .B(zreg[38]), .A(start), .Z(\zin[0][38] ) );
  ANDN U196 ( .B(zreg[389]), .A(start), .Z(\zin[0][389] ) );
  ANDN U197 ( .B(zreg[388]), .A(start), .Z(\zin[0][388] ) );
  ANDN U198 ( .B(zreg[387]), .A(start), .Z(\zin[0][387] ) );
  ANDN U199 ( .B(zreg[386]), .A(start), .Z(\zin[0][386] ) );
  ANDN U200 ( .B(zreg[385]), .A(start), .Z(\zin[0][385] ) );
  ANDN U201 ( .B(zreg[384]), .A(start), .Z(\zin[0][384] ) );
  ANDN U202 ( .B(zreg[383]), .A(start), .Z(\zin[0][383] ) );
  ANDN U203 ( .B(zreg[382]), .A(start), .Z(\zin[0][382] ) );
  ANDN U204 ( .B(zreg[381]), .A(start), .Z(\zin[0][381] ) );
  ANDN U205 ( .B(zreg[380]), .A(start), .Z(\zin[0][380] ) );
  ANDN U206 ( .B(zreg[37]), .A(start), .Z(\zin[0][37] ) );
  ANDN U207 ( .B(zreg[379]), .A(start), .Z(\zin[0][379] ) );
  ANDN U208 ( .B(zreg[378]), .A(start), .Z(\zin[0][378] ) );
  ANDN U209 ( .B(zreg[377]), .A(start), .Z(\zin[0][377] ) );
  ANDN U210 ( .B(zreg[376]), .A(start), .Z(\zin[0][376] ) );
  ANDN U211 ( .B(zreg[375]), .A(start), .Z(\zin[0][375] ) );
  ANDN U212 ( .B(zreg[374]), .A(start), .Z(\zin[0][374] ) );
  ANDN U213 ( .B(zreg[373]), .A(start), .Z(\zin[0][373] ) );
  ANDN U214 ( .B(zreg[372]), .A(start), .Z(\zin[0][372] ) );
  ANDN U215 ( .B(zreg[371]), .A(start), .Z(\zin[0][371] ) );
  ANDN U216 ( .B(zreg[370]), .A(start), .Z(\zin[0][370] ) );
  ANDN U217 ( .B(zreg[36]), .A(start), .Z(\zin[0][36] ) );
  ANDN U218 ( .B(zreg[369]), .A(start), .Z(\zin[0][369] ) );
  ANDN U219 ( .B(zreg[368]), .A(start), .Z(\zin[0][368] ) );
  ANDN U220 ( .B(zreg[367]), .A(start), .Z(\zin[0][367] ) );
  ANDN U221 ( .B(zreg[366]), .A(start), .Z(\zin[0][366] ) );
  ANDN U222 ( .B(zreg[365]), .A(start), .Z(\zin[0][365] ) );
  ANDN U223 ( .B(zreg[364]), .A(start), .Z(\zin[0][364] ) );
  ANDN U224 ( .B(zreg[363]), .A(start), .Z(\zin[0][363] ) );
  ANDN U225 ( .B(zreg[362]), .A(start), .Z(\zin[0][362] ) );
  ANDN U226 ( .B(zreg[361]), .A(start), .Z(\zin[0][361] ) );
  ANDN U227 ( .B(zreg[360]), .A(start), .Z(\zin[0][360] ) );
  ANDN U228 ( .B(zreg[35]), .A(start), .Z(\zin[0][35] ) );
  ANDN U229 ( .B(zreg[359]), .A(start), .Z(\zin[0][359] ) );
  ANDN U230 ( .B(zreg[358]), .A(start), .Z(\zin[0][358] ) );
  ANDN U231 ( .B(zreg[357]), .A(start), .Z(\zin[0][357] ) );
  ANDN U232 ( .B(zreg[356]), .A(start), .Z(\zin[0][356] ) );
  ANDN U233 ( .B(zreg[355]), .A(start), .Z(\zin[0][355] ) );
  ANDN U234 ( .B(zreg[354]), .A(start), .Z(\zin[0][354] ) );
  ANDN U235 ( .B(zreg[353]), .A(start), .Z(\zin[0][353] ) );
  ANDN U236 ( .B(zreg[352]), .A(start), .Z(\zin[0][352] ) );
  ANDN U237 ( .B(zreg[351]), .A(start), .Z(\zin[0][351] ) );
  ANDN U238 ( .B(zreg[350]), .A(start), .Z(\zin[0][350] ) );
  ANDN U239 ( .B(zreg[34]), .A(start), .Z(\zin[0][34] ) );
  ANDN U240 ( .B(zreg[349]), .A(start), .Z(\zin[0][349] ) );
  ANDN U241 ( .B(zreg[348]), .A(start), .Z(\zin[0][348] ) );
  ANDN U242 ( .B(zreg[347]), .A(start), .Z(\zin[0][347] ) );
  ANDN U243 ( .B(zreg[346]), .A(start), .Z(\zin[0][346] ) );
  ANDN U244 ( .B(zreg[345]), .A(start), .Z(\zin[0][345] ) );
  ANDN U245 ( .B(zreg[344]), .A(start), .Z(\zin[0][344] ) );
  ANDN U246 ( .B(zreg[343]), .A(start), .Z(\zin[0][343] ) );
  ANDN U247 ( .B(zreg[342]), .A(start), .Z(\zin[0][342] ) );
  ANDN U248 ( .B(zreg[341]), .A(start), .Z(\zin[0][341] ) );
  ANDN U249 ( .B(zreg[340]), .A(start), .Z(\zin[0][340] ) );
  ANDN U250 ( .B(zreg[33]), .A(start), .Z(\zin[0][33] ) );
  ANDN U251 ( .B(zreg[339]), .A(start), .Z(\zin[0][339] ) );
  ANDN U252 ( .B(zreg[338]), .A(start), .Z(\zin[0][338] ) );
  ANDN U253 ( .B(zreg[337]), .A(start), .Z(\zin[0][337] ) );
  ANDN U254 ( .B(zreg[336]), .A(start), .Z(\zin[0][336] ) );
  ANDN U255 ( .B(zreg[335]), .A(start), .Z(\zin[0][335] ) );
  ANDN U256 ( .B(zreg[334]), .A(start), .Z(\zin[0][334] ) );
  ANDN U257 ( .B(zreg[333]), .A(start), .Z(\zin[0][333] ) );
  ANDN U258 ( .B(zreg[332]), .A(start), .Z(\zin[0][332] ) );
  ANDN U259 ( .B(zreg[331]), .A(start), .Z(\zin[0][331] ) );
  ANDN U260 ( .B(zreg[330]), .A(start), .Z(\zin[0][330] ) );
  ANDN U261 ( .B(zreg[32]), .A(start), .Z(\zin[0][32] ) );
  ANDN U262 ( .B(zreg[329]), .A(start), .Z(\zin[0][329] ) );
  ANDN U263 ( .B(zreg[328]), .A(start), .Z(\zin[0][328] ) );
  ANDN U264 ( .B(zreg[327]), .A(start), .Z(\zin[0][327] ) );
  ANDN U265 ( .B(zreg[326]), .A(start), .Z(\zin[0][326] ) );
  ANDN U266 ( .B(zreg[325]), .A(start), .Z(\zin[0][325] ) );
  ANDN U267 ( .B(zreg[324]), .A(start), .Z(\zin[0][324] ) );
  ANDN U268 ( .B(zreg[323]), .A(start), .Z(\zin[0][323] ) );
  ANDN U269 ( .B(zreg[322]), .A(start), .Z(\zin[0][322] ) );
  ANDN U270 ( .B(zreg[321]), .A(start), .Z(\zin[0][321] ) );
  ANDN U271 ( .B(zreg[320]), .A(start), .Z(\zin[0][320] ) );
  ANDN U272 ( .B(zreg[31]), .A(start), .Z(\zin[0][31] ) );
  ANDN U273 ( .B(zreg[319]), .A(start), .Z(\zin[0][319] ) );
  ANDN U274 ( .B(zreg[318]), .A(start), .Z(\zin[0][318] ) );
  ANDN U275 ( .B(zreg[317]), .A(start), .Z(\zin[0][317] ) );
  ANDN U276 ( .B(zreg[316]), .A(start), .Z(\zin[0][316] ) );
  ANDN U277 ( .B(zreg[315]), .A(start), .Z(\zin[0][315] ) );
  ANDN U278 ( .B(zreg[314]), .A(start), .Z(\zin[0][314] ) );
  ANDN U279 ( .B(zreg[313]), .A(start), .Z(\zin[0][313] ) );
  ANDN U280 ( .B(zreg[312]), .A(start), .Z(\zin[0][312] ) );
  ANDN U281 ( .B(zreg[311]), .A(start), .Z(\zin[0][311] ) );
  ANDN U282 ( .B(zreg[310]), .A(start), .Z(\zin[0][310] ) );
  ANDN U283 ( .B(zreg[30]), .A(start), .Z(\zin[0][30] ) );
  ANDN U284 ( .B(zreg[309]), .A(start), .Z(\zin[0][309] ) );
  ANDN U285 ( .B(zreg[308]), .A(start), .Z(\zin[0][308] ) );
  ANDN U286 ( .B(zreg[307]), .A(start), .Z(\zin[0][307] ) );
  ANDN U287 ( .B(zreg[306]), .A(start), .Z(\zin[0][306] ) );
  ANDN U288 ( .B(zreg[305]), .A(start), .Z(\zin[0][305] ) );
  ANDN U289 ( .B(zreg[304]), .A(start), .Z(\zin[0][304] ) );
  ANDN U290 ( .B(zreg[303]), .A(start), .Z(\zin[0][303] ) );
  ANDN U291 ( .B(zreg[302]), .A(start), .Z(\zin[0][302] ) );
  ANDN U292 ( .B(zreg[301]), .A(start), .Z(\zin[0][301] ) );
  ANDN U293 ( .B(zreg[300]), .A(start), .Z(\zin[0][300] ) );
  ANDN U294 ( .B(zreg[2]), .A(start), .Z(\zin[0][2] ) );
  ANDN U295 ( .B(zreg[29]), .A(start), .Z(\zin[0][29] ) );
  ANDN U296 ( .B(zreg[299]), .A(start), .Z(\zin[0][299] ) );
  ANDN U297 ( .B(zreg[298]), .A(start), .Z(\zin[0][298] ) );
  ANDN U298 ( .B(zreg[297]), .A(start), .Z(\zin[0][297] ) );
  ANDN U299 ( .B(zreg[296]), .A(start), .Z(\zin[0][296] ) );
  ANDN U300 ( .B(zreg[295]), .A(start), .Z(\zin[0][295] ) );
  ANDN U301 ( .B(zreg[294]), .A(start), .Z(\zin[0][294] ) );
  ANDN U302 ( .B(zreg[293]), .A(start), .Z(\zin[0][293] ) );
  ANDN U303 ( .B(zreg[292]), .A(start), .Z(\zin[0][292] ) );
  ANDN U304 ( .B(zreg[291]), .A(start), .Z(\zin[0][291] ) );
  ANDN U305 ( .B(zreg[290]), .A(start), .Z(\zin[0][290] ) );
  ANDN U306 ( .B(zreg[28]), .A(start), .Z(\zin[0][28] ) );
  ANDN U307 ( .B(zreg[289]), .A(start), .Z(\zin[0][289] ) );
  ANDN U308 ( .B(zreg[288]), .A(start), .Z(\zin[0][288] ) );
  ANDN U309 ( .B(zreg[287]), .A(start), .Z(\zin[0][287] ) );
  ANDN U310 ( .B(zreg[286]), .A(start), .Z(\zin[0][286] ) );
  ANDN U311 ( .B(zreg[285]), .A(start), .Z(\zin[0][285] ) );
  ANDN U312 ( .B(zreg[284]), .A(start), .Z(\zin[0][284] ) );
  ANDN U313 ( .B(zreg[283]), .A(start), .Z(\zin[0][283] ) );
  ANDN U314 ( .B(zreg[282]), .A(start), .Z(\zin[0][282] ) );
  ANDN U315 ( .B(zreg[281]), .A(start), .Z(\zin[0][281] ) );
  ANDN U316 ( .B(zreg[280]), .A(start), .Z(\zin[0][280] ) );
  ANDN U317 ( .B(zreg[27]), .A(start), .Z(\zin[0][27] ) );
  ANDN U318 ( .B(zreg[279]), .A(start), .Z(\zin[0][279] ) );
  ANDN U319 ( .B(zreg[278]), .A(start), .Z(\zin[0][278] ) );
  ANDN U320 ( .B(zreg[277]), .A(start), .Z(\zin[0][277] ) );
  ANDN U321 ( .B(zreg[276]), .A(start), .Z(\zin[0][276] ) );
  ANDN U322 ( .B(zreg[275]), .A(start), .Z(\zin[0][275] ) );
  ANDN U323 ( .B(zreg[274]), .A(start), .Z(\zin[0][274] ) );
  ANDN U324 ( .B(zreg[273]), .A(start), .Z(\zin[0][273] ) );
  ANDN U325 ( .B(zreg[272]), .A(start), .Z(\zin[0][272] ) );
  ANDN U326 ( .B(zreg[271]), .A(start), .Z(\zin[0][271] ) );
  ANDN U327 ( .B(zreg[270]), .A(start), .Z(\zin[0][270] ) );
  ANDN U328 ( .B(zreg[26]), .A(start), .Z(\zin[0][26] ) );
  ANDN U329 ( .B(zreg[269]), .A(start), .Z(\zin[0][269] ) );
  ANDN U330 ( .B(zreg[268]), .A(start), .Z(\zin[0][268] ) );
  ANDN U331 ( .B(zreg[267]), .A(start), .Z(\zin[0][267] ) );
  ANDN U332 ( .B(zreg[266]), .A(start), .Z(\zin[0][266] ) );
  ANDN U333 ( .B(zreg[265]), .A(start), .Z(\zin[0][265] ) );
  ANDN U334 ( .B(zreg[264]), .A(start), .Z(\zin[0][264] ) );
  ANDN U335 ( .B(zreg[263]), .A(start), .Z(\zin[0][263] ) );
  ANDN U336 ( .B(zreg[262]), .A(start), .Z(\zin[0][262] ) );
  ANDN U337 ( .B(zreg[261]), .A(start), .Z(\zin[0][261] ) );
  ANDN U338 ( .B(zreg[260]), .A(start), .Z(\zin[0][260] ) );
  ANDN U339 ( .B(zreg[25]), .A(start), .Z(\zin[0][25] ) );
  ANDN U340 ( .B(zreg[259]), .A(start), .Z(\zin[0][259] ) );
  ANDN U341 ( .B(zreg[258]), .A(start), .Z(\zin[0][258] ) );
  ANDN U342 ( .B(zreg[257]), .A(start), .Z(\zin[0][257] ) );
  ANDN U343 ( .B(zreg[256]), .A(start), .Z(\zin[0][256] ) );
  ANDN U344 ( .B(zreg[255]), .A(start), .Z(\zin[0][255] ) );
  ANDN U345 ( .B(zreg[254]), .A(start), .Z(\zin[0][254] ) );
  ANDN U346 ( .B(zreg[253]), .A(start), .Z(\zin[0][253] ) );
  ANDN U347 ( .B(zreg[252]), .A(start), .Z(\zin[0][252] ) );
  ANDN U348 ( .B(zreg[251]), .A(start), .Z(\zin[0][251] ) );
  ANDN U349 ( .B(zreg[250]), .A(start), .Z(\zin[0][250] ) );
  ANDN U350 ( .B(zreg[24]), .A(start), .Z(\zin[0][24] ) );
  ANDN U351 ( .B(zreg[249]), .A(start), .Z(\zin[0][249] ) );
  ANDN U352 ( .B(zreg[248]), .A(start), .Z(\zin[0][248] ) );
  ANDN U353 ( .B(zreg[247]), .A(start), .Z(\zin[0][247] ) );
  ANDN U354 ( .B(zreg[246]), .A(start), .Z(\zin[0][246] ) );
  ANDN U355 ( .B(zreg[245]), .A(start), .Z(\zin[0][245] ) );
  ANDN U356 ( .B(zreg[244]), .A(start), .Z(\zin[0][244] ) );
  ANDN U357 ( .B(zreg[243]), .A(start), .Z(\zin[0][243] ) );
  ANDN U358 ( .B(zreg[242]), .A(start), .Z(\zin[0][242] ) );
  ANDN U359 ( .B(zreg[241]), .A(start), .Z(\zin[0][241] ) );
  ANDN U360 ( .B(zreg[240]), .A(start), .Z(\zin[0][240] ) );
  ANDN U361 ( .B(zreg[23]), .A(start), .Z(\zin[0][23] ) );
  ANDN U362 ( .B(zreg[239]), .A(start), .Z(\zin[0][239] ) );
  ANDN U363 ( .B(zreg[238]), .A(start), .Z(\zin[0][238] ) );
  ANDN U364 ( .B(zreg[237]), .A(start), .Z(\zin[0][237] ) );
  ANDN U365 ( .B(zreg[236]), .A(start), .Z(\zin[0][236] ) );
  ANDN U366 ( .B(zreg[235]), .A(start), .Z(\zin[0][235] ) );
  ANDN U367 ( .B(zreg[234]), .A(start), .Z(\zin[0][234] ) );
  ANDN U368 ( .B(zreg[233]), .A(start), .Z(\zin[0][233] ) );
  ANDN U369 ( .B(zreg[232]), .A(start), .Z(\zin[0][232] ) );
  ANDN U370 ( .B(zreg[231]), .A(start), .Z(\zin[0][231] ) );
  ANDN U371 ( .B(zreg[230]), .A(start), .Z(\zin[0][230] ) );
  ANDN U372 ( .B(zreg[22]), .A(start), .Z(\zin[0][22] ) );
  ANDN U373 ( .B(zreg[229]), .A(start), .Z(\zin[0][229] ) );
  ANDN U374 ( .B(zreg[228]), .A(start), .Z(\zin[0][228] ) );
  ANDN U375 ( .B(zreg[227]), .A(start), .Z(\zin[0][227] ) );
  ANDN U376 ( .B(zreg[226]), .A(start), .Z(\zin[0][226] ) );
  ANDN U377 ( .B(zreg[225]), .A(start), .Z(\zin[0][225] ) );
  ANDN U378 ( .B(zreg[224]), .A(start), .Z(\zin[0][224] ) );
  ANDN U379 ( .B(zreg[223]), .A(start), .Z(\zin[0][223] ) );
  ANDN U380 ( .B(zreg[222]), .A(start), .Z(\zin[0][222] ) );
  ANDN U381 ( .B(zreg[221]), .A(start), .Z(\zin[0][221] ) );
  ANDN U382 ( .B(zreg[220]), .A(start), .Z(\zin[0][220] ) );
  ANDN U383 ( .B(zreg[21]), .A(start), .Z(\zin[0][21] ) );
  ANDN U384 ( .B(zreg[219]), .A(start), .Z(\zin[0][219] ) );
  ANDN U385 ( .B(zreg[218]), .A(start), .Z(\zin[0][218] ) );
  ANDN U386 ( .B(zreg[217]), .A(start), .Z(\zin[0][217] ) );
  ANDN U387 ( .B(zreg[216]), .A(start), .Z(\zin[0][216] ) );
  ANDN U388 ( .B(zreg[215]), .A(start), .Z(\zin[0][215] ) );
  ANDN U389 ( .B(zreg[214]), .A(start), .Z(\zin[0][214] ) );
  ANDN U390 ( .B(zreg[213]), .A(start), .Z(\zin[0][213] ) );
  ANDN U391 ( .B(zreg[212]), .A(start), .Z(\zin[0][212] ) );
  ANDN U392 ( .B(zreg[211]), .A(start), .Z(\zin[0][211] ) );
  ANDN U393 ( .B(zreg[210]), .A(start), .Z(\zin[0][210] ) );
  ANDN U394 ( .B(zreg[20]), .A(start), .Z(\zin[0][20] ) );
  ANDN U395 ( .B(zreg[209]), .A(start), .Z(\zin[0][209] ) );
  ANDN U396 ( .B(zreg[208]), .A(start), .Z(\zin[0][208] ) );
  ANDN U397 ( .B(zreg[207]), .A(start), .Z(\zin[0][207] ) );
  ANDN U398 ( .B(zreg[206]), .A(start), .Z(\zin[0][206] ) );
  ANDN U399 ( .B(zreg[205]), .A(start), .Z(\zin[0][205] ) );
  ANDN U400 ( .B(zreg[204]), .A(start), .Z(\zin[0][204] ) );
  ANDN U401 ( .B(zreg[203]), .A(start), .Z(\zin[0][203] ) );
  ANDN U402 ( .B(zreg[202]), .A(start), .Z(\zin[0][202] ) );
  ANDN U403 ( .B(zreg[201]), .A(start), .Z(\zin[0][201] ) );
  ANDN U404 ( .B(zreg[200]), .A(start), .Z(\zin[0][200] ) );
  ANDN U405 ( .B(zreg[1]), .A(start), .Z(\zin[0][1] ) );
  ANDN U406 ( .B(zreg[19]), .A(start), .Z(\zin[0][19] ) );
  ANDN U407 ( .B(zreg[199]), .A(start), .Z(\zin[0][199] ) );
  ANDN U408 ( .B(zreg[198]), .A(start), .Z(\zin[0][198] ) );
  ANDN U409 ( .B(zreg[197]), .A(start), .Z(\zin[0][197] ) );
  ANDN U410 ( .B(zreg[196]), .A(start), .Z(\zin[0][196] ) );
  ANDN U411 ( .B(zreg[195]), .A(start), .Z(\zin[0][195] ) );
  ANDN U412 ( .B(zreg[194]), .A(start), .Z(\zin[0][194] ) );
  ANDN U413 ( .B(zreg[193]), .A(start), .Z(\zin[0][193] ) );
  ANDN U414 ( .B(zreg[192]), .A(start), .Z(\zin[0][192] ) );
  ANDN U415 ( .B(zreg[191]), .A(start), .Z(\zin[0][191] ) );
  ANDN U416 ( .B(zreg[190]), .A(start), .Z(\zin[0][190] ) );
  ANDN U417 ( .B(zreg[18]), .A(start), .Z(\zin[0][18] ) );
  ANDN U418 ( .B(zreg[189]), .A(start), .Z(\zin[0][189] ) );
  ANDN U419 ( .B(zreg[188]), .A(start), .Z(\zin[0][188] ) );
  ANDN U420 ( .B(zreg[187]), .A(start), .Z(\zin[0][187] ) );
  ANDN U421 ( .B(zreg[186]), .A(start), .Z(\zin[0][186] ) );
  ANDN U422 ( .B(zreg[185]), .A(start), .Z(\zin[0][185] ) );
  ANDN U423 ( .B(zreg[184]), .A(start), .Z(\zin[0][184] ) );
  ANDN U424 ( .B(zreg[183]), .A(start), .Z(\zin[0][183] ) );
  ANDN U425 ( .B(zreg[182]), .A(start), .Z(\zin[0][182] ) );
  ANDN U426 ( .B(zreg[181]), .A(start), .Z(\zin[0][181] ) );
  ANDN U427 ( .B(zreg[180]), .A(start), .Z(\zin[0][180] ) );
  ANDN U428 ( .B(zreg[17]), .A(start), .Z(\zin[0][17] ) );
  ANDN U429 ( .B(zreg[179]), .A(start), .Z(\zin[0][179] ) );
  ANDN U430 ( .B(zreg[178]), .A(start), .Z(\zin[0][178] ) );
  ANDN U431 ( .B(zreg[177]), .A(start), .Z(\zin[0][177] ) );
  ANDN U432 ( .B(zreg[176]), .A(start), .Z(\zin[0][176] ) );
  ANDN U433 ( .B(zreg[175]), .A(start), .Z(\zin[0][175] ) );
  ANDN U434 ( .B(zreg[174]), .A(start), .Z(\zin[0][174] ) );
  ANDN U435 ( .B(zreg[173]), .A(start), .Z(\zin[0][173] ) );
  ANDN U436 ( .B(zreg[172]), .A(start), .Z(\zin[0][172] ) );
  ANDN U437 ( .B(zreg[171]), .A(start), .Z(\zin[0][171] ) );
  ANDN U438 ( .B(zreg[170]), .A(start), .Z(\zin[0][170] ) );
  ANDN U439 ( .B(zreg[16]), .A(start), .Z(\zin[0][16] ) );
  ANDN U440 ( .B(zreg[169]), .A(start), .Z(\zin[0][169] ) );
  ANDN U441 ( .B(zreg[168]), .A(start), .Z(\zin[0][168] ) );
  ANDN U442 ( .B(zreg[167]), .A(start), .Z(\zin[0][167] ) );
  ANDN U443 ( .B(zreg[166]), .A(start), .Z(\zin[0][166] ) );
  ANDN U444 ( .B(zreg[165]), .A(start), .Z(\zin[0][165] ) );
  ANDN U445 ( .B(zreg[164]), .A(start), .Z(\zin[0][164] ) );
  ANDN U446 ( .B(zreg[163]), .A(start), .Z(\zin[0][163] ) );
  ANDN U447 ( .B(zreg[162]), .A(start), .Z(\zin[0][162] ) );
  ANDN U448 ( .B(zreg[161]), .A(start), .Z(\zin[0][161] ) );
  ANDN U449 ( .B(zreg[160]), .A(start), .Z(\zin[0][160] ) );
  ANDN U450 ( .B(zreg[15]), .A(start), .Z(\zin[0][15] ) );
  ANDN U451 ( .B(zreg[159]), .A(start), .Z(\zin[0][159] ) );
  ANDN U452 ( .B(zreg[158]), .A(start), .Z(\zin[0][158] ) );
  ANDN U453 ( .B(zreg[157]), .A(start), .Z(\zin[0][157] ) );
  ANDN U454 ( .B(zreg[156]), .A(start), .Z(\zin[0][156] ) );
  ANDN U455 ( .B(zreg[155]), .A(start), .Z(\zin[0][155] ) );
  ANDN U456 ( .B(zreg[154]), .A(start), .Z(\zin[0][154] ) );
  ANDN U457 ( .B(zreg[153]), .A(start), .Z(\zin[0][153] ) );
  ANDN U458 ( .B(zreg[152]), .A(start), .Z(\zin[0][152] ) );
  ANDN U459 ( .B(zreg[151]), .A(start), .Z(\zin[0][151] ) );
  ANDN U460 ( .B(zreg[150]), .A(start), .Z(\zin[0][150] ) );
  ANDN U461 ( .B(zreg[14]), .A(start), .Z(\zin[0][14] ) );
  ANDN U462 ( .B(zreg[149]), .A(start), .Z(\zin[0][149] ) );
  ANDN U463 ( .B(zreg[148]), .A(start), .Z(\zin[0][148] ) );
  ANDN U464 ( .B(zreg[147]), .A(start), .Z(\zin[0][147] ) );
  ANDN U465 ( .B(zreg[146]), .A(start), .Z(\zin[0][146] ) );
  ANDN U466 ( .B(zreg[145]), .A(start), .Z(\zin[0][145] ) );
  ANDN U467 ( .B(zreg[144]), .A(start), .Z(\zin[0][144] ) );
  ANDN U468 ( .B(zreg[143]), .A(start), .Z(\zin[0][143] ) );
  ANDN U469 ( .B(zreg[142]), .A(start), .Z(\zin[0][142] ) );
  ANDN U470 ( .B(zreg[141]), .A(start), .Z(\zin[0][141] ) );
  ANDN U471 ( .B(zreg[140]), .A(start), .Z(\zin[0][140] ) );
  ANDN U472 ( .B(zreg[13]), .A(start), .Z(\zin[0][13] ) );
  ANDN U473 ( .B(zreg[139]), .A(start), .Z(\zin[0][139] ) );
  ANDN U474 ( .B(zreg[138]), .A(start), .Z(\zin[0][138] ) );
  ANDN U475 ( .B(zreg[137]), .A(start), .Z(\zin[0][137] ) );
  ANDN U476 ( .B(zreg[136]), .A(start), .Z(\zin[0][136] ) );
  ANDN U477 ( .B(zreg[135]), .A(start), .Z(\zin[0][135] ) );
  ANDN U478 ( .B(zreg[134]), .A(start), .Z(\zin[0][134] ) );
  ANDN U479 ( .B(zreg[133]), .A(start), .Z(\zin[0][133] ) );
  ANDN U480 ( .B(zreg[132]), .A(start), .Z(\zin[0][132] ) );
  ANDN U481 ( .B(zreg[131]), .A(start), .Z(\zin[0][131] ) );
  ANDN U482 ( .B(zreg[130]), .A(start), .Z(\zin[0][130] ) );
  ANDN U483 ( .B(zreg[12]), .A(start), .Z(\zin[0][12] ) );
  ANDN U484 ( .B(zreg[129]), .A(start), .Z(\zin[0][129] ) );
  ANDN U485 ( .B(zreg[128]), .A(start), .Z(\zin[0][128] ) );
  ANDN U486 ( .B(zreg[127]), .A(start), .Z(\zin[0][127] ) );
  ANDN U487 ( .B(zreg[126]), .A(start), .Z(\zin[0][126] ) );
  ANDN U488 ( .B(zreg[125]), .A(start), .Z(\zin[0][125] ) );
  ANDN U489 ( .B(zreg[124]), .A(start), .Z(\zin[0][124] ) );
  ANDN U490 ( .B(zreg[123]), .A(start), .Z(\zin[0][123] ) );
  ANDN U491 ( .B(zreg[122]), .A(start), .Z(\zin[0][122] ) );
  ANDN U492 ( .B(zreg[121]), .A(start), .Z(\zin[0][121] ) );
  ANDN U493 ( .B(zreg[120]), .A(start), .Z(\zin[0][120] ) );
  ANDN U494 ( .B(zreg[11]), .A(start), .Z(\zin[0][11] ) );
  ANDN U495 ( .B(zreg[119]), .A(start), .Z(\zin[0][119] ) );
  ANDN U496 ( .B(zreg[118]), .A(start), .Z(\zin[0][118] ) );
  ANDN U497 ( .B(zreg[117]), .A(start), .Z(\zin[0][117] ) );
  ANDN U498 ( .B(zreg[116]), .A(start), .Z(\zin[0][116] ) );
  ANDN U499 ( .B(zreg[115]), .A(start), .Z(\zin[0][115] ) );
  ANDN U500 ( .B(zreg[114]), .A(start), .Z(\zin[0][114] ) );
  ANDN U501 ( .B(zreg[113]), .A(start), .Z(\zin[0][113] ) );
  ANDN U502 ( .B(zreg[112]), .A(start), .Z(\zin[0][112] ) );
  ANDN U503 ( .B(zreg[111]), .A(start), .Z(\zin[0][111] ) );
  ANDN U504 ( .B(zreg[110]), .A(start), .Z(\zin[0][110] ) );
  ANDN U505 ( .B(zreg[10]), .A(start), .Z(\zin[0][10] ) );
  ANDN U506 ( .B(zreg[109]), .A(start), .Z(\zin[0][109] ) );
  ANDN U507 ( .B(zreg[108]), .A(start), .Z(\zin[0][108] ) );
  ANDN U508 ( .B(zreg[107]), .A(start), .Z(\zin[0][107] ) );
  ANDN U509 ( .B(zreg[106]), .A(start), .Z(\zin[0][106] ) );
  ANDN U510 ( .B(zreg[105]), .A(start), .Z(\zin[0][105] ) );
  ANDN U511 ( .B(zreg[104]), .A(start), .Z(\zin[0][104] ) );
  ANDN U512 ( .B(zreg[103]), .A(start), .Z(\zin[0][103] ) );
  ANDN U513 ( .B(zreg[102]), .A(start), .Z(\zin[0][102] ) );
  ANDN U514 ( .B(zreg[101]), .A(start), .Z(\zin[0][101] ) );
  ANDN U515 ( .B(zreg[100]), .A(start), .Z(\zin[0][100] ) );
  ANDN U516 ( .B(zreg[0]), .A(start), .Z(\zin[0][0] ) );
  NAND U517 ( .A(n1), .B(n2), .Z(xin[9]) );
  NANDN U518 ( .A(start), .B(xreg[9]), .Z(n2) );
  NAND U519 ( .A(x[9]), .B(start), .Z(n1) );
  NAND U520 ( .A(n3), .B(n4), .Z(xin[99]) );
  NANDN U521 ( .A(start), .B(xreg[99]), .Z(n4) );
  NAND U522 ( .A(x[99]), .B(start), .Z(n3) );
  NAND U523 ( .A(n5), .B(n6), .Z(xin[98]) );
  NANDN U524 ( .A(start), .B(xreg[98]), .Z(n6) );
  NAND U525 ( .A(x[98]), .B(start), .Z(n5) );
  NAND U526 ( .A(n7), .B(n8), .Z(xin[97]) );
  NANDN U527 ( .A(start), .B(xreg[97]), .Z(n8) );
  NAND U528 ( .A(x[97]), .B(start), .Z(n7) );
  NAND U529 ( .A(n9), .B(n10), .Z(xin[96]) );
  NANDN U530 ( .A(start), .B(xreg[96]), .Z(n10) );
  NAND U531 ( .A(x[96]), .B(start), .Z(n9) );
  NAND U532 ( .A(n11), .B(n12), .Z(xin[95]) );
  NANDN U533 ( .A(start), .B(xreg[95]), .Z(n12) );
  NAND U534 ( .A(x[95]), .B(start), .Z(n11) );
  NAND U535 ( .A(n13), .B(n14), .Z(xin[94]) );
  NANDN U536 ( .A(start), .B(xreg[94]), .Z(n14) );
  NAND U537 ( .A(x[94]), .B(start), .Z(n13) );
  NAND U538 ( .A(n15), .B(n16), .Z(xin[93]) );
  NANDN U539 ( .A(start), .B(xreg[93]), .Z(n16) );
  NAND U540 ( .A(x[93]), .B(start), .Z(n15) );
  NAND U541 ( .A(n17), .B(n18), .Z(xin[92]) );
  NANDN U542 ( .A(start), .B(xreg[92]), .Z(n18) );
  NAND U543 ( .A(x[92]), .B(start), .Z(n17) );
  NAND U544 ( .A(n19), .B(n20), .Z(xin[91]) );
  NANDN U545 ( .A(start), .B(xreg[91]), .Z(n20) );
  NAND U546 ( .A(x[91]), .B(start), .Z(n19) );
  NAND U547 ( .A(n21), .B(n22), .Z(xin[90]) );
  NANDN U548 ( .A(start), .B(xreg[90]), .Z(n22) );
  NAND U549 ( .A(x[90]), .B(start), .Z(n21) );
  NAND U550 ( .A(n23), .B(n24), .Z(xin[8]) );
  NANDN U551 ( .A(start), .B(xreg[8]), .Z(n24) );
  NAND U552 ( .A(x[8]), .B(start), .Z(n23) );
  NAND U553 ( .A(n25), .B(n26), .Z(xin[89]) );
  NANDN U554 ( .A(start), .B(xreg[89]), .Z(n26) );
  NAND U555 ( .A(x[89]), .B(start), .Z(n25) );
  NAND U556 ( .A(n27), .B(n28), .Z(xin[88]) );
  NANDN U557 ( .A(start), .B(xreg[88]), .Z(n28) );
  NAND U558 ( .A(x[88]), .B(start), .Z(n27) );
  NAND U559 ( .A(n29), .B(n30), .Z(xin[87]) );
  NANDN U560 ( .A(start), .B(xreg[87]), .Z(n30) );
  NAND U561 ( .A(x[87]), .B(start), .Z(n29) );
  NAND U562 ( .A(n31), .B(n32), .Z(xin[86]) );
  NANDN U563 ( .A(start), .B(xreg[86]), .Z(n32) );
  NAND U564 ( .A(x[86]), .B(start), .Z(n31) );
  NAND U565 ( .A(n33), .B(n34), .Z(xin[85]) );
  NANDN U566 ( .A(start), .B(xreg[85]), .Z(n34) );
  NAND U567 ( .A(x[85]), .B(start), .Z(n33) );
  NAND U568 ( .A(n35), .B(n36), .Z(xin[84]) );
  NANDN U569 ( .A(start), .B(xreg[84]), .Z(n36) );
  NAND U570 ( .A(x[84]), .B(start), .Z(n35) );
  NAND U571 ( .A(n37), .B(n38), .Z(xin[83]) );
  NANDN U572 ( .A(start), .B(xreg[83]), .Z(n38) );
  NAND U573 ( .A(x[83]), .B(start), .Z(n37) );
  NAND U574 ( .A(n39), .B(n40), .Z(xin[82]) );
  NANDN U575 ( .A(start), .B(xreg[82]), .Z(n40) );
  NAND U576 ( .A(x[82]), .B(start), .Z(n39) );
  NAND U577 ( .A(n41), .B(n42), .Z(xin[81]) );
  NANDN U578 ( .A(start), .B(xreg[81]), .Z(n42) );
  NAND U579 ( .A(x[81]), .B(start), .Z(n41) );
  NAND U580 ( .A(n43), .B(n44), .Z(xin[80]) );
  NANDN U581 ( .A(start), .B(xreg[80]), .Z(n44) );
  NAND U582 ( .A(x[80]), .B(start), .Z(n43) );
  NAND U583 ( .A(n45), .B(n46), .Z(xin[7]) );
  NANDN U584 ( .A(start), .B(xreg[7]), .Z(n46) );
  NAND U585 ( .A(x[7]), .B(start), .Z(n45) );
  NAND U586 ( .A(n47), .B(n48), .Z(xin[79]) );
  NANDN U587 ( .A(start), .B(xreg[79]), .Z(n48) );
  NAND U588 ( .A(x[79]), .B(start), .Z(n47) );
  NAND U589 ( .A(n49), .B(n50), .Z(xin[78]) );
  NANDN U590 ( .A(start), .B(xreg[78]), .Z(n50) );
  NAND U591 ( .A(x[78]), .B(start), .Z(n49) );
  NAND U592 ( .A(n51), .B(n52), .Z(xin[77]) );
  NANDN U593 ( .A(start), .B(xreg[77]), .Z(n52) );
  NAND U594 ( .A(x[77]), .B(start), .Z(n51) );
  NAND U595 ( .A(n53), .B(n54), .Z(xin[76]) );
  NANDN U596 ( .A(start), .B(xreg[76]), .Z(n54) );
  NAND U597 ( .A(x[76]), .B(start), .Z(n53) );
  NAND U598 ( .A(n55), .B(n56), .Z(xin[75]) );
  NANDN U599 ( .A(start), .B(xreg[75]), .Z(n56) );
  NAND U600 ( .A(x[75]), .B(start), .Z(n55) );
  NAND U601 ( .A(n57), .B(n58), .Z(xin[74]) );
  NANDN U602 ( .A(start), .B(xreg[74]), .Z(n58) );
  NAND U603 ( .A(x[74]), .B(start), .Z(n57) );
  NAND U604 ( .A(n59), .B(n60), .Z(xin[73]) );
  NANDN U605 ( .A(start), .B(xreg[73]), .Z(n60) );
  NAND U606 ( .A(x[73]), .B(start), .Z(n59) );
  NAND U607 ( .A(n61), .B(n62), .Z(xin[72]) );
  NANDN U608 ( .A(start), .B(xreg[72]), .Z(n62) );
  NAND U609 ( .A(x[72]), .B(start), .Z(n61) );
  NAND U610 ( .A(n63), .B(n64), .Z(xin[71]) );
  NANDN U611 ( .A(start), .B(xreg[71]), .Z(n64) );
  NAND U612 ( .A(x[71]), .B(start), .Z(n63) );
  NAND U613 ( .A(n65), .B(n66), .Z(xin[70]) );
  NANDN U614 ( .A(start), .B(xreg[70]), .Z(n66) );
  NAND U615 ( .A(x[70]), .B(start), .Z(n65) );
  NAND U616 ( .A(n67), .B(n68), .Z(xin[6]) );
  NANDN U617 ( .A(start), .B(xreg[6]), .Z(n68) );
  NAND U618 ( .A(x[6]), .B(start), .Z(n67) );
  NAND U619 ( .A(n69), .B(n70), .Z(xin[69]) );
  NANDN U620 ( .A(start), .B(xreg[69]), .Z(n70) );
  NAND U621 ( .A(x[69]), .B(start), .Z(n69) );
  NAND U622 ( .A(n71), .B(n72), .Z(xin[68]) );
  NANDN U623 ( .A(start), .B(xreg[68]), .Z(n72) );
  NAND U624 ( .A(x[68]), .B(start), .Z(n71) );
  NAND U625 ( .A(n73), .B(n74), .Z(xin[67]) );
  NANDN U626 ( .A(start), .B(xreg[67]), .Z(n74) );
  NAND U627 ( .A(x[67]), .B(start), .Z(n73) );
  NAND U628 ( .A(n75), .B(n76), .Z(xin[66]) );
  NANDN U629 ( .A(start), .B(xreg[66]), .Z(n76) );
  NAND U630 ( .A(x[66]), .B(start), .Z(n75) );
  NAND U631 ( .A(n77), .B(n78), .Z(xin[65]) );
  NANDN U632 ( .A(start), .B(xreg[65]), .Z(n78) );
  NAND U633 ( .A(x[65]), .B(start), .Z(n77) );
  NAND U634 ( .A(n79), .B(n80), .Z(xin[64]) );
  NANDN U635 ( .A(start), .B(xreg[64]), .Z(n80) );
  NAND U636 ( .A(x[64]), .B(start), .Z(n79) );
  NAND U637 ( .A(n81), .B(n82), .Z(xin[63]) );
  NANDN U638 ( .A(start), .B(xreg[63]), .Z(n82) );
  NAND U639 ( .A(x[63]), .B(start), .Z(n81) );
  NAND U640 ( .A(n83), .B(n84), .Z(xin[62]) );
  NANDN U641 ( .A(start), .B(xreg[62]), .Z(n84) );
  NAND U642 ( .A(x[62]), .B(start), .Z(n83) );
  NAND U643 ( .A(n85), .B(n86), .Z(xin[61]) );
  NANDN U644 ( .A(start), .B(xreg[61]), .Z(n86) );
  NAND U645 ( .A(x[61]), .B(start), .Z(n85) );
  NAND U646 ( .A(n87), .B(n88), .Z(xin[60]) );
  NANDN U647 ( .A(start), .B(xreg[60]), .Z(n88) );
  NAND U648 ( .A(x[60]), .B(start), .Z(n87) );
  NAND U649 ( .A(n89), .B(n90), .Z(xin[5]) );
  NANDN U650 ( .A(start), .B(xreg[5]), .Z(n90) );
  NAND U651 ( .A(x[5]), .B(start), .Z(n89) );
  NAND U652 ( .A(n91), .B(n92), .Z(xin[59]) );
  NANDN U653 ( .A(start), .B(xreg[59]), .Z(n92) );
  NAND U654 ( .A(x[59]), .B(start), .Z(n91) );
  NAND U655 ( .A(n93), .B(n94), .Z(xin[58]) );
  NANDN U656 ( .A(start), .B(xreg[58]), .Z(n94) );
  NAND U657 ( .A(x[58]), .B(start), .Z(n93) );
  NAND U658 ( .A(n95), .B(n96), .Z(xin[57]) );
  NANDN U659 ( .A(start), .B(xreg[57]), .Z(n96) );
  NAND U660 ( .A(x[57]), .B(start), .Z(n95) );
  NAND U661 ( .A(n97), .B(n98), .Z(xin[56]) );
  NANDN U662 ( .A(start), .B(xreg[56]), .Z(n98) );
  NAND U663 ( .A(x[56]), .B(start), .Z(n97) );
  NAND U664 ( .A(n99), .B(n100), .Z(xin[55]) );
  NANDN U665 ( .A(start), .B(xreg[55]), .Z(n100) );
  NAND U666 ( .A(x[55]), .B(start), .Z(n99) );
  NAND U667 ( .A(n101), .B(n102), .Z(xin[54]) );
  NANDN U668 ( .A(start), .B(xreg[54]), .Z(n102) );
  NAND U669 ( .A(x[54]), .B(start), .Z(n101) );
  NAND U670 ( .A(n103), .B(n104), .Z(xin[53]) );
  NANDN U671 ( .A(start), .B(xreg[53]), .Z(n104) );
  NAND U672 ( .A(x[53]), .B(start), .Z(n103) );
  NAND U673 ( .A(n105), .B(n106), .Z(xin[52]) );
  NANDN U674 ( .A(start), .B(xreg[52]), .Z(n106) );
  NAND U675 ( .A(x[52]), .B(start), .Z(n105) );
  NAND U676 ( .A(n107), .B(n108), .Z(xin[51]) );
  NANDN U677 ( .A(start), .B(xreg[51]), .Z(n108) );
  NAND U678 ( .A(x[51]), .B(start), .Z(n107) );
  NAND U679 ( .A(n109), .B(n110), .Z(xin[511]) );
  NANDN U680 ( .A(start), .B(xreg[511]), .Z(n110) );
  NAND U681 ( .A(x[511]), .B(start), .Z(n109) );
  NAND U682 ( .A(n111), .B(n112), .Z(xin[510]) );
  NANDN U683 ( .A(start), .B(xreg[510]), .Z(n112) );
  NAND U684 ( .A(x[510]), .B(start), .Z(n111) );
  NAND U685 ( .A(n113), .B(n114), .Z(xin[50]) );
  NANDN U686 ( .A(start), .B(xreg[50]), .Z(n114) );
  NAND U687 ( .A(x[50]), .B(start), .Z(n113) );
  NAND U688 ( .A(n115), .B(n116), .Z(xin[509]) );
  NANDN U689 ( .A(start), .B(xreg[509]), .Z(n116) );
  NAND U690 ( .A(x[509]), .B(start), .Z(n115) );
  NAND U691 ( .A(n117), .B(n118), .Z(xin[508]) );
  NANDN U692 ( .A(start), .B(xreg[508]), .Z(n118) );
  NAND U693 ( .A(x[508]), .B(start), .Z(n117) );
  NAND U694 ( .A(n119), .B(n120), .Z(xin[507]) );
  NANDN U695 ( .A(start), .B(xreg[507]), .Z(n120) );
  NAND U696 ( .A(x[507]), .B(start), .Z(n119) );
  NAND U697 ( .A(n121), .B(n122), .Z(xin[506]) );
  NANDN U698 ( .A(start), .B(xreg[506]), .Z(n122) );
  NAND U699 ( .A(x[506]), .B(start), .Z(n121) );
  NAND U700 ( .A(n123), .B(n124), .Z(xin[505]) );
  NANDN U701 ( .A(start), .B(xreg[505]), .Z(n124) );
  NAND U702 ( .A(x[505]), .B(start), .Z(n123) );
  NAND U703 ( .A(n125), .B(n126), .Z(xin[504]) );
  NANDN U704 ( .A(start), .B(xreg[504]), .Z(n126) );
  NAND U705 ( .A(x[504]), .B(start), .Z(n125) );
  NAND U706 ( .A(n127), .B(n128), .Z(xin[503]) );
  NANDN U707 ( .A(start), .B(xreg[503]), .Z(n128) );
  NAND U708 ( .A(x[503]), .B(start), .Z(n127) );
  NAND U709 ( .A(n129), .B(n130), .Z(xin[502]) );
  NANDN U710 ( .A(start), .B(xreg[502]), .Z(n130) );
  NAND U711 ( .A(x[502]), .B(start), .Z(n129) );
  NAND U712 ( .A(n131), .B(n132), .Z(xin[501]) );
  NANDN U713 ( .A(start), .B(xreg[501]), .Z(n132) );
  NAND U714 ( .A(x[501]), .B(start), .Z(n131) );
  NAND U715 ( .A(n133), .B(n134), .Z(xin[500]) );
  NANDN U716 ( .A(start), .B(xreg[500]), .Z(n134) );
  NAND U717 ( .A(x[500]), .B(start), .Z(n133) );
  NAND U718 ( .A(n135), .B(n136), .Z(xin[4]) );
  NANDN U719 ( .A(start), .B(xreg[4]), .Z(n136) );
  NAND U720 ( .A(x[4]), .B(start), .Z(n135) );
  NAND U721 ( .A(n137), .B(n138), .Z(xin[49]) );
  NANDN U722 ( .A(start), .B(xreg[49]), .Z(n138) );
  NAND U723 ( .A(x[49]), .B(start), .Z(n137) );
  NAND U724 ( .A(n139), .B(n140), .Z(xin[499]) );
  NANDN U725 ( .A(start), .B(xreg[499]), .Z(n140) );
  NAND U726 ( .A(x[499]), .B(start), .Z(n139) );
  NAND U727 ( .A(n141), .B(n142), .Z(xin[498]) );
  NANDN U728 ( .A(start), .B(xreg[498]), .Z(n142) );
  NAND U729 ( .A(x[498]), .B(start), .Z(n141) );
  NAND U730 ( .A(n143), .B(n144), .Z(xin[497]) );
  NANDN U731 ( .A(start), .B(xreg[497]), .Z(n144) );
  NAND U732 ( .A(x[497]), .B(start), .Z(n143) );
  NAND U733 ( .A(n145), .B(n146), .Z(xin[496]) );
  NANDN U734 ( .A(start), .B(xreg[496]), .Z(n146) );
  NAND U735 ( .A(x[496]), .B(start), .Z(n145) );
  NAND U736 ( .A(n147), .B(n148), .Z(xin[495]) );
  NANDN U737 ( .A(start), .B(xreg[495]), .Z(n148) );
  NAND U738 ( .A(x[495]), .B(start), .Z(n147) );
  NAND U739 ( .A(n149), .B(n150), .Z(xin[494]) );
  NANDN U740 ( .A(start), .B(xreg[494]), .Z(n150) );
  NAND U741 ( .A(x[494]), .B(start), .Z(n149) );
  NAND U742 ( .A(n151), .B(n152), .Z(xin[493]) );
  NANDN U743 ( .A(start), .B(xreg[493]), .Z(n152) );
  NAND U744 ( .A(x[493]), .B(start), .Z(n151) );
  NAND U745 ( .A(n153), .B(n154), .Z(xin[492]) );
  NANDN U746 ( .A(start), .B(xreg[492]), .Z(n154) );
  NAND U747 ( .A(x[492]), .B(start), .Z(n153) );
  NAND U748 ( .A(n155), .B(n156), .Z(xin[491]) );
  NANDN U749 ( .A(start), .B(xreg[491]), .Z(n156) );
  NAND U750 ( .A(x[491]), .B(start), .Z(n155) );
  NAND U751 ( .A(n157), .B(n158), .Z(xin[490]) );
  NANDN U752 ( .A(start), .B(xreg[490]), .Z(n158) );
  NAND U753 ( .A(x[490]), .B(start), .Z(n157) );
  NAND U754 ( .A(n159), .B(n160), .Z(xin[48]) );
  NANDN U755 ( .A(start), .B(xreg[48]), .Z(n160) );
  NAND U756 ( .A(x[48]), .B(start), .Z(n159) );
  NAND U757 ( .A(n161), .B(n162), .Z(xin[489]) );
  NANDN U758 ( .A(start), .B(xreg[489]), .Z(n162) );
  NAND U759 ( .A(x[489]), .B(start), .Z(n161) );
  NAND U760 ( .A(n163), .B(n164), .Z(xin[488]) );
  NANDN U761 ( .A(start), .B(xreg[488]), .Z(n164) );
  NAND U762 ( .A(x[488]), .B(start), .Z(n163) );
  NAND U763 ( .A(n165), .B(n166), .Z(xin[487]) );
  NANDN U764 ( .A(start), .B(xreg[487]), .Z(n166) );
  NAND U765 ( .A(x[487]), .B(start), .Z(n165) );
  NAND U766 ( .A(n167), .B(n168), .Z(xin[486]) );
  NANDN U767 ( .A(start), .B(xreg[486]), .Z(n168) );
  NAND U768 ( .A(x[486]), .B(start), .Z(n167) );
  NAND U769 ( .A(n169), .B(n170), .Z(xin[485]) );
  NANDN U770 ( .A(start), .B(xreg[485]), .Z(n170) );
  NAND U771 ( .A(x[485]), .B(start), .Z(n169) );
  NAND U772 ( .A(n171), .B(n172), .Z(xin[484]) );
  NANDN U773 ( .A(start), .B(xreg[484]), .Z(n172) );
  NAND U774 ( .A(x[484]), .B(start), .Z(n171) );
  NAND U775 ( .A(n173), .B(n174), .Z(xin[483]) );
  NANDN U776 ( .A(start), .B(xreg[483]), .Z(n174) );
  NAND U777 ( .A(x[483]), .B(start), .Z(n173) );
  NAND U778 ( .A(n175), .B(n176), .Z(xin[482]) );
  NANDN U779 ( .A(start), .B(xreg[482]), .Z(n176) );
  NAND U780 ( .A(x[482]), .B(start), .Z(n175) );
  NAND U781 ( .A(n177), .B(n178), .Z(xin[481]) );
  NANDN U782 ( .A(start), .B(xreg[481]), .Z(n178) );
  NAND U783 ( .A(x[481]), .B(start), .Z(n177) );
  NAND U784 ( .A(n179), .B(n180), .Z(xin[480]) );
  NANDN U785 ( .A(start), .B(xreg[480]), .Z(n180) );
  NAND U786 ( .A(x[480]), .B(start), .Z(n179) );
  NAND U787 ( .A(n181), .B(n182), .Z(xin[47]) );
  NANDN U788 ( .A(start), .B(xreg[47]), .Z(n182) );
  NAND U789 ( .A(x[47]), .B(start), .Z(n181) );
  NAND U790 ( .A(n183), .B(n184), .Z(xin[479]) );
  NANDN U791 ( .A(start), .B(xreg[479]), .Z(n184) );
  NAND U792 ( .A(x[479]), .B(start), .Z(n183) );
  NAND U793 ( .A(n185), .B(n186), .Z(xin[478]) );
  NANDN U794 ( .A(start), .B(xreg[478]), .Z(n186) );
  NAND U795 ( .A(x[478]), .B(start), .Z(n185) );
  NAND U796 ( .A(n187), .B(n188), .Z(xin[477]) );
  NANDN U797 ( .A(start), .B(xreg[477]), .Z(n188) );
  NAND U798 ( .A(x[477]), .B(start), .Z(n187) );
  NAND U799 ( .A(n189), .B(n190), .Z(xin[476]) );
  NANDN U800 ( .A(start), .B(xreg[476]), .Z(n190) );
  NAND U801 ( .A(x[476]), .B(start), .Z(n189) );
  NAND U802 ( .A(n191), .B(n192), .Z(xin[475]) );
  NANDN U803 ( .A(start), .B(xreg[475]), .Z(n192) );
  NAND U804 ( .A(x[475]), .B(start), .Z(n191) );
  NAND U805 ( .A(n193), .B(n194), .Z(xin[474]) );
  NANDN U806 ( .A(start), .B(xreg[474]), .Z(n194) );
  NAND U807 ( .A(x[474]), .B(start), .Z(n193) );
  NAND U808 ( .A(n195), .B(n196), .Z(xin[473]) );
  NANDN U809 ( .A(start), .B(xreg[473]), .Z(n196) );
  NAND U810 ( .A(x[473]), .B(start), .Z(n195) );
  NAND U811 ( .A(n197), .B(n198), .Z(xin[472]) );
  NANDN U812 ( .A(start), .B(xreg[472]), .Z(n198) );
  NAND U813 ( .A(x[472]), .B(start), .Z(n197) );
  NAND U814 ( .A(n199), .B(n200), .Z(xin[471]) );
  NANDN U815 ( .A(start), .B(xreg[471]), .Z(n200) );
  NAND U816 ( .A(x[471]), .B(start), .Z(n199) );
  NAND U817 ( .A(n201), .B(n202), .Z(xin[470]) );
  NANDN U818 ( .A(start), .B(xreg[470]), .Z(n202) );
  NAND U819 ( .A(x[470]), .B(start), .Z(n201) );
  NAND U820 ( .A(n203), .B(n204), .Z(xin[46]) );
  NANDN U821 ( .A(start), .B(xreg[46]), .Z(n204) );
  NAND U822 ( .A(x[46]), .B(start), .Z(n203) );
  NAND U823 ( .A(n205), .B(n206), .Z(xin[469]) );
  NANDN U824 ( .A(start), .B(xreg[469]), .Z(n206) );
  NAND U825 ( .A(x[469]), .B(start), .Z(n205) );
  NAND U826 ( .A(n207), .B(n208), .Z(xin[468]) );
  NANDN U827 ( .A(start), .B(xreg[468]), .Z(n208) );
  NAND U828 ( .A(x[468]), .B(start), .Z(n207) );
  NAND U829 ( .A(n209), .B(n210), .Z(xin[467]) );
  NANDN U830 ( .A(start), .B(xreg[467]), .Z(n210) );
  NAND U831 ( .A(x[467]), .B(start), .Z(n209) );
  NAND U832 ( .A(n211), .B(n212), .Z(xin[466]) );
  NANDN U833 ( .A(start), .B(xreg[466]), .Z(n212) );
  NAND U834 ( .A(x[466]), .B(start), .Z(n211) );
  NAND U835 ( .A(n213), .B(n214), .Z(xin[465]) );
  NANDN U836 ( .A(start), .B(xreg[465]), .Z(n214) );
  NAND U837 ( .A(x[465]), .B(start), .Z(n213) );
  NAND U838 ( .A(n215), .B(n216), .Z(xin[464]) );
  NANDN U839 ( .A(start), .B(xreg[464]), .Z(n216) );
  NAND U840 ( .A(x[464]), .B(start), .Z(n215) );
  NAND U841 ( .A(n217), .B(n218), .Z(xin[463]) );
  NANDN U842 ( .A(start), .B(xreg[463]), .Z(n218) );
  NAND U843 ( .A(x[463]), .B(start), .Z(n217) );
  NAND U844 ( .A(n219), .B(n220), .Z(xin[462]) );
  NANDN U845 ( .A(start), .B(xreg[462]), .Z(n220) );
  NAND U846 ( .A(x[462]), .B(start), .Z(n219) );
  NAND U847 ( .A(n221), .B(n222), .Z(xin[461]) );
  NANDN U848 ( .A(start), .B(xreg[461]), .Z(n222) );
  NAND U849 ( .A(x[461]), .B(start), .Z(n221) );
  NAND U850 ( .A(n223), .B(n224), .Z(xin[460]) );
  NANDN U851 ( .A(start), .B(xreg[460]), .Z(n224) );
  NAND U852 ( .A(x[460]), .B(start), .Z(n223) );
  NAND U853 ( .A(n225), .B(n226), .Z(xin[45]) );
  NANDN U854 ( .A(start), .B(xreg[45]), .Z(n226) );
  NAND U855 ( .A(x[45]), .B(start), .Z(n225) );
  NAND U856 ( .A(n227), .B(n228), .Z(xin[459]) );
  NANDN U857 ( .A(start), .B(xreg[459]), .Z(n228) );
  NAND U858 ( .A(x[459]), .B(start), .Z(n227) );
  NAND U859 ( .A(n229), .B(n230), .Z(xin[458]) );
  NANDN U860 ( .A(start), .B(xreg[458]), .Z(n230) );
  NAND U861 ( .A(x[458]), .B(start), .Z(n229) );
  NAND U862 ( .A(n231), .B(n232), .Z(xin[457]) );
  NANDN U863 ( .A(start), .B(xreg[457]), .Z(n232) );
  NAND U864 ( .A(x[457]), .B(start), .Z(n231) );
  NAND U865 ( .A(n233), .B(n234), .Z(xin[456]) );
  NANDN U866 ( .A(start), .B(xreg[456]), .Z(n234) );
  NAND U867 ( .A(x[456]), .B(start), .Z(n233) );
  NAND U868 ( .A(n235), .B(n236), .Z(xin[455]) );
  NANDN U869 ( .A(start), .B(xreg[455]), .Z(n236) );
  NAND U870 ( .A(x[455]), .B(start), .Z(n235) );
  NAND U871 ( .A(n237), .B(n238), .Z(xin[454]) );
  NANDN U872 ( .A(start), .B(xreg[454]), .Z(n238) );
  NAND U873 ( .A(x[454]), .B(start), .Z(n237) );
  NAND U874 ( .A(n239), .B(n240), .Z(xin[453]) );
  NANDN U875 ( .A(start), .B(xreg[453]), .Z(n240) );
  NAND U876 ( .A(x[453]), .B(start), .Z(n239) );
  NAND U877 ( .A(n241), .B(n242), .Z(xin[452]) );
  NANDN U878 ( .A(start), .B(xreg[452]), .Z(n242) );
  NAND U879 ( .A(x[452]), .B(start), .Z(n241) );
  NAND U880 ( .A(n243), .B(n244), .Z(xin[451]) );
  NANDN U881 ( .A(start), .B(xreg[451]), .Z(n244) );
  NAND U882 ( .A(x[451]), .B(start), .Z(n243) );
  NAND U883 ( .A(n245), .B(n246), .Z(xin[450]) );
  NANDN U884 ( .A(start), .B(xreg[450]), .Z(n246) );
  NAND U885 ( .A(x[450]), .B(start), .Z(n245) );
  NAND U886 ( .A(n247), .B(n248), .Z(xin[44]) );
  NANDN U887 ( .A(start), .B(xreg[44]), .Z(n248) );
  NAND U888 ( .A(x[44]), .B(start), .Z(n247) );
  NAND U889 ( .A(n249), .B(n250), .Z(xin[449]) );
  NANDN U890 ( .A(start), .B(xreg[449]), .Z(n250) );
  NAND U891 ( .A(x[449]), .B(start), .Z(n249) );
  NAND U892 ( .A(n251), .B(n252), .Z(xin[448]) );
  NANDN U893 ( .A(start), .B(xreg[448]), .Z(n252) );
  NAND U894 ( .A(x[448]), .B(start), .Z(n251) );
  NAND U895 ( .A(n253), .B(n254), .Z(xin[447]) );
  NANDN U896 ( .A(start), .B(xreg[447]), .Z(n254) );
  NAND U897 ( .A(x[447]), .B(start), .Z(n253) );
  NAND U898 ( .A(n255), .B(n256), .Z(xin[446]) );
  NANDN U899 ( .A(start), .B(xreg[446]), .Z(n256) );
  NAND U900 ( .A(x[446]), .B(start), .Z(n255) );
  NAND U901 ( .A(n257), .B(n258), .Z(xin[445]) );
  NANDN U902 ( .A(start), .B(xreg[445]), .Z(n258) );
  NAND U903 ( .A(x[445]), .B(start), .Z(n257) );
  NAND U904 ( .A(n259), .B(n260), .Z(xin[444]) );
  NANDN U905 ( .A(start), .B(xreg[444]), .Z(n260) );
  NAND U906 ( .A(x[444]), .B(start), .Z(n259) );
  NAND U907 ( .A(n261), .B(n262), .Z(xin[443]) );
  NANDN U908 ( .A(start), .B(xreg[443]), .Z(n262) );
  NAND U909 ( .A(x[443]), .B(start), .Z(n261) );
  NAND U910 ( .A(n263), .B(n264), .Z(xin[442]) );
  NANDN U911 ( .A(start), .B(xreg[442]), .Z(n264) );
  NAND U912 ( .A(x[442]), .B(start), .Z(n263) );
  NAND U913 ( .A(n265), .B(n266), .Z(xin[441]) );
  NANDN U914 ( .A(start), .B(xreg[441]), .Z(n266) );
  NAND U915 ( .A(x[441]), .B(start), .Z(n265) );
  NAND U916 ( .A(n267), .B(n268), .Z(xin[440]) );
  NANDN U917 ( .A(start), .B(xreg[440]), .Z(n268) );
  NAND U918 ( .A(x[440]), .B(start), .Z(n267) );
  NAND U919 ( .A(n269), .B(n270), .Z(xin[43]) );
  NANDN U920 ( .A(start), .B(xreg[43]), .Z(n270) );
  NAND U921 ( .A(x[43]), .B(start), .Z(n269) );
  NAND U922 ( .A(n271), .B(n272), .Z(xin[439]) );
  NANDN U923 ( .A(start), .B(xreg[439]), .Z(n272) );
  NAND U924 ( .A(x[439]), .B(start), .Z(n271) );
  NAND U925 ( .A(n273), .B(n274), .Z(xin[438]) );
  NANDN U926 ( .A(start), .B(xreg[438]), .Z(n274) );
  NAND U927 ( .A(x[438]), .B(start), .Z(n273) );
  NAND U928 ( .A(n275), .B(n276), .Z(xin[437]) );
  NANDN U929 ( .A(start), .B(xreg[437]), .Z(n276) );
  NAND U930 ( .A(x[437]), .B(start), .Z(n275) );
  NAND U931 ( .A(n277), .B(n278), .Z(xin[436]) );
  NANDN U932 ( .A(start), .B(xreg[436]), .Z(n278) );
  NAND U933 ( .A(x[436]), .B(start), .Z(n277) );
  NAND U934 ( .A(n279), .B(n280), .Z(xin[435]) );
  NANDN U935 ( .A(start), .B(xreg[435]), .Z(n280) );
  NAND U936 ( .A(x[435]), .B(start), .Z(n279) );
  NAND U937 ( .A(n281), .B(n282), .Z(xin[434]) );
  NANDN U938 ( .A(start), .B(xreg[434]), .Z(n282) );
  NAND U939 ( .A(x[434]), .B(start), .Z(n281) );
  NAND U940 ( .A(n283), .B(n284), .Z(xin[433]) );
  NANDN U941 ( .A(start), .B(xreg[433]), .Z(n284) );
  NAND U942 ( .A(x[433]), .B(start), .Z(n283) );
  NAND U943 ( .A(n285), .B(n286), .Z(xin[432]) );
  NANDN U944 ( .A(start), .B(xreg[432]), .Z(n286) );
  NAND U945 ( .A(x[432]), .B(start), .Z(n285) );
  NAND U946 ( .A(n287), .B(n288), .Z(xin[431]) );
  NANDN U947 ( .A(start), .B(xreg[431]), .Z(n288) );
  NAND U948 ( .A(x[431]), .B(start), .Z(n287) );
  NAND U949 ( .A(n289), .B(n290), .Z(xin[430]) );
  NANDN U950 ( .A(start), .B(xreg[430]), .Z(n290) );
  NAND U951 ( .A(x[430]), .B(start), .Z(n289) );
  NAND U952 ( .A(n291), .B(n292), .Z(xin[42]) );
  NANDN U953 ( .A(start), .B(xreg[42]), .Z(n292) );
  NAND U954 ( .A(x[42]), .B(start), .Z(n291) );
  NAND U955 ( .A(n293), .B(n294), .Z(xin[429]) );
  NANDN U956 ( .A(start), .B(xreg[429]), .Z(n294) );
  NAND U957 ( .A(x[429]), .B(start), .Z(n293) );
  NAND U958 ( .A(n295), .B(n296), .Z(xin[428]) );
  NANDN U959 ( .A(start), .B(xreg[428]), .Z(n296) );
  NAND U960 ( .A(x[428]), .B(start), .Z(n295) );
  NAND U961 ( .A(n297), .B(n298), .Z(xin[427]) );
  NANDN U962 ( .A(start), .B(xreg[427]), .Z(n298) );
  NAND U963 ( .A(x[427]), .B(start), .Z(n297) );
  NAND U964 ( .A(n299), .B(n300), .Z(xin[426]) );
  NANDN U965 ( .A(start), .B(xreg[426]), .Z(n300) );
  NAND U966 ( .A(x[426]), .B(start), .Z(n299) );
  NAND U967 ( .A(n301), .B(n302), .Z(xin[425]) );
  NANDN U968 ( .A(start), .B(xreg[425]), .Z(n302) );
  NAND U969 ( .A(x[425]), .B(start), .Z(n301) );
  NAND U970 ( .A(n303), .B(n304), .Z(xin[424]) );
  NANDN U971 ( .A(start), .B(xreg[424]), .Z(n304) );
  NAND U972 ( .A(x[424]), .B(start), .Z(n303) );
  NAND U973 ( .A(n305), .B(n306), .Z(xin[423]) );
  NANDN U974 ( .A(start), .B(xreg[423]), .Z(n306) );
  NAND U975 ( .A(x[423]), .B(start), .Z(n305) );
  NAND U976 ( .A(n307), .B(n308), .Z(xin[422]) );
  NANDN U977 ( .A(start), .B(xreg[422]), .Z(n308) );
  NAND U978 ( .A(x[422]), .B(start), .Z(n307) );
  NAND U979 ( .A(n309), .B(n310), .Z(xin[421]) );
  NANDN U980 ( .A(start), .B(xreg[421]), .Z(n310) );
  NAND U981 ( .A(x[421]), .B(start), .Z(n309) );
  NAND U982 ( .A(n311), .B(n312), .Z(xin[420]) );
  NANDN U983 ( .A(start), .B(xreg[420]), .Z(n312) );
  NAND U984 ( .A(x[420]), .B(start), .Z(n311) );
  NAND U985 ( .A(n313), .B(n314), .Z(xin[41]) );
  NANDN U986 ( .A(start), .B(xreg[41]), .Z(n314) );
  NAND U987 ( .A(x[41]), .B(start), .Z(n313) );
  NAND U988 ( .A(n315), .B(n316), .Z(xin[419]) );
  NANDN U989 ( .A(start), .B(xreg[419]), .Z(n316) );
  NAND U990 ( .A(x[419]), .B(start), .Z(n315) );
  NAND U991 ( .A(n317), .B(n318), .Z(xin[418]) );
  NANDN U992 ( .A(start), .B(xreg[418]), .Z(n318) );
  NAND U993 ( .A(x[418]), .B(start), .Z(n317) );
  NAND U994 ( .A(n319), .B(n320), .Z(xin[417]) );
  NANDN U995 ( .A(start), .B(xreg[417]), .Z(n320) );
  NAND U996 ( .A(x[417]), .B(start), .Z(n319) );
  NAND U997 ( .A(n321), .B(n322), .Z(xin[416]) );
  NANDN U998 ( .A(start), .B(xreg[416]), .Z(n322) );
  NAND U999 ( .A(x[416]), .B(start), .Z(n321) );
  NAND U1000 ( .A(n323), .B(n324), .Z(xin[415]) );
  NANDN U1001 ( .A(start), .B(xreg[415]), .Z(n324) );
  NAND U1002 ( .A(x[415]), .B(start), .Z(n323) );
  NAND U1003 ( .A(n325), .B(n326), .Z(xin[414]) );
  NANDN U1004 ( .A(start), .B(xreg[414]), .Z(n326) );
  NAND U1005 ( .A(x[414]), .B(start), .Z(n325) );
  NAND U1006 ( .A(n327), .B(n328), .Z(xin[413]) );
  NANDN U1007 ( .A(start), .B(xreg[413]), .Z(n328) );
  NAND U1008 ( .A(x[413]), .B(start), .Z(n327) );
  NAND U1009 ( .A(n329), .B(n330), .Z(xin[412]) );
  NANDN U1010 ( .A(start), .B(xreg[412]), .Z(n330) );
  NAND U1011 ( .A(x[412]), .B(start), .Z(n329) );
  NAND U1012 ( .A(n331), .B(n332), .Z(xin[411]) );
  NANDN U1013 ( .A(start), .B(xreg[411]), .Z(n332) );
  NAND U1014 ( .A(x[411]), .B(start), .Z(n331) );
  NAND U1015 ( .A(n333), .B(n334), .Z(xin[410]) );
  NANDN U1016 ( .A(start), .B(xreg[410]), .Z(n334) );
  NAND U1017 ( .A(x[410]), .B(start), .Z(n333) );
  NAND U1018 ( .A(n335), .B(n336), .Z(xin[40]) );
  NANDN U1019 ( .A(start), .B(xreg[40]), .Z(n336) );
  NAND U1020 ( .A(x[40]), .B(start), .Z(n335) );
  NAND U1021 ( .A(n337), .B(n338), .Z(xin[409]) );
  NANDN U1022 ( .A(start), .B(xreg[409]), .Z(n338) );
  NAND U1023 ( .A(x[409]), .B(start), .Z(n337) );
  NAND U1024 ( .A(n339), .B(n340), .Z(xin[408]) );
  NANDN U1025 ( .A(start), .B(xreg[408]), .Z(n340) );
  NAND U1026 ( .A(x[408]), .B(start), .Z(n339) );
  NAND U1027 ( .A(n341), .B(n342), .Z(xin[407]) );
  NANDN U1028 ( .A(start), .B(xreg[407]), .Z(n342) );
  NAND U1029 ( .A(x[407]), .B(start), .Z(n341) );
  NAND U1030 ( .A(n343), .B(n344), .Z(xin[406]) );
  NANDN U1031 ( .A(start), .B(xreg[406]), .Z(n344) );
  NAND U1032 ( .A(x[406]), .B(start), .Z(n343) );
  NAND U1033 ( .A(n345), .B(n346), .Z(xin[405]) );
  NANDN U1034 ( .A(start), .B(xreg[405]), .Z(n346) );
  NAND U1035 ( .A(x[405]), .B(start), .Z(n345) );
  NAND U1036 ( .A(n347), .B(n348), .Z(xin[404]) );
  NANDN U1037 ( .A(start), .B(xreg[404]), .Z(n348) );
  NAND U1038 ( .A(x[404]), .B(start), .Z(n347) );
  NAND U1039 ( .A(n349), .B(n350), .Z(xin[403]) );
  NANDN U1040 ( .A(start), .B(xreg[403]), .Z(n350) );
  NAND U1041 ( .A(x[403]), .B(start), .Z(n349) );
  NAND U1042 ( .A(n351), .B(n352), .Z(xin[402]) );
  NANDN U1043 ( .A(start), .B(xreg[402]), .Z(n352) );
  NAND U1044 ( .A(x[402]), .B(start), .Z(n351) );
  NAND U1045 ( .A(n353), .B(n354), .Z(xin[401]) );
  NANDN U1046 ( .A(start), .B(xreg[401]), .Z(n354) );
  NAND U1047 ( .A(x[401]), .B(start), .Z(n353) );
  NAND U1048 ( .A(n355), .B(n356), .Z(xin[400]) );
  NANDN U1049 ( .A(start), .B(xreg[400]), .Z(n356) );
  NAND U1050 ( .A(x[400]), .B(start), .Z(n355) );
  NAND U1051 ( .A(n357), .B(n358), .Z(xin[3]) );
  NANDN U1052 ( .A(start), .B(xreg[3]), .Z(n358) );
  NAND U1053 ( .A(x[3]), .B(start), .Z(n357) );
  NAND U1054 ( .A(n359), .B(n360), .Z(xin[39]) );
  NANDN U1055 ( .A(start), .B(xreg[39]), .Z(n360) );
  NAND U1056 ( .A(x[39]), .B(start), .Z(n359) );
  NAND U1057 ( .A(n361), .B(n362), .Z(xin[399]) );
  NANDN U1058 ( .A(start), .B(xreg[399]), .Z(n362) );
  NAND U1059 ( .A(x[399]), .B(start), .Z(n361) );
  NAND U1060 ( .A(n363), .B(n364), .Z(xin[398]) );
  NANDN U1061 ( .A(start), .B(xreg[398]), .Z(n364) );
  NAND U1062 ( .A(x[398]), .B(start), .Z(n363) );
  NAND U1063 ( .A(n365), .B(n366), .Z(xin[397]) );
  NANDN U1064 ( .A(start), .B(xreg[397]), .Z(n366) );
  NAND U1065 ( .A(x[397]), .B(start), .Z(n365) );
  NAND U1066 ( .A(n367), .B(n368), .Z(xin[396]) );
  NANDN U1067 ( .A(start), .B(xreg[396]), .Z(n368) );
  NAND U1068 ( .A(x[396]), .B(start), .Z(n367) );
  NAND U1069 ( .A(n369), .B(n370), .Z(xin[395]) );
  NANDN U1070 ( .A(start), .B(xreg[395]), .Z(n370) );
  NAND U1071 ( .A(x[395]), .B(start), .Z(n369) );
  NAND U1072 ( .A(n371), .B(n372), .Z(xin[394]) );
  NANDN U1073 ( .A(start), .B(xreg[394]), .Z(n372) );
  NAND U1074 ( .A(x[394]), .B(start), .Z(n371) );
  NAND U1075 ( .A(n373), .B(n374), .Z(xin[393]) );
  NANDN U1076 ( .A(start), .B(xreg[393]), .Z(n374) );
  NAND U1077 ( .A(x[393]), .B(start), .Z(n373) );
  NAND U1078 ( .A(n375), .B(n376), .Z(xin[392]) );
  NANDN U1079 ( .A(start), .B(xreg[392]), .Z(n376) );
  NAND U1080 ( .A(x[392]), .B(start), .Z(n375) );
  NAND U1081 ( .A(n377), .B(n378), .Z(xin[391]) );
  NANDN U1082 ( .A(start), .B(xreg[391]), .Z(n378) );
  NAND U1083 ( .A(x[391]), .B(start), .Z(n377) );
  NAND U1084 ( .A(n379), .B(n380), .Z(xin[390]) );
  NANDN U1085 ( .A(start), .B(xreg[390]), .Z(n380) );
  NAND U1086 ( .A(x[390]), .B(start), .Z(n379) );
  NAND U1087 ( .A(n381), .B(n382), .Z(xin[38]) );
  NANDN U1088 ( .A(start), .B(xreg[38]), .Z(n382) );
  NAND U1089 ( .A(x[38]), .B(start), .Z(n381) );
  NAND U1090 ( .A(n383), .B(n384), .Z(xin[389]) );
  NANDN U1091 ( .A(start), .B(xreg[389]), .Z(n384) );
  NAND U1092 ( .A(x[389]), .B(start), .Z(n383) );
  NAND U1093 ( .A(n385), .B(n386), .Z(xin[388]) );
  NANDN U1094 ( .A(start), .B(xreg[388]), .Z(n386) );
  NAND U1095 ( .A(x[388]), .B(start), .Z(n385) );
  NAND U1096 ( .A(n387), .B(n388), .Z(xin[387]) );
  NANDN U1097 ( .A(start), .B(xreg[387]), .Z(n388) );
  NAND U1098 ( .A(x[387]), .B(start), .Z(n387) );
  NAND U1099 ( .A(n389), .B(n390), .Z(xin[386]) );
  NANDN U1100 ( .A(start), .B(xreg[386]), .Z(n390) );
  NAND U1101 ( .A(x[386]), .B(start), .Z(n389) );
  NAND U1102 ( .A(n391), .B(n392), .Z(xin[385]) );
  NANDN U1103 ( .A(start), .B(xreg[385]), .Z(n392) );
  NAND U1104 ( .A(x[385]), .B(start), .Z(n391) );
  NAND U1105 ( .A(n393), .B(n394), .Z(xin[384]) );
  NANDN U1106 ( .A(start), .B(xreg[384]), .Z(n394) );
  NAND U1107 ( .A(x[384]), .B(start), .Z(n393) );
  NAND U1108 ( .A(n395), .B(n396), .Z(xin[383]) );
  NANDN U1109 ( .A(start), .B(xreg[383]), .Z(n396) );
  NAND U1110 ( .A(x[383]), .B(start), .Z(n395) );
  NAND U1111 ( .A(n397), .B(n398), .Z(xin[382]) );
  NANDN U1112 ( .A(start), .B(xreg[382]), .Z(n398) );
  NAND U1113 ( .A(x[382]), .B(start), .Z(n397) );
  NAND U1114 ( .A(n399), .B(n400), .Z(xin[381]) );
  NANDN U1115 ( .A(start), .B(xreg[381]), .Z(n400) );
  NAND U1116 ( .A(x[381]), .B(start), .Z(n399) );
  NAND U1117 ( .A(n401), .B(n402), .Z(xin[380]) );
  NANDN U1118 ( .A(start), .B(xreg[380]), .Z(n402) );
  NAND U1119 ( .A(x[380]), .B(start), .Z(n401) );
  NAND U1120 ( .A(n403), .B(n404), .Z(xin[37]) );
  NANDN U1121 ( .A(start), .B(xreg[37]), .Z(n404) );
  NAND U1122 ( .A(x[37]), .B(start), .Z(n403) );
  NAND U1123 ( .A(n405), .B(n406), .Z(xin[379]) );
  NANDN U1124 ( .A(start), .B(xreg[379]), .Z(n406) );
  NAND U1125 ( .A(x[379]), .B(start), .Z(n405) );
  NAND U1126 ( .A(n407), .B(n408), .Z(xin[378]) );
  NANDN U1127 ( .A(start), .B(xreg[378]), .Z(n408) );
  NAND U1128 ( .A(x[378]), .B(start), .Z(n407) );
  NAND U1129 ( .A(n409), .B(n410), .Z(xin[377]) );
  NANDN U1130 ( .A(start), .B(xreg[377]), .Z(n410) );
  NAND U1131 ( .A(x[377]), .B(start), .Z(n409) );
  NAND U1132 ( .A(n411), .B(n412), .Z(xin[376]) );
  NANDN U1133 ( .A(start), .B(xreg[376]), .Z(n412) );
  NAND U1134 ( .A(x[376]), .B(start), .Z(n411) );
  NAND U1135 ( .A(n413), .B(n414), .Z(xin[375]) );
  NANDN U1136 ( .A(start), .B(xreg[375]), .Z(n414) );
  NAND U1137 ( .A(x[375]), .B(start), .Z(n413) );
  NAND U1138 ( .A(n415), .B(n416), .Z(xin[374]) );
  NANDN U1139 ( .A(start), .B(xreg[374]), .Z(n416) );
  NAND U1140 ( .A(x[374]), .B(start), .Z(n415) );
  NAND U1141 ( .A(n417), .B(n418), .Z(xin[373]) );
  NANDN U1142 ( .A(start), .B(xreg[373]), .Z(n418) );
  NAND U1143 ( .A(x[373]), .B(start), .Z(n417) );
  NAND U1144 ( .A(n419), .B(n420), .Z(xin[372]) );
  NANDN U1145 ( .A(start), .B(xreg[372]), .Z(n420) );
  NAND U1146 ( .A(x[372]), .B(start), .Z(n419) );
  NAND U1147 ( .A(n421), .B(n422), .Z(xin[371]) );
  NANDN U1148 ( .A(start), .B(xreg[371]), .Z(n422) );
  NAND U1149 ( .A(x[371]), .B(start), .Z(n421) );
  NAND U1150 ( .A(n423), .B(n424), .Z(xin[370]) );
  NANDN U1151 ( .A(start), .B(xreg[370]), .Z(n424) );
  NAND U1152 ( .A(x[370]), .B(start), .Z(n423) );
  NAND U1153 ( .A(n425), .B(n426), .Z(xin[36]) );
  NANDN U1154 ( .A(start), .B(xreg[36]), .Z(n426) );
  NAND U1155 ( .A(x[36]), .B(start), .Z(n425) );
  NAND U1156 ( .A(n427), .B(n428), .Z(xin[369]) );
  NANDN U1157 ( .A(start), .B(xreg[369]), .Z(n428) );
  NAND U1158 ( .A(x[369]), .B(start), .Z(n427) );
  NAND U1159 ( .A(n429), .B(n430), .Z(xin[368]) );
  NANDN U1160 ( .A(start), .B(xreg[368]), .Z(n430) );
  NAND U1161 ( .A(x[368]), .B(start), .Z(n429) );
  NAND U1162 ( .A(n431), .B(n432), .Z(xin[367]) );
  NANDN U1163 ( .A(start), .B(xreg[367]), .Z(n432) );
  NAND U1164 ( .A(x[367]), .B(start), .Z(n431) );
  NAND U1165 ( .A(n433), .B(n434), .Z(xin[366]) );
  NANDN U1166 ( .A(start), .B(xreg[366]), .Z(n434) );
  NAND U1167 ( .A(x[366]), .B(start), .Z(n433) );
  NAND U1168 ( .A(n435), .B(n436), .Z(xin[365]) );
  NANDN U1169 ( .A(start), .B(xreg[365]), .Z(n436) );
  NAND U1170 ( .A(x[365]), .B(start), .Z(n435) );
  NAND U1171 ( .A(n437), .B(n438), .Z(xin[364]) );
  NANDN U1172 ( .A(start), .B(xreg[364]), .Z(n438) );
  NAND U1173 ( .A(x[364]), .B(start), .Z(n437) );
  NAND U1174 ( .A(n439), .B(n440), .Z(xin[363]) );
  NANDN U1175 ( .A(start), .B(xreg[363]), .Z(n440) );
  NAND U1176 ( .A(x[363]), .B(start), .Z(n439) );
  NAND U1177 ( .A(n441), .B(n442), .Z(xin[362]) );
  NANDN U1178 ( .A(start), .B(xreg[362]), .Z(n442) );
  NAND U1179 ( .A(x[362]), .B(start), .Z(n441) );
  NAND U1180 ( .A(n443), .B(n444), .Z(xin[361]) );
  NANDN U1181 ( .A(start), .B(xreg[361]), .Z(n444) );
  NAND U1182 ( .A(x[361]), .B(start), .Z(n443) );
  NAND U1183 ( .A(n445), .B(n446), .Z(xin[360]) );
  NANDN U1184 ( .A(start), .B(xreg[360]), .Z(n446) );
  NAND U1185 ( .A(x[360]), .B(start), .Z(n445) );
  NAND U1186 ( .A(n447), .B(n448), .Z(xin[35]) );
  NANDN U1187 ( .A(start), .B(xreg[35]), .Z(n448) );
  NAND U1188 ( .A(x[35]), .B(start), .Z(n447) );
  NAND U1189 ( .A(n449), .B(n450), .Z(xin[359]) );
  NANDN U1190 ( .A(start), .B(xreg[359]), .Z(n450) );
  NAND U1191 ( .A(x[359]), .B(start), .Z(n449) );
  NAND U1192 ( .A(n451), .B(n452), .Z(xin[358]) );
  NANDN U1193 ( .A(start), .B(xreg[358]), .Z(n452) );
  NAND U1194 ( .A(x[358]), .B(start), .Z(n451) );
  NAND U1195 ( .A(n453), .B(n454), .Z(xin[357]) );
  NANDN U1196 ( .A(start), .B(xreg[357]), .Z(n454) );
  NAND U1197 ( .A(x[357]), .B(start), .Z(n453) );
  NAND U1198 ( .A(n455), .B(n456), .Z(xin[356]) );
  NANDN U1199 ( .A(start), .B(xreg[356]), .Z(n456) );
  NAND U1200 ( .A(x[356]), .B(start), .Z(n455) );
  NAND U1201 ( .A(n457), .B(n458), .Z(xin[355]) );
  NANDN U1202 ( .A(start), .B(xreg[355]), .Z(n458) );
  NAND U1203 ( .A(x[355]), .B(start), .Z(n457) );
  NAND U1204 ( .A(n459), .B(n460), .Z(xin[354]) );
  NANDN U1205 ( .A(start), .B(xreg[354]), .Z(n460) );
  NAND U1206 ( .A(x[354]), .B(start), .Z(n459) );
  NAND U1207 ( .A(n461), .B(n462), .Z(xin[353]) );
  NANDN U1208 ( .A(start), .B(xreg[353]), .Z(n462) );
  NAND U1209 ( .A(x[353]), .B(start), .Z(n461) );
  NAND U1210 ( .A(n463), .B(n464), .Z(xin[352]) );
  NANDN U1211 ( .A(start), .B(xreg[352]), .Z(n464) );
  NAND U1212 ( .A(x[352]), .B(start), .Z(n463) );
  NAND U1213 ( .A(n465), .B(n466), .Z(xin[351]) );
  NANDN U1214 ( .A(start), .B(xreg[351]), .Z(n466) );
  NAND U1215 ( .A(x[351]), .B(start), .Z(n465) );
  NAND U1216 ( .A(n467), .B(n468), .Z(xin[350]) );
  NANDN U1217 ( .A(start), .B(xreg[350]), .Z(n468) );
  NAND U1218 ( .A(x[350]), .B(start), .Z(n467) );
  NAND U1219 ( .A(n469), .B(n470), .Z(xin[34]) );
  NANDN U1220 ( .A(start), .B(xreg[34]), .Z(n470) );
  NAND U1221 ( .A(x[34]), .B(start), .Z(n469) );
  NAND U1222 ( .A(n471), .B(n472), .Z(xin[349]) );
  NANDN U1223 ( .A(start), .B(xreg[349]), .Z(n472) );
  NAND U1224 ( .A(x[349]), .B(start), .Z(n471) );
  NAND U1225 ( .A(n473), .B(n474), .Z(xin[348]) );
  NANDN U1226 ( .A(start), .B(xreg[348]), .Z(n474) );
  NAND U1227 ( .A(x[348]), .B(start), .Z(n473) );
  NAND U1228 ( .A(n475), .B(n476), .Z(xin[347]) );
  NANDN U1229 ( .A(start), .B(xreg[347]), .Z(n476) );
  NAND U1230 ( .A(x[347]), .B(start), .Z(n475) );
  NAND U1231 ( .A(n477), .B(n478), .Z(xin[346]) );
  NANDN U1232 ( .A(start), .B(xreg[346]), .Z(n478) );
  NAND U1233 ( .A(x[346]), .B(start), .Z(n477) );
  NAND U1234 ( .A(n479), .B(n480), .Z(xin[345]) );
  NANDN U1235 ( .A(start), .B(xreg[345]), .Z(n480) );
  NAND U1236 ( .A(x[345]), .B(start), .Z(n479) );
  NAND U1237 ( .A(n481), .B(n482), .Z(xin[344]) );
  NANDN U1238 ( .A(start), .B(xreg[344]), .Z(n482) );
  NAND U1239 ( .A(x[344]), .B(start), .Z(n481) );
  NAND U1240 ( .A(n483), .B(n484), .Z(xin[343]) );
  NANDN U1241 ( .A(start), .B(xreg[343]), .Z(n484) );
  NAND U1242 ( .A(x[343]), .B(start), .Z(n483) );
  NAND U1243 ( .A(n485), .B(n486), .Z(xin[342]) );
  NANDN U1244 ( .A(start), .B(xreg[342]), .Z(n486) );
  NAND U1245 ( .A(x[342]), .B(start), .Z(n485) );
  NAND U1246 ( .A(n487), .B(n488), .Z(xin[341]) );
  NANDN U1247 ( .A(start), .B(xreg[341]), .Z(n488) );
  NAND U1248 ( .A(x[341]), .B(start), .Z(n487) );
  NAND U1249 ( .A(n489), .B(n490), .Z(xin[340]) );
  NANDN U1250 ( .A(start), .B(xreg[340]), .Z(n490) );
  NAND U1251 ( .A(x[340]), .B(start), .Z(n489) );
  NAND U1252 ( .A(n491), .B(n492), .Z(xin[33]) );
  NANDN U1253 ( .A(start), .B(xreg[33]), .Z(n492) );
  NAND U1254 ( .A(x[33]), .B(start), .Z(n491) );
  NAND U1255 ( .A(n493), .B(n494), .Z(xin[339]) );
  NANDN U1256 ( .A(start), .B(xreg[339]), .Z(n494) );
  NAND U1257 ( .A(x[339]), .B(start), .Z(n493) );
  NAND U1258 ( .A(n495), .B(n496), .Z(xin[338]) );
  NANDN U1259 ( .A(start), .B(xreg[338]), .Z(n496) );
  NAND U1260 ( .A(x[338]), .B(start), .Z(n495) );
  NAND U1261 ( .A(n497), .B(n498), .Z(xin[337]) );
  NANDN U1262 ( .A(start), .B(xreg[337]), .Z(n498) );
  NAND U1263 ( .A(x[337]), .B(start), .Z(n497) );
  NAND U1264 ( .A(n499), .B(n500), .Z(xin[336]) );
  NANDN U1265 ( .A(start), .B(xreg[336]), .Z(n500) );
  NAND U1266 ( .A(x[336]), .B(start), .Z(n499) );
  NAND U1267 ( .A(n501), .B(n502), .Z(xin[335]) );
  NANDN U1268 ( .A(start), .B(xreg[335]), .Z(n502) );
  NAND U1269 ( .A(x[335]), .B(start), .Z(n501) );
  NAND U1270 ( .A(n503), .B(n504), .Z(xin[334]) );
  NANDN U1271 ( .A(start), .B(xreg[334]), .Z(n504) );
  NAND U1272 ( .A(x[334]), .B(start), .Z(n503) );
  NAND U1273 ( .A(n505), .B(n506), .Z(xin[333]) );
  NANDN U1274 ( .A(start), .B(xreg[333]), .Z(n506) );
  NAND U1275 ( .A(x[333]), .B(start), .Z(n505) );
  NAND U1276 ( .A(n507), .B(n508), .Z(xin[332]) );
  NANDN U1277 ( .A(start), .B(xreg[332]), .Z(n508) );
  NAND U1278 ( .A(x[332]), .B(start), .Z(n507) );
  NAND U1279 ( .A(n509), .B(n510), .Z(xin[331]) );
  NANDN U1280 ( .A(start), .B(xreg[331]), .Z(n510) );
  NAND U1281 ( .A(x[331]), .B(start), .Z(n509) );
  NAND U1282 ( .A(n511), .B(n512), .Z(xin[330]) );
  NANDN U1283 ( .A(start), .B(xreg[330]), .Z(n512) );
  NAND U1284 ( .A(x[330]), .B(start), .Z(n511) );
  NAND U1285 ( .A(n513), .B(n514), .Z(xin[32]) );
  NANDN U1286 ( .A(start), .B(xreg[32]), .Z(n514) );
  NAND U1287 ( .A(x[32]), .B(start), .Z(n513) );
  NAND U1288 ( .A(n515), .B(n516), .Z(xin[329]) );
  NANDN U1289 ( .A(start), .B(xreg[329]), .Z(n516) );
  NAND U1290 ( .A(x[329]), .B(start), .Z(n515) );
  NAND U1291 ( .A(n517), .B(n518), .Z(xin[328]) );
  NANDN U1292 ( .A(start), .B(xreg[328]), .Z(n518) );
  NAND U1293 ( .A(x[328]), .B(start), .Z(n517) );
  NAND U1294 ( .A(n519), .B(n520), .Z(xin[327]) );
  NANDN U1295 ( .A(start), .B(xreg[327]), .Z(n520) );
  NAND U1296 ( .A(x[327]), .B(start), .Z(n519) );
  NAND U1297 ( .A(n521), .B(n522), .Z(xin[326]) );
  NANDN U1298 ( .A(start), .B(xreg[326]), .Z(n522) );
  NAND U1299 ( .A(x[326]), .B(start), .Z(n521) );
  NAND U1300 ( .A(n523), .B(n524), .Z(xin[325]) );
  NANDN U1301 ( .A(start), .B(xreg[325]), .Z(n524) );
  NAND U1302 ( .A(x[325]), .B(start), .Z(n523) );
  NAND U1303 ( .A(n525), .B(n526), .Z(xin[324]) );
  NANDN U1304 ( .A(start), .B(xreg[324]), .Z(n526) );
  NAND U1305 ( .A(x[324]), .B(start), .Z(n525) );
  NAND U1306 ( .A(n527), .B(n528), .Z(xin[323]) );
  NANDN U1307 ( .A(start), .B(xreg[323]), .Z(n528) );
  NAND U1308 ( .A(x[323]), .B(start), .Z(n527) );
  NAND U1309 ( .A(n529), .B(n530), .Z(xin[322]) );
  NANDN U1310 ( .A(start), .B(xreg[322]), .Z(n530) );
  NAND U1311 ( .A(x[322]), .B(start), .Z(n529) );
  NAND U1312 ( .A(n531), .B(n532), .Z(xin[321]) );
  NANDN U1313 ( .A(start), .B(xreg[321]), .Z(n532) );
  NAND U1314 ( .A(x[321]), .B(start), .Z(n531) );
  NAND U1315 ( .A(n533), .B(n534), .Z(xin[320]) );
  NANDN U1316 ( .A(start), .B(xreg[320]), .Z(n534) );
  NAND U1317 ( .A(x[320]), .B(start), .Z(n533) );
  NAND U1318 ( .A(n535), .B(n536), .Z(xin[31]) );
  NANDN U1319 ( .A(start), .B(xreg[31]), .Z(n536) );
  NAND U1320 ( .A(x[31]), .B(start), .Z(n535) );
  NAND U1321 ( .A(n537), .B(n538), .Z(xin[319]) );
  NANDN U1322 ( .A(start), .B(xreg[319]), .Z(n538) );
  NAND U1323 ( .A(x[319]), .B(start), .Z(n537) );
  NAND U1324 ( .A(n539), .B(n540), .Z(xin[318]) );
  NANDN U1325 ( .A(start), .B(xreg[318]), .Z(n540) );
  NAND U1326 ( .A(x[318]), .B(start), .Z(n539) );
  NAND U1327 ( .A(n541), .B(n542), .Z(xin[317]) );
  NANDN U1328 ( .A(start), .B(xreg[317]), .Z(n542) );
  NAND U1329 ( .A(x[317]), .B(start), .Z(n541) );
  NAND U1330 ( .A(n543), .B(n544), .Z(xin[316]) );
  NANDN U1331 ( .A(start), .B(xreg[316]), .Z(n544) );
  NAND U1332 ( .A(x[316]), .B(start), .Z(n543) );
  NAND U1333 ( .A(n545), .B(n546), .Z(xin[315]) );
  NANDN U1334 ( .A(start), .B(xreg[315]), .Z(n546) );
  NAND U1335 ( .A(x[315]), .B(start), .Z(n545) );
  NAND U1336 ( .A(n547), .B(n548), .Z(xin[314]) );
  NANDN U1337 ( .A(start), .B(xreg[314]), .Z(n548) );
  NAND U1338 ( .A(x[314]), .B(start), .Z(n547) );
  NAND U1339 ( .A(n549), .B(n550), .Z(xin[313]) );
  NANDN U1340 ( .A(start), .B(xreg[313]), .Z(n550) );
  NAND U1341 ( .A(x[313]), .B(start), .Z(n549) );
  NAND U1342 ( .A(n551), .B(n552), .Z(xin[312]) );
  NANDN U1343 ( .A(start), .B(xreg[312]), .Z(n552) );
  NAND U1344 ( .A(x[312]), .B(start), .Z(n551) );
  NAND U1345 ( .A(n553), .B(n554), .Z(xin[311]) );
  NANDN U1346 ( .A(start), .B(xreg[311]), .Z(n554) );
  NAND U1347 ( .A(x[311]), .B(start), .Z(n553) );
  NAND U1348 ( .A(n555), .B(n556), .Z(xin[310]) );
  NANDN U1349 ( .A(start), .B(xreg[310]), .Z(n556) );
  NAND U1350 ( .A(x[310]), .B(start), .Z(n555) );
  NAND U1351 ( .A(n557), .B(n558), .Z(xin[30]) );
  NANDN U1352 ( .A(start), .B(xreg[30]), .Z(n558) );
  NAND U1353 ( .A(x[30]), .B(start), .Z(n557) );
  NAND U1354 ( .A(n559), .B(n560), .Z(xin[309]) );
  NANDN U1355 ( .A(start), .B(xreg[309]), .Z(n560) );
  NAND U1356 ( .A(x[309]), .B(start), .Z(n559) );
  NAND U1357 ( .A(n561), .B(n562), .Z(xin[308]) );
  NANDN U1358 ( .A(start), .B(xreg[308]), .Z(n562) );
  NAND U1359 ( .A(x[308]), .B(start), .Z(n561) );
  NAND U1360 ( .A(n563), .B(n564), .Z(xin[307]) );
  NANDN U1361 ( .A(start), .B(xreg[307]), .Z(n564) );
  NAND U1362 ( .A(x[307]), .B(start), .Z(n563) );
  NAND U1363 ( .A(n565), .B(n566), .Z(xin[306]) );
  NANDN U1364 ( .A(start), .B(xreg[306]), .Z(n566) );
  NAND U1365 ( .A(x[306]), .B(start), .Z(n565) );
  NAND U1366 ( .A(n567), .B(n568), .Z(xin[305]) );
  NANDN U1367 ( .A(start), .B(xreg[305]), .Z(n568) );
  NAND U1368 ( .A(x[305]), .B(start), .Z(n567) );
  NAND U1369 ( .A(n569), .B(n570), .Z(xin[304]) );
  NANDN U1370 ( .A(start), .B(xreg[304]), .Z(n570) );
  NAND U1371 ( .A(x[304]), .B(start), .Z(n569) );
  NAND U1372 ( .A(n571), .B(n572), .Z(xin[303]) );
  NANDN U1373 ( .A(start), .B(xreg[303]), .Z(n572) );
  NAND U1374 ( .A(x[303]), .B(start), .Z(n571) );
  NAND U1375 ( .A(n573), .B(n574), .Z(xin[302]) );
  NANDN U1376 ( .A(start), .B(xreg[302]), .Z(n574) );
  NAND U1377 ( .A(x[302]), .B(start), .Z(n573) );
  NAND U1378 ( .A(n575), .B(n576), .Z(xin[301]) );
  NANDN U1379 ( .A(start), .B(xreg[301]), .Z(n576) );
  NAND U1380 ( .A(x[301]), .B(start), .Z(n575) );
  NAND U1381 ( .A(n577), .B(n578), .Z(xin[300]) );
  NANDN U1382 ( .A(start), .B(xreg[300]), .Z(n578) );
  NAND U1383 ( .A(x[300]), .B(start), .Z(n577) );
  NAND U1384 ( .A(n579), .B(n580), .Z(xin[2]) );
  NANDN U1385 ( .A(start), .B(xreg[2]), .Z(n580) );
  NAND U1386 ( .A(x[2]), .B(start), .Z(n579) );
  NAND U1387 ( .A(n581), .B(n582), .Z(xin[29]) );
  NANDN U1388 ( .A(start), .B(xreg[29]), .Z(n582) );
  NAND U1389 ( .A(x[29]), .B(start), .Z(n581) );
  NAND U1390 ( .A(n583), .B(n584), .Z(xin[299]) );
  NANDN U1391 ( .A(start), .B(xreg[299]), .Z(n584) );
  NAND U1392 ( .A(x[299]), .B(start), .Z(n583) );
  NAND U1393 ( .A(n585), .B(n586), .Z(xin[298]) );
  NANDN U1394 ( .A(start), .B(xreg[298]), .Z(n586) );
  NAND U1395 ( .A(x[298]), .B(start), .Z(n585) );
  NAND U1396 ( .A(n587), .B(n588), .Z(xin[297]) );
  NANDN U1397 ( .A(start), .B(xreg[297]), .Z(n588) );
  NAND U1398 ( .A(x[297]), .B(start), .Z(n587) );
  NAND U1399 ( .A(n589), .B(n590), .Z(xin[296]) );
  NANDN U1400 ( .A(start), .B(xreg[296]), .Z(n590) );
  NAND U1401 ( .A(x[296]), .B(start), .Z(n589) );
  NAND U1402 ( .A(n591), .B(n592), .Z(xin[295]) );
  NANDN U1403 ( .A(start), .B(xreg[295]), .Z(n592) );
  NAND U1404 ( .A(x[295]), .B(start), .Z(n591) );
  NAND U1405 ( .A(n593), .B(n594), .Z(xin[294]) );
  NANDN U1406 ( .A(start), .B(xreg[294]), .Z(n594) );
  NAND U1407 ( .A(x[294]), .B(start), .Z(n593) );
  NAND U1408 ( .A(n595), .B(n596), .Z(xin[293]) );
  NANDN U1409 ( .A(start), .B(xreg[293]), .Z(n596) );
  NAND U1410 ( .A(x[293]), .B(start), .Z(n595) );
  NAND U1411 ( .A(n597), .B(n598), .Z(xin[292]) );
  NANDN U1412 ( .A(start), .B(xreg[292]), .Z(n598) );
  NAND U1413 ( .A(x[292]), .B(start), .Z(n597) );
  NAND U1414 ( .A(n599), .B(n600), .Z(xin[291]) );
  NANDN U1415 ( .A(start), .B(xreg[291]), .Z(n600) );
  NAND U1416 ( .A(x[291]), .B(start), .Z(n599) );
  NAND U1417 ( .A(n601), .B(n602), .Z(xin[290]) );
  NANDN U1418 ( .A(start), .B(xreg[290]), .Z(n602) );
  NAND U1419 ( .A(x[290]), .B(start), .Z(n601) );
  NAND U1420 ( .A(n603), .B(n604), .Z(xin[28]) );
  NANDN U1421 ( .A(start), .B(xreg[28]), .Z(n604) );
  NAND U1422 ( .A(x[28]), .B(start), .Z(n603) );
  NAND U1423 ( .A(n605), .B(n606), .Z(xin[289]) );
  NANDN U1424 ( .A(start), .B(xreg[289]), .Z(n606) );
  NAND U1425 ( .A(x[289]), .B(start), .Z(n605) );
  NAND U1426 ( .A(n607), .B(n608), .Z(xin[288]) );
  NANDN U1427 ( .A(start), .B(xreg[288]), .Z(n608) );
  NAND U1428 ( .A(x[288]), .B(start), .Z(n607) );
  NAND U1429 ( .A(n609), .B(n610), .Z(xin[287]) );
  NANDN U1430 ( .A(start), .B(xreg[287]), .Z(n610) );
  NAND U1431 ( .A(x[287]), .B(start), .Z(n609) );
  NAND U1432 ( .A(n611), .B(n612), .Z(xin[286]) );
  NANDN U1433 ( .A(start), .B(xreg[286]), .Z(n612) );
  NAND U1434 ( .A(x[286]), .B(start), .Z(n611) );
  NAND U1435 ( .A(n613), .B(n614), .Z(xin[285]) );
  NANDN U1436 ( .A(start), .B(xreg[285]), .Z(n614) );
  NAND U1437 ( .A(x[285]), .B(start), .Z(n613) );
  NAND U1438 ( .A(n615), .B(n616), .Z(xin[284]) );
  NANDN U1439 ( .A(start), .B(xreg[284]), .Z(n616) );
  NAND U1440 ( .A(x[284]), .B(start), .Z(n615) );
  NAND U1441 ( .A(n617), .B(n618), .Z(xin[283]) );
  NANDN U1442 ( .A(start), .B(xreg[283]), .Z(n618) );
  NAND U1443 ( .A(x[283]), .B(start), .Z(n617) );
  NAND U1444 ( .A(n619), .B(n620), .Z(xin[282]) );
  NANDN U1445 ( .A(start), .B(xreg[282]), .Z(n620) );
  NAND U1446 ( .A(x[282]), .B(start), .Z(n619) );
  NAND U1447 ( .A(n621), .B(n622), .Z(xin[281]) );
  NANDN U1448 ( .A(start), .B(xreg[281]), .Z(n622) );
  NAND U1449 ( .A(x[281]), .B(start), .Z(n621) );
  NAND U1450 ( .A(n623), .B(n624), .Z(xin[280]) );
  NANDN U1451 ( .A(start), .B(xreg[280]), .Z(n624) );
  NAND U1452 ( .A(x[280]), .B(start), .Z(n623) );
  NAND U1453 ( .A(n625), .B(n626), .Z(xin[27]) );
  NANDN U1454 ( .A(start), .B(xreg[27]), .Z(n626) );
  NAND U1455 ( .A(x[27]), .B(start), .Z(n625) );
  NAND U1456 ( .A(n627), .B(n628), .Z(xin[279]) );
  NANDN U1457 ( .A(start), .B(xreg[279]), .Z(n628) );
  NAND U1458 ( .A(x[279]), .B(start), .Z(n627) );
  NAND U1459 ( .A(n629), .B(n630), .Z(xin[278]) );
  NANDN U1460 ( .A(start), .B(xreg[278]), .Z(n630) );
  NAND U1461 ( .A(x[278]), .B(start), .Z(n629) );
  NAND U1462 ( .A(n631), .B(n632), .Z(xin[277]) );
  NANDN U1463 ( .A(start), .B(xreg[277]), .Z(n632) );
  NAND U1464 ( .A(x[277]), .B(start), .Z(n631) );
  NAND U1465 ( .A(n633), .B(n634), .Z(xin[276]) );
  NANDN U1466 ( .A(start), .B(xreg[276]), .Z(n634) );
  NAND U1467 ( .A(x[276]), .B(start), .Z(n633) );
  NAND U1468 ( .A(n635), .B(n636), .Z(xin[275]) );
  NANDN U1469 ( .A(start), .B(xreg[275]), .Z(n636) );
  NAND U1470 ( .A(x[275]), .B(start), .Z(n635) );
  NAND U1471 ( .A(n637), .B(n638), .Z(xin[274]) );
  NANDN U1472 ( .A(start), .B(xreg[274]), .Z(n638) );
  NAND U1473 ( .A(x[274]), .B(start), .Z(n637) );
  NAND U1474 ( .A(n639), .B(n640), .Z(xin[273]) );
  NANDN U1475 ( .A(start), .B(xreg[273]), .Z(n640) );
  NAND U1476 ( .A(x[273]), .B(start), .Z(n639) );
  NAND U1477 ( .A(n641), .B(n642), .Z(xin[272]) );
  NANDN U1478 ( .A(start), .B(xreg[272]), .Z(n642) );
  NAND U1479 ( .A(x[272]), .B(start), .Z(n641) );
  NAND U1480 ( .A(n643), .B(n644), .Z(xin[271]) );
  NANDN U1481 ( .A(start), .B(xreg[271]), .Z(n644) );
  NAND U1482 ( .A(x[271]), .B(start), .Z(n643) );
  NAND U1483 ( .A(n645), .B(n646), .Z(xin[270]) );
  NANDN U1484 ( .A(start), .B(xreg[270]), .Z(n646) );
  NAND U1485 ( .A(x[270]), .B(start), .Z(n645) );
  NAND U1486 ( .A(n647), .B(n648), .Z(xin[26]) );
  NANDN U1487 ( .A(start), .B(xreg[26]), .Z(n648) );
  NAND U1488 ( .A(x[26]), .B(start), .Z(n647) );
  NAND U1489 ( .A(n649), .B(n650), .Z(xin[269]) );
  NANDN U1490 ( .A(start), .B(xreg[269]), .Z(n650) );
  NAND U1491 ( .A(x[269]), .B(start), .Z(n649) );
  NAND U1492 ( .A(n651), .B(n652), .Z(xin[268]) );
  NANDN U1493 ( .A(start), .B(xreg[268]), .Z(n652) );
  NAND U1494 ( .A(x[268]), .B(start), .Z(n651) );
  NAND U1495 ( .A(n653), .B(n654), .Z(xin[267]) );
  NANDN U1496 ( .A(start), .B(xreg[267]), .Z(n654) );
  NAND U1497 ( .A(x[267]), .B(start), .Z(n653) );
  NAND U1498 ( .A(n655), .B(n656), .Z(xin[266]) );
  NANDN U1499 ( .A(start), .B(xreg[266]), .Z(n656) );
  NAND U1500 ( .A(x[266]), .B(start), .Z(n655) );
  NAND U1501 ( .A(n657), .B(n658), .Z(xin[265]) );
  NANDN U1502 ( .A(start), .B(xreg[265]), .Z(n658) );
  NAND U1503 ( .A(x[265]), .B(start), .Z(n657) );
  NAND U1504 ( .A(n659), .B(n660), .Z(xin[264]) );
  NANDN U1505 ( .A(start), .B(xreg[264]), .Z(n660) );
  NAND U1506 ( .A(x[264]), .B(start), .Z(n659) );
  NAND U1507 ( .A(n661), .B(n662), .Z(xin[263]) );
  NANDN U1508 ( .A(start), .B(xreg[263]), .Z(n662) );
  NAND U1509 ( .A(x[263]), .B(start), .Z(n661) );
  NAND U1510 ( .A(n663), .B(n664), .Z(xin[262]) );
  NANDN U1511 ( .A(start), .B(xreg[262]), .Z(n664) );
  NAND U1512 ( .A(x[262]), .B(start), .Z(n663) );
  NAND U1513 ( .A(n665), .B(n666), .Z(xin[261]) );
  NANDN U1514 ( .A(start), .B(xreg[261]), .Z(n666) );
  NAND U1515 ( .A(x[261]), .B(start), .Z(n665) );
  NAND U1516 ( .A(n667), .B(n668), .Z(xin[260]) );
  NANDN U1517 ( .A(start), .B(xreg[260]), .Z(n668) );
  NAND U1518 ( .A(x[260]), .B(start), .Z(n667) );
  NAND U1519 ( .A(n669), .B(n670), .Z(xin[25]) );
  NANDN U1520 ( .A(start), .B(xreg[25]), .Z(n670) );
  NAND U1521 ( .A(x[25]), .B(start), .Z(n669) );
  NAND U1522 ( .A(n671), .B(n672), .Z(xin[259]) );
  NANDN U1523 ( .A(start), .B(xreg[259]), .Z(n672) );
  NAND U1524 ( .A(x[259]), .B(start), .Z(n671) );
  NAND U1525 ( .A(n673), .B(n674), .Z(xin[258]) );
  NANDN U1526 ( .A(start), .B(xreg[258]), .Z(n674) );
  NAND U1527 ( .A(x[258]), .B(start), .Z(n673) );
  NAND U1528 ( .A(n675), .B(n676), .Z(xin[257]) );
  NANDN U1529 ( .A(start), .B(xreg[257]), .Z(n676) );
  NAND U1530 ( .A(x[257]), .B(start), .Z(n675) );
  NAND U1531 ( .A(n677), .B(n678), .Z(xin[256]) );
  NANDN U1532 ( .A(start), .B(xreg[256]), .Z(n678) );
  NAND U1533 ( .A(x[256]), .B(start), .Z(n677) );
  NAND U1534 ( .A(n679), .B(n680), .Z(xin[255]) );
  NANDN U1535 ( .A(start), .B(xreg[255]), .Z(n680) );
  NAND U1536 ( .A(x[255]), .B(start), .Z(n679) );
  NAND U1537 ( .A(n681), .B(n682), .Z(xin[254]) );
  NANDN U1538 ( .A(start), .B(xreg[254]), .Z(n682) );
  NAND U1539 ( .A(x[254]), .B(start), .Z(n681) );
  NAND U1540 ( .A(n683), .B(n684), .Z(xin[253]) );
  NANDN U1541 ( .A(start), .B(xreg[253]), .Z(n684) );
  NAND U1542 ( .A(x[253]), .B(start), .Z(n683) );
  NAND U1543 ( .A(n685), .B(n686), .Z(xin[252]) );
  NANDN U1544 ( .A(start), .B(xreg[252]), .Z(n686) );
  NAND U1545 ( .A(x[252]), .B(start), .Z(n685) );
  NAND U1546 ( .A(n687), .B(n688), .Z(xin[251]) );
  NANDN U1547 ( .A(start), .B(xreg[251]), .Z(n688) );
  NAND U1548 ( .A(x[251]), .B(start), .Z(n687) );
  NAND U1549 ( .A(n689), .B(n690), .Z(xin[250]) );
  NANDN U1550 ( .A(start), .B(xreg[250]), .Z(n690) );
  NAND U1551 ( .A(x[250]), .B(start), .Z(n689) );
  NAND U1552 ( .A(n691), .B(n692), .Z(xin[24]) );
  NANDN U1553 ( .A(start), .B(xreg[24]), .Z(n692) );
  NAND U1554 ( .A(x[24]), .B(start), .Z(n691) );
  NAND U1555 ( .A(n693), .B(n694), .Z(xin[249]) );
  NANDN U1556 ( .A(start), .B(xreg[249]), .Z(n694) );
  NAND U1557 ( .A(x[249]), .B(start), .Z(n693) );
  NAND U1558 ( .A(n695), .B(n696), .Z(xin[248]) );
  NANDN U1559 ( .A(start), .B(xreg[248]), .Z(n696) );
  NAND U1560 ( .A(x[248]), .B(start), .Z(n695) );
  NAND U1561 ( .A(n697), .B(n698), .Z(xin[247]) );
  NANDN U1562 ( .A(start), .B(xreg[247]), .Z(n698) );
  NAND U1563 ( .A(x[247]), .B(start), .Z(n697) );
  NAND U1564 ( .A(n699), .B(n700), .Z(xin[246]) );
  NANDN U1565 ( .A(start), .B(xreg[246]), .Z(n700) );
  NAND U1566 ( .A(x[246]), .B(start), .Z(n699) );
  NAND U1567 ( .A(n701), .B(n702), .Z(xin[245]) );
  NANDN U1568 ( .A(start), .B(xreg[245]), .Z(n702) );
  NAND U1569 ( .A(x[245]), .B(start), .Z(n701) );
  NAND U1570 ( .A(n703), .B(n704), .Z(xin[244]) );
  NANDN U1571 ( .A(start), .B(xreg[244]), .Z(n704) );
  NAND U1572 ( .A(x[244]), .B(start), .Z(n703) );
  NAND U1573 ( .A(n705), .B(n706), .Z(xin[243]) );
  NANDN U1574 ( .A(start), .B(xreg[243]), .Z(n706) );
  NAND U1575 ( .A(x[243]), .B(start), .Z(n705) );
  NAND U1576 ( .A(n707), .B(n708), .Z(xin[242]) );
  NANDN U1577 ( .A(start), .B(xreg[242]), .Z(n708) );
  NAND U1578 ( .A(x[242]), .B(start), .Z(n707) );
  NAND U1579 ( .A(n709), .B(n710), .Z(xin[241]) );
  NANDN U1580 ( .A(start), .B(xreg[241]), .Z(n710) );
  NAND U1581 ( .A(x[241]), .B(start), .Z(n709) );
  NAND U1582 ( .A(n711), .B(n712), .Z(xin[240]) );
  NANDN U1583 ( .A(start), .B(xreg[240]), .Z(n712) );
  NAND U1584 ( .A(x[240]), .B(start), .Z(n711) );
  NAND U1585 ( .A(n713), .B(n714), .Z(xin[23]) );
  NANDN U1586 ( .A(start), .B(xreg[23]), .Z(n714) );
  NAND U1587 ( .A(x[23]), .B(start), .Z(n713) );
  NAND U1588 ( .A(n715), .B(n716), .Z(xin[239]) );
  NANDN U1589 ( .A(start), .B(xreg[239]), .Z(n716) );
  NAND U1590 ( .A(x[239]), .B(start), .Z(n715) );
  NAND U1591 ( .A(n717), .B(n718), .Z(xin[238]) );
  NANDN U1592 ( .A(start), .B(xreg[238]), .Z(n718) );
  NAND U1593 ( .A(x[238]), .B(start), .Z(n717) );
  NAND U1594 ( .A(n719), .B(n720), .Z(xin[237]) );
  NANDN U1595 ( .A(start), .B(xreg[237]), .Z(n720) );
  NAND U1596 ( .A(x[237]), .B(start), .Z(n719) );
  NAND U1597 ( .A(n721), .B(n722), .Z(xin[236]) );
  NANDN U1598 ( .A(start), .B(xreg[236]), .Z(n722) );
  NAND U1599 ( .A(x[236]), .B(start), .Z(n721) );
  NAND U1600 ( .A(n723), .B(n724), .Z(xin[235]) );
  NANDN U1601 ( .A(start), .B(xreg[235]), .Z(n724) );
  NAND U1602 ( .A(x[235]), .B(start), .Z(n723) );
  NAND U1603 ( .A(n725), .B(n726), .Z(xin[234]) );
  NANDN U1604 ( .A(start), .B(xreg[234]), .Z(n726) );
  NAND U1605 ( .A(x[234]), .B(start), .Z(n725) );
  NAND U1606 ( .A(n727), .B(n728), .Z(xin[233]) );
  NANDN U1607 ( .A(start), .B(xreg[233]), .Z(n728) );
  NAND U1608 ( .A(x[233]), .B(start), .Z(n727) );
  NAND U1609 ( .A(n729), .B(n730), .Z(xin[232]) );
  NANDN U1610 ( .A(start), .B(xreg[232]), .Z(n730) );
  NAND U1611 ( .A(x[232]), .B(start), .Z(n729) );
  NAND U1612 ( .A(n731), .B(n732), .Z(xin[231]) );
  NANDN U1613 ( .A(start), .B(xreg[231]), .Z(n732) );
  NAND U1614 ( .A(x[231]), .B(start), .Z(n731) );
  NAND U1615 ( .A(n733), .B(n734), .Z(xin[230]) );
  NANDN U1616 ( .A(start), .B(xreg[230]), .Z(n734) );
  NAND U1617 ( .A(x[230]), .B(start), .Z(n733) );
  NAND U1618 ( .A(n735), .B(n736), .Z(xin[22]) );
  NANDN U1619 ( .A(start), .B(xreg[22]), .Z(n736) );
  NAND U1620 ( .A(x[22]), .B(start), .Z(n735) );
  NAND U1621 ( .A(n737), .B(n738), .Z(xin[229]) );
  NANDN U1622 ( .A(start), .B(xreg[229]), .Z(n738) );
  NAND U1623 ( .A(x[229]), .B(start), .Z(n737) );
  NAND U1624 ( .A(n739), .B(n740), .Z(xin[228]) );
  NANDN U1625 ( .A(start), .B(xreg[228]), .Z(n740) );
  NAND U1626 ( .A(x[228]), .B(start), .Z(n739) );
  NAND U1627 ( .A(n741), .B(n742), .Z(xin[227]) );
  NANDN U1628 ( .A(start), .B(xreg[227]), .Z(n742) );
  NAND U1629 ( .A(x[227]), .B(start), .Z(n741) );
  NAND U1630 ( .A(n743), .B(n744), .Z(xin[226]) );
  NANDN U1631 ( .A(start), .B(xreg[226]), .Z(n744) );
  NAND U1632 ( .A(x[226]), .B(start), .Z(n743) );
  NAND U1633 ( .A(n745), .B(n746), .Z(xin[225]) );
  NANDN U1634 ( .A(start), .B(xreg[225]), .Z(n746) );
  NAND U1635 ( .A(x[225]), .B(start), .Z(n745) );
  NAND U1636 ( .A(n747), .B(n748), .Z(xin[224]) );
  NANDN U1637 ( .A(start), .B(xreg[224]), .Z(n748) );
  NAND U1638 ( .A(x[224]), .B(start), .Z(n747) );
  NAND U1639 ( .A(n749), .B(n750), .Z(xin[223]) );
  NANDN U1640 ( .A(start), .B(xreg[223]), .Z(n750) );
  NAND U1641 ( .A(x[223]), .B(start), .Z(n749) );
  NAND U1642 ( .A(n751), .B(n752), .Z(xin[222]) );
  NANDN U1643 ( .A(start), .B(xreg[222]), .Z(n752) );
  NAND U1644 ( .A(x[222]), .B(start), .Z(n751) );
  NAND U1645 ( .A(n753), .B(n754), .Z(xin[221]) );
  NANDN U1646 ( .A(start), .B(xreg[221]), .Z(n754) );
  NAND U1647 ( .A(x[221]), .B(start), .Z(n753) );
  NAND U1648 ( .A(n755), .B(n756), .Z(xin[220]) );
  NANDN U1649 ( .A(start), .B(xreg[220]), .Z(n756) );
  NAND U1650 ( .A(x[220]), .B(start), .Z(n755) );
  NAND U1651 ( .A(n757), .B(n758), .Z(xin[21]) );
  NANDN U1652 ( .A(start), .B(xreg[21]), .Z(n758) );
  NAND U1653 ( .A(x[21]), .B(start), .Z(n757) );
  NAND U1654 ( .A(n759), .B(n760), .Z(xin[219]) );
  NANDN U1655 ( .A(start), .B(xreg[219]), .Z(n760) );
  NAND U1656 ( .A(x[219]), .B(start), .Z(n759) );
  NAND U1657 ( .A(n761), .B(n762), .Z(xin[218]) );
  NANDN U1658 ( .A(start), .B(xreg[218]), .Z(n762) );
  NAND U1659 ( .A(x[218]), .B(start), .Z(n761) );
  NAND U1660 ( .A(n763), .B(n764), .Z(xin[217]) );
  NANDN U1661 ( .A(start), .B(xreg[217]), .Z(n764) );
  NAND U1662 ( .A(x[217]), .B(start), .Z(n763) );
  NAND U1663 ( .A(n765), .B(n766), .Z(xin[216]) );
  NANDN U1664 ( .A(start), .B(xreg[216]), .Z(n766) );
  NAND U1665 ( .A(x[216]), .B(start), .Z(n765) );
  NAND U1666 ( .A(n767), .B(n768), .Z(xin[215]) );
  NANDN U1667 ( .A(start), .B(xreg[215]), .Z(n768) );
  NAND U1668 ( .A(x[215]), .B(start), .Z(n767) );
  NAND U1669 ( .A(n769), .B(n770), .Z(xin[214]) );
  NANDN U1670 ( .A(start), .B(xreg[214]), .Z(n770) );
  NAND U1671 ( .A(x[214]), .B(start), .Z(n769) );
  NAND U1672 ( .A(n771), .B(n772), .Z(xin[213]) );
  NANDN U1673 ( .A(start), .B(xreg[213]), .Z(n772) );
  NAND U1674 ( .A(x[213]), .B(start), .Z(n771) );
  NAND U1675 ( .A(n773), .B(n774), .Z(xin[212]) );
  NANDN U1676 ( .A(start), .B(xreg[212]), .Z(n774) );
  NAND U1677 ( .A(x[212]), .B(start), .Z(n773) );
  NAND U1678 ( .A(n775), .B(n776), .Z(xin[211]) );
  NANDN U1679 ( .A(start), .B(xreg[211]), .Z(n776) );
  NAND U1680 ( .A(x[211]), .B(start), .Z(n775) );
  NAND U1681 ( .A(n777), .B(n778), .Z(xin[210]) );
  NANDN U1682 ( .A(start), .B(xreg[210]), .Z(n778) );
  NAND U1683 ( .A(x[210]), .B(start), .Z(n777) );
  NAND U1684 ( .A(n779), .B(n780), .Z(xin[20]) );
  NANDN U1685 ( .A(start), .B(xreg[20]), .Z(n780) );
  NAND U1686 ( .A(x[20]), .B(start), .Z(n779) );
  NAND U1687 ( .A(n781), .B(n782), .Z(xin[209]) );
  NANDN U1688 ( .A(start), .B(xreg[209]), .Z(n782) );
  NAND U1689 ( .A(x[209]), .B(start), .Z(n781) );
  NAND U1690 ( .A(n783), .B(n784), .Z(xin[208]) );
  NANDN U1691 ( .A(start), .B(xreg[208]), .Z(n784) );
  NAND U1692 ( .A(x[208]), .B(start), .Z(n783) );
  NAND U1693 ( .A(n785), .B(n786), .Z(xin[207]) );
  NANDN U1694 ( .A(start), .B(xreg[207]), .Z(n786) );
  NAND U1695 ( .A(x[207]), .B(start), .Z(n785) );
  NAND U1696 ( .A(n787), .B(n788), .Z(xin[206]) );
  NANDN U1697 ( .A(start), .B(xreg[206]), .Z(n788) );
  NAND U1698 ( .A(x[206]), .B(start), .Z(n787) );
  NAND U1699 ( .A(n789), .B(n790), .Z(xin[205]) );
  NANDN U1700 ( .A(start), .B(xreg[205]), .Z(n790) );
  NAND U1701 ( .A(x[205]), .B(start), .Z(n789) );
  NAND U1702 ( .A(n791), .B(n792), .Z(xin[204]) );
  NANDN U1703 ( .A(start), .B(xreg[204]), .Z(n792) );
  NAND U1704 ( .A(x[204]), .B(start), .Z(n791) );
  NAND U1705 ( .A(n793), .B(n794), .Z(xin[203]) );
  NANDN U1706 ( .A(start), .B(xreg[203]), .Z(n794) );
  NAND U1707 ( .A(x[203]), .B(start), .Z(n793) );
  NAND U1708 ( .A(n795), .B(n796), .Z(xin[202]) );
  NANDN U1709 ( .A(start), .B(xreg[202]), .Z(n796) );
  NAND U1710 ( .A(x[202]), .B(start), .Z(n795) );
  NAND U1711 ( .A(n797), .B(n798), .Z(xin[201]) );
  NANDN U1712 ( .A(start), .B(xreg[201]), .Z(n798) );
  NAND U1713 ( .A(x[201]), .B(start), .Z(n797) );
  NAND U1714 ( .A(n799), .B(n800), .Z(xin[200]) );
  NANDN U1715 ( .A(start), .B(xreg[200]), .Z(n800) );
  NAND U1716 ( .A(x[200]), .B(start), .Z(n799) );
  NAND U1717 ( .A(n801), .B(n802), .Z(xin[1]) );
  NANDN U1718 ( .A(start), .B(xreg[1]), .Z(n802) );
  NAND U1719 ( .A(x[1]), .B(start), .Z(n801) );
  NAND U1720 ( .A(n803), .B(n804), .Z(xin[19]) );
  NANDN U1721 ( .A(start), .B(xreg[19]), .Z(n804) );
  NAND U1722 ( .A(x[19]), .B(start), .Z(n803) );
  NAND U1723 ( .A(n805), .B(n806), .Z(xin[199]) );
  NANDN U1724 ( .A(start), .B(xreg[199]), .Z(n806) );
  NAND U1725 ( .A(x[199]), .B(start), .Z(n805) );
  NAND U1726 ( .A(n807), .B(n808), .Z(xin[198]) );
  NANDN U1727 ( .A(start), .B(xreg[198]), .Z(n808) );
  NAND U1728 ( .A(x[198]), .B(start), .Z(n807) );
  NAND U1729 ( .A(n809), .B(n810), .Z(xin[197]) );
  NANDN U1730 ( .A(start), .B(xreg[197]), .Z(n810) );
  NAND U1731 ( .A(x[197]), .B(start), .Z(n809) );
  NAND U1732 ( .A(n811), .B(n812), .Z(xin[196]) );
  NANDN U1733 ( .A(start), .B(xreg[196]), .Z(n812) );
  NAND U1734 ( .A(x[196]), .B(start), .Z(n811) );
  NAND U1735 ( .A(n813), .B(n814), .Z(xin[195]) );
  NANDN U1736 ( .A(start), .B(xreg[195]), .Z(n814) );
  NAND U1737 ( .A(x[195]), .B(start), .Z(n813) );
  NAND U1738 ( .A(n815), .B(n816), .Z(xin[194]) );
  NANDN U1739 ( .A(start), .B(xreg[194]), .Z(n816) );
  NAND U1740 ( .A(x[194]), .B(start), .Z(n815) );
  NAND U1741 ( .A(n817), .B(n818), .Z(xin[193]) );
  NANDN U1742 ( .A(start), .B(xreg[193]), .Z(n818) );
  NAND U1743 ( .A(x[193]), .B(start), .Z(n817) );
  NAND U1744 ( .A(n819), .B(n820), .Z(xin[192]) );
  NANDN U1745 ( .A(start), .B(xreg[192]), .Z(n820) );
  NAND U1746 ( .A(x[192]), .B(start), .Z(n819) );
  NAND U1747 ( .A(n821), .B(n822), .Z(xin[191]) );
  NANDN U1748 ( .A(start), .B(xreg[191]), .Z(n822) );
  NAND U1749 ( .A(x[191]), .B(start), .Z(n821) );
  NAND U1750 ( .A(n823), .B(n824), .Z(xin[190]) );
  NANDN U1751 ( .A(start), .B(xreg[190]), .Z(n824) );
  NAND U1752 ( .A(x[190]), .B(start), .Z(n823) );
  NAND U1753 ( .A(n825), .B(n826), .Z(xin[18]) );
  NANDN U1754 ( .A(start), .B(xreg[18]), .Z(n826) );
  NAND U1755 ( .A(x[18]), .B(start), .Z(n825) );
  NAND U1756 ( .A(n827), .B(n828), .Z(xin[189]) );
  NANDN U1757 ( .A(start), .B(xreg[189]), .Z(n828) );
  NAND U1758 ( .A(x[189]), .B(start), .Z(n827) );
  NAND U1759 ( .A(n829), .B(n830), .Z(xin[188]) );
  NANDN U1760 ( .A(start), .B(xreg[188]), .Z(n830) );
  NAND U1761 ( .A(x[188]), .B(start), .Z(n829) );
  NAND U1762 ( .A(n831), .B(n832), .Z(xin[187]) );
  NANDN U1763 ( .A(start), .B(xreg[187]), .Z(n832) );
  NAND U1764 ( .A(x[187]), .B(start), .Z(n831) );
  NAND U1765 ( .A(n833), .B(n834), .Z(xin[186]) );
  NANDN U1766 ( .A(start), .B(xreg[186]), .Z(n834) );
  NAND U1767 ( .A(x[186]), .B(start), .Z(n833) );
  NAND U1768 ( .A(n835), .B(n836), .Z(xin[185]) );
  NANDN U1769 ( .A(start), .B(xreg[185]), .Z(n836) );
  NAND U1770 ( .A(x[185]), .B(start), .Z(n835) );
  NAND U1771 ( .A(n837), .B(n838), .Z(xin[184]) );
  NANDN U1772 ( .A(start), .B(xreg[184]), .Z(n838) );
  NAND U1773 ( .A(x[184]), .B(start), .Z(n837) );
  NAND U1774 ( .A(n839), .B(n840), .Z(xin[183]) );
  NANDN U1775 ( .A(start), .B(xreg[183]), .Z(n840) );
  NAND U1776 ( .A(x[183]), .B(start), .Z(n839) );
  NAND U1777 ( .A(n841), .B(n842), .Z(xin[182]) );
  NANDN U1778 ( .A(start), .B(xreg[182]), .Z(n842) );
  NAND U1779 ( .A(x[182]), .B(start), .Z(n841) );
  NAND U1780 ( .A(n843), .B(n844), .Z(xin[181]) );
  NANDN U1781 ( .A(start), .B(xreg[181]), .Z(n844) );
  NAND U1782 ( .A(x[181]), .B(start), .Z(n843) );
  NAND U1783 ( .A(n845), .B(n846), .Z(xin[180]) );
  NANDN U1784 ( .A(start), .B(xreg[180]), .Z(n846) );
  NAND U1785 ( .A(x[180]), .B(start), .Z(n845) );
  NAND U1786 ( .A(n847), .B(n848), .Z(xin[17]) );
  NANDN U1787 ( .A(start), .B(xreg[17]), .Z(n848) );
  NAND U1788 ( .A(x[17]), .B(start), .Z(n847) );
  NAND U1789 ( .A(n849), .B(n850), .Z(xin[179]) );
  NANDN U1790 ( .A(start), .B(xreg[179]), .Z(n850) );
  NAND U1791 ( .A(x[179]), .B(start), .Z(n849) );
  NAND U1792 ( .A(n851), .B(n852), .Z(xin[178]) );
  NANDN U1793 ( .A(start), .B(xreg[178]), .Z(n852) );
  NAND U1794 ( .A(x[178]), .B(start), .Z(n851) );
  NAND U1795 ( .A(n853), .B(n854), .Z(xin[177]) );
  NANDN U1796 ( .A(start), .B(xreg[177]), .Z(n854) );
  NAND U1797 ( .A(x[177]), .B(start), .Z(n853) );
  NAND U1798 ( .A(n855), .B(n856), .Z(xin[176]) );
  NANDN U1799 ( .A(start), .B(xreg[176]), .Z(n856) );
  NAND U1800 ( .A(x[176]), .B(start), .Z(n855) );
  NAND U1801 ( .A(n857), .B(n858), .Z(xin[175]) );
  NANDN U1802 ( .A(start), .B(xreg[175]), .Z(n858) );
  NAND U1803 ( .A(x[175]), .B(start), .Z(n857) );
  NAND U1804 ( .A(n859), .B(n860), .Z(xin[174]) );
  NANDN U1805 ( .A(start), .B(xreg[174]), .Z(n860) );
  NAND U1806 ( .A(x[174]), .B(start), .Z(n859) );
  NAND U1807 ( .A(n861), .B(n862), .Z(xin[173]) );
  NANDN U1808 ( .A(start), .B(xreg[173]), .Z(n862) );
  NAND U1809 ( .A(x[173]), .B(start), .Z(n861) );
  NAND U1810 ( .A(n863), .B(n864), .Z(xin[172]) );
  NANDN U1811 ( .A(start), .B(xreg[172]), .Z(n864) );
  NAND U1812 ( .A(x[172]), .B(start), .Z(n863) );
  NAND U1813 ( .A(n865), .B(n866), .Z(xin[171]) );
  NANDN U1814 ( .A(start), .B(xreg[171]), .Z(n866) );
  NAND U1815 ( .A(x[171]), .B(start), .Z(n865) );
  NAND U1816 ( .A(n867), .B(n868), .Z(xin[170]) );
  NANDN U1817 ( .A(start), .B(xreg[170]), .Z(n868) );
  NAND U1818 ( .A(x[170]), .B(start), .Z(n867) );
  NAND U1819 ( .A(n869), .B(n870), .Z(xin[16]) );
  NANDN U1820 ( .A(start), .B(xreg[16]), .Z(n870) );
  NAND U1821 ( .A(x[16]), .B(start), .Z(n869) );
  NAND U1822 ( .A(n871), .B(n872), .Z(xin[169]) );
  NANDN U1823 ( .A(start), .B(xreg[169]), .Z(n872) );
  NAND U1824 ( .A(x[169]), .B(start), .Z(n871) );
  NAND U1825 ( .A(n873), .B(n874), .Z(xin[168]) );
  NANDN U1826 ( .A(start), .B(xreg[168]), .Z(n874) );
  NAND U1827 ( .A(x[168]), .B(start), .Z(n873) );
  NAND U1828 ( .A(n875), .B(n876), .Z(xin[167]) );
  NANDN U1829 ( .A(start), .B(xreg[167]), .Z(n876) );
  NAND U1830 ( .A(x[167]), .B(start), .Z(n875) );
  NAND U1831 ( .A(n877), .B(n878), .Z(xin[166]) );
  NANDN U1832 ( .A(start), .B(xreg[166]), .Z(n878) );
  NAND U1833 ( .A(x[166]), .B(start), .Z(n877) );
  NAND U1834 ( .A(n879), .B(n880), .Z(xin[165]) );
  NANDN U1835 ( .A(start), .B(xreg[165]), .Z(n880) );
  NAND U1836 ( .A(x[165]), .B(start), .Z(n879) );
  NAND U1837 ( .A(n881), .B(n882), .Z(xin[164]) );
  NANDN U1838 ( .A(start), .B(xreg[164]), .Z(n882) );
  NAND U1839 ( .A(x[164]), .B(start), .Z(n881) );
  NAND U1840 ( .A(n883), .B(n884), .Z(xin[163]) );
  NANDN U1841 ( .A(start), .B(xreg[163]), .Z(n884) );
  NAND U1842 ( .A(x[163]), .B(start), .Z(n883) );
  NAND U1843 ( .A(n885), .B(n886), .Z(xin[162]) );
  NANDN U1844 ( .A(start), .B(xreg[162]), .Z(n886) );
  NAND U1845 ( .A(x[162]), .B(start), .Z(n885) );
  NAND U1846 ( .A(n887), .B(n888), .Z(xin[161]) );
  NANDN U1847 ( .A(start), .B(xreg[161]), .Z(n888) );
  NAND U1848 ( .A(x[161]), .B(start), .Z(n887) );
  NAND U1849 ( .A(n889), .B(n890), .Z(xin[160]) );
  NANDN U1850 ( .A(start), .B(xreg[160]), .Z(n890) );
  NAND U1851 ( .A(x[160]), .B(start), .Z(n889) );
  NAND U1852 ( .A(n891), .B(n892), .Z(xin[15]) );
  NANDN U1853 ( .A(start), .B(xreg[15]), .Z(n892) );
  NAND U1854 ( .A(x[15]), .B(start), .Z(n891) );
  NAND U1855 ( .A(n893), .B(n894), .Z(xin[159]) );
  NANDN U1856 ( .A(start), .B(xreg[159]), .Z(n894) );
  NAND U1857 ( .A(x[159]), .B(start), .Z(n893) );
  NAND U1858 ( .A(n895), .B(n896), .Z(xin[158]) );
  NANDN U1859 ( .A(start), .B(xreg[158]), .Z(n896) );
  NAND U1860 ( .A(x[158]), .B(start), .Z(n895) );
  NAND U1861 ( .A(n897), .B(n898), .Z(xin[157]) );
  NANDN U1862 ( .A(start), .B(xreg[157]), .Z(n898) );
  NAND U1863 ( .A(x[157]), .B(start), .Z(n897) );
  NAND U1864 ( .A(n899), .B(n900), .Z(xin[156]) );
  NANDN U1865 ( .A(start), .B(xreg[156]), .Z(n900) );
  NAND U1866 ( .A(x[156]), .B(start), .Z(n899) );
  NAND U1867 ( .A(n901), .B(n902), .Z(xin[155]) );
  NANDN U1868 ( .A(start), .B(xreg[155]), .Z(n902) );
  NAND U1869 ( .A(x[155]), .B(start), .Z(n901) );
  NAND U1870 ( .A(n903), .B(n904), .Z(xin[154]) );
  NANDN U1871 ( .A(start), .B(xreg[154]), .Z(n904) );
  NAND U1872 ( .A(x[154]), .B(start), .Z(n903) );
  NAND U1873 ( .A(n905), .B(n906), .Z(xin[153]) );
  NANDN U1874 ( .A(start), .B(xreg[153]), .Z(n906) );
  NAND U1875 ( .A(x[153]), .B(start), .Z(n905) );
  NAND U1876 ( .A(n907), .B(n908), .Z(xin[152]) );
  NANDN U1877 ( .A(start), .B(xreg[152]), .Z(n908) );
  NAND U1878 ( .A(x[152]), .B(start), .Z(n907) );
  NAND U1879 ( .A(n909), .B(n910), .Z(xin[151]) );
  NANDN U1880 ( .A(start), .B(xreg[151]), .Z(n910) );
  NAND U1881 ( .A(x[151]), .B(start), .Z(n909) );
  NAND U1882 ( .A(n911), .B(n912), .Z(xin[150]) );
  NANDN U1883 ( .A(start), .B(xreg[150]), .Z(n912) );
  NAND U1884 ( .A(x[150]), .B(start), .Z(n911) );
  NAND U1885 ( .A(n913), .B(n914), .Z(xin[14]) );
  NANDN U1886 ( .A(start), .B(xreg[14]), .Z(n914) );
  NAND U1887 ( .A(x[14]), .B(start), .Z(n913) );
  NAND U1888 ( .A(n915), .B(n916), .Z(xin[149]) );
  NANDN U1889 ( .A(start), .B(xreg[149]), .Z(n916) );
  NAND U1890 ( .A(x[149]), .B(start), .Z(n915) );
  NAND U1891 ( .A(n917), .B(n918), .Z(xin[148]) );
  NANDN U1892 ( .A(start), .B(xreg[148]), .Z(n918) );
  NAND U1893 ( .A(x[148]), .B(start), .Z(n917) );
  NAND U1894 ( .A(n919), .B(n920), .Z(xin[147]) );
  NANDN U1895 ( .A(start), .B(xreg[147]), .Z(n920) );
  NAND U1896 ( .A(x[147]), .B(start), .Z(n919) );
  NAND U1897 ( .A(n921), .B(n922), .Z(xin[146]) );
  NANDN U1898 ( .A(start), .B(xreg[146]), .Z(n922) );
  NAND U1899 ( .A(x[146]), .B(start), .Z(n921) );
  NAND U1900 ( .A(n923), .B(n924), .Z(xin[145]) );
  NANDN U1901 ( .A(start), .B(xreg[145]), .Z(n924) );
  NAND U1902 ( .A(x[145]), .B(start), .Z(n923) );
  NAND U1903 ( .A(n925), .B(n926), .Z(xin[144]) );
  NANDN U1904 ( .A(start), .B(xreg[144]), .Z(n926) );
  NAND U1905 ( .A(x[144]), .B(start), .Z(n925) );
  NAND U1906 ( .A(n927), .B(n928), .Z(xin[143]) );
  NANDN U1907 ( .A(start), .B(xreg[143]), .Z(n928) );
  NAND U1908 ( .A(x[143]), .B(start), .Z(n927) );
  NAND U1909 ( .A(n929), .B(n930), .Z(xin[142]) );
  NANDN U1910 ( .A(start), .B(xreg[142]), .Z(n930) );
  NAND U1911 ( .A(x[142]), .B(start), .Z(n929) );
  NAND U1912 ( .A(n931), .B(n932), .Z(xin[141]) );
  NANDN U1913 ( .A(start), .B(xreg[141]), .Z(n932) );
  NAND U1914 ( .A(x[141]), .B(start), .Z(n931) );
  NAND U1915 ( .A(n933), .B(n934), .Z(xin[140]) );
  NANDN U1916 ( .A(start), .B(xreg[140]), .Z(n934) );
  NAND U1917 ( .A(x[140]), .B(start), .Z(n933) );
  NAND U1918 ( .A(n935), .B(n936), .Z(xin[13]) );
  NANDN U1919 ( .A(start), .B(xreg[13]), .Z(n936) );
  NAND U1920 ( .A(x[13]), .B(start), .Z(n935) );
  NAND U1921 ( .A(n937), .B(n938), .Z(xin[139]) );
  NANDN U1922 ( .A(start), .B(xreg[139]), .Z(n938) );
  NAND U1923 ( .A(x[139]), .B(start), .Z(n937) );
  NAND U1924 ( .A(n939), .B(n940), .Z(xin[138]) );
  NANDN U1925 ( .A(start), .B(xreg[138]), .Z(n940) );
  NAND U1926 ( .A(x[138]), .B(start), .Z(n939) );
  NAND U1927 ( .A(n941), .B(n942), .Z(xin[137]) );
  NANDN U1928 ( .A(start), .B(xreg[137]), .Z(n942) );
  NAND U1929 ( .A(x[137]), .B(start), .Z(n941) );
  NAND U1930 ( .A(n943), .B(n944), .Z(xin[136]) );
  NANDN U1931 ( .A(start), .B(xreg[136]), .Z(n944) );
  NAND U1932 ( .A(x[136]), .B(start), .Z(n943) );
  NAND U1933 ( .A(n945), .B(n946), .Z(xin[135]) );
  NANDN U1934 ( .A(start), .B(xreg[135]), .Z(n946) );
  NAND U1935 ( .A(x[135]), .B(start), .Z(n945) );
  NAND U1936 ( .A(n947), .B(n948), .Z(xin[134]) );
  NANDN U1937 ( .A(start), .B(xreg[134]), .Z(n948) );
  NAND U1938 ( .A(x[134]), .B(start), .Z(n947) );
  NAND U1939 ( .A(n949), .B(n950), .Z(xin[133]) );
  NANDN U1940 ( .A(start), .B(xreg[133]), .Z(n950) );
  NAND U1941 ( .A(x[133]), .B(start), .Z(n949) );
  NAND U1942 ( .A(n951), .B(n952), .Z(xin[132]) );
  NANDN U1943 ( .A(start), .B(xreg[132]), .Z(n952) );
  NAND U1944 ( .A(x[132]), .B(start), .Z(n951) );
  NAND U1945 ( .A(n953), .B(n954), .Z(xin[131]) );
  NANDN U1946 ( .A(start), .B(xreg[131]), .Z(n954) );
  NAND U1947 ( .A(x[131]), .B(start), .Z(n953) );
  NAND U1948 ( .A(n955), .B(n956), .Z(xin[130]) );
  NANDN U1949 ( .A(start), .B(xreg[130]), .Z(n956) );
  NAND U1950 ( .A(x[130]), .B(start), .Z(n955) );
  NAND U1951 ( .A(n957), .B(n958), .Z(xin[12]) );
  NANDN U1952 ( .A(start), .B(xreg[12]), .Z(n958) );
  NAND U1953 ( .A(x[12]), .B(start), .Z(n957) );
  NAND U1954 ( .A(n959), .B(n960), .Z(xin[129]) );
  NANDN U1955 ( .A(start), .B(xreg[129]), .Z(n960) );
  NAND U1956 ( .A(x[129]), .B(start), .Z(n959) );
  NAND U1957 ( .A(n961), .B(n962), .Z(xin[128]) );
  NANDN U1958 ( .A(start), .B(xreg[128]), .Z(n962) );
  NAND U1959 ( .A(x[128]), .B(start), .Z(n961) );
  NAND U1960 ( .A(n963), .B(n964), .Z(xin[127]) );
  NANDN U1961 ( .A(start), .B(xreg[127]), .Z(n964) );
  NAND U1962 ( .A(x[127]), .B(start), .Z(n963) );
  NAND U1963 ( .A(n965), .B(n966), .Z(xin[126]) );
  NANDN U1964 ( .A(start), .B(xreg[126]), .Z(n966) );
  NAND U1965 ( .A(x[126]), .B(start), .Z(n965) );
  NAND U1966 ( .A(n967), .B(n968), .Z(xin[125]) );
  NANDN U1967 ( .A(start), .B(xreg[125]), .Z(n968) );
  NAND U1968 ( .A(x[125]), .B(start), .Z(n967) );
  NAND U1969 ( .A(n969), .B(n970), .Z(xin[124]) );
  NANDN U1970 ( .A(start), .B(xreg[124]), .Z(n970) );
  NAND U1971 ( .A(x[124]), .B(start), .Z(n969) );
  NAND U1972 ( .A(n971), .B(n972), .Z(xin[123]) );
  NANDN U1973 ( .A(start), .B(xreg[123]), .Z(n972) );
  NAND U1974 ( .A(x[123]), .B(start), .Z(n971) );
  NAND U1975 ( .A(n973), .B(n974), .Z(xin[122]) );
  NANDN U1976 ( .A(start), .B(xreg[122]), .Z(n974) );
  NAND U1977 ( .A(x[122]), .B(start), .Z(n973) );
  NAND U1978 ( .A(n975), .B(n976), .Z(xin[121]) );
  NANDN U1979 ( .A(start), .B(xreg[121]), .Z(n976) );
  NAND U1980 ( .A(x[121]), .B(start), .Z(n975) );
  NAND U1981 ( .A(n977), .B(n978), .Z(xin[120]) );
  NANDN U1982 ( .A(start), .B(xreg[120]), .Z(n978) );
  NAND U1983 ( .A(x[120]), .B(start), .Z(n977) );
  NAND U1984 ( .A(n979), .B(n980), .Z(xin[11]) );
  NANDN U1985 ( .A(start), .B(xreg[11]), .Z(n980) );
  NAND U1986 ( .A(x[11]), .B(start), .Z(n979) );
  NAND U1987 ( .A(n981), .B(n982), .Z(xin[119]) );
  NANDN U1988 ( .A(start), .B(xreg[119]), .Z(n982) );
  NAND U1989 ( .A(x[119]), .B(start), .Z(n981) );
  NAND U1990 ( .A(n983), .B(n984), .Z(xin[118]) );
  NANDN U1991 ( .A(start), .B(xreg[118]), .Z(n984) );
  NAND U1992 ( .A(x[118]), .B(start), .Z(n983) );
  NAND U1993 ( .A(n985), .B(n986), .Z(xin[117]) );
  NANDN U1994 ( .A(start), .B(xreg[117]), .Z(n986) );
  NAND U1995 ( .A(x[117]), .B(start), .Z(n985) );
  NAND U1996 ( .A(n987), .B(n988), .Z(xin[116]) );
  NANDN U1997 ( .A(start), .B(xreg[116]), .Z(n988) );
  NAND U1998 ( .A(x[116]), .B(start), .Z(n987) );
  NAND U1999 ( .A(n989), .B(n990), .Z(xin[115]) );
  NANDN U2000 ( .A(start), .B(xreg[115]), .Z(n990) );
  NAND U2001 ( .A(x[115]), .B(start), .Z(n989) );
  NAND U2002 ( .A(n991), .B(n992), .Z(xin[114]) );
  NANDN U2003 ( .A(start), .B(xreg[114]), .Z(n992) );
  NAND U2004 ( .A(x[114]), .B(start), .Z(n991) );
  NAND U2005 ( .A(n993), .B(n994), .Z(xin[113]) );
  NANDN U2006 ( .A(start), .B(xreg[113]), .Z(n994) );
  NAND U2007 ( .A(x[113]), .B(start), .Z(n993) );
  NAND U2008 ( .A(n995), .B(n996), .Z(xin[112]) );
  NANDN U2009 ( .A(start), .B(xreg[112]), .Z(n996) );
  NAND U2010 ( .A(x[112]), .B(start), .Z(n995) );
  NAND U2011 ( .A(n997), .B(n998), .Z(xin[111]) );
  NANDN U2012 ( .A(start), .B(xreg[111]), .Z(n998) );
  NAND U2013 ( .A(x[111]), .B(start), .Z(n997) );
  NAND U2014 ( .A(n999), .B(n1000), .Z(xin[110]) );
  NANDN U2015 ( .A(start), .B(xreg[110]), .Z(n1000) );
  NAND U2016 ( .A(x[110]), .B(start), .Z(n999) );
  NAND U2017 ( .A(n1001), .B(n1002), .Z(xin[10]) );
  NANDN U2018 ( .A(start), .B(xreg[10]), .Z(n1002) );
  NAND U2019 ( .A(x[10]), .B(start), .Z(n1001) );
  NAND U2020 ( .A(n1003), .B(n1004), .Z(xin[109]) );
  NANDN U2021 ( .A(start), .B(xreg[109]), .Z(n1004) );
  NAND U2022 ( .A(x[109]), .B(start), .Z(n1003) );
  NAND U2023 ( .A(n1005), .B(n1006), .Z(xin[108]) );
  NANDN U2024 ( .A(start), .B(xreg[108]), .Z(n1006) );
  NAND U2025 ( .A(x[108]), .B(start), .Z(n1005) );
  NAND U2026 ( .A(n1007), .B(n1008), .Z(xin[107]) );
  NANDN U2027 ( .A(start), .B(xreg[107]), .Z(n1008) );
  NAND U2028 ( .A(x[107]), .B(start), .Z(n1007) );
  NAND U2029 ( .A(n1009), .B(n1010), .Z(xin[106]) );
  NANDN U2030 ( .A(start), .B(xreg[106]), .Z(n1010) );
  NAND U2031 ( .A(x[106]), .B(start), .Z(n1009) );
  NAND U2032 ( .A(n1011), .B(n1012), .Z(xin[105]) );
  NANDN U2033 ( .A(start), .B(xreg[105]), .Z(n1012) );
  NAND U2034 ( .A(x[105]), .B(start), .Z(n1011) );
  NAND U2035 ( .A(n1013), .B(n1014), .Z(xin[104]) );
  NANDN U2036 ( .A(start), .B(xreg[104]), .Z(n1014) );
  NAND U2037 ( .A(x[104]), .B(start), .Z(n1013) );
  NAND U2038 ( .A(n1015), .B(n1016), .Z(xin[103]) );
  NANDN U2039 ( .A(start), .B(xreg[103]), .Z(n1016) );
  NAND U2040 ( .A(x[103]), .B(start), .Z(n1015) );
  NAND U2041 ( .A(n1017), .B(n1018), .Z(xin[102]) );
  NANDN U2042 ( .A(start), .B(xreg[102]), .Z(n1018) );
  NAND U2043 ( .A(x[102]), .B(start), .Z(n1017) );
  NAND U2044 ( .A(n1019), .B(n1020), .Z(xin[101]) );
  NANDN U2045 ( .A(start), .B(xreg[101]), .Z(n1020) );
  NAND U2046 ( .A(x[101]), .B(start), .Z(n1019) );
  NAND U2047 ( .A(n1021), .B(n1022), .Z(xin[100]) );
  NANDN U2048 ( .A(start), .B(xreg[100]), .Z(n1022) );
  NAND U2049 ( .A(x[100]), .B(start), .Z(n1021) );
  AND U2050 ( .A(x[0]), .B(start), .Z(n1023) );
endmodule


module modexp_2N_NN_N512_CC524288 ( clk, rst, m, e, n, c );
  input [511:0] m;
  input [511:0] e;
  input [511:0] n;
  output [511:0] c;
  input clk, rst;
  wire   init, mul_pow, first_one, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
         n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
         n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
         n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
         n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
         n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
         n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
         n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
         n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
         n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
         n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
         n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
         n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
         n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
         n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
         n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
         n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
         n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
         n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
         n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
         n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
         n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
         n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
         n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
         n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
         n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
         n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
         n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
         n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
         n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
         n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
         n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429,
         n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
         n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
         n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
         n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
         n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
         n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
         n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
         n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
         n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
         n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
         n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
         n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
         n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
         n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
         n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
         n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
         n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
         n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
         n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
         n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
         n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
         n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
         n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
         n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
         n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
         n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
         n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
         n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
         n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
         n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
         n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
         n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
         n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
         n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
         n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
         n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019,
         n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029,
         n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
         n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
         n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
         n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
         n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
         n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
         n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
         n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
         n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
         n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
         n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
         n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
         n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
         n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
         n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
         n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
         n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
         n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
         n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239,
         n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
         n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259,
         n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269,
         n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
         n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289,
         n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299,
         n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309,
         n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319,
         n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329,
         n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339,
         n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349,
         n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359,
         n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369,
         n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379,
         n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389,
         n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399,
         n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409,
         n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419,
         n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429,
         n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439,
         n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449,
         n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459,
         n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469,
         n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479,
         n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489,
         n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499,
         n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509,
         n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519,
         n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529,
         n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539,
         n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549,
         n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559,
         n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569,
         n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579,
         n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
         n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
         n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
         n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
         n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
         n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
         n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
         n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
         n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
         n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
         n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
         n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
         n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
         n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
         n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
         n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
         n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
         n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
         n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
         n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951,
         n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
         n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967,
         n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975,
         n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983,
         n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
         n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999,
         n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
         n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015,
         n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023,
         n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
         n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
         n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047,
         n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055,
         n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063,
         n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071,
         n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079,
         n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087,
         n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095,
         n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103,
         n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111,
         n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119,
         n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127,
         n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135,
         n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143,
         n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151,
         n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159,
         n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167,
         n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175,
         n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183,
         n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191,
         n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199,
         n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207,
         n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215,
         n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223,
         n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231,
         n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239,
         n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247,
         n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255,
         n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263,
         n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271,
         n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279,
         n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287,
         n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295,
         n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303,
         n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311,
         n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319,
         n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327,
         n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335,
         n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343,
         n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351,
         n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359,
         n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367,
         n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375,
         n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383,
         n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391,
         n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399,
         n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407,
         n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415,
         n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423,
         n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431,
         n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439,
         n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447,
         n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455,
         n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463,
         n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471,
         n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479,
         n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487,
         n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495,
         n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503,
         n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511,
         n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519,
         n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527,
         n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535,
         n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543,
         n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551,
         n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559,
         n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567,
         n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575,
         n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583,
         n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591,
         n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599,
         n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607,
         n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615,
         n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623,
         n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631,
         n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639,
         n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647,
         n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655,
         n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663,
         n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671,
         n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679,
         n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687,
         n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695,
         n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703,
         n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711,
         n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719,
         n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727,
         n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735,
         n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743,
         n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751,
         n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759,
         n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767,
         n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775,
         n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783,
         n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791,
         n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799,
         n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807,
         n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815,
         n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823,
         n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831,
         n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839,
         n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847,
         n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855,
         n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863,
         n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871,
         n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879,
         n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887,
         n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895,
         n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903,
         n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911,
         n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919,
         n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927,
         n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935,
         n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943,
         n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951,
         n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959,
         n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967,
         n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975,
         n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983,
         n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991,
         n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999,
         n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007,
         n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015,
         n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023,
         n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031,
         n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039,
         n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047,
         n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055,
         n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063,
         n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071,
         n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079,
         n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087,
         n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095,
         n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103,
         n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111,
         n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119,
         n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127,
         n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135,
         n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143,
         n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151,
         n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159,
         n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167,
         n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175,
         n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183,
         n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191,
         n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199,
         n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207,
         n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215,
         n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223,
         n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231,
         n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239,
         n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247,
         n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255,
         n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263,
         n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271,
         n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279,
         n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287,
         n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295,
         n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303,
         n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311,
         n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319,
         n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327,
         n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335,
         n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343,
         n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351,
         n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359,
         n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367,
         n14368, n14369, n14370, n14371, n14372;
  wire   [511:0] start_in;
  wire   [511:0] start_reg;
  wire   [511:0] ereg;
  wire   [511:0] o;
  wire   [511:0] creg;
  wire   [511:0] x;
  wire   [511:0] y;

  DFF init_reg ( .D(1'b1), .CLK(clk), .RST(rst), .Q(init) );
  DFF \start_reg_reg[0]  ( .D(n14372), .CLK(clk), .RST(rst), .Q(start_reg[0])
         );
  DFF \start_reg_reg[1]  ( .D(start_in[0]), .CLK(clk), .RST(rst), .Q(
        start_reg[1]) );
  DFF \start_reg_reg[2]  ( .D(start_in[1]), .CLK(clk), .RST(rst), .Q(
        start_reg[2]) );
  DFF \start_reg_reg[3]  ( .D(start_in[2]), .CLK(clk), .RST(rst), .Q(
        start_reg[3]) );
  DFF \start_reg_reg[4]  ( .D(start_in[3]), .CLK(clk), .RST(rst), .Q(
        start_reg[4]) );
  DFF \start_reg_reg[5]  ( .D(start_in[4]), .CLK(clk), .RST(rst), .Q(
        start_reg[5]) );
  DFF \start_reg_reg[6]  ( .D(start_in[5]), .CLK(clk), .RST(rst), .Q(
        start_reg[6]) );
  DFF \start_reg_reg[7]  ( .D(start_in[6]), .CLK(clk), .RST(rst), .Q(
        start_reg[7]) );
  DFF \start_reg_reg[8]  ( .D(start_in[7]), .CLK(clk), .RST(rst), .Q(
        start_reg[8]) );
  DFF \start_reg_reg[9]  ( .D(start_in[8]), .CLK(clk), .RST(rst), .Q(
        start_reg[9]) );
  DFF \start_reg_reg[10]  ( .D(start_in[9]), .CLK(clk), .RST(rst), .Q(
        start_reg[10]) );
  DFF \start_reg_reg[11]  ( .D(start_in[10]), .CLK(clk), .RST(rst), .Q(
        start_reg[11]) );
  DFF \start_reg_reg[12]  ( .D(start_in[11]), .CLK(clk), .RST(rst), .Q(
        start_reg[12]) );
  DFF \start_reg_reg[13]  ( .D(start_in[12]), .CLK(clk), .RST(rst), .Q(
        start_reg[13]) );
  DFF \start_reg_reg[14]  ( .D(start_in[13]), .CLK(clk), .RST(rst), .Q(
        start_reg[14]) );
  DFF \start_reg_reg[15]  ( .D(start_in[14]), .CLK(clk), .RST(rst), .Q(
        start_reg[15]) );
  DFF \start_reg_reg[16]  ( .D(start_in[15]), .CLK(clk), .RST(rst), .Q(
        start_reg[16]) );
  DFF \start_reg_reg[17]  ( .D(start_in[16]), .CLK(clk), .RST(rst), .Q(
        start_reg[17]) );
  DFF \start_reg_reg[18]  ( .D(start_in[17]), .CLK(clk), .RST(rst), .Q(
        start_reg[18]) );
  DFF \start_reg_reg[19]  ( .D(start_in[18]), .CLK(clk), .RST(rst), .Q(
        start_reg[19]) );
  DFF \start_reg_reg[20]  ( .D(start_in[19]), .CLK(clk), .RST(rst), .Q(
        start_reg[20]) );
  DFF \start_reg_reg[21]  ( .D(start_in[20]), .CLK(clk), .RST(rst), .Q(
        start_reg[21]) );
  DFF \start_reg_reg[22]  ( .D(start_in[21]), .CLK(clk), .RST(rst), .Q(
        start_reg[22]) );
  DFF \start_reg_reg[23]  ( .D(start_in[22]), .CLK(clk), .RST(rst), .Q(
        start_reg[23]) );
  DFF \start_reg_reg[24]  ( .D(start_in[23]), .CLK(clk), .RST(rst), .Q(
        start_reg[24]) );
  DFF \start_reg_reg[25]  ( .D(start_in[24]), .CLK(clk), .RST(rst), .Q(
        start_reg[25]) );
  DFF \start_reg_reg[26]  ( .D(start_in[25]), .CLK(clk), .RST(rst), .Q(
        start_reg[26]) );
  DFF \start_reg_reg[27]  ( .D(start_in[26]), .CLK(clk), .RST(rst), .Q(
        start_reg[27]) );
  DFF \start_reg_reg[28]  ( .D(start_in[27]), .CLK(clk), .RST(rst), .Q(
        start_reg[28]) );
  DFF \start_reg_reg[29]  ( .D(start_in[28]), .CLK(clk), .RST(rst), .Q(
        start_reg[29]) );
  DFF \start_reg_reg[30]  ( .D(start_in[29]), .CLK(clk), .RST(rst), .Q(
        start_reg[30]) );
  DFF \start_reg_reg[31]  ( .D(start_in[30]), .CLK(clk), .RST(rst), .Q(
        start_reg[31]) );
  DFF \start_reg_reg[32]  ( .D(start_in[31]), .CLK(clk), .RST(rst), .Q(
        start_reg[32]) );
  DFF \start_reg_reg[33]  ( .D(start_in[32]), .CLK(clk), .RST(rst), .Q(
        start_reg[33]) );
  DFF \start_reg_reg[34]  ( .D(start_in[33]), .CLK(clk), .RST(rst), .Q(
        start_reg[34]) );
  DFF \start_reg_reg[35]  ( .D(start_in[34]), .CLK(clk), .RST(rst), .Q(
        start_reg[35]) );
  DFF \start_reg_reg[36]  ( .D(start_in[35]), .CLK(clk), .RST(rst), .Q(
        start_reg[36]) );
  DFF \start_reg_reg[37]  ( .D(start_in[36]), .CLK(clk), .RST(rst), .Q(
        start_reg[37]) );
  DFF \start_reg_reg[38]  ( .D(start_in[37]), .CLK(clk), .RST(rst), .Q(
        start_reg[38]) );
  DFF \start_reg_reg[39]  ( .D(start_in[38]), .CLK(clk), .RST(rst), .Q(
        start_reg[39]) );
  DFF \start_reg_reg[40]  ( .D(start_in[39]), .CLK(clk), .RST(rst), .Q(
        start_reg[40]) );
  DFF \start_reg_reg[41]  ( .D(start_in[40]), .CLK(clk), .RST(rst), .Q(
        start_reg[41]) );
  DFF \start_reg_reg[42]  ( .D(start_in[41]), .CLK(clk), .RST(rst), .Q(
        start_reg[42]) );
  DFF \start_reg_reg[43]  ( .D(start_in[42]), .CLK(clk), .RST(rst), .Q(
        start_reg[43]) );
  DFF \start_reg_reg[44]  ( .D(start_in[43]), .CLK(clk), .RST(rst), .Q(
        start_reg[44]) );
  DFF \start_reg_reg[45]  ( .D(start_in[44]), .CLK(clk), .RST(rst), .Q(
        start_reg[45]) );
  DFF \start_reg_reg[46]  ( .D(start_in[45]), .CLK(clk), .RST(rst), .Q(
        start_reg[46]) );
  DFF \start_reg_reg[47]  ( .D(start_in[46]), .CLK(clk), .RST(rst), .Q(
        start_reg[47]) );
  DFF \start_reg_reg[48]  ( .D(start_in[47]), .CLK(clk), .RST(rst), .Q(
        start_reg[48]) );
  DFF \start_reg_reg[49]  ( .D(start_in[48]), .CLK(clk), .RST(rst), .Q(
        start_reg[49]) );
  DFF \start_reg_reg[50]  ( .D(start_in[49]), .CLK(clk), .RST(rst), .Q(
        start_reg[50]) );
  DFF \start_reg_reg[51]  ( .D(start_in[50]), .CLK(clk), .RST(rst), .Q(
        start_reg[51]) );
  DFF \start_reg_reg[52]  ( .D(start_in[51]), .CLK(clk), .RST(rst), .Q(
        start_reg[52]) );
  DFF \start_reg_reg[53]  ( .D(start_in[52]), .CLK(clk), .RST(rst), .Q(
        start_reg[53]) );
  DFF \start_reg_reg[54]  ( .D(start_in[53]), .CLK(clk), .RST(rst), .Q(
        start_reg[54]) );
  DFF \start_reg_reg[55]  ( .D(start_in[54]), .CLK(clk), .RST(rst), .Q(
        start_reg[55]) );
  DFF \start_reg_reg[56]  ( .D(start_in[55]), .CLK(clk), .RST(rst), .Q(
        start_reg[56]) );
  DFF \start_reg_reg[57]  ( .D(start_in[56]), .CLK(clk), .RST(rst), .Q(
        start_reg[57]) );
  DFF \start_reg_reg[58]  ( .D(start_in[57]), .CLK(clk), .RST(rst), .Q(
        start_reg[58]) );
  DFF \start_reg_reg[59]  ( .D(start_in[58]), .CLK(clk), .RST(rst), .Q(
        start_reg[59]) );
  DFF \start_reg_reg[60]  ( .D(start_in[59]), .CLK(clk), .RST(rst), .Q(
        start_reg[60]) );
  DFF \start_reg_reg[61]  ( .D(start_in[60]), .CLK(clk), .RST(rst), .Q(
        start_reg[61]) );
  DFF \start_reg_reg[62]  ( .D(start_in[61]), .CLK(clk), .RST(rst), .Q(
        start_reg[62]) );
  DFF \start_reg_reg[63]  ( .D(start_in[62]), .CLK(clk), .RST(rst), .Q(
        start_reg[63]) );
  DFF \start_reg_reg[64]  ( .D(start_in[63]), .CLK(clk), .RST(rst), .Q(
        start_reg[64]) );
  DFF \start_reg_reg[65]  ( .D(start_in[64]), .CLK(clk), .RST(rst), .Q(
        start_reg[65]) );
  DFF \start_reg_reg[66]  ( .D(start_in[65]), .CLK(clk), .RST(rst), .Q(
        start_reg[66]) );
  DFF \start_reg_reg[67]  ( .D(start_in[66]), .CLK(clk), .RST(rst), .Q(
        start_reg[67]) );
  DFF \start_reg_reg[68]  ( .D(start_in[67]), .CLK(clk), .RST(rst), .Q(
        start_reg[68]) );
  DFF \start_reg_reg[69]  ( .D(start_in[68]), .CLK(clk), .RST(rst), .Q(
        start_reg[69]) );
  DFF \start_reg_reg[70]  ( .D(start_in[69]), .CLK(clk), .RST(rst), .Q(
        start_reg[70]) );
  DFF \start_reg_reg[71]  ( .D(start_in[70]), .CLK(clk), .RST(rst), .Q(
        start_reg[71]) );
  DFF \start_reg_reg[72]  ( .D(start_in[71]), .CLK(clk), .RST(rst), .Q(
        start_reg[72]) );
  DFF \start_reg_reg[73]  ( .D(start_in[72]), .CLK(clk), .RST(rst), .Q(
        start_reg[73]) );
  DFF \start_reg_reg[74]  ( .D(start_in[73]), .CLK(clk), .RST(rst), .Q(
        start_reg[74]) );
  DFF \start_reg_reg[75]  ( .D(start_in[74]), .CLK(clk), .RST(rst), .Q(
        start_reg[75]) );
  DFF \start_reg_reg[76]  ( .D(start_in[75]), .CLK(clk), .RST(rst), .Q(
        start_reg[76]) );
  DFF \start_reg_reg[77]  ( .D(start_in[76]), .CLK(clk), .RST(rst), .Q(
        start_reg[77]) );
  DFF \start_reg_reg[78]  ( .D(start_in[77]), .CLK(clk), .RST(rst), .Q(
        start_reg[78]) );
  DFF \start_reg_reg[79]  ( .D(start_in[78]), .CLK(clk), .RST(rst), .Q(
        start_reg[79]) );
  DFF \start_reg_reg[80]  ( .D(start_in[79]), .CLK(clk), .RST(rst), .Q(
        start_reg[80]) );
  DFF \start_reg_reg[81]  ( .D(start_in[80]), .CLK(clk), .RST(rst), .Q(
        start_reg[81]) );
  DFF \start_reg_reg[82]  ( .D(start_in[81]), .CLK(clk), .RST(rst), .Q(
        start_reg[82]) );
  DFF \start_reg_reg[83]  ( .D(start_in[82]), .CLK(clk), .RST(rst), .Q(
        start_reg[83]) );
  DFF \start_reg_reg[84]  ( .D(start_in[83]), .CLK(clk), .RST(rst), .Q(
        start_reg[84]) );
  DFF \start_reg_reg[85]  ( .D(start_in[84]), .CLK(clk), .RST(rst), .Q(
        start_reg[85]) );
  DFF \start_reg_reg[86]  ( .D(start_in[85]), .CLK(clk), .RST(rst), .Q(
        start_reg[86]) );
  DFF \start_reg_reg[87]  ( .D(start_in[86]), .CLK(clk), .RST(rst), .Q(
        start_reg[87]) );
  DFF \start_reg_reg[88]  ( .D(start_in[87]), .CLK(clk), .RST(rst), .Q(
        start_reg[88]) );
  DFF \start_reg_reg[89]  ( .D(start_in[88]), .CLK(clk), .RST(rst), .Q(
        start_reg[89]) );
  DFF \start_reg_reg[90]  ( .D(start_in[89]), .CLK(clk), .RST(rst), .Q(
        start_reg[90]) );
  DFF \start_reg_reg[91]  ( .D(start_in[90]), .CLK(clk), .RST(rst), .Q(
        start_reg[91]) );
  DFF \start_reg_reg[92]  ( .D(start_in[91]), .CLK(clk), .RST(rst), .Q(
        start_reg[92]) );
  DFF \start_reg_reg[93]  ( .D(start_in[92]), .CLK(clk), .RST(rst), .Q(
        start_reg[93]) );
  DFF \start_reg_reg[94]  ( .D(start_in[93]), .CLK(clk), .RST(rst), .Q(
        start_reg[94]) );
  DFF \start_reg_reg[95]  ( .D(start_in[94]), .CLK(clk), .RST(rst), .Q(
        start_reg[95]) );
  DFF \start_reg_reg[96]  ( .D(start_in[95]), .CLK(clk), .RST(rst), .Q(
        start_reg[96]) );
  DFF \start_reg_reg[97]  ( .D(start_in[96]), .CLK(clk), .RST(rst), .Q(
        start_reg[97]) );
  DFF \start_reg_reg[98]  ( .D(start_in[97]), .CLK(clk), .RST(rst), .Q(
        start_reg[98]) );
  DFF \start_reg_reg[99]  ( .D(start_in[98]), .CLK(clk), .RST(rst), .Q(
        start_reg[99]) );
  DFF \start_reg_reg[100]  ( .D(start_in[99]), .CLK(clk), .RST(rst), .Q(
        start_reg[100]) );
  DFF \start_reg_reg[101]  ( .D(start_in[100]), .CLK(clk), .RST(rst), .Q(
        start_reg[101]) );
  DFF \start_reg_reg[102]  ( .D(start_in[101]), .CLK(clk), .RST(rst), .Q(
        start_reg[102]) );
  DFF \start_reg_reg[103]  ( .D(start_in[102]), .CLK(clk), .RST(rst), .Q(
        start_reg[103]) );
  DFF \start_reg_reg[104]  ( .D(start_in[103]), .CLK(clk), .RST(rst), .Q(
        start_reg[104]) );
  DFF \start_reg_reg[105]  ( .D(start_in[104]), .CLK(clk), .RST(rst), .Q(
        start_reg[105]) );
  DFF \start_reg_reg[106]  ( .D(start_in[105]), .CLK(clk), .RST(rst), .Q(
        start_reg[106]) );
  DFF \start_reg_reg[107]  ( .D(start_in[106]), .CLK(clk), .RST(rst), .Q(
        start_reg[107]) );
  DFF \start_reg_reg[108]  ( .D(start_in[107]), .CLK(clk), .RST(rst), .Q(
        start_reg[108]) );
  DFF \start_reg_reg[109]  ( .D(start_in[108]), .CLK(clk), .RST(rst), .Q(
        start_reg[109]) );
  DFF \start_reg_reg[110]  ( .D(start_in[109]), .CLK(clk), .RST(rst), .Q(
        start_reg[110]) );
  DFF \start_reg_reg[111]  ( .D(start_in[110]), .CLK(clk), .RST(rst), .Q(
        start_reg[111]) );
  DFF \start_reg_reg[112]  ( .D(start_in[111]), .CLK(clk), .RST(rst), .Q(
        start_reg[112]) );
  DFF \start_reg_reg[113]  ( .D(start_in[112]), .CLK(clk), .RST(rst), .Q(
        start_reg[113]) );
  DFF \start_reg_reg[114]  ( .D(start_in[113]), .CLK(clk), .RST(rst), .Q(
        start_reg[114]) );
  DFF \start_reg_reg[115]  ( .D(start_in[114]), .CLK(clk), .RST(rst), .Q(
        start_reg[115]) );
  DFF \start_reg_reg[116]  ( .D(start_in[115]), .CLK(clk), .RST(rst), .Q(
        start_reg[116]) );
  DFF \start_reg_reg[117]  ( .D(start_in[116]), .CLK(clk), .RST(rst), .Q(
        start_reg[117]) );
  DFF \start_reg_reg[118]  ( .D(start_in[117]), .CLK(clk), .RST(rst), .Q(
        start_reg[118]) );
  DFF \start_reg_reg[119]  ( .D(start_in[118]), .CLK(clk), .RST(rst), .Q(
        start_reg[119]) );
  DFF \start_reg_reg[120]  ( .D(start_in[119]), .CLK(clk), .RST(rst), .Q(
        start_reg[120]) );
  DFF \start_reg_reg[121]  ( .D(start_in[120]), .CLK(clk), .RST(rst), .Q(
        start_reg[121]) );
  DFF \start_reg_reg[122]  ( .D(start_in[121]), .CLK(clk), .RST(rst), .Q(
        start_reg[122]) );
  DFF \start_reg_reg[123]  ( .D(start_in[122]), .CLK(clk), .RST(rst), .Q(
        start_reg[123]) );
  DFF \start_reg_reg[124]  ( .D(start_in[123]), .CLK(clk), .RST(rst), .Q(
        start_reg[124]) );
  DFF \start_reg_reg[125]  ( .D(start_in[124]), .CLK(clk), .RST(rst), .Q(
        start_reg[125]) );
  DFF \start_reg_reg[126]  ( .D(start_in[125]), .CLK(clk), .RST(rst), .Q(
        start_reg[126]) );
  DFF \start_reg_reg[127]  ( .D(start_in[126]), .CLK(clk), .RST(rst), .Q(
        start_reg[127]) );
  DFF \start_reg_reg[128]  ( .D(start_in[127]), .CLK(clk), .RST(rst), .Q(
        start_reg[128]) );
  DFF \start_reg_reg[129]  ( .D(start_in[128]), .CLK(clk), .RST(rst), .Q(
        start_reg[129]) );
  DFF \start_reg_reg[130]  ( .D(start_in[129]), .CLK(clk), .RST(rst), .Q(
        start_reg[130]) );
  DFF \start_reg_reg[131]  ( .D(start_in[130]), .CLK(clk), .RST(rst), .Q(
        start_reg[131]) );
  DFF \start_reg_reg[132]  ( .D(start_in[131]), .CLK(clk), .RST(rst), .Q(
        start_reg[132]) );
  DFF \start_reg_reg[133]  ( .D(start_in[132]), .CLK(clk), .RST(rst), .Q(
        start_reg[133]) );
  DFF \start_reg_reg[134]  ( .D(start_in[133]), .CLK(clk), .RST(rst), .Q(
        start_reg[134]) );
  DFF \start_reg_reg[135]  ( .D(start_in[134]), .CLK(clk), .RST(rst), .Q(
        start_reg[135]) );
  DFF \start_reg_reg[136]  ( .D(start_in[135]), .CLK(clk), .RST(rst), .Q(
        start_reg[136]) );
  DFF \start_reg_reg[137]  ( .D(start_in[136]), .CLK(clk), .RST(rst), .Q(
        start_reg[137]) );
  DFF \start_reg_reg[138]  ( .D(start_in[137]), .CLK(clk), .RST(rst), .Q(
        start_reg[138]) );
  DFF \start_reg_reg[139]  ( .D(start_in[138]), .CLK(clk), .RST(rst), .Q(
        start_reg[139]) );
  DFF \start_reg_reg[140]  ( .D(start_in[139]), .CLK(clk), .RST(rst), .Q(
        start_reg[140]) );
  DFF \start_reg_reg[141]  ( .D(start_in[140]), .CLK(clk), .RST(rst), .Q(
        start_reg[141]) );
  DFF \start_reg_reg[142]  ( .D(start_in[141]), .CLK(clk), .RST(rst), .Q(
        start_reg[142]) );
  DFF \start_reg_reg[143]  ( .D(start_in[142]), .CLK(clk), .RST(rst), .Q(
        start_reg[143]) );
  DFF \start_reg_reg[144]  ( .D(start_in[143]), .CLK(clk), .RST(rst), .Q(
        start_reg[144]) );
  DFF \start_reg_reg[145]  ( .D(start_in[144]), .CLK(clk), .RST(rst), .Q(
        start_reg[145]) );
  DFF \start_reg_reg[146]  ( .D(start_in[145]), .CLK(clk), .RST(rst), .Q(
        start_reg[146]) );
  DFF \start_reg_reg[147]  ( .D(start_in[146]), .CLK(clk), .RST(rst), .Q(
        start_reg[147]) );
  DFF \start_reg_reg[148]  ( .D(start_in[147]), .CLK(clk), .RST(rst), .Q(
        start_reg[148]) );
  DFF \start_reg_reg[149]  ( .D(start_in[148]), .CLK(clk), .RST(rst), .Q(
        start_reg[149]) );
  DFF \start_reg_reg[150]  ( .D(start_in[149]), .CLK(clk), .RST(rst), .Q(
        start_reg[150]) );
  DFF \start_reg_reg[151]  ( .D(start_in[150]), .CLK(clk), .RST(rst), .Q(
        start_reg[151]) );
  DFF \start_reg_reg[152]  ( .D(start_in[151]), .CLK(clk), .RST(rst), .Q(
        start_reg[152]) );
  DFF \start_reg_reg[153]  ( .D(start_in[152]), .CLK(clk), .RST(rst), .Q(
        start_reg[153]) );
  DFF \start_reg_reg[154]  ( .D(start_in[153]), .CLK(clk), .RST(rst), .Q(
        start_reg[154]) );
  DFF \start_reg_reg[155]  ( .D(start_in[154]), .CLK(clk), .RST(rst), .Q(
        start_reg[155]) );
  DFF \start_reg_reg[156]  ( .D(start_in[155]), .CLK(clk), .RST(rst), .Q(
        start_reg[156]) );
  DFF \start_reg_reg[157]  ( .D(start_in[156]), .CLK(clk), .RST(rst), .Q(
        start_reg[157]) );
  DFF \start_reg_reg[158]  ( .D(start_in[157]), .CLK(clk), .RST(rst), .Q(
        start_reg[158]) );
  DFF \start_reg_reg[159]  ( .D(start_in[158]), .CLK(clk), .RST(rst), .Q(
        start_reg[159]) );
  DFF \start_reg_reg[160]  ( .D(start_in[159]), .CLK(clk), .RST(rst), .Q(
        start_reg[160]) );
  DFF \start_reg_reg[161]  ( .D(start_in[160]), .CLK(clk), .RST(rst), .Q(
        start_reg[161]) );
  DFF \start_reg_reg[162]  ( .D(start_in[161]), .CLK(clk), .RST(rst), .Q(
        start_reg[162]) );
  DFF \start_reg_reg[163]  ( .D(start_in[162]), .CLK(clk), .RST(rst), .Q(
        start_reg[163]) );
  DFF \start_reg_reg[164]  ( .D(start_in[163]), .CLK(clk), .RST(rst), .Q(
        start_reg[164]) );
  DFF \start_reg_reg[165]  ( .D(start_in[164]), .CLK(clk), .RST(rst), .Q(
        start_reg[165]) );
  DFF \start_reg_reg[166]  ( .D(start_in[165]), .CLK(clk), .RST(rst), .Q(
        start_reg[166]) );
  DFF \start_reg_reg[167]  ( .D(start_in[166]), .CLK(clk), .RST(rst), .Q(
        start_reg[167]) );
  DFF \start_reg_reg[168]  ( .D(start_in[167]), .CLK(clk), .RST(rst), .Q(
        start_reg[168]) );
  DFF \start_reg_reg[169]  ( .D(start_in[168]), .CLK(clk), .RST(rst), .Q(
        start_reg[169]) );
  DFF \start_reg_reg[170]  ( .D(start_in[169]), .CLK(clk), .RST(rst), .Q(
        start_reg[170]) );
  DFF \start_reg_reg[171]  ( .D(start_in[170]), .CLK(clk), .RST(rst), .Q(
        start_reg[171]) );
  DFF \start_reg_reg[172]  ( .D(start_in[171]), .CLK(clk), .RST(rst), .Q(
        start_reg[172]) );
  DFF \start_reg_reg[173]  ( .D(start_in[172]), .CLK(clk), .RST(rst), .Q(
        start_reg[173]) );
  DFF \start_reg_reg[174]  ( .D(start_in[173]), .CLK(clk), .RST(rst), .Q(
        start_reg[174]) );
  DFF \start_reg_reg[175]  ( .D(start_in[174]), .CLK(clk), .RST(rst), .Q(
        start_reg[175]) );
  DFF \start_reg_reg[176]  ( .D(start_in[175]), .CLK(clk), .RST(rst), .Q(
        start_reg[176]) );
  DFF \start_reg_reg[177]  ( .D(start_in[176]), .CLK(clk), .RST(rst), .Q(
        start_reg[177]) );
  DFF \start_reg_reg[178]  ( .D(start_in[177]), .CLK(clk), .RST(rst), .Q(
        start_reg[178]) );
  DFF \start_reg_reg[179]  ( .D(start_in[178]), .CLK(clk), .RST(rst), .Q(
        start_reg[179]) );
  DFF \start_reg_reg[180]  ( .D(start_in[179]), .CLK(clk), .RST(rst), .Q(
        start_reg[180]) );
  DFF \start_reg_reg[181]  ( .D(start_in[180]), .CLK(clk), .RST(rst), .Q(
        start_reg[181]) );
  DFF \start_reg_reg[182]  ( .D(start_in[181]), .CLK(clk), .RST(rst), .Q(
        start_reg[182]) );
  DFF \start_reg_reg[183]  ( .D(start_in[182]), .CLK(clk), .RST(rst), .Q(
        start_reg[183]) );
  DFF \start_reg_reg[184]  ( .D(start_in[183]), .CLK(clk), .RST(rst), .Q(
        start_reg[184]) );
  DFF \start_reg_reg[185]  ( .D(start_in[184]), .CLK(clk), .RST(rst), .Q(
        start_reg[185]) );
  DFF \start_reg_reg[186]  ( .D(start_in[185]), .CLK(clk), .RST(rst), .Q(
        start_reg[186]) );
  DFF \start_reg_reg[187]  ( .D(start_in[186]), .CLK(clk), .RST(rst), .Q(
        start_reg[187]) );
  DFF \start_reg_reg[188]  ( .D(start_in[187]), .CLK(clk), .RST(rst), .Q(
        start_reg[188]) );
  DFF \start_reg_reg[189]  ( .D(start_in[188]), .CLK(clk), .RST(rst), .Q(
        start_reg[189]) );
  DFF \start_reg_reg[190]  ( .D(start_in[189]), .CLK(clk), .RST(rst), .Q(
        start_reg[190]) );
  DFF \start_reg_reg[191]  ( .D(start_in[190]), .CLK(clk), .RST(rst), .Q(
        start_reg[191]) );
  DFF \start_reg_reg[192]  ( .D(start_in[191]), .CLK(clk), .RST(rst), .Q(
        start_reg[192]) );
  DFF \start_reg_reg[193]  ( .D(start_in[192]), .CLK(clk), .RST(rst), .Q(
        start_reg[193]) );
  DFF \start_reg_reg[194]  ( .D(start_in[193]), .CLK(clk), .RST(rst), .Q(
        start_reg[194]) );
  DFF \start_reg_reg[195]  ( .D(start_in[194]), .CLK(clk), .RST(rst), .Q(
        start_reg[195]) );
  DFF \start_reg_reg[196]  ( .D(start_in[195]), .CLK(clk), .RST(rst), .Q(
        start_reg[196]) );
  DFF \start_reg_reg[197]  ( .D(start_in[196]), .CLK(clk), .RST(rst), .Q(
        start_reg[197]) );
  DFF \start_reg_reg[198]  ( .D(start_in[197]), .CLK(clk), .RST(rst), .Q(
        start_reg[198]) );
  DFF \start_reg_reg[199]  ( .D(start_in[198]), .CLK(clk), .RST(rst), .Q(
        start_reg[199]) );
  DFF \start_reg_reg[200]  ( .D(start_in[199]), .CLK(clk), .RST(rst), .Q(
        start_reg[200]) );
  DFF \start_reg_reg[201]  ( .D(start_in[200]), .CLK(clk), .RST(rst), .Q(
        start_reg[201]) );
  DFF \start_reg_reg[202]  ( .D(start_in[201]), .CLK(clk), .RST(rst), .Q(
        start_reg[202]) );
  DFF \start_reg_reg[203]  ( .D(start_in[202]), .CLK(clk), .RST(rst), .Q(
        start_reg[203]) );
  DFF \start_reg_reg[204]  ( .D(start_in[203]), .CLK(clk), .RST(rst), .Q(
        start_reg[204]) );
  DFF \start_reg_reg[205]  ( .D(start_in[204]), .CLK(clk), .RST(rst), .Q(
        start_reg[205]) );
  DFF \start_reg_reg[206]  ( .D(start_in[205]), .CLK(clk), .RST(rst), .Q(
        start_reg[206]) );
  DFF \start_reg_reg[207]  ( .D(start_in[206]), .CLK(clk), .RST(rst), .Q(
        start_reg[207]) );
  DFF \start_reg_reg[208]  ( .D(start_in[207]), .CLK(clk), .RST(rst), .Q(
        start_reg[208]) );
  DFF \start_reg_reg[209]  ( .D(start_in[208]), .CLK(clk), .RST(rst), .Q(
        start_reg[209]) );
  DFF \start_reg_reg[210]  ( .D(start_in[209]), .CLK(clk), .RST(rst), .Q(
        start_reg[210]) );
  DFF \start_reg_reg[211]  ( .D(start_in[210]), .CLK(clk), .RST(rst), .Q(
        start_reg[211]) );
  DFF \start_reg_reg[212]  ( .D(start_in[211]), .CLK(clk), .RST(rst), .Q(
        start_reg[212]) );
  DFF \start_reg_reg[213]  ( .D(start_in[212]), .CLK(clk), .RST(rst), .Q(
        start_reg[213]) );
  DFF \start_reg_reg[214]  ( .D(start_in[213]), .CLK(clk), .RST(rst), .Q(
        start_reg[214]) );
  DFF \start_reg_reg[215]  ( .D(start_in[214]), .CLK(clk), .RST(rst), .Q(
        start_reg[215]) );
  DFF \start_reg_reg[216]  ( .D(start_in[215]), .CLK(clk), .RST(rst), .Q(
        start_reg[216]) );
  DFF \start_reg_reg[217]  ( .D(start_in[216]), .CLK(clk), .RST(rst), .Q(
        start_reg[217]) );
  DFF \start_reg_reg[218]  ( .D(start_in[217]), .CLK(clk), .RST(rst), .Q(
        start_reg[218]) );
  DFF \start_reg_reg[219]  ( .D(start_in[218]), .CLK(clk), .RST(rst), .Q(
        start_reg[219]) );
  DFF \start_reg_reg[220]  ( .D(start_in[219]), .CLK(clk), .RST(rst), .Q(
        start_reg[220]) );
  DFF \start_reg_reg[221]  ( .D(start_in[220]), .CLK(clk), .RST(rst), .Q(
        start_reg[221]) );
  DFF \start_reg_reg[222]  ( .D(start_in[221]), .CLK(clk), .RST(rst), .Q(
        start_reg[222]) );
  DFF \start_reg_reg[223]  ( .D(start_in[222]), .CLK(clk), .RST(rst), .Q(
        start_reg[223]) );
  DFF \start_reg_reg[224]  ( .D(start_in[223]), .CLK(clk), .RST(rst), .Q(
        start_reg[224]) );
  DFF \start_reg_reg[225]  ( .D(start_in[224]), .CLK(clk), .RST(rst), .Q(
        start_reg[225]) );
  DFF \start_reg_reg[226]  ( .D(start_in[225]), .CLK(clk), .RST(rst), .Q(
        start_reg[226]) );
  DFF \start_reg_reg[227]  ( .D(start_in[226]), .CLK(clk), .RST(rst), .Q(
        start_reg[227]) );
  DFF \start_reg_reg[228]  ( .D(start_in[227]), .CLK(clk), .RST(rst), .Q(
        start_reg[228]) );
  DFF \start_reg_reg[229]  ( .D(start_in[228]), .CLK(clk), .RST(rst), .Q(
        start_reg[229]) );
  DFF \start_reg_reg[230]  ( .D(start_in[229]), .CLK(clk), .RST(rst), .Q(
        start_reg[230]) );
  DFF \start_reg_reg[231]  ( .D(start_in[230]), .CLK(clk), .RST(rst), .Q(
        start_reg[231]) );
  DFF \start_reg_reg[232]  ( .D(start_in[231]), .CLK(clk), .RST(rst), .Q(
        start_reg[232]) );
  DFF \start_reg_reg[233]  ( .D(start_in[232]), .CLK(clk), .RST(rst), .Q(
        start_reg[233]) );
  DFF \start_reg_reg[234]  ( .D(start_in[233]), .CLK(clk), .RST(rst), .Q(
        start_reg[234]) );
  DFF \start_reg_reg[235]  ( .D(start_in[234]), .CLK(clk), .RST(rst), .Q(
        start_reg[235]) );
  DFF \start_reg_reg[236]  ( .D(start_in[235]), .CLK(clk), .RST(rst), .Q(
        start_reg[236]) );
  DFF \start_reg_reg[237]  ( .D(start_in[236]), .CLK(clk), .RST(rst), .Q(
        start_reg[237]) );
  DFF \start_reg_reg[238]  ( .D(start_in[237]), .CLK(clk), .RST(rst), .Q(
        start_reg[238]) );
  DFF \start_reg_reg[239]  ( .D(start_in[238]), .CLK(clk), .RST(rst), .Q(
        start_reg[239]) );
  DFF \start_reg_reg[240]  ( .D(start_in[239]), .CLK(clk), .RST(rst), .Q(
        start_reg[240]) );
  DFF \start_reg_reg[241]  ( .D(start_in[240]), .CLK(clk), .RST(rst), .Q(
        start_reg[241]) );
  DFF \start_reg_reg[242]  ( .D(start_in[241]), .CLK(clk), .RST(rst), .Q(
        start_reg[242]) );
  DFF \start_reg_reg[243]  ( .D(start_in[242]), .CLK(clk), .RST(rst), .Q(
        start_reg[243]) );
  DFF \start_reg_reg[244]  ( .D(start_in[243]), .CLK(clk), .RST(rst), .Q(
        start_reg[244]) );
  DFF \start_reg_reg[245]  ( .D(start_in[244]), .CLK(clk), .RST(rst), .Q(
        start_reg[245]) );
  DFF \start_reg_reg[246]  ( .D(start_in[245]), .CLK(clk), .RST(rst), .Q(
        start_reg[246]) );
  DFF \start_reg_reg[247]  ( .D(start_in[246]), .CLK(clk), .RST(rst), .Q(
        start_reg[247]) );
  DFF \start_reg_reg[248]  ( .D(start_in[247]), .CLK(clk), .RST(rst), .Q(
        start_reg[248]) );
  DFF \start_reg_reg[249]  ( .D(start_in[248]), .CLK(clk), .RST(rst), .Q(
        start_reg[249]) );
  DFF \start_reg_reg[250]  ( .D(start_in[249]), .CLK(clk), .RST(rst), .Q(
        start_reg[250]) );
  DFF \start_reg_reg[251]  ( .D(start_in[250]), .CLK(clk), .RST(rst), .Q(
        start_reg[251]) );
  DFF \start_reg_reg[252]  ( .D(start_in[251]), .CLK(clk), .RST(rst), .Q(
        start_reg[252]) );
  DFF \start_reg_reg[253]  ( .D(start_in[252]), .CLK(clk), .RST(rst), .Q(
        start_reg[253]) );
  DFF \start_reg_reg[254]  ( .D(start_in[253]), .CLK(clk), .RST(rst), .Q(
        start_reg[254]) );
  DFF \start_reg_reg[255]  ( .D(start_in[254]), .CLK(clk), .RST(rst), .Q(
        start_reg[255]) );
  DFF \start_reg_reg[256]  ( .D(start_in[255]), .CLK(clk), .RST(rst), .Q(
        start_reg[256]) );
  DFF \start_reg_reg[257]  ( .D(start_in[256]), .CLK(clk), .RST(rst), .Q(
        start_reg[257]) );
  DFF \start_reg_reg[258]  ( .D(start_in[257]), .CLK(clk), .RST(rst), .Q(
        start_reg[258]) );
  DFF \start_reg_reg[259]  ( .D(start_in[258]), .CLK(clk), .RST(rst), .Q(
        start_reg[259]) );
  DFF \start_reg_reg[260]  ( .D(start_in[259]), .CLK(clk), .RST(rst), .Q(
        start_reg[260]) );
  DFF \start_reg_reg[261]  ( .D(start_in[260]), .CLK(clk), .RST(rst), .Q(
        start_reg[261]) );
  DFF \start_reg_reg[262]  ( .D(start_in[261]), .CLK(clk), .RST(rst), .Q(
        start_reg[262]) );
  DFF \start_reg_reg[263]  ( .D(start_in[262]), .CLK(clk), .RST(rst), .Q(
        start_reg[263]) );
  DFF \start_reg_reg[264]  ( .D(start_in[263]), .CLK(clk), .RST(rst), .Q(
        start_reg[264]) );
  DFF \start_reg_reg[265]  ( .D(start_in[264]), .CLK(clk), .RST(rst), .Q(
        start_reg[265]) );
  DFF \start_reg_reg[266]  ( .D(start_in[265]), .CLK(clk), .RST(rst), .Q(
        start_reg[266]) );
  DFF \start_reg_reg[267]  ( .D(start_in[266]), .CLK(clk), .RST(rst), .Q(
        start_reg[267]) );
  DFF \start_reg_reg[268]  ( .D(start_in[267]), .CLK(clk), .RST(rst), .Q(
        start_reg[268]) );
  DFF \start_reg_reg[269]  ( .D(start_in[268]), .CLK(clk), .RST(rst), .Q(
        start_reg[269]) );
  DFF \start_reg_reg[270]  ( .D(start_in[269]), .CLK(clk), .RST(rst), .Q(
        start_reg[270]) );
  DFF \start_reg_reg[271]  ( .D(start_in[270]), .CLK(clk), .RST(rst), .Q(
        start_reg[271]) );
  DFF \start_reg_reg[272]  ( .D(start_in[271]), .CLK(clk), .RST(rst), .Q(
        start_reg[272]) );
  DFF \start_reg_reg[273]  ( .D(start_in[272]), .CLK(clk), .RST(rst), .Q(
        start_reg[273]) );
  DFF \start_reg_reg[274]  ( .D(start_in[273]), .CLK(clk), .RST(rst), .Q(
        start_reg[274]) );
  DFF \start_reg_reg[275]  ( .D(start_in[274]), .CLK(clk), .RST(rst), .Q(
        start_reg[275]) );
  DFF \start_reg_reg[276]  ( .D(start_in[275]), .CLK(clk), .RST(rst), .Q(
        start_reg[276]) );
  DFF \start_reg_reg[277]  ( .D(start_in[276]), .CLK(clk), .RST(rst), .Q(
        start_reg[277]) );
  DFF \start_reg_reg[278]  ( .D(start_in[277]), .CLK(clk), .RST(rst), .Q(
        start_reg[278]) );
  DFF \start_reg_reg[279]  ( .D(start_in[278]), .CLK(clk), .RST(rst), .Q(
        start_reg[279]) );
  DFF \start_reg_reg[280]  ( .D(start_in[279]), .CLK(clk), .RST(rst), .Q(
        start_reg[280]) );
  DFF \start_reg_reg[281]  ( .D(start_in[280]), .CLK(clk), .RST(rst), .Q(
        start_reg[281]) );
  DFF \start_reg_reg[282]  ( .D(start_in[281]), .CLK(clk), .RST(rst), .Q(
        start_reg[282]) );
  DFF \start_reg_reg[283]  ( .D(start_in[282]), .CLK(clk), .RST(rst), .Q(
        start_reg[283]) );
  DFF \start_reg_reg[284]  ( .D(start_in[283]), .CLK(clk), .RST(rst), .Q(
        start_reg[284]) );
  DFF \start_reg_reg[285]  ( .D(start_in[284]), .CLK(clk), .RST(rst), .Q(
        start_reg[285]) );
  DFF \start_reg_reg[286]  ( .D(start_in[285]), .CLK(clk), .RST(rst), .Q(
        start_reg[286]) );
  DFF \start_reg_reg[287]  ( .D(start_in[286]), .CLK(clk), .RST(rst), .Q(
        start_reg[287]) );
  DFF \start_reg_reg[288]  ( .D(start_in[287]), .CLK(clk), .RST(rst), .Q(
        start_reg[288]) );
  DFF \start_reg_reg[289]  ( .D(start_in[288]), .CLK(clk), .RST(rst), .Q(
        start_reg[289]) );
  DFF \start_reg_reg[290]  ( .D(start_in[289]), .CLK(clk), .RST(rst), .Q(
        start_reg[290]) );
  DFF \start_reg_reg[291]  ( .D(start_in[290]), .CLK(clk), .RST(rst), .Q(
        start_reg[291]) );
  DFF \start_reg_reg[292]  ( .D(start_in[291]), .CLK(clk), .RST(rst), .Q(
        start_reg[292]) );
  DFF \start_reg_reg[293]  ( .D(start_in[292]), .CLK(clk), .RST(rst), .Q(
        start_reg[293]) );
  DFF \start_reg_reg[294]  ( .D(start_in[293]), .CLK(clk), .RST(rst), .Q(
        start_reg[294]) );
  DFF \start_reg_reg[295]  ( .D(start_in[294]), .CLK(clk), .RST(rst), .Q(
        start_reg[295]) );
  DFF \start_reg_reg[296]  ( .D(start_in[295]), .CLK(clk), .RST(rst), .Q(
        start_reg[296]) );
  DFF \start_reg_reg[297]  ( .D(start_in[296]), .CLK(clk), .RST(rst), .Q(
        start_reg[297]) );
  DFF \start_reg_reg[298]  ( .D(start_in[297]), .CLK(clk), .RST(rst), .Q(
        start_reg[298]) );
  DFF \start_reg_reg[299]  ( .D(start_in[298]), .CLK(clk), .RST(rst), .Q(
        start_reg[299]) );
  DFF \start_reg_reg[300]  ( .D(start_in[299]), .CLK(clk), .RST(rst), .Q(
        start_reg[300]) );
  DFF \start_reg_reg[301]  ( .D(start_in[300]), .CLK(clk), .RST(rst), .Q(
        start_reg[301]) );
  DFF \start_reg_reg[302]  ( .D(start_in[301]), .CLK(clk), .RST(rst), .Q(
        start_reg[302]) );
  DFF \start_reg_reg[303]  ( .D(start_in[302]), .CLK(clk), .RST(rst), .Q(
        start_reg[303]) );
  DFF \start_reg_reg[304]  ( .D(start_in[303]), .CLK(clk), .RST(rst), .Q(
        start_reg[304]) );
  DFF \start_reg_reg[305]  ( .D(start_in[304]), .CLK(clk), .RST(rst), .Q(
        start_reg[305]) );
  DFF \start_reg_reg[306]  ( .D(start_in[305]), .CLK(clk), .RST(rst), .Q(
        start_reg[306]) );
  DFF \start_reg_reg[307]  ( .D(start_in[306]), .CLK(clk), .RST(rst), .Q(
        start_reg[307]) );
  DFF \start_reg_reg[308]  ( .D(start_in[307]), .CLK(clk), .RST(rst), .Q(
        start_reg[308]) );
  DFF \start_reg_reg[309]  ( .D(start_in[308]), .CLK(clk), .RST(rst), .Q(
        start_reg[309]) );
  DFF \start_reg_reg[310]  ( .D(start_in[309]), .CLK(clk), .RST(rst), .Q(
        start_reg[310]) );
  DFF \start_reg_reg[311]  ( .D(start_in[310]), .CLK(clk), .RST(rst), .Q(
        start_reg[311]) );
  DFF \start_reg_reg[312]  ( .D(start_in[311]), .CLK(clk), .RST(rst), .Q(
        start_reg[312]) );
  DFF \start_reg_reg[313]  ( .D(start_in[312]), .CLK(clk), .RST(rst), .Q(
        start_reg[313]) );
  DFF \start_reg_reg[314]  ( .D(start_in[313]), .CLK(clk), .RST(rst), .Q(
        start_reg[314]) );
  DFF \start_reg_reg[315]  ( .D(start_in[314]), .CLK(clk), .RST(rst), .Q(
        start_reg[315]) );
  DFF \start_reg_reg[316]  ( .D(start_in[315]), .CLK(clk), .RST(rst), .Q(
        start_reg[316]) );
  DFF \start_reg_reg[317]  ( .D(start_in[316]), .CLK(clk), .RST(rst), .Q(
        start_reg[317]) );
  DFF \start_reg_reg[318]  ( .D(start_in[317]), .CLK(clk), .RST(rst), .Q(
        start_reg[318]) );
  DFF \start_reg_reg[319]  ( .D(start_in[318]), .CLK(clk), .RST(rst), .Q(
        start_reg[319]) );
  DFF \start_reg_reg[320]  ( .D(start_in[319]), .CLK(clk), .RST(rst), .Q(
        start_reg[320]) );
  DFF \start_reg_reg[321]  ( .D(start_in[320]), .CLK(clk), .RST(rst), .Q(
        start_reg[321]) );
  DFF \start_reg_reg[322]  ( .D(start_in[321]), .CLK(clk), .RST(rst), .Q(
        start_reg[322]) );
  DFF \start_reg_reg[323]  ( .D(start_in[322]), .CLK(clk), .RST(rst), .Q(
        start_reg[323]) );
  DFF \start_reg_reg[324]  ( .D(start_in[323]), .CLK(clk), .RST(rst), .Q(
        start_reg[324]) );
  DFF \start_reg_reg[325]  ( .D(start_in[324]), .CLK(clk), .RST(rst), .Q(
        start_reg[325]) );
  DFF \start_reg_reg[326]  ( .D(start_in[325]), .CLK(clk), .RST(rst), .Q(
        start_reg[326]) );
  DFF \start_reg_reg[327]  ( .D(start_in[326]), .CLK(clk), .RST(rst), .Q(
        start_reg[327]) );
  DFF \start_reg_reg[328]  ( .D(start_in[327]), .CLK(clk), .RST(rst), .Q(
        start_reg[328]) );
  DFF \start_reg_reg[329]  ( .D(start_in[328]), .CLK(clk), .RST(rst), .Q(
        start_reg[329]) );
  DFF \start_reg_reg[330]  ( .D(start_in[329]), .CLK(clk), .RST(rst), .Q(
        start_reg[330]) );
  DFF \start_reg_reg[331]  ( .D(start_in[330]), .CLK(clk), .RST(rst), .Q(
        start_reg[331]) );
  DFF \start_reg_reg[332]  ( .D(start_in[331]), .CLK(clk), .RST(rst), .Q(
        start_reg[332]) );
  DFF \start_reg_reg[333]  ( .D(start_in[332]), .CLK(clk), .RST(rst), .Q(
        start_reg[333]) );
  DFF \start_reg_reg[334]  ( .D(start_in[333]), .CLK(clk), .RST(rst), .Q(
        start_reg[334]) );
  DFF \start_reg_reg[335]  ( .D(start_in[334]), .CLK(clk), .RST(rst), .Q(
        start_reg[335]) );
  DFF \start_reg_reg[336]  ( .D(start_in[335]), .CLK(clk), .RST(rst), .Q(
        start_reg[336]) );
  DFF \start_reg_reg[337]  ( .D(start_in[336]), .CLK(clk), .RST(rst), .Q(
        start_reg[337]) );
  DFF \start_reg_reg[338]  ( .D(start_in[337]), .CLK(clk), .RST(rst), .Q(
        start_reg[338]) );
  DFF \start_reg_reg[339]  ( .D(start_in[338]), .CLK(clk), .RST(rst), .Q(
        start_reg[339]) );
  DFF \start_reg_reg[340]  ( .D(start_in[339]), .CLK(clk), .RST(rst), .Q(
        start_reg[340]) );
  DFF \start_reg_reg[341]  ( .D(start_in[340]), .CLK(clk), .RST(rst), .Q(
        start_reg[341]) );
  DFF \start_reg_reg[342]  ( .D(start_in[341]), .CLK(clk), .RST(rst), .Q(
        start_reg[342]) );
  DFF \start_reg_reg[343]  ( .D(start_in[342]), .CLK(clk), .RST(rst), .Q(
        start_reg[343]) );
  DFF \start_reg_reg[344]  ( .D(start_in[343]), .CLK(clk), .RST(rst), .Q(
        start_reg[344]) );
  DFF \start_reg_reg[345]  ( .D(start_in[344]), .CLK(clk), .RST(rst), .Q(
        start_reg[345]) );
  DFF \start_reg_reg[346]  ( .D(start_in[345]), .CLK(clk), .RST(rst), .Q(
        start_reg[346]) );
  DFF \start_reg_reg[347]  ( .D(start_in[346]), .CLK(clk), .RST(rst), .Q(
        start_reg[347]) );
  DFF \start_reg_reg[348]  ( .D(start_in[347]), .CLK(clk), .RST(rst), .Q(
        start_reg[348]) );
  DFF \start_reg_reg[349]  ( .D(start_in[348]), .CLK(clk), .RST(rst), .Q(
        start_reg[349]) );
  DFF \start_reg_reg[350]  ( .D(start_in[349]), .CLK(clk), .RST(rst), .Q(
        start_reg[350]) );
  DFF \start_reg_reg[351]  ( .D(start_in[350]), .CLK(clk), .RST(rst), .Q(
        start_reg[351]) );
  DFF \start_reg_reg[352]  ( .D(start_in[351]), .CLK(clk), .RST(rst), .Q(
        start_reg[352]) );
  DFF \start_reg_reg[353]  ( .D(start_in[352]), .CLK(clk), .RST(rst), .Q(
        start_reg[353]) );
  DFF \start_reg_reg[354]  ( .D(start_in[353]), .CLK(clk), .RST(rst), .Q(
        start_reg[354]) );
  DFF \start_reg_reg[355]  ( .D(start_in[354]), .CLK(clk), .RST(rst), .Q(
        start_reg[355]) );
  DFF \start_reg_reg[356]  ( .D(start_in[355]), .CLK(clk), .RST(rst), .Q(
        start_reg[356]) );
  DFF \start_reg_reg[357]  ( .D(start_in[356]), .CLK(clk), .RST(rst), .Q(
        start_reg[357]) );
  DFF \start_reg_reg[358]  ( .D(start_in[357]), .CLK(clk), .RST(rst), .Q(
        start_reg[358]) );
  DFF \start_reg_reg[359]  ( .D(start_in[358]), .CLK(clk), .RST(rst), .Q(
        start_reg[359]) );
  DFF \start_reg_reg[360]  ( .D(start_in[359]), .CLK(clk), .RST(rst), .Q(
        start_reg[360]) );
  DFF \start_reg_reg[361]  ( .D(start_in[360]), .CLK(clk), .RST(rst), .Q(
        start_reg[361]) );
  DFF \start_reg_reg[362]  ( .D(start_in[361]), .CLK(clk), .RST(rst), .Q(
        start_reg[362]) );
  DFF \start_reg_reg[363]  ( .D(start_in[362]), .CLK(clk), .RST(rst), .Q(
        start_reg[363]) );
  DFF \start_reg_reg[364]  ( .D(start_in[363]), .CLK(clk), .RST(rst), .Q(
        start_reg[364]) );
  DFF \start_reg_reg[365]  ( .D(start_in[364]), .CLK(clk), .RST(rst), .Q(
        start_reg[365]) );
  DFF \start_reg_reg[366]  ( .D(start_in[365]), .CLK(clk), .RST(rst), .Q(
        start_reg[366]) );
  DFF \start_reg_reg[367]  ( .D(start_in[366]), .CLK(clk), .RST(rst), .Q(
        start_reg[367]) );
  DFF \start_reg_reg[368]  ( .D(start_in[367]), .CLK(clk), .RST(rst), .Q(
        start_reg[368]) );
  DFF \start_reg_reg[369]  ( .D(start_in[368]), .CLK(clk), .RST(rst), .Q(
        start_reg[369]) );
  DFF \start_reg_reg[370]  ( .D(start_in[369]), .CLK(clk), .RST(rst), .Q(
        start_reg[370]) );
  DFF \start_reg_reg[371]  ( .D(start_in[370]), .CLK(clk), .RST(rst), .Q(
        start_reg[371]) );
  DFF \start_reg_reg[372]  ( .D(start_in[371]), .CLK(clk), .RST(rst), .Q(
        start_reg[372]) );
  DFF \start_reg_reg[373]  ( .D(start_in[372]), .CLK(clk), .RST(rst), .Q(
        start_reg[373]) );
  DFF \start_reg_reg[374]  ( .D(start_in[373]), .CLK(clk), .RST(rst), .Q(
        start_reg[374]) );
  DFF \start_reg_reg[375]  ( .D(start_in[374]), .CLK(clk), .RST(rst), .Q(
        start_reg[375]) );
  DFF \start_reg_reg[376]  ( .D(start_in[375]), .CLK(clk), .RST(rst), .Q(
        start_reg[376]) );
  DFF \start_reg_reg[377]  ( .D(start_in[376]), .CLK(clk), .RST(rst), .Q(
        start_reg[377]) );
  DFF \start_reg_reg[378]  ( .D(start_in[377]), .CLK(clk), .RST(rst), .Q(
        start_reg[378]) );
  DFF \start_reg_reg[379]  ( .D(start_in[378]), .CLK(clk), .RST(rst), .Q(
        start_reg[379]) );
  DFF \start_reg_reg[380]  ( .D(start_in[379]), .CLK(clk), .RST(rst), .Q(
        start_reg[380]) );
  DFF \start_reg_reg[381]  ( .D(start_in[380]), .CLK(clk), .RST(rst), .Q(
        start_reg[381]) );
  DFF \start_reg_reg[382]  ( .D(start_in[381]), .CLK(clk), .RST(rst), .Q(
        start_reg[382]) );
  DFF \start_reg_reg[383]  ( .D(start_in[382]), .CLK(clk), .RST(rst), .Q(
        start_reg[383]) );
  DFF \start_reg_reg[384]  ( .D(start_in[383]), .CLK(clk), .RST(rst), .Q(
        start_reg[384]) );
  DFF \start_reg_reg[385]  ( .D(start_in[384]), .CLK(clk), .RST(rst), .Q(
        start_reg[385]) );
  DFF \start_reg_reg[386]  ( .D(start_in[385]), .CLK(clk), .RST(rst), .Q(
        start_reg[386]) );
  DFF \start_reg_reg[387]  ( .D(start_in[386]), .CLK(clk), .RST(rst), .Q(
        start_reg[387]) );
  DFF \start_reg_reg[388]  ( .D(start_in[387]), .CLK(clk), .RST(rst), .Q(
        start_reg[388]) );
  DFF \start_reg_reg[389]  ( .D(start_in[388]), .CLK(clk), .RST(rst), .Q(
        start_reg[389]) );
  DFF \start_reg_reg[390]  ( .D(start_in[389]), .CLK(clk), .RST(rst), .Q(
        start_reg[390]) );
  DFF \start_reg_reg[391]  ( .D(start_in[390]), .CLK(clk), .RST(rst), .Q(
        start_reg[391]) );
  DFF \start_reg_reg[392]  ( .D(start_in[391]), .CLK(clk), .RST(rst), .Q(
        start_reg[392]) );
  DFF \start_reg_reg[393]  ( .D(start_in[392]), .CLK(clk), .RST(rst), .Q(
        start_reg[393]) );
  DFF \start_reg_reg[394]  ( .D(start_in[393]), .CLK(clk), .RST(rst), .Q(
        start_reg[394]) );
  DFF \start_reg_reg[395]  ( .D(start_in[394]), .CLK(clk), .RST(rst), .Q(
        start_reg[395]) );
  DFF \start_reg_reg[396]  ( .D(start_in[395]), .CLK(clk), .RST(rst), .Q(
        start_reg[396]) );
  DFF \start_reg_reg[397]  ( .D(start_in[396]), .CLK(clk), .RST(rst), .Q(
        start_reg[397]) );
  DFF \start_reg_reg[398]  ( .D(start_in[397]), .CLK(clk), .RST(rst), .Q(
        start_reg[398]) );
  DFF \start_reg_reg[399]  ( .D(start_in[398]), .CLK(clk), .RST(rst), .Q(
        start_reg[399]) );
  DFF \start_reg_reg[400]  ( .D(start_in[399]), .CLK(clk), .RST(rst), .Q(
        start_reg[400]) );
  DFF \start_reg_reg[401]  ( .D(start_in[400]), .CLK(clk), .RST(rst), .Q(
        start_reg[401]) );
  DFF \start_reg_reg[402]  ( .D(start_in[401]), .CLK(clk), .RST(rst), .Q(
        start_reg[402]) );
  DFF \start_reg_reg[403]  ( .D(start_in[402]), .CLK(clk), .RST(rst), .Q(
        start_reg[403]) );
  DFF \start_reg_reg[404]  ( .D(start_in[403]), .CLK(clk), .RST(rst), .Q(
        start_reg[404]) );
  DFF \start_reg_reg[405]  ( .D(start_in[404]), .CLK(clk), .RST(rst), .Q(
        start_reg[405]) );
  DFF \start_reg_reg[406]  ( .D(start_in[405]), .CLK(clk), .RST(rst), .Q(
        start_reg[406]) );
  DFF \start_reg_reg[407]  ( .D(start_in[406]), .CLK(clk), .RST(rst), .Q(
        start_reg[407]) );
  DFF \start_reg_reg[408]  ( .D(start_in[407]), .CLK(clk), .RST(rst), .Q(
        start_reg[408]) );
  DFF \start_reg_reg[409]  ( .D(start_in[408]), .CLK(clk), .RST(rst), .Q(
        start_reg[409]) );
  DFF \start_reg_reg[410]  ( .D(start_in[409]), .CLK(clk), .RST(rst), .Q(
        start_reg[410]) );
  DFF \start_reg_reg[411]  ( .D(start_in[410]), .CLK(clk), .RST(rst), .Q(
        start_reg[411]) );
  DFF \start_reg_reg[412]  ( .D(start_in[411]), .CLK(clk), .RST(rst), .Q(
        start_reg[412]) );
  DFF \start_reg_reg[413]  ( .D(start_in[412]), .CLK(clk), .RST(rst), .Q(
        start_reg[413]) );
  DFF \start_reg_reg[414]  ( .D(start_in[413]), .CLK(clk), .RST(rst), .Q(
        start_reg[414]) );
  DFF \start_reg_reg[415]  ( .D(start_in[414]), .CLK(clk), .RST(rst), .Q(
        start_reg[415]) );
  DFF \start_reg_reg[416]  ( .D(start_in[415]), .CLK(clk), .RST(rst), .Q(
        start_reg[416]) );
  DFF \start_reg_reg[417]  ( .D(start_in[416]), .CLK(clk), .RST(rst), .Q(
        start_reg[417]) );
  DFF \start_reg_reg[418]  ( .D(start_in[417]), .CLK(clk), .RST(rst), .Q(
        start_reg[418]) );
  DFF \start_reg_reg[419]  ( .D(start_in[418]), .CLK(clk), .RST(rst), .Q(
        start_reg[419]) );
  DFF \start_reg_reg[420]  ( .D(start_in[419]), .CLK(clk), .RST(rst), .Q(
        start_reg[420]) );
  DFF \start_reg_reg[421]  ( .D(start_in[420]), .CLK(clk), .RST(rst), .Q(
        start_reg[421]) );
  DFF \start_reg_reg[422]  ( .D(start_in[421]), .CLK(clk), .RST(rst), .Q(
        start_reg[422]) );
  DFF \start_reg_reg[423]  ( .D(start_in[422]), .CLK(clk), .RST(rst), .Q(
        start_reg[423]) );
  DFF \start_reg_reg[424]  ( .D(start_in[423]), .CLK(clk), .RST(rst), .Q(
        start_reg[424]) );
  DFF \start_reg_reg[425]  ( .D(start_in[424]), .CLK(clk), .RST(rst), .Q(
        start_reg[425]) );
  DFF \start_reg_reg[426]  ( .D(start_in[425]), .CLK(clk), .RST(rst), .Q(
        start_reg[426]) );
  DFF \start_reg_reg[427]  ( .D(start_in[426]), .CLK(clk), .RST(rst), .Q(
        start_reg[427]) );
  DFF \start_reg_reg[428]  ( .D(start_in[427]), .CLK(clk), .RST(rst), .Q(
        start_reg[428]) );
  DFF \start_reg_reg[429]  ( .D(start_in[428]), .CLK(clk), .RST(rst), .Q(
        start_reg[429]) );
  DFF \start_reg_reg[430]  ( .D(start_in[429]), .CLK(clk), .RST(rst), .Q(
        start_reg[430]) );
  DFF \start_reg_reg[431]  ( .D(start_in[430]), .CLK(clk), .RST(rst), .Q(
        start_reg[431]) );
  DFF \start_reg_reg[432]  ( .D(start_in[431]), .CLK(clk), .RST(rst), .Q(
        start_reg[432]) );
  DFF \start_reg_reg[433]  ( .D(start_in[432]), .CLK(clk), .RST(rst), .Q(
        start_reg[433]) );
  DFF \start_reg_reg[434]  ( .D(start_in[433]), .CLK(clk), .RST(rst), .Q(
        start_reg[434]) );
  DFF \start_reg_reg[435]  ( .D(start_in[434]), .CLK(clk), .RST(rst), .Q(
        start_reg[435]) );
  DFF \start_reg_reg[436]  ( .D(start_in[435]), .CLK(clk), .RST(rst), .Q(
        start_reg[436]) );
  DFF \start_reg_reg[437]  ( .D(start_in[436]), .CLK(clk), .RST(rst), .Q(
        start_reg[437]) );
  DFF \start_reg_reg[438]  ( .D(start_in[437]), .CLK(clk), .RST(rst), .Q(
        start_reg[438]) );
  DFF \start_reg_reg[439]  ( .D(start_in[438]), .CLK(clk), .RST(rst), .Q(
        start_reg[439]) );
  DFF \start_reg_reg[440]  ( .D(start_in[439]), .CLK(clk), .RST(rst), .Q(
        start_reg[440]) );
  DFF \start_reg_reg[441]  ( .D(start_in[440]), .CLK(clk), .RST(rst), .Q(
        start_reg[441]) );
  DFF \start_reg_reg[442]  ( .D(start_in[441]), .CLK(clk), .RST(rst), .Q(
        start_reg[442]) );
  DFF \start_reg_reg[443]  ( .D(start_in[442]), .CLK(clk), .RST(rst), .Q(
        start_reg[443]) );
  DFF \start_reg_reg[444]  ( .D(start_in[443]), .CLK(clk), .RST(rst), .Q(
        start_reg[444]) );
  DFF \start_reg_reg[445]  ( .D(start_in[444]), .CLK(clk), .RST(rst), .Q(
        start_reg[445]) );
  DFF \start_reg_reg[446]  ( .D(start_in[445]), .CLK(clk), .RST(rst), .Q(
        start_reg[446]) );
  DFF \start_reg_reg[447]  ( .D(start_in[446]), .CLK(clk), .RST(rst), .Q(
        start_reg[447]) );
  DFF \start_reg_reg[448]  ( .D(start_in[447]), .CLK(clk), .RST(rst), .Q(
        start_reg[448]) );
  DFF \start_reg_reg[449]  ( .D(start_in[448]), .CLK(clk), .RST(rst), .Q(
        start_reg[449]) );
  DFF \start_reg_reg[450]  ( .D(start_in[449]), .CLK(clk), .RST(rst), .Q(
        start_reg[450]) );
  DFF \start_reg_reg[451]  ( .D(start_in[450]), .CLK(clk), .RST(rst), .Q(
        start_reg[451]) );
  DFF \start_reg_reg[452]  ( .D(start_in[451]), .CLK(clk), .RST(rst), .Q(
        start_reg[452]) );
  DFF \start_reg_reg[453]  ( .D(start_in[452]), .CLK(clk), .RST(rst), .Q(
        start_reg[453]) );
  DFF \start_reg_reg[454]  ( .D(start_in[453]), .CLK(clk), .RST(rst), .Q(
        start_reg[454]) );
  DFF \start_reg_reg[455]  ( .D(start_in[454]), .CLK(clk), .RST(rst), .Q(
        start_reg[455]) );
  DFF \start_reg_reg[456]  ( .D(start_in[455]), .CLK(clk), .RST(rst), .Q(
        start_reg[456]) );
  DFF \start_reg_reg[457]  ( .D(start_in[456]), .CLK(clk), .RST(rst), .Q(
        start_reg[457]) );
  DFF \start_reg_reg[458]  ( .D(start_in[457]), .CLK(clk), .RST(rst), .Q(
        start_reg[458]) );
  DFF \start_reg_reg[459]  ( .D(start_in[458]), .CLK(clk), .RST(rst), .Q(
        start_reg[459]) );
  DFF \start_reg_reg[460]  ( .D(start_in[459]), .CLK(clk), .RST(rst), .Q(
        start_reg[460]) );
  DFF \start_reg_reg[461]  ( .D(start_in[460]), .CLK(clk), .RST(rst), .Q(
        start_reg[461]) );
  DFF \start_reg_reg[462]  ( .D(start_in[461]), .CLK(clk), .RST(rst), .Q(
        start_reg[462]) );
  DFF \start_reg_reg[463]  ( .D(start_in[462]), .CLK(clk), .RST(rst), .Q(
        start_reg[463]) );
  DFF \start_reg_reg[464]  ( .D(start_in[463]), .CLK(clk), .RST(rst), .Q(
        start_reg[464]) );
  DFF \start_reg_reg[465]  ( .D(start_in[464]), .CLK(clk), .RST(rst), .Q(
        start_reg[465]) );
  DFF \start_reg_reg[466]  ( .D(start_in[465]), .CLK(clk), .RST(rst), .Q(
        start_reg[466]) );
  DFF \start_reg_reg[467]  ( .D(start_in[466]), .CLK(clk), .RST(rst), .Q(
        start_reg[467]) );
  DFF \start_reg_reg[468]  ( .D(start_in[467]), .CLK(clk), .RST(rst), .Q(
        start_reg[468]) );
  DFF \start_reg_reg[469]  ( .D(start_in[468]), .CLK(clk), .RST(rst), .Q(
        start_reg[469]) );
  DFF \start_reg_reg[470]  ( .D(start_in[469]), .CLK(clk), .RST(rst), .Q(
        start_reg[470]) );
  DFF \start_reg_reg[471]  ( .D(start_in[470]), .CLK(clk), .RST(rst), .Q(
        start_reg[471]) );
  DFF \start_reg_reg[472]  ( .D(start_in[471]), .CLK(clk), .RST(rst), .Q(
        start_reg[472]) );
  DFF \start_reg_reg[473]  ( .D(start_in[472]), .CLK(clk), .RST(rst), .Q(
        start_reg[473]) );
  DFF \start_reg_reg[474]  ( .D(start_in[473]), .CLK(clk), .RST(rst), .Q(
        start_reg[474]) );
  DFF \start_reg_reg[475]  ( .D(start_in[474]), .CLK(clk), .RST(rst), .Q(
        start_reg[475]) );
  DFF \start_reg_reg[476]  ( .D(start_in[475]), .CLK(clk), .RST(rst), .Q(
        start_reg[476]) );
  DFF \start_reg_reg[477]  ( .D(start_in[476]), .CLK(clk), .RST(rst), .Q(
        start_reg[477]) );
  DFF \start_reg_reg[478]  ( .D(start_in[477]), .CLK(clk), .RST(rst), .Q(
        start_reg[478]) );
  DFF \start_reg_reg[479]  ( .D(start_in[478]), .CLK(clk), .RST(rst), .Q(
        start_reg[479]) );
  DFF \start_reg_reg[480]  ( .D(start_in[479]), .CLK(clk), .RST(rst), .Q(
        start_reg[480]) );
  DFF \start_reg_reg[481]  ( .D(start_in[480]), .CLK(clk), .RST(rst), .Q(
        start_reg[481]) );
  DFF \start_reg_reg[482]  ( .D(start_in[481]), .CLK(clk), .RST(rst), .Q(
        start_reg[482]) );
  DFF \start_reg_reg[483]  ( .D(start_in[482]), .CLK(clk), .RST(rst), .Q(
        start_reg[483]) );
  DFF \start_reg_reg[484]  ( .D(start_in[483]), .CLK(clk), .RST(rst), .Q(
        start_reg[484]) );
  DFF \start_reg_reg[485]  ( .D(start_in[484]), .CLK(clk), .RST(rst), .Q(
        start_reg[485]) );
  DFF \start_reg_reg[486]  ( .D(start_in[485]), .CLK(clk), .RST(rst), .Q(
        start_reg[486]) );
  DFF \start_reg_reg[487]  ( .D(start_in[486]), .CLK(clk), .RST(rst), .Q(
        start_reg[487]) );
  DFF \start_reg_reg[488]  ( .D(start_in[487]), .CLK(clk), .RST(rst), .Q(
        start_reg[488]) );
  DFF \start_reg_reg[489]  ( .D(start_in[488]), .CLK(clk), .RST(rst), .Q(
        start_reg[489]) );
  DFF \start_reg_reg[490]  ( .D(start_in[489]), .CLK(clk), .RST(rst), .Q(
        start_reg[490]) );
  DFF \start_reg_reg[491]  ( .D(start_in[490]), .CLK(clk), .RST(rst), .Q(
        start_reg[491]) );
  DFF \start_reg_reg[492]  ( .D(start_in[491]), .CLK(clk), .RST(rst), .Q(
        start_reg[492]) );
  DFF \start_reg_reg[493]  ( .D(start_in[492]), .CLK(clk), .RST(rst), .Q(
        start_reg[493]) );
  DFF \start_reg_reg[494]  ( .D(start_in[493]), .CLK(clk), .RST(rst), .Q(
        start_reg[494]) );
  DFF \start_reg_reg[495]  ( .D(start_in[494]), .CLK(clk), .RST(rst), .Q(
        start_reg[495]) );
  DFF \start_reg_reg[496]  ( .D(start_in[495]), .CLK(clk), .RST(rst), .Q(
        start_reg[496]) );
  DFF \start_reg_reg[497]  ( .D(start_in[496]), .CLK(clk), .RST(rst), .Q(
        start_reg[497]) );
  DFF \start_reg_reg[498]  ( .D(start_in[497]), .CLK(clk), .RST(rst), .Q(
        start_reg[498]) );
  DFF \start_reg_reg[499]  ( .D(start_in[498]), .CLK(clk), .RST(rst), .Q(
        start_reg[499]) );
  DFF \start_reg_reg[500]  ( .D(start_in[499]), .CLK(clk), .RST(rst), .Q(
        start_reg[500]) );
  DFF \start_reg_reg[501]  ( .D(start_in[500]), .CLK(clk), .RST(rst), .Q(
        start_reg[501]) );
  DFF \start_reg_reg[502]  ( .D(start_in[501]), .CLK(clk), .RST(rst), .Q(
        start_reg[502]) );
  DFF \start_reg_reg[503]  ( .D(start_in[502]), .CLK(clk), .RST(rst), .Q(
        start_reg[503]) );
  DFF \start_reg_reg[504]  ( .D(start_in[503]), .CLK(clk), .RST(rst), .Q(
        start_reg[504]) );
  DFF \start_reg_reg[505]  ( .D(start_in[504]), .CLK(clk), .RST(rst), .Q(
        start_reg[505]) );
  DFF \start_reg_reg[506]  ( .D(start_in[505]), .CLK(clk), .RST(rst), .Q(
        start_reg[506]) );
  DFF \start_reg_reg[507]  ( .D(start_in[506]), .CLK(clk), .RST(rst), .Q(
        start_reg[507]) );
  DFF \start_reg_reg[508]  ( .D(start_in[507]), .CLK(clk), .RST(rst), .Q(
        start_reg[508]) );
  DFF \start_reg_reg[509]  ( .D(start_in[508]), .CLK(clk), .RST(rst), .Q(
        start_reg[509]) );
  DFF \start_reg_reg[510]  ( .D(start_in[509]), .CLK(clk), .RST(rst), .Q(
        start_reg[510]) );
  DFF \start_reg_reg[511]  ( .D(start_in[510]), .CLK(clk), .RST(rst), .Q(
        start_reg[511]) );
  DFF mul_pow_reg ( .D(n7699), .CLK(clk), .RST(rst), .Q(mul_pow) );
  DFF \ereg_reg[0]  ( .D(n7698), .CLK(clk), .RST(rst), .Q(ereg[0]) );
  DFF \ereg_reg[1]  ( .D(n7697), .CLK(clk), .RST(rst), .Q(ereg[1]) );
  DFF \ereg_reg[2]  ( .D(n7696), .CLK(clk), .RST(rst), .Q(ereg[2]) );
  DFF \ereg_reg[3]  ( .D(n7695), .CLK(clk), .RST(rst), .Q(ereg[3]) );
  DFF \ereg_reg[4]  ( .D(n7694), .CLK(clk), .RST(rst), .Q(ereg[4]) );
  DFF \ereg_reg[5]  ( .D(n7693), .CLK(clk), .RST(rst), .Q(ereg[5]) );
  DFF \ereg_reg[6]  ( .D(n7692), .CLK(clk), .RST(rst), .Q(ereg[6]) );
  DFF \ereg_reg[7]  ( .D(n7691), .CLK(clk), .RST(rst), .Q(ereg[7]) );
  DFF \ereg_reg[8]  ( .D(n7690), .CLK(clk), .RST(rst), .Q(ereg[8]) );
  DFF \ereg_reg[9]  ( .D(n7689), .CLK(clk), .RST(rst), .Q(ereg[9]) );
  DFF \ereg_reg[10]  ( .D(n7688), .CLK(clk), .RST(rst), .Q(ereg[10]) );
  DFF \ereg_reg[11]  ( .D(n7687), .CLK(clk), .RST(rst), .Q(ereg[11]) );
  DFF \ereg_reg[12]  ( .D(n7686), .CLK(clk), .RST(rst), .Q(ereg[12]) );
  DFF \ereg_reg[13]  ( .D(n7685), .CLK(clk), .RST(rst), .Q(ereg[13]) );
  DFF \ereg_reg[14]  ( .D(n7684), .CLK(clk), .RST(rst), .Q(ereg[14]) );
  DFF \ereg_reg[15]  ( .D(n7683), .CLK(clk), .RST(rst), .Q(ereg[15]) );
  DFF \ereg_reg[16]  ( .D(n7682), .CLK(clk), .RST(rst), .Q(ereg[16]) );
  DFF \ereg_reg[17]  ( .D(n7681), .CLK(clk), .RST(rst), .Q(ereg[17]) );
  DFF \ereg_reg[18]  ( .D(n7680), .CLK(clk), .RST(rst), .Q(ereg[18]) );
  DFF \ereg_reg[19]  ( .D(n7679), .CLK(clk), .RST(rst), .Q(ereg[19]) );
  DFF \ereg_reg[20]  ( .D(n7678), .CLK(clk), .RST(rst), .Q(ereg[20]) );
  DFF \ereg_reg[21]  ( .D(n7677), .CLK(clk), .RST(rst), .Q(ereg[21]) );
  DFF \ereg_reg[22]  ( .D(n7676), .CLK(clk), .RST(rst), .Q(ereg[22]) );
  DFF \ereg_reg[23]  ( .D(n7675), .CLK(clk), .RST(rst), .Q(ereg[23]) );
  DFF \ereg_reg[24]  ( .D(n7674), .CLK(clk), .RST(rst), .Q(ereg[24]) );
  DFF \ereg_reg[25]  ( .D(n7673), .CLK(clk), .RST(rst), .Q(ereg[25]) );
  DFF \ereg_reg[26]  ( .D(n7672), .CLK(clk), .RST(rst), .Q(ereg[26]) );
  DFF \ereg_reg[27]  ( .D(n7671), .CLK(clk), .RST(rst), .Q(ereg[27]) );
  DFF \ereg_reg[28]  ( .D(n7670), .CLK(clk), .RST(rst), .Q(ereg[28]) );
  DFF \ereg_reg[29]  ( .D(n7669), .CLK(clk), .RST(rst), .Q(ereg[29]) );
  DFF \ereg_reg[30]  ( .D(n7668), .CLK(clk), .RST(rst), .Q(ereg[30]) );
  DFF \ereg_reg[31]  ( .D(n7667), .CLK(clk), .RST(rst), .Q(ereg[31]) );
  DFF \ereg_reg[32]  ( .D(n7666), .CLK(clk), .RST(rst), .Q(ereg[32]) );
  DFF \ereg_reg[33]  ( .D(n7665), .CLK(clk), .RST(rst), .Q(ereg[33]) );
  DFF \ereg_reg[34]  ( .D(n7664), .CLK(clk), .RST(rst), .Q(ereg[34]) );
  DFF \ereg_reg[35]  ( .D(n7663), .CLK(clk), .RST(rst), .Q(ereg[35]) );
  DFF \ereg_reg[36]  ( .D(n7662), .CLK(clk), .RST(rst), .Q(ereg[36]) );
  DFF \ereg_reg[37]  ( .D(n7661), .CLK(clk), .RST(rst), .Q(ereg[37]) );
  DFF \ereg_reg[38]  ( .D(n7660), .CLK(clk), .RST(rst), .Q(ereg[38]) );
  DFF \ereg_reg[39]  ( .D(n7659), .CLK(clk), .RST(rst), .Q(ereg[39]) );
  DFF \ereg_reg[40]  ( .D(n7658), .CLK(clk), .RST(rst), .Q(ereg[40]) );
  DFF \ereg_reg[41]  ( .D(n7657), .CLK(clk), .RST(rst), .Q(ereg[41]) );
  DFF \ereg_reg[42]  ( .D(n7656), .CLK(clk), .RST(rst), .Q(ereg[42]) );
  DFF \ereg_reg[43]  ( .D(n7655), .CLK(clk), .RST(rst), .Q(ereg[43]) );
  DFF \ereg_reg[44]  ( .D(n7654), .CLK(clk), .RST(rst), .Q(ereg[44]) );
  DFF \ereg_reg[45]  ( .D(n7653), .CLK(clk), .RST(rst), .Q(ereg[45]) );
  DFF \ereg_reg[46]  ( .D(n7652), .CLK(clk), .RST(rst), .Q(ereg[46]) );
  DFF \ereg_reg[47]  ( .D(n7651), .CLK(clk), .RST(rst), .Q(ereg[47]) );
  DFF \ereg_reg[48]  ( .D(n7650), .CLK(clk), .RST(rst), .Q(ereg[48]) );
  DFF \ereg_reg[49]  ( .D(n7649), .CLK(clk), .RST(rst), .Q(ereg[49]) );
  DFF \ereg_reg[50]  ( .D(n7648), .CLK(clk), .RST(rst), .Q(ereg[50]) );
  DFF \ereg_reg[51]  ( .D(n7647), .CLK(clk), .RST(rst), .Q(ereg[51]) );
  DFF \ereg_reg[52]  ( .D(n7646), .CLK(clk), .RST(rst), .Q(ereg[52]) );
  DFF \ereg_reg[53]  ( .D(n7645), .CLK(clk), .RST(rst), .Q(ereg[53]) );
  DFF \ereg_reg[54]  ( .D(n7644), .CLK(clk), .RST(rst), .Q(ereg[54]) );
  DFF \ereg_reg[55]  ( .D(n7643), .CLK(clk), .RST(rst), .Q(ereg[55]) );
  DFF \ereg_reg[56]  ( .D(n7642), .CLK(clk), .RST(rst), .Q(ereg[56]) );
  DFF \ereg_reg[57]  ( .D(n7641), .CLK(clk), .RST(rst), .Q(ereg[57]) );
  DFF \ereg_reg[58]  ( .D(n7640), .CLK(clk), .RST(rst), .Q(ereg[58]) );
  DFF \ereg_reg[59]  ( .D(n7639), .CLK(clk), .RST(rst), .Q(ereg[59]) );
  DFF \ereg_reg[60]  ( .D(n7638), .CLK(clk), .RST(rst), .Q(ereg[60]) );
  DFF \ereg_reg[61]  ( .D(n7637), .CLK(clk), .RST(rst), .Q(ereg[61]) );
  DFF \ereg_reg[62]  ( .D(n7636), .CLK(clk), .RST(rst), .Q(ereg[62]) );
  DFF \ereg_reg[63]  ( .D(n7635), .CLK(clk), .RST(rst), .Q(ereg[63]) );
  DFF \ereg_reg[64]  ( .D(n7634), .CLK(clk), .RST(rst), .Q(ereg[64]) );
  DFF \ereg_reg[65]  ( .D(n7633), .CLK(clk), .RST(rst), .Q(ereg[65]) );
  DFF \ereg_reg[66]  ( .D(n7632), .CLK(clk), .RST(rst), .Q(ereg[66]) );
  DFF \ereg_reg[67]  ( .D(n7631), .CLK(clk), .RST(rst), .Q(ereg[67]) );
  DFF \ereg_reg[68]  ( .D(n7630), .CLK(clk), .RST(rst), .Q(ereg[68]) );
  DFF \ereg_reg[69]  ( .D(n7629), .CLK(clk), .RST(rst), .Q(ereg[69]) );
  DFF \ereg_reg[70]  ( .D(n7628), .CLK(clk), .RST(rst), .Q(ereg[70]) );
  DFF \ereg_reg[71]  ( .D(n7627), .CLK(clk), .RST(rst), .Q(ereg[71]) );
  DFF \ereg_reg[72]  ( .D(n7626), .CLK(clk), .RST(rst), .Q(ereg[72]) );
  DFF \ereg_reg[73]  ( .D(n7625), .CLK(clk), .RST(rst), .Q(ereg[73]) );
  DFF \ereg_reg[74]  ( .D(n7624), .CLK(clk), .RST(rst), .Q(ereg[74]) );
  DFF \ereg_reg[75]  ( .D(n7623), .CLK(clk), .RST(rst), .Q(ereg[75]) );
  DFF \ereg_reg[76]  ( .D(n7622), .CLK(clk), .RST(rst), .Q(ereg[76]) );
  DFF \ereg_reg[77]  ( .D(n7621), .CLK(clk), .RST(rst), .Q(ereg[77]) );
  DFF \ereg_reg[78]  ( .D(n7620), .CLK(clk), .RST(rst), .Q(ereg[78]) );
  DFF \ereg_reg[79]  ( .D(n7619), .CLK(clk), .RST(rst), .Q(ereg[79]) );
  DFF \ereg_reg[80]  ( .D(n7618), .CLK(clk), .RST(rst), .Q(ereg[80]) );
  DFF \ereg_reg[81]  ( .D(n7617), .CLK(clk), .RST(rst), .Q(ereg[81]) );
  DFF \ereg_reg[82]  ( .D(n7616), .CLK(clk), .RST(rst), .Q(ereg[82]) );
  DFF \ereg_reg[83]  ( .D(n7615), .CLK(clk), .RST(rst), .Q(ereg[83]) );
  DFF \ereg_reg[84]  ( .D(n7614), .CLK(clk), .RST(rst), .Q(ereg[84]) );
  DFF \ereg_reg[85]  ( .D(n7613), .CLK(clk), .RST(rst), .Q(ereg[85]) );
  DFF \ereg_reg[86]  ( .D(n7612), .CLK(clk), .RST(rst), .Q(ereg[86]) );
  DFF \ereg_reg[87]  ( .D(n7611), .CLK(clk), .RST(rst), .Q(ereg[87]) );
  DFF \ereg_reg[88]  ( .D(n7610), .CLK(clk), .RST(rst), .Q(ereg[88]) );
  DFF \ereg_reg[89]  ( .D(n7609), .CLK(clk), .RST(rst), .Q(ereg[89]) );
  DFF \ereg_reg[90]  ( .D(n7608), .CLK(clk), .RST(rst), .Q(ereg[90]) );
  DFF \ereg_reg[91]  ( .D(n7607), .CLK(clk), .RST(rst), .Q(ereg[91]) );
  DFF \ereg_reg[92]  ( .D(n7606), .CLK(clk), .RST(rst), .Q(ereg[92]) );
  DFF \ereg_reg[93]  ( .D(n7605), .CLK(clk), .RST(rst), .Q(ereg[93]) );
  DFF \ereg_reg[94]  ( .D(n7604), .CLK(clk), .RST(rst), .Q(ereg[94]) );
  DFF \ereg_reg[95]  ( .D(n7603), .CLK(clk), .RST(rst), .Q(ereg[95]) );
  DFF \ereg_reg[96]  ( .D(n7602), .CLK(clk), .RST(rst), .Q(ereg[96]) );
  DFF \ereg_reg[97]  ( .D(n7601), .CLK(clk), .RST(rst), .Q(ereg[97]) );
  DFF \ereg_reg[98]  ( .D(n7600), .CLK(clk), .RST(rst), .Q(ereg[98]) );
  DFF \ereg_reg[99]  ( .D(n7599), .CLK(clk), .RST(rst), .Q(ereg[99]) );
  DFF \ereg_reg[100]  ( .D(n7598), .CLK(clk), .RST(rst), .Q(ereg[100]) );
  DFF \ereg_reg[101]  ( .D(n7597), .CLK(clk), .RST(rst), .Q(ereg[101]) );
  DFF \ereg_reg[102]  ( .D(n7596), .CLK(clk), .RST(rst), .Q(ereg[102]) );
  DFF \ereg_reg[103]  ( .D(n7595), .CLK(clk), .RST(rst), .Q(ereg[103]) );
  DFF \ereg_reg[104]  ( .D(n7594), .CLK(clk), .RST(rst), .Q(ereg[104]) );
  DFF \ereg_reg[105]  ( .D(n7593), .CLK(clk), .RST(rst), .Q(ereg[105]) );
  DFF \ereg_reg[106]  ( .D(n7592), .CLK(clk), .RST(rst), .Q(ereg[106]) );
  DFF \ereg_reg[107]  ( .D(n7591), .CLK(clk), .RST(rst), .Q(ereg[107]) );
  DFF \ereg_reg[108]  ( .D(n7590), .CLK(clk), .RST(rst), .Q(ereg[108]) );
  DFF \ereg_reg[109]  ( .D(n7589), .CLK(clk), .RST(rst), .Q(ereg[109]) );
  DFF \ereg_reg[110]  ( .D(n7588), .CLK(clk), .RST(rst), .Q(ereg[110]) );
  DFF \ereg_reg[111]  ( .D(n7587), .CLK(clk), .RST(rst), .Q(ereg[111]) );
  DFF \ereg_reg[112]  ( .D(n7586), .CLK(clk), .RST(rst), .Q(ereg[112]) );
  DFF \ereg_reg[113]  ( .D(n7585), .CLK(clk), .RST(rst), .Q(ereg[113]) );
  DFF \ereg_reg[114]  ( .D(n7584), .CLK(clk), .RST(rst), .Q(ereg[114]) );
  DFF \ereg_reg[115]  ( .D(n7583), .CLK(clk), .RST(rst), .Q(ereg[115]) );
  DFF \ereg_reg[116]  ( .D(n7582), .CLK(clk), .RST(rst), .Q(ereg[116]) );
  DFF \ereg_reg[117]  ( .D(n7581), .CLK(clk), .RST(rst), .Q(ereg[117]) );
  DFF \ereg_reg[118]  ( .D(n7580), .CLK(clk), .RST(rst), .Q(ereg[118]) );
  DFF \ereg_reg[119]  ( .D(n7579), .CLK(clk), .RST(rst), .Q(ereg[119]) );
  DFF \ereg_reg[120]  ( .D(n7578), .CLK(clk), .RST(rst), .Q(ereg[120]) );
  DFF \ereg_reg[121]  ( .D(n7577), .CLK(clk), .RST(rst), .Q(ereg[121]) );
  DFF \ereg_reg[122]  ( .D(n7576), .CLK(clk), .RST(rst), .Q(ereg[122]) );
  DFF \ereg_reg[123]  ( .D(n7575), .CLK(clk), .RST(rst), .Q(ereg[123]) );
  DFF \ereg_reg[124]  ( .D(n7574), .CLK(clk), .RST(rst), .Q(ereg[124]) );
  DFF \ereg_reg[125]  ( .D(n7573), .CLK(clk), .RST(rst), .Q(ereg[125]) );
  DFF \ereg_reg[126]  ( .D(n7572), .CLK(clk), .RST(rst), .Q(ereg[126]) );
  DFF \ereg_reg[127]  ( .D(n7571), .CLK(clk), .RST(rst), .Q(ereg[127]) );
  DFF \ereg_reg[128]  ( .D(n7570), .CLK(clk), .RST(rst), .Q(ereg[128]) );
  DFF \ereg_reg[129]  ( .D(n7569), .CLK(clk), .RST(rst), .Q(ereg[129]) );
  DFF \ereg_reg[130]  ( .D(n7568), .CLK(clk), .RST(rst), .Q(ereg[130]) );
  DFF \ereg_reg[131]  ( .D(n7567), .CLK(clk), .RST(rst), .Q(ereg[131]) );
  DFF \ereg_reg[132]  ( .D(n7566), .CLK(clk), .RST(rst), .Q(ereg[132]) );
  DFF \ereg_reg[133]  ( .D(n7565), .CLK(clk), .RST(rst), .Q(ereg[133]) );
  DFF \ereg_reg[134]  ( .D(n7564), .CLK(clk), .RST(rst), .Q(ereg[134]) );
  DFF \ereg_reg[135]  ( .D(n7563), .CLK(clk), .RST(rst), .Q(ereg[135]) );
  DFF \ereg_reg[136]  ( .D(n7562), .CLK(clk), .RST(rst), .Q(ereg[136]) );
  DFF \ereg_reg[137]  ( .D(n7561), .CLK(clk), .RST(rst), .Q(ereg[137]) );
  DFF \ereg_reg[138]  ( .D(n7560), .CLK(clk), .RST(rst), .Q(ereg[138]) );
  DFF \ereg_reg[139]  ( .D(n7559), .CLK(clk), .RST(rst), .Q(ereg[139]) );
  DFF \ereg_reg[140]  ( .D(n7558), .CLK(clk), .RST(rst), .Q(ereg[140]) );
  DFF \ereg_reg[141]  ( .D(n7557), .CLK(clk), .RST(rst), .Q(ereg[141]) );
  DFF \ereg_reg[142]  ( .D(n7556), .CLK(clk), .RST(rst), .Q(ereg[142]) );
  DFF \ereg_reg[143]  ( .D(n7555), .CLK(clk), .RST(rst), .Q(ereg[143]) );
  DFF \ereg_reg[144]  ( .D(n7554), .CLK(clk), .RST(rst), .Q(ereg[144]) );
  DFF \ereg_reg[145]  ( .D(n7553), .CLK(clk), .RST(rst), .Q(ereg[145]) );
  DFF \ereg_reg[146]  ( .D(n7552), .CLK(clk), .RST(rst), .Q(ereg[146]) );
  DFF \ereg_reg[147]  ( .D(n7551), .CLK(clk), .RST(rst), .Q(ereg[147]) );
  DFF \ereg_reg[148]  ( .D(n7550), .CLK(clk), .RST(rst), .Q(ereg[148]) );
  DFF \ereg_reg[149]  ( .D(n7549), .CLK(clk), .RST(rst), .Q(ereg[149]) );
  DFF \ereg_reg[150]  ( .D(n7548), .CLK(clk), .RST(rst), .Q(ereg[150]) );
  DFF \ereg_reg[151]  ( .D(n7547), .CLK(clk), .RST(rst), .Q(ereg[151]) );
  DFF \ereg_reg[152]  ( .D(n7546), .CLK(clk), .RST(rst), .Q(ereg[152]) );
  DFF \ereg_reg[153]  ( .D(n7545), .CLK(clk), .RST(rst), .Q(ereg[153]) );
  DFF \ereg_reg[154]  ( .D(n7544), .CLK(clk), .RST(rst), .Q(ereg[154]) );
  DFF \ereg_reg[155]  ( .D(n7543), .CLK(clk), .RST(rst), .Q(ereg[155]) );
  DFF \ereg_reg[156]  ( .D(n7542), .CLK(clk), .RST(rst), .Q(ereg[156]) );
  DFF \ereg_reg[157]  ( .D(n7541), .CLK(clk), .RST(rst), .Q(ereg[157]) );
  DFF \ereg_reg[158]  ( .D(n7540), .CLK(clk), .RST(rst), .Q(ereg[158]) );
  DFF \ereg_reg[159]  ( .D(n7539), .CLK(clk), .RST(rst), .Q(ereg[159]) );
  DFF \ereg_reg[160]  ( .D(n7538), .CLK(clk), .RST(rst), .Q(ereg[160]) );
  DFF \ereg_reg[161]  ( .D(n7537), .CLK(clk), .RST(rst), .Q(ereg[161]) );
  DFF \ereg_reg[162]  ( .D(n7536), .CLK(clk), .RST(rst), .Q(ereg[162]) );
  DFF \ereg_reg[163]  ( .D(n7535), .CLK(clk), .RST(rst), .Q(ereg[163]) );
  DFF \ereg_reg[164]  ( .D(n7534), .CLK(clk), .RST(rst), .Q(ereg[164]) );
  DFF \ereg_reg[165]  ( .D(n7533), .CLK(clk), .RST(rst), .Q(ereg[165]) );
  DFF \ereg_reg[166]  ( .D(n7532), .CLK(clk), .RST(rst), .Q(ereg[166]) );
  DFF \ereg_reg[167]  ( .D(n7531), .CLK(clk), .RST(rst), .Q(ereg[167]) );
  DFF \ereg_reg[168]  ( .D(n7530), .CLK(clk), .RST(rst), .Q(ereg[168]) );
  DFF \ereg_reg[169]  ( .D(n7529), .CLK(clk), .RST(rst), .Q(ereg[169]) );
  DFF \ereg_reg[170]  ( .D(n7528), .CLK(clk), .RST(rst), .Q(ereg[170]) );
  DFF \ereg_reg[171]  ( .D(n7527), .CLK(clk), .RST(rst), .Q(ereg[171]) );
  DFF \ereg_reg[172]  ( .D(n7526), .CLK(clk), .RST(rst), .Q(ereg[172]) );
  DFF \ereg_reg[173]  ( .D(n7525), .CLK(clk), .RST(rst), .Q(ereg[173]) );
  DFF \ereg_reg[174]  ( .D(n7524), .CLK(clk), .RST(rst), .Q(ereg[174]) );
  DFF \ereg_reg[175]  ( .D(n7523), .CLK(clk), .RST(rst), .Q(ereg[175]) );
  DFF \ereg_reg[176]  ( .D(n7522), .CLK(clk), .RST(rst), .Q(ereg[176]) );
  DFF \ereg_reg[177]  ( .D(n7521), .CLK(clk), .RST(rst), .Q(ereg[177]) );
  DFF \ereg_reg[178]  ( .D(n7520), .CLK(clk), .RST(rst), .Q(ereg[178]) );
  DFF \ereg_reg[179]  ( .D(n7519), .CLK(clk), .RST(rst), .Q(ereg[179]) );
  DFF \ereg_reg[180]  ( .D(n7518), .CLK(clk), .RST(rst), .Q(ereg[180]) );
  DFF \ereg_reg[181]  ( .D(n7517), .CLK(clk), .RST(rst), .Q(ereg[181]) );
  DFF \ereg_reg[182]  ( .D(n7516), .CLK(clk), .RST(rst), .Q(ereg[182]) );
  DFF \ereg_reg[183]  ( .D(n7515), .CLK(clk), .RST(rst), .Q(ereg[183]) );
  DFF \ereg_reg[184]  ( .D(n7514), .CLK(clk), .RST(rst), .Q(ereg[184]) );
  DFF \ereg_reg[185]  ( .D(n7513), .CLK(clk), .RST(rst), .Q(ereg[185]) );
  DFF \ereg_reg[186]  ( .D(n7512), .CLK(clk), .RST(rst), .Q(ereg[186]) );
  DFF \ereg_reg[187]  ( .D(n7511), .CLK(clk), .RST(rst), .Q(ereg[187]) );
  DFF \ereg_reg[188]  ( .D(n7510), .CLK(clk), .RST(rst), .Q(ereg[188]) );
  DFF \ereg_reg[189]  ( .D(n7509), .CLK(clk), .RST(rst), .Q(ereg[189]) );
  DFF \ereg_reg[190]  ( .D(n7508), .CLK(clk), .RST(rst), .Q(ereg[190]) );
  DFF \ereg_reg[191]  ( .D(n7507), .CLK(clk), .RST(rst), .Q(ereg[191]) );
  DFF \ereg_reg[192]  ( .D(n7506), .CLK(clk), .RST(rst), .Q(ereg[192]) );
  DFF \ereg_reg[193]  ( .D(n7505), .CLK(clk), .RST(rst), .Q(ereg[193]) );
  DFF \ereg_reg[194]  ( .D(n7504), .CLK(clk), .RST(rst), .Q(ereg[194]) );
  DFF \ereg_reg[195]  ( .D(n7503), .CLK(clk), .RST(rst), .Q(ereg[195]) );
  DFF \ereg_reg[196]  ( .D(n7502), .CLK(clk), .RST(rst), .Q(ereg[196]) );
  DFF \ereg_reg[197]  ( .D(n7501), .CLK(clk), .RST(rst), .Q(ereg[197]) );
  DFF \ereg_reg[198]  ( .D(n7500), .CLK(clk), .RST(rst), .Q(ereg[198]) );
  DFF \ereg_reg[199]  ( .D(n7499), .CLK(clk), .RST(rst), .Q(ereg[199]) );
  DFF \ereg_reg[200]  ( .D(n7498), .CLK(clk), .RST(rst), .Q(ereg[200]) );
  DFF \ereg_reg[201]  ( .D(n7497), .CLK(clk), .RST(rst), .Q(ereg[201]) );
  DFF \ereg_reg[202]  ( .D(n7496), .CLK(clk), .RST(rst), .Q(ereg[202]) );
  DFF \ereg_reg[203]  ( .D(n7495), .CLK(clk), .RST(rst), .Q(ereg[203]) );
  DFF \ereg_reg[204]  ( .D(n7494), .CLK(clk), .RST(rst), .Q(ereg[204]) );
  DFF \ereg_reg[205]  ( .D(n7493), .CLK(clk), .RST(rst), .Q(ereg[205]) );
  DFF \ereg_reg[206]  ( .D(n7492), .CLK(clk), .RST(rst), .Q(ereg[206]) );
  DFF \ereg_reg[207]  ( .D(n7491), .CLK(clk), .RST(rst), .Q(ereg[207]) );
  DFF \ereg_reg[208]  ( .D(n7490), .CLK(clk), .RST(rst), .Q(ereg[208]) );
  DFF \ereg_reg[209]  ( .D(n7489), .CLK(clk), .RST(rst), .Q(ereg[209]) );
  DFF \ereg_reg[210]  ( .D(n7488), .CLK(clk), .RST(rst), .Q(ereg[210]) );
  DFF \ereg_reg[211]  ( .D(n7487), .CLK(clk), .RST(rst), .Q(ereg[211]) );
  DFF \ereg_reg[212]  ( .D(n7486), .CLK(clk), .RST(rst), .Q(ereg[212]) );
  DFF \ereg_reg[213]  ( .D(n7485), .CLK(clk), .RST(rst), .Q(ereg[213]) );
  DFF \ereg_reg[214]  ( .D(n7484), .CLK(clk), .RST(rst), .Q(ereg[214]) );
  DFF \ereg_reg[215]  ( .D(n7483), .CLK(clk), .RST(rst), .Q(ereg[215]) );
  DFF \ereg_reg[216]  ( .D(n7482), .CLK(clk), .RST(rst), .Q(ereg[216]) );
  DFF \ereg_reg[217]  ( .D(n7481), .CLK(clk), .RST(rst), .Q(ereg[217]) );
  DFF \ereg_reg[218]  ( .D(n7480), .CLK(clk), .RST(rst), .Q(ereg[218]) );
  DFF \ereg_reg[219]  ( .D(n7479), .CLK(clk), .RST(rst), .Q(ereg[219]) );
  DFF \ereg_reg[220]  ( .D(n7478), .CLK(clk), .RST(rst), .Q(ereg[220]) );
  DFF \ereg_reg[221]  ( .D(n7477), .CLK(clk), .RST(rst), .Q(ereg[221]) );
  DFF \ereg_reg[222]  ( .D(n7476), .CLK(clk), .RST(rst), .Q(ereg[222]) );
  DFF \ereg_reg[223]  ( .D(n7475), .CLK(clk), .RST(rst), .Q(ereg[223]) );
  DFF \ereg_reg[224]  ( .D(n7474), .CLK(clk), .RST(rst), .Q(ereg[224]) );
  DFF \ereg_reg[225]  ( .D(n7473), .CLK(clk), .RST(rst), .Q(ereg[225]) );
  DFF \ereg_reg[226]  ( .D(n7472), .CLK(clk), .RST(rst), .Q(ereg[226]) );
  DFF \ereg_reg[227]  ( .D(n7471), .CLK(clk), .RST(rst), .Q(ereg[227]) );
  DFF \ereg_reg[228]  ( .D(n7470), .CLK(clk), .RST(rst), .Q(ereg[228]) );
  DFF \ereg_reg[229]  ( .D(n7469), .CLK(clk), .RST(rst), .Q(ereg[229]) );
  DFF \ereg_reg[230]  ( .D(n7468), .CLK(clk), .RST(rst), .Q(ereg[230]) );
  DFF \ereg_reg[231]  ( .D(n7467), .CLK(clk), .RST(rst), .Q(ereg[231]) );
  DFF \ereg_reg[232]  ( .D(n7466), .CLK(clk), .RST(rst), .Q(ereg[232]) );
  DFF \ereg_reg[233]  ( .D(n7465), .CLK(clk), .RST(rst), .Q(ereg[233]) );
  DFF \ereg_reg[234]  ( .D(n7464), .CLK(clk), .RST(rst), .Q(ereg[234]) );
  DFF \ereg_reg[235]  ( .D(n7463), .CLK(clk), .RST(rst), .Q(ereg[235]) );
  DFF \ereg_reg[236]  ( .D(n7462), .CLK(clk), .RST(rst), .Q(ereg[236]) );
  DFF \ereg_reg[237]  ( .D(n7461), .CLK(clk), .RST(rst), .Q(ereg[237]) );
  DFF \ereg_reg[238]  ( .D(n7460), .CLK(clk), .RST(rst), .Q(ereg[238]) );
  DFF \ereg_reg[239]  ( .D(n7459), .CLK(clk), .RST(rst), .Q(ereg[239]) );
  DFF \ereg_reg[240]  ( .D(n7458), .CLK(clk), .RST(rst), .Q(ereg[240]) );
  DFF \ereg_reg[241]  ( .D(n7457), .CLK(clk), .RST(rst), .Q(ereg[241]) );
  DFF \ereg_reg[242]  ( .D(n7456), .CLK(clk), .RST(rst), .Q(ereg[242]) );
  DFF \ereg_reg[243]  ( .D(n7455), .CLK(clk), .RST(rst), .Q(ereg[243]) );
  DFF \ereg_reg[244]  ( .D(n7454), .CLK(clk), .RST(rst), .Q(ereg[244]) );
  DFF \ereg_reg[245]  ( .D(n7453), .CLK(clk), .RST(rst), .Q(ereg[245]) );
  DFF \ereg_reg[246]  ( .D(n7452), .CLK(clk), .RST(rst), .Q(ereg[246]) );
  DFF \ereg_reg[247]  ( .D(n7451), .CLK(clk), .RST(rst), .Q(ereg[247]) );
  DFF \ereg_reg[248]  ( .D(n7450), .CLK(clk), .RST(rst), .Q(ereg[248]) );
  DFF \ereg_reg[249]  ( .D(n7449), .CLK(clk), .RST(rst), .Q(ereg[249]) );
  DFF \ereg_reg[250]  ( .D(n7448), .CLK(clk), .RST(rst), .Q(ereg[250]) );
  DFF \ereg_reg[251]  ( .D(n7447), .CLK(clk), .RST(rst), .Q(ereg[251]) );
  DFF \ereg_reg[252]  ( .D(n7446), .CLK(clk), .RST(rst), .Q(ereg[252]) );
  DFF \ereg_reg[253]  ( .D(n7445), .CLK(clk), .RST(rst), .Q(ereg[253]) );
  DFF \ereg_reg[254]  ( .D(n7444), .CLK(clk), .RST(rst), .Q(ereg[254]) );
  DFF \ereg_reg[255]  ( .D(n7443), .CLK(clk), .RST(rst), .Q(ereg[255]) );
  DFF \ereg_reg[256]  ( .D(n7442), .CLK(clk), .RST(rst), .Q(ereg[256]) );
  DFF \ereg_reg[257]  ( .D(n7441), .CLK(clk), .RST(rst), .Q(ereg[257]) );
  DFF \ereg_reg[258]  ( .D(n7440), .CLK(clk), .RST(rst), .Q(ereg[258]) );
  DFF \ereg_reg[259]  ( .D(n7439), .CLK(clk), .RST(rst), .Q(ereg[259]) );
  DFF \ereg_reg[260]  ( .D(n7438), .CLK(clk), .RST(rst), .Q(ereg[260]) );
  DFF \ereg_reg[261]  ( .D(n7437), .CLK(clk), .RST(rst), .Q(ereg[261]) );
  DFF \ereg_reg[262]  ( .D(n7436), .CLK(clk), .RST(rst), .Q(ereg[262]) );
  DFF \ereg_reg[263]  ( .D(n7435), .CLK(clk), .RST(rst), .Q(ereg[263]) );
  DFF \ereg_reg[264]  ( .D(n7434), .CLK(clk), .RST(rst), .Q(ereg[264]) );
  DFF \ereg_reg[265]  ( .D(n7433), .CLK(clk), .RST(rst), .Q(ereg[265]) );
  DFF \ereg_reg[266]  ( .D(n7432), .CLK(clk), .RST(rst), .Q(ereg[266]) );
  DFF \ereg_reg[267]  ( .D(n7431), .CLK(clk), .RST(rst), .Q(ereg[267]) );
  DFF \ereg_reg[268]  ( .D(n7430), .CLK(clk), .RST(rst), .Q(ereg[268]) );
  DFF \ereg_reg[269]  ( .D(n7429), .CLK(clk), .RST(rst), .Q(ereg[269]) );
  DFF \ereg_reg[270]  ( .D(n7428), .CLK(clk), .RST(rst), .Q(ereg[270]) );
  DFF \ereg_reg[271]  ( .D(n7427), .CLK(clk), .RST(rst), .Q(ereg[271]) );
  DFF \ereg_reg[272]  ( .D(n7426), .CLK(clk), .RST(rst), .Q(ereg[272]) );
  DFF \ereg_reg[273]  ( .D(n7425), .CLK(clk), .RST(rst), .Q(ereg[273]) );
  DFF \ereg_reg[274]  ( .D(n7424), .CLK(clk), .RST(rst), .Q(ereg[274]) );
  DFF \ereg_reg[275]  ( .D(n7423), .CLK(clk), .RST(rst), .Q(ereg[275]) );
  DFF \ereg_reg[276]  ( .D(n7422), .CLK(clk), .RST(rst), .Q(ereg[276]) );
  DFF \ereg_reg[277]  ( .D(n7421), .CLK(clk), .RST(rst), .Q(ereg[277]) );
  DFF \ereg_reg[278]  ( .D(n7420), .CLK(clk), .RST(rst), .Q(ereg[278]) );
  DFF \ereg_reg[279]  ( .D(n7419), .CLK(clk), .RST(rst), .Q(ereg[279]) );
  DFF \ereg_reg[280]  ( .D(n7418), .CLK(clk), .RST(rst), .Q(ereg[280]) );
  DFF \ereg_reg[281]  ( .D(n7417), .CLK(clk), .RST(rst), .Q(ereg[281]) );
  DFF \ereg_reg[282]  ( .D(n7416), .CLK(clk), .RST(rst), .Q(ereg[282]) );
  DFF \ereg_reg[283]  ( .D(n7415), .CLK(clk), .RST(rst), .Q(ereg[283]) );
  DFF \ereg_reg[284]  ( .D(n7414), .CLK(clk), .RST(rst), .Q(ereg[284]) );
  DFF \ereg_reg[285]  ( .D(n7413), .CLK(clk), .RST(rst), .Q(ereg[285]) );
  DFF \ereg_reg[286]  ( .D(n7412), .CLK(clk), .RST(rst), .Q(ereg[286]) );
  DFF \ereg_reg[287]  ( .D(n7411), .CLK(clk), .RST(rst), .Q(ereg[287]) );
  DFF \ereg_reg[288]  ( .D(n7410), .CLK(clk), .RST(rst), .Q(ereg[288]) );
  DFF \ereg_reg[289]  ( .D(n7409), .CLK(clk), .RST(rst), .Q(ereg[289]) );
  DFF \ereg_reg[290]  ( .D(n7408), .CLK(clk), .RST(rst), .Q(ereg[290]) );
  DFF \ereg_reg[291]  ( .D(n7407), .CLK(clk), .RST(rst), .Q(ereg[291]) );
  DFF \ereg_reg[292]  ( .D(n7406), .CLK(clk), .RST(rst), .Q(ereg[292]) );
  DFF \ereg_reg[293]  ( .D(n7405), .CLK(clk), .RST(rst), .Q(ereg[293]) );
  DFF \ereg_reg[294]  ( .D(n7404), .CLK(clk), .RST(rst), .Q(ereg[294]) );
  DFF \ereg_reg[295]  ( .D(n7403), .CLK(clk), .RST(rst), .Q(ereg[295]) );
  DFF \ereg_reg[296]  ( .D(n7402), .CLK(clk), .RST(rst), .Q(ereg[296]) );
  DFF \ereg_reg[297]  ( .D(n7401), .CLK(clk), .RST(rst), .Q(ereg[297]) );
  DFF \ereg_reg[298]  ( .D(n7400), .CLK(clk), .RST(rst), .Q(ereg[298]) );
  DFF \ereg_reg[299]  ( .D(n7399), .CLK(clk), .RST(rst), .Q(ereg[299]) );
  DFF \ereg_reg[300]  ( .D(n7398), .CLK(clk), .RST(rst), .Q(ereg[300]) );
  DFF \ereg_reg[301]  ( .D(n7397), .CLK(clk), .RST(rst), .Q(ereg[301]) );
  DFF \ereg_reg[302]  ( .D(n7396), .CLK(clk), .RST(rst), .Q(ereg[302]) );
  DFF \ereg_reg[303]  ( .D(n7395), .CLK(clk), .RST(rst), .Q(ereg[303]) );
  DFF \ereg_reg[304]  ( .D(n7394), .CLK(clk), .RST(rst), .Q(ereg[304]) );
  DFF \ereg_reg[305]  ( .D(n7393), .CLK(clk), .RST(rst), .Q(ereg[305]) );
  DFF \ereg_reg[306]  ( .D(n7392), .CLK(clk), .RST(rst), .Q(ereg[306]) );
  DFF \ereg_reg[307]  ( .D(n7391), .CLK(clk), .RST(rst), .Q(ereg[307]) );
  DFF \ereg_reg[308]  ( .D(n7390), .CLK(clk), .RST(rst), .Q(ereg[308]) );
  DFF \ereg_reg[309]  ( .D(n7389), .CLK(clk), .RST(rst), .Q(ereg[309]) );
  DFF \ereg_reg[310]  ( .D(n7388), .CLK(clk), .RST(rst), .Q(ereg[310]) );
  DFF \ereg_reg[311]  ( .D(n7387), .CLK(clk), .RST(rst), .Q(ereg[311]) );
  DFF \ereg_reg[312]  ( .D(n7386), .CLK(clk), .RST(rst), .Q(ereg[312]) );
  DFF \ereg_reg[313]  ( .D(n7385), .CLK(clk), .RST(rst), .Q(ereg[313]) );
  DFF \ereg_reg[314]  ( .D(n7384), .CLK(clk), .RST(rst), .Q(ereg[314]) );
  DFF \ereg_reg[315]  ( .D(n7383), .CLK(clk), .RST(rst), .Q(ereg[315]) );
  DFF \ereg_reg[316]  ( .D(n7382), .CLK(clk), .RST(rst), .Q(ereg[316]) );
  DFF \ereg_reg[317]  ( .D(n7381), .CLK(clk), .RST(rst), .Q(ereg[317]) );
  DFF \ereg_reg[318]  ( .D(n7380), .CLK(clk), .RST(rst), .Q(ereg[318]) );
  DFF \ereg_reg[319]  ( .D(n7379), .CLK(clk), .RST(rst), .Q(ereg[319]) );
  DFF \ereg_reg[320]  ( .D(n7378), .CLK(clk), .RST(rst), .Q(ereg[320]) );
  DFF \ereg_reg[321]  ( .D(n7377), .CLK(clk), .RST(rst), .Q(ereg[321]) );
  DFF \ereg_reg[322]  ( .D(n7376), .CLK(clk), .RST(rst), .Q(ereg[322]) );
  DFF \ereg_reg[323]  ( .D(n7375), .CLK(clk), .RST(rst), .Q(ereg[323]) );
  DFF \ereg_reg[324]  ( .D(n7374), .CLK(clk), .RST(rst), .Q(ereg[324]) );
  DFF \ereg_reg[325]  ( .D(n7373), .CLK(clk), .RST(rst), .Q(ereg[325]) );
  DFF \ereg_reg[326]  ( .D(n7372), .CLK(clk), .RST(rst), .Q(ereg[326]) );
  DFF \ereg_reg[327]  ( .D(n7371), .CLK(clk), .RST(rst), .Q(ereg[327]) );
  DFF \ereg_reg[328]  ( .D(n7370), .CLK(clk), .RST(rst), .Q(ereg[328]) );
  DFF \ereg_reg[329]  ( .D(n7369), .CLK(clk), .RST(rst), .Q(ereg[329]) );
  DFF \ereg_reg[330]  ( .D(n7368), .CLK(clk), .RST(rst), .Q(ereg[330]) );
  DFF \ereg_reg[331]  ( .D(n7367), .CLK(clk), .RST(rst), .Q(ereg[331]) );
  DFF \ereg_reg[332]  ( .D(n7366), .CLK(clk), .RST(rst), .Q(ereg[332]) );
  DFF \ereg_reg[333]  ( .D(n7365), .CLK(clk), .RST(rst), .Q(ereg[333]) );
  DFF \ereg_reg[334]  ( .D(n7364), .CLK(clk), .RST(rst), .Q(ereg[334]) );
  DFF \ereg_reg[335]  ( .D(n7363), .CLK(clk), .RST(rst), .Q(ereg[335]) );
  DFF \ereg_reg[336]  ( .D(n7362), .CLK(clk), .RST(rst), .Q(ereg[336]) );
  DFF \ereg_reg[337]  ( .D(n7361), .CLK(clk), .RST(rst), .Q(ereg[337]) );
  DFF \ereg_reg[338]  ( .D(n7360), .CLK(clk), .RST(rst), .Q(ereg[338]) );
  DFF \ereg_reg[339]  ( .D(n7359), .CLK(clk), .RST(rst), .Q(ereg[339]) );
  DFF \ereg_reg[340]  ( .D(n7358), .CLK(clk), .RST(rst), .Q(ereg[340]) );
  DFF \ereg_reg[341]  ( .D(n7357), .CLK(clk), .RST(rst), .Q(ereg[341]) );
  DFF \ereg_reg[342]  ( .D(n7356), .CLK(clk), .RST(rst), .Q(ereg[342]) );
  DFF \ereg_reg[343]  ( .D(n7355), .CLK(clk), .RST(rst), .Q(ereg[343]) );
  DFF \ereg_reg[344]  ( .D(n7354), .CLK(clk), .RST(rst), .Q(ereg[344]) );
  DFF \ereg_reg[345]  ( .D(n7353), .CLK(clk), .RST(rst), .Q(ereg[345]) );
  DFF \ereg_reg[346]  ( .D(n7352), .CLK(clk), .RST(rst), .Q(ereg[346]) );
  DFF \ereg_reg[347]  ( .D(n7351), .CLK(clk), .RST(rst), .Q(ereg[347]) );
  DFF \ereg_reg[348]  ( .D(n7350), .CLK(clk), .RST(rst), .Q(ereg[348]) );
  DFF \ereg_reg[349]  ( .D(n7349), .CLK(clk), .RST(rst), .Q(ereg[349]) );
  DFF \ereg_reg[350]  ( .D(n7348), .CLK(clk), .RST(rst), .Q(ereg[350]) );
  DFF \ereg_reg[351]  ( .D(n7347), .CLK(clk), .RST(rst), .Q(ereg[351]) );
  DFF \ereg_reg[352]  ( .D(n7346), .CLK(clk), .RST(rst), .Q(ereg[352]) );
  DFF \ereg_reg[353]  ( .D(n7345), .CLK(clk), .RST(rst), .Q(ereg[353]) );
  DFF \ereg_reg[354]  ( .D(n7344), .CLK(clk), .RST(rst), .Q(ereg[354]) );
  DFF \ereg_reg[355]  ( .D(n7343), .CLK(clk), .RST(rst), .Q(ereg[355]) );
  DFF \ereg_reg[356]  ( .D(n7342), .CLK(clk), .RST(rst), .Q(ereg[356]) );
  DFF \ereg_reg[357]  ( .D(n7341), .CLK(clk), .RST(rst), .Q(ereg[357]) );
  DFF \ereg_reg[358]  ( .D(n7340), .CLK(clk), .RST(rst), .Q(ereg[358]) );
  DFF \ereg_reg[359]  ( .D(n7339), .CLK(clk), .RST(rst), .Q(ereg[359]) );
  DFF \ereg_reg[360]  ( .D(n7338), .CLK(clk), .RST(rst), .Q(ereg[360]) );
  DFF \ereg_reg[361]  ( .D(n7337), .CLK(clk), .RST(rst), .Q(ereg[361]) );
  DFF \ereg_reg[362]  ( .D(n7336), .CLK(clk), .RST(rst), .Q(ereg[362]) );
  DFF \ereg_reg[363]  ( .D(n7335), .CLK(clk), .RST(rst), .Q(ereg[363]) );
  DFF \ereg_reg[364]  ( .D(n7334), .CLK(clk), .RST(rst), .Q(ereg[364]) );
  DFF \ereg_reg[365]  ( .D(n7333), .CLK(clk), .RST(rst), .Q(ereg[365]) );
  DFF \ereg_reg[366]  ( .D(n7332), .CLK(clk), .RST(rst), .Q(ereg[366]) );
  DFF \ereg_reg[367]  ( .D(n7331), .CLK(clk), .RST(rst), .Q(ereg[367]) );
  DFF \ereg_reg[368]  ( .D(n7330), .CLK(clk), .RST(rst), .Q(ereg[368]) );
  DFF \ereg_reg[369]  ( .D(n7329), .CLK(clk), .RST(rst), .Q(ereg[369]) );
  DFF \ereg_reg[370]  ( .D(n7328), .CLK(clk), .RST(rst), .Q(ereg[370]) );
  DFF \ereg_reg[371]  ( .D(n7327), .CLK(clk), .RST(rst), .Q(ereg[371]) );
  DFF \ereg_reg[372]  ( .D(n7326), .CLK(clk), .RST(rst), .Q(ereg[372]) );
  DFF \ereg_reg[373]  ( .D(n7325), .CLK(clk), .RST(rst), .Q(ereg[373]) );
  DFF \ereg_reg[374]  ( .D(n7324), .CLK(clk), .RST(rst), .Q(ereg[374]) );
  DFF \ereg_reg[375]  ( .D(n7323), .CLK(clk), .RST(rst), .Q(ereg[375]) );
  DFF \ereg_reg[376]  ( .D(n7322), .CLK(clk), .RST(rst), .Q(ereg[376]) );
  DFF \ereg_reg[377]  ( .D(n7321), .CLK(clk), .RST(rst), .Q(ereg[377]) );
  DFF \ereg_reg[378]  ( .D(n7320), .CLK(clk), .RST(rst), .Q(ereg[378]) );
  DFF \ereg_reg[379]  ( .D(n7319), .CLK(clk), .RST(rst), .Q(ereg[379]) );
  DFF \ereg_reg[380]  ( .D(n7318), .CLK(clk), .RST(rst), .Q(ereg[380]) );
  DFF \ereg_reg[381]  ( .D(n7317), .CLK(clk), .RST(rst), .Q(ereg[381]) );
  DFF \ereg_reg[382]  ( .D(n7316), .CLK(clk), .RST(rst), .Q(ereg[382]) );
  DFF \ereg_reg[383]  ( .D(n7315), .CLK(clk), .RST(rst), .Q(ereg[383]) );
  DFF \ereg_reg[384]  ( .D(n7314), .CLK(clk), .RST(rst), .Q(ereg[384]) );
  DFF \ereg_reg[385]  ( .D(n7313), .CLK(clk), .RST(rst), .Q(ereg[385]) );
  DFF \ereg_reg[386]  ( .D(n7312), .CLK(clk), .RST(rst), .Q(ereg[386]) );
  DFF \ereg_reg[387]  ( .D(n7311), .CLK(clk), .RST(rst), .Q(ereg[387]) );
  DFF \ereg_reg[388]  ( .D(n7310), .CLK(clk), .RST(rst), .Q(ereg[388]) );
  DFF \ereg_reg[389]  ( .D(n7309), .CLK(clk), .RST(rst), .Q(ereg[389]) );
  DFF \ereg_reg[390]  ( .D(n7308), .CLK(clk), .RST(rst), .Q(ereg[390]) );
  DFF \ereg_reg[391]  ( .D(n7307), .CLK(clk), .RST(rst), .Q(ereg[391]) );
  DFF \ereg_reg[392]  ( .D(n7306), .CLK(clk), .RST(rst), .Q(ereg[392]) );
  DFF \ereg_reg[393]  ( .D(n7305), .CLK(clk), .RST(rst), .Q(ereg[393]) );
  DFF \ereg_reg[394]  ( .D(n7304), .CLK(clk), .RST(rst), .Q(ereg[394]) );
  DFF \ereg_reg[395]  ( .D(n7303), .CLK(clk), .RST(rst), .Q(ereg[395]) );
  DFF \ereg_reg[396]  ( .D(n7302), .CLK(clk), .RST(rst), .Q(ereg[396]) );
  DFF \ereg_reg[397]  ( .D(n7301), .CLK(clk), .RST(rst), .Q(ereg[397]) );
  DFF \ereg_reg[398]  ( .D(n7300), .CLK(clk), .RST(rst), .Q(ereg[398]) );
  DFF \ereg_reg[399]  ( .D(n7299), .CLK(clk), .RST(rst), .Q(ereg[399]) );
  DFF \ereg_reg[400]  ( .D(n7298), .CLK(clk), .RST(rst), .Q(ereg[400]) );
  DFF \ereg_reg[401]  ( .D(n7297), .CLK(clk), .RST(rst), .Q(ereg[401]) );
  DFF \ereg_reg[402]  ( .D(n7296), .CLK(clk), .RST(rst), .Q(ereg[402]) );
  DFF \ereg_reg[403]  ( .D(n7295), .CLK(clk), .RST(rst), .Q(ereg[403]) );
  DFF \ereg_reg[404]  ( .D(n7294), .CLK(clk), .RST(rst), .Q(ereg[404]) );
  DFF \ereg_reg[405]  ( .D(n7293), .CLK(clk), .RST(rst), .Q(ereg[405]) );
  DFF \ereg_reg[406]  ( .D(n7292), .CLK(clk), .RST(rst), .Q(ereg[406]) );
  DFF \ereg_reg[407]  ( .D(n7291), .CLK(clk), .RST(rst), .Q(ereg[407]) );
  DFF \ereg_reg[408]  ( .D(n7290), .CLK(clk), .RST(rst), .Q(ereg[408]) );
  DFF \ereg_reg[409]  ( .D(n7289), .CLK(clk), .RST(rst), .Q(ereg[409]) );
  DFF \ereg_reg[410]  ( .D(n7288), .CLK(clk), .RST(rst), .Q(ereg[410]) );
  DFF \ereg_reg[411]  ( .D(n7287), .CLK(clk), .RST(rst), .Q(ereg[411]) );
  DFF \ereg_reg[412]  ( .D(n7286), .CLK(clk), .RST(rst), .Q(ereg[412]) );
  DFF \ereg_reg[413]  ( .D(n7285), .CLK(clk), .RST(rst), .Q(ereg[413]) );
  DFF \ereg_reg[414]  ( .D(n7284), .CLK(clk), .RST(rst), .Q(ereg[414]) );
  DFF \ereg_reg[415]  ( .D(n7283), .CLK(clk), .RST(rst), .Q(ereg[415]) );
  DFF \ereg_reg[416]  ( .D(n7282), .CLK(clk), .RST(rst), .Q(ereg[416]) );
  DFF \ereg_reg[417]  ( .D(n7281), .CLK(clk), .RST(rst), .Q(ereg[417]) );
  DFF \ereg_reg[418]  ( .D(n7280), .CLK(clk), .RST(rst), .Q(ereg[418]) );
  DFF \ereg_reg[419]  ( .D(n7279), .CLK(clk), .RST(rst), .Q(ereg[419]) );
  DFF \ereg_reg[420]  ( .D(n7278), .CLK(clk), .RST(rst), .Q(ereg[420]) );
  DFF \ereg_reg[421]  ( .D(n7277), .CLK(clk), .RST(rst), .Q(ereg[421]) );
  DFF \ereg_reg[422]  ( .D(n7276), .CLK(clk), .RST(rst), .Q(ereg[422]) );
  DFF \ereg_reg[423]  ( .D(n7275), .CLK(clk), .RST(rst), .Q(ereg[423]) );
  DFF \ereg_reg[424]  ( .D(n7274), .CLK(clk), .RST(rst), .Q(ereg[424]) );
  DFF \ereg_reg[425]  ( .D(n7273), .CLK(clk), .RST(rst), .Q(ereg[425]) );
  DFF \ereg_reg[426]  ( .D(n7272), .CLK(clk), .RST(rst), .Q(ereg[426]) );
  DFF \ereg_reg[427]  ( .D(n7271), .CLK(clk), .RST(rst), .Q(ereg[427]) );
  DFF \ereg_reg[428]  ( .D(n7270), .CLK(clk), .RST(rst), .Q(ereg[428]) );
  DFF \ereg_reg[429]  ( .D(n7269), .CLK(clk), .RST(rst), .Q(ereg[429]) );
  DFF \ereg_reg[430]  ( .D(n7268), .CLK(clk), .RST(rst), .Q(ereg[430]) );
  DFF \ereg_reg[431]  ( .D(n7267), .CLK(clk), .RST(rst), .Q(ereg[431]) );
  DFF \ereg_reg[432]  ( .D(n7266), .CLK(clk), .RST(rst), .Q(ereg[432]) );
  DFF \ereg_reg[433]  ( .D(n7265), .CLK(clk), .RST(rst), .Q(ereg[433]) );
  DFF \ereg_reg[434]  ( .D(n7264), .CLK(clk), .RST(rst), .Q(ereg[434]) );
  DFF \ereg_reg[435]  ( .D(n7263), .CLK(clk), .RST(rst), .Q(ereg[435]) );
  DFF \ereg_reg[436]  ( .D(n7262), .CLK(clk), .RST(rst), .Q(ereg[436]) );
  DFF \ereg_reg[437]  ( .D(n7261), .CLK(clk), .RST(rst), .Q(ereg[437]) );
  DFF \ereg_reg[438]  ( .D(n7260), .CLK(clk), .RST(rst), .Q(ereg[438]) );
  DFF \ereg_reg[439]  ( .D(n7259), .CLK(clk), .RST(rst), .Q(ereg[439]) );
  DFF \ereg_reg[440]  ( .D(n7258), .CLK(clk), .RST(rst), .Q(ereg[440]) );
  DFF \ereg_reg[441]  ( .D(n7257), .CLK(clk), .RST(rst), .Q(ereg[441]) );
  DFF \ereg_reg[442]  ( .D(n7256), .CLK(clk), .RST(rst), .Q(ereg[442]) );
  DFF \ereg_reg[443]  ( .D(n7255), .CLK(clk), .RST(rst), .Q(ereg[443]) );
  DFF \ereg_reg[444]  ( .D(n7254), .CLK(clk), .RST(rst), .Q(ereg[444]) );
  DFF \ereg_reg[445]  ( .D(n7253), .CLK(clk), .RST(rst), .Q(ereg[445]) );
  DFF \ereg_reg[446]  ( .D(n7252), .CLK(clk), .RST(rst), .Q(ereg[446]) );
  DFF \ereg_reg[447]  ( .D(n7251), .CLK(clk), .RST(rst), .Q(ereg[447]) );
  DFF \ereg_reg[448]  ( .D(n7250), .CLK(clk), .RST(rst), .Q(ereg[448]) );
  DFF \ereg_reg[449]  ( .D(n7249), .CLK(clk), .RST(rst), .Q(ereg[449]) );
  DFF \ereg_reg[450]  ( .D(n7248), .CLK(clk), .RST(rst), .Q(ereg[450]) );
  DFF \ereg_reg[451]  ( .D(n7247), .CLK(clk), .RST(rst), .Q(ereg[451]) );
  DFF \ereg_reg[452]  ( .D(n7246), .CLK(clk), .RST(rst), .Q(ereg[452]) );
  DFF \ereg_reg[453]  ( .D(n7245), .CLK(clk), .RST(rst), .Q(ereg[453]) );
  DFF \ereg_reg[454]  ( .D(n7244), .CLK(clk), .RST(rst), .Q(ereg[454]) );
  DFF \ereg_reg[455]  ( .D(n7243), .CLK(clk), .RST(rst), .Q(ereg[455]) );
  DFF \ereg_reg[456]  ( .D(n7242), .CLK(clk), .RST(rst), .Q(ereg[456]) );
  DFF \ereg_reg[457]  ( .D(n7241), .CLK(clk), .RST(rst), .Q(ereg[457]) );
  DFF \ereg_reg[458]  ( .D(n7240), .CLK(clk), .RST(rst), .Q(ereg[458]) );
  DFF \ereg_reg[459]  ( .D(n7239), .CLK(clk), .RST(rst), .Q(ereg[459]) );
  DFF \ereg_reg[460]  ( .D(n7238), .CLK(clk), .RST(rst), .Q(ereg[460]) );
  DFF \ereg_reg[461]  ( .D(n7237), .CLK(clk), .RST(rst), .Q(ereg[461]) );
  DFF \ereg_reg[462]  ( .D(n7236), .CLK(clk), .RST(rst), .Q(ereg[462]) );
  DFF \ereg_reg[463]  ( .D(n7235), .CLK(clk), .RST(rst), .Q(ereg[463]) );
  DFF \ereg_reg[464]  ( .D(n7234), .CLK(clk), .RST(rst), .Q(ereg[464]) );
  DFF \ereg_reg[465]  ( .D(n7233), .CLK(clk), .RST(rst), .Q(ereg[465]) );
  DFF \ereg_reg[466]  ( .D(n7232), .CLK(clk), .RST(rst), .Q(ereg[466]) );
  DFF \ereg_reg[467]  ( .D(n7231), .CLK(clk), .RST(rst), .Q(ereg[467]) );
  DFF \ereg_reg[468]  ( .D(n7230), .CLK(clk), .RST(rst), .Q(ereg[468]) );
  DFF \ereg_reg[469]  ( .D(n7229), .CLK(clk), .RST(rst), .Q(ereg[469]) );
  DFF \ereg_reg[470]  ( .D(n7228), .CLK(clk), .RST(rst), .Q(ereg[470]) );
  DFF \ereg_reg[471]  ( .D(n7227), .CLK(clk), .RST(rst), .Q(ereg[471]) );
  DFF \ereg_reg[472]  ( .D(n7226), .CLK(clk), .RST(rst), .Q(ereg[472]) );
  DFF \ereg_reg[473]  ( .D(n7225), .CLK(clk), .RST(rst), .Q(ereg[473]) );
  DFF \ereg_reg[474]  ( .D(n7224), .CLK(clk), .RST(rst), .Q(ereg[474]) );
  DFF \ereg_reg[475]  ( .D(n7223), .CLK(clk), .RST(rst), .Q(ereg[475]) );
  DFF \ereg_reg[476]  ( .D(n7222), .CLK(clk), .RST(rst), .Q(ereg[476]) );
  DFF \ereg_reg[477]  ( .D(n7221), .CLK(clk), .RST(rst), .Q(ereg[477]) );
  DFF \ereg_reg[478]  ( .D(n7220), .CLK(clk), .RST(rst), .Q(ereg[478]) );
  DFF \ereg_reg[479]  ( .D(n7219), .CLK(clk), .RST(rst), .Q(ereg[479]) );
  DFF \ereg_reg[480]  ( .D(n7218), .CLK(clk), .RST(rst), .Q(ereg[480]) );
  DFF \ereg_reg[481]  ( .D(n7217), .CLK(clk), .RST(rst), .Q(ereg[481]) );
  DFF \ereg_reg[482]  ( .D(n7216), .CLK(clk), .RST(rst), .Q(ereg[482]) );
  DFF \ereg_reg[483]  ( .D(n7215), .CLK(clk), .RST(rst), .Q(ereg[483]) );
  DFF \ereg_reg[484]  ( .D(n7214), .CLK(clk), .RST(rst), .Q(ereg[484]) );
  DFF \ereg_reg[485]  ( .D(n7213), .CLK(clk), .RST(rst), .Q(ereg[485]) );
  DFF \ereg_reg[486]  ( .D(n7212), .CLK(clk), .RST(rst), .Q(ereg[486]) );
  DFF \ereg_reg[487]  ( .D(n7211), .CLK(clk), .RST(rst), .Q(ereg[487]) );
  DFF \ereg_reg[488]  ( .D(n7210), .CLK(clk), .RST(rst), .Q(ereg[488]) );
  DFF \ereg_reg[489]  ( .D(n7209), .CLK(clk), .RST(rst), .Q(ereg[489]) );
  DFF \ereg_reg[490]  ( .D(n7208), .CLK(clk), .RST(rst), .Q(ereg[490]) );
  DFF \ereg_reg[491]  ( .D(n7207), .CLK(clk), .RST(rst), .Q(ereg[491]) );
  DFF \ereg_reg[492]  ( .D(n7206), .CLK(clk), .RST(rst), .Q(ereg[492]) );
  DFF \ereg_reg[493]  ( .D(n7205), .CLK(clk), .RST(rst), .Q(ereg[493]) );
  DFF \ereg_reg[494]  ( .D(n7204), .CLK(clk), .RST(rst), .Q(ereg[494]) );
  DFF \ereg_reg[495]  ( .D(n7203), .CLK(clk), .RST(rst), .Q(ereg[495]) );
  DFF \ereg_reg[496]  ( .D(n7202), .CLK(clk), .RST(rst), .Q(ereg[496]) );
  DFF \ereg_reg[497]  ( .D(n7201), .CLK(clk), .RST(rst), .Q(ereg[497]) );
  DFF \ereg_reg[498]  ( .D(n7200), .CLK(clk), .RST(rst), .Q(ereg[498]) );
  DFF \ereg_reg[499]  ( .D(n7199), .CLK(clk), .RST(rst), .Q(ereg[499]) );
  DFF \ereg_reg[500]  ( .D(n7198), .CLK(clk), .RST(rst), .Q(ereg[500]) );
  DFF \ereg_reg[501]  ( .D(n7197), .CLK(clk), .RST(rst), .Q(ereg[501]) );
  DFF \ereg_reg[502]  ( .D(n7196), .CLK(clk), .RST(rst), .Q(ereg[502]) );
  DFF \ereg_reg[503]  ( .D(n7195), .CLK(clk), .RST(rst), .Q(ereg[503]) );
  DFF \ereg_reg[504]  ( .D(n7194), .CLK(clk), .RST(rst), .Q(ereg[504]) );
  DFF \ereg_reg[505]  ( .D(n7193), .CLK(clk), .RST(rst), .Q(ereg[505]) );
  DFF \ereg_reg[506]  ( .D(n7192), .CLK(clk), .RST(rst), .Q(ereg[506]) );
  DFF \ereg_reg[507]  ( .D(n7191), .CLK(clk), .RST(rst), .Q(ereg[507]) );
  DFF \ereg_reg[508]  ( .D(n7190), .CLK(clk), .RST(rst), .Q(ereg[508]) );
  DFF \ereg_reg[509]  ( .D(n7189), .CLK(clk), .RST(rst), .Q(ereg[509]) );
  DFF \ereg_reg[510]  ( .D(n7188), .CLK(clk), .RST(rst), .Q(ereg[510]) );
  DFF \ereg_reg[511]  ( .D(n7187), .CLK(clk), .RST(rst), .Q(ereg[511]) );
  DFF first_one_reg ( .D(n6674), .CLK(clk), .RST(rst), .Q(first_one) );
  DFF \creg_reg[0]  ( .D(n7185), .CLK(clk), .RST(rst), .Q(creg[0]) );
  DFF \creg_reg[1]  ( .D(n7184), .CLK(clk), .RST(rst), .Q(creg[1]) );
  DFF \creg_reg[2]  ( .D(n7183), .CLK(clk), .RST(rst), .Q(creg[2]) );
  DFF \creg_reg[3]  ( .D(n7182), .CLK(clk), .RST(rst), .Q(creg[3]) );
  DFF \creg_reg[4]  ( .D(n7181), .CLK(clk), .RST(rst), .Q(creg[4]) );
  DFF \creg_reg[5]  ( .D(n7180), .CLK(clk), .RST(rst), .Q(creg[5]) );
  DFF \creg_reg[6]  ( .D(n7179), .CLK(clk), .RST(rst), .Q(creg[6]) );
  DFF \creg_reg[7]  ( .D(n7178), .CLK(clk), .RST(rst), .Q(creg[7]) );
  DFF \creg_reg[8]  ( .D(n7177), .CLK(clk), .RST(rst), .Q(creg[8]) );
  DFF \creg_reg[9]  ( .D(n7176), .CLK(clk), .RST(rst), .Q(creg[9]) );
  DFF \creg_reg[10]  ( .D(n7175), .CLK(clk), .RST(rst), .Q(creg[10]) );
  DFF \creg_reg[11]  ( .D(n7174), .CLK(clk), .RST(rst), .Q(creg[11]) );
  DFF \creg_reg[12]  ( .D(n7173), .CLK(clk), .RST(rst), .Q(creg[12]) );
  DFF \creg_reg[13]  ( .D(n7172), .CLK(clk), .RST(rst), .Q(creg[13]) );
  DFF \creg_reg[14]  ( .D(n7171), .CLK(clk), .RST(rst), .Q(creg[14]) );
  DFF \creg_reg[15]  ( .D(n7170), .CLK(clk), .RST(rst), .Q(creg[15]) );
  DFF \creg_reg[16]  ( .D(n7169), .CLK(clk), .RST(rst), .Q(creg[16]) );
  DFF \creg_reg[17]  ( .D(n7168), .CLK(clk), .RST(rst), .Q(creg[17]) );
  DFF \creg_reg[18]  ( .D(n7167), .CLK(clk), .RST(rst), .Q(creg[18]) );
  DFF \creg_reg[19]  ( .D(n7166), .CLK(clk), .RST(rst), .Q(creg[19]) );
  DFF \creg_reg[20]  ( .D(n7165), .CLK(clk), .RST(rst), .Q(creg[20]) );
  DFF \creg_reg[21]  ( .D(n7164), .CLK(clk), .RST(rst), .Q(creg[21]) );
  DFF \creg_reg[22]  ( .D(n7163), .CLK(clk), .RST(rst), .Q(creg[22]) );
  DFF \creg_reg[23]  ( .D(n7162), .CLK(clk), .RST(rst), .Q(creg[23]) );
  DFF \creg_reg[24]  ( .D(n7161), .CLK(clk), .RST(rst), .Q(creg[24]) );
  DFF \creg_reg[25]  ( .D(n7160), .CLK(clk), .RST(rst), .Q(creg[25]) );
  DFF \creg_reg[26]  ( .D(n7159), .CLK(clk), .RST(rst), .Q(creg[26]) );
  DFF \creg_reg[27]  ( .D(n7158), .CLK(clk), .RST(rst), .Q(creg[27]) );
  DFF \creg_reg[28]  ( .D(n7157), .CLK(clk), .RST(rst), .Q(creg[28]) );
  DFF \creg_reg[29]  ( .D(n7156), .CLK(clk), .RST(rst), .Q(creg[29]) );
  DFF \creg_reg[30]  ( .D(n7155), .CLK(clk), .RST(rst), .Q(creg[30]) );
  DFF \creg_reg[31]  ( .D(n7154), .CLK(clk), .RST(rst), .Q(creg[31]) );
  DFF \creg_reg[32]  ( .D(n7153), .CLK(clk), .RST(rst), .Q(creg[32]) );
  DFF \creg_reg[33]  ( .D(n7152), .CLK(clk), .RST(rst), .Q(creg[33]) );
  DFF \creg_reg[34]  ( .D(n7151), .CLK(clk), .RST(rst), .Q(creg[34]) );
  DFF \creg_reg[35]  ( .D(n7150), .CLK(clk), .RST(rst), .Q(creg[35]) );
  DFF \creg_reg[36]  ( .D(n7149), .CLK(clk), .RST(rst), .Q(creg[36]) );
  DFF \creg_reg[37]  ( .D(n7148), .CLK(clk), .RST(rst), .Q(creg[37]) );
  DFF \creg_reg[38]  ( .D(n7147), .CLK(clk), .RST(rst), .Q(creg[38]) );
  DFF \creg_reg[39]  ( .D(n7146), .CLK(clk), .RST(rst), .Q(creg[39]) );
  DFF \creg_reg[40]  ( .D(n7145), .CLK(clk), .RST(rst), .Q(creg[40]) );
  DFF \creg_reg[41]  ( .D(n7144), .CLK(clk), .RST(rst), .Q(creg[41]) );
  DFF \creg_reg[42]  ( .D(n7143), .CLK(clk), .RST(rst), .Q(creg[42]) );
  DFF \creg_reg[43]  ( .D(n7142), .CLK(clk), .RST(rst), .Q(creg[43]) );
  DFF \creg_reg[44]  ( .D(n7141), .CLK(clk), .RST(rst), .Q(creg[44]) );
  DFF \creg_reg[45]  ( .D(n7140), .CLK(clk), .RST(rst), .Q(creg[45]) );
  DFF \creg_reg[46]  ( .D(n7139), .CLK(clk), .RST(rst), .Q(creg[46]) );
  DFF \creg_reg[47]  ( .D(n7138), .CLK(clk), .RST(rst), .Q(creg[47]) );
  DFF \creg_reg[48]  ( .D(n7137), .CLK(clk), .RST(rst), .Q(creg[48]) );
  DFF \creg_reg[49]  ( .D(n7136), .CLK(clk), .RST(rst), .Q(creg[49]) );
  DFF \creg_reg[50]  ( .D(n7135), .CLK(clk), .RST(rst), .Q(creg[50]) );
  DFF \creg_reg[51]  ( .D(n7134), .CLK(clk), .RST(rst), .Q(creg[51]) );
  DFF \creg_reg[52]  ( .D(n7133), .CLK(clk), .RST(rst), .Q(creg[52]) );
  DFF \creg_reg[53]  ( .D(n7132), .CLK(clk), .RST(rst), .Q(creg[53]) );
  DFF \creg_reg[54]  ( .D(n7131), .CLK(clk), .RST(rst), .Q(creg[54]) );
  DFF \creg_reg[55]  ( .D(n7130), .CLK(clk), .RST(rst), .Q(creg[55]) );
  DFF \creg_reg[56]  ( .D(n7129), .CLK(clk), .RST(rst), .Q(creg[56]) );
  DFF \creg_reg[57]  ( .D(n7128), .CLK(clk), .RST(rst), .Q(creg[57]) );
  DFF \creg_reg[58]  ( .D(n7127), .CLK(clk), .RST(rst), .Q(creg[58]) );
  DFF \creg_reg[59]  ( .D(n7126), .CLK(clk), .RST(rst), .Q(creg[59]) );
  DFF \creg_reg[60]  ( .D(n7125), .CLK(clk), .RST(rst), .Q(creg[60]) );
  DFF \creg_reg[61]  ( .D(n7124), .CLK(clk), .RST(rst), .Q(creg[61]) );
  DFF \creg_reg[62]  ( .D(n7123), .CLK(clk), .RST(rst), .Q(creg[62]) );
  DFF \creg_reg[63]  ( .D(n7122), .CLK(clk), .RST(rst), .Q(creg[63]) );
  DFF \creg_reg[64]  ( .D(n7121), .CLK(clk), .RST(rst), .Q(creg[64]) );
  DFF \creg_reg[65]  ( .D(n7120), .CLK(clk), .RST(rst), .Q(creg[65]) );
  DFF \creg_reg[66]  ( .D(n7119), .CLK(clk), .RST(rst), .Q(creg[66]) );
  DFF \creg_reg[67]  ( .D(n7118), .CLK(clk), .RST(rst), .Q(creg[67]) );
  DFF \creg_reg[68]  ( .D(n7117), .CLK(clk), .RST(rst), .Q(creg[68]) );
  DFF \creg_reg[69]  ( .D(n7116), .CLK(clk), .RST(rst), .Q(creg[69]) );
  DFF \creg_reg[70]  ( .D(n7115), .CLK(clk), .RST(rst), .Q(creg[70]) );
  DFF \creg_reg[71]  ( .D(n7114), .CLK(clk), .RST(rst), .Q(creg[71]) );
  DFF \creg_reg[72]  ( .D(n7113), .CLK(clk), .RST(rst), .Q(creg[72]) );
  DFF \creg_reg[73]  ( .D(n7112), .CLK(clk), .RST(rst), .Q(creg[73]) );
  DFF \creg_reg[74]  ( .D(n7111), .CLK(clk), .RST(rst), .Q(creg[74]) );
  DFF \creg_reg[75]  ( .D(n7110), .CLK(clk), .RST(rst), .Q(creg[75]) );
  DFF \creg_reg[76]  ( .D(n7109), .CLK(clk), .RST(rst), .Q(creg[76]) );
  DFF \creg_reg[77]  ( .D(n7108), .CLK(clk), .RST(rst), .Q(creg[77]) );
  DFF \creg_reg[78]  ( .D(n7107), .CLK(clk), .RST(rst), .Q(creg[78]) );
  DFF \creg_reg[79]  ( .D(n7106), .CLK(clk), .RST(rst), .Q(creg[79]) );
  DFF \creg_reg[80]  ( .D(n7105), .CLK(clk), .RST(rst), .Q(creg[80]) );
  DFF \creg_reg[81]  ( .D(n7104), .CLK(clk), .RST(rst), .Q(creg[81]) );
  DFF \creg_reg[82]  ( .D(n7103), .CLK(clk), .RST(rst), .Q(creg[82]) );
  DFF \creg_reg[83]  ( .D(n7102), .CLK(clk), .RST(rst), .Q(creg[83]) );
  DFF \creg_reg[84]  ( .D(n7101), .CLK(clk), .RST(rst), .Q(creg[84]) );
  DFF \creg_reg[85]  ( .D(n7100), .CLK(clk), .RST(rst), .Q(creg[85]) );
  DFF \creg_reg[86]  ( .D(n7099), .CLK(clk), .RST(rst), .Q(creg[86]) );
  DFF \creg_reg[87]  ( .D(n7098), .CLK(clk), .RST(rst), .Q(creg[87]) );
  DFF \creg_reg[88]  ( .D(n7097), .CLK(clk), .RST(rst), .Q(creg[88]) );
  DFF \creg_reg[89]  ( .D(n7096), .CLK(clk), .RST(rst), .Q(creg[89]) );
  DFF \creg_reg[90]  ( .D(n7095), .CLK(clk), .RST(rst), .Q(creg[90]) );
  DFF \creg_reg[91]  ( .D(n7094), .CLK(clk), .RST(rst), .Q(creg[91]) );
  DFF \creg_reg[92]  ( .D(n7093), .CLK(clk), .RST(rst), .Q(creg[92]) );
  DFF \creg_reg[93]  ( .D(n7092), .CLK(clk), .RST(rst), .Q(creg[93]) );
  DFF \creg_reg[94]  ( .D(n7091), .CLK(clk), .RST(rst), .Q(creg[94]) );
  DFF \creg_reg[95]  ( .D(n7090), .CLK(clk), .RST(rst), .Q(creg[95]) );
  DFF \creg_reg[96]  ( .D(n7089), .CLK(clk), .RST(rst), .Q(creg[96]) );
  DFF \creg_reg[97]  ( .D(n7088), .CLK(clk), .RST(rst), .Q(creg[97]) );
  DFF \creg_reg[98]  ( .D(n7087), .CLK(clk), .RST(rst), .Q(creg[98]) );
  DFF \creg_reg[99]  ( .D(n7086), .CLK(clk), .RST(rst), .Q(creg[99]) );
  DFF \creg_reg[100]  ( .D(n7085), .CLK(clk), .RST(rst), .Q(creg[100]) );
  DFF \creg_reg[101]  ( .D(n7084), .CLK(clk), .RST(rst), .Q(creg[101]) );
  DFF \creg_reg[102]  ( .D(n7083), .CLK(clk), .RST(rst), .Q(creg[102]) );
  DFF \creg_reg[103]  ( .D(n7082), .CLK(clk), .RST(rst), .Q(creg[103]) );
  DFF \creg_reg[104]  ( .D(n7081), .CLK(clk), .RST(rst), .Q(creg[104]) );
  DFF \creg_reg[105]  ( .D(n7080), .CLK(clk), .RST(rst), .Q(creg[105]) );
  DFF \creg_reg[106]  ( .D(n7079), .CLK(clk), .RST(rst), .Q(creg[106]) );
  DFF \creg_reg[107]  ( .D(n7078), .CLK(clk), .RST(rst), .Q(creg[107]) );
  DFF \creg_reg[108]  ( .D(n7077), .CLK(clk), .RST(rst), .Q(creg[108]) );
  DFF \creg_reg[109]  ( .D(n7076), .CLK(clk), .RST(rst), .Q(creg[109]) );
  DFF \creg_reg[110]  ( .D(n7075), .CLK(clk), .RST(rst), .Q(creg[110]) );
  DFF \creg_reg[111]  ( .D(n7074), .CLK(clk), .RST(rst), .Q(creg[111]) );
  DFF \creg_reg[112]  ( .D(n7073), .CLK(clk), .RST(rst), .Q(creg[112]) );
  DFF \creg_reg[113]  ( .D(n7072), .CLK(clk), .RST(rst), .Q(creg[113]) );
  DFF \creg_reg[114]  ( .D(n7071), .CLK(clk), .RST(rst), .Q(creg[114]) );
  DFF \creg_reg[115]  ( .D(n7070), .CLK(clk), .RST(rst), .Q(creg[115]) );
  DFF \creg_reg[116]  ( .D(n7069), .CLK(clk), .RST(rst), .Q(creg[116]) );
  DFF \creg_reg[117]  ( .D(n7068), .CLK(clk), .RST(rst), .Q(creg[117]) );
  DFF \creg_reg[118]  ( .D(n7067), .CLK(clk), .RST(rst), .Q(creg[118]) );
  DFF \creg_reg[119]  ( .D(n7066), .CLK(clk), .RST(rst), .Q(creg[119]) );
  DFF \creg_reg[120]  ( .D(n7065), .CLK(clk), .RST(rst), .Q(creg[120]) );
  DFF \creg_reg[121]  ( .D(n7064), .CLK(clk), .RST(rst), .Q(creg[121]) );
  DFF \creg_reg[122]  ( .D(n7063), .CLK(clk), .RST(rst), .Q(creg[122]) );
  DFF \creg_reg[123]  ( .D(n7062), .CLK(clk), .RST(rst), .Q(creg[123]) );
  DFF \creg_reg[124]  ( .D(n7061), .CLK(clk), .RST(rst), .Q(creg[124]) );
  DFF \creg_reg[125]  ( .D(n7060), .CLK(clk), .RST(rst), .Q(creg[125]) );
  DFF \creg_reg[126]  ( .D(n7059), .CLK(clk), .RST(rst), .Q(creg[126]) );
  DFF \creg_reg[127]  ( .D(n7058), .CLK(clk), .RST(rst), .Q(creg[127]) );
  DFF \creg_reg[128]  ( .D(n7057), .CLK(clk), .RST(rst), .Q(creg[128]) );
  DFF \creg_reg[129]  ( .D(n7056), .CLK(clk), .RST(rst), .Q(creg[129]) );
  DFF \creg_reg[130]  ( .D(n7055), .CLK(clk), .RST(rst), .Q(creg[130]) );
  DFF \creg_reg[131]  ( .D(n7054), .CLK(clk), .RST(rst), .Q(creg[131]) );
  DFF \creg_reg[132]  ( .D(n7053), .CLK(clk), .RST(rst), .Q(creg[132]) );
  DFF \creg_reg[133]  ( .D(n7052), .CLK(clk), .RST(rst), .Q(creg[133]) );
  DFF \creg_reg[134]  ( .D(n7051), .CLK(clk), .RST(rst), .Q(creg[134]) );
  DFF \creg_reg[135]  ( .D(n7050), .CLK(clk), .RST(rst), .Q(creg[135]) );
  DFF \creg_reg[136]  ( .D(n7049), .CLK(clk), .RST(rst), .Q(creg[136]) );
  DFF \creg_reg[137]  ( .D(n7048), .CLK(clk), .RST(rst), .Q(creg[137]) );
  DFF \creg_reg[138]  ( .D(n7047), .CLK(clk), .RST(rst), .Q(creg[138]) );
  DFF \creg_reg[139]  ( .D(n7046), .CLK(clk), .RST(rst), .Q(creg[139]) );
  DFF \creg_reg[140]  ( .D(n7045), .CLK(clk), .RST(rst), .Q(creg[140]) );
  DFF \creg_reg[141]  ( .D(n7044), .CLK(clk), .RST(rst), .Q(creg[141]) );
  DFF \creg_reg[142]  ( .D(n7043), .CLK(clk), .RST(rst), .Q(creg[142]) );
  DFF \creg_reg[143]  ( .D(n7042), .CLK(clk), .RST(rst), .Q(creg[143]) );
  DFF \creg_reg[144]  ( .D(n7041), .CLK(clk), .RST(rst), .Q(creg[144]) );
  DFF \creg_reg[145]  ( .D(n7040), .CLK(clk), .RST(rst), .Q(creg[145]) );
  DFF \creg_reg[146]  ( .D(n7039), .CLK(clk), .RST(rst), .Q(creg[146]) );
  DFF \creg_reg[147]  ( .D(n7038), .CLK(clk), .RST(rst), .Q(creg[147]) );
  DFF \creg_reg[148]  ( .D(n7037), .CLK(clk), .RST(rst), .Q(creg[148]) );
  DFF \creg_reg[149]  ( .D(n7036), .CLK(clk), .RST(rst), .Q(creg[149]) );
  DFF \creg_reg[150]  ( .D(n7035), .CLK(clk), .RST(rst), .Q(creg[150]) );
  DFF \creg_reg[151]  ( .D(n7034), .CLK(clk), .RST(rst), .Q(creg[151]) );
  DFF \creg_reg[152]  ( .D(n7033), .CLK(clk), .RST(rst), .Q(creg[152]) );
  DFF \creg_reg[153]  ( .D(n7032), .CLK(clk), .RST(rst), .Q(creg[153]) );
  DFF \creg_reg[154]  ( .D(n7031), .CLK(clk), .RST(rst), .Q(creg[154]) );
  DFF \creg_reg[155]  ( .D(n7030), .CLK(clk), .RST(rst), .Q(creg[155]) );
  DFF \creg_reg[156]  ( .D(n7029), .CLK(clk), .RST(rst), .Q(creg[156]) );
  DFF \creg_reg[157]  ( .D(n7028), .CLK(clk), .RST(rst), .Q(creg[157]) );
  DFF \creg_reg[158]  ( .D(n7027), .CLK(clk), .RST(rst), .Q(creg[158]) );
  DFF \creg_reg[159]  ( .D(n7026), .CLK(clk), .RST(rst), .Q(creg[159]) );
  DFF \creg_reg[160]  ( .D(n7025), .CLK(clk), .RST(rst), .Q(creg[160]) );
  DFF \creg_reg[161]  ( .D(n7024), .CLK(clk), .RST(rst), .Q(creg[161]) );
  DFF \creg_reg[162]  ( .D(n7023), .CLK(clk), .RST(rst), .Q(creg[162]) );
  DFF \creg_reg[163]  ( .D(n7022), .CLK(clk), .RST(rst), .Q(creg[163]) );
  DFF \creg_reg[164]  ( .D(n7021), .CLK(clk), .RST(rst), .Q(creg[164]) );
  DFF \creg_reg[165]  ( .D(n7020), .CLK(clk), .RST(rst), .Q(creg[165]) );
  DFF \creg_reg[166]  ( .D(n7019), .CLK(clk), .RST(rst), .Q(creg[166]) );
  DFF \creg_reg[167]  ( .D(n7018), .CLK(clk), .RST(rst), .Q(creg[167]) );
  DFF \creg_reg[168]  ( .D(n7017), .CLK(clk), .RST(rst), .Q(creg[168]) );
  DFF \creg_reg[169]  ( .D(n7016), .CLK(clk), .RST(rst), .Q(creg[169]) );
  DFF \creg_reg[170]  ( .D(n7015), .CLK(clk), .RST(rst), .Q(creg[170]) );
  DFF \creg_reg[171]  ( .D(n7014), .CLK(clk), .RST(rst), .Q(creg[171]) );
  DFF \creg_reg[172]  ( .D(n7013), .CLK(clk), .RST(rst), .Q(creg[172]) );
  DFF \creg_reg[173]  ( .D(n7012), .CLK(clk), .RST(rst), .Q(creg[173]) );
  DFF \creg_reg[174]  ( .D(n7011), .CLK(clk), .RST(rst), .Q(creg[174]) );
  DFF \creg_reg[175]  ( .D(n7010), .CLK(clk), .RST(rst), .Q(creg[175]) );
  DFF \creg_reg[176]  ( .D(n7009), .CLK(clk), .RST(rst), .Q(creg[176]) );
  DFF \creg_reg[177]  ( .D(n7008), .CLK(clk), .RST(rst), .Q(creg[177]) );
  DFF \creg_reg[178]  ( .D(n7007), .CLK(clk), .RST(rst), .Q(creg[178]) );
  DFF \creg_reg[179]  ( .D(n7006), .CLK(clk), .RST(rst), .Q(creg[179]) );
  DFF \creg_reg[180]  ( .D(n7005), .CLK(clk), .RST(rst), .Q(creg[180]) );
  DFF \creg_reg[181]  ( .D(n7004), .CLK(clk), .RST(rst), .Q(creg[181]) );
  DFF \creg_reg[182]  ( .D(n7003), .CLK(clk), .RST(rst), .Q(creg[182]) );
  DFF \creg_reg[183]  ( .D(n7002), .CLK(clk), .RST(rst), .Q(creg[183]) );
  DFF \creg_reg[184]  ( .D(n7001), .CLK(clk), .RST(rst), .Q(creg[184]) );
  DFF \creg_reg[185]  ( .D(n7000), .CLK(clk), .RST(rst), .Q(creg[185]) );
  DFF \creg_reg[186]  ( .D(n6999), .CLK(clk), .RST(rst), .Q(creg[186]) );
  DFF \creg_reg[187]  ( .D(n6998), .CLK(clk), .RST(rst), .Q(creg[187]) );
  DFF \creg_reg[188]  ( .D(n6997), .CLK(clk), .RST(rst), .Q(creg[188]) );
  DFF \creg_reg[189]  ( .D(n6996), .CLK(clk), .RST(rst), .Q(creg[189]) );
  DFF \creg_reg[190]  ( .D(n6995), .CLK(clk), .RST(rst), .Q(creg[190]) );
  DFF \creg_reg[191]  ( .D(n6994), .CLK(clk), .RST(rst), .Q(creg[191]) );
  DFF \creg_reg[192]  ( .D(n6993), .CLK(clk), .RST(rst), .Q(creg[192]) );
  DFF \creg_reg[193]  ( .D(n6992), .CLK(clk), .RST(rst), .Q(creg[193]) );
  DFF \creg_reg[194]  ( .D(n6991), .CLK(clk), .RST(rst), .Q(creg[194]) );
  DFF \creg_reg[195]  ( .D(n6990), .CLK(clk), .RST(rst), .Q(creg[195]) );
  DFF \creg_reg[196]  ( .D(n6989), .CLK(clk), .RST(rst), .Q(creg[196]) );
  DFF \creg_reg[197]  ( .D(n6988), .CLK(clk), .RST(rst), .Q(creg[197]) );
  DFF \creg_reg[198]  ( .D(n6987), .CLK(clk), .RST(rst), .Q(creg[198]) );
  DFF \creg_reg[199]  ( .D(n6986), .CLK(clk), .RST(rst), .Q(creg[199]) );
  DFF \creg_reg[200]  ( .D(n6985), .CLK(clk), .RST(rst), .Q(creg[200]) );
  DFF \creg_reg[201]  ( .D(n6984), .CLK(clk), .RST(rst), .Q(creg[201]) );
  DFF \creg_reg[202]  ( .D(n6983), .CLK(clk), .RST(rst), .Q(creg[202]) );
  DFF \creg_reg[203]  ( .D(n6982), .CLK(clk), .RST(rst), .Q(creg[203]) );
  DFF \creg_reg[204]  ( .D(n6981), .CLK(clk), .RST(rst), .Q(creg[204]) );
  DFF \creg_reg[205]  ( .D(n6980), .CLK(clk), .RST(rst), .Q(creg[205]) );
  DFF \creg_reg[206]  ( .D(n6979), .CLK(clk), .RST(rst), .Q(creg[206]) );
  DFF \creg_reg[207]  ( .D(n6978), .CLK(clk), .RST(rst), .Q(creg[207]) );
  DFF \creg_reg[208]  ( .D(n6977), .CLK(clk), .RST(rst), .Q(creg[208]) );
  DFF \creg_reg[209]  ( .D(n6976), .CLK(clk), .RST(rst), .Q(creg[209]) );
  DFF \creg_reg[210]  ( .D(n6975), .CLK(clk), .RST(rst), .Q(creg[210]) );
  DFF \creg_reg[211]  ( .D(n6974), .CLK(clk), .RST(rst), .Q(creg[211]) );
  DFF \creg_reg[212]  ( .D(n6973), .CLK(clk), .RST(rst), .Q(creg[212]) );
  DFF \creg_reg[213]  ( .D(n6972), .CLK(clk), .RST(rst), .Q(creg[213]) );
  DFF \creg_reg[214]  ( .D(n6971), .CLK(clk), .RST(rst), .Q(creg[214]) );
  DFF \creg_reg[215]  ( .D(n6970), .CLK(clk), .RST(rst), .Q(creg[215]) );
  DFF \creg_reg[216]  ( .D(n6969), .CLK(clk), .RST(rst), .Q(creg[216]) );
  DFF \creg_reg[217]  ( .D(n6968), .CLK(clk), .RST(rst), .Q(creg[217]) );
  DFF \creg_reg[218]  ( .D(n6967), .CLK(clk), .RST(rst), .Q(creg[218]) );
  DFF \creg_reg[219]  ( .D(n6966), .CLK(clk), .RST(rst), .Q(creg[219]) );
  DFF \creg_reg[220]  ( .D(n6965), .CLK(clk), .RST(rst), .Q(creg[220]) );
  DFF \creg_reg[221]  ( .D(n6964), .CLK(clk), .RST(rst), .Q(creg[221]) );
  DFF \creg_reg[222]  ( .D(n6963), .CLK(clk), .RST(rst), .Q(creg[222]) );
  DFF \creg_reg[223]  ( .D(n6962), .CLK(clk), .RST(rst), .Q(creg[223]) );
  DFF \creg_reg[224]  ( .D(n6961), .CLK(clk), .RST(rst), .Q(creg[224]) );
  DFF \creg_reg[225]  ( .D(n6960), .CLK(clk), .RST(rst), .Q(creg[225]) );
  DFF \creg_reg[226]  ( .D(n6959), .CLK(clk), .RST(rst), .Q(creg[226]) );
  DFF \creg_reg[227]  ( .D(n6958), .CLK(clk), .RST(rst), .Q(creg[227]) );
  DFF \creg_reg[228]  ( .D(n6957), .CLK(clk), .RST(rst), .Q(creg[228]) );
  DFF \creg_reg[229]  ( .D(n6956), .CLK(clk), .RST(rst), .Q(creg[229]) );
  DFF \creg_reg[230]  ( .D(n6955), .CLK(clk), .RST(rst), .Q(creg[230]) );
  DFF \creg_reg[231]  ( .D(n6954), .CLK(clk), .RST(rst), .Q(creg[231]) );
  DFF \creg_reg[232]  ( .D(n6953), .CLK(clk), .RST(rst), .Q(creg[232]) );
  DFF \creg_reg[233]  ( .D(n6952), .CLK(clk), .RST(rst), .Q(creg[233]) );
  DFF \creg_reg[234]  ( .D(n6951), .CLK(clk), .RST(rst), .Q(creg[234]) );
  DFF \creg_reg[235]  ( .D(n6950), .CLK(clk), .RST(rst), .Q(creg[235]) );
  DFF \creg_reg[236]  ( .D(n6949), .CLK(clk), .RST(rst), .Q(creg[236]) );
  DFF \creg_reg[237]  ( .D(n6948), .CLK(clk), .RST(rst), .Q(creg[237]) );
  DFF \creg_reg[238]  ( .D(n6947), .CLK(clk), .RST(rst), .Q(creg[238]) );
  DFF \creg_reg[239]  ( .D(n6946), .CLK(clk), .RST(rst), .Q(creg[239]) );
  DFF \creg_reg[240]  ( .D(n6945), .CLK(clk), .RST(rst), .Q(creg[240]) );
  DFF \creg_reg[241]  ( .D(n6944), .CLK(clk), .RST(rst), .Q(creg[241]) );
  DFF \creg_reg[242]  ( .D(n6943), .CLK(clk), .RST(rst), .Q(creg[242]) );
  DFF \creg_reg[243]  ( .D(n6942), .CLK(clk), .RST(rst), .Q(creg[243]) );
  DFF \creg_reg[244]  ( .D(n6941), .CLK(clk), .RST(rst), .Q(creg[244]) );
  DFF \creg_reg[245]  ( .D(n6940), .CLK(clk), .RST(rst), .Q(creg[245]) );
  DFF \creg_reg[246]  ( .D(n6939), .CLK(clk), .RST(rst), .Q(creg[246]) );
  DFF \creg_reg[247]  ( .D(n6938), .CLK(clk), .RST(rst), .Q(creg[247]) );
  DFF \creg_reg[248]  ( .D(n6937), .CLK(clk), .RST(rst), .Q(creg[248]) );
  DFF \creg_reg[249]  ( .D(n6936), .CLK(clk), .RST(rst), .Q(creg[249]) );
  DFF \creg_reg[250]  ( .D(n6935), .CLK(clk), .RST(rst), .Q(creg[250]) );
  DFF \creg_reg[251]  ( .D(n6934), .CLK(clk), .RST(rst), .Q(creg[251]) );
  DFF \creg_reg[252]  ( .D(n6933), .CLK(clk), .RST(rst), .Q(creg[252]) );
  DFF \creg_reg[253]  ( .D(n6932), .CLK(clk), .RST(rst), .Q(creg[253]) );
  DFF \creg_reg[254]  ( .D(n6931), .CLK(clk), .RST(rst), .Q(creg[254]) );
  DFF \creg_reg[255]  ( .D(n6930), .CLK(clk), .RST(rst), .Q(creg[255]) );
  DFF \creg_reg[256]  ( .D(n6929), .CLK(clk), .RST(rst), .Q(creg[256]) );
  DFF \creg_reg[257]  ( .D(n6928), .CLK(clk), .RST(rst), .Q(creg[257]) );
  DFF \creg_reg[258]  ( .D(n6927), .CLK(clk), .RST(rst), .Q(creg[258]) );
  DFF \creg_reg[259]  ( .D(n6926), .CLK(clk), .RST(rst), .Q(creg[259]) );
  DFF \creg_reg[260]  ( .D(n6925), .CLK(clk), .RST(rst), .Q(creg[260]) );
  DFF \creg_reg[261]  ( .D(n6924), .CLK(clk), .RST(rst), .Q(creg[261]) );
  DFF \creg_reg[262]  ( .D(n6923), .CLK(clk), .RST(rst), .Q(creg[262]) );
  DFF \creg_reg[263]  ( .D(n6922), .CLK(clk), .RST(rst), .Q(creg[263]) );
  DFF \creg_reg[264]  ( .D(n6921), .CLK(clk), .RST(rst), .Q(creg[264]) );
  DFF \creg_reg[265]  ( .D(n6920), .CLK(clk), .RST(rst), .Q(creg[265]) );
  DFF \creg_reg[266]  ( .D(n6919), .CLK(clk), .RST(rst), .Q(creg[266]) );
  DFF \creg_reg[267]  ( .D(n6918), .CLK(clk), .RST(rst), .Q(creg[267]) );
  DFF \creg_reg[268]  ( .D(n6917), .CLK(clk), .RST(rst), .Q(creg[268]) );
  DFF \creg_reg[269]  ( .D(n6916), .CLK(clk), .RST(rst), .Q(creg[269]) );
  DFF \creg_reg[270]  ( .D(n6915), .CLK(clk), .RST(rst), .Q(creg[270]) );
  DFF \creg_reg[271]  ( .D(n6914), .CLK(clk), .RST(rst), .Q(creg[271]) );
  DFF \creg_reg[272]  ( .D(n6913), .CLK(clk), .RST(rst), .Q(creg[272]) );
  DFF \creg_reg[273]  ( .D(n6912), .CLK(clk), .RST(rst), .Q(creg[273]) );
  DFF \creg_reg[274]  ( .D(n6911), .CLK(clk), .RST(rst), .Q(creg[274]) );
  DFF \creg_reg[275]  ( .D(n6910), .CLK(clk), .RST(rst), .Q(creg[275]) );
  DFF \creg_reg[276]  ( .D(n6909), .CLK(clk), .RST(rst), .Q(creg[276]) );
  DFF \creg_reg[277]  ( .D(n6908), .CLK(clk), .RST(rst), .Q(creg[277]) );
  DFF \creg_reg[278]  ( .D(n6907), .CLK(clk), .RST(rst), .Q(creg[278]) );
  DFF \creg_reg[279]  ( .D(n6906), .CLK(clk), .RST(rst), .Q(creg[279]) );
  DFF \creg_reg[280]  ( .D(n6905), .CLK(clk), .RST(rst), .Q(creg[280]) );
  DFF \creg_reg[281]  ( .D(n6904), .CLK(clk), .RST(rst), .Q(creg[281]) );
  DFF \creg_reg[282]  ( .D(n6903), .CLK(clk), .RST(rst), .Q(creg[282]) );
  DFF \creg_reg[283]  ( .D(n6902), .CLK(clk), .RST(rst), .Q(creg[283]) );
  DFF \creg_reg[284]  ( .D(n6901), .CLK(clk), .RST(rst), .Q(creg[284]) );
  DFF \creg_reg[285]  ( .D(n6900), .CLK(clk), .RST(rst), .Q(creg[285]) );
  DFF \creg_reg[286]  ( .D(n6899), .CLK(clk), .RST(rst), .Q(creg[286]) );
  DFF \creg_reg[287]  ( .D(n6898), .CLK(clk), .RST(rst), .Q(creg[287]) );
  DFF \creg_reg[288]  ( .D(n6897), .CLK(clk), .RST(rst), .Q(creg[288]) );
  DFF \creg_reg[289]  ( .D(n6896), .CLK(clk), .RST(rst), .Q(creg[289]) );
  DFF \creg_reg[290]  ( .D(n6895), .CLK(clk), .RST(rst), .Q(creg[290]) );
  DFF \creg_reg[291]  ( .D(n6894), .CLK(clk), .RST(rst), .Q(creg[291]) );
  DFF \creg_reg[292]  ( .D(n6893), .CLK(clk), .RST(rst), .Q(creg[292]) );
  DFF \creg_reg[293]  ( .D(n6892), .CLK(clk), .RST(rst), .Q(creg[293]) );
  DFF \creg_reg[294]  ( .D(n6891), .CLK(clk), .RST(rst), .Q(creg[294]) );
  DFF \creg_reg[295]  ( .D(n6890), .CLK(clk), .RST(rst), .Q(creg[295]) );
  DFF \creg_reg[296]  ( .D(n6889), .CLK(clk), .RST(rst), .Q(creg[296]) );
  DFF \creg_reg[297]  ( .D(n6888), .CLK(clk), .RST(rst), .Q(creg[297]) );
  DFF \creg_reg[298]  ( .D(n6887), .CLK(clk), .RST(rst), .Q(creg[298]) );
  DFF \creg_reg[299]  ( .D(n6886), .CLK(clk), .RST(rst), .Q(creg[299]) );
  DFF \creg_reg[300]  ( .D(n6885), .CLK(clk), .RST(rst), .Q(creg[300]) );
  DFF \creg_reg[301]  ( .D(n6884), .CLK(clk), .RST(rst), .Q(creg[301]) );
  DFF \creg_reg[302]  ( .D(n6883), .CLK(clk), .RST(rst), .Q(creg[302]) );
  DFF \creg_reg[303]  ( .D(n6882), .CLK(clk), .RST(rst), .Q(creg[303]) );
  DFF \creg_reg[304]  ( .D(n6881), .CLK(clk), .RST(rst), .Q(creg[304]) );
  DFF \creg_reg[305]  ( .D(n6880), .CLK(clk), .RST(rst), .Q(creg[305]) );
  DFF \creg_reg[306]  ( .D(n6879), .CLK(clk), .RST(rst), .Q(creg[306]) );
  DFF \creg_reg[307]  ( .D(n6878), .CLK(clk), .RST(rst), .Q(creg[307]) );
  DFF \creg_reg[308]  ( .D(n6877), .CLK(clk), .RST(rst), .Q(creg[308]) );
  DFF \creg_reg[309]  ( .D(n6876), .CLK(clk), .RST(rst), .Q(creg[309]) );
  DFF \creg_reg[310]  ( .D(n6875), .CLK(clk), .RST(rst), .Q(creg[310]) );
  DFF \creg_reg[311]  ( .D(n6874), .CLK(clk), .RST(rst), .Q(creg[311]) );
  DFF \creg_reg[312]  ( .D(n6873), .CLK(clk), .RST(rst), .Q(creg[312]) );
  DFF \creg_reg[313]  ( .D(n6872), .CLK(clk), .RST(rst), .Q(creg[313]) );
  DFF \creg_reg[314]  ( .D(n6871), .CLK(clk), .RST(rst), .Q(creg[314]) );
  DFF \creg_reg[315]  ( .D(n6870), .CLK(clk), .RST(rst), .Q(creg[315]) );
  DFF \creg_reg[316]  ( .D(n6869), .CLK(clk), .RST(rst), .Q(creg[316]) );
  DFF \creg_reg[317]  ( .D(n6868), .CLK(clk), .RST(rst), .Q(creg[317]) );
  DFF \creg_reg[318]  ( .D(n6867), .CLK(clk), .RST(rst), .Q(creg[318]) );
  DFF \creg_reg[319]  ( .D(n6866), .CLK(clk), .RST(rst), .Q(creg[319]) );
  DFF \creg_reg[320]  ( .D(n6865), .CLK(clk), .RST(rst), .Q(creg[320]) );
  DFF \creg_reg[321]  ( .D(n6864), .CLK(clk), .RST(rst), .Q(creg[321]) );
  DFF \creg_reg[322]  ( .D(n6863), .CLK(clk), .RST(rst), .Q(creg[322]) );
  DFF \creg_reg[323]  ( .D(n6862), .CLK(clk), .RST(rst), .Q(creg[323]) );
  DFF \creg_reg[324]  ( .D(n6861), .CLK(clk), .RST(rst), .Q(creg[324]) );
  DFF \creg_reg[325]  ( .D(n6860), .CLK(clk), .RST(rst), .Q(creg[325]) );
  DFF \creg_reg[326]  ( .D(n6859), .CLK(clk), .RST(rst), .Q(creg[326]) );
  DFF \creg_reg[327]  ( .D(n6858), .CLK(clk), .RST(rst), .Q(creg[327]) );
  DFF \creg_reg[328]  ( .D(n6857), .CLK(clk), .RST(rst), .Q(creg[328]) );
  DFF \creg_reg[329]  ( .D(n6856), .CLK(clk), .RST(rst), .Q(creg[329]) );
  DFF \creg_reg[330]  ( .D(n6855), .CLK(clk), .RST(rst), .Q(creg[330]) );
  DFF \creg_reg[331]  ( .D(n6854), .CLK(clk), .RST(rst), .Q(creg[331]) );
  DFF \creg_reg[332]  ( .D(n6853), .CLK(clk), .RST(rst), .Q(creg[332]) );
  DFF \creg_reg[333]  ( .D(n6852), .CLK(clk), .RST(rst), .Q(creg[333]) );
  DFF \creg_reg[334]  ( .D(n6851), .CLK(clk), .RST(rst), .Q(creg[334]) );
  DFF \creg_reg[335]  ( .D(n6850), .CLK(clk), .RST(rst), .Q(creg[335]) );
  DFF \creg_reg[336]  ( .D(n6849), .CLK(clk), .RST(rst), .Q(creg[336]) );
  DFF \creg_reg[337]  ( .D(n6848), .CLK(clk), .RST(rst), .Q(creg[337]) );
  DFF \creg_reg[338]  ( .D(n6847), .CLK(clk), .RST(rst), .Q(creg[338]) );
  DFF \creg_reg[339]  ( .D(n6846), .CLK(clk), .RST(rst), .Q(creg[339]) );
  DFF \creg_reg[340]  ( .D(n6845), .CLK(clk), .RST(rst), .Q(creg[340]) );
  DFF \creg_reg[341]  ( .D(n6844), .CLK(clk), .RST(rst), .Q(creg[341]) );
  DFF \creg_reg[342]  ( .D(n6843), .CLK(clk), .RST(rst), .Q(creg[342]) );
  DFF \creg_reg[343]  ( .D(n6842), .CLK(clk), .RST(rst), .Q(creg[343]) );
  DFF \creg_reg[344]  ( .D(n6841), .CLK(clk), .RST(rst), .Q(creg[344]) );
  DFF \creg_reg[345]  ( .D(n6840), .CLK(clk), .RST(rst), .Q(creg[345]) );
  DFF \creg_reg[346]  ( .D(n6839), .CLK(clk), .RST(rst), .Q(creg[346]) );
  DFF \creg_reg[347]  ( .D(n6838), .CLK(clk), .RST(rst), .Q(creg[347]) );
  DFF \creg_reg[348]  ( .D(n6837), .CLK(clk), .RST(rst), .Q(creg[348]) );
  DFF \creg_reg[349]  ( .D(n6836), .CLK(clk), .RST(rst), .Q(creg[349]) );
  DFF \creg_reg[350]  ( .D(n6835), .CLK(clk), .RST(rst), .Q(creg[350]) );
  DFF \creg_reg[351]  ( .D(n6834), .CLK(clk), .RST(rst), .Q(creg[351]) );
  DFF \creg_reg[352]  ( .D(n6833), .CLK(clk), .RST(rst), .Q(creg[352]) );
  DFF \creg_reg[353]  ( .D(n6832), .CLK(clk), .RST(rst), .Q(creg[353]) );
  DFF \creg_reg[354]  ( .D(n6831), .CLK(clk), .RST(rst), .Q(creg[354]) );
  DFF \creg_reg[355]  ( .D(n6830), .CLK(clk), .RST(rst), .Q(creg[355]) );
  DFF \creg_reg[356]  ( .D(n6829), .CLK(clk), .RST(rst), .Q(creg[356]) );
  DFF \creg_reg[357]  ( .D(n6828), .CLK(clk), .RST(rst), .Q(creg[357]) );
  DFF \creg_reg[358]  ( .D(n6827), .CLK(clk), .RST(rst), .Q(creg[358]) );
  DFF \creg_reg[359]  ( .D(n6826), .CLK(clk), .RST(rst), .Q(creg[359]) );
  DFF \creg_reg[360]  ( .D(n6825), .CLK(clk), .RST(rst), .Q(creg[360]) );
  DFF \creg_reg[361]  ( .D(n6824), .CLK(clk), .RST(rst), .Q(creg[361]) );
  DFF \creg_reg[362]  ( .D(n6823), .CLK(clk), .RST(rst), .Q(creg[362]) );
  DFF \creg_reg[363]  ( .D(n6822), .CLK(clk), .RST(rst), .Q(creg[363]) );
  DFF \creg_reg[364]  ( .D(n6821), .CLK(clk), .RST(rst), .Q(creg[364]) );
  DFF \creg_reg[365]  ( .D(n6820), .CLK(clk), .RST(rst), .Q(creg[365]) );
  DFF \creg_reg[366]  ( .D(n6819), .CLK(clk), .RST(rst), .Q(creg[366]) );
  DFF \creg_reg[367]  ( .D(n6818), .CLK(clk), .RST(rst), .Q(creg[367]) );
  DFF \creg_reg[368]  ( .D(n6817), .CLK(clk), .RST(rst), .Q(creg[368]) );
  DFF \creg_reg[369]  ( .D(n6816), .CLK(clk), .RST(rst), .Q(creg[369]) );
  DFF \creg_reg[370]  ( .D(n6815), .CLK(clk), .RST(rst), .Q(creg[370]) );
  DFF \creg_reg[371]  ( .D(n6814), .CLK(clk), .RST(rst), .Q(creg[371]) );
  DFF \creg_reg[372]  ( .D(n6813), .CLK(clk), .RST(rst), .Q(creg[372]) );
  DFF \creg_reg[373]  ( .D(n6812), .CLK(clk), .RST(rst), .Q(creg[373]) );
  DFF \creg_reg[374]  ( .D(n6811), .CLK(clk), .RST(rst), .Q(creg[374]) );
  DFF \creg_reg[375]  ( .D(n6810), .CLK(clk), .RST(rst), .Q(creg[375]) );
  DFF \creg_reg[376]  ( .D(n6809), .CLK(clk), .RST(rst), .Q(creg[376]) );
  DFF \creg_reg[377]  ( .D(n6808), .CLK(clk), .RST(rst), .Q(creg[377]) );
  DFF \creg_reg[378]  ( .D(n6807), .CLK(clk), .RST(rst), .Q(creg[378]) );
  DFF \creg_reg[379]  ( .D(n6806), .CLK(clk), .RST(rst), .Q(creg[379]) );
  DFF \creg_reg[380]  ( .D(n6805), .CLK(clk), .RST(rst), .Q(creg[380]) );
  DFF \creg_reg[381]  ( .D(n6804), .CLK(clk), .RST(rst), .Q(creg[381]) );
  DFF \creg_reg[382]  ( .D(n6803), .CLK(clk), .RST(rst), .Q(creg[382]) );
  DFF \creg_reg[383]  ( .D(n6802), .CLK(clk), .RST(rst), .Q(creg[383]) );
  DFF \creg_reg[384]  ( .D(n6801), .CLK(clk), .RST(rst), .Q(creg[384]) );
  DFF \creg_reg[385]  ( .D(n6800), .CLK(clk), .RST(rst), .Q(creg[385]) );
  DFF \creg_reg[386]  ( .D(n6799), .CLK(clk), .RST(rst), .Q(creg[386]) );
  DFF \creg_reg[387]  ( .D(n6798), .CLK(clk), .RST(rst), .Q(creg[387]) );
  DFF \creg_reg[388]  ( .D(n6797), .CLK(clk), .RST(rst), .Q(creg[388]) );
  DFF \creg_reg[389]  ( .D(n6796), .CLK(clk), .RST(rst), .Q(creg[389]) );
  DFF \creg_reg[390]  ( .D(n6795), .CLK(clk), .RST(rst), .Q(creg[390]) );
  DFF \creg_reg[391]  ( .D(n6794), .CLK(clk), .RST(rst), .Q(creg[391]) );
  DFF \creg_reg[392]  ( .D(n6793), .CLK(clk), .RST(rst), .Q(creg[392]) );
  DFF \creg_reg[393]  ( .D(n6792), .CLK(clk), .RST(rst), .Q(creg[393]) );
  DFF \creg_reg[394]  ( .D(n6791), .CLK(clk), .RST(rst), .Q(creg[394]) );
  DFF \creg_reg[395]  ( .D(n6790), .CLK(clk), .RST(rst), .Q(creg[395]) );
  DFF \creg_reg[396]  ( .D(n6789), .CLK(clk), .RST(rst), .Q(creg[396]) );
  DFF \creg_reg[397]  ( .D(n6788), .CLK(clk), .RST(rst), .Q(creg[397]) );
  DFF \creg_reg[398]  ( .D(n6787), .CLK(clk), .RST(rst), .Q(creg[398]) );
  DFF \creg_reg[399]  ( .D(n6786), .CLK(clk), .RST(rst), .Q(creg[399]) );
  DFF \creg_reg[400]  ( .D(n6785), .CLK(clk), .RST(rst), .Q(creg[400]) );
  DFF \creg_reg[401]  ( .D(n6784), .CLK(clk), .RST(rst), .Q(creg[401]) );
  DFF \creg_reg[402]  ( .D(n6783), .CLK(clk), .RST(rst), .Q(creg[402]) );
  DFF \creg_reg[403]  ( .D(n6782), .CLK(clk), .RST(rst), .Q(creg[403]) );
  DFF \creg_reg[404]  ( .D(n6781), .CLK(clk), .RST(rst), .Q(creg[404]) );
  DFF \creg_reg[405]  ( .D(n6780), .CLK(clk), .RST(rst), .Q(creg[405]) );
  DFF \creg_reg[406]  ( .D(n6779), .CLK(clk), .RST(rst), .Q(creg[406]) );
  DFF \creg_reg[407]  ( .D(n6778), .CLK(clk), .RST(rst), .Q(creg[407]) );
  DFF \creg_reg[408]  ( .D(n6777), .CLK(clk), .RST(rst), .Q(creg[408]) );
  DFF \creg_reg[409]  ( .D(n6776), .CLK(clk), .RST(rst), .Q(creg[409]) );
  DFF \creg_reg[410]  ( .D(n6775), .CLK(clk), .RST(rst), .Q(creg[410]) );
  DFF \creg_reg[411]  ( .D(n6774), .CLK(clk), .RST(rst), .Q(creg[411]) );
  DFF \creg_reg[412]  ( .D(n6773), .CLK(clk), .RST(rst), .Q(creg[412]) );
  DFF \creg_reg[413]  ( .D(n6772), .CLK(clk), .RST(rst), .Q(creg[413]) );
  DFF \creg_reg[414]  ( .D(n6771), .CLK(clk), .RST(rst), .Q(creg[414]) );
  DFF \creg_reg[415]  ( .D(n6770), .CLK(clk), .RST(rst), .Q(creg[415]) );
  DFF \creg_reg[416]  ( .D(n6769), .CLK(clk), .RST(rst), .Q(creg[416]) );
  DFF \creg_reg[417]  ( .D(n6768), .CLK(clk), .RST(rst), .Q(creg[417]) );
  DFF \creg_reg[418]  ( .D(n6767), .CLK(clk), .RST(rst), .Q(creg[418]) );
  DFF \creg_reg[419]  ( .D(n6766), .CLK(clk), .RST(rst), .Q(creg[419]) );
  DFF \creg_reg[420]  ( .D(n6765), .CLK(clk), .RST(rst), .Q(creg[420]) );
  DFF \creg_reg[421]  ( .D(n6764), .CLK(clk), .RST(rst), .Q(creg[421]) );
  DFF \creg_reg[422]  ( .D(n6763), .CLK(clk), .RST(rst), .Q(creg[422]) );
  DFF \creg_reg[423]  ( .D(n6762), .CLK(clk), .RST(rst), .Q(creg[423]) );
  DFF \creg_reg[424]  ( .D(n6761), .CLK(clk), .RST(rst), .Q(creg[424]) );
  DFF \creg_reg[425]  ( .D(n6760), .CLK(clk), .RST(rst), .Q(creg[425]) );
  DFF \creg_reg[426]  ( .D(n6759), .CLK(clk), .RST(rst), .Q(creg[426]) );
  DFF \creg_reg[427]  ( .D(n6758), .CLK(clk), .RST(rst), .Q(creg[427]) );
  DFF \creg_reg[428]  ( .D(n6757), .CLK(clk), .RST(rst), .Q(creg[428]) );
  DFF \creg_reg[429]  ( .D(n6756), .CLK(clk), .RST(rst), .Q(creg[429]) );
  DFF \creg_reg[430]  ( .D(n6755), .CLK(clk), .RST(rst), .Q(creg[430]) );
  DFF \creg_reg[431]  ( .D(n6754), .CLK(clk), .RST(rst), .Q(creg[431]) );
  DFF \creg_reg[432]  ( .D(n6753), .CLK(clk), .RST(rst), .Q(creg[432]) );
  DFF \creg_reg[433]  ( .D(n6752), .CLK(clk), .RST(rst), .Q(creg[433]) );
  DFF \creg_reg[434]  ( .D(n6751), .CLK(clk), .RST(rst), .Q(creg[434]) );
  DFF \creg_reg[435]  ( .D(n6750), .CLK(clk), .RST(rst), .Q(creg[435]) );
  DFF \creg_reg[436]  ( .D(n6749), .CLK(clk), .RST(rst), .Q(creg[436]) );
  DFF \creg_reg[437]  ( .D(n6748), .CLK(clk), .RST(rst), .Q(creg[437]) );
  DFF \creg_reg[438]  ( .D(n6747), .CLK(clk), .RST(rst), .Q(creg[438]) );
  DFF \creg_reg[439]  ( .D(n6746), .CLK(clk), .RST(rst), .Q(creg[439]) );
  DFF \creg_reg[440]  ( .D(n6745), .CLK(clk), .RST(rst), .Q(creg[440]) );
  DFF \creg_reg[441]  ( .D(n6744), .CLK(clk), .RST(rst), .Q(creg[441]) );
  DFF \creg_reg[442]  ( .D(n6743), .CLK(clk), .RST(rst), .Q(creg[442]) );
  DFF \creg_reg[443]  ( .D(n6742), .CLK(clk), .RST(rst), .Q(creg[443]) );
  DFF \creg_reg[444]  ( .D(n6741), .CLK(clk), .RST(rst), .Q(creg[444]) );
  DFF \creg_reg[445]  ( .D(n6740), .CLK(clk), .RST(rst), .Q(creg[445]) );
  DFF \creg_reg[446]  ( .D(n6739), .CLK(clk), .RST(rst), .Q(creg[446]) );
  DFF \creg_reg[447]  ( .D(n6738), .CLK(clk), .RST(rst), .Q(creg[447]) );
  DFF \creg_reg[448]  ( .D(n6737), .CLK(clk), .RST(rst), .Q(creg[448]) );
  DFF \creg_reg[449]  ( .D(n6736), .CLK(clk), .RST(rst), .Q(creg[449]) );
  DFF \creg_reg[450]  ( .D(n6735), .CLK(clk), .RST(rst), .Q(creg[450]) );
  DFF \creg_reg[451]  ( .D(n6734), .CLK(clk), .RST(rst), .Q(creg[451]) );
  DFF \creg_reg[452]  ( .D(n6733), .CLK(clk), .RST(rst), .Q(creg[452]) );
  DFF \creg_reg[453]  ( .D(n6732), .CLK(clk), .RST(rst), .Q(creg[453]) );
  DFF \creg_reg[454]  ( .D(n6731), .CLK(clk), .RST(rst), .Q(creg[454]) );
  DFF \creg_reg[455]  ( .D(n6730), .CLK(clk), .RST(rst), .Q(creg[455]) );
  DFF \creg_reg[456]  ( .D(n6729), .CLK(clk), .RST(rst), .Q(creg[456]) );
  DFF \creg_reg[457]  ( .D(n6728), .CLK(clk), .RST(rst), .Q(creg[457]) );
  DFF \creg_reg[458]  ( .D(n6727), .CLK(clk), .RST(rst), .Q(creg[458]) );
  DFF \creg_reg[459]  ( .D(n6726), .CLK(clk), .RST(rst), .Q(creg[459]) );
  DFF \creg_reg[460]  ( .D(n6725), .CLK(clk), .RST(rst), .Q(creg[460]) );
  DFF \creg_reg[461]  ( .D(n6724), .CLK(clk), .RST(rst), .Q(creg[461]) );
  DFF \creg_reg[462]  ( .D(n6723), .CLK(clk), .RST(rst), .Q(creg[462]) );
  DFF \creg_reg[463]  ( .D(n6722), .CLK(clk), .RST(rst), .Q(creg[463]) );
  DFF \creg_reg[464]  ( .D(n6721), .CLK(clk), .RST(rst), .Q(creg[464]) );
  DFF \creg_reg[465]  ( .D(n6720), .CLK(clk), .RST(rst), .Q(creg[465]) );
  DFF \creg_reg[466]  ( .D(n6719), .CLK(clk), .RST(rst), .Q(creg[466]) );
  DFF \creg_reg[467]  ( .D(n6718), .CLK(clk), .RST(rst), .Q(creg[467]) );
  DFF \creg_reg[468]  ( .D(n6717), .CLK(clk), .RST(rst), .Q(creg[468]) );
  DFF \creg_reg[469]  ( .D(n6716), .CLK(clk), .RST(rst), .Q(creg[469]) );
  DFF \creg_reg[470]  ( .D(n6715), .CLK(clk), .RST(rst), .Q(creg[470]) );
  DFF \creg_reg[471]  ( .D(n6714), .CLK(clk), .RST(rst), .Q(creg[471]) );
  DFF \creg_reg[472]  ( .D(n6713), .CLK(clk), .RST(rst), .Q(creg[472]) );
  DFF \creg_reg[473]  ( .D(n6712), .CLK(clk), .RST(rst), .Q(creg[473]) );
  DFF \creg_reg[474]  ( .D(n6711), .CLK(clk), .RST(rst), .Q(creg[474]) );
  DFF \creg_reg[475]  ( .D(n6710), .CLK(clk), .RST(rst), .Q(creg[475]) );
  DFF \creg_reg[476]  ( .D(n6709), .CLK(clk), .RST(rst), .Q(creg[476]) );
  DFF \creg_reg[477]  ( .D(n6708), .CLK(clk), .RST(rst), .Q(creg[477]) );
  DFF \creg_reg[478]  ( .D(n6707), .CLK(clk), .RST(rst), .Q(creg[478]) );
  DFF \creg_reg[479]  ( .D(n6706), .CLK(clk), .RST(rst), .Q(creg[479]) );
  DFF \creg_reg[480]  ( .D(n6705), .CLK(clk), .RST(rst), .Q(creg[480]) );
  DFF \creg_reg[481]  ( .D(n6704), .CLK(clk), .RST(rst), .Q(creg[481]) );
  DFF \creg_reg[482]  ( .D(n6703), .CLK(clk), .RST(rst), .Q(creg[482]) );
  DFF \creg_reg[483]  ( .D(n6702), .CLK(clk), .RST(rst), .Q(creg[483]) );
  DFF \creg_reg[484]  ( .D(n6701), .CLK(clk), .RST(rst), .Q(creg[484]) );
  DFF \creg_reg[485]  ( .D(n6700), .CLK(clk), .RST(rst), .Q(creg[485]) );
  DFF \creg_reg[486]  ( .D(n6699), .CLK(clk), .RST(rst), .Q(creg[486]) );
  DFF \creg_reg[487]  ( .D(n6698), .CLK(clk), .RST(rst), .Q(creg[487]) );
  DFF \creg_reg[488]  ( .D(n6697), .CLK(clk), .RST(rst), .Q(creg[488]) );
  DFF \creg_reg[489]  ( .D(n6696), .CLK(clk), .RST(rst), .Q(creg[489]) );
  DFF \creg_reg[490]  ( .D(n6695), .CLK(clk), .RST(rst), .Q(creg[490]) );
  DFF \creg_reg[491]  ( .D(n6694), .CLK(clk), .RST(rst), .Q(creg[491]) );
  DFF \creg_reg[492]  ( .D(n6693), .CLK(clk), .RST(rst), .Q(creg[492]) );
  DFF \creg_reg[493]  ( .D(n6692), .CLK(clk), .RST(rst), .Q(creg[493]) );
  DFF \creg_reg[494]  ( .D(n6691), .CLK(clk), .RST(rst), .Q(creg[494]) );
  DFF \creg_reg[495]  ( .D(n6690), .CLK(clk), .RST(rst), .Q(creg[495]) );
  DFF \creg_reg[496]  ( .D(n6689), .CLK(clk), .RST(rst), .Q(creg[496]) );
  DFF \creg_reg[497]  ( .D(n6688), .CLK(clk), .RST(rst), .Q(creg[497]) );
  DFF \creg_reg[498]  ( .D(n6687), .CLK(clk), .RST(rst), .Q(creg[498]) );
  DFF \creg_reg[499]  ( .D(n6686), .CLK(clk), .RST(rst), .Q(creg[499]) );
  DFF \creg_reg[500]  ( .D(n6685), .CLK(clk), .RST(rst), .Q(creg[500]) );
  DFF \creg_reg[501]  ( .D(n6684), .CLK(clk), .RST(rst), .Q(creg[501]) );
  DFF \creg_reg[502]  ( .D(n6683), .CLK(clk), .RST(rst), .Q(creg[502]) );
  DFF \creg_reg[503]  ( .D(n6682), .CLK(clk), .RST(rst), .Q(creg[503]) );
  DFF \creg_reg[504]  ( .D(n6681), .CLK(clk), .RST(rst), .Q(creg[504]) );
  DFF \creg_reg[505]  ( .D(n6680), .CLK(clk), .RST(rst), .Q(creg[505]) );
  DFF \creg_reg[506]  ( .D(n6679), .CLK(clk), .RST(rst), .Q(creg[506]) );
  DFF \creg_reg[507]  ( .D(n6678), .CLK(clk), .RST(rst), .Q(creg[507]) );
  DFF \creg_reg[508]  ( .D(n6677), .CLK(clk), .RST(rst), .Q(creg[508]) );
  DFF \creg_reg[509]  ( .D(n6676), .CLK(clk), .RST(rst), .Q(creg[509]) );
  DFF \creg_reg[510]  ( .D(n6675), .CLK(clk), .RST(rst), .Q(creg[510]) );
  DFF \creg_reg[511]  ( .D(n7186), .CLK(clk), .RST(rst), .Q(creg[511]) );
  modmult_N512_CC512 modmult_1 ( .clk(clk), .rst(rst), .start(start_in[0]), 
        .x(x), .y(y), .n(n), .o(o) );
  NAND U9750 ( .A(n7700), .B(n7701), .Z(y[9]) );
  NAND U9751 ( .A(n7702), .B(m[9]), .Z(n7701) );
  NAND U9752 ( .A(n7703), .B(creg[9]), .Z(n7700) );
  NAND U9753 ( .A(n7704), .B(n7705), .Z(y[99]) );
  NAND U9754 ( .A(n7702), .B(m[99]), .Z(n7705) );
  NAND U9755 ( .A(n7703), .B(creg[99]), .Z(n7704) );
  NAND U9756 ( .A(n7706), .B(n7707), .Z(y[98]) );
  NAND U9757 ( .A(n7702), .B(m[98]), .Z(n7707) );
  NAND U9758 ( .A(n7703), .B(creg[98]), .Z(n7706) );
  NAND U9759 ( .A(n7708), .B(n7709), .Z(y[97]) );
  NAND U9760 ( .A(n7702), .B(m[97]), .Z(n7709) );
  NAND U9761 ( .A(n7703), .B(creg[97]), .Z(n7708) );
  NAND U9762 ( .A(n7710), .B(n7711), .Z(y[96]) );
  NAND U9763 ( .A(n7702), .B(m[96]), .Z(n7711) );
  NAND U9764 ( .A(n7703), .B(creg[96]), .Z(n7710) );
  NAND U9765 ( .A(n7712), .B(n7713), .Z(y[95]) );
  NAND U9766 ( .A(n7702), .B(m[95]), .Z(n7713) );
  NAND U9767 ( .A(n7703), .B(creg[95]), .Z(n7712) );
  NAND U9768 ( .A(n7714), .B(n7715), .Z(y[94]) );
  NAND U9769 ( .A(n7702), .B(m[94]), .Z(n7715) );
  NAND U9770 ( .A(n7703), .B(creg[94]), .Z(n7714) );
  NAND U9771 ( .A(n7716), .B(n7717), .Z(y[93]) );
  NAND U9772 ( .A(n7702), .B(m[93]), .Z(n7717) );
  NAND U9773 ( .A(n7703), .B(creg[93]), .Z(n7716) );
  NAND U9774 ( .A(n7718), .B(n7719), .Z(y[92]) );
  NAND U9775 ( .A(n7702), .B(m[92]), .Z(n7719) );
  NAND U9776 ( .A(n7703), .B(creg[92]), .Z(n7718) );
  NAND U9777 ( .A(n7720), .B(n7721), .Z(y[91]) );
  NAND U9778 ( .A(n7702), .B(m[91]), .Z(n7721) );
  NAND U9779 ( .A(n7703), .B(creg[91]), .Z(n7720) );
  NAND U9780 ( .A(n7722), .B(n7723), .Z(y[90]) );
  NAND U9781 ( .A(n7702), .B(m[90]), .Z(n7723) );
  NAND U9782 ( .A(n7703), .B(creg[90]), .Z(n7722) );
  NAND U9783 ( .A(n7724), .B(n7725), .Z(y[8]) );
  NAND U9784 ( .A(n7702), .B(m[8]), .Z(n7725) );
  NAND U9785 ( .A(n7703), .B(creg[8]), .Z(n7724) );
  NAND U9786 ( .A(n7726), .B(n7727), .Z(y[89]) );
  NAND U9787 ( .A(n7702), .B(m[89]), .Z(n7727) );
  NAND U9788 ( .A(n7703), .B(creg[89]), .Z(n7726) );
  NAND U9789 ( .A(n7728), .B(n7729), .Z(y[88]) );
  NAND U9790 ( .A(n7702), .B(m[88]), .Z(n7729) );
  NAND U9791 ( .A(n7703), .B(creg[88]), .Z(n7728) );
  NAND U9792 ( .A(n7730), .B(n7731), .Z(y[87]) );
  NAND U9793 ( .A(n7702), .B(m[87]), .Z(n7731) );
  NAND U9794 ( .A(n7703), .B(creg[87]), .Z(n7730) );
  NAND U9795 ( .A(n7732), .B(n7733), .Z(y[86]) );
  NAND U9796 ( .A(n7702), .B(m[86]), .Z(n7733) );
  NAND U9797 ( .A(n7703), .B(creg[86]), .Z(n7732) );
  NAND U9798 ( .A(n7734), .B(n7735), .Z(y[85]) );
  NAND U9799 ( .A(n7702), .B(m[85]), .Z(n7735) );
  NAND U9800 ( .A(n7703), .B(creg[85]), .Z(n7734) );
  NAND U9801 ( .A(n7736), .B(n7737), .Z(y[84]) );
  NAND U9802 ( .A(n7702), .B(m[84]), .Z(n7737) );
  NAND U9803 ( .A(n7703), .B(creg[84]), .Z(n7736) );
  NAND U9804 ( .A(n7738), .B(n7739), .Z(y[83]) );
  NAND U9805 ( .A(n7702), .B(m[83]), .Z(n7739) );
  NAND U9806 ( .A(n7703), .B(creg[83]), .Z(n7738) );
  NAND U9807 ( .A(n7740), .B(n7741), .Z(y[82]) );
  NAND U9808 ( .A(n7702), .B(m[82]), .Z(n7741) );
  NAND U9809 ( .A(n7703), .B(creg[82]), .Z(n7740) );
  NAND U9810 ( .A(n7742), .B(n7743), .Z(y[81]) );
  NAND U9811 ( .A(n7702), .B(m[81]), .Z(n7743) );
  NAND U9812 ( .A(n7703), .B(creg[81]), .Z(n7742) );
  NAND U9813 ( .A(n7744), .B(n7745), .Z(y[80]) );
  NAND U9814 ( .A(n7702), .B(m[80]), .Z(n7745) );
  NAND U9815 ( .A(n7703), .B(creg[80]), .Z(n7744) );
  NAND U9816 ( .A(n7746), .B(n7747), .Z(y[7]) );
  NAND U9817 ( .A(n7702), .B(m[7]), .Z(n7747) );
  NAND U9818 ( .A(n7703), .B(creg[7]), .Z(n7746) );
  NAND U9819 ( .A(n7748), .B(n7749), .Z(y[79]) );
  NAND U9820 ( .A(n7702), .B(m[79]), .Z(n7749) );
  NAND U9821 ( .A(n7703), .B(creg[79]), .Z(n7748) );
  NAND U9822 ( .A(n7750), .B(n7751), .Z(y[78]) );
  NAND U9823 ( .A(n7702), .B(m[78]), .Z(n7751) );
  NAND U9824 ( .A(n7703), .B(creg[78]), .Z(n7750) );
  NAND U9825 ( .A(n7752), .B(n7753), .Z(y[77]) );
  NAND U9826 ( .A(n7702), .B(m[77]), .Z(n7753) );
  NAND U9827 ( .A(n7703), .B(creg[77]), .Z(n7752) );
  NAND U9828 ( .A(n7754), .B(n7755), .Z(y[76]) );
  NAND U9829 ( .A(n7702), .B(m[76]), .Z(n7755) );
  NAND U9830 ( .A(n7703), .B(creg[76]), .Z(n7754) );
  NAND U9831 ( .A(n7756), .B(n7757), .Z(y[75]) );
  NAND U9832 ( .A(n7702), .B(m[75]), .Z(n7757) );
  NAND U9833 ( .A(n7703), .B(creg[75]), .Z(n7756) );
  NAND U9834 ( .A(n7758), .B(n7759), .Z(y[74]) );
  NAND U9835 ( .A(n7702), .B(m[74]), .Z(n7759) );
  NAND U9836 ( .A(n7703), .B(creg[74]), .Z(n7758) );
  NAND U9837 ( .A(n7760), .B(n7761), .Z(y[73]) );
  NAND U9838 ( .A(n7702), .B(m[73]), .Z(n7761) );
  NAND U9839 ( .A(n7703), .B(creg[73]), .Z(n7760) );
  NAND U9840 ( .A(n7762), .B(n7763), .Z(y[72]) );
  NAND U9841 ( .A(n7702), .B(m[72]), .Z(n7763) );
  NAND U9842 ( .A(n7703), .B(creg[72]), .Z(n7762) );
  NAND U9843 ( .A(n7764), .B(n7765), .Z(y[71]) );
  NAND U9844 ( .A(n7702), .B(m[71]), .Z(n7765) );
  NAND U9845 ( .A(n7703), .B(creg[71]), .Z(n7764) );
  NAND U9846 ( .A(n7766), .B(n7767), .Z(y[70]) );
  NAND U9847 ( .A(n7702), .B(m[70]), .Z(n7767) );
  NAND U9848 ( .A(n7703), .B(creg[70]), .Z(n7766) );
  NAND U9849 ( .A(n7768), .B(n7769), .Z(y[6]) );
  NAND U9850 ( .A(n7702), .B(m[6]), .Z(n7769) );
  NAND U9851 ( .A(n7703), .B(creg[6]), .Z(n7768) );
  NAND U9852 ( .A(n7770), .B(n7771), .Z(y[69]) );
  NAND U9853 ( .A(n7702), .B(m[69]), .Z(n7771) );
  NAND U9854 ( .A(n7703), .B(creg[69]), .Z(n7770) );
  NAND U9855 ( .A(n7772), .B(n7773), .Z(y[68]) );
  NAND U9856 ( .A(n7702), .B(m[68]), .Z(n7773) );
  NAND U9857 ( .A(n7703), .B(creg[68]), .Z(n7772) );
  NAND U9858 ( .A(n7774), .B(n7775), .Z(y[67]) );
  NAND U9859 ( .A(n7702), .B(m[67]), .Z(n7775) );
  NAND U9860 ( .A(n7703), .B(creg[67]), .Z(n7774) );
  NAND U9861 ( .A(n7776), .B(n7777), .Z(y[66]) );
  NAND U9862 ( .A(n7702), .B(m[66]), .Z(n7777) );
  NAND U9863 ( .A(n7703), .B(creg[66]), .Z(n7776) );
  NAND U9864 ( .A(n7778), .B(n7779), .Z(y[65]) );
  NAND U9865 ( .A(n7702), .B(m[65]), .Z(n7779) );
  NAND U9866 ( .A(n7703), .B(creg[65]), .Z(n7778) );
  NAND U9867 ( .A(n7780), .B(n7781), .Z(y[64]) );
  NAND U9868 ( .A(n7702), .B(m[64]), .Z(n7781) );
  NAND U9869 ( .A(n7703), .B(creg[64]), .Z(n7780) );
  NAND U9870 ( .A(n7782), .B(n7783), .Z(y[63]) );
  NAND U9871 ( .A(n7702), .B(m[63]), .Z(n7783) );
  NAND U9872 ( .A(n7703), .B(creg[63]), .Z(n7782) );
  NAND U9873 ( .A(n7784), .B(n7785), .Z(y[62]) );
  NAND U9874 ( .A(n7702), .B(m[62]), .Z(n7785) );
  NAND U9875 ( .A(n7703), .B(creg[62]), .Z(n7784) );
  NAND U9876 ( .A(n7786), .B(n7787), .Z(y[61]) );
  NAND U9877 ( .A(n7702), .B(m[61]), .Z(n7787) );
  NAND U9878 ( .A(n7703), .B(creg[61]), .Z(n7786) );
  NAND U9879 ( .A(n7788), .B(n7789), .Z(y[60]) );
  NAND U9880 ( .A(n7702), .B(m[60]), .Z(n7789) );
  NAND U9881 ( .A(n7703), .B(creg[60]), .Z(n7788) );
  NAND U9882 ( .A(n7790), .B(n7791), .Z(y[5]) );
  NAND U9883 ( .A(n7702), .B(m[5]), .Z(n7791) );
  NAND U9884 ( .A(n7703), .B(creg[5]), .Z(n7790) );
  NAND U9885 ( .A(n7792), .B(n7793), .Z(y[59]) );
  NAND U9886 ( .A(n7702), .B(m[59]), .Z(n7793) );
  NAND U9887 ( .A(n7703), .B(creg[59]), .Z(n7792) );
  NAND U9888 ( .A(n7794), .B(n7795), .Z(y[58]) );
  NAND U9889 ( .A(n7702), .B(m[58]), .Z(n7795) );
  NAND U9890 ( .A(n7703), .B(creg[58]), .Z(n7794) );
  NAND U9891 ( .A(n7796), .B(n7797), .Z(y[57]) );
  NAND U9892 ( .A(n7702), .B(m[57]), .Z(n7797) );
  NAND U9893 ( .A(n7703), .B(creg[57]), .Z(n7796) );
  NAND U9894 ( .A(n7798), .B(n7799), .Z(y[56]) );
  NAND U9895 ( .A(n7702), .B(m[56]), .Z(n7799) );
  NAND U9896 ( .A(n7703), .B(creg[56]), .Z(n7798) );
  NAND U9897 ( .A(n7800), .B(n7801), .Z(y[55]) );
  NAND U9898 ( .A(n7702), .B(m[55]), .Z(n7801) );
  NAND U9899 ( .A(n7703), .B(creg[55]), .Z(n7800) );
  NAND U9900 ( .A(n7802), .B(n7803), .Z(y[54]) );
  NAND U9901 ( .A(n7702), .B(m[54]), .Z(n7803) );
  NAND U9902 ( .A(n7703), .B(creg[54]), .Z(n7802) );
  NAND U9903 ( .A(n7804), .B(n7805), .Z(y[53]) );
  NAND U9904 ( .A(n7702), .B(m[53]), .Z(n7805) );
  NAND U9905 ( .A(n7703), .B(creg[53]), .Z(n7804) );
  NAND U9906 ( .A(n7806), .B(n7807), .Z(y[52]) );
  NAND U9907 ( .A(n7702), .B(m[52]), .Z(n7807) );
  NAND U9908 ( .A(n7703), .B(creg[52]), .Z(n7806) );
  NAND U9909 ( .A(n7808), .B(n7809), .Z(y[51]) );
  NAND U9910 ( .A(n7702), .B(m[51]), .Z(n7809) );
  NAND U9911 ( .A(n7703), .B(creg[51]), .Z(n7808) );
  NAND U9912 ( .A(n7810), .B(n7811), .Z(y[511]) );
  NAND U9913 ( .A(n7702), .B(m[511]), .Z(n7811) );
  NAND U9914 ( .A(n7703), .B(creg[511]), .Z(n7810) );
  NAND U9915 ( .A(n7812), .B(n7813), .Z(y[510]) );
  NAND U9916 ( .A(n7702), .B(m[510]), .Z(n7813) );
  NAND U9917 ( .A(n7703), .B(creg[510]), .Z(n7812) );
  NAND U9918 ( .A(n7814), .B(n7815), .Z(y[50]) );
  NAND U9919 ( .A(n7702), .B(m[50]), .Z(n7815) );
  NAND U9920 ( .A(n7703), .B(creg[50]), .Z(n7814) );
  NAND U9921 ( .A(n7816), .B(n7817), .Z(y[509]) );
  NAND U9922 ( .A(n7702), .B(m[509]), .Z(n7817) );
  NAND U9923 ( .A(n7703), .B(creg[509]), .Z(n7816) );
  NAND U9924 ( .A(n7818), .B(n7819), .Z(y[508]) );
  NAND U9925 ( .A(n7702), .B(m[508]), .Z(n7819) );
  NAND U9926 ( .A(n7703), .B(creg[508]), .Z(n7818) );
  NAND U9927 ( .A(n7820), .B(n7821), .Z(y[507]) );
  NAND U9928 ( .A(n7702), .B(m[507]), .Z(n7821) );
  NAND U9929 ( .A(n7703), .B(creg[507]), .Z(n7820) );
  NAND U9930 ( .A(n7822), .B(n7823), .Z(y[506]) );
  NAND U9931 ( .A(n7702), .B(m[506]), .Z(n7823) );
  NAND U9932 ( .A(n7703), .B(creg[506]), .Z(n7822) );
  NAND U9933 ( .A(n7824), .B(n7825), .Z(y[505]) );
  NAND U9934 ( .A(n7702), .B(m[505]), .Z(n7825) );
  NAND U9935 ( .A(n7703), .B(creg[505]), .Z(n7824) );
  NAND U9936 ( .A(n7826), .B(n7827), .Z(y[504]) );
  NAND U9937 ( .A(n7702), .B(m[504]), .Z(n7827) );
  NAND U9938 ( .A(n7703), .B(creg[504]), .Z(n7826) );
  NAND U9939 ( .A(n7828), .B(n7829), .Z(y[503]) );
  NAND U9940 ( .A(n7702), .B(m[503]), .Z(n7829) );
  NAND U9941 ( .A(n7703), .B(creg[503]), .Z(n7828) );
  NAND U9942 ( .A(n7830), .B(n7831), .Z(y[502]) );
  NAND U9943 ( .A(n7702), .B(m[502]), .Z(n7831) );
  NAND U9944 ( .A(n7703), .B(creg[502]), .Z(n7830) );
  NAND U9945 ( .A(n7832), .B(n7833), .Z(y[501]) );
  NAND U9946 ( .A(n7702), .B(m[501]), .Z(n7833) );
  NAND U9947 ( .A(n7703), .B(creg[501]), .Z(n7832) );
  NAND U9948 ( .A(n7834), .B(n7835), .Z(y[500]) );
  NAND U9949 ( .A(n7702), .B(m[500]), .Z(n7835) );
  NAND U9950 ( .A(n7703), .B(creg[500]), .Z(n7834) );
  NAND U9951 ( .A(n7836), .B(n7837), .Z(y[4]) );
  NAND U9952 ( .A(n7702), .B(m[4]), .Z(n7837) );
  NAND U9953 ( .A(n7703), .B(creg[4]), .Z(n7836) );
  NAND U9954 ( .A(n7838), .B(n7839), .Z(y[49]) );
  NAND U9955 ( .A(n7702), .B(m[49]), .Z(n7839) );
  NAND U9956 ( .A(n7703), .B(creg[49]), .Z(n7838) );
  NAND U9957 ( .A(n7840), .B(n7841), .Z(y[499]) );
  NAND U9958 ( .A(n7702), .B(m[499]), .Z(n7841) );
  NAND U9959 ( .A(n7703), .B(creg[499]), .Z(n7840) );
  NAND U9960 ( .A(n7842), .B(n7843), .Z(y[498]) );
  NAND U9961 ( .A(n7702), .B(m[498]), .Z(n7843) );
  NAND U9962 ( .A(n7703), .B(creg[498]), .Z(n7842) );
  NAND U9963 ( .A(n7844), .B(n7845), .Z(y[497]) );
  NAND U9964 ( .A(n7702), .B(m[497]), .Z(n7845) );
  NAND U9965 ( .A(n7703), .B(creg[497]), .Z(n7844) );
  NAND U9966 ( .A(n7846), .B(n7847), .Z(y[496]) );
  NAND U9967 ( .A(n7702), .B(m[496]), .Z(n7847) );
  NAND U9968 ( .A(n7703), .B(creg[496]), .Z(n7846) );
  NAND U9969 ( .A(n7848), .B(n7849), .Z(y[495]) );
  NAND U9970 ( .A(n7702), .B(m[495]), .Z(n7849) );
  NAND U9971 ( .A(n7703), .B(creg[495]), .Z(n7848) );
  NAND U9972 ( .A(n7850), .B(n7851), .Z(y[494]) );
  NAND U9973 ( .A(n7702), .B(m[494]), .Z(n7851) );
  NAND U9974 ( .A(n7703), .B(creg[494]), .Z(n7850) );
  NAND U9975 ( .A(n7852), .B(n7853), .Z(y[493]) );
  NAND U9976 ( .A(n7702), .B(m[493]), .Z(n7853) );
  NAND U9977 ( .A(n7703), .B(creg[493]), .Z(n7852) );
  NAND U9978 ( .A(n7854), .B(n7855), .Z(y[492]) );
  NAND U9979 ( .A(n7702), .B(m[492]), .Z(n7855) );
  NAND U9980 ( .A(n7703), .B(creg[492]), .Z(n7854) );
  NAND U9981 ( .A(n7856), .B(n7857), .Z(y[491]) );
  NAND U9982 ( .A(n7702), .B(m[491]), .Z(n7857) );
  NAND U9983 ( .A(n7703), .B(creg[491]), .Z(n7856) );
  NAND U9984 ( .A(n7858), .B(n7859), .Z(y[490]) );
  NAND U9985 ( .A(n7702), .B(m[490]), .Z(n7859) );
  NAND U9986 ( .A(n7703), .B(creg[490]), .Z(n7858) );
  NAND U9987 ( .A(n7860), .B(n7861), .Z(y[48]) );
  NAND U9988 ( .A(n7702), .B(m[48]), .Z(n7861) );
  NAND U9989 ( .A(n7703), .B(creg[48]), .Z(n7860) );
  NAND U9990 ( .A(n7862), .B(n7863), .Z(y[489]) );
  NAND U9991 ( .A(n7702), .B(m[489]), .Z(n7863) );
  NAND U9992 ( .A(n7703), .B(creg[489]), .Z(n7862) );
  NAND U9993 ( .A(n7864), .B(n7865), .Z(y[488]) );
  NAND U9994 ( .A(n7702), .B(m[488]), .Z(n7865) );
  NAND U9995 ( .A(n7703), .B(creg[488]), .Z(n7864) );
  NAND U9996 ( .A(n7866), .B(n7867), .Z(y[487]) );
  NAND U9997 ( .A(n7702), .B(m[487]), .Z(n7867) );
  NAND U9998 ( .A(n7703), .B(creg[487]), .Z(n7866) );
  NAND U9999 ( .A(n7868), .B(n7869), .Z(y[486]) );
  NAND U10000 ( .A(n7702), .B(m[486]), .Z(n7869) );
  NAND U10001 ( .A(n7703), .B(creg[486]), .Z(n7868) );
  NAND U10002 ( .A(n7870), .B(n7871), .Z(y[485]) );
  NAND U10003 ( .A(n7702), .B(m[485]), .Z(n7871) );
  NAND U10004 ( .A(n7703), .B(creg[485]), .Z(n7870) );
  NAND U10005 ( .A(n7872), .B(n7873), .Z(y[484]) );
  NAND U10006 ( .A(n7702), .B(m[484]), .Z(n7873) );
  NAND U10007 ( .A(n7703), .B(creg[484]), .Z(n7872) );
  NAND U10008 ( .A(n7874), .B(n7875), .Z(y[483]) );
  NAND U10009 ( .A(n7702), .B(m[483]), .Z(n7875) );
  NAND U10010 ( .A(n7703), .B(creg[483]), .Z(n7874) );
  NAND U10011 ( .A(n7876), .B(n7877), .Z(y[482]) );
  NAND U10012 ( .A(n7702), .B(m[482]), .Z(n7877) );
  NAND U10013 ( .A(n7703), .B(creg[482]), .Z(n7876) );
  NAND U10014 ( .A(n7878), .B(n7879), .Z(y[481]) );
  NAND U10015 ( .A(n7702), .B(m[481]), .Z(n7879) );
  NAND U10016 ( .A(n7703), .B(creg[481]), .Z(n7878) );
  NAND U10017 ( .A(n7880), .B(n7881), .Z(y[480]) );
  NAND U10018 ( .A(n7702), .B(m[480]), .Z(n7881) );
  NAND U10019 ( .A(n7703), .B(creg[480]), .Z(n7880) );
  NAND U10020 ( .A(n7882), .B(n7883), .Z(y[47]) );
  NAND U10021 ( .A(n7702), .B(m[47]), .Z(n7883) );
  NAND U10022 ( .A(n7703), .B(creg[47]), .Z(n7882) );
  NAND U10023 ( .A(n7884), .B(n7885), .Z(y[479]) );
  NAND U10024 ( .A(n7702), .B(m[479]), .Z(n7885) );
  NAND U10025 ( .A(n7703), .B(creg[479]), .Z(n7884) );
  NAND U10026 ( .A(n7886), .B(n7887), .Z(y[478]) );
  NAND U10027 ( .A(n7702), .B(m[478]), .Z(n7887) );
  NAND U10028 ( .A(n7703), .B(creg[478]), .Z(n7886) );
  NAND U10029 ( .A(n7888), .B(n7889), .Z(y[477]) );
  NAND U10030 ( .A(n7702), .B(m[477]), .Z(n7889) );
  NAND U10031 ( .A(n7703), .B(creg[477]), .Z(n7888) );
  NAND U10032 ( .A(n7890), .B(n7891), .Z(y[476]) );
  NAND U10033 ( .A(n7702), .B(m[476]), .Z(n7891) );
  NAND U10034 ( .A(n7703), .B(creg[476]), .Z(n7890) );
  NAND U10035 ( .A(n7892), .B(n7893), .Z(y[475]) );
  NAND U10036 ( .A(n7702), .B(m[475]), .Z(n7893) );
  NAND U10037 ( .A(n7703), .B(creg[475]), .Z(n7892) );
  NAND U10038 ( .A(n7894), .B(n7895), .Z(y[474]) );
  NAND U10039 ( .A(n7702), .B(m[474]), .Z(n7895) );
  NAND U10040 ( .A(n7703), .B(creg[474]), .Z(n7894) );
  NAND U10041 ( .A(n7896), .B(n7897), .Z(y[473]) );
  NAND U10042 ( .A(n7702), .B(m[473]), .Z(n7897) );
  NAND U10043 ( .A(n7703), .B(creg[473]), .Z(n7896) );
  NAND U10044 ( .A(n7898), .B(n7899), .Z(y[472]) );
  NAND U10045 ( .A(n7702), .B(m[472]), .Z(n7899) );
  NAND U10046 ( .A(n7703), .B(creg[472]), .Z(n7898) );
  NAND U10047 ( .A(n7900), .B(n7901), .Z(y[471]) );
  NAND U10048 ( .A(n7702), .B(m[471]), .Z(n7901) );
  NAND U10049 ( .A(n7703), .B(creg[471]), .Z(n7900) );
  NAND U10050 ( .A(n7902), .B(n7903), .Z(y[470]) );
  NAND U10051 ( .A(n7702), .B(m[470]), .Z(n7903) );
  NAND U10052 ( .A(n7703), .B(creg[470]), .Z(n7902) );
  NAND U10053 ( .A(n7904), .B(n7905), .Z(y[46]) );
  NAND U10054 ( .A(n7702), .B(m[46]), .Z(n7905) );
  NAND U10055 ( .A(n7703), .B(creg[46]), .Z(n7904) );
  NAND U10056 ( .A(n7906), .B(n7907), .Z(y[469]) );
  NAND U10057 ( .A(n7702), .B(m[469]), .Z(n7907) );
  NAND U10058 ( .A(n7703), .B(creg[469]), .Z(n7906) );
  NAND U10059 ( .A(n7908), .B(n7909), .Z(y[468]) );
  NAND U10060 ( .A(n7702), .B(m[468]), .Z(n7909) );
  NAND U10061 ( .A(n7703), .B(creg[468]), .Z(n7908) );
  NAND U10062 ( .A(n7910), .B(n7911), .Z(y[467]) );
  NAND U10063 ( .A(n7702), .B(m[467]), .Z(n7911) );
  NAND U10064 ( .A(n7703), .B(creg[467]), .Z(n7910) );
  NAND U10065 ( .A(n7912), .B(n7913), .Z(y[466]) );
  NAND U10066 ( .A(n7702), .B(m[466]), .Z(n7913) );
  NAND U10067 ( .A(n7703), .B(creg[466]), .Z(n7912) );
  NAND U10068 ( .A(n7914), .B(n7915), .Z(y[465]) );
  NAND U10069 ( .A(n7702), .B(m[465]), .Z(n7915) );
  NAND U10070 ( .A(n7703), .B(creg[465]), .Z(n7914) );
  NAND U10071 ( .A(n7916), .B(n7917), .Z(y[464]) );
  NAND U10072 ( .A(n7702), .B(m[464]), .Z(n7917) );
  NAND U10073 ( .A(n7703), .B(creg[464]), .Z(n7916) );
  NAND U10074 ( .A(n7918), .B(n7919), .Z(y[463]) );
  NAND U10075 ( .A(n7702), .B(m[463]), .Z(n7919) );
  NAND U10076 ( .A(n7703), .B(creg[463]), .Z(n7918) );
  NAND U10077 ( .A(n7920), .B(n7921), .Z(y[462]) );
  NAND U10078 ( .A(n7702), .B(m[462]), .Z(n7921) );
  NAND U10079 ( .A(n7703), .B(creg[462]), .Z(n7920) );
  NAND U10080 ( .A(n7922), .B(n7923), .Z(y[461]) );
  NAND U10081 ( .A(n7702), .B(m[461]), .Z(n7923) );
  NAND U10082 ( .A(n7703), .B(creg[461]), .Z(n7922) );
  NAND U10083 ( .A(n7924), .B(n7925), .Z(y[460]) );
  NAND U10084 ( .A(n7702), .B(m[460]), .Z(n7925) );
  NAND U10085 ( .A(n7703), .B(creg[460]), .Z(n7924) );
  NAND U10086 ( .A(n7926), .B(n7927), .Z(y[45]) );
  NAND U10087 ( .A(n7702), .B(m[45]), .Z(n7927) );
  NAND U10088 ( .A(n7703), .B(creg[45]), .Z(n7926) );
  NAND U10089 ( .A(n7928), .B(n7929), .Z(y[459]) );
  NAND U10090 ( .A(n7702), .B(m[459]), .Z(n7929) );
  NAND U10091 ( .A(n7703), .B(creg[459]), .Z(n7928) );
  NAND U10092 ( .A(n7930), .B(n7931), .Z(y[458]) );
  NAND U10093 ( .A(n7702), .B(m[458]), .Z(n7931) );
  NAND U10094 ( .A(n7703), .B(creg[458]), .Z(n7930) );
  NAND U10095 ( .A(n7932), .B(n7933), .Z(y[457]) );
  NAND U10096 ( .A(n7702), .B(m[457]), .Z(n7933) );
  NAND U10097 ( .A(n7703), .B(creg[457]), .Z(n7932) );
  NAND U10098 ( .A(n7934), .B(n7935), .Z(y[456]) );
  NAND U10099 ( .A(n7702), .B(m[456]), .Z(n7935) );
  NAND U10100 ( .A(n7703), .B(creg[456]), .Z(n7934) );
  NAND U10101 ( .A(n7936), .B(n7937), .Z(y[455]) );
  NAND U10102 ( .A(n7702), .B(m[455]), .Z(n7937) );
  NAND U10103 ( .A(n7703), .B(creg[455]), .Z(n7936) );
  NAND U10104 ( .A(n7938), .B(n7939), .Z(y[454]) );
  NAND U10105 ( .A(n7702), .B(m[454]), .Z(n7939) );
  NAND U10106 ( .A(n7703), .B(creg[454]), .Z(n7938) );
  NAND U10107 ( .A(n7940), .B(n7941), .Z(y[453]) );
  NAND U10108 ( .A(n7702), .B(m[453]), .Z(n7941) );
  NAND U10109 ( .A(n7703), .B(creg[453]), .Z(n7940) );
  NAND U10110 ( .A(n7942), .B(n7943), .Z(y[452]) );
  NAND U10111 ( .A(n7702), .B(m[452]), .Z(n7943) );
  NAND U10112 ( .A(n7703), .B(creg[452]), .Z(n7942) );
  NAND U10113 ( .A(n7944), .B(n7945), .Z(y[451]) );
  NAND U10114 ( .A(n7702), .B(m[451]), .Z(n7945) );
  NAND U10115 ( .A(n7703), .B(creg[451]), .Z(n7944) );
  NAND U10116 ( .A(n7946), .B(n7947), .Z(y[450]) );
  NAND U10117 ( .A(n7702), .B(m[450]), .Z(n7947) );
  NAND U10118 ( .A(n7703), .B(creg[450]), .Z(n7946) );
  NAND U10119 ( .A(n7948), .B(n7949), .Z(y[44]) );
  NAND U10120 ( .A(n7702), .B(m[44]), .Z(n7949) );
  NAND U10121 ( .A(n7703), .B(creg[44]), .Z(n7948) );
  NAND U10122 ( .A(n7950), .B(n7951), .Z(y[449]) );
  NAND U10123 ( .A(n7702), .B(m[449]), .Z(n7951) );
  NAND U10124 ( .A(n7703), .B(creg[449]), .Z(n7950) );
  NAND U10125 ( .A(n7952), .B(n7953), .Z(y[448]) );
  NAND U10126 ( .A(n7702), .B(m[448]), .Z(n7953) );
  NAND U10127 ( .A(n7703), .B(creg[448]), .Z(n7952) );
  NAND U10128 ( .A(n7954), .B(n7955), .Z(y[447]) );
  NAND U10129 ( .A(n7702), .B(m[447]), .Z(n7955) );
  NAND U10130 ( .A(n7703), .B(creg[447]), .Z(n7954) );
  NAND U10131 ( .A(n7956), .B(n7957), .Z(y[446]) );
  NAND U10132 ( .A(n7702), .B(m[446]), .Z(n7957) );
  NAND U10133 ( .A(n7703), .B(creg[446]), .Z(n7956) );
  NAND U10134 ( .A(n7958), .B(n7959), .Z(y[445]) );
  NAND U10135 ( .A(n7702), .B(m[445]), .Z(n7959) );
  NAND U10136 ( .A(n7703), .B(creg[445]), .Z(n7958) );
  NAND U10137 ( .A(n7960), .B(n7961), .Z(y[444]) );
  NAND U10138 ( .A(n7702), .B(m[444]), .Z(n7961) );
  NAND U10139 ( .A(n7703), .B(creg[444]), .Z(n7960) );
  NAND U10140 ( .A(n7962), .B(n7963), .Z(y[443]) );
  NAND U10141 ( .A(n7702), .B(m[443]), .Z(n7963) );
  NAND U10142 ( .A(n7703), .B(creg[443]), .Z(n7962) );
  NAND U10143 ( .A(n7964), .B(n7965), .Z(y[442]) );
  NAND U10144 ( .A(n7702), .B(m[442]), .Z(n7965) );
  NAND U10145 ( .A(n7703), .B(creg[442]), .Z(n7964) );
  NAND U10146 ( .A(n7966), .B(n7967), .Z(y[441]) );
  NAND U10147 ( .A(n7702), .B(m[441]), .Z(n7967) );
  NAND U10148 ( .A(n7703), .B(creg[441]), .Z(n7966) );
  NAND U10149 ( .A(n7968), .B(n7969), .Z(y[440]) );
  NAND U10150 ( .A(n7702), .B(m[440]), .Z(n7969) );
  NAND U10151 ( .A(n7703), .B(creg[440]), .Z(n7968) );
  NAND U10152 ( .A(n7970), .B(n7971), .Z(y[43]) );
  NAND U10153 ( .A(n7702), .B(m[43]), .Z(n7971) );
  NAND U10154 ( .A(n7703), .B(creg[43]), .Z(n7970) );
  NAND U10155 ( .A(n7972), .B(n7973), .Z(y[439]) );
  NAND U10156 ( .A(n7702), .B(m[439]), .Z(n7973) );
  NAND U10157 ( .A(n7703), .B(creg[439]), .Z(n7972) );
  NAND U10158 ( .A(n7974), .B(n7975), .Z(y[438]) );
  NAND U10159 ( .A(n7702), .B(m[438]), .Z(n7975) );
  NAND U10160 ( .A(n7703), .B(creg[438]), .Z(n7974) );
  NAND U10161 ( .A(n7976), .B(n7977), .Z(y[437]) );
  NAND U10162 ( .A(n7702), .B(m[437]), .Z(n7977) );
  NAND U10163 ( .A(n7703), .B(creg[437]), .Z(n7976) );
  NAND U10164 ( .A(n7978), .B(n7979), .Z(y[436]) );
  NAND U10165 ( .A(n7702), .B(m[436]), .Z(n7979) );
  NAND U10166 ( .A(n7703), .B(creg[436]), .Z(n7978) );
  NAND U10167 ( .A(n7980), .B(n7981), .Z(y[435]) );
  NAND U10168 ( .A(n7702), .B(m[435]), .Z(n7981) );
  NAND U10169 ( .A(n7703), .B(creg[435]), .Z(n7980) );
  NAND U10170 ( .A(n7982), .B(n7983), .Z(y[434]) );
  NAND U10171 ( .A(n7702), .B(m[434]), .Z(n7983) );
  NAND U10172 ( .A(n7703), .B(creg[434]), .Z(n7982) );
  NAND U10173 ( .A(n7984), .B(n7985), .Z(y[433]) );
  NAND U10174 ( .A(n7702), .B(m[433]), .Z(n7985) );
  NAND U10175 ( .A(n7703), .B(creg[433]), .Z(n7984) );
  NAND U10176 ( .A(n7986), .B(n7987), .Z(y[432]) );
  NAND U10177 ( .A(n7702), .B(m[432]), .Z(n7987) );
  NAND U10178 ( .A(n7703), .B(creg[432]), .Z(n7986) );
  NAND U10179 ( .A(n7988), .B(n7989), .Z(y[431]) );
  NAND U10180 ( .A(n7702), .B(m[431]), .Z(n7989) );
  NAND U10181 ( .A(n7703), .B(creg[431]), .Z(n7988) );
  NAND U10182 ( .A(n7990), .B(n7991), .Z(y[430]) );
  NAND U10183 ( .A(n7702), .B(m[430]), .Z(n7991) );
  NAND U10184 ( .A(n7703), .B(creg[430]), .Z(n7990) );
  NAND U10185 ( .A(n7992), .B(n7993), .Z(y[42]) );
  NAND U10186 ( .A(n7702), .B(m[42]), .Z(n7993) );
  NAND U10187 ( .A(n7703), .B(creg[42]), .Z(n7992) );
  NAND U10188 ( .A(n7994), .B(n7995), .Z(y[429]) );
  NAND U10189 ( .A(n7702), .B(m[429]), .Z(n7995) );
  NAND U10190 ( .A(n7703), .B(creg[429]), .Z(n7994) );
  NAND U10191 ( .A(n7996), .B(n7997), .Z(y[428]) );
  NAND U10192 ( .A(n7702), .B(m[428]), .Z(n7997) );
  NAND U10193 ( .A(n7703), .B(creg[428]), .Z(n7996) );
  NAND U10194 ( .A(n7998), .B(n7999), .Z(y[427]) );
  NAND U10195 ( .A(n7702), .B(m[427]), .Z(n7999) );
  NAND U10196 ( .A(n7703), .B(creg[427]), .Z(n7998) );
  NAND U10197 ( .A(n8000), .B(n8001), .Z(y[426]) );
  NAND U10198 ( .A(n7702), .B(m[426]), .Z(n8001) );
  NAND U10199 ( .A(n7703), .B(creg[426]), .Z(n8000) );
  NAND U10200 ( .A(n8002), .B(n8003), .Z(y[425]) );
  NAND U10201 ( .A(n7702), .B(m[425]), .Z(n8003) );
  NAND U10202 ( .A(n7703), .B(creg[425]), .Z(n8002) );
  NAND U10203 ( .A(n8004), .B(n8005), .Z(y[424]) );
  NAND U10204 ( .A(n7702), .B(m[424]), .Z(n8005) );
  NAND U10205 ( .A(n7703), .B(creg[424]), .Z(n8004) );
  NAND U10206 ( .A(n8006), .B(n8007), .Z(y[423]) );
  NAND U10207 ( .A(n7702), .B(m[423]), .Z(n8007) );
  NAND U10208 ( .A(n7703), .B(creg[423]), .Z(n8006) );
  NAND U10209 ( .A(n8008), .B(n8009), .Z(y[422]) );
  NAND U10210 ( .A(n7702), .B(m[422]), .Z(n8009) );
  NAND U10211 ( .A(n7703), .B(creg[422]), .Z(n8008) );
  NAND U10212 ( .A(n8010), .B(n8011), .Z(y[421]) );
  NAND U10213 ( .A(n7702), .B(m[421]), .Z(n8011) );
  NAND U10214 ( .A(n7703), .B(creg[421]), .Z(n8010) );
  NAND U10215 ( .A(n8012), .B(n8013), .Z(y[420]) );
  NAND U10216 ( .A(n7702), .B(m[420]), .Z(n8013) );
  NAND U10217 ( .A(n7703), .B(creg[420]), .Z(n8012) );
  NAND U10218 ( .A(n8014), .B(n8015), .Z(y[41]) );
  NAND U10219 ( .A(n7702), .B(m[41]), .Z(n8015) );
  NAND U10220 ( .A(n7703), .B(creg[41]), .Z(n8014) );
  NAND U10221 ( .A(n8016), .B(n8017), .Z(y[419]) );
  NAND U10222 ( .A(n7702), .B(m[419]), .Z(n8017) );
  NAND U10223 ( .A(n7703), .B(creg[419]), .Z(n8016) );
  NAND U10224 ( .A(n8018), .B(n8019), .Z(y[418]) );
  NAND U10225 ( .A(n7702), .B(m[418]), .Z(n8019) );
  NAND U10226 ( .A(n7703), .B(creg[418]), .Z(n8018) );
  NAND U10227 ( .A(n8020), .B(n8021), .Z(y[417]) );
  NAND U10228 ( .A(n7702), .B(m[417]), .Z(n8021) );
  NAND U10229 ( .A(n7703), .B(creg[417]), .Z(n8020) );
  NAND U10230 ( .A(n8022), .B(n8023), .Z(y[416]) );
  NAND U10231 ( .A(n7702), .B(m[416]), .Z(n8023) );
  NAND U10232 ( .A(n7703), .B(creg[416]), .Z(n8022) );
  NAND U10233 ( .A(n8024), .B(n8025), .Z(y[415]) );
  NAND U10234 ( .A(n7702), .B(m[415]), .Z(n8025) );
  NAND U10235 ( .A(n7703), .B(creg[415]), .Z(n8024) );
  NAND U10236 ( .A(n8026), .B(n8027), .Z(y[414]) );
  NAND U10237 ( .A(n7702), .B(m[414]), .Z(n8027) );
  NAND U10238 ( .A(n7703), .B(creg[414]), .Z(n8026) );
  NAND U10239 ( .A(n8028), .B(n8029), .Z(y[413]) );
  NAND U10240 ( .A(n7702), .B(m[413]), .Z(n8029) );
  NAND U10241 ( .A(n7703), .B(creg[413]), .Z(n8028) );
  NAND U10242 ( .A(n8030), .B(n8031), .Z(y[412]) );
  NAND U10243 ( .A(n7702), .B(m[412]), .Z(n8031) );
  NAND U10244 ( .A(n7703), .B(creg[412]), .Z(n8030) );
  NAND U10245 ( .A(n8032), .B(n8033), .Z(y[411]) );
  NAND U10246 ( .A(n7702), .B(m[411]), .Z(n8033) );
  NAND U10247 ( .A(n7703), .B(creg[411]), .Z(n8032) );
  NAND U10248 ( .A(n8034), .B(n8035), .Z(y[410]) );
  NAND U10249 ( .A(n7702), .B(m[410]), .Z(n8035) );
  NAND U10250 ( .A(n7703), .B(creg[410]), .Z(n8034) );
  NAND U10251 ( .A(n8036), .B(n8037), .Z(y[40]) );
  NAND U10252 ( .A(n7702), .B(m[40]), .Z(n8037) );
  NAND U10253 ( .A(n7703), .B(creg[40]), .Z(n8036) );
  NAND U10254 ( .A(n8038), .B(n8039), .Z(y[409]) );
  NAND U10255 ( .A(n7702), .B(m[409]), .Z(n8039) );
  NAND U10256 ( .A(n7703), .B(creg[409]), .Z(n8038) );
  NAND U10257 ( .A(n8040), .B(n8041), .Z(y[408]) );
  NAND U10258 ( .A(n7702), .B(m[408]), .Z(n8041) );
  NAND U10259 ( .A(n7703), .B(creg[408]), .Z(n8040) );
  NAND U10260 ( .A(n8042), .B(n8043), .Z(y[407]) );
  NAND U10261 ( .A(n7702), .B(m[407]), .Z(n8043) );
  NAND U10262 ( .A(n7703), .B(creg[407]), .Z(n8042) );
  NAND U10263 ( .A(n8044), .B(n8045), .Z(y[406]) );
  NAND U10264 ( .A(n7702), .B(m[406]), .Z(n8045) );
  NAND U10265 ( .A(n7703), .B(creg[406]), .Z(n8044) );
  NAND U10266 ( .A(n8046), .B(n8047), .Z(y[405]) );
  NAND U10267 ( .A(n7702), .B(m[405]), .Z(n8047) );
  NAND U10268 ( .A(n7703), .B(creg[405]), .Z(n8046) );
  NAND U10269 ( .A(n8048), .B(n8049), .Z(y[404]) );
  NAND U10270 ( .A(n7702), .B(m[404]), .Z(n8049) );
  NAND U10271 ( .A(n7703), .B(creg[404]), .Z(n8048) );
  NAND U10272 ( .A(n8050), .B(n8051), .Z(y[403]) );
  NAND U10273 ( .A(n7702), .B(m[403]), .Z(n8051) );
  NAND U10274 ( .A(n7703), .B(creg[403]), .Z(n8050) );
  NAND U10275 ( .A(n8052), .B(n8053), .Z(y[402]) );
  NAND U10276 ( .A(n7702), .B(m[402]), .Z(n8053) );
  NAND U10277 ( .A(n7703), .B(creg[402]), .Z(n8052) );
  NAND U10278 ( .A(n8054), .B(n8055), .Z(y[401]) );
  NAND U10279 ( .A(n7702), .B(m[401]), .Z(n8055) );
  NAND U10280 ( .A(n7703), .B(creg[401]), .Z(n8054) );
  NAND U10281 ( .A(n8056), .B(n8057), .Z(y[400]) );
  NAND U10282 ( .A(n7702), .B(m[400]), .Z(n8057) );
  NAND U10283 ( .A(n7703), .B(creg[400]), .Z(n8056) );
  NAND U10284 ( .A(n8058), .B(n8059), .Z(y[3]) );
  NAND U10285 ( .A(n7702), .B(m[3]), .Z(n8059) );
  NAND U10286 ( .A(n7703), .B(creg[3]), .Z(n8058) );
  NAND U10287 ( .A(n8060), .B(n8061), .Z(y[39]) );
  NAND U10288 ( .A(n7702), .B(m[39]), .Z(n8061) );
  NAND U10289 ( .A(n7703), .B(creg[39]), .Z(n8060) );
  NAND U10290 ( .A(n8062), .B(n8063), .Z(y[399]) );
  NAND U10291 ( .A(n7702), .B(m[399]), .Z(n8063) );
  NAND U10292 ( .A(n7703), .B(creg[399]), .Z(n8062) );
  NAND U10293 ( .A(n8064), .B(n8065), .Z(y[398]) );
  NAND U10294 ( .A(n7702), .B(m[398]), .Z(n8065) );
  NAND U10295 ( .A(n7703), .B(creg[398]), .Z(n8064) );
  NAND U10296 ( .A(n8066), .B(n8067), .Z(y[397]) );
  NAND U10297 ( .A(n7702), .B(m[397]), .Z(n8067) );
  NAND U10298 ( .A(n7703), .B(creg[397]), .Z(n8066) );
  NAND U10299 ( .A(n8068), .B(n8069), .Z(y[396]) );
  NAND U10300 ( .A(n7702), .B(m[396]), .Z(n8069) );
  NAND U10301 ( .A(n7703), .B(creg[396]), .Z(n8068) );
  NAND U10302 ( .A(n8070), .B(n8071), .Z(y[395]) );
  NAND U10303 ( .A(n7702), .B(m[395]), .Z(n8071) );
  NAND U10304 ( .A(n7703), .B(creg[395]), .Z(n8070) );
  NAND U10305 ( .A(n8072), .B(n8073), .Z(y[394]) );
  NAND U10306 ( .A(n7702), .B(m[394]), .Z(n8073) );
  NAND U10307 ( .A(n7703), .B(creg[394]), .Z(n8072) );
  NAND U10308 ( .A(n8074), .B(n8075), .Z(y[393]) );
  NAND U10309 ( .A(n7702), .B(m[393]), .Z(n8075) );
  NAND U10310 ( .A(n7703), .B(creg[393]), .Z(n8074) );
  NAND U10311 ( .A(n8076), .B(n8077), .Z(y[392]) );
  NAND U10312 ( .A(n7702), .B(m[392]), .Z(n8077) );
  NAND U10313 ( .A(n7703), .B(creg[392]), .Z(n8076) );
  NAND U10314 ( .A(n8078), .B(n8079), .Z(y[391]) );
  NAND U10315 ( .A(n7702), .B(m[391]), .Z(n8079) );
  NAND U10316 ( .A(n7703), .B(creg[391]), .Z(n8078) );
  NAND U10317 ( .A(n8080), .B(n8081), .Z(y[390]) );
  NAND U10318 ( .A(n7702), .B(m[390]), .Z(n8081) );
  NAND U10319 ( .A(n7703), .B(creg[390]), .Z(n8080) );
  NAND U10320 ( .A(n8082), .B(n8083), .Z(y[38]) );
  NAND U10321 ( .A(n7702), .B(m[38]), .Z(n8083) );
  NAND U10322 ( .A(n7703), .B(creg[38]), .Z(n8082) );
  NAND U10323 ( .A(n8084), .B(n8085), .Z(y[389]) );
  NAND U10324 ( .A(n7702), .B(m[389]), .Z(n8085) );
  NAND U10325 ( .A(n7703), .B(creg[389]), .Z(n8084) );
  NAND U10326 ( .A(n8086), .B(n8087), .Z(y[388]) );
  NAND U10327 ( .A(n7702), .B(m[388]), .Z(n8087) );
  NAND U10328 ( .A(n7703), .B(creg[388]), .Z(n8086) );
  NAND U10329 ( .A(n8088), .B(n8089), .Z(y[387]) );
  NAND U10330 ( .A(n7702), .B(m[387]), .Z(n8089) );
  NAND U10331 ( .A(n7703), .B(creg[387]), .Z(n8088) );
  NAND U10332 ( .A(n8090), .B(n8091), .Z(y[386]) );
  NAND U10333 ( .A(n7702), .B(m[386]), .Z(n8091) );
  NAND U10334 ( .A(n7703), .B(creg[386]), .Z(n8090) );
  NAND U10335 ( .A(n8092), .B(n8093), .Z(y[385]) );
  NAND U10336 ( .A(n7702), .B(m[385]), .Z(n8093) );
  NAND U10337 ( .A(n7703), .B(creg[385]), .Z(n8092) );
  NAND U10338 ( .A(n8094), .B(n8095), .Z(y[384]) );
  NAND U10339 ( .A(n7702), .B(m[384]), .Z(n8095) );
  NAND U10340 ( .A(n7703), .B(creg[384]), .Z(n8094) );
  NAND U10341 ( .A(n8096), .B(n8097), .Z(y[383]) );
  NAND U10342 ( .A(n7702), .B(m[383]), .Z(n8097) );
  NAND U10343 ( .A(n7703), .B(creg[383]), .Z(n8096) );
  NAND U10344 ( .A(n8098), .B(n8099), .Z(y[382]) );
  NAND U10345 ( .A(n7702), .B(m[382]), .Z(n8099) );
  NAND U10346 ( .A(n7703), .B(creg[382]), .Z(n8098) );
  NAND U10347 ( .A(n8100), .B(n8101), .Z(y[381]) );
  NAND U10348 ( .A(n7702), .B(m[381]), .Z(n8101) );
  NAND U10349 ( .A(n7703), .B(creg[381]), .Z(n8100) );
  NAND U10350 ( .A(n8102), .B(n8103), .Z(y[380]) );
  NAND U10351 ( .A(n7702), .B(m[380]), .Z(n8103) );
  NAND U10352 ( .A(n7703), .B(creg[380]), .Z(n8102) );
  NAND U10353 ( .A(n8104), .B(n8105), .Z(y[37]) );
  NAND U10354 ( .A(n7702), .B(m[37]), .Z(n8105) );
  NAND U10355 ( .A(n7703), .B(creg[37]), .Z(n8104) );
  NAND U10356 ( .A(n8106), .B(n8107), .Z(y[379]) );
  NAND U10357 ( .A(n7702), .B(m[379]), .Z(n8107) );
  NAND U10358 ( .A(n7703), .B(creg[379]), .Z(n8106) );
  NAND U10359 ( .A(n8108), .B(n8109), .Z(y[378]) );
  NAND U10360 ( .A(n7702), .B(m[378]), .Z(n8109) );
  NAND U10361 ( .A(n7703), .B(creg[378]), .Z(n8108) );
  NAND U10362 ( .A(n8110), .B(n8111), .Z(y[377]) );
  NAND U10363 ( .A(n7702), .B(m[377]), .Z(n8111) );
  NAND U10364 ( .A(n7703), .B(creg[377]), .Z(n8110) );
  NAND U10365 ( .A(n8112), .B(n8113), .Z(y[376]) );
  NAND U10366 ( .A(n7702), .B(m[376]), .Z(n8113) );
  NAND U10367 ( .A(n7703), .B(creg[376]), .Z(n8112) );
  NAND U10368 ( .A(n8114), .B(n8115), .Z(y[375]) );
  NAND U10369 ( .A(n7702), .B(m[375]), .Z(n8115) );
  NAND U10370 ( .A(n7703), .B(creg[375]), .Z(n8114) );
  NAND U10371 ( .A(n8116), .B(n8117), .Z(y[374]) );
  NAND U10372 ( .A(n7702), .B(m[374]), .Z(n8117) );
  NAND U10373 ( .A(n7703), .B(creg[374]), .Z(n8116) );
  NAND U10374 ( .A(n8118), .B(n8119), .Z(y[373]) );
  NAND U10375 ( .A(n7702), .B(m[373]), .Z(n8119) );
  NAND U10376 ( .A(n7703), .B(creg[373]), .Z(n8118) );
  NAND U10377 ( .A(n8120), .B(n8121), .Z(y[372]) );
  NAND U10378 ( .A(n7702), .B(m[372]), .Z(n8121) );
  NAND U10379 ( .A(n7703), .B(creg[372]), .Z(n8120) );
  NAND U10380 ( .A(n8122), .B(n8123), .Z(y[371]) );
  NAND U10381 ( .A(n7702), .B(m[371]), .Z(n8123) );
  NAND U10382 ( .A(n7703), .B(creg[371]), .Z(n8122) );
  NAND U10383 ( .A(n8124), .B(n8125), .Z(y[370]) );
  NAND U10384 ( .A(n7702), .B(m[370]), .Z(n8125) );
  NAND U10385 ( .A(n7703), .B(creg[370]), .Z(n8124) );
  NAND U10386 ( .A(n8126), .B(n8127), .Z(y[36]) );
  NAND U10387 ( .A(n7702), .B(m[36]), .Z(n8127) );
  NAND U10388 ( .A(n7703), .B(creg[36]), .Z(n8126) );
  NAND U10389 ( .A(n8128), .B(n8129), .Z(y[369]) );
  NAND U10390 ( .A(n7702), .B(m[369]), .Z(n8129) );
  NAND U10391 ( .A(n7703), .B(creg[369]), .Z(n8128) );
  NAND U10392 ( .A(n8130), .B(n8131), .Z(y[368]) );
  NAND U10393 ( .A(n7702), .B(m[368]), .Z(n8131) );
  NAND U10394 ( .A(n7703), .B(creg[368]), .Z(n8130) );
  NAND U10395 ( .A(n8132), .B(n8133), .Z(y[367]) );
  NAND U10396 ( .A(n7702), .B(m[367]), .Z(n8133) );
  NAND U10397 ( .A(n7703), .B(creg[367]), .Z(n8132) );
  NAND U10398 ( .A(n8134), .B(n8135), .Z(y[366]) );
  NAND U10399 ( .A(n7702), .B(m[366]), .Z(n8135) );
  NAND U10400 ( .A(n7703), .B(creg[366]), .Z(n8134) );
  NAND U10401 ( .A(n8136), .B(n8137), .Z(y[365]) );
  NAND U10402 ( .A(n7702), .B(m[365]), .Z(n8137) );
  NAND U10403 ( .A(n7703), .B(creg[365]), .Z(n8136) );
  NAND U10404 ( .A(n8138), .B(n8139), .Z(y[364]) );
  NAND U10405 ( .A(n7702), .B(m[364]), .Z(n8139) );
  NAND U10406 ( .A(n7703), .B(creg[364]), .Z(n8138) );
  NAND U10407 ( .A(n8140), .B(n8141), .Z(y[363]) );
  NAND U10408 ( .A(n7702), .B(m[363]), .Z(n8141) );
  NAND U10409 ( .A(n7703), .B(creg[363]), .Z(n8140) );
  NAND U10410 ( .A(n8142), .B(n8143), .Z(y[362]) );
  NAND U10411 ( .A(n7702), .B(m[362]), .Z(n8143) );
  NAND U10412 ( .A(n7703), .B(creg[362]), .Z(n8142) );
  NAND U10413 ( .A(n8144), .B(n8145), .Z(y[361]) );
  NAND U10414 ( .A(n7702), .B(m[361]), .Z(n8145) );
  NAND U10415 ( .A(n7703), .B(creg[361]), .Z(n8144) );
  NAND U10416 ( .A(n8146), .B(n8147), .Z(y[360]) );
  NAND U10417 ( .A(n7702), .B(m[360]), .Z(n8147) );
  NAND U10418 ( .A(n7703), .B(creg[360]), .Z(n8146) );
  NAND U10419 ( .A(n8148), .B(n8149), .Z(y[35]) );
  NAND U10420 ( .A(n7702), .B(m[35]), .Z(n8149) );
  NAND U10421 ( .A(n7703), .B(creg[35]), .Z(n8148) );
  NAND U10422 ( .A(n8150), .B(n8151), .Z(y[359]) );
  NAND U10423 ( .A(n7702), .B(m[359]), .Z(n8151) );
  NAND U10424 ( .A(n7703), .B(creg[359]), .Z(n8150) );
  NAND U10425 ( .A(n8152), .B(n8153), .Z(y[358]) );
  NAND U10426 ( .A(n7702), .B(m[358]), .Z(n8153) );
  NAND U10427 ( .A(n7703), .B(creg[358]), .Z(n8152) );
  NAND U10428 ( .A(n8154), .B(n8155), .Z(y[357]) );
  NAND U10429 ( .A(n7702), .B(m[357]), .Z(n8155) );
  NAND U10430 ( .A(n7703), .B(creg[357]), .Z(n8154) );
  NAND U10431 ( .A(n8156), .B(n8157), .Z(y[356]) );
  NAND U10432 ( .A(n7702), .B(m[356]), .Z(n8157) );
  NAND U10433 ( .A(n7703), .B(creg[356]), .Z(n8156) );
  NAND U10434 ( .A(n8158), .B(n8159), .Z(y[355]) );
  NAND U10435 ( .A(n7702), .B(m[355]), .Z(n8159) );
  NAND U10436 ( .A(n7703), .B(creg[355]), .Z(n8158) );
  NAND U10437 ( .A(n8160), .B(n8161), .Z(y[354]) );
  NAND U10438 ( .A(n7702), .B(m[354]), .Z(n8161) );
  NAND U10439 ( .A(n7703), .B(creg[354]), .Z(n8160) );
  NAND U10440 ( .A(n8162), .B(n8163), .Z(y[353]) );
  NAND U10441 ( .A(n7702), .B(m[353]), .Z(n8163) );
  NAND U10442 ( .A(n7703), .B(creg[353]), .Z(n8162) );
  NAND U10443 ( .A(n8164), .B(n8165), .Z(y[352]) );
  NAND U10444 ( .A(n7702), .B(m[352]), .Z(n8165) );
  NAND U10445 ( .A(n7703), .B(creg[352]), .Z(n8164) );
  NAND U10446 ( .A(n8166), .B(n8167), .Z(y[351]) );
  NAND U10447 ( .A(n7702), .B(m[351]), .Z(n8167) );
  NAND U10448 ( .A(n7703), .B(creg[351]), .Z(n8166) );
  NAND U10449 ( .A(n8168), .B(n8169), .Z(y[350]) );
  NAND U10450 ( .A(n7702), .B(m[350]), .Z(n8169) );
  NAND U10451 ( .A(n7703), .B(creg[350]), .Z(n8168) );
  NAND U10452 ( .A(n8170), .B(n8171), .Z(y[34]) );
  NAND U10453 ( .A(n7702), .B(m[34]), .Z(n8171) );
  NAND U10454 ( .A(n7703), .B(creg[34]), .Z(n8170) );
  NAND U10455 ( .A(n8172), .B(n8173), .Z(y[349]) );
  NAND U10456 ( .A(n7702), .B(m[349]), .Z(n8173) );
  NAND U10457 ( .A(n7703), .B(creg[349]), .Z(n8172) );
  NAND U10458 ( .A(n8174), .B(n8175), .Z(y[348]) );
  NAND U10459 ( .A(n7702), .B(m[348]), .Z(n8175) );
  NAND U10460 ( .A(n7703), .B(creg[348]), .Z(n8174) );
  NAND U10461 ( .A(n8176), .B(n8177), .Z(y[347]) );
  NAND U10462 ( .A(n7702), .B(m[347]), .Z(n8177) );
  NAND U10463 ( .A(n7703), .B(creg[347]), .Z(n8176) );
  NAND U10464 ( .A(n8178), .B(n8179), .Z(y[346]) );
  NAND U10465 ( .A(n7702), .B(m[346]), .Z(n8179) );
  NAND U10466 ( .A(n7703), .B(creg[346]), .Z(n8178) );
  NAND U10467 ( .A(n8180), .B(n8181), .Z(y[345]) );
  NAND U10468 ( .A(n7702), .B(m[345]), .Z(n8181) );
  NAND U10469 ( .A(n7703), .B(creg[345]), .Z(n8180) );
  NAND U10470 ( .A(n8182), .B(n8183), .Z(y[344]) );
  NAND U10471 ( .A(n7702), .B(m[344]), .Z(n8183) );
  NAND U10472 ( .A(n7703), .B(creg[344]), .Z(n8182) );
  NAND U10473 ( .A(n8184), .B(n8185), .Z(y[343]) );
  NAND U10474 ( .A(n7702), .B(m[343]), .Z(n8185) );
  NAND U10475 ( .A(n7703), .B(creg[343]), .Z(n8184) );
  NAND U10476 ( .A(n8186), .B(n8187), .Z(y[342]) );
  NAND U10477 ( .A(n7702), .B(m[342]), .Z(n8187) );
  NAND U10478 ( .A(n7703), .B(creg[342]), .Z(n8186) );
  NAND U10479 ( .A(n8188), .B(n8189), .Z(y[341]) );
  NAND U10480 ( .A(n7702), .B(m[341]), .Z(n8189) );
  NAND U10481 ( .A(n7703), .B(creg[341]), .Z(n8188) );
  NAND U10482 ( .A(n8190), .B(n8191), .Z(y[340]) );
  NAND U10483 ( .A(n7702), .B(m[340]), .Z(n8191) );
  NAND U10484 ( .A(n7703), .B(creg[340]), .Z(n8190) );
  NAND U10485 ( .A(n8192), .B(n8193), .Z(y[33]) );
  NAND U10486 ( .A(n7702), .B(m[33]), .Z(n8193) );
  NAND U10487 ( .A(n7703), .B(creg[33]), .Z(n8192) );
  NAND U10488 ( .A(n8194), .B(n8195), .Z(y[339]) );
  NAND U10489 ( .A(n7702), .B(m[339]), .Z(n8195) );
  NAND U10490 ( .A(n7703), .B(creg[339]), .Z(n8194) );
  NAND U10491 ( .A(n8196), .B(n8197), .Z(y[338]) );
  NAND U10492 ( .A(n7702), .B(m[338]), .Z(n8197) );
  NAND U10493 ( .A(n7703), .B(creg[338]), .Z(n8196) );
  NAND U10494 ( .A(n8198), .B(n8199), .Z(y[337]) );
  NAND U10495 ( .A(n7702), .B(m[337]), .Z(n8199) );
  NAND U10496 ( .A(n7703), .B(creg[337]), .Z(n8198) );
  NAND U10497 ( .A(n8200), .B(n8201), .Z(y[336]) );
  NAND U10498 ( .A(n7702), .B(m[336]), .Z(n8201) );
  NAND U10499 ( .A(n7703), .B(creg[336]), .Z(n8200) );
  NAND U10500 ( .A(n8202), .B(n8203), .Z(y[335]) );
  NAND U10501 ( .A(n7702), .B(m[335]), .Z(n8203) );
  NAND U10502 ( .A(n7703), .B(creg[335]), .Z(n8202) );
  NAND U10503 ( .A(n8204), .B(n8205), .Z(y[334]) );
  NAND U10504 ( .A(n7702), .B(m[334]), .Z(n8205) );
  NAND U10505 ( .A(n7703), .B(creg[334]), .Z(n8204) );
  NAND U10506 ( .A(n8206), .B(n8207), .Z(y[333]) );
  NAND U10507 ( .A(n7702), .B(m[333]), .Z(n8207) );
  NAND U10508 ( .A(n7703), .B(creg[333]), .Z(n8206) );
  NAND U10509 ( .A(n8208), .B(n8209), .Z(y[332]) );
  NAND U10510 ( .A(n7702), .B(m[332]), .Z(n8209) );
  NAND U10511 ( .A(n7703), .B(creg[332]), .Z(n8208) );
  NAND U10512 ( .A(n8210), .B(n8211), .Z(y[331]) );
  NAND U10513 ( .A(n7702), .B(m[331]), .Z(n8211) );
  NAND U10514 ( .A(n7703), .B(creg[331]), .Z(n8210) );
  NAND U10515 ( .A(n8212), .B(n8213), .Z(y[330]) );
  NAND U10516 ( .A(n7702), .B(m[330]), .Z(n8213) );
  NAND U10517 ( .A(n7703), .B(creg[330]), .Z(n8212) );
  NAND U10518 ( .A(n8214), .B(n8215), .Z(y[32]) );
  NAND U10519 ( .A(n7702), .B(m[32]), .Z(n8215) );
  NAND U10520 ( .A(n7703), .B(creg[32]), .Z(n8214) );
  NAND U10521 ( .A(n8216), .B(n8217), .Z(y[329]) );
  NAND U10522 ( .A(n7702), .B(m[329]), .Z(n8217) );
  NAND U10523 ( .A(n7703), .B(creg[329]), .Z(n8216) );
  NAND U10524 ( .A(n8218), .B(n8219), .Z(y[328]) );
  NAND U10525 ( .A(n7702), .B(m[328]), .Z(n8219) );
  NAND U10526 ( .A(n7703), .B(creg[328]), .Z(n8218) );
  NAND U10527 ( .A(n8220), .B(n8221), .Z(y[327]) );
  NAND U10528 ( .A(n7702), .B(m[327]), .Z(n8221) );
  NAND U10529 ( .A(n7703), .B(creg[327]), .Z(n8220) );
  NAND U10530 ( .A(n8222), .B(n8223), .Z(y[326]) );
  NAND U10531 ( .A(n7702), .B(m[326]), .Z(n8223) );
  NAND U10532 ( .A(n7703), .B(creg[326]), .Z(n8222) );
  NAND U10533 ( .A(n8224), .B(n8225), .Z(y[325]) );
  NAND U10534 ( .A(n7702), .B(m[325]), .Z(n8225) );
  NAND U10535 ( .A(n7703), .B(creg[325]), .Z(n8224) );
  NAND U10536 ( .A(n8226), .B(n8227), .Z(y[324]) );
  NAND U10537 ( .A(n7702), .B(m[324]), .Z(n8227) );
  NAND U10538 ( .A(n7703), .B(creg[324]), .Z(n8226) );
  NAND U10539 ( .A(n8228), .B(n8229), .Z(y[323]) );
  NAND U10540 ( .A(n7702), .B(m[323]), .Z(n8229) );
  NAND U10541 ( .A(n7703), .B(creg[323]), .Z(n8228) );
  NAND U10542 ( .A(n8230), .B(n8231), .Z(y[322]) );
  NAND U10543 ( .A(n7702), .B(m[322]), .Z(n8231) );
  NAND U10544 ( .A(n7703), .B(creg[322]), .Z(n8230) );
  NAND U10545 ( .A(n8232), .B(n8233), .Z(y[321]) );
  NAND U10546 ( .A(n7702), .B(m[321]), .Z(n8233) );
  NAND U10547 ( .A(n7703), .B(creg[321]), .Z(n8232) );
  NAND U10548 ( .A(n8234), .B(n8235), .Z(y[320]) );
  NAND U10549 ( .A(n7702), .B(m[320]), .Z(n8235) );
  NAND U10550 ( .A(n7703), .B(creg[320]), .Z(n8234) );
  NAND U10551 ( .A(n8236), .B(n8237), .Z(y[31]) );
  NAND U10552 ( .A(n7702), .B(m[31]), .Z(n8237) );
  NAND U10553 ( .A(n7703), .B(creg[31]), .Z(n8236) );
  NAND U10554 ( .A(n8238), .B(n8239), .Z(y[319]) );
  NAND U10555 ( .A(n7702), .B(m[319]), .Z(n8239) );
  NAND U10556 ( .A(n7703), .B(creg[319]), .Z(n8238) );
  NAND U10557 ( .A(n8240), .B(n8241), .Z(y[318]) );
  NAND U10558 ( .A(n7702), .B(m[318]), .Z(n8241) );
  NAND U10559 ( .A(n7703), .B(creg[318]), .Z(n8240) );
  NAND U10560 ( .A(n8242), .B(n8243), .Z(y[317]) );
  NAND U10561 ( .A(n7702), .B(m[317]), .Z(n8243) );
  NAND U10562 ( .A(n7703), .B(creg[317]), .Z(n8242) );
  NAND U10563 ( .A(n8244), .B(n8245), .Z(y[316]) );
  NAND U10564 ( .A(n7702), .B(m[316]), .Z(n8245) );
  NAND U10565 ( .A(n7703), .B(creg[316]), .Z(n8244) );
  NAND U10566 ( .A(n8246), .B(n8247), .Z(y[315]) );
  NAND U10567 ( .A(n7702), .B(m[315]), .Z(n8247) );
  NAND U10568 ( .A(n7703), .B(creg[315]), .Z(n8246) );
  NAND U10569 ( .A(n8248), .B(n8249), .Z(y[314]) );
  NAND U10570 ( .A(n7702), .B(m[314]), .Z(n8249) );
  NAND U10571 ( .A(n7703), .B(creg[314]), .Z(n8248) );
  NAND U10572 ( .A(n8250), .B(n8251), .Z(y[313]) );
  NAND U10573 ( .A(n7702), .B(m[313]), .Z(n8251) );
  NAND U10574 ( .A(n7703), .B(creg[313]), .Z(n8250) );
  NAND U10575 ( .A(n8252), .B(n8253), .Z(y[312]) );
  NAND U10576 ( .A(n7702), .B(m[312]), .Z(n8253) );
  NAND U10577 ( .A(n7703), .B(creg[312]), .Z(n8252) );
  NAND U10578 ( .A(n8254), .B(n8255), .Z(y[311]) );
  NAND U10579 ( .A(n7702), .B(m[311]), .Z(n8255) );
  NAND U10580 ( .A(n7703), .B(creg[311]), .Z(n8254) );
  NAND U10581 ( .A(n8256), .B(n8257), .Z(y[310]) );
  NAND U10582 ( .A(n7702), .B(m[310]), .Z(n8257) );
  NAND U10583 ( .A(n7703), .B(creg[310]), .Z(n8256) );
  NAND U10584 ( .A(n8258), .B(n8259), .Z(y[30]) );
  NAND U10585 ( .A(n7702), .B(m[30]), .Z(n8259) );
  NAND U10586 ( .A(n7703), .B(creg[30]), .Z(n8258) );
  NAND U10587 ( .A(n8260), .B(n8261), .Z(y[309]) );
  NAND U10588 ( .A(n7702), .B(m[309]), .Z(n8261) );
  NAND U10589 ( .A(n7703), .B(creg[309]), .Z(n8260) );
  NAND U10590 ( .A(n8262), .B(n8263), .Z(y[308]) );
  NAND U10591 ( .A(n7702), .B(m[308]), .Z(n8263) );
  NAND U10592 ( .A(n7703), .B(creg[308]), .Z(n8262) );
  NAND U10593 ( .A(n8264), .B(n8265), .Z(y[307]) );
  NAND U10594 ( .A(n7702), .B(m[307]), .Z(n8265) );
  NAND U10595 ( .A(n7703), .B(creg[307]), .Z(n8264) );
  NAND U10596 ( .A(n8266), .B(n8267), .Z(y[306]) );
  NAND U10597 ( .A(n7702), .B(m[306]), .Z(n8267) );
  NAND U10598 ( .A(n7703), .B(creg[306]), .Z(n8266) );
  NAND U10599 ( .A(n8268), .B(n8269), .Z(y[305]) );
  NAND U10600 ( .A(n7702), .B(m[305]), .Z(n8269) );
  NAND U10601 ( .A(n7703), .B(creg[305]), .Z(n8268) );
  NAND U10602 ( .A(n8270), .B(n8271), .Z(y[304]) );
  NAND U10603 ( .A(n7702), .B(m[304]), .Z(n8271) );
  NAND U10604 ( .A(n7703), .B(creg[304]), .Z(n8270) );
  NAND U10605 ( .A(n8272), .B(n8273), .Z(y[303]) );
  NAND U10606 ( .A(n7702), .B(m[303]), .Z(n8273) );
  NAND U10607 ( .A(n7703), .B(creg[303]), .Z(n8272) );
  NAND U10608 ( .A(n8274), .B(n8275), .Z(y[302]) );
  NAND U10609 ( .A(n7702), .B(m[302]), .Z(n8275) );
  NAND U10610 ( .A(n7703), .B(creg[302]), .Z(n8274) );
  NAND U10611 ( .A(n8276), .B(n8277), .Z(y[301]) );
  NAND U10612 ( .A(n7702), .B(m[301]), .Z(n8277) );
  NAND U10613 ( .A(n7703), .B(creg[301]), .Z(n8276) );
  NAND U10614 ( .A(n8278), .B(n8279), .Z(y[300]) );
  NAND U10615 ( .A(n7702), .B(m[300]), .Z(n8279) );
  NAND U10616 ( .A(n7703), .B(creg[300]), .Z(n8278) );
  NAND U10617 ( .A(n8280), .B(n8281), .Z(y[2]) );
  NAND U10618 ( .A(n7702), .B(m[2]), .Z(n8281) );
  NAND U10619 ( .A(n7703), .B(creg[2]), .Z(n8280) );
  NAND U10620 ( .A(n8282), .B(n8283), .Z(y[29]) );
  NAND U10621 ( .A(n7702), .B(m[29]), .Z(n8283) );
  NAND U10622 ( .A(n7703), .B(creg[29]), .Z(n8282) );
  NAND U10623 ( .A(n8284), .B(n8285), .Z(y[299]) );
  NAND U10624 ( .A(n7702), .B(m[299]), .Z(n8285) );
  NAND U10625 ( .A(n7703), .B(creg[299]), .Z(n8284) );
  NAND U10626 ( .A(n8286), .B(n8287), .Z(y[298]) );
  NAND U10627 ( .A(n7702), .B(m[298]), .Z(n8287) );
  NAND U10628 ( .A(n7703), .B(creg[298]), .Z(n8286) );
  NAND U10629 ( .A(n8288), .B(n8289), .Z(y[297]) );
  NAND U10630 ( .A(n7702), .B(m[297]), .Z(n8289) );
  NAND U10631 ( .A(n7703), .B(creg[297]), .Z(n8288) );
  NAND U10632 ( .A(n8290), .B(n8291), .Z(y[296]) );
  NAND U10633 ( .A(n7702), .B(m[296]), .Z(n8291) );
  NAND U10634 ( .A(n7703), .B(creg[296]), .Z(n8290) );
  NAND U10635 ( .A(n8292), .B(n8293), .Z(y[295]) );
  NAND U10636 ( .A(n7702), .B(m[295]), .Z(n8293) );
  NAND U10637 ( .A(n7703), .B(creg[295]), .Z(n8292) );
  NAND U10638 ( .A(n8294), .B(n8295), .Z(y[294]) );
  NAND U10639 ( .A(n7702), .B(m[294]), .Z(n8295) );
  NAND U10640 ( .A(n7703), .B(creg[294]), .Z(n8294) );
  NAND U10641 ( .A(n8296), .B(n8297), .Z(y[293]) );
  NAND U10642 ( .A(n7702), .B(m[293]), .Z(n8297) );
  NAND U10643 ( .A(n7703), .B(creg[293]), .Z(n8296) );
  NAND U10644 ( .A(n8298), .B(n8299), .Z(y[292]) );
  NAND U10645 ( .A(n7702), .B(m[292]), .Z(n8299) );
  NAND U10646 ( .A(n7703), .B(creg[292]), .Z(n8298) );
  NAND U10647 ( .A(n8300), .B(n8301), .Z(y[291]) );
  NAND U10648 ( .A(n7702), .B(m[291]), .Z(n8301) );
  NAND U10649 ( .A(n7703), .B(creg[291]), .Z(n8300) );
  NAND U10650 ( .A(n8302), .B(n8303), .Z(y[290]) );
  NAND U10651 ( .A(n7702), .B(m[290]), .Z(n8303) );
  NAND U10652 ( .A(n7703), .B(creg[290]), .Z(n8302) );
  NAND U10653 ( .A(n8304), .B(n8305), .Z(y[28]) );
  NAND U10654 ( .A(n7702), .B(m[28]), .Z(n8305) );
  NAND U10655 ( .A(n7703), .B(creg[28]), .Z(n8304) );
  NAND U10656 ( .A(n8306), .B(n8307), .Z(y[289]) );
  NAND U10657 ( .A(n7702), .B(m[289]), .Z(n8307) );
  NAND U10658 ( .A(n7703), .B(creg[289]), .Z(n8306) );
  NAND U10659 ( .A(n8308), .B(n8309), .Z(y[288]) );
  NAND U10660 ( .A(n7702), .B(m[288]), .Z(n8309) );
  NAND U10661 ( .A(n7703), .B(creg[288]), .Z(n8308) );
  NAND U10662 ( .A(n8310), .B(n8311), .Z(y[287]) );
  NAND U10663 ( .A(n7702), .B(m[287]), .Z(n8311) );
  NAND U10664 ( .A(n7703), .B(creg[287]), .Z(n8310) );
  NAND U10665 ( .A(n8312), .B(n8313), .Z(y[286]) );
  NAND U10666 ( .A(n7702), .B(m[286]), .Z(n8313) );
  NAND U10667 ( .A(n7703), .B(creg[286]), .Z(n8312) );
  NAND U10668 ( .A(n8314), .B(n8315), .Z(y[285]) );
  NAND U10669 ( .A(n7702), .B(m[285]), .Z(n8315) );
  NAND U10670 ( .A(n7703), .B(creg[285]), .Z(n8314) );
  NAND U10671 ( .A(n8316), .B(n8317), .Z(y[284]) );
  NAND U10672 ( .A(n7702), .B(m[284]), .Z(n8317) );
  NAND U10673 ( .A(n7703), .B(creg[284]), .Z(n8316) );
  NAND U10674 ( .A(n8318), .B(n8319), .Z(y[283]) );
  NAND U10675 ( .A(n7702), .B(m[283]), .Z(n8319) );
  NAND U10676 ( .A(n7703), .B(creg[283]), .Z(n8318) );
  NAND U10677 ( .A(n8320), .B(n8321), .Z(y[282]) );
  NAND U10678 ( .A(n7702), .B(m[282]), .Z(n8321) );
  NAND U10679 ( .A(n7703), .B(creg[282]), .Z(n8320) );
  NAND U10680 ( .A(n8322), .B(n8323), .Z(y[281]) );
  NAND U10681 ( .A(n7702), .B(m[281]), .Z(n8323) );
  NAND U10682 ( .A(n7703), .B(creg[281]), .Z(n8322) );
  NAND U10683 ( .A(n8324), .B(n8325), .Z(y[280]) );
  NAND U10684 ( .A(n7702), .B(m[280]), .Z(n8325) );
  NAND U10685 ( .A(n7703), .B(creg[280]), .Z(n8324) );
  NAND U10686 ( .A(n8326), .B(n8327), .Z(y[27]) );
  NAND U10687 ( .A(n7702), .B(m[27]), .Z(n8327) );
  NAND U10688 ( .A(n7703), .B(creg[27]), .Z(n8326) );
  NAND U10689 ( .A(n8328), .B(n8329), .Z(y[279]) );
  NAND U10690 ( .A(n7702), .B(m[279]), .Z(n8329) );
  NAND U10691 ( .A(n7703), .B(creg[279]), .Z(n8328) );
  NAND U10692 ( .A(n8330), .B(n8331), .Z(y[278]) );
  NAND U10693 ( .A(n7702), .B(m[278]), .Z(n8331) );
  NAND U10694 ( .A(n7703), .B(creg[278]), .Z(n8330) );
  NAND U10695 ( .A(n8332), .B(n8333), .Z(y[277]) );
  NAND U10696 ( .A(n7702), .B(m[277]), .Z(n8333) );
  NAND U10697 ( .A(n7703), .B(creg[277]), .Z(n8332) );
  NAND U10698 ( .A(n8334), .B(n8335), .Z(y[276]) );
  NAND U10699 ( .A(n7702), .B(m[276]), .Z(n8335) );
  NAND U10700 ( .A(n7703), .B(creg[276]), .Z(n8334) );
  NAND U10701 ( .A(n8336), .B(n8337), .Z(y[275]) );
  NAND U10702 ( .A(n7702), .B(m[275]), .Z(n8337) );
  NAND U10703 ( .A(n7703), .B(creg[275]), .Z(n8336) );
  NAND U10704 ( .A(n8338), .B(n8339), .Z(y[274]) );
  NAND U10705 ( .A(n7702), .B(m[274]), .Z(n8339) );
  NAND U10706 ( .A(n7703), .B(creg[274]), .Z(n8338) );
  NAND U10707 ( .A(n8340), .B(n8341), .Z(y[273]) );
  NAND U10708 ( .A(n7702), .B(m[273]), .Z(n8341) );
  NAND U10709 ( .A(n7703), .B(creg[273]), .Z(n8340) );
  NAND U10710 ( .A(n8342), .B(n8343), .Z(y[272]) );
  NAND U10711 ( .A(n7702), .B(m[272]), .Z(n8343) );
  NAND U10712 ( .A(n7703), .B(creg[272]), .Z(n8342) );
  NAND U10713 ( .A(n8344), .B(n8345), .Z(y[271]) );
  NAND U10714 ( .A(n7702), .B(m[271]), .Z(n8345) );
  NAND U10715 ( .A(n7703), .B(creg[271]), .Z(n8344) );
  NAND U10716 ( .A(n8346), .B(n8347), .Z(y[270]) );
  NAND U10717 ( .A(n7702), .B(m[270]), .Z(n8347) );
  NAND U10718 ( .A(n7703), .B(creg[270]), .Z(n8346) );
  NAND U10719 ( .A(n8348), .B(n8349), .Z(y[26]) );
  NAND U10720 ( .A(n7702), .B(m[26]), .Z(n8349) );
  NAND U10721 ( .A(n7703), .B(creg[26]), .Z(n8348) );
  NAND U10722 ( .A(n8350), .B(n8351), .Z(y[269]) );
  NAND U10723 ( .A(n7702), .B(m[269]), .Z(n8351) );
  NAND U10724 ( .A(n7703), .B(creg[269]), .Z(n8350) );
  NAND U10725 ( .A(n8352), .B(n8353), .Z(y[268]) );
  NAND U10726 ( .A(n7702), .B(m[268]), .Z(n8353) );
  NAND U10727 ( .A(n7703), .B(creg[268]), .Z(n8352) );
  NAND U10728 ( .A(n8354), .B(n8355), .Z(y[267]) );
  NAND U10729 ( .A(n7702), .B(m[267]), .Z(n8355) );
  NAND U10730 ( .A(n7703), .B(creg[267]), .Z(n8354) );
  NAND U10731 ( .A(n8356), .B(n8357), .Z(y[266]) );
  NAND U10732 ( .A(n7702), .B(m[266]), .Z(n8357) );
  NAND U10733 ( .A(n7703), .B(creg[266]), .Z(n8356) );
  NAND U10734 ( .A(n8358), .B(n8359), .Z(y[265]) );
  NAND U10735 ( .A(n7702), .B(m[265]), .Z(n8359) );
  NAND U10736 ( .A(n7703), .B(creg[265]), .Z(n8358) );
  NAND U10737 ( .A(n8360), .B(n8361), .Z(y[264]) );
  NAND U10738 ( .A(n7702), .B(m[264]), .Z(n8361) );
  NAND U10739 ( .A(n7703), .B(creg[264]), .Z(n8360) );
  NAND U10740 ( .A(n8362), .B(n8363), .Z(y[263]) );
  NAND U10741 ( .A(n7702), .B(m[263]), .Z(n8363) );
  NAND U10742 ( .A(n7703), .B(creg[263]), .Z(n8362) );
  NAND U10743 ( .A(n8364), .B(n8365), .Z(y[262]) );
  NAND U10744 ( .A(n7702), .B(m[262]), .Z(n8365) );
  NAND U10745 ( .A(n7703), .B(creg[262]), .Z(n8364) );
  NAND U10746 ( .A(n8366), .B(n8367), .Z(y[261]) );
  NAND U10747 ( .A(n7702), .B(m[261]), .Z(n8367) );
  NAND U10748 ( .A(n7703), .B(creg[261]), .Z(n8366) );
  NAND U10749 ( .A(n8368), .B(n8369), .Z(y[260]) );
  NAND U10750 ( .A(n7702), .B(m[260]), .Z(n8369) );
  NAND U10751 ( .A(n7703), .B(creg[260]), .Z(n8368) );
  NAND U10752 ( .A(n8370), .B(n8371), .Z(y[25]) );
  NAND U10753 ( .A(n7702), .B(m[25]), .Z(n8371) );
  NAND U10754 ( .A(n7703), .B(creg[25]), .Z(n8370) );
  NAND U10755 ( .A(n8372), .B(n8373), .Z(y[259]) );
  NAND U10756 ( .A(n7702), .B(m[259]), .Z(n8373) );
  NAND U10757 ( .A(n7703), .B(creg[259]), .Z(n8372) );
  NAND U10758 ( .A(n8374), .B(n8375), .Z(y[258]) );
  NAND U10759 ( .A(n7702), .B(m[258]), .Z(n8375) );
  NAND U10760 ( .A(n7703), .B(creg[258]), .Z(n8374) );
  NAND U10761 ( .A(n8376), .B(n8377), .Z(y[257]) );
  NAND U10762 ( .A(n7702), .B(m[257]), .Z(n8377) );
  NAND U10763 ( .A(n7703), .B(creg[257]), .Z(n8376) );
  NAND U10764 ( .A(n8378), .B(n8379), .Z(y[256]) );
  NAND U10765 ( .A(n7702), .B(m[256]), .Z(n8379) );
  NAND U10766 ( .A(n7703), .B(creg[256]), .Z(n8378) );
  NAND U10767 ( .A(n8380), .B(n8381), .Z(y[255]) );
  NAND U10768 ( .A(n7702), .B(m[255]), .Z(n8381) );
  NAND U10769 ( .A(n7703), .B(creg[255]), .Z(n8380) );
  NAND U10770 ( .A(n8382), .B(n8383), .Z(y[254]) );
  NAND U10771 ( .A(n7702), .B(m[254]), .Z(n8383) );
  NAND U10772 ( .A(n7703), .B(creg[254]), .Z(n8382) );
  NAND U10773 ( .A(n8384), .B(n8385), .Z(y[253]) );
  NAND U10774 ( .A(n7702), .B(m[253]), .Z(n8385) );
  NAND U10775 ( .A(n7703), .B(creg[253]), .Z(n8384) );
  NAND U10776 ( .A(n8386), .B(n8387), .Z(y[252]) );
  NAND U10777 ( .A(n7702), .B(m[252]), .Z(n8387) );
  NAND U10778 ( .A(n7703), .B(creg[252]), .Z(n8386) );
  NAND U10779 ( .A(n8388), .B(n8389), .Z(y[251]) );
  NAND U10780 ( .A(n7702), .B(m[251]), .Z(n8389) );
  NAND U10781 ( .A(n7703), .B(creg[251]), .Z(n8388) );
  NAND U10782 ( .A(n8390), .B(n8391), .Z(y[250]) );
  NAND U10783 ( .A(n7702), .B(m[250]), .Z(n8391) );
  NAND U10784 ( .A(n7703), .B(creg[250]), .Z(n8390) );
  NAND U10785 ( .A(n8392), .B(n8393), .Z(y[24]) );
  NAND U10786 ( .A(n7702), .B(m[24]), .Z(n8393) );
  NAND U10787 ( .A(n7703), .B(creg[24]), .Z(n8392) );
  NAND U10788 ( .A(n8394), .B(n8395), .Z(y[249]) );
  NAND U10789 ( .A(n7702), .B(m[249]), .Z(n8395) );
  NAND U10790 ( .A(n7703), .B(creg[249]), .Z(n8394) );
  NAND U10791 ( .A(n8396), .B(n8397), .Z(y[248]) );
  NAND U10792 ( .A(n7702), .B(m[248]), .Z(n8397) );
  NAND U10793 ( .A(n7703), .B(creg[248]), .Z(n8396) );
  NAND U10794 ( .A(n8398), .B(n8399), .Z(y[247]) );
  NAND U10795 ( .A(n7702), .B(m[247]), .Z(n8399) );
  NAND U10796 ( .A(n7703), .B(creg[247]), .Z(n8398) );
  NAND U10797 ( .A(n8400), .B(n8401), .Z(y[246]) );
  NAND U10798 ( .A(n7702), .B(m[246]), .Z(n8401) );
  NAND U10799 ( .A(n7703), .B(creg[246]), .Z(n8400) );
  NAND U10800 ( .A(n8402), .B(n8403), .Z(y[245]) );
  NAND U10801 ( .A(n7702), .B(m[245]), .Z(n8403) );
  NAND U10802 ( .A(n7703), .B(creg[245]), .Z(n8402) );
  NAND U10803 ( .A(n8404), .B(n8405), .Z(y[244]) );
  NAND U10804 ( .A(n7702), .B(m[244]), .Z(n8405) );
  NAND U10805 ( .A(n7703), .B(creg[244]), .Z(n8404) );
  NAND U10806 ( .A(n8406), .B(n8407), .Z(y[243]) );
  NAND U10807 ( .A(n7702), .B(m[243]), .Z(n8407) );
  NAND U10808 ( .A(n7703), .B(creg[243]), .Z(n8406) );
  NAND U10809 ( .A(n8408), .B(n8409), .Z(y[242]) );
  NAND U10810 ( .A(n7702), .B(m[242]), .Z(n8409) );
  NAND U10811 ( .A(n7703), .B(creg[242]), .Z(n8408) );
  NAND U10812 ( .A(n8410), .B(n8411), .Z(y[241]) );
  NAND U10813 ( .A(n7702), .B(m[241]), .Z(n8411) );
  NAND U10814 ( .A(n7703), .B(creg[241]), .Z(n8410) );
  NAND U10815 ( .A(n8412), .B(n8413), .Z(y[240]) );
  NAND U10816 ( .A(n7702), .B(m[240]), .Z(n8413) );
  NAND U10817 ( .A(n7703), .B(creg[240]), .Z(n8412) );
  NAND U10818 ( .A(n8414), .B(n8415), .Z(y[23]) );
  NAND U10819 ( .A(n7702), .B(m[23]), .Z(n8415) );
  NAND U10820 ( .A(n7703), .B(creg[23]), .Z(n8414) );
  NAND U10821 ( .A(n8416), .B(n8417), .Z(y[239]) );
  NAND U10822 ( .A(n7702), .B(m[239]), .Z(n8417) );
  NAND U10823 ( .A(n7703), .B(creg[239]), .Z(n8416) );
  NAND U10824 ( .A(n8418), .B(n8419), .Z(y[238]) );
  NAND U10825 ( .A(n7702), .B(m[238]), .Z(n8419) );
  NAND U10826 ( .A(n7703), .B(creg[238]), .Z(n8418) );
  NAND U10827 ( .A(n8420), .B(n8421), .Z(y[237]) );
  NAND U10828 ( .A(n7702), .B(m[237]), .Z(n8421) );
  NAND U10829 ( .A(n7703), .B(creg[237]), .Z(n8420) );
  NAND U10830 ( .A(n8422), .B(n8423), .Z(y[236]) );
  NAND U10831 ( .A(n7702), .B(m[236]), .Z(n8423) );
  NAND U10832 ( .A(n7703), .B(creg[236]), .Z(n8422) );
  NAND U10833 ( .A(n8424), .B(n8425), .Z(y[235]) );
  NAND U10834 ( .A(n7702), .B(m[235]), .Z(n8425) );
  NAND U10835 ( .A(n7703), .B(creg[235]), .Z(n8424) );
  NAND U10836 ( .A(n8426), .B(n8427), .Z(y[234]) );
  NAND U10837 ( .A(n7702), .B(m[234]), .Z(n8427) );
  NAND U10838 ( .A(n7703), .B(creg[234]), .Z(n8426) );
  NAND U10839 ( .A(n8428), .B(n8429), .Z(y[233]) );
  NAND U10840 ( .A(n7702), .B(m[233]), .Z(n8429) );
  NAND U10841 ( .A(n7703), .B(creg[233]), .Z(n8428) );
  NAND U10842 ( .A(n8430), .B(n8431), .Z(y[232]) );
  NAND U10843 ( .A(n7702), .B(m[232]), .Z(n8431) );
  NAND U10844 ( .A(n7703), .B(creg[232]), .Z(n8430) );
  NAND U10845 ( .A(n8432), .B(n8433), .Z(y[231]) );
  NAND U10846 ( .A(n7702), .B(m[231]), .Z(n8433) );
  NAND U10847 ( .A(n7703), .B(creg[231]), .Z(n8432) );
  NAND U10848 ( .A(n8434), .B(n8435), .Z(y[230]) );
  NAND U10849 ( .A(n7702), .B(m[230]), .Z(n8435) );
  NAND U10850 ( .A(n7703), .B(creg[230]), .Z(n8434) );
  NAND U10851 ( .A(n8436), .B(n8437), .Z(y[22]) );
  NAND U10852 ( .A(n7702), .B(m[22]), .Z(n8437) );
  NAND U10853 ( .A(n7703), .B(creg[22]), .Z(n8436) );
  NAND U10854 ( .A(n8438), .B(n8439), .Z(y[229]) );
  NAND U10855 ( .A(n7702), .B(m[229]), .Z(n8439) );
  NAND U10856 ( .A(n7703), .B(creg[229]), .Z(n8438) );
  NAND U10857 ( .A(n8440), .B(n8441), .Z(y[228]) );
  NAND U10858 ( .A(n7702), .B(m[228]), .Z(n8441) );
  NAND U10859 ( .A(n7703), .B(creg[228]), .Z(n8440) );
  NAND U10860 ( .A(n8442), .B(n8443), .Z(y[227]) );
  NAND U10861 ( .A(n7702), .B(m[227]), .Z(n8443) );
  NAND U10862 ( .A(n7703), .B(creg[227]), .Z(n8442) );
  NAND U10863 ( .A(n8444), .B(n8445), .Z(y[226]) );
  NAND U10864 ( .A(n7702), .B(m[226]), .Z(n8445) );
  NAND U10865 ( .A(n7703), .B(creg[226]), .Z(n8444) );
  NAND U10866 ( .A(n8446), .B(n8447), .Z(y[225]) );
  NAND U10867 ( .A(n7702), .B(m[225]), .Z(n8447) );
  NAND U10868 ( .A(n7703), .B(creg[225]), .Z(n8446) );
  NAND U10869 ( .A(n8448), .B(n8449), .Z(y[224]) );
  NAND U10870 ( .A(n7702), .B(m[224]), .Z(n8449) );
  NAND U10871 ( .A(n7703), .B(creg[224]), .Z(n8448) );
  NAND U10872 ( .A(n8450), .B(n8451), .Z(y[223]) );
  NAND U10873 ( .A(n7702), .B(m[223]), .Z(n8451) );
  NAND U10874 ( .A(n7703), .B(creg[223]), .Z(n8450) );
  NAND U10875 ( .A(n8452), .B(n8453), .Z(y[222]) );
  NAND U10876 ( .A(n7702), .B(m[222]), .Z(n8453) );
  NAND U10877 ( .A(n7703), .B(creg[222]), .Z(n8452) );
  NAND U10878 ( .A(n8454), .B(n8455), .Z(y[221]) );
  NAND U10879 ( .A(n7702), .B(m[221]), .Z(n8455) );
  NAND U10880 ( .A(n7703), .B(creg[221]), .Z(n8454) );
  NAND U10881 ( .A(n8456), .B(n8457), .Z(y[220]) );
  NAND U10882 ( .A(n7702), .B(m[220]), .Z(n8457) );
  NAND U10883 ( .A(n7703), .B(creg[220]), .Z(n8456) );
  NAND U10884 ( .A(n8458), .B(n8459), .Z(y[21]) );
  NAND U10885 ( .A(n7702), .B(m[21]), .Z(n8459) );
  NAND U10886 ( .A(n7703), .B(creg[21]), .Z(n8458) );
  NAND U10887 ( .A(n8460), .B(n8461), .Z(y[219]) );
  NAND U10888 ( .A(n7702), .B(m[219]), .Z(n8461) );
  NAND U10889 ( .A(n7703), .B(creg[219]), .Z(n8460) );
  NAND U10890 ( .A(n8462), .B(n8463), .Z(y[218]) );
  NAND U10891 ( .A(n7702), .B(m[218]), .Z(n8463) );
  NAND U10892 ( .A(n7703), .B(creg[218]), .Z(n8462) );
  NAND U10893 ( .A(n8464), .B(n8465), .Z(y[217]) );
  NAND U10894 ( .A(n7702), .B(m[217]), .Z(n8465) );
  NAND U10895 ( .A(n7703), .B(creg[217]), .Z(n8464) );
  NAND U10896 ( .A(n8466), .B(n8467), .Z(y[216]) );
  NAND U10897 ( .A(n7702), .B(m[216]), .Z(n8467) );
  NAND U10898 ( .A(n7703), .B(creg[216]), .Z(n8466) );
  NAND U10899 ( .A(n8468), .B(n8469), .Z(y[215]) );
  NAND U10900 ( .A(n7702), .B(m[215]), .Z(n8469) );
  NAND U10901 ( .A(n7703), .B(creg[215]), .Z(n8468) );
  NAND U10902 ( .A(n8470), .B(n8471), .Z(y[214]) );
  NAND U10903 ( .A(n7702), .B(m[214]), .Z(n8471) );
  NAND U10904 ( .A(n7703), .B(creg[214]), .Z(n8470) );
  NAND U10905 ( .A(n8472), .B(n8473), .Z(y[213]) );
  NAND U10906 ( .A(n7702), .B(m[213]), .Z(n8473) );
  NAND U10907 ( .A(n7703), .B(creg[213]), .Z(n8472) );
  NAND U10908 ( .A(n8474), .B(n8475), .Z(y[212]) );
  NAND U10909 ( .A(n7702), .B(m[212]), .Z(n8475) );
  NAND U10910 ( .A(n7703), .B(creg[212]), .Z(n8474) );
  NAND U10911 ( .A(n8476), .B(n8477), .Z(y[211]) );
  NAND U10912 ( .A(n7702), .B(m[211]), .Z(n8477) );
  NAND U10913 ( .A(n7703), .B(creg[211]), .Z(n8476) );
  NAND U10914 ( .A(n8478), .B(n8479), .Z(y[210]) );
  NAND U10915 ( .A(n7702), .B(m[210]), .Z(n8479) );
  NAND U10916 ( .A(n7703), .B(creg[210]), .Z(n8478) );
  NAND U10917 ( .A(n8480), .B(n8481), .Z(y[20]) );
  NAND U10918 ( .A(n7702), .B(m[20]), .Z(n8481) );
  NAND U10919 ( .A(n7703), .B(creg[20]), .Z(n8480) );
  NAND U10920 ( .A(n8482), .B(n8483), .Z(y[209]) );
  NAND U10921 ( .A(n7702), .B(m[209]), .Z(n8483) );
  NAND U10922 ( .A(n7703), .B(creg[209]), .Z(n8482) );
  NAND U10923 ( .A(n8484), .B(n8485), .Z(y[208]) );
  NAND U10924 ( .A(n7702), .B(m[208]), .Z(n8485) );
  NAND U10925 ( .A(n7703), .B(creg[208]), .Z(n8484) );
  NAND U10926 ( .A(n8486), .B(n8487), .Z(y[207]) );
  NAND U10927 ( .A(n7702), .B(m[207]), .Z(n8487) );
  NAND U10928 ( .A(n7703), .B(creg[207]), .Z(n8486) );
  NAND U10929 ( .A(n8488), .B(n8489), .Z(y[206]) );
  NAND U10930 ( .A(n7702), .B(m[206]), .Z(n8489) );
  NAND U10931 ( .A(n7703), .B(creg[206]), .Z(n8488) );
  NAND U10932 ( .A(n8490), .B(n8491), .Z(y[205]) );
  NAND U10933 ( .A(n7702), .B(m[205]), .Z(n8491) );
  NAND U10934 ( .A(n7703), .B(creg[205]), .Z(n8490) );
  NAND U10935 ( .A(n8492), .B(n8493), .Z(y[204]) );
  NAND U10936 ( .A(n7702), .B(m[204]), .Z(n8493) );
  NAND U10937 ( .A(n7703), .B(creg[204]), .Z(n8492) );
  NAND U10938 ( .A(n8494), .B(n8495), .Z(y[203]) );
  NAND U10939 ( .A(n7702), .B(m[203]), .Z(n8495) );
  NAND U10940 ( .A(n7703), .B(creg[203]), .Z(n8494) );
  NAND U10941 ( .A(n8496), .B(n8497), .Z(y[202]) );
  NAND U10942 ( .A(n7702), .B(m[202]), .Z(n8497) );
  NAND U10943 ( .A(n7703), .B(creg[202]), .Z(n8496) );
  NAND U10944 ( .A(n8498), .B(n8499), .Z(y[201]) );
  NAND U10945 ( .A(n7702), .B(m[201]), .Z(n8499) );
  NAND U10946 ( .A(n7703), .B(creg[201]), .Z(n8498) );
  NAND U10947 ( .A(n8500), .B(n8501), .Z(y[200]) );
  NAND U10948 ( .A(n7702), .B(m[200]), .Z(n8501) );
  NAND U10949 ( .A(n7703), .B(creg[200]), .Z(n8500) );
  NAND U10950 ( .A(n8502), .B(n8503), .Z(y[1]) );
  NAND U10951 ( .A(n7702), .B(m[1]), .Z(n8503) );
  NAND U10952 ( .A(n7703), .B(creg[1]), .Z(n8502) );
  NAND U10953 ( .A(n8504), .B(n8505), .Z(y[19]) );
  NAND U10954 ( .A(n7702), .B(m[19]), .Z(n8505) );
  NAND U10955 ( .A(n7703), .B(creg[19]), .Z(n8504) );
  NAND U10956 ( .A(n8506), .B(n8507), .Z(y[199]) );
  NAND U10957 ( .A(n7702), .B(m[199]), .Z(n8507) );
  NAND U10958 ( .A(n7703), .B(creg[199]), .Z(n8506) );
  NAND U10959 ( .A(n8508), .B(n8509), .Z(y[198]) );
  NAND U10960 ( .A(n7702), .B(m[198]), .Z(n8509) );
  NAND U10961 ( .A(n7703), .B(creg[198]), .Z(n8508) );
  NAND U10962 ( .A(n8510), .B(n8511), .Z(y[197]) );
  NAND U10963 ( .A(n7702), .B(m[197]), .Z(n8511) );
  NAND U10964 ( .A(n7703), .B(creg[197]), .Z(n8510) );
  NAND U10965 ( .A(n8512), .B(n8513), .Z(y[196]) );
  NAND U10966 ( .A(n7702), .B(m[196]), .Z(n8513) );
  NAND U10967 ( .A(n7703), .B(creg[196]), .Z(n8512) );
  NAND U10968 ( .A(n8514), .B(n8515), .Z(y[195]) );
  NAND U10969 ( .A(n7702), .B(m[195]), .Z(n8515) );
  NAND U10970 ( .A(n7703), .B(creg[195]), .Z(n8514) );
  NAND U10971 ( .A(n8516), .B(n8517), .Z(y[194]) );
  NAND U10972 ( .A(n7702), .B(m[194]), .Z(n8517) );
  NAND U10973 ( .A(n7703), .B(creg[194]), .Z(n8516) );
  NAND U10974 ( .A(n8518), .B(n8519), .Z(y[193]) );
  NAND U10975 ( .A(n7702), .B(m[193]), .Z(n8519) );
  NAND U10976 ( .A(n7703), .B(creg[193]), .Z(n8518) );
  NAND U10977 ( .A(n8520), .B(n8521), .Z(y[192]) );
  NAND U10978 ( .A(n7702), .B(m[192]), .Z(n8521) );
  NAND U10979 ( .A(n7703), .B(creg[192]), .Z(n8520) );
  NAND U10980 ( .A(n8522), .B(n8523), .Z(y[191]) );
  NAND U10981 ( .A(n7702), .B(m[191]), .Z(n8523) );
  NAND U10982 ( .A(n7703), .B(creg[191]), .Z(n8522) );
  NAND U10983 ( .A(n8524), .B(n8525), .Z(y[190]) );
  NAND U10984 ( .A(n7702), .B(m[190]), .Z(n8525) );
  NAND U10985 ( .A(n7703), .B(creg[190]), .Z(n8524) );
  NAND U10986 ( .A(n8526), .B(n8527), .Z(y[18]) );
  NAND U10987 ( .A(n7702), .B(m[18]), .Z(n8527) );
  NAND U10988 ( .A(n7703), .B(creg[18]), .Z(n8526) );
  NAND U10989 ( .A(n8528), .B(n8529), .Z(y[189]) );
  NAND U10990 ( .A(n7702), .B(m[189]), .Z(n8529) );
  NAND U10991 ( .A(n7703), .B(creg[189]), .Z(n8528) );
  NAND U10992 ( .A(n8530), .B(n8531), .Z(y[188]) );
  NAND U10993 ( .A(n7702), .B(m[188]), .Z(n8531) );
  NAND U10994 ( .A(n7703), .B(creg[188]), .Z(n8530) );
  NAND U10995 ( .A(n8532), .B(n8533), .Z(y[187]) );
  NAND U10996 ( .A(n7702), .B(m[187]), .Z(n8533) );
  NAND U10997 ( .A(n7703), .B(creg[187]), .Z(n8532) );
  NAND U10998 ( .A(n8534), .B(n8535), .Z(y[186]) );
  NAND U10999 ( .A(n7702), .B(m[186]), .Z(n8535) );
  NAND U11000 ( .A(n7703), .B(creg[186]), .Z(n8534) );
  NAND U11001 ( .A(n8536), .B(n8537), .Z(y[185]) );
  NAND U11002 ( .A(n7702), .B(m[185]), .Z(n8537) );
  NAND U11003 ( .A(n7703), .B(creg[185]), .Z(n8536) );
  NAND U11004 ( .A(n8538), .B(n8539), .Z(y[184]) );
  NAND U11005 ( .A(n7702), .B(m[184]), .Z(n8539) );
  NAND U11006 ( .A(n7703), .B(creg[184]), .Z(n8538) );
  NAND U11007 ( .A(n8540), .B(n8541), .Z(y[183]) );
  NAND U11008 ( .A(n7702), .B(m[183]), .Z(n8541) );
  NAND U11009 ( .A(n7703), .B(creg[183]), .Z(n8540) );
  NAND U11010 ( .A(n8542), .B(n8543), .Z(y[182]) );
  NAND U11011 ( .A(n7702), .B(m[182]), .Z(n8543) );
  NAND U11012 ( .A(n7703), .B(creg[182]), .Z(n8542) );
  NAND U11013 ( .A(n8544), .B(n8545), .Z(y[181]) );
  NAND U11014 ( .A(n7702), .B(m[181]), .Z(n8545) );
  NAND U11015 ( .A(n7703), .B(creg[181]), .Z(n8544) );
  NAND U11016 ( .A(n8546), .B(n8547), .Z(y[180]) );
  NAND U11017 ( .A(n7702), .B(m[180]), .Z(n8547) );
  NAND U11018 ( .A(n7703), .B(creg[180]), .Z(n8546) );
  NAND U11019 ( .A(n8548), .B(n8549), .Z(y[17]) );
  NAND U11020 ( .A(n7702), .B(m[17]), .Z(n8549) );
  NAND U11021 ( .A(n7703), .B(creg[17]), .Z(n8548) );
  NAND U11022 ( .A(n8550), .B(n8551), .Z(y[179]) );
  NAND U11023 ( .A(n7702), .B(m[179]), .Z(n8551) );
  NAND U11024 ( .A(n7703), .B(creg[179]), .Z(n8550) );
  NAND U11025 ( .A(n8552), .B(n8553), .Z(y[178]) );
  NAND U11026 ( .A(n7702), .B(m[178]), .Z(n8553) );
  NAND U11027 ( .A(n7703), .B(creg[178]), .Z(n8552) );
  NAND U11028 ( .A(n8554), .B(n8555), .Z(y[177]) );
  NAND U11029 ( .A(n7702), .B(m[177]), .Z(n8555) );
  NAND U11030 ( .A(n7703), .B(creg[177]), .Z(n8554) );
  NAND U11031 ( .A(n8556), .B(n8557), .Z(y[176]) );
  NAND U11032 ( .A(n7702), .B(m[176]), .Z(n8557) );
  NAND U11033 ( .A(n7703), .B(creg[176]), .Z(n8556) );
  NAND U11034 ( .A(n8558), .B(n8559), .Z(y[175]) );
  NAND U11035 ( .A(n7702), .B(m[175]), .Z(n8559) );
  NAND U11036 ( .A(n7703), .B(creg[175]), .Z(n8558) );
  NAND U11037 ( .A(n8560), .B(n8561), .Z(y[174]) );
  NAND U11038 ( .A(n7702), .B(m[174]), .Z(n8561) );
  NAND U11039 ( .A(n7703), .B(creg[174]), .Z(n8560) );
  NAND U11040 ( .A(n8562), .B(n8563), .Z(y[173]) );
  NAND U11041 ( .A(n7702), .B(m[173]), .Z(n8563) );
  NAND U11042 ( .A(n7703), .B(creg[173]), .Z(n8562) );
  NAND U11043 ( .A(n8564), .B(n8565), .Z(y[172]) );
  NAND U11044 ( .A(n7702), .B(m[172]), .Z(n8565) );
  NAND U11045 ( .A(n7703), .B(creg[172]), .Z(n8564) );
  NAND U11046 ( .A(n8566), .B(n8567), .Z(y[171]) );
  NAND U11047 ( .A(n7702), .B(m[171]), .Z(n8567) );
  NAND U11048 ( .A(n7703), .B(creg[171]), .Z(n8566) );
  NAND U11049 ( .A(n8568), .B(n8569), .Z(y[170]) );
  NAND U11050 ( .A(n7702), .B(m[170]), .Z(n8569) );
  NAND U11051 ( .A(n7703), .B(creg[170]), .Z(n8568) );
  NAND U11052 ( .A(n8570), .B(n8571), .Z(y[16]) );
  NAND U11053 ( .A(n7702), .B(m[16]), .Z(n8571) );
  NAND U11054 ( .A(n7703), .B(creg[16]), .Z(n8570) );
  NAND U11055 ( .A(n8572), .B(n8573), .Z(y[169]) );
  NAND U11056 ( .A(n7702), .B(m[169]), .Z(n8573) );
  NAND U11057 ( .A(n7703), .B(creg[169]), .Z(n8572) );
  NAND U11058 ( .A(n8574), .B(n8575), .Z(y[168]) );
  NAND U11059 ( .A(n7702), .B(m[168]), .Z(n8575) );
  NAND U11060 ( .A(n7703), .B(creg[168]), .Z(n8574) );
  NAND U11061 ( .A(n8576), .B(n8577), .Z(y[167]) );
  NAND U11062 ( .A(n7702), .B(m[167]), .Z(n8577) );
  NAND U11063 ( .A(n7703), .B(creg[167]), .Z(n8576) );
  NAND U11064 ( .A(n8578), .B(n8579), .Z(y[166]) );
  NAND U11065 ( .A(n7702), .B(m[166]), .Z(n8579) );
  NAND U11066 ( .A(n7703), .B(creg[166]), .Z(n8578) );
  NAND U11067 ( .A(n8580), .B(n8581), .Z(y[165]) );
  NAND U11068 ( .A(n7702), .B(m[165]), .Z(n8581) );
  NAND U11069 ( .A(n7703), .B(creg[165]), .Z(n8580) );
  NAND U11070 ( .A(n8582), .B(n8583), .Z(y[164]) );
  NAND U11071 ( .A(n7702), .B(m[164]), .Z(n8583) );
  NAND U11072 ( .A(n7703), .B(creg[164]), .Z(n8582) );
  NAND U11073 ( .A(n8584), .B(n8585), .Z(y[163]) );
  NAND U11074 ( .A(n7702), .B(m[163]), .Z(n8585) );
  NAND U11075 ( .A(n7703), .B(creg[163]), .Z(n8584) );
  NAND U11076 ( .A(n8586), .B(n8587), .Z(y[162]) );
  NAND U11077 ( .A(n7702), .B(m[162]), .Z(n8587) );
  NAND U11078 ( .A(n7703), .B(creg[162]), .Z(n8586) );
  NAND U11079 ( .A(n8588), .B(n8589), .Z(y[161]) );
  NAND U11080 ( .A(n7702), .B(m[161]), .Z(n8589) );
  NAND U11081 ( .A(n7703), .B(creg[161]), .Z(n8588) );
  NAND U11082 ( .A(n8590), .B(n8591), .Z(y[160]) );
  NAND U11083 ( .A(n7702), .B(m[160]), .Z(n8591) );
  NAND U11084 ( .A(n7703), .B(creg[160]), .Z(n8590) );
  NAND U11085 ( .A(n8592), .B(n8593), .Z(y[15]) );
  NAND U11086 ( .A(n7702), .B(m[15]), .Z(n8593) );
  NAND U11087 ( .A(n7703), .B(creg[15]), .Z(n8592) );
  NAND U11088 ( .A(n8594), .B(n8595), .Z(y[159]) );
  NAND U11089 ( .A(n7702), .B(m[159]), .Z(n8595) );
  NAND U11090 ( .A(n7703), .B(creg[159]), .Z(n8594) );
  NAND U11091 ( .A(n8596), .B(n8597), .Z(y[158]) );
  NAND U11092 ( .A(n7702), .B(m[158]), .Z(n8597) );
  NAND U11093 ( .A(n7703), .B(creg[158]), .Z(n8596) );
  NAND U11094 ( .A(n8598), .B(n8599), .Z(y[157]) );
  NAND U11095 ( .A(n7702), .B(m[157]), .Z(n8599) );
  NAND U11096 ( .A(n7703), .B(creg[157]), .Z(n8598) );
  NAND U11097 ( .A(n8600), .B(n8601), .Z(y[156]) );
  NAND U11098 ( .A(n7702), .B(m[156]), .Z(n8601) );
  NAND U11099 ( .A(n7703), .B(creg[156]), .Z(n8600) );
  NAND U11100 ( .A(n8602), .B(n8603), .Z(y[155]) );
  NAND U11101 ( .A(n7702), .B(m[155]), .Z(n8603) );
  NAND U11102 ( .A(n7703), .B(creg[155]), .Z(n8602) );
  NAND U11103 ( .A(n8604), .B(n8605), .Z(y[154]) );
  NAND U11104 ( .A(n7702), .B(m[154]), .Z(n8605) );
  NAND U11105 ( .A(n7703), .B(creg[154]), .Z(n8604) );
  NAND U11106 ( .A(n8606), .B(n8607), .Z(y[153]) );
  NAND U11107 ( .A(n7702), .B(m[153]), .Z(n8607) );
  NAND U11108 ( .A(n7703), .B(creg[153]), .Z(n8606) );
  NAND U11109 ( .A(n8608), .B(n8609), .Z(y[152]) );
  NAND U11110 ( .A(n7702), .B(m[152]), .Z(n8609) );
  NAND U11111 ( .A(n7703), .B(creg[152]), .Z(n8608) );
  NAND U11112 ( .A(n8610), .B(n8611), .Z(y[151]) );
  NAND U11113 ( .A(n7702), .B(m[151]), .Z(n8611) );
  NAND U11114 ( .A(n7703), .B(creg[151]), .Z(n8610) );
  NAND U11115 ( .A(n8612), .B(n8613), .Z(y[150]) );
  NAND U11116 ( .A(n7702), .B(m[150]), .Z(n8613) );
  NAND U11117 ( .A(n7703), .B(creg[150]), .Z(n8612) );
  NAND U11118 ( .A(n8614), .B(n8615), .Z(y[14]) );
  NAND U11119 ( .A(n7702), .B(m[14]), .Z(n8615) );
  NAND U11120 ( .A(n7703), .B(creg[14]), .Z(n8614) );
  NAND U11121 ( .A(n8616), .B(n8617), .Z(y[149]) );
  NAND U11122 ( .A(n7702), .B(m[149]), .Z(n8617) );
  NAND U11123 ( .A(n7703), .B(creg[149]), .Z(n8616) );
  NAND U11124 ( .A(n8618), .B(n8619), .Z(y[148]) );
  NAND U11125 ( .A(n7702), .B(m[148]), .Z(n8619) );
  NAND U11126 ( .A(n7703), .B(creg[148]), .Z(n8618) );
  NAND U11127 ( .A(n8620), .B(n8621), .Z(y[147]) );
  NAND U11128 ( .A(n7702), .B(m[147]), .Z(n8621) );
  NAND U11129 ( .A(n7703), .B(creg[147]), .Z(n8620) );
  NAND U11130 ( .A(n8622), .B(n8623), .Z(y[146]) );
  NAND U11131 ( .A(n7702), .B(m[146]), .Z(n8623) );
  NAND U11132 ( .A(n7703), .B(creg[146]), .Z(n8622) );
  NAND U11133 ( .A(n8624), .B(n8625), .Z(y[145]) );
  NAND U11134 ( .A(n7702), .B(m[145]), .Z(n8625) );
  NAND U11135 ( .A(n7703), .B(creg[145]), .Z(n8624) );
  NAND U11136 ( .A(n8626), .B(n8627), .Z(y[144]) );
  NAND U11137 ( .A(n7702), .B(m[144]), .Z(n8627) );
  NAND U11138 ( .A(n7703), .B(creg[144]), .Z(n8626) );
  NAND U11139 ( .A(n8628), .B(n8629), .Z(y[143]) );
  NAND U11140 ( .A(n7702), .B(m[143]), .Z(n8629) );
  NAND U11141 ( .A(n7703), .B(creg[143]), .Z(n8628) );
  NAND U11142 ( .A(n8630), .B(n8631), .Z(y[142]) );
  NAND U11143 ( .A(n7702), .B(m[142]), .Z(n8631) );
  NAND U11144 ( .A(n7703), .B(creg[142]), .Z(n8630) );
  NAND U11145 ( .A(n8632), .B(n8633), .Z(y[141]) );
  NAND U11146 ( .A(n7702), .B(m[141]), .Z(n8633) );
  NAND U11147 ( .A(n7703), .B(creg[141]), .Z(n8632) );
  NAND U11148 ( .A(n8634), .B(n8635), .Z(y[140]) );
  NAND U11149 ( .A(n7702), .B(m[140]), .Z(n8635) );
  NAND U11150 ( .A(n7703), .B(creg[140]), .Z(n8634) );
  NAND U11151 ( .A(n8636), .B(n8637), .Z(y[13]) );
  NAND U11152 ( .A(n7702), .B(m[13]), .Z(n8637) );
  NAND U11153 ( .A(n7703), .B(creg[13]), .Z(n8636) );
  NAND U11154 ( .A(n8638), .B(n8639), .Z(y[139]) );
  NAND U11155 ( .A(n7702), .B(m[139]), .Z(n8639) );
  NAND U11156 ( .A(n7703), .B(creg[139]), .Z(n8638) );
  NAND U11157 ( .A(n8640), .B(n8641), .Z(y[138]) );
  NAND U11158 ( .A(n7702), .B(m[138]), .Z(n8641) );
  NAND U11159 ( .A(n7703), .B(creg[138]), .Z(n8640) );
  NAND U11160 ( .A(n8642), .B(n8643), .Z(y[137]) );
  NAND U11161 ( .A(n7702), .B(m[137]), .Z(n8643) );
  NAND U11162 ( .A(n7703), .B(creg[137]), .Z(n8642) );
  NAND U11163 ( .A(n8644), .B(n8645), .Z(y[136]) );
  NAND U11164 ( .A(n7702), .B(m[136]), .Z(n8645) );
  NAND U11165 ( .A(n7703), .B(creg[136]), .Z(n8644) );
  NAND U11166 ( .A(n8646), .B(n8647), .Z(y[135]) );
  NAND U11167 ( .A(n7702), .B(m[135]), .Z(n8647) );
  NAND U11168 ( .A(n7703), .B(creg[135]), .Z(n8646) );
  NAND U11169 ( .A(n8648), .B(n8649), .Z(y[134]) );
  NAND U11170 ( .A(n7702), .B(m[134]), .Z(n8649) );
  NAND U11171 ( .A(n7703), .B(creg[134]), .Z(n8648) );
  NAND U11172 ( .A(n8650), .B(n8651), .Z(y[133]) );
  NAND U11173 ( .A(n7702), .B(m[133]), .Z(n8651) );
  NAND U11174 ( .A(n7703), .B(creg[133]), .Z(n8650) );
  NAND U11175 ( .A(n8652), .B(n8653), .Z(y[132]) );
  NAND U11176 ( .A(n7702), .B(m[132]), .Z(n8653) );
  NAND U11177 ( .A(n7703), .B(creg[132]), .Z(n8652) );
  NAND U11178 ( .A(n8654), .B(n8655), .Z(y[131]) );
  NAND U11179 ( .A(n7702), .B(m[131]), .Z(n8655) );
  NAND U11180 ( .A(n7703), .B(creg[131]), .Z(n8654) );
  NAND U11181 ( .A(n8656), .B(n8657), .Z(y[130]) );
  NAND U11182 ( .A(n7702), .B(m[130]), .Z(n8657) );
  NAND U11183 ( .A(n7703), .B(creg[130]), .Z(n8656) );
  NAND U11184 ( .A(n8658), .B(n8659), .Z(y[12]) );
  NAND U11185 ( .A(n7702), .B(m[12]), .Z(n8659) );
  NAND U11186 ( .A(n7703), .B(creg[12]), .Z(n8658) );
  NAND U11187 ( .A(n8660), .B(n8661), .Z(y[129]) );
  NAND U11188 ( .A(n7702), .B(m[129]), .Z(n8661) );
  NAND U11189 ( .A(n7703), .B(creg[129]), .Z(n8660) );
  NAND U11190 ( .A(n8662), .B(n8663), .Z(y[128]) );
  NAND U11191 ( .A(n7702), .B(m[128]), .Z(n8663) );
  NAND U11192 ( .A(n7703), .B(creg[128]), .Z(n8662) );
  NAND U11193 ( .A(n8664), .B(n8665), .Z(y[127]) );
  NAND U11194 ( .A(n7702), .B(m[127]), .Z(n8665) );
  NAND U11195 ( .A(n7703), .B(creg[127]), .Z(n8664) );
  NAND U11196 ( .A(n8666), .B(n8667), .Z(y[126]) );
  NAND U11197 ( .A(n7702), .B(m[126]), .Z(n8667) );
  NAND U11198 ( .A(n7703), .B(creg[126]), .Z(n8666) );
  NAND U11199 ( .A(n8668), .B(n8669), .Z(y[125]) );
  NAND U11200 ( .A(n7702), .B(m[125]), .Z(n8669) );
  NAND U11201 ( .A(n7703), .B(creg[125]), .Z(n8668) );
  NAND U11202 ( .A(n8670), .B(n8671), .Z(y[124]) );
  NAND U11203 ( .A(n7702), .B(m[124]), .Z(n8671) );
  NAND U11204 ( .A(n7703), .B(creg[124]), .Z(n8670) );
  NAND U11205 ( .A(n8672), .B(n8673), .Z(y[123]) );
  NAND U11206 ( .A(n7702), .B(m[123]), .Z(n8673) );
  NAND U11207 ( .A(n7703), .B(creg[123]), .Z(n8672) );
  NAND U11208 ( .A(n8674), .B(n8675), .Z(y[122]) );
  NAND U11209 ( .A(n7702), .B(m[122]), .Z(n8675) );
  NAND U11210 ( .A(n7703), .B(creg[122]), .Z(n8674) );
  NAND U11211 ( .A(n8676), .B(n8677), .Z(y[121]) );
  NAND U11212 ( .A(n7702), .B(m[121]), .Z(n8677) );
  NAND U11213 ( .A(n7703), .B(creg[121]), .Z(n8676) );
  NAND U11214 ( .A(n8678), .B(n8679), .Z(y[120]) );
  NAND U11215 ( .A(n7702), .B(m[120]), .Z(n8679) );
  NAND U11216 ( .A(n7703), .B(creg[120]), .Z(n8678) );
  NAND U11217 ( .A(n8680), .B(n8681), .Z(y[11]) );
  NAND U11218 ( .A(n7702), .B(m[11]), .Z(n8681) );
  NAND U11219 ( .A(n7703), .B(creg[11]), .Z(n8680) );
  NAND U11220 ( .A(n8682), .B(n8683), .Z(y[119]) );
  NAND U11221 ( .A(n7702), .B(m[119]), .Z(n8683) );
  NAND U11222 ( .A(n7703), .B(creg[119]), .Z(n8682) );
  NAND U11223 ( .A(n8684), .B(n8685), .Z(y[118]) );
  NAND U11224 ( .A(n7702), .B(m[118]), .Z(n8685) );
  NAND U11225 ( .A(n7703), .B(creg[118]), .Z(n8684) );
  NAND U11226 ( .A(n8686), .B(n8687), .Z(y[117]) );
  NAND U11227 ( .A(n7702), .B(m[117]), .Z(n8687) );
  NAND U11228 ( .A(n7703), .B(creg[117]), .Z(n8686) );
  NAND U11229 ( .A(n8688), .B(n8689), .Z(y[116]) );
  NAND U11230 ( .A(n7702), .B(m[116]), .Z(n8689) );
  NAND U11231 ( .A(n7703), .B(creg[116]), .Z(n8688) );
  NAND U11232 ( .A(n8690), .B(n8691), .Z(y[115]) );
  NAND U11233 ( .A(n7702), .B(m[115]), .Z(n8691) );
  NAND U11234 ( .A(n7703), .B(creg[115]), .Z(n8690) );
  NAND U11235 ( .A(n8692), .B(n8693), .Z(y[114]) );
  NAND U11236 ( .A(n7702), .B(m[114]), .Z(n8693) );
  NAND U11237 ( .A(n7703), .B(creg[114]), .Z(n8692) );
  NAND U11238 ( .A(n8694), .B(n8695), .Z(y[113]) );
  NAND U11239 ( .A(n7702), .B(m[113]), .Z(n8695) );
  NAND U11240 ( .A(n7703), .B(creg[113]), .Z(n8694) );
  NAND U11241 ( .A(n8696), .B(n8697), .Z(y[112]) );
  NAND U11242 ( .A(n7702), .B(m[112]), .Z(n8697) );
  NAND U11243 ( .A(n7703), .B(creg[112]), .Z(n8696) );
  NAND U11244 ( .A(n8698), .B(n8699), .Z(y[111]) );
  NAND U11245 ( .A(n7702), .B(m[111]), .Z(n8699) );
  NAND U11246 ( .A(n7703), .B(creg[111]), .Z(n8698) );
  NAND U11247 ( .A(n8700), .B(n8701), .Z(y[110]) );
  NAND U11248 ( .A(n7702), .B(m[110]), .Z(n8701) );
  NAND U11249 ( .A(n7703), .B(creg[110]), .Z(n8700) );
  NAND U11250 ( .A(n8702), .B(n8703), .Z(y[10]) );
  NAND U11251 ( .A(n7702), .B(m[10]), .Z(n8703) );
  NAND U11252 ( .A(n7703), .B(creg[10]), .Z(n8702) );
  NAND U11253 ( .A(n8704), .B(n8705), .Z(y[109]) );
  NAND U11254 ( .A(n7702), .B(m[109]), .Z(n8705) );
  NAND U11255 ( .A(n7703), .B(creg[109]), .Z(n8704) );
  NAND U11256 ( .A(n8706), .B(n8707), .Z(y[108]) );
  NAND U11257 ( .A(n7702), .B(m[108]), .Z(n8707) );
  NAND U11258 ( .A(n7703), .B(creg[108]), .Z(n8706) );
  NAND U11259 ( .A(n8708), .B(n8709), .Z(y[107]) );
  NAND U11260 ( .A(n7702), .B(m[107]), .Z(n8709) );
  NAND U11261 ( .A(n7703), .B(creg[107]), .Z(n8708) );
  NAND U11262 ( .A(n8710), .B(n8711), .Z(y[106]) );
  NAND U11263 ( .A(n7702), .B(m[106]), .Z(n8711) );
  NAND U11264 ( .A(n7703), .B(creg[106]), .Z(n8710) );
  NAND U11265 ( .A(n8712), .B(n8713), .Z(y[105]) );
  NAND U11266 ( .A(n7702), .B(m[105]), .Z(n8713) );
  NAND U11267 ( .A(n7703), .B(creg[105]), .Z(n8712) );
  NAND U11268 ( .A(n8714), .B(n8715), .Z(y[104]) );
  NAND U11269 ( .A(n7702), .B(m[104]), .Z(n8715) );
  NAND U11270 ( .A(n7703), .B(creg[104]), .Z(n8714) );
  NAND U11271 ( .A(n8716), .B(n8717), .Z(y[103]) );
  NAND U11272 ( .A(n7702), .B(m[103]), .Z(n8717) );
  NAND U11273 ( .A(n7703), .B(creg[103]), .Z(n8716) );
  NAND U11274 ( .A(n8718), .B(n8719), .Z(y[102]) );
  NAND U11275 ( .A(n7702), .B(m[102]), .Z(n8719) );
  NAND U11276 ( .A(n7703), .B(creg[102]), .Z(n8718) );
  NAND U11277 ( .A(n8720), .B(n8721), .Z(y[101]) );
  NAND U11278 ( .A(n7702), .B(m[101]), .Z(n8721) );
  NAND U11279 ( .A(n7703), .B(creg[101]), .Z(n8720) );
  NAND U11280 ( .A(n8722), .B(n8723), .Z(y[100]) );
  NAND U11281 ( .A(n7702), .B(m[100]), .Z(n8723) );
  NAND U11282 ( .A(n7703), .B(creg[100]), .Z(n8722) );
  NAND U11283 ( .A(n8724), .B(n8725), .Z(y[0]) );
  NAND U11284 ( .A(n7702), .B(m[0]), .Z(n8725) );
  NAND U11285 ( .A(n7703), .B(creg[0]), .Z(n8724) );
  NAND U11286 ( .A(n8726), .B(n8727), .Z(x[9]) );
  NAND U11287 ( .A(creg[9]), .B(init), .Z(n8726) );
  NAND U11288 ( .A(n8728), .B(n8729), .Z(x[99]) );
  NAND U11289 ( .A(creg[99]), .B(init), .Z(n8728) );
  NAND U11290 ( .A(n8730), .B(n8731), .Z(x[98]) );
  NAND U11291 ( .A(creg[98]), .B(init), .Z(n8730) );
  NAND U11292 ( .A(n8732), .B(n8733), .Z(x[97]) );
  NAND U11293 ( .A(creg[97]), .B(init), .Z(n8732) );
  NAND U11294 ( .A(n8734), .B(n8735), .Z(x[96]) );
  NAND U11295 ( .A(creg[96]), .B(init), .Z(n8734) );
  NAND U11296 ( .A(n8736), .B(n8737), .Z(x[95]) );
  NAND U11297 ( .A(creg[95]), .B(init), .Z(n8736) );
  NAND U11298 ( .A(n8738), .B(n8739), .Z(x[94]) );
  NAND U11299 ( .A(creg[94]), .B(init), .Z(n8738) );
  NAND U11300 ( .A(n8740), .B(n8741), .Z(x[93]) );
  NAND U11301 ( .A(creg[93]), .B(init), .Z(n8740) );
  NAND U11302 ( .A(n8742), .B(n8743), .Z(x[92]) );
  NAND U11303 ( .A(creg[92]), .B(init), .Z(n8742) );
  NAND U11304 ( .A(n8744), .B(n8745), .Z(x[91]) );
  NAND U11305 ( .A(creg[91]), .B(init), .Z(n8744) );
  NAND U11306 ( .A(n8746), .B(n8747), .Z(x[90]) );
  NAND U11307 ( .A(creg[90]), .B(init), .Z(n8746) );
  NAND U11308 ( .A(n8748), .B(n8749), .Z(x[8]) );
  NAND U11309 ( .A(creg[8]), .B(init), .Z(n8748) );
  NAND U11310 ( .A(n8750), .B(n8751), .Z(x[89]) );
  NAND U11311 ( .A(creg[89]), .B(init), .Z(n8750) );
  NAND U11312 ( .A(n8752), .B(n8753), .Z(x[88]) );
  NAND U11313 ( .A(creg[88]), .B(init), .Z(n8752) );
  NAND U11314 ( .A(n8754), .B(n8755), .Z(x[87]) );
  NAND U11315 ( .A(creg[87]), .B(init), .Z(n8754) );
  NAND U11316 ( .A(n8756), .B(n8757), .Z(x[86]) );
  NAND U11317 ( .A(creg[86]), .B(init), .Z(n8756) );
  NAND U11318 ( .A(n8758), .B(n8759), .Z(x[85]) );
  NAND U11319 ( .A(creg[85]), .B(init), .Z(n8758) );
  NAND U11320 ( .A(n8760), .B(n8761), .Z(x[84]) );
  NAND U11321 ( .A(creg[84]), .B(init), .Z(n8760) );
  NAND U11322 ( .A(n8762), .B(n8763), .Z(x[83]) );
  NAND U11323 ( .A(creg[83]), .B(init), .Z(n8762) );
  NAND U11324 ( .A(n8764), .B(n8765), .Z(x[82]) );
  NAND U11325 ( .A(creg[82]), .B(init), .Z(n8764) );
  NAND U11326 ( .A(n8766), .B(n8767), .Z(x[81]) );
  NAND U11327 ( .A(creg[81]), .B(init), .Z(n8766) );
  NAND U11328 ( .A(n8768), .B(n8769), .Z(x[80]) );
  NAND U11329 ( .A(creg[80]), .B(init), .Z(n8768) );
  NAND U11330 ( .A(n8770), .B(n8771), .Z(x[7]) );
  NAND U11331 ( .A(creg[7]), .B(init), .Z(n8770) );
  NAND U11332 ( .A(n8772), .B(n8773), .Z(x[79]) );
  NAND U11333 ( .A(creg[79]), .B(init), .Z(n8772) );
  NAND U11334 ( .A(n8774), .B(n8775), .Z(x[78]) );
  NAND U11335 ( .A(creg[78]), .B(init), .Z(n8774) );
  NAND U11336 ( .A(n8776), .B(n8777), .Z(x[77]) );
  NAND U11337 ( .A(creg[77]), .B(init), .Z(n8776) );
  NAND U11338 ( .A(n8778), .B(n8779), .Z(x[76]) );
  NAND U11339 ( .A(creg[76]), .B(init), .Z(n8778) );
  NAND U11340 ( .A(n8780), .B(n8781), .Z(x[75]) );
  NAND U11341 ( .A(creg[75]), .B(init), .Z(n8780) );
  NAND U11342 ( .A(n8782), .B(n8783), .Z(x[74]) );
  NAND U11343 ( .A(creg[74]), .B(init), .Z(n8782) );
  NAND U11344 ( .A(n8784), .B(n8785), .Z(x[73]) );
  NAND U11345 ( .A(creg[73]), .B(init), .Z(n8784) );
  NAND U11346 ( .A(n8786), .B(n8787), .Z(x[72]) );
  NAND U11347 ( .A(creg[72]), .B(init), .Z(n8786) );
  NAND U11348 ( .A(n8788), .B(n8789), .Z(x[71]) );
  NAND U11349 ( .A(creg[71]), .B(init), .Z(n8788) );
  NAND U11350 ( .A(n8790), .B(n8791), .Z(x[70]) );
  NAND U11351 ( .A(creg[70]), .B(init), .Z(n8790) );
  NAND U11352 ( .A(n8792), .B(n8793), .Z(x[6]) );
  NAND U11353 ( .A(creg[6]), .B(init), .Z(n8792) );
  NAND U11354 ( .A(n8794), .B(n8795), .Z(x[69]) );
  NAND U11355 ( .A(creg[69]), .B(init), .Z(n8794) );
  NAND U11356 ( .A(n8796), .B(n8797), .Z(x[68]) );
  NAND U11357 ( .A(creg[68]), .B(init), .Z(n8796) );
  NAND U11358 ( .A(n8798), .B(n8799), .Z(x[67]) );
  NAND U11359 ( .A(creg[67]), .B(init), .Z(n8798) );
  NAND U11360 ( .A(n8800), .B(n8801), .Z(x[66]) );
  NAND U11361 ( .A(creg[66]), .B(init), .Z(n8800) );
  NAND U11362 ( .A(n8802), .B(n8803), .Z(x[65]) );
  NAND U11363 ( .A(creg[65]), .B(init), .Z(n8802) );
  NAND U11364 ( .A(n8804), .B(n8805), .Z(x[64]) );
  NAND U11365 ( .A(creg[64]), .B(init), .Z(n8804) );
  NAND U11366 ( .A(n8806), .B(n8807), .Z(x[63]) );
  NAND U11367 ( .A(creg[63]), .B(init), .Z(n8806) );
  NAND U11368 ( .A(n8808), .B(n8809), .Z(x[62]) );
  NAND U11369 ( .A(creg[62]), .B(init), .Z(n8808) );
  NAND U11370 ( .A(n8810), .B(n8811), .Z(x[61]) );
  NAND U11371 ( .A(creg[61]), .B(init), .Z(n8810) );
  NAND U11372 ( .A(n8812), .B(n8813), .Z(x[60]) );
  NAND U11373 ( .A(creg[60]), .B(init), .Z(n8812) );
  NAND U11374 ( .A(n8814), .B(n8815), .Z(x[5]) );
  NAND U11375 ( .A(creg[5]), .B(init), .Z(n8814) );
  NAND U11376 ( .A(n8816), .B(n8817), .Z(x[59]) );
  NAND U11377 ( .A(creg[59]), .B(init), .Z(n8816) );
  NAND U11378 ( .A(n8818), .B(n8819), .Z(x[58]) );
  NAND U11379 ( .A(creg[58]), .B(init), .Z(n8818) );
  NAND U11380 ( .A(n8820), .B(n8821), .Z(x[57]) );
  NAND U11381 ( .A(creg[57]), .B(init), .Z(n8820) );
  NAND U11382 ( .A(n8822), .B(n8823), .Z(x[56]) );
  NAND U11383 ( .A(creg[56]), .B(init), .Z(n8822) );
  NAND U11384 ( .A(n8824), .B(n8825), .Z(x[55]) );
  NAND U11385 ( .A(creg[55]), .B(init), .Z(n8824) );
  NAND U11386 ( .A(n8826), .B(n8827), .Z(x[54]) );
  NAND U11387 ( .A(creg[54]), .B(init), .Z(n8826) );
  NAND U11388 ( .A(n8828), .B(n8829), .Z(x[53]) );
  NAND U11389 ( .A(creg[53]), .B(init), .Z(n8828) );
  NAND U11390 ( .A(n8830), .B(n8831), .Z(x[52]) );
  NAND U11391 ( .A(creg[52]), .B(init), .Z(n8830) );
  NAND U11392 ( .A(n8832), .B(n8833), .Z(x[51]) );
  NAND U11393 ( .A(creg[51]), .B(init), .Z(n8832) );
  NAND U11394 ( .A(n8834), .B(n8835), .Z(x[511]) );
  NAND U11395 ( .A(creg[511]), .B(init), .Z(n8834) );
  NAND U11396 ( .A(n8836), .B(n8837), .Z(x[510]) );
  NAND U11397 ( .A(creg[510]), .B(init), .Z(n8836) );
  NAND U11398 ( .A(n8838), .B(n8839), .Z(x[50]) );
  NAND U11399 ( .A(creg[50]), .B(init), .Z(n8838) );
  NAND U11400 ( .A(n8840), .B(n8841), .Z(x[509]) );
  NAND U11401 ( .A(creg[509]), .B(init), .Z(n8840) );
  NAND U11402 ( .A(n8842), .B(n8843), .Z(x[508]) );
  NAND U11403 ( .A(creg[508]), .B(init), .Z(n8842) );
  NAND U11404 ( .A(n8844), .B(n8845), .Z(x[507]) );
  NAND U11405 ( .A(creg[507]), .B(init), .Z(n8844) );
  NAND U11406 ( .A(n8846), .B(n8847), .Z(x[506]) );
  NAND U11407 ( .A(creg[506]), .B(init), .Z(n8846) );
  NAND U11408 ( .A(n8848), .B(n8849), .Z(x[505]) );
  NAND U11409 ( .A(creg[505]), .B(init), .Z(n8848) );
  NAND U11410 ( .A(n8850), .B(n8851), .Z(x[504]) );
  NAND U11411 ( .A(creg[504]), .B(init), .Z(n8850) );
  NAND U11412 ( .A(n8852), .B(n8853), .Z(x[503]) );
  NAND U11413 ( .A(creg[503]), .B(init), .Z(n8852) );
  NAND U11414 ( .A(n8854), .B(n8855), .Z(x[502]) );
  NAND U11415 ( .A(creg[502]), .B(init), .Z(n8854) );
  NAND U11416 ( .A(n8856), .B(n8857), .Z(x[501]) );
  NAND U11417 ( .A(creg[501]), .B(init), .Z(n8856) );
  NAND U11418 ( .A(n8858), .B(n8859), .Z(x[500]) );
  NAND U11419 ( .A(creg[500]), .B(init), .Z(n8858) );
  NAND U11420 ( .A(n8860), .B(n8861), .Z(x[4]) );
  NAND U11421 ( .A(creg[4]), .B(init), .Z(n8860) );
  NAND U11422 ( .A(n8862), .B(n8863), .Z(x[49]) );
  NAND U11423 ( .A(creg[49]), .B(init), .Z(n8862) );
  NAND U11424 ( .A(n8864), .B(n8865), .Z(x[499]) );
  NAND U11425 ( .A(creg[499]), .B(init), .Z(n8864) );
  NAND U11426 ( .A(n8866), .B(n8867), .Z(x[498]) );
  NAND U11427 ( .A(creg[498]), .B(init), .Z(n8866) );
  NAND U11428 ( .A(n8868), .B(n8869), .Z(x[497]) );
  NAND U11429 ( .A(creg[497]), .B(init), .Z(n8868) );
  NAND U11430 ( .A(n8870), .B(n8871), .Z(x[496]) );
  NAND U11431 ( .A(creg[496]), .B(init), .Z(n8870) );
  NAND U11432 ( .A(n8872), .B(n8873), .Z(x[495]) );
  NAND U11433 ( .A(creg[495]), .B(init), .Z(n8872) );
  NAND U11434 ( .A(n8874), .B(n8875), .Z(x[494]) );
  NAND U11435 ( .A(creg[494]), .B(init), .Z(n8874) );
  NAND U11436 ( .A(n8876), .B(n8877), .Z(x[493]) );
  NAND U11437 ( .A(creg[493]), .B(init), .Z(n8876) );
  NAND U11438 ( .A(n8878), .B(n8879), .Z(x[492]) );
  NAND U11439 ( .A(creg[492]), .B(init), .Z(n8878) );
  NAND U11440 ( .A(n8880), .B(n8881), .Z(x[491]) );
  NAND U11441 ( .A(creg[491]), .B(init), .Z(n8880) );
  NAND U11442 ( .A(n8882), .B(n8883), .Z(x[490]) );
  NAND U11443 ( .A(creg[490]), .B(init), .Z(n8882) );
  NAND U11444 ( .A(n8884), .B(n8885), .Z(x[48]) );
  NAND U11445 ( .A(creg[48]), .B(init), .Z(n8884) );
  NAND U11446 ( .A(n8886), .B(n8887), .Z(x[489]) );
  NAND U11447 ( .A(creg[489]), .B(init), .Z(n8886) );
  NAND U11448 ( .A(n8888), .B(n8889), .Z(x[488]) );
  NAND U11449 ( .A(creg[488]), .B(init), .Z(n8888) );
  NAND U11450 ( .A(n8890), .B(n8891), .Z(x[487]) );
  NAND U11451 ( .A(creg[487]), .B(init), .Z(n8890) );
  NAND U11452 ( .A(n8892), .B(n8893), .Z(x[486]) );
  NAND U11453 ( .A(creg[486]), .B(init), .Z(n8892) );
  NAND U11454 ( .A(n8894), .B(n8895), .Z(x[485]) );
  NAND U11455 ( .A(creg[485]), .B(init), .Z(n8894) );
  NAND U11456 ( .A(n8896), .B(n8897), .Z(x[484]) );
  NAND U11457 ( .A(creg[484]), .B(init), .Z(n8896) );
  NAND U11458 ( .A(n8898), .B(n8899), .Z(x[483]) );
  NAND U11459 ( .A(creg[483]), .B(init), .Z(n8898) );
  NAND U11460 ( .A(n8900), .B(n8901), .Z(x[482]) );
  NAND U11461 ( .A(creg[482]), .B(init), .Z(n8900) );
  NAND U11462 ( .A(n8902), .B(n8903), .Z(x[481]) );
  NAND U11463 ( .A(creg[481]), .B(init), .Z(n8902) );
  NAND U11464 ( .A(n8904), .B(n8905), .Z(x[480]) );
  NAND U11465 ( .A(creg[480]), .B(init), .Z(n8904) );
  NAND U11466 ( .A(n8906), .B(n8907), .Z(x[47]) );
  NAND U11467 ( .A(creg[47]), .B(init), .Z(n8906) );
  NAND U11468 ( .A(n8908), .B(n8909), .Z(x[479]) );
  NAND U11469 ( .A(creg[479]), .B(init), .Z(n8908) );
  NAND U11470 ( .A(n8910), .B(n8911), .Z(x[478]) );
  NAND U11471 ( .A(creg[478]), .B(init), .Z(n8910) );
  NAND U11472 ( .A(n8912), .B(n8913), .Z(x[477]) );
  NAND U11473 ( .A(creg[477]), .B(init), .Z(n8912) );
  NAND U11474 ( .A(n8914), .B(n8915), .Z(x[476]) );
  NAND U11475 ( .A(creg[476]), .B(init), .Z(n8914) );
  NAND U11476 ( .A(n8916), .B(n8917), .Z(x[475]) );
  NAND U11477 ( .A(creg[475]), .B(init), .Z(n8916) );
  NAND U11478 ( .A(n8918), .B(n8919), .Z(x[474]) );
  NAND U11479 ( .A(creg[474]), .B(init), .Z(n8918) );
  NAND U11480 ( .A(n8920), .B(n8921), .Z(x[473]) );
  NAND U11481 ( .A(creg[473]), .B(init), .Z(n8920) );
  NAND U11482 ( .A(n8922), .B(n8923), .Z(x[472]) );
  NAND U11483 ( .A(creg[472]), .B(init), .Z(n8922) );
  NAND U11484 ( .A(n8924), .B(n8925), .Z(x[471]) );
  NAND U11485 ( .A(creg[471]), .B(init), .Z(n8924) );
  NAND U11486 ( .A(n8926), .B(n8927), .Z(x[470]) );
  NAND U11487 ( .A(creg[470]), .B(init), .Z(n8926) );
  NAND U11488 ( .A(n8928), .B(n8929), .Z(x[46]) );
  NAND U11489 ( .A(creg[46]), .B(init), .Z(n8928) );
  NAND U11490 ( .A(n8930), .B(n8931), .Z(x[469]) );
  NAND U11491 ( .A(creg[469]), .B(init), .Z(n8930) );
  NAND U11492 ( .A(n8932), .B(n8933), .Z(x[468]) );
  NAND U11493 ( .A(creg[468]), .B(init), .Z(n8932) );
  NAND U11494 ( .A(n8934), .B(n8935), .Z(x[467]) );
  NAND U11495 ( .A(creg[467]), .B(init), .Z(n8934) );
  NAND U11496 ( .A(n8936), .B(n8937), .Z(x[466]) );
  NAND U11497 ( .A(creg[466]), .B(init), .Z(n8936) );
  NAND U11498 ( .A(n8938), .B(n8939), .Z(x[465]) );
  NAND U11499 ( .A(creg[465]), .B(init), .Z(n8938) );
  NAND U11500 ( .A(n8940), .B(n8941), .Z(x[464]) );
  NAND U11501 ( .A(creg[464]), .B(init), .Z(n8940) );
  NAND U11502 ( .A(n8942), .B(n8943), .Z(x[463]) );
  NAND U11503 ( .A(creg[463]), .B(init), .Z(n8942) );
  NAND U11504 ( .A(n8944), .B(n8945), .Z(x[462]) );
  NAND U11505 ( .A(creg[462]), .B(init), .Z(n8944) );
  NAND U11506 ( .A(n8946), .B(n8947), .Z(x[461]) );
  NAND U11507 ( .A(creg[461]), .B(init), .Z(n8946) );
  NAND U11508 ( .A(n8948), .B(n8949), .Z(x[460]) );
  NAND U11509 ( .A(creg[460]), .B(init), .Z(n8948) );
  NAND U11510 ( .A(n8950), .B(n8951), .Z(x[45]) );
  NAND U11511 ( .A(creg[45]), .B(init), .Z(n8950) );
  NAND U11512 ( .A(n8952), .B(n8953), .Z(x[459]) );
  NAND U11513 ( .A(creg[459]), .B(init), .Z(n8952) );
  NAND U11514 ( .A(n8954), .B(n8955), .Z(x[458]) );
  NAND U11515 ( .A(creg[458]), .B(init), .Z(n8954) );
  NAND U11516 ( .A(n8956), .B(n8957), .Z(x[457]) );
  NAND U11517 ( .A(creg[457]), .B(init), .Z(n8956) );
  NAND U11518 ( .A(n8958), .B(n8959), .Z(x[456]) );
  NAND U11519 ( .A(creg[456]), .B(init), .Z(n8958) );
  NAND U11520 ( .A(n8960), .B(n8961), .Z(x[455]) );
  NAND U11521 ( .A(creg[455]), .B(init), .Z(n8960) );
  NAND U11522 ( .A(n8962), .B(n8963), .Z(x[454]) );
  NAND U11523 ( .A(creg[454]), .B(init), .Z(n8962) );
  NAND U11524 ( .A(n8964), .B(n8965), .Z(x[453]) );
  NAND U11525 ( .A(creg[453]), .B(init), .Z(n8964) );
  NAND U11526 ( .A(n8966), .B(n8967), .Z(x[452]) );
  NAND U11527 ( .A(creg[452]), .B(init), .Z(n8966) );
  NAND U11528 ( .A(n8968), .B(n8969), .Z(x[451]) );
  NAND U11529 ( .A(creg[451]), .B(init), .Z(n8968) );
  NAND U11530 ( .A(n8970), .B(n8971), .Z(x[450]) );
  NAND U11531 ( .A(creg[450]), .B(init), .Z(n8970) );
  NAND U11532 ( .A(n8972), .B(n8973), .Z(x[44]) );
  NAND U11533 ( .A(creg[44]), .B(init), .Z(n8972) );
  NAND U11534 ( .A(n8974), .B(n8975), .Z(x[449]) );
  NAND U11535 ( .A(creg[449]), .B(init), .Z(n8974) );
  NAND U11536 ( .A(n8976), .B(n8977), .Z(x[448]) );
  NAND U11537 ( .A(creg[448]), .B(init), .Z(n8976) );
  NAND U11538 ( .A(n8978), .B(n8979), .Z(x[447]) );
  NAND U11539 ( .A(creg[447]), .B(init), .Z(n8978) );
  NAND U11540 ( .A(n8980), .B(n8981), .Z(x[446]) );
  NAND U11541 ( .A(creg[446]), .B(init), .Z(n8980) );
  NAND U11542 ( .A(n8982), .B(n8983), .Z(x[445]) );
  NAND U11543 ( .A(creg[445]), .B(init), .Z(n8982) );
  NAND U11544 ( .A(n8984), .B(n8985), .Z(x[444]) );
  NAND U11545 ( .A(creg[444]), .B(init), .Z(n8984) );
  NAND U11546 ( .A(n8986), .B(n8987), .Z(x[443]) );
  NAND U11547 ( .A(creg[443]), .B(init), .Z(n8986) );
  NAND U11548 ( .A(n8988), .B(n8989), .Z(x[442]) );
  NAND U11549 ( .A(creg[442]), .B(init), .Z(n8988) );
  NAND U11550 ( .A(n8990), .B(n8991), .Z(x[441]) );
  NAND U11551 ( .A(creg[441]), .B(init), .Z(n8990) );
  NAND U11552 ( .A(n8992), .B(n8993), .Z(x[440]) );
  NAND U11553 ( .A(creg[440]), .B(init), .Z(n8992) );
  NAND U11554 ( .A(n8994), .B(n8995), .Z(x[43]) );
  NAND U11555 ( .A(creg[43]), .B(init), .Z(n8994) );
  NAND U11556 ( .A(n8996), .B(n8997), .Z(x[439]) );
  NAND U11557 ( .A(creg[439]), .B(init), .Z(n8996) );
  NAND U11558 ( .A(n8998), .B(n8999), .Z(x[438]) );
  NAND U11559 ( .A(creg[438]), .B(init), .Z(n8998) );
  NAND U11560 ( .A(n9000), .B(n9001), .Z(x[437]) );
  NAND U11561 ( .A(creg[437]), .B(init), .Z(n9000) );
  NAND U11562 ( .A(n9002), .B(n9003), .Z(x[436]) );
  NAND U11563 ( .A(creg[436]), .B(init), .Z(n9002) );
  NAND U11564 ( .A(n9004), .B(n9005), .Z(x[435]) );
  NAND U11565 ( .A(creg[435]), .B(init), .Z(n9004) );
  NAND U11566 ( .A(n9006), .B(n9007), .Z(x[434]) );
  NAND U11567 ( .A(creg[434]), .B(init), .Z(n9006) );
  NAND U11568 ( .A(n9008), .B(n9009), .Z(x[433]) );
  NAND U11569 ( .A(creg[433]), .B(init), .Z(n9008) );
  NAND U11570 ( .A(n9010), .B(n9011), .Z(x[432]) );
  NAND U11571 ( .A(creg[432]), .B(init), .Z(n9010) );
  NAND U11572 ( .A(n9012), .B(n9013), .Z(x[431]) );
  NAND U11573 ( .A(creg[431]), .B(init), .Z(n9012) );
  NAND U11574 ( .A(n9014), .B(n9015), .Z(x[430]) );
  NAND U11575 ( .A(creg[430]), .B(init), .Z(n9014) );
  NAND U11576 ( .A(n9016), .B(n9017), .Z(x[42]) );
  NAND U11577 ( .A(creg[42]), .B(init), .Z(n9016) );
  NAND U11578 ( .A(n9018), .B(n9019), .Z(x[429]) );
  NAND U11579 ( .A(creg[429]), .B(init), .Z(n9018) );
  NAND U11580 ( .A(n9020), .B(n9021), .Z(x[428]) );
  NAND U11581 ( .A(creg[428]), .B(init), .Z(n9020) );
  NAND U11582 ( .A(n9022), .B(n9023), .Z(x[427]) );
  NAND U11583 ( .A(creg[427]), .B(init), .Z(n9022) );
  NAND U11584 ( .A(n9024), .B(n9025), .Z(x[426]) );
  NAND U11585 ( .A(creg[426]), .B(init), .Z(n9024) );
  NAND U11586 ( .A(n9026), .B(n9027), .Z(x[425]) );
  NAND U11587 ( .A(creg[425]), .B(init), .Z(n9026) );
  NAND U11588 ( .A(n9028), .B(n9029), .Z(x[424]) );
  NAND U11589 ( .A(creg[424]), .B(init), .Z(n9028) );
  NAND U11590 ( .A(n9030), .B(n9031), .Z(x[423]) );
  NAND U11591 ( .A(creg[423]), .B(init), .Z(n9030) );
  NAND U11592 ( .A(n9032), .B(n9033), .Z(x[422]) );
  NAND U11593 ( .A(creg[422]), .B(init), .Z(n9032) );
  NAND U11594 ( .A(n9034), .B(n9035), .Z(x[421]) );
  NAND U11595 ( .A(creg[421]), .B(init), .Z(n9034) );
  NAND U11596 ( .A(n9036), .B(n9037), .Z(x[420]) );
  NAND U11597 ( .A(creg[420]), .B(init), .Z(n9036) );
  NAND U11598 ( .A(n9038), .B(n9039), .Z(x[41]) );
  NAND U11599 ( .A(creg[41]), .B(init), .Z(n9038) );
  NAND U11600 ( .A(n9040), .B(n9041), .Z(x[419]) );
  NAND U11601 ( .A(creg[419]), .B(init), .Z(n9040) );
  NAND U11602 ( .A(n9042), .B(n9043), .Z(x[418]) );
  NAND U11603 ( .A(creg[418]), .B(init), .Z(n9042) );
  NAND U11604 ( .A(n9044), .B(n9045), .Z(x[417]) );
  NAND U11605 ( .A(creg[417]), .B(init), .Z(n9044) );
  NAND U11606 ( .A(n9046), .B(n9047), .Z(x[416]) );
  NAND U11607 ( .A(creg[416]), .B(init), .Z(n9046) );
  NAND U11608 ( .A(n9048), .B(n9049), .Z(x[415]) );
  NAND U11609 ( .A(creg[415]), .B(init), .Z(n9048) );
  NAND U11610 ( .A(n9050), .B(n9051), .Z(x[414]) );
  NAND U11611 ( .A(creg[414]), .B(init), .Z(n9050) );
  NAND U11612 ( .A(n9052), .B(n9053), .Z(x[413]) );
  NAND U11613 ( .A(creg[413]), .B(init), .Z(n9052) );
  NAND U11614 ( .A(n9054), .B(n9055), .Z(x[412]) );
  NAND U11615 ( .A(creg[412]), .B(init), .Z(n9054) );
  NAND U11616 ( .A(n9056), .B(n9057), .Z(x[411]) );
  NAND U11617 ( .A(creg[411]), .B(init), .Z(n9056) );
  NAND U11618 ( .A(n9058), .B(n9059), .Z(x[410]) );
  NAND U11619 ( .A(creg[410]), .B(init), .Z(n9058) );
  NAND U11620 ( .A(n9060), .B(n9061), .Z(x[40]) );
  NAND U11621 ( .A(creg[40]), .B(init), .Z(n9060) );
  NAND U11622 ( .A(n9062), .B(n9063), .Z(x[409]) );
  NAND U11623 ( .A(creg[409]), .B(init), .Z(n9062) );
  NAND U11624 ( .A(n9064), .B(n9065), .Z(x[408]) );
  NAND U11625 ( .A(creg[408]), .B(init), .Z(n9064) );
  NAND U11626 ( .A(n9066), .B(n9067), .Z(x[407]) );
  NAND U11627 ( .A(creg[407]), .B(init), .Z(n9066) );
  NAND U11628 ( .A(n9068), .B(n9069), .Z(x[406]) );
  NAND U11629 ( .A(creg[406]), .B(init), .Z(n9068) );
  NAND U11630 ( .A(n9070), .B(n9071), .Z(x[405]) );
  NAND U11631 ( .A(creg[405]), .B(init), .Z(n9070) );
  NAND U11632 ( .A(n9072), .B(n9073), .Z(x[404]) );
  NAND U11633 ( .A(creg[404]), .B(init), .Z(n9072) );
  NAND U11634 ( .A(n9074), .B(n9075), .Z(x[403]) );
  NAND U11635 ( .A(creg[403]), .B(init), .Z(n9074) );
  NAND U11636 ( .A(n9076), .B(n9077), .Z(x[402]) );
  NAND U11637 ( .A(creg[402]), .B(init), .Z(n9076) );
  NAND U11638 ( .A(n9078), .B(n9079), .Z(x[401]) );
  NAND U11639 ( .A(creg[401]), .B(init), .Z(n9078) );
  NAND U11640 ( .A(n9080), .B(n9081), .Z(x[400]) );
  NAND U11641 ( .A(creg[400]), .B(init), .Z(n9080) );
  NAND U11642 ( .A(n9082), .B(n9083), .Z(x[3]) );
  NAND U11643 ( .A(creg[3]), .B(init), .Z(n9082) );
  NAND U11644 ( .A(n9084), .B(n9085), .Z(x[39]) );
  NAND U11645 ( .A(creg[39]), .B(init), .Z(n9084) );
  NAND U11646 ( .A(n9086), .B(n9087), .Z(x[399]) );
  NAND U11647 ( .A(creg[399]), .B(init), .Z(n9086) );
  NAND U11648 ( .A(n9088), .B(n9089), .Z(x[398]) );
  NAND U11649 ( .A(creg[398]), .B(init), .Z(n9088) );
  NAND U11650 ( .A(n9090), .B(n9091), .Z(x[397]) );
  NAND U11651 ( .A(creg[397]), .B(init), .Z(n9090) );
  NAND U11652 ( .A(n9092), .B(n9093), .Z(x[396]) );
  NAND U11653 ( .A(creg[396]), .B(init), .Z(n9092) );
  NAND U11654 ( .A(n9094), .B(n9095), .Z(x[395]) );
  NAND U11655 ( .A(creg[395]), .B(init), .Z(n9094) );
  NAND U11656 ( .A(n9096), .B(n9097), .Z(x[394]) );
  NAND U11657 ( .A(creg[394]), .B(init), .Z(n9096) );
  NAND U11658 ( .A(n9098), .B(n9099), .Z(x[393]) );
  NAND U11659 ( .A(creg[393]), .B(init), .Z(n9098) );
  NAND U11660 ( .A(n9100), .B(n9101), .Z(x[392]) );
  NAND U11661 ( .A(creg[392]), .B(init), .Z(n9100) );
  NAND U11662 ( .A(n9102), .B(n9103), .Z(x[391]) );
  NAND U11663 ( .A(creg[391]), .B(init), .Z(n9102) );
  NAND U11664 ( .A(n9104), .B(n9105), .Z(x[390]) );
  NAND U11665 ( .A(creg[390]), .B(init), .Z(n9104) );
  NAND U11666 ( .A(n9106), .B(n9107), .Z(x[38]) );
  NAND U11667 ( .A(creg[38]), .B(init), .Z(n9106) );
  NAND U11668 ( .A(n9108), .B(n9109), .Z(x[389]) );
  NAND U11669 ( .A(creg[389]), .B(init), .Z(n9108) );
  NAND U11670 ( .A(n9110), .B(n9111), .Z(x[388]) );
  NAND U11671 ( .A(creg[388]), .B(init), .Z(n9110) );
  NAND U11672 ( .A(n9112), .B(n9113), .Z(x[387]) );
  NAND U11673 ( .A(creg[387]), .B(init), .Z(n9112) );
  NAND U11674 ( .A(n9114), .B(n9115), .Z(x[386]) );
  NAND U11675 ( .A(creg[386]), .B(init), .Z(n9114) );
  NAND U11676 ( .A(n9116), .B(n9117), .Z(x[385]) );
  NAND U11677 ( .A(creg[385]), .B(init), .Z(n9116) );
  NAND U11678 ( .A(n9118), .B(n9119), .Z(x[384]) );
  NAND U11679 ( .A(creg[384]), .B(init), .Z(n9118) );
  NAND U11680 ( .A(n9120), .B(n9121), .Z(x[383]) );
  NAND U11681 ( .A(creg[383]), .B(init), .Z(n9120) );
  NAND U11682 ( .A(n9122), .B(n9123), .Z(x[382]) );
  NAND U11683 ( .A(creg[382]), .B(init), .Z(n9122) );
  NAND U11684 ( .A(n9124), .B(n9125), .Z(x[381]) );
  NAND U11685 ( .A(creg[381]), .B(init), .Z(n9124) );
  NAND U11686 ( .A(n9126), .B(n9127), .Z(x[380]) );
  NAND U11687 ( .A(creg[380]), .B(init), .Z(n9126) );
  NAND U11688 ( .A(n9128), .B(n9129), .Z(x[37]) );
  NAND U11689 ( .A(creg[37]), .B(init), .Z(n9128) );
  NAND U11690 ( .A(n9130), .B(n9131), .Z(x[379]) );
  NAND U11691 ( .A(creg[379]), .B(init), .Z(n9130) );
  NAND U11692 ( .A(n9132), .B(n9133), .Z(x[378]) );
  NAND U11693 ( .A(creg[378]), .B(init), .Z(n9132) );
  NAND U11694 ( .A(n9134), .B(n9135), .Z(x[377]) );
  NAND U11695 ( .A(creg[377]), .B(init), .Z(n9134) );
  NAND U11696 ( .A(n9136), .B(n9137), .Z(x[376]) );
  NAND U11697 ( .A(creg[376]), .B(init), .Z(n9136) );
  NAND U11698 ( .A(n9138), .B(n9139), .Z(x[375]) );
  NAND U11699 ( .A(creg[375]), .B(init), .Z(n9138) );
  NAND U11700 ( .A(n9140), .B(n9141), .Z(x[374]) );
  NAND U11701 ( .A(creg[374]), .B(init), .Z(n9140) );
  NAND U11702 ( .A(n9142), .B(n9143), .Z(x[373]) );
  NAND U11703 ( .A(creg[373]), .B(init), .Z(n9142) );
  NAND U11704 ( .A(n9144), .B(n9145), .Z(x[372]) );
  NAND U11705 ( .A(creg[372]), .B(init), .Z(n9144) );
  NAND U11706 ( .A(n9146), .B(n9147), .Z(x[371]) );
  NAND U11707 ( .A(creg[371]), .B(init), .Z(n9146) );
  NAND U11708 ( .A(n9148), .B(n9149), .Z(x[370]) );
  NAND U11709 ( .A(creg[370]), .B(init), .Z(n9148) );
  NAND U11710 ( .A(n9150), .B(n9151), .Z(x[36]) );
  NAND U11711 ( .A(creg[36]), .B(init), .Z(n9150) );
  NAND U11712 ( .A(n9152), .B(n9153), .Z(x[369]) );
  NAND U11713 ( .A(creg[369]), .B(init), .Z(n9152) );
  NAND U11714 ( .A(n9154), .B(n9155), .Z(x[368]) );
  NAND U11715 ( .A(creg[368]), .B(init), .Z(n9154) );
  NAND U11716 ( .A(n9156), .B(n9157), .Z(x[367]) );
  NAND U11717 ( .A(creg[367]), .B(init), .Z(n9156) );
  NAND U11718 ( .A(n9158), .B(n9159), .Z(x[366]) );
  NAND U11719 ( .A(creg[366]), .B(init), .Z(n9158) );
  NAND U11720 ( .A(n9160), .B(n9161), .Z(x[365]) );
  NAND U11721 ( .A(creg[365]), .B(init), .Z(n9160) );
  NAND U11722 ( .A(n9162), .B(n9163), .Z(x[364]) );
  NAND U11723 ( .A(creg[364]), .B(init), .Z(n9162) );
  NAND U11724 ( .A(n9164), .B(n9165), .Z(x[363]) );
  NAND U11725 ( .A(creg[363]), .B(init), .Z(n9164) );
  NAND U11726 ( .A(n9166), .B(n9167), .Z(x[362]) );
  NAND U11727 ( .A(creg[362]), .B(init), .Z(n9166) );
  NAND U11728 ( .A(n9168), .B(n9169), .Z(x[361]) );
  NAND U11729 ( .A(creg[361]), .B(init), .Z(n9168) );
  NAND U11730 ( .A(n9170), .B(n9171), .Z(x[360]) );
  NAND U11731 ( .A(creg[360]), .B(init), .Z(n9170) );
  NAND U11732 ( .A(n9172), .B(n9173), .Z(x[35]) );
  NAND U11733 ( .A(creg[35]), .B(init), .Z(n9172) );
  NAND U11734 ( .A(n9174), .B(n9175), .Z(x[359]) );
  NAND U11735 ( .A(creg[359]), .B(init), .Z(n9174) );
  NAND U11736 ( .A(n9176), .B(n9177), .Z(x[358]) );
  NAND U11737 ( .A(creg[358]), .B(init), .Z(n9176) );
  NAND U11738 ( .A(n9178), .B(n9179), .Z(x[357]) );
  NAND U11739 ( .A(creg[357]), .B(init), .Z(n9178) );
  NAND U11740 ( .A(n9180), .B(n9181), .Z(x[356]) );
  NAND U11741 ( .A(creg[356]), .B(init), .Z(n9180) );
  NAND U11742 ( .A(n9182), .B(n9183), .Z(x[355]) );
  NAND U11743 ( .A(creg[355]), .B(init), .Z(n9182) );
  NAND U11744 ( .A(n9184), .B(n9185), .Z(x[354]) );
  NAND U11745 ( .A(creg[354]), .B(init), .Z(n9184) );
  NAND U11746 ( .A(n9186), .B(n9187), .Z(x[353]) );
  NAND U11747 ( .A(creg[353]), .B(init), .Z(n9186) );
  NAND U11748 ( .A(n9188), .B(n9189), .Z(x[352]) );
  NAND U11749 ( .A(creg[352]), .B(init), .Z(n9188) );
  NAND U11750 ( .A(n9190), .B(n9191), .Z(x[351]) );
  NAND U11751 ( .A(creg[351]), .B(init), .Z(n9190) );
  NAND U11752 ( .A(n9192), .B(n9193), .Z(x[350]) );
  NAND U11753 ( .A(creg[350]), .B(init), .Z(n9192) );
  NAND U11754 ( .A(n9194), .B(n9195), .Z(x[34]) );
  NAND U11755 ( .A(creg[34]), .B(init), .Z(n9194) );
  NAND U11756 ( .A(n9196), .B(n9197), .Z(x[349]) );
  NAND U11757 ( .A(creg[349]), .B(init), .Z(n9196) );
  NAND U11758 ( .A(n9198), .B(n9199), .Z(x[348]) );
  NAND U11759 ( .A(creg[348]), .B(init), .Z(n9198) );
  NAND U11760 ( .A(n9200), .B(n9201), .Z(x[347]) );
  NAND U11761 ( .A(creg[347]), .B(init), .Z(n9200) );
  NAND U11762 ( .A(n9202), .B(n9203), .Z(x[346]) );
  NAND U11763 ( .A(creg[346]), .B(init), .Z(n9202) );
  NAND U11764 ( .A(n9204), .B(n9205), .Z(x[345]) );
  NAND U11765 ( .A(creg[345]), .B(init), .Z(n9204) );
  NAND U11766 ( .A(n9206), .B(n9207), .Z(x[344]) );
  NAND U11767 ( .A(creg[344]), .B(init), .Z(n9206) );
  NAND U11768 ( .A(n9208), .B(n9209), .Z(x[343]) );
  NAND U11769 ( .A(creg[343]), .B(init), .Z(n9208) );
  NAND U11770 ( .A(n9210), .B(n9211), .Z(x[342]) );
  NAND U11771 ( .A(creg[342]), .B(init), .Z(n9210) );
  NAND U11772 ( .A(n9212), .B(n9213), .Z(x[341]) );
  NAND U11773 ( .A(creg[341]), .B(init), .Z(n9212) );
  NAND U11774 ( .A(n9214), .B(n9215), .Z(x[340]) );
  NAND U11775 ( .A(creg[340]), .B(init), .Z(n9214) );
  NAND U11776 ( .A(n9216), .B(n9217), .Z(x[33]) );
  NAND U11777 ( .A(creg[33]), .B(init), .Z(n9216) );
  NAND U11778 ( .A(n9218), .B(n9219), .Z(x[339]) );
  NAND U11779 ( .A(creg[339]), .B(init), .Z(n9218) );
  NAND U11780 ( .A(n9220), .B(n9221), .Z(x[338]) );
  NAND U11781 ( .A(creg[338]), .B(init), .Z(n9220) );
  NAND U11782 ( .A(n9222), .B(n9223), .Z(x[337]) );
  NAND U11783 ( .A(creg[337]), .B(init), .Z(n9222) );
  NAND U11784 ( .A(n9224), .B(n9225), .Z(x[336]) );
  NAND U11785 ( .A(creg[336]), .B(init), .Z(n9224) );
  NAND U11786 ( .A(n9226), .B(n9227), .Z(x[335]) );
  NAND U11787 ( .A(creg[335]), .B(init), .Z(n9226) );
  NAND U11788 ( .A(n9228), .B(n9229), .Z(x[334]) );
  NAND U11789 ( .A(creg[334]), .B(init), .Z(n9228) );
  NAND U11790 ( .A(n9230), .B(n9231), .Z(x[333]) );
  NAND U11791 ( .A(creg[333]), .B(init), .Z(n9230) );
  NAND U11792 ( .A(n9232), .B(n9233), .Z(x[332]) );
  NAND U11793 ( .A(creg[332]), .B(init), .Z(n9232) );
  NAND U11794 ( .A(n9234), .B(n9235), .Z(x[331]) );
  NAND U11795 ( .A(creg[331]), .B(init), .Z(n9234) );
  NAND U11796 ( .A(n9236), .B(n9237), .Z(x[330]) );
  NAND U11797 ( .A(creg[330]), .B(init), .Z(n9236) );
  NAND U11798 ( .A(n9238), .B(n9239), .Z(x[32]) );
  NAND U11799 ( .A(creg[32]), .B(init), .Z(n9238) );
  NAND U11800 ( .A(n9240), .B(n9241), .Z(x[329]) );
  NAND U11801 ( .A(creg[329]), .B(init), .Z(n9240) );
  NAND U11802 ( .A(n9242), .B(n9243), .Z(x[328]) );
  NAND U11803 ( .A(creg[328]), .B(init), .Z(n9242) );
  NAND U11804 ( .A(n9244), .B(n9245), .Z(x[327]) );
  NAND U11805 ( .A(creg[327]), .B(init), .Z(n9244) );
  NAND U11806 ( .A(n9246), .B(n9247), .Z(x[326]) );
  NAND U11807 ( .A(creg[326]), .B(init), .Z(n9246) );
  NAND U11808 ( .A(n9248), .B(n9249), .Z(x[325]) );
  NAND U11809 ( .A(creg[325]), .B(init), .Z(n9248) );
  NAND U11810 ( .A(n9250), .B(n9251), .Z(x[324]) );
  NAND U11811 ( .A(creg[324]), .B(init), .Z(n9250) );
  NAND U11812 ( .A(n9252), .B(n9253), .Z(x[323]) );
  NAND U11813 ( .A(creg[323]), .B(init), .Z(n9252) );
  NAND U11814 ( .A(n9254), .B(n9255), .Z(x[322]) );
  NAND U11815 ( .A(creg[322]), .B(init), .Z(n9254) );
  NAND U11816 ( .A(n9256), .B(n9257), .Z(x[321]) );
  NAND U11817 ( .A(creg[321]), .B(init), .Z(n9256) );
  NAND U11818 ( .A(n9258), .B(n9259), .Z(x[320]) );
  NAND U11819 ( .A(creg[320]), .B(init), .Z(n9258) );
  NAND U11820 ( .A(n9260), .B(n9261), .Z(x[31]) );
  NAND U11821 ( .A(creg[31]), .B(init), .Z(n9260) );
  NAND U11822 ( .A(n9262), .B(n9263), .Z(x[319]) );
  NAND U11823 ( .A(creg[319]), .B(init), .Z(n9262) );
  NAND U11824 ( .A(n9264), .B(n9265), .Z(x[318]) );
  NAND U11825 ( .A(creg[318]), .B(init), .Z(n9264) );
  NAND U11826 ( .A(n9266), .B(n9267), .Z(x[317]) );
  NAND U11827 ( .A(creg[317]), .B(init), .Z(n9266) );
  NAND U11828 ( .A(n9268), .B(n9269), .Z(x[316]) );
  NAND U11829 ( .A(creg[316]), .B(init), .Z(n9268) );
  NAND U11830 ( .A(n9270), .B(n9271), .Z(x[315]) );
  NAND U11831 ( .A(creg[315]), .B(init), .Z(n9270) );
  NAND U11832 ( .A(n9272), .B(n9273), .Z(x[314]) );
  NAND U11833 ( .A(creg[314]), .B(init), .Z(n9272) );
  NAND U11834 ( .A(n9274), .B(n9275), .Z(x[313]) );
  NAND U11835 ( .A(creg[313]), .B(init), .Z(n9274) );
  NAND U11836 ( .A(n9276), .B(n9277), .Z(x[312]) );
  NAND U11837 ( .A(creg[312]), .B(init), .Z(n9276) );
  NAND U11838 ( .A(n9278), .B(n9279), .Z(x[311]) );
  NAND U11839 ( .A(creg[311]), .B(init), .Z(n9278) );
  NAND U11840 ( .A(n9280), .B(n9281), .Z(x[310]) );
  NAND U11841 ( .A(creg[310]), .B(init), .Z(n9280) );
  NAND U11842 ( .A(n9282), .B(n9283), .Z(x[30]) );
  NAND U11843 ( .A(creg[30]), .B(init), .Z(n9282) );
  NAND U11844 ( .A(n9284), .B(n9285), .Z(x[309]) );
  NAND U11845 ( .A(creg[309]), .B(init), .Z(n9284) );
  NAND U11846 ( .A(n9286), .B(n9287), .Z(x[308]) );
  NAND U11847 ( .A(creg[308]), .B(init), .Z(n9286) );
  NAND U11848 ( .A(n9288), .B(n9289), .Z(x[307]) );
  NAND U11849 ( .A(creg[307]), .B(init), .Z(n9288) );
  NAND U11850 ( .A(n9290), .B(n9291), .Z(x[306]) );
  NAND U11851 ( .A(creg[306]), .B(init), .Z(n9290) );
  NAND U11852 ( .A(n9292), .B(n9293), .Z(x[305]) );
  NAND U11853 ( .A(creg[305]), .B(init), .Z(n9292) );
  NAND U11854 ( .A(n9294), .B(n9295), .Z(x[304]) );
  NAND U11855 ( .A(creg[304]), .B(init), .Z(n9294) );
  NAND U11856 ( .A(n9296), .B(n9297), .Z(x[303]) );
  NAND U11857 ( .A(creg[303]), .B(init), .Z(n9296) );
  NAND U11858 ( .A(n9298), .B(n9299), .Z(x[302]) );
  NAND U11859 ( .A(creg[302]), .B(init), .Z(n9298) );
  NAND U11860 ( .A(n9300), .B(n9301), .Z(x[301]) );
  NAND U11861 ( .A(creg[301]), .B(init), .Z(n9300) );
  NAND U11862 ( .A(n9302), .B(n9303), .Z(x[300]) );
  NAND U11863 ( .A(creg[300]), .B(init), .Z(n9302) );
  NAND U11864 ( .A(n9304), .B(n9305), .Z(x[2]) );
  NAND U11865 ( .A(creg[2]), .B(init), .Z(n9304) );
  NAND U11866 ( .A(n9306), .B(n9307), .Z(x[29]) );
  NAND U11867 ( .A(creg[29]), .B(init), .Z(n9306) );
  NAND U11868 ( .A(n9308), .B(n9309), .Z(x[299]) );
  NAND U11869 ( .A(creg[299]), .B(init), .Z(n9308) );
  NAND U11870 ( .A(n9310), .B(n9311), .Z(x[298]) );
  NAND U11871 ( .A(creg[298]), .B(init), .Z(n9310) );
  NAND U11872 ( .A(n9312), .B(n9313), .Z(x[297]) );
  NAND U11873 ( .A(creg[297]), .B(init), .Z(n9312) );
  NAND U11874 ( .A(n9314), .B(n9315), .Z(x[296]) );
  NAND U11875 ( .A(creg[296]), .B(init), .Z(n9314) );
  NAND U11876 ( .A(n9316), .B(n9317), .Z(x[295]) );
  NAND U11877 ( .A(creg[295]), .B(init), .Z(n9316) );
  NAND U11878 ( .A(n9318), .B(n9319), .Z(x[294]) );
  NAND U11879 ( .A(creg[294]), .B(init), .Z(n9318) );
  NAND U11880 ( .A(n9320), .B(n9321), .Z(x[293]) );
  NAND U11881 ( .A(creg[293]), .B(init), .Z(n9320) );
  NAND U11882 ( .A(n9322), .B(n9323), .Z(x[292]) );
  NAND U11883 ( .A(creg[292]), .B(init), .Z(n9322) );
  NAND U11884 ( .A(n9324), .B(n9325), .Z(x[291]) );
  NAND U11885 ( .A(creg[291]), .B(init), .Z(n9324) );
  NAND U11886 ( .A(n9326), .B(n9327), .Z(x[290]) );
  NAND U11887 ( .A(creg[290]), .B(init), .Z(n9326) );
  NAND U11888 ( .A(n9328), .B(n9329), .Z(x[28]) );
  NAND U11889 ( .A(creg[28]), .B(init), .Z(n9328) );
  NAND U11890 ( .A(n9330), .B(n9331), .Z(x[289]) );
  NAND U11891 ( .A(creg[289]), .B(init), .Z(n9330) );
  NAND U11892 ( .A(n9332), .B(n9333), .Z(x[288]) );
  NAND U11893 ( .A(creg[288]), .B(init), .Z(n9332) );
  NAND U11894 ( .A(n9334), .B(n9335), .Z(x[287]) );
  NAND U11895 ( .A(creg[287]), .B(init), .Z(n9334) );
  NAND U11896 ( .A(n9336), .B(n9337), .Z(x[286]) );
  NAND U11897 ( .A(creg[286]), .B(init), .Z(n9336) );
  NAND U11898 ( .A(n9338), .B(n9339), .Z(x[285]) );
  NAND U11899 ( .A(creg[285]), .B(init), .Z(n9338) );
  NAND U11900 ( .A(n9340), .B(n9341), .Z(x[284]) );
  NAND U11901 ( .A(creg[284]), .B(init), .Z(n9340) );
  NAND U11902 ( .A(n9342), .B(n9343), .Z(x[283]) );
  NAND U11903 ( .A(creg[283]), .B(init), .Z(n9342) );
  NAND U11904 ( .A(n9344), .B(n9345), .Z(x[282]) );
  NAND U11905 ( .A(creg[282]), .B(init), .Z(n9344) );
  NAND U11906 ( .A(n9346), .B(n9347), .Z(x[281]) );
  NAND U11907 ( .A(creg[281]), .B(init), .Z(n9346) );
  NAND U11908 ( .A(n9348), .B(n9349), .Z(x[280]) );
  NAND U11909 ( .A(creg[280]), .B(init), .Z(n9348) );
  NAND U11910 ( .A(n9350), .B(n9351), .Z(x[27]) );
  NAND U11911 ( .A(creg[27]), .B(init), .Z(n9350) );
  NAND U11912 ( .A(n9352), .B(n9353), .Z(x[279]) );
  NAND U11913 ( .A(creg[279]), .B(init), .Z(n9352) );
  NAND U11914 ( .A(n9354), .B(n9355), .Z(x[278]) );
  NAND U11915 ( .A(creg[278]), .B(init), .Z(n9354) );
  NAND U11916 ( .A(n9356), .B(n9357), .Z(x[277]) );
  NAND U11917 ( .A(creg[277]), .B(init), .Z(n9356) );
  NAND U11918 ( .A(n9358), .B(n9359), .Z(x[276]) );
  NAND U11919 ( .A(creg[276]), .B(init), .Z(n9358) );
  NAND U11920 ( .A(n9360), .B(n9361), .Z(x[275]) );
  NAND U11921 ( .A(creg[275]), .B(init), .Z(n9360) );
  NAND U11922 ( .A(n9362), .B(n9363), .Z(x[274]) );
  NAND U11923 ( .A(creg[274]), .B(init), .Z(n9362) );
  NAND U11924 ( .A(n9364), .B(n9365), .Z(x[273]) );
  NAND U11925 ( .A(creg[273]), .B(init), .Z(n9364) );
  NAND U11926 ( .A(n9366), .B(n9367), .Z(x[272]) );
  NAND U11927 ( .A(creg[272]), .B(init), .Z(n9366) );
  NAND U11928 ( .A(n9368), .B(n9369), .Z(x[271]) );
  NAND U11929 ( .A(creg[271]), .B(init), .Z(n9368) );
  NAND U11930 ( .A(n9370), .B(n9371), .Z(x[270]) );
  NAND U11931 ( .A(creg[270]), .B(init), .Z(n9370) );
  NAND U11932 ( .A(n9372), .B(n9373), .Z(x[26]) );
  NAND U11933 ( .A(creg[26]), .B(init), .Z(n9372) );
  NAND U11934 ( .A(n9374), .B(n9375), .Z(x[269]) );
  NAND U11935 ( .A(creg[269]), .B(init), .Z(n9374) );
  NAND U11936 ( .A(n9376), .B(n9377), .Z(x[268]) );
  NAND U11937 ( .A(creg[268]), .B(init), .Z(n9376) );
  NAND U11938 ( .A(n9378), .B(n9379), .Z(x[267]) );
  NAND U11939 ( .A(creg[267]), .B(init), .Z(n9378) );
  NAND U11940 ( .A(n9380), .B(n9381), .Z(x[266]) );
  NAND U11941 ( .A(creg[266]), .B(init), .Z(n9380) );
  NAND U11942 ( .A(n9382), .B(n9383), .Z(x[265]) );
  NAND U11943 ( .A(creg[265]), .B(init), .Z(n9382) );
  NAND U11944 ( .A(n9384), .B(n9385), .Z(x[264]) );
  NAND U11945 ( .A(creg[264]), .B(init), .Z(n9384) );
  NAND U11946 ( .A(n9386), .B(n9387), .Z(x[263]) );
  NAND U11947 ( .A(creg[263]), .B(init), .Z(n9386) );
  NAND U11948 ( .A(n9388), .B(n9389), .Z(x[262]) );
  NAND U11949 ( .A(creg[262]), .B(init), .Z(n9388) );
  NAND U11950 ( .A(n9390), .B(n9391), .Z(x[261]) );
  NAND U11951 ( .A(creg[261]), .B(init), .Z(n9390) );
  NAND U11952 ( .A(n9392), .B(n9393), .Z(x[260]) );
  NAND U11953 ( .A(creg[260]), .B(init), .Z(n9392) );
  NAND U11954 ( .A(n9394), .B(n9395), .Z(x[25]) );
  NAND U11955 ( .A(creg[25]), .B(init), .Z(n9394) );
  NAND U11956 ( .A(n9396), .B(n9397), .Z(x[259]) );
  NAND U11957 ( .A(creg[259]), .B(init), .Z(n9396) );
  NAND U11958 ( .A(n9398), .B(n9399), .Z(x[258]) );
  NAND U11959 ( .A(creg[258]), .B(init), .Z(n9398) );
  NAND U11960 ( .A(n9400), .B(n9401), .Z(x[257]) );
  NAND U11961 ( .A(creg[257]), .B(init), .Z(n9400) );
  NAND U11962 ( .A(n9402), .B(n9403), .Z(x[256]) );
  NAND U11963 ( .A(creg[256]), .B(init), .Z(n9402) );
  NAND U11964 ( .A(n9404), .B(n9405), .Z(x[255]) );
  NAND U11965 ( .A(creg[255]), .B(init), .Z(n9404) );
  NAND U11966 ( .A(n9406), .B(n9407), .Z(x[254]) );
  NAND U11967 ( .A(creg[254]), .B(init), .Z(n9406) );
  NAND U11968 ( .A(n9408), .B(n9409), .Z(x[253]) );
  NAND U11969 ( .A(creg[253]), .B(init), .Z(n9408) );
  NAND U11970 ( .A(n9410), .B(n9411), .Z(x[252]) );
  NAND U11971 ( .A(creg[252]), .B(init), .Z(n9410) );
  NAND U11972 ( .A(n9412), .B(n9413), .Z(x[251]) );
  NAND U11973 ( .A(creg[251]), .B(init), .Z(n9412) );
  NAND U11974 ( .A(n9414), .B(n9415), .Z(x[250]) );
  NAND U11975 ( .A(creg[250]), .B(init), .Z(n9414) );
  NAND U11976 ( .A(n9416), .B(n9417), .Z(x[24]) );
  NAND U11977 ( .A(creg[24]), .B(init), .Z(n9416) );
  NAND U11978 ( .A(n9418), .B(n9419), .Z(x[249]) );
  NAND U11979 ( .A(creg[249]), .B(init), .Z(n9418) );
  NAND U11980 ( .A(n9420), .B(n9421), .Z(x[248]) );
  NAND U11981 ( .A(creg[248]), .B(init), .Z(n9420) );
  NAND U11982 ( .A(n9422), .B(n9423), .Z(x[247]) );
  NAND U11983 ( .A(creg[247]), .B(init), .Z(n9422) );
  NAND U11984 ( .A(n9424), .B(n9425), .Z(x[246]) );
  NAND U11985 ( .A(creg[246]), .B(init), .Z(n9424) );
  NAND U11986 ( .A(n9426), .B(n9427), .Z(x[245]) );
  NAND U11987 ( .A(creg[245]), .B(init), .Z(n9426) );
  NAND U11988 ( .A(n9428), .B(n9429), .Z(x[244]) );
  NAND U11989 ( .A(creg[244]), .B(init), .Z(n9428) );
  NAND U11990 ( .A(n9430), .B(n9431), .Z(x[243]) );
  NAND U11991 ( .A(creg[243]), .B(init), .Z(n9430) );
  NAND U11992 ( .A(n9432), .B(n9433), .Z(x[242]) );
  NAND U11993 ( .A(creg[242]), .B(init), .Z(n9432) );
  NAND U11994 ( .A(n9434), .B(n9435), .Z(x[241]) );
  NAND U11995 ( .A(creg[241]), .B(init), .Z(n9434) );
  NAND U11996 ( .A(n9436), .B(n9437), .Z(x[240]) );
  NAND U11997 ( .A(creg[240]), .B(init), .Z(n9436) );
  NAND U11998 ( .A(n9438), .B(n9439), .Z(x[23]) );
  NAND U11999 ( .A(creg[23]), .B(init), .Z(n9438) );
  NAND U12000 ( .A(n9440), .B(n9441), .Z(x[239]) );
  NAND U12001 ( .A(creg[239]), .B(init), .Z(n9440) );
  NAND U12002 ( .A(n9442), .B(n9443), .Z(x[238]) );
  NAND U12003 ( .A(creg[238]), .B(init), .Z(n9442) );
  NAND U12004 ( .A(n9444), .B(n9445), .Z(x[237]) );
  NAND U12005 ( .A(creg[237]), .B(init), .Z(n9444) );
  NAND U12006 ( .A(n9446), .B(n9447), .Z(x[236]) );
  NAND U12007 ( .A(creg[236]), .B(init), .Z(n9446) );
  NAND U12008 ( .A(n9448), .B(n9449), .Z(x[235]) );
  NAND U12009 ( .A(creg[235]), .B(init), .Z(n9448) );
  NAND U12010 ( .A(n9450), .B(n9451), .Z(x[234]) );
  NAND U12011 ( .A(creg[234]), .B(init), .Z(n9450) );
  NAND U12012 ( .A(n9452), .B(n9453), .Z(x[233]) );
  NAND U12013 ( .A(creg[233]), .B(init), .Z(n9452) );
  NAND U12014 ( .A(n9454), .B(n9455), .Z(x[232]) );
  NAND U12015 ( .A(creg[232]), .B(init), .Z(n9454) );
  NAND U12016 ( .A(n9456), .B(n9457), .Z(x[231]) );
  NAND U12017 ( .A(creg[231]), .B(init), .Z(n9456) );
  NAND U12018 ( .A(n9458), .B(n9459), .Z(x[230]) );
  NAND U12019 ( .A(creg[230]), .B(init), .Z(n9458) );
  NAND U12020 ( .A(n9460), .B(n9461), .Z(x[22]) );
  NAND U12021 ( .A(creg[22]), .B(init), .Z(n9460) );
  NAND U12022 ( .A(n9462), .B(n9463), .Z(x[229]) );
  NAND U12023 ( .A(creg[229]), .B(init), .Z(n9462) );
  NAND U12024 ( .A(n9464), .B(n9465), .Z(x[228]) );
  NAND U12025 ( .A(creg[228]), .B(init), .Z(n9464) );
  NAND U12026 ( .A(n9466), .B(n9467), .Z(x[227]) );
  NAND U12027 ( .A(creg[227]), .B(init), .Z(n9466) );
  NAND U12028 ( .A(n9468), .B(n9469), .Z(x[226]) );
  NAND U12029 ( .A(creg[226]), .B(init), .Z(n9468) );
  NAND U12030 ( .A(n9470), .B(n9471), .Z(x[225]) );
  NAND U12031 ( .A(creg[225]), .B(init), .Z(n9470) );
  NAND U12032 ( .A(n9472), .B(n9473), .Z(x[224]) );
  NAND U12033 ( .A(creg[224]), .B(init), .Z(n9472) );
  NAND U12034 ( .A(n9474), .B(n9475), .Z(x[223]) );
  NAND U12035 ( .A(creg[223]), .B(init), .Z(n9474) );
  NAND U12036 ( .A(n9476), .B(n9477), .Z(x[222]) );
  NAND U12037 ( .A(creg[222]), .B(init), .Z(n9476) );
  NAND U12038 ( .A(n9478), .B(n9479), .Z(x[221]) );
  NAND U12039 ( .A(creg[221]), .B(init), .Z(n9478) );
  NAND U12040 ( .A(n9480), .B(n9481), .Z(x[220]) );
  NAND U12041 ( .A(creg[220]), .B(init), .Z(n9480) );
  NAND U12042 ( .A(n9482), .B(n9483), .Z(x[21]) );
  NAND U12043 ( .A(creg[21]), .B(init), .Z(n9482) );
  NAND U12044 ( .A(n9484), .B(n9485), .Z(x[219]) );
  NAND U12045 ( .A(creg[219]), .B(init), .Z(n9484) );
  NAND U12046 ( .A(n9486), .B(n9487), .Z(x[218]) );
  NAND U12047 ( .A(creg[218]), .B(init), .Z(n9486) );
  NAND U12048 ( .A(n9488), .B(n9489), .Z(x[217]) );
  NAND U12049 ( .A(creg[217]), .B(init), .Z(n9488) );
  NAND U12050 ( .A(n9490), .B(n9491), .Z(x[216]) );
  NAND U12051 ( .A(creg[216]), .B(init), .Z(n9490) );
  NAND U12052 ( .A(n9492), .B(n9493), .Z(x[215]) );
  NAND U12053 ( .A(creg[215]), .B(init), .Z(n9492) );
  NAND U12054 ( .A(n9494), .B(n9495), .Z(x[214]) );
  NAND U12055 ( .A(creg[214]), .B(init), .Z(n9494) );
  NAND U12056 ( .A(n9496), .B(n9497), .Z(x[213]) );
  NAND U12057 ( .A(creg[213]), .B(init), .Z(n9496) );
  NAND U12058 ( .A(n9498), .B(n9499), .Z(x[212]) );
  NAND U12059 ( .A(creg[212]), .B(init), .Z(n9498) );
  NAND U12060 ( .A(n9500), .B(n9501), .Z(x[211]) );
  NAND U12061 ( .A(creg[211]), .B(init), .Z(n9500) );
  NAND U12062 ( .A(n9502), .B(n9503), .Z(x[210]) );
  NAND U12063 ( .A(creg[210]), .B(init), .Z(n9502) );
  NAND U12064 ( .A(n9504), .B(n9505), .Z(x[20]) );
  NAND U12065 ( .A(creg[20]), .B(init), .Z(n9504) );
  NAND U12066 ( .A(n9506), .B(n9507), .Z(x[209]) );
  NAND U12067 ( .A(creg[209]), .B(init), .Z(n9506) );
  NAND U12068 ( .A(n9508), .B(n9509), .Z(x[208]) );
  NAND U12069 ( .A(creg[208]), .B(init), .Z(n9508) );
  NAND U12070 ( .A(n9510), .B(n9511), .Z(x[207]) );
  NAND U12071 ( .A(creg[207]), .B(init), .Z(n9510) );
  NAND U12072 ( .A(n9512), .B(n9513), .Z(x[206]) );
  NAND U12073 ( .A(creg[206]), .B(init), .Z(n9512) );
  NAND U12074 ( .A(n9514), .B(n9515), .Z(x[205]) );
  NAND U12075 ( .A(creg[205]), .B(init), .Z(n9514) );
  NAND U12076 ( .A(n9516), .B(n9517), .Z(x[204]) );
  NAND U12077 ( .A(creg[204]), .B(init), .Z(n9516) );
  NAND U12078 ( .A(n9518), .B(n9519), .Z(x[203]) );
  NAND U12079 ( .A(creg[203]), .B(init), .Z(n9518) );
  NAND U12080 ( .A(n9520), .B(n9521), .Z(x[202]) );
  NAND U12081 ( .A(creg[202]), .B(init), .Z(n9520) );
  NAND U12082 ( .A(n9522), .B(n9523), .Z(x[201]) );
  NAND U12083 ( .A(creg[201]), .B(init), .Z(n9522) );
  NAND U12084 ( .A(n9524), .B(n9525), .Z(x[200]) );
  NAND U12085 ( .A(creg[200]), .B(init), .Z(n9524) );
  NAND U12086 ( .A(n9526), .B(n9527), .Z(x[1]) );
  NAND U12087 ( .A(creg[1]), .B(init), .Z(n9526) );
  NAND U12088 ( .A(n9528), .B(n9529), .Z(x[19]) );
  NAND U12089 ( .A(creg[19]), .B(init), .Z(n9528) );
  NAND U12090 ( .A(n9530), .B(n9531), .Z(x[199]) );
  NAND U12091 ( .A(creg[199]), .B(init), .Z(n9530) );
  NAND U12092 ( .A(n9532), .B(n9533), .Z(x[198]) );
  NAND U12093 ( .A(creg[198]), .B(init), .Z(n9532) );
  NAND U12094 ( .A(n9534), .B(n9535), .Z(x[197]) );
  NAND U12095 ( .A(creg[197]), .B(init), .Z(n9534) );
  NAND U12096 ( .A(n9536), .B(n9537), .Z(x[196]) );
  NAND U12097 ( .A(creg[196]), .B(init), .Z(n9536) );
  NAND U12098 ( .A(n9538), .B(n9539), .Z(x[195]) );
  NAND U12099 ( .A(creg[195]), .B(init), .Z(n9538) );
  NAND U12100 ( .A(n9540), .B(n9541), .Z(x[194]) );
  NAND U12101 ( .A(creg[194]), .B(init), .Z(n9540) );
  NAND U12102 ( .A(n9542), .B(n9543), .Z(x[193]) );
  NAND U12103 ( .A(creg[193]), .B(init), .Z(n9542) );
  NAND U12104 ( .A(n9544), .B(n9545), .Z(x[192]) );
  NAND U12105 ( .A(creg[192]), .B(init), .Z(n9544) );
  NAND U12106 ( .A(n9546), .B(n9547), .Z(x[191]) );
  NAND U12107 ( .A(creg[191]), .B(init), .Z(n9546) );
  NAND U12108 ( .A(n9548), .B(n9549), .Z(x[190]) );
  NAND U12109 ( .A(creg[190]), .B(init), .Z(n9548) );
  NAND U12110 ( .A(n9550), .B(n9551), .Z(x[18]) );
  NAND U12111 ( .A(creg[18]), .B(init), .Z(n9550) );
  NAND U12112 ( .A(n9552), .B(n9553), .Z(x[189]) );
  NAND U12113 ( .A(creg[189]), .B(init), .Z(n9552) );
  NAND U12114 ( .A(n9554), .B(n9555), .Z(x[188]) );
  NAND U12115 ( .A(creg[188]), .B(init), .Z(n9554) );
  NAND U12116 ( .A(n9556), .B(n9557), .Z(x[187]) );
  NAND U12117 ( .A(creg[187]), .B(init), .Z(n9556) );
  NAND U12118 ( .A(n9558), .B(n9559), .Z(x[186]) );
  NAND U12119 ( .A(creg[186]), .B(init), .Z(n9558) );
  NAND U12120 ( .A(n9560), .B(n9561), .Z(x[185]) );
  NAND U12121 ( .A(creg[185]), .B(init), .Z(n9560) );
  NAND U12122 ( .A(n9562), .B(n9563), .Z(x[184]) );
  NAND U12123 ( .A(creg[184]), .B(init), .Z(n9562) );
  NAND U12124 ( .A(n9564), .B(n9565), .Z(x[183]) );
  NAND U12125 ( .A(creg[183]), .B(init), .Z(n9564) );
  NAND U12126 ( .A(n9566), .B(n9567), .Z(x[182]) );
  NAND U12127 ( .A(creg[182]), .B(init), .Z(n9566) );
  NAND U12128 ( .A(n9568), .B(n9569), .Z(x[181]) );
  NAND U12129 ( .A(creg[181]), .B(init), .Z(n9568) );
  NAND U12130 ( .A(n9570), .B(n9571), .Z(x[180]) );
  NAND U12131 ( .A(creg[180]), .B(init), .Z(n9570) );
  NAND U12132 ( .A(n9572), .B(n9573), .Z(x[17]) );
  NAND U12133 ( .A(creg[17]), .B(init), .Z(n9572) );
  NAND U12134 ( .A(n9574), .B(n9575), .Z(x[179]) );
  NAND U12135 ( .A(creg[179]), .B(init), .Z(n9574) );
  NAND U12136 ( .A(n9576), .B(n9577), .Z(x[178]) );
  NAND U12137 ( .A(creg[178]), .B(init), .Z(n9576) );
  NAND U12138 ( .A(n9578), .B(n9579), .Z(x[177]) );
  NAND U12139 ( .A(creg[177]), .B(init), .Z(n9578) );
  NAND U12140 ( .A(n9580), .B(n9581), .Z(x[176]) );
  NAND U12141 ( .A(creg[176]), .B(init), .Z(n9580) );
  NAND U12142 ( .A(n9582), .B(n9583), .Z(x[175]) );
  NAND U12143 ( .A(creg[175]), .B(init), .Z(n9582) );
  NAND U12144 ( .A(n9584), .B(n9585), .Z(x[174]) );
  NAND U12145 ( .A(creg[174]), .B(init), .Z(n9584) );
  NAND U12146 ( .A(n9586), .B(n9587), .Z(x[173]) );
  NAND U12147 ( .A(creg[173]), .B(init), .Z(n9586) );
  NAND U12148 ( .A(n9588), .B(n9589), .Z(x[172]) );
  NAND U12149 ( .A(creg[172]), .B(init), .Z(n9588) );
  NAND U12150 ( .A(n9590), .B(n9591), .Z(x[171]) );
  NAND U12151 ( .A(creg[171]), .B(init), .Z(n9590) );
  NAND U12152 ( .A(n9592), .B(n9593), .Z(x[170]) );
  NAND U12153 ( .A(creg[170]), .B(init), .Z(n9592) );
  NAND U12154 ( .A(n9594), .B(n9595), .Z(x[16]) );
  NAND U12155 ( .A(creg[16]), .B(init), .Z(n9594) );
  NAND U12156 ( .A(n9596), .B(n9597), .Z(x[169]) );
  NAND U12157 ( .A(creg[169]), .B(init), .Z(n9596) );
  NAND U12158 ( .A(n9598), .B(n9599), .Z(x[168]) );
  NAND U12159 ( .A(creg[168]), .B(init), .Z(n9598) );
  NAND U12160 ( .A(n9600), .B(n9601), .Z(x[167]) );
  NAND U12161 ( .A(creg[167]), .B(init), .Z(n9600) );
  NAND U12162 ( .A(n9602), .B(n9603), .Z(x[166]) );
  NAND U12163 ( .A(creg[166]), .B(init), .Z(n9602) );
  NAND U12164 ( .A(n9604), .B(n9605), .Z(x[165]) );
  NAND U12165 ( .A(creg[165]), .B(init), .Z(n9604) );
  NAND U12166 ( .A(n9606), .B(n9607), .Z(x[164]) );
  NAND U12167 ( .A(creg[164]), .B(init), .Z(n9606) );
  NAND U12168 ( .A(n9608), .B(n9609), .Z(x[163]) );
  NAND U12169 ( .A(creg[163]), .B(init), .Z(n9608) );
  NAND U12170 ( .A(n9610), .B(n9611), .Z(x[162]) );
  NAND U12171 ( .A(creg[162]), .B(init), .Z(n9610) );
  NAND U12172 ( .A(n9612), .B(n9613), .Z(x[161]) );
  NAND U12173 ( .A(creg[161]), .B(init), .Z(n9612) );
  NAND U12174 ( .A(n9614), .B(n9615), .Z(x[160]) );
  NAND U12175 ( .A(creg[160]), .B(init), .Z(n9614) );
  NAND U12176 ( .A(n9616), .B(n9617), .Z(x[15]) );
  NAND U12177 ( .A(creg[15]), .B(init), .Z(n9616) );
  NAND U12178 ( .A(n9618), .B(n9619), .Z(x[159]) );
  NAND U12179 ( .A(creg[159]), .B(init), .Z(n9618) );
  NAND U12180 ( .A(n9620), .B(n9621), .Z(x[158]) );
  NAND U12181 ( .A(creg[158]), .B(init), .Z(n9620) );
  NAND U12182 ( .A(n9622), .B(n9623), .Z(x[157]) );
  NAND U12183 ( .A(creg[157]), .B(init), .Z(n9622) );
  NAND U12184 ( .A(n9624), .B(n9625), .Z(x[156]) );
  NAND U12185 ( .A(creg[156]), .B(init), .Z(n9624) );
  NAND U12186 ( .A(n9626), .B(n9627), .Z(x[155]) );
  NAND U12187 ( .A(creg[155]), .B(init), .Z(n9626) );
  NAND U12188 ( .A(n9628), .B(n9629), .Z(x[154]) );
  NAND U12189 ( .A(creg[154]), .B(init), .Z(n9628) );
  NAND U12190 ( .A(n9630), .B(n9631), .Z(x[153]) );
  NAND U12191 ( .A(creg[153]), .B(init), .Z(n9630) );
  NAND U12192 ( .A(n9632), .B(n9633), .Z(x[152]) );
  NAND U12193 ( .A(creg[152]), .B(init), .Z(n9632) );
  NAND U12194 ( .A(n9634), .B(n9635), .Z(x[151]) );
  NAND U12195 ( .A(creg[151]), .B(init), .Z(n9634) );
  NAND U12196 ( .A(n9636), .B(n9637), .Z(x[150]) );
  NAND U12197 ( .A(creg[150]), .B(init), .Z(n9636) );
  NAND U12198 ( .A(n9638), .B(n9639), .Z(x[14]) );
  NAND U12199 ( .A(creg[14]), .B(init), .Z(n9638) );
  NAND U12200 ( .A(n9640), .B(n9641), .Z(x[149]) );
  NAND U12201 ( .A(creg[149]), .B(init), .Z(n9640) );
  NAND U12202 ( .A(n9642), .B(n9643), .Z(x[148]) );
  NAND U12203 ( .A(creg[148]), .B(init), .Z(n9642) );
  NAND U12204 ( .A(n9644), .B(n9645), .Z(x[147]) );
  NAND U12205 ( .A(creg[147]), .B(init), .Z(n9644) );
  NAND U12206 ( .A(n9646), .B(n9647), .Z(x[146]) );
  NAND U12207 ( .A(creg[146]), .B(init), .Z(n9646) );
  NAND U12208 ( .A(n9648), .B(n9649), .Z(x[145]) );
  NAND U12209 ( .A(creg[145]), .B(init), .Z(n9648) );
  NAND U12210 ( .A(n9650), .B(n9651), .Z(x[144]) );
  NAND U12211 ( .A(creg[144]), .B(init), .Z(n9650) );
  NAND U12212 ( .A(n9652), .B(n9653), .Z(x[143]) );
  NAND U12213 ( .A(creg[143]), .B(init), .Z(n9652) );
  NAND U12214 ( .A(n9654), .B(n9655), .Z(x[142]) );
  NAND U12215 ( .A(creg[142]), .B(init), .Z(n9654) );
  NAND U12216 ( .A(n9656), .B(n9657), .Z(x[141]) );
  NAND U12217 ( .A(creg[141]), .B(init), .Z(n9656) );
  NAND U12218 ( .A(n9658), .B(n9659), .Z(x[140]) );
  NAND U12219 ( .A(creg[140]), .B(init), .Z(n9658) );
  NAND U12220 ( .A(n9660), .B(n9661), .Z(x[13]) );
  NAND U12221 ( .A(creg[13]), .B(init), .Z(n9660) );
  NAND U12222 ( .A(n9662), .B(n9663), .Z(x[139]) );
  NAND U12223 ( .A(creg[139]), .B(init), .Z(n9662) );
  NAND U12224 ( .A(n9664), .B(n9665), .Z(x[138]) );
  NAND U12225 ( .A(creg[138]), .B(init), .Z(n9664) );
  NAND U12226 ( .A(n9666), .B(n9667), .Z(x[137]) );
  NAND U12227 ( .A(creg[137]), .B(init), .Z(n9666) );
  NAND U12228 ( .A(n9668), .B(n9669), .Z(x[136]) );
  NAND U12229 ( .A(creg[136]), .B(init), .Z(n9668) );
  NAND U12230 ( .A(n9670), .B(n9671), .Z(x[135]) );
  NAND U12231 ( .A(creg[135]), .B(init), .Z(n9670) );
  NAND U12232 ( .A(n9672), .B(n9673), .Z(x[134]) );
  NAND U12233 ( .A(creg[134]), .B(init), .Z(n9672) );
  NAND U12234 ( .A(n9674), .B(n9675), .Z(x[133]) );
  NAND U12235 ( .A(creg[133]), .B(init), .Z(n9674) );
  NAND U12236 ( .A(n9676), .B(n9677), .Z(x[132]) );
  NAND U12237 ( .A(creg[132]), .B(init), .Z(n9676) );
  NAND U12238 ( .A(n9678), .B(n9679), .Z(x[131]) );
  NAND U12239 ( .A(creg[131]), .B(init), .Z(n9678) );
  NAND U12240 ( .A(n9680), .B(n9681), .Z(x[130]) );
  NAND U12241 ( .A(creg[130]), .B(init), .Z(n9680) );
  NAND U12242 ( .A(n9682), .B(n9683), .Z(x[12]) );
  NAND U12243 ( .A(creg[12]), .B(init), .Z(n9682) );
  NAND U12244 ( .A(n9684), .B(n9685), .Z(x[129]) );
  NAND U12245 ( .A(creg[129]), .B(init), .Z(n9684) );
  NAND U12246 ( .A(n9686), .B(n9687), .Z(x[128]) );
  NAND U12247 ( .A(creg[128]), .B(init), .Z(n9686) );
  NAND U12248 ( .A(n9688), .B(n9689), .Z(x[127]) );
  NAND U12249 ( .A(creg[127]), .B(init), .Z(n9688) );
  NAND U12250 ( .A(n9690), .B(n9691), .Z(x[126]) );
  NAND U12251 ( .A(creg[126]), .B(init), .Z(n9690) );
  NAND U12252 ( .A(n9692), .B(n9693), .Z(x[125]) );
  NAND U12253 ( .A(creg[125]), .B(init), .Z(n9692) );
  NAND U12254 ( .A(n9694), .B(n9695), .Z(x[124]) );
  NAND U12255 ( .A(creg[124]), .B(init), .Z(n9694) );
  NAND U12256 ( .A(n9696), .B(n9697), .Z(x[123]) );
  NAND U12257 ( .A(creg[123]), .B(init), .Z(n9696) );
  NAND U12258 ( .A(n9698), .B(n9699), .Z(x[122]) );
  NAND U12259 ( .A(creg[122]), .B(init), .Z(n9698) );
  NAND U12260 ( .A(n9700), .B(n9701), .Z(x[121]) );
  NAND U12261 ( .A(creg[121]), .B(init), .Z(n9700) );
  NAND U12262 ( .A(n9702), .B(n9703), .Z(x[120]) );
  NAND U12263 ( .A(creg[120]), .B(init), .Z(n9702) );
  NAND U12264 ( .A(n9704), .B(n9705), .Z(x[11]) );
  NAND U12265 ( .A(creg[11]), .B(init), .Z(n9704) );
  NAND U12266 ( .A(n9706), .B(n9707), .Z(x[119]) );
  NAND U12267 ( .A(creg[119]), .B(init), .Z(n9706) );
  NAND U12268 ( .A(n9708), .B(n9709), .Z(x[118]) );
  NAND U12269 ( .A(creg[118]), .B(init), .Z(n9708) );
  NAND U12270 ( .A(n9710), .B(n9711), .Z(x[117]) );
  NAND U12271 ( .A(creg[117]), .B(init), .Z(n9710) );
  NAND U12272 ( .A(n9712), .B(n9713), .Z(x[116]) );
  NAND U12273 ( .A(creg[116]), .B(init), .Z(n9712) );
  NAND U12274 ( .A(n9714), .B(n9715), .Z(x[115]) );
  NAND U12275 ( .A(creg[115]), .B(init), .Z(n9714) );
  NAND U12276 ( .A(n9716), .B(n9717), .Z(x[114]) );
  NAND U12277 ( .A(creg[114]), .B(init), .Z(n9716) );
  NAND U12278 ( .A(n9718), .B(n9719), .Z(x[113]) );
  NAND U12279 ( .A(creg[113]), .B(init), .Z(n9718) );
  NAND U12280 ( .A(n9720), .B(n9721), .Z(x[112]) );
  NAND U12281 ( .A(creg[112]), .B(init), .Z(n9720) );
  NAND U12282 ( .A(n9722), .B(n9723), .Z(x[111]) );
  NAND U12283 ( .A(creg[111]), .B(init), .Z(n9722) );
  NAND U12284 ( .A(n9724), .B(n9725), .Z(x[110]) );
  NAND U12285 ( .A(creg[110]), .B(init), .Z(n9724) );
  NAND U12286 ( .A(n9726), .B(n9727), .Z(x[10]) );
  NAND U12287 ( .A(creg[10]), .B(init), .Z(n9726) );
  NAND U12288 ( .A(n9728), .B(n9729), .Z(x[109]) );
  NAND U12289 ( .A(creg[109]), .B(init), .Z(n9728) );
  NAND U12290 ( .A(n9730), .B(n9731), .Z(x[108]) );
  NAND U12291 ( .A(creg[108]), .B(init), .Z(n9730) );
  NAND U12292 ( .A(n9732), .B(n9733), .Z(x[107]) );
  NAND U12293 ( .A(creg[107]), .B(init), .Z(n9732) );
  NAND U12294 ( .A(n9734), .B(n9735), .Z(x[106]) );
  NAND U12295 ( .A(creg[106]), .B(init), .Z(n9734) );
  NAND U12296 ( .A(n9736), .B(n9737), .Z(x[105]) );
  NAND U12297 ( .A(creg[105]), .B(init), .Z(n9736) );
  NAND U12298 ( .A(n9738), .B(n9739), .Z(x[104]) );
  NAND U12299 ( .A(creg[104]), .B(init), .Z(n9738) );
  NAND U12300 ( .A(n9740), .B(n9741), .Z(x[103]) );
  NAND U12301 ( .A(creg[103]), .B(init), .Z(n9740) );
  NAND U12302 ( .A(n9742), .B(n9743), .Z(x[102]) );
  NAND U12303 ( .A(creg[102]), .B(init), .Z(n9742) );
  NAND U12304 ( .A(n9744), .B(n9745), .Z(x[101]) );
  NAND U12305 ( .A(creg[101]), .B(init), .Z(n9744) );
  NAND U12306 ( .A(n9746), .B(n9747), .Z(x[100]) );
  NAND U12307 ( .A(creg[100]), .B(init), .Z(n9746) );
  NAND U12308 ( .A(n9748), .B(n9749), .Z(x[0]) );
  NAND U12309 ( .A(creg[0]), .B(init), .Z(n9748) );
  AND U12310 ( .A(start_reg[9]), .B(init), .Z(start_in[9]) );
  AND U12311 ( .A(start_reg[99]), .B(init), .Z(start_in[99]) );
  AND U12312 ( .A(start_reg[98]), .B(init), .Z(start_in[98]) );
  AND U12313 ( .A(start_reg[97]), .B(init), .Z(start_in[97]) );
  AND U12314 ( .A(start_reg[96]), .B(init), .Z(start_in[96]) );
  AND U12315 ( .A(start_reg[95]), .B(init), .Z(start_in[95]) );
  AND U12316 ( .A(start_reg[94]), .B(init), .Z(start_in[94]) );
  AND U12317 ( .A(start_reg[93]), .B(init), .Z(start_in[93]) );
  AND U12318 ( .A(start_reg[92]), .B(init), .Z(start_in[92]) );
  AND U12319 ( .A(start_reg[91]), .B(init), .Z(start_in[91]) );
  AND U12320 ( .A(start_reg[90]), .B(init), .Z(start_in[90]) );
  AND U12321 ( .A(start_reg[8]), .B(init), .Z(start_in[8]) );
  AND U12322 ( .A(start_reg[89]), .B(init), .Z(start_in[89]) );
  AND U12323 ( .A(start_reg[88]), .B(init), .Z(start_in[88]) );
  AND U12324 ( .A(start_reg[87]), .B(init), .Z(start_in[87]) );
  AND U12325 ( .A(start_reg[86]), .B(init), .Z(start_in[86]) );
  AND U12326 ( .A(start_reg[85]), .B(init), .Z(start_in[85]) );
  AND U12327 ( .A(start_reg[84]), .B(init), .Z(start_in[84]) );
  AND U12328 ( .A(start_reg[83]), .B(init), .Z(start_in[83]) );
  AND U12329 ( .A(start_reg[82]), .B(init), .Z(start_in[82]) );
  AND U12330 ( .A(start_reg[81]), .B(init), .Z(start_in[81]) );
  AND U12331 ( .A(start_reg[80]), .B(init), .Z(start_in[80]) );
  AND U12332 ( .A(start_reg[7]), .B(init), .Z(start_in[7]) );
  AND U12333 ( .A(start_reg[79]), .B(init), .Z(start_in[79]) );
  AND U12334 ( .A(start_reg[78]), .B(init), .Z(start_in[78]) );
  AND U12335 ( .A(start_reg[77]), .B(init), .Z(start_in[77]) );
  AND U12336 ( .A(start_reg[76]), .B(init), .Z(start_in[76]) );
  AND U12337 ( .A(start_reg[75]), .B(init), .Z(start_in[75]) );
  AND U12338 ( .A(start_reg[74]), .B(init), .Z(start_in[74]) );
  AND U12339 ( .A(start_reg[73]), .B(init), .Z(start_in[73]) );
  AND U12340 ( .A(start_reg[72]), .B(init), .Z(start_in[72]) );
  AND U12341 ( .A(start_reg[71]), .B(init), .Z(start_in[71]) );
  AND U12342 ( .A(start_reg[70]), .B(init), .Z(start_in[70]) );
  AND U12343 ( .A(start_reg[6]), .B(init), .Z(start_in[6]) );
  AND U12344 ( .A(start_reg[69]), .B(init), .Z(start_in[69]) );
  AND U12345 ( .A(start_reg[68]), .B(init), .Z(start_in[68]) );
  AND U12346 ( .A(start_reg[67]), .B(init), .Z(start_in[67]) );
  AND U12347 ( .A(start_reg[66]), .B(init), .Z(start_in[66]) );
  AND U12348 ( .A(start_reg[65]), .B(init), .Z(start_in[65]) );
  AND U12349 ( .A(start_reg[64]), .B(init), .Z(start_in[64]) );
  AND U12350 ( .A(start_reg[63]), .B(init), .Z(start_in[63]) );
  AND U12351 ( .A(start_reg[62]), .B(init), .Z(start_in[62]) );
  AND U12352 ( .A(start_reg[61]), .B(init), .Z(start_in[61]) );
  AND U12353 ( .A(start_reg[60]), .B(init), .Z(start_in[60]) );
  AND U12354 ( .A(start_reg[5]), .B(init), .Z(start_in[5]) );
  AND U12355 ( .A(start_reg[59]), .B(init), .Z(start_in[59]) );
  AND U12356 ( .A(start_reg[58]), .B(init), .Z(start_in[58]) );
  AND U12357 ( .A(start_reg[57]), .B(init), .Z(start_in[57]) );
  AND U12358 ( .A(start_reg[56]), .B(init), .Z(start_in[56]) );
  AND U12359 ( .A(start_reg[55]), .B(init), .Z(start_in[55]) );
  AND U12360 ( .A(start_reg[54]), .B(init), .Z(start_in[54]) );
  AND U12361 ( .A(start_reg[53]), .B(init), .Z(start_in[53]) );
  AND U12362 ( .A(start_reg[52]), .B(init), .Z(start_in[52]) );
  AND U12363 ( .A(start_reg[51]), .B(init), .Z(start_in[51]) );
  AND U12364 ( .A(start_reg[510]), .B(init), .Z(start_in[510]) );
  AND U12365 ( .A(start_reg[50]), .B(init), .Z(start_in[50]) );
  AND U12366 ( .A(start_reg[509]), .B(init), .Z(start_in[509]) );
  AND U12367 ( .A(start_reg[508]), .B(init), .Z(start_in[508]) );
  AND U12368 ( .A(start_reg[507]), .B(init), .Z(start_in[507]) );
  AND U12369 ( .A(start_reg[506]), .B(init), .Z(start_in[506]) );
  AND U12370 ( .A(start_reg[505]), .B(init), .Z(start_in[505]) );
  AND U12371 ( .A(start_reg[504]), .B(init), .Z(start_in[504]) );
  AND U12372 ( .A(start_reg[503]), .B(init), .Z(start_in[503]) );
  AND U12373 ( .A(start_reg[502]), .B(init), .Z(start_in[502]) );
  AND U12374 ( .A(start_reg[501]), .B(init), .Z(start_in[501]) );
  AND U12375 ( .A(start_reg[500]), .B(init), .Z(start_in[500]) );
  AND U12376 ( .A(start_reg[4]), .B(init), .Z(start_in[4]) );
  AND U12377 ( .A(start_reg[49]), .B(init), .Z(start_in[49]) );
  AND U12378 ( .A(start_reg[499]), .B(init), .Z(start_in[499]) );
  AND U12379 ( .A(start_reg[498]), .B(init), .Z(start_in[498]) );
  AND U12380 ( .A(start_reg[497]), .B(init), .Z(start_in[497]) );
  AND U12381 ( .A(start_reg[496]), .B(init), .Z(start_in[496]) );
  AND U12382 ( .A(start_reg[495]), .B(init), .Z(start_in[495]) );
  AND U12383 ( .A(start_reg[494]), .B(init), .Z(start_in[494]) );
  AND U12384 ( .A(start_reg[493]), .B(init), .Z(start_in[493]) );
  AND U12385 ( .A(start_reg[492]), .B(init), .Z(start_in[492]) );
  AND U12386 ( .A(start_reg[491]), .B(init), .Z(start_in[491]) );
  AND U12387 ( .A(start_reg[490]), .B(init), .Z(start_in[490]) );
  AND U12388 ( .A(start_reg[48]), .B(init), .Z(start_in[48]) );
  AND U12389 ( .A(start_reg[489]), .B(init), .Z(start_in[489]) );
  AND U12390 ( .A(start_reg[488]), .B(init), .Z(start_in[488]) );
  AND U12391 ( .A(start_reg[487]), .B(init), .Z(start_in[487]) );
  AND U12392 ( .A(start_reg[486]), .B(init), .Z(start_in[486]) );
  AND U12393 ( .A(start_reg[485]), .B(init), .Z(start_in[485]) );
  AND U12394 ( .A(start_reg[484]), .B(init), .Z(start_in[484]) );
  AND U12395 ( .A(start_reg[483]), .B(init), .Z(start_in[483]) );
  AND U12396 ( .A(start_reg[482]), .B(init), .Z(start_in[482]) );
  AND U12397 ( .A(start_reg[481]), .B(init), .Z(start_in[481]) );
  AND U12398 ( .A(start_reg[480]), .B(init), .Z(start_in[480]) );
  AND U12399 ( .A(start_reg[47]), .B(init), .Z(start_in[47]) );
  AND U12400 ( .A(start_reg[479]), .B(init), .Z(start_in[479]) );
  AND U12401 ( .A(start_reg[478]), .B(init), .Z(start_in[478]) );
  AND U12402 ( .A(start_reg[477]), .B(init), .Z(start_in[477]) );
  AND U12403 ( .A(start_reg[476]), .B(init), .Z(start_in[476]) );
  AND U12404 ( .A(start_reg[475]), .B(init), .Z(start_in[475]) );
  AND U12405 ( .A(start_reg[474]), .B(init), .Z(start_in[474]) );
  AND U12406 ( .A(start_reg[473]), .B(init), .Z(start_in[473]) );
  AND U12407 ( .A(start_reg[472]), .B(init), .Z(start_in[472]) );
  AND U12408 ( .A(start_reg[471]), .B(init), .Z(start_in[471]) );
  AND U12409 ( .A(start_reg[470]), .B(init), .Z(start_in[470]) );
  AND U12410 ( .A(start_reg[46]), .B(init), .Z(start_in[46]) );
  AND U12411 ( .A(start_reg[469]), .B(init), .Z(start_in[469]) );
  AND U12412 ( .A(start_reg[468]), .B(init), .Z(start_in[468]) );
  AND U12413 ( .A(start_reg[467]), .B(init), .Z(start_in[467]) );
  AND U12414 ( .A(start_reg[466]), .B(init), .Z(start_in[466]) );
  AND U12415 ( .A(start_reg[465]), .B(init), .Z(start_in[465]) );
  AND U12416 ( .A(start_reg[464]), .B(init), .Z(start_in[464]) );
  AND U12417 ( .A(start_reg[463]), .B(init), .Z(start_in[463]) );
  AND U12418 ( .A(start_reg[462]), .B(init), .Z(start_in[462]) );
  AND U12419 ( .A(start_reg[461]), .B(init), .Z(start_in[461]) );
  AND U12420 ( .A(start_reg[460]), .B(init), .Z(start_in[460]) );
  AND U12421 ( .A(start_reg[45]), .B(init), .Z(start_in[45]) );
  AND U12422 ( .A(start_reg[459]), .B(init), .Z(start_in[459]) );
  AND U12423 ( .A(start_reg[458]), .B(init), .Z(start_in[458]) );
  AND U12424 ( .A(start_reg[457]), .B(init), .Z(start_in[457]) );
  AND U12425 ( .A(start_reg[456]), .B(init), .Z(start_in[456]) );
  AND U12426 ( .A(start_reg[455]), .B(init), .Z(start_in[455]) );
  AND U12427 ( .A(start_reg[454]), .B(init), .Z(start_in[454]) );
  AND U12428 ( .A(start_reg[453]), .B(init), .Z(start_in[453]) );
  AND U12429 ( .A(start_reg[452]), .B(init), .Z(start_in[452]) );
  AND U12430 ( .A(start_reg[451]), .B(init), .Z(start_in[451]) );
  AND U12431 ( .A(start_reg[450]), .B(init), .Z(start_in[450]) );
  AND U12432 ( .A(start_reg[44]), .B(init), .Z(start_in[44]) );
  AND U12433 ( .A(start_reg[449]), .B(init), .Z(start_in[449]) );
  AND U12434 ( .A(start_reg[448]), .B(init), .Z(start_in[448]) );
  AND U12435 ( .A(start_reg[447]), .B(init), .Z(start_in[447]) );
  AND U12436 ( .A(start_reg[446]), .B(init), .Z(start_in[446]) );
  AND U12437 ( .A(start_reg[445]), .B(init), .Z(start_in[445]) );
  AND U12438 ( .A(start_reg[444]), .B(init), .Z(start_in[444]) );
  AND U12439 ( .A(start_reg[443]), .B(init), .Z(start_in[443]) );
  AND U12440 ( .A(start_reg[442]), .B(init), .Z(start_in[442]) );
  AND U12441 ( .A(start_reg[441]), .B(init), .Z(start_in[441]) );
  AND U12442 ( .A(start_reg[440]), .B(init), .Z(start_in[440]) );
  AND U12443 ( .A(start_reg[43]), .B(init), .Z(start_in[43]) );
  AND U12444 ( .A(start_reg[439]), .B(init), .Z(start_in[439]) );
  AND U12445 ( .A(start_reg[438]), .B(init), .Z(start_in[438]) );
  AND U12446 ( .A(start_reg[437]), .B(init), .Z(start_in[437]) );
  AND U12447 ( .A(start_reg[436]), .B(init), .Z(start_in[436]) );
  AND U12448 ( .A(start_reg[435]), .B(init), .Z(start_in[435]) );
  AND U12449 ( .A(start_reg[434]), .B(init), .Z(start_in[434]) );
  AND U12450 ( .A(start_reg[433]), .B(init), .Z(start_in[433]) );
  AND U12451 ( .A(start_reg[432]), .B(init), .Z(start_in[432]) );
  AND U12452 ( .A(start_reg[431]), .B(init), .Z(start_in[431]) );
  AND U12453 ( .A(start_reg[430]), .B(init), .Z(start_in[430]) );
  AND U12454 ( .A(start_reg[42]), .B(init), .Z(start_in[42]) );
  AND U12455 ( .A(start_reg[429]), .B(init), .Z(start_in[429]) );
  AND U12456 ( .A(start_reg[428]), .B(init), .Z(start_in[428]) );
  AND U12457 ( .A(start_reg[427]), .B(init), .Z(start_in[427]) );
  AND U12458 ( .A(start_reg[426]), .B(init), .Z(start_in[426]) );
  AND U12459 ( .A(start_reg[425]), .B(init), .Z(start_in[425]) );
  AND U12460 ( .A(start_reg[424]), .B(init), .Z(start_in[424]) );
  AND U12461 ( .A(start_reg[423]), .B(init), .Z(start_in[423]) );
  AND U12462 ( .A(start_reg[422]), .B(init), .Z(start_in[422]) );
  AND U12463 ( .A(start_reg[421]), .B(init), .Z(start_in[421]) );
  AND U12464 ( .A(start_reg[420]), .B(init), .Z(start_in[420]) );
  AND U12465 ( .A(start_reg[41]), .B(init), .Z(start_in[41]) );
  AND U12466 ( .A(start_reg[419]), .B(init), .Z(start_in[419]) );
  AND U12467 ( .A(start_reg[418]), .B(init), .Z(start_in[418]) );
  AND U12468 ( .A(start_reg[417]), .B(init), .Z(start_in[417]) );
  AND U12469 ( .A(start_reg[416]), .B(init), .Z(start_in[416]) );
  AND U12470 ( .A(start_reg[415]), .B(init), .Z(start_in[415]) );
  AND U12471 ( .A(start_reg[414]), .B(init), .Z(start_in[414]) );
  AND U12472 ( .A(start_reg[413]), .B(init), .Z(start_in[413]) );
  AND U12473 ( .A(start_reg[412]), .B(init), .Z(start_in[412]) );
  AND U12474 ( .A(start_reg[411]), .B(init), .Z(start_in[411]) );
  AND U12475 ( .A(start_reg[410]), .B(init), .Z(start_in[410]) );
  AND U12476 ( .A(start_reg[40]), .B(init), .Z(start_in[40]) );
  AND U12477 ( .A(start_reg[409]), .B(init), .Z(start_in[409]) );
  AND U12478 ( .A(start_reg[408]), .B(init), .Z(start_in[408]) );
  AND U12479 ( .A(start_reg[407]), .B(init), .Z(start_in[407]) );
  AND U12480 ( .A(start_reg[406]), .B(init), .Z(start_in[406]) );
  AND U12481 ( .A(start_reg[405]), .B(init), .Z(start_in[405]) );
  AND U12482 ( .A(start_reg[404]), .B(init), .Z(start_in[404]) );
  AND U12483 ( .A(start_reg[403]), .B(init), .Z(start_in[403]) );
  AND U12484 ( .A(start_reg[402]), .B(init), .Z(start_in[402]) );
  AND U12485 ( .A(start_reg[401]), .B(init), .Z(start_in[401]) );
  AND U12486 ( .A(start_reg[400]), .B(init), .Z(start_in[400]) );
  AND U12487 ( .A(start_reg[3]), .B(init), .Z(start_in[3]) );
  AND U12488 ( .A(start_reg[39]), .B(init), .Z(start_in[39]) );
  AND U12489 ( .A(start_reg[399]), .B(init), .Z(start_in[399]) );
  AND U12490 ( .A(start_reg[398]), .B(init), .Z(start_in[398]) );
  AND U12491 ( .A(start_reg[397]), .B(init), .Z(start_in[397]) );
  AND U12492 ( .A(start_reg[396]), .B(init), .Z(start_in[396]) );
  AND U12493 ( .A(start_reg[395]), .B(init), .Z(start_in[395]) );
  AND U12494 ( .A(start_reg[394]), .B(init), .Z(start_in[394]) );
  AND U12495 ( .A(start_reg[393]), .B(init), .Z(start_in[393]) );
  AND U12496 ( .A(start_reg[392]), .B(init), .Z(start_in[392]) );
  AND U12497 ( .A(start_reg[391]), .B(init), .Z(start_in[391]) );
  AND U12498 ( .A(start_reg[390]), .B(init), .Z(start_in[390]) );
  AND U12499 ( .A(start_reg[38]), .B(init), .Z(start_in[38]) );
  AND U12500 ( .A(start_reg[389]), .B(init), .Z(start_in[389]) );
  AND U12501 ( .A(start_reg[388]), .B(init), .Z(start_in[388]) );
  AND U12502 ( .A(start_reg[387]), .B(init), .Z(start_in[387]) );
  AND U12503 ( .A(start_reg[386]), .B(init), .Z(start_in[386]) );
  AND U12504 ( .A(start_reg[385]), .B(init), .Z(start_in[385]) );
  AND U12505 ( .A(start_reg[384]), .B(init), .Z(start_in[384]) );
  AND U12506 ( .A(start_reg[383]), .B(init), .Z(start_in[383]) );
  AND U12507 ( .A(start_reg[382]), .B(init), .Z(start_in[382]) );
  AND U12508 ( .A(start_reg[381]), .B(init), .Z(start_in[381]) );
  AND U12509 ( .A(start_reg[380]), .B(init), .Z(start_in[380]) );
  AND U12510 ( .A(start_reg[37]), .B(init), .Z(start_in[37]) );
  AND U12511 ( .A(start_reg[379]), .B(init), .Z(start_in[379]) );
  AND U12512 ( .A(start_reg[378]), .B(init), .Z(start_in[378]) );
  AND U12513 ( .A(start_reg[377]), .B(init), .Z(start_in[377]) );
  AND U12514 ( .A(start_reg[376]), .B(init), .Z(start_in[376]) );
  AND U12515 ( .A(start_reg[375]), .B(init), .Z(start_in[375]) );
  AND U12516 ( .A(start_reg[374]), .B(init), .Z(start_in[374]) );
  AND U12517 ( .A(start_reg[373]), .B(init), .Z(start_in[373]) );
  AND U12518 ( .A(start_reg[372]), .B(init), .Z(start_in[372]) );
  AND U12519 ( .A(start_reg[371]), .B(init), .Z(start_in[371]) );
  AND U12520 ( .A(start_reg[370]), .B(init), .Z(start_in[370]) );
  AND U12521 ( .A(start_reg[36]), .B(init), .Z(start_in[36]) );
  AND U12522 ( .A(start_reg[369]), .B(init), .Z(start_in[369]) );
  AND U12523 ( .A(start_reg[368]), .B(init), .Z(start_in[368]) );
  AND U12524 ( .A(start_reg[367]), .B(init), .Z(start_in[367]) );
  AND U12525 ( .A(start_reg[366]), .B(init), .Z(start_in[366]) );
  AND U12526 ( .A(start_reg[365]), .B(init), .Z(start_in[365]) );
  AND U12527 ( .A(start_reg[364]), .B(init), .Z(start_in[364]) );
  AND U12528 ( .A(start_reg[363]), .B(init), .Z(start_in[363]) );
  AND U12529 ( .A(start_reg[362]), .B(init), .Z(start_in[362]) );
  AND U12530 ( .A(start_reg[361]), .B(init), .Z(start_in[361]) );
  AND U12531 ( .A(start_reg[360]), .B(init), .Z(start_in[360]) );
  AND U12532 ( .A(start_reg[35]), .B(init), .Z(start_in[35]) );
  AND U12533 ( .A(start_reg[359]), .B(init), .Z(start_in[359]) );
  AND U12534 ( .A(start_reg[358]), .B(init), .Z(start_in[358]) );
  AND U12535 ( .A(start_reg[357]), .B(init), .Z(start_in[357]) );
  AND U12536 ( .A(start_reg[356]), .B(init), .Z(start_in[356]) );
  AND U12537 ( .A(start_reg[355]), .B(init), .Z(start_in[355]) );
  AND U12538 ( .A(start_reg[354]), .B(init), .Z(start_in[354]) );
  AND U12539 ( .A(start_reg[353]), .B(init), .Z(start_in[353]) );
  AND U12540 ( .A(start_reg[352]), .B(init), .Z(start_in[352]) );
  AND U12541 ( .A(start_reg[351]), .B(init), .Z(start_in[351]) );
  AND U12542 ( .A(start_reg[350]), .B(init), .Z(start_in[350]) );
  AND U12543 ( .A(start_reg[34]), .B(init), .Z(start_in[34]) );
  AND U12544 ( .A(start_reg[349]), .B(init), .Z(start_in[349]) );
  AND U12545 ( .A(start_reg[348]), .B(init), .Z(start_in[348]) );
  AND U12546 ( .A(start_reg[347]), .B(init), .Z(start_in[347]) );
  AND U12547 ( .A(start_reg[346]), .B(init), .Z(start_in[346]) );
  AND U12548 ( .A(start_reg[345]), .B(init), .Z(start_in[345]) );
  AND U12549 ( .A(start_reg[344]), .B(init), .Z(start_in[344]) );
  AND U12550 ( .A(start_reg[343]), .B(init), .Z(start_in[343]) );
  AND U12551 ( .A(start_reg[342]), .B(init), .Z(start_in[342]) );
  AND U12552 ( .A(start_reg[341]), .B(init), .Z(start_in[341]) );
  AND U12553 ( .A(start_reg[340]), .B(init), .Z(start_in[340]) );
  AND U12554 ( .A(start_reg[33]), .B(init), .Z(start_in[33]) );
  AND U12555 ( .A(start_reg[339]), .B(init), .Z(start_in[339]) );
  AND U12556 ( .A(start_reg[338]), .B(init), .Z(start_in[338]) );
  AND U12557 ( .A(start_reg[337]), .B(init), .Z(start_in[337]) );
  AND U12558 ( .A(start_reg[336]), .B(init), .Z(start_in[336]) );
  AND U12559 ( .A(start_reg[335]), .B(init), .Z(start_in[335]) );
  AND U12560 ( .A(start_reg[334]), .B(init), .Z(start_in[334]) );
  AND U12561 ( .A(start_reg[333]), .B(init), .Z(start_in[333]) );
  AND U12562 ( .A(start_reg[332]), .B(init), .Z(start_in[332]) );
  AND U12563 ( .A(start_reg[331]), .B(init), .Z(start_in[331]) );
  AND U12564 ( .A(start_reg[330]), .B(init), .Z(start_in[330]) );
  AND U12565 ( .A(start_reg[32]), .B(init), .Z(start_in[32]) );
  AND U12566 ( .A(start_reg[329]), .B(init), .Z(start_in[329]) );
  AND U12567 ( .A(start_reg[328]), .B(init), .Z(start_in[328]) );
  AND U12568 ( .A(start_reg[327]), .B(init), .Z(start_in[327]) );
  AND U12569 ( .A(start_reg[326]), .B(init), .Z(start_in[326]) );
  AND U12570 ( .A(start_reg[325]), .B(init), .Z(start_in[325]) );
  AND U12571 ( .A(start_reg[324]), .B(init), .Z(start_in[324]) );
  AND U12572 ( .A(start_reg[323]), .B(init), .Z(start_in[323]) );
  AND U12573 ( .A(start_reg[322]), .B(init), .Z(start_in[322]) );
  AND U12574 ( .A(start_reg[321]), .B(init), .Z(start_in[321]) );
  AND U12575 ( .A(start_reg[320]), .B(init), .Z(start_in[320]) );
  AND U12576 ( .A(start_reg[31]), .B(init), .Z(start_in[31]) );
  AND U12577 ( .A(start_reg[319]), .B(init), .Z(start_in[319]) );
  AND U12578 ( .A(start_reg[318]), .B(init), .Z(start_in[318]) );
  AND U12579 ( .A(start_reg[317]), .B(init), .Z(start_in[317]) );
  AND U12580 ( .A(start_reg[316]), .B(init), .Z(start_in[316]) );
  AND U12581 ( .A(start_reg[315]), .B(init), .Z(start_in[315]) );
  AND U12582 ( .A(start_reg[314]), .B(init), .Z(start_in[314]) );
  AND U12583 ( .A(start_reg[313]), .B(init), .Z(start_in[313]) );
  AND U12584 ( .A(start_reg[312]), .B(init), .Z(start_in[312]) );
  AND U12585 ( .A(start_reg[311]), .B(init), .Z(start_in[311]) );
  AND U12586 ( .A(start_reg[310]), .B(init), .Z(start_in[310]) );
  AND U12587 ( .A(start_reg[30]), .B(init), .Z(start_in[30]) );
  AND U12588 ( .A(start_reg[309]), .B(init), .Z(start_in[309]) );
  AND U12589 ( .A(start_reg[308]), .B(init), .Z(start_in[308]) );
  AND U12590 ( .A(start_reg[307]), .B(init), .Z(start_in[307]) );
  AND U12591 ( .A(start_reg[306]), .B(init), .Z(start_in[306]) );
  AND U12592 ( .A(start_reg[305]), .B(init), .Z(start_in[305]) );
  AND U12593 ( .A(start_reg[304]), .B(init), .Z(start_in[304]) );
  AND U12594 ( .A(start_reg[303]), .B(init), .Z(start_in[303]) );
  AND U12595 ( .A(start_reg[302]), .B(init), .Z(start_in[302]) );
  AND U12596 ( .A(start_reg[301]), .B(init), .Z(start_in[301]) );
  AND U12597 ( .A(start_reg[300]), .B(init), .Z(start_in[300]) );
  AND U12598 ( .A(start_reg[2]), .B(init), .Z(start_in[2]) );
  AND U12599 ( .A(start_reg[29]), .B(init), .Z(start_in[29]) );
  AND U12600 ( .A(start_reg[299]), .B(init), .Z(start_in[299]) );
  AND U12601 ( .A(start_reg[298]), .B(init), .Z(start_in[298]) );
  AND U12602 ( .A(start_reg[297]), .B(init), .Z(start_in[297]) );
  AND U12603 ( .A(start_reg[296]), .B(init), .Z(start_in[296]) );
  AND U12604 ( .A(start_reg[295]), .B(init), .Z(start_in[295]) );
  AND U12605 ( .A(start_reg[294]), .B(init), .Z(start_in[294]) );
  AND U12606 ( .A(start_reg[293]), .B(init), .Z(start_in[293]) );
  AND U12607 ( .A(start_reg[292]), .B(init), .Z(start_in[292]) );
  AND U12608 ( .A(start_reg[291]), .B(init), .Z(start_in[291]) );
  AND U12609 ( .A(start_reg[290]), .B(init), .Z(start_in[290]) );
  AND U12610 ( .A(start_reg[28]), .B(init), .Z(start_in[28]) );
  AND U12611 ( .A(start_reg[289]), .B(init), .Z(start_in[289]) );
  AND U12612 ( .A(start_reg[288]), .B(init), .Z(start_in[288]) );
  AND U12613 ( .A(start_reg[287]), .B(init), .Z(start_in[287]) );
  AND U12614 ( .A(start_reg[286]), .B(init), .Z(start_in[286]) );
  AND U12615 ( .A(start_reg[285]), .B(init), .Z(start_in[285]) );
  AND U12616 ( .A(start_reg[284]), .B(init), .Z(start_in[284]) );
  AND U12617 ( .A(start_reg[283]), .B(init), .Z(start_in[283]) );
  AND U12618 ( .A(start_reg[282]), .B(init), .Z(start_in[282]) );
  AND U12619 ( .A(start_reg[281]), .B(init), .Z(start_in[281]) );
  AND U12620 ( .A(start_reg[280]), .B(init), .Z(start_in[280]) );
  AND U12621 ( .A(start_reg[27]), .B(init), .Z(start_in[27]) );
  AND U12622 ( .A(start_reg[279]), .B(init), .Z(start_in[279]) );
  AND U12623 ( .A(start_reg[278]), .B(init), .Z(start_in[278]) );
  AND U12624 ( .A(start_reg[277]), .B(init), .Z(start_in[277]) );
  AND U12625 ( .A(start_reg[276]), .B(init), .Z(start_in[276]) );
  AND U12626 ( .A(start_reg[275]), .B(init), .Z(start_in[275]) );
  AND U12627 ( .A(start_reg[274]), .B(init), .Z(start_in[274]) );
  AND U12628 ( .A(start_reg[273]), .B(init), .Z(start_in[273]) );
  AND U12629 ( .A(start_reg[272]), .B(init), .Z(start_in[272]) );
  AND U12630 ( .A(start_reg[271]), .B(init), .Z(start_in[271]) );
  AND U12631 ( .A(start_reg[270]), .B(init), .Z(start_in[270]) );
  AND U12632 ( .A(start_reg[26]), .B(init), .Z(start_in[26]) );
  AND U12633 ( .A(start_reg[269]), .B(init), .Z(start_in[269]) );
  AND U12634 ( .A(start_reg[268]), .B(init), .Z(start_in[268]) );
  AND U12635 ( .A(start_reg[267]), .B(init), .Z(start_in[267]) );
  AND U12636 ( .A(start_reg[266]), .B(init), .Z(start_in[266]) );
  AND U12637 ( .A(start_reg[265]), .B(init), .Z(start_in[265]) );
  AND U12638 ( .A(start_reg[264]), .B(init), .Z(start_in[264]) );
  AND U12639 ( .A(start_reg[263]), .B(init), .Z(start_in[263]) );
  AND U12640 ( .A(start_reg[262]), .B(init), .Z(start_in[262]) );
  AND U12641 ( .A(start_reg[261]), .B(init), .Z(start_in[261]) );
  AND U12642 ( .A(start_reg[260]), .B(init), .Z(start_in[260]) );
  AND U12643 ( .A(start_reg[25]), .B(init), .Z(start_in[25]) );
  AND U12644 ( .A(start_reg[259]), .B(init), .Z(start_in[259]) );
  AND U12645 ( .A(start_reg[258]), .B(init), .Z(start_in[258]) );
  AND U12646 ( .A(start_reg[257]), .B(init), .Z(start_in[257]) );
  AND U12647 ( .A(start_reg[256]), .B(init), .Z(start_in[256]) );
  AND U12648 ( .A(start_reg[255]), .B(init), .Z(start_in[255]) );
  AND U12649 ( .A(start_reg[254]), .B(init), .Z(start_in[254]) );
  AND U12650 ( .A(start_reg[253]), .B(init), .Z(start_in[253]) );
  AND U12651 ( .A(start_reg[252]), .B(init), .Z(start_in[252]) );
  AND U12652 ( .A(start_reg[251]), .B(init), .Z(start_in[251]) );
  AND U12653 ( .A(start_reg[250]), .B(init), .Z(start_in[250]) );
  AND U12654 ( .A(start_reg[24]), .B(init), .Z(start_in[24]) );
  AND U12655 ( .A(start_reg[249]), .B(init), .Z(start_in[249]) );
  AND U12656 ( .A(start_reg[248]), .B(init), .Z(start_in[248]) );
  AND U12657 ( .A(start_reg[247]), .B(init), .Z(start_in[247]) );
  AND U12658 ( .A(start_reg[246]), .B(init), .Z(start_in[246]) );
  AND U12659 ( .A(start_reg[245]), .B(init), .Z(start_in[245]) );
  AND U12660 ( .A(start_reg[244]), .B(init), .Z(start_in[244]) );
  AND U12661 ( .A(start_reg[243]), .B(init), .Z(start_in[243]) );
  AND U12662 ( .A(start_reg[242]), .B(init), .Z(start_in[242]) );
  AND U12663 ( .A(start_reg[241]), .B(init), .Z(start_in[241]) );
  AND U12664 ( .A(start_reg[240]), .B(init), .Z(start_in[240]) );
  AND U12665 ( .A(start_reg[23]), .B(init), .Z(start_in[23]) );
  AND U12666 ( .A(start_reg[239]), .B(init), .Z(start_in[239]) );
  AND U12667 ( .A(start_reg[238]), .B(init), .Z(start_in[238]) );
  AND U12668 ( .A(start_reg[237]), .B(init), .Z(start_in[237]) );
  AND U12669 ( .A(start_reg[236]), .B(init), .Z(start_in[236]) );
  AND U12670 ( .A(start_reg[235]), .B(init), .Z(start_in[235]) );
  AND U12671 ( .A(start_reg[234]), .B(init), .Z(start_in[234]) );
  AND U12672 ( .A(start_reg[233]), .B(init), .Z(start_in[233]) );
  AND U12673 ( .A(start_reg[232]), .B(init), .Z(start_in[232]) );
  AND U12674 ( .A(start_reg[231]), .B(init), .Z(start_in[231]) );
  AND U12675 ( .A(start_reg[230]), .B(init), .Z(start_in[230]) );
  AND U12676 ( .A(start_reg[22]), .B(init), .Z(start_in[22]) );
  AND U12677 ( .A(start_reg[229]), .B(init), .Z(start_in[229]) );
  AND U12678 ( .A(start_reg[228]), .B(init), .Z(start_in[228]) );
  AND U12679 ( .A(start_reg[227]), .B(init), .Z(start_in[227]) );
  AND U12680 ( .A(start_reg[226]), .B(init), .Z(start_in[226]) );
  AND U12681 ( .A(start_reg[225]), .B(init), .Z(start_in[225]) );
  AND U12682 ( .A(start_reg[224]), .B(init), .Z(start_in[224]) );
  AND U12683 ( .A(start_reg[223]), .B(init), .Z(start_in[223]) );
  AND U12684 ( .A(start_reg[222]), .B(init), .Z(start_in[222]) );
  AND U12685 ( .A(start_reg[221]), .B(init), .Z(start_in[221]) );
  AND U12686 ( .A(start_reg[220]), .B(init), .Z(start_in[220]) );
  AND U12687 ( .A(start_reg[21]), .B(init), .Z(start_in[21]) );
  AND U12688 ( .A(start_reg[219]), .B(init), .Z(start_in[219]) );
  AND U12689 ( .A(start_reg[218]), .B(init), .Z(start_in[218]) );
  AND U12690 ( .A(start_reg[217]), .B(init), .Z(start_in[217]) );
  AND U12691 ( .A(start_reg[216]), .B(init), .Z(start_in[216]) );
  AND U12692 ( .A(start_reg[215]), .B(init), .Z(start_in[215]) );
  AND U12693 ( .A(start_reg[214]), .B(init), .Z(start_in[214]) );
  AND U12694 ( .A(start_reg[213]), .B(init), .Z(start_in[213]) );
  AND U12695 ( .A(start_reg[212]), .B(init), .Z(start_in[212]) );
  AND U12696 ( .A(start_reg[211]), .B(init), .Z(start_in[211]) );
  AND U12697 ( .A(start_reg[210]), .B(init), .Z(start_in[210]) );
  AND U12698 ( .A(start_reg[20]), .B(init), .Z(start_in[20]) );
  AND U12699 ( .A(start_reg[209]), .B(init), .Z(start_in[209]) );
  AND U12700 ( .A(start_reg[208]), .B(init), .Z(start_in[208]) );
  AND U12701 ( .A(start_reg[207]), .B(init), .Z(start_in[207]) );
  AND U12702 ( .A(start_reg[206]), .B(init), .Z(start_in[206]) );
  AND U12703 ( .A(start_reg[205]), .B(init), .Z(start_in[205]) );
  AND U12704 ( .A(start_reg[204]), .B(init), .Z(start_in[204]) );
  AND U12705 ( .A(start_reg[203]), .B(init), .Z(start_in[203]) );
  AND U12706 ( .A(start_reg[202]), .B(init), .Z(start_in[202]) );
  AND U12707 ( .A(start_reg[201]), .B(init), .Z(start_in[201]) );
  AND U12708 ( .A(start_reg[200]), .B(init), .Z(start_in[200]) );
  AND U12709 ( .A(start_reg[1]), .B(init), .Z(start_in[1]) );
  AND U12710 ( .A(start_reg[19]), .B(init), .Z(start_in[19]) );
  AND U12711 ( .A(start_reg[199]), .B(init), .Z(start_in[199]) );
  AND U12712 ( .A(start_reg[198]), .B(init), .Z(start_in[198]) );
  AND U12713 ( .A(start_reg[197]), .B(init), .Z(start_in[197]) );
  AND U12714 ( .A(start_reg[196]), .B(init), .Z(start_in[196]) );
  AND U12715 ( .A(start_reg[195]), .B(init), .Z(start_in[195]) );
  AND U12716 ( .A(start_reg[194]), .B(init), .Z(start_in[194]) );
  AND U12717 ( .A(start_reg[193]), .B(init), .Z(start_in[193]) );
  AND U12718 ( .A(start_reg[192]), .B(init), .Z(start_in[192]) );
  AND U12719 ( .A(start_reg[191]), .B(init), .Z(start_in[191]) );
  AND U12720 ( .A(start_reg[190]), .B(init), .Z(start_in[190]) );
  AND U12721 ( .A(start_reg[18]), .B(init), .Z(start_in[18]) );
  AND U12722 ( .A(start_reg[189]), .B(init), .Z(start_in[189]) );
  AND U12723 ( .A(start_reg[188]), .B(init), .Z(start_in[188]) );
  AND U12724 ( .A(start_reg[187]), .B(init), .Z(start_in[187]) );
  AND U12725 ( .A(start_reg[186]), .B(init), .Z(start_in[186]) );
  AND U12726 ( .A(start_reg[185]), .B(init), .Z(start_in[185]) );
  AND U12727 ( .A(start_reg[184]), .B(init), .Z(start_in[184]) );
  AND U12728 ( .A(start_reg[183]), .B(init), .Z(start_in[183]) );
  AND U12729 ( .A(start_reg[182]), .B(init), .Z(start_in[182]) );
  AND U12730 ( .A(start_reg[181]), .B(init), .Z(start_in[181]) );
  AND U12731 ( .A(start_reg[180]), .B(init), .Z(start_in[180]) );
  AND U12732 ( .A(start_reg[17]), .B(init), .Z(start_in[17]) );
  AND U12733 ( .A(start_reg[179]), .B(init), .Z(start_in[179]) );
  AND U12734 ( .A(start_reg[178]), .B(init), .Z(start_in[178]) );
  AND U12735 ( .A(start_reg[177]), .B(init), .Z(start_in[177]) );
  AND U12736 ( .A(start_reg[176]), .B(init), .Z(start_in[176]) );
  AND U12737 ( .A(start_reg[175]), .B(init), .Z(start_in[175]) );
  AND U12738 ( .A(start_reg[174]), .B(init), .Z(start_in[174]) );
  AND U12739 ( .A(start_reg[173]), .B(init), .Z(start_in[173]) );
  AND U12740 ( .A(start_reg[172]), .B(init), .Z(start_in[172]) );
  AND U12741 ( .A(start_reg[171]), .B(init), .Z(start_in[171]) );
  AND U12742 ( .A(start_reg[170]), .B(init), .Z(start_in[170]) );
  AND U12743 ( .A(start_reg[16]), .B(init), .Z(start_in[16]) );
  AND U12744 ( .A(start_reg[169]), .B(init), .Z(start_in[169]) );
  AND U12745 ( .A(start_reg[168]), .B(init), .Z(start_in[168]) );
  AND U12746 ( .A(start_reg[167]), .B(init), .Z(start_in[167]) );
  AND U12747 ( .A(start_reg[166]), .B(init), .Z(start_in[166]) );
  AND U12748 ( .A(start_reg[165]), .B(init), .Z(start_in[165]) );
  AND U12749 ( .A(start_reg[164]), .B(init), .Z(start_in[164]) );
  AND U12750 ( .A(start_reg[163]), .B(init), .Z(start_in[163]) );
  AND U12751 ( .A(start_reg[162]), .B(init), .Z(start_in[162]) );
  AND U12752 ( .A(start_reg[161]), .B(init), .Z(start_in[161]) );
  AND U12753 ( .A(start_reg[160]), .B(init), .Z(start_in[160]) );
  AND U12754 ( .A(start_reg[15]), .B(init), .Z(start_in[15]) );
  AND U12755 ( .A(start_reg[159]), .B(init), .Z(start_in[159]) );
  AND U12756 ( .A(start_reg[158]), .B(init), .Z(start_in[158]) );
  AND U12757 ( .A(start_reg[157]), .B(init), .Z(start_in[157]) );
  AND U12758 ( .A(start_reg[156]), .B(init), .Z(start_in[156]) );
  AND U12759 ( .A(start_reg[155]), .B(init), .Z(start_in[155]) );
  AND U12760 ( .A(start_reg[154]), .B(init), .Z(start_in[154]) );
  AND U12761 ( .A(start_reg[153]), .B(init), .Z(start_in[153]) );
  AND U12762 ( .A(start_reg[152]), .B(init), .Z(start_in[152]) );
  AND U12763 ( .A(start_reg[151]), .B(init), .Z(start_in[151]) );
  AND U12764 ( .A(start_reg[150]), .B(init), .Z(start_in[150]) );
  AND U12765 ( .A(start_reg[14]), .B(init), .Z(start_in[14]) );
  AND U12766 ( .A(start_reg[149]), .B(init), .Z(start_in[149]) );
  AND U12767 ( .A(start_reg[148]), .B(init), .Z(start_in[148]) );
  AND U12768 ( .A(start_reg[147]), .B(init), .Z(start_in[147]) );
  AND U12769 ( .A(start_reg[146]), .B(init), .Z(start_in[146]) );
  AND U12770 ( .A(start_reg[145]), .B(init), .Z(start_in[145]) );
  AND U12771 ( .A(start_reg[144]), .B(init), .Z(start_in[144]) );
  AND U12772 ( .A(start_reg[143]), .B(init), .Z(start_in[143]) );
  AND U12773 ( .A(start_reg[142]), .B(init), .Z(start_in[142]) );
  AND U12774 ( .A(start_reg[141]), .B(init), .Z(start_in[141]) );
  AND U12775 ( .A(start_reg[140]), .B(init), .Z(start_in[140]) );
  AND U12776 ( .A(start_reg[13]), .B(init), .Z(start_in[13]) );
  AND U12777 ( .A(start_reg[139]), .B(init), .Z(start_in[139]) );
  AND U12778 ( .A(start_reg[138]), .B(init), .Z(start_in[138]) );
  AND U12779 ( .A(start_reg[137]), .B(init), .Z(start_in[137]) );
  AND U12780 ( .A(start_reg[136]), .B(init), .Z(start_in[136]) );
  AND U12781 ( .A(start_reg[135]), .B(init), .Z(start_in[135]) );
  AND U12782 ( .A(start_reg[134]), .B(init), .Z(start_in[134]) );
  AND U12783 ( .A(start_reg[133]), .B(init), .Z(start_in[133]) );
  AND U12784 ( .A(start_reg[132]), .B(init), .Z(start_in[132]) );
  AND U12785 ( .A(start_reg[131]), .B(init), .Z(start_in[131]) );
  AND U12786 ( .A(start_reg[130]), .B(init), .Z(start_in[130]) );
  AND U12787 ( .A(start_reg[12]), .B(init), .Z(start_in[12]) );
  AND U12788 ( .A(start_reg[129]), .B(init), .Z(start_in[129]) );
  AND U12789 ( .A(start_reg[128]), .B(init), .Z(start_in[128]) );
  AND U12790 ( .A(start_reg[127]), .B(init), .Z(start_in[127]) );
  AND U12791 ( .A(start_reg[126]), .B(init), .Z(start_in[126]) );
  AND U12792 ( .A(start_reg[125]), .B(init), .Z(start_in[125]) );
  AND U12793 ( .A(start_reg[124]), .B(init), .Z(start_in[124]) );
  AND U12794 ( .A(start_reg[123]), .B(init), .Z(start_in[123]) );
  AND U12795 ( .A(start_reg[122]), .B(init), .Z(start_in[122]) );
  AND U12796 ( .A(start_reg[121]), .B(init), .Z(start_in[121]) );
  AND U12797 ( .A(start_reg[120]), .B(init), .Z(start_in[120]) );
  AND U12798 ( .A(start_reg[11]), .B(init), .Z(start_in[11]) );
  AND U12799 ( .A(start_reg[119]), .B(init), .Z(start_in[119]) );
  AND U12800 ( .A(start_reg[118]), .B(init), .Z(start_in[118]) );
  AND U12801 ( .A(start_reg[117]), .B(init), .Z(start_in[117]) );
  AND U12802 ( .A(start_reg[116]), .B(init), .Z(start_in[116]) );
  AND U12803 ( .A(start_reg[115]), .B(init), .Z(start_in[115]) );
  AND U12804 ( .A(start_reg[114]), .B(init), .Z(start_in[114]) );
  AND U12805 ( .A(start_reg[113]), .B(init), .Z(start_in[113]) );
  AND U12806 ( .A(start_reg[112]), .B(init), .Z(start_in[112]) );
  AND U12807 ( .A(start_reg[111]), .B(init), .Z(start_in[111]) );
  AND U12808 ( .A(start_reg[110]), .B(init), .Z(start_in[110]) );
  AND U12809 ( .A(start_reg[10]), .B(init), .Z(start_in[10]) );
  AND U12810 ( .A(start_reg[109]), .B(init), .Z(start_in[109]) );
  AND U12811 ( .A(start_reg[108]), .B(init), .Z(start_in[108]) );
  AND U12812 ( .A(start_reg[107]), .B(init), .Z(start_in[107]) );
  AND U12813 ( .A(start_reg[106]), .B(init), .Z(start_in[106]) );
  AND U12814 ( .A(start_reg[105]), .B(init), .Z(start_in[105]) );
  AND U12815 ( .A(start_reg[104]), .B(init), .Z(start_in[104]) );
  AND U12816 ( .A(start_reg[103]), .B(init), .Z(start_in[103]) );
  AND U12817 ( .A(start_reg[102]), .B(init), .Z(start_in[102]) );
  AND U12818 ( .A(start_reg[101]), .B(init), .Z(start_in[101]) );
  AND U12819 ( .A(start_reg[100]), .B(init), .Z(start_in[100]) );
  NANDN U12820 ( .A(start_reg[0]), .B(init), .Z(start_in[0]) );
  NAND U12821 ( .A(n9750), .B(n9751), .Z(n7699) );
  NAND U12822 ( .A(n7703), .B(start_reg[511]), .Z(n9751) );
  IV U12823 ( .A(n7702), .Z(n7703) );
  NANDN U12824 ( .A(n14372), .B(mul_pow), .Z(n9750) );
  NAND U12825 ( .A(n9752), .B(n9753), .Z(n7698) );
  NANDN U12826 ( .A(n9754), .B(ereg[0]), .Z(n9753) );
  NANDN U12827 ( .A(init), .B(e[0]), .Z(n9752) );
  NAND U12828 ( .A(n9755), .B(n9756), .Z(n7697) );
  NANDN U12829 ( .A(init), .B(e[1]), .Z(n9756) );
  AND U12830 ( .A(n9757), .B(n9758), .Z(n9755) );
  NAND U12831 ( .A(n9759), .B(ereg[0]), .Z(n9758) );
  NANDN U12832 ( .A(n9754), .B(ereg[1]), .Z(n9757) );
  NAND U12833 ( .A(n9760), .B(n9761), .Z(n7696) );
  NANDN U12834 ( .A(init), .B(e[2]), .Z(n9761) );
  AND U12835 ( .A(n9762), .B(n9763), .Z(n9760) );
  NAND U12836 ( .A(ereg[1]), .B(n9759), .Z(n9763) );
  NANDN U12837 ( .A(n9754), .B(ereg[2]), .Z(n9762) );
  NAND U12838 ( .A(n9764), .B(n9765), .Z(n7695) );
  NANDN U12839 ( .A(init), .B(e[3]), .Z(n9765) );
  AND U12840 ( .A(n9766), .B(n9767), .Z(n9764) );
  NAND U12841 ( .A(ereg[2]), .B(n9759), .Z(n9767) );
  NANDN U12842 ( .A(n9754), .B(ereg[3]), .Z(n9766) );
  NAND U12843 ( .A(n9768), .B(n9769), .Z(n7694) );
  NANDN U12844 ( .A(init), .B(e[4]), .Z(n9769) );
  AND U12845 ( .A(n9770), .B(n9771), .Z(n9768) );
  NAND U12846 ( .A(ereg[3]), .B(n9759), .Z(n9771) );
  NANDN U12847 ( .A(n9754), .B(ereg[4]), .Z(n9770) );
  NAND U12848 ( .A(n9772), .B(n9773), .Z(n7693) );
  NANDN U12849 ( .A(init), .B(e[5]), .Z(n9773) );
  AND U12850 ( .A(n9774), .B(n9775), .Z(n9772) );
  NAND U12851 ( .A(ereg[4]), .B(n9759), .Z(n9775) );
  NANDN U12852 ( .A(n9754), .B(ereg[5]), .Z(n9774) );
  NAND U12853 ( .A(n9776), .B(n9777), .Z(n7692) );
  NANDN U12854 ( .A(init), .B(e[6]), .Z(n9777) );
  AND U12855 ( .A(n9778), .B(n9779), .Z(n9776) );
  NAND U12856 ( .A(ereg[5]), .B(n9759), .Z(n9779) );
  NANDN U12857 ( .A(n9754), .B(ereg[6]), .Z(n9778) );
  NAND U12858 ( .A(n9780), .B(n9781), .Z(n7691) );
  NANDN U12859 ( .A(init), .B(e[7]), .Z(n9781) );
  AND U12860 ( .A(n9782), .B(n9783), .Z(n9780) );
  NAND U12861 ( .A(ereg[6]), .B(n9759), .Z(n9783) );
  NANDN U12862 ( .A(n9754), .B(ereg[7]), .Z(n9782) );
  NAND U12863 ( .A(n9784), .B(n9785), .Z(n7690) );
  NANDN U12864 ( .A(init), .B(e[8]), .Z(n9785) );
  AND U12865 ( .A(n9786), .B(n9787), .Z(n9784) );
  NAND U12866 ( .A(ereg[7]), .B(n9759), .Z(n9787) );
  NANDN U12867 ( .A(n9754), .B(ereg[8]), .Z(n9786) );
  NAND U12868 ( .A(n9788), .B(n9789), .Z(n7689) );
  NANDN U12869 ( .A(init), .B(e[9]), .Z(n9789) );
  AND U12870 ( .A(n9790), .B(n9791), .Z(n9788) );
  NAND U12871 ( .A(ereg[8]), .B(n9759), .Z(n9791) );
  NANDN U12872 ( .A(n9754), .B(ereg[9]), .Z(n9790) );
  NAND U12873 ( .A(n9792), .B(n9793), .Z(n7688) );
  NANDN U12874 ( .A(init), .B(e[10]), .Z(n9793) );
  AND U12875 ( .A(n9794), .B(n9795), .Z(n9792) );
  NAND U12876 ( .A(ereg[9]), .B(n9759), .Z(n9795) );
  NANDN U12877 ( .A(n9754), .B(ereg[10]), .Z(n9794) );
  NAND U12878 ( .A(n9796), .B(n9797), .Z(n7687) );
  NANDN U12879 ( .A(init), .B(e[11]), .Z(n9797) );
  AND U12880 ( .A(n9798), .B(n9799), .Z(n9796) );
  NAND U12881 ( .A(ereg[10]), .B(n9759), .Z(n9799) );
  NANDN U12882 ( .A(n9754), .B(ereg[11]), .Z(n9798) );
  NAND U12883 ( .A(n9800), .B(n9801), .Z(n7686) );
  NANDN U12884 ( .A(init), .B(e[12]), .Z(n9801) );
  AND U12885 ( .A(n9802), .B(n9803), .Z(n9800) );
  NAND U12886 ( .A(ereg[11]), .B(n9759), .Z(n9803) );
  NANDN U12887 ( .A(n9754), .B(ereg[12]), .Z(n9802) );
  NAND U12888 ( .A(n9804), .B(n9805), .Z(n7685) );
  NANDN U12889 ( .A(init), .B(e[13]), .Z(n9805) );
  AND U12890 ( .A(n9806), .B(n9807), .Z(n9804) );
  NAND U12891 ( .A(ereg[12]), .B(n9759), .Z(n9807) );
  NANDN U12892 ( .A(n9754), .B(ereg[13]), .Z(n9806) );
  NAND U12893 ( .A(n9808), .B(n9809), .Z(n7684) );
  NANDN U12894 ( .A(init), .B(e[14]), .Z(n9809) );
  AND U12895 ( .A(n9810), .B(n9811), .Z(n9808) );
  NAND U12896 ( .A(ereg[13]), .B(n9759), .Z(n9811) );
  NANDN U12897 ( .A(n9754), .B(ereg[14]), .Z(n9810) );
  NAND U12898 ( .A(n9812), .B(n9813), .Z(n7683) );
  NANDN U12899 ( .A(init), .B(e[15]), .Z(n9813) );
  AND U12900 ( .A(n9814), .B(n9815), .Z(n9812) );
  NAND U12901 ( .A(ereg[14]), .B(n9759), .Z(n9815) );
  NANDN U12902 ( .A(n9754), .B(ereg[15]), .Z(n9814) );
  NAND U12903 ( .A(n9816), .B(n9817), .Z(n7682) );
  NANDN U12904 ( .A(init), .B(e[16]), .Z(n9817) );
  AND U12905 ( .A(n9818), .B(n9819), .Z(n9816) );
  NAND U12906 ( .A(ereg[15]), .B(n9759), .Z(n9819) );
  NANDN U12907 ( .A(n9754), .B(ereg[16]), .Z(n9818) );
  NAND U12908 ( .A(n9820), .B(n9821), .Z(n7681) );
  NANDN U12909 ( .A(init), .B(e[17]), .Z(n9821) );
  AND U12910 ( .A(n9822), .B(n9823), .Z(n9820) );
  NAND U12911 ( .A(ereg[16]), .B(n9759), .Z(n9823) );
  NANDN U12912 ( .A(n9754), .B(ereg[17]), .Z(n9822) );
  NAND U12913 ( .A(n9824), .B(n9825), .Z(n7680) );
  NANDN U12914 ( .A(init), .B(e[18]), .Z(n9825) );
  AND U12915 ( .A(n9826), .B(n9827), .Z(n9824) );
  NAND U12916 ( .A(ereg[17]), .B(n9759), .Z(n9827) );
  NANDN U12917 ( .A(n9754), .B(ereg[18]), .Z(n9826) );
  NAND U12918 ( .A(n9828), .B(n9829), .Z(n7679) );
  NANDN U12919 ( .A(init), .B(e[19]), .Z(n9829) );
  AND U12920 ( .A(n9830), .B(n9831), .Z(n9828) );
  NAND U12921 ( .A(ereg[18]), .B(n9759), .Z(n9831) );
  NANDN U12922 ( .A(n9754), .B(ereg[19]), .Z(n9830) );
  NAND U12923 ( .A(n9832), .B(n9833), .Z(n7678) );
  NANDN U12924 ( .A(init), .B(e[20]), .Z(n9833) );
  AND U12925 ( .A(n9834), .B(n9835), .Z(n9832) );
  NAND U12926 ( .A(ereg[19]), .B(n9759), .Z(n9835) );
  NANDN U12927 ( .A(n9754), .B(ereg[20]), .Z(n9834) );
  NAND U12928 ( .A(n9836), .B(n9837), .Z(n7677) );
  NANDN U12929 ( .A(init), .B(e[21]), .Z(n9837) );
  AND U12930 ( .A(n9838), .B(n9839), .Z(n9836) );
  NAND U12931 ( .A(ereg[20]), .B(n9759), .Z(n9839) );
  NANDN U12932 ( .A(n9754), .B(ereg[21]), .Z(n9838) );
  NAND U12933 ( .A(n9840), .B(n9841), .Z(n7676) );
  NANDN U12934 ( .A(init), .B(e[22]), .Z(n9841) );
  AND U12935 ( .A(n9842), .B(n9843), .Z(n9840) );
  NAND U12936 ( .A(ereg[21]), .B(n9759), .Z(n9843) );
  NANDN U12937 ( .A(n9754), .B(ereg[22]), .Z(n9842) );
  NAND U12938 ( .A(n9844), .B(n9845), .Z(n7675) );
  NANDN U12939 ( .A(init), .B(e[23]), .Z(n9845) );
  AND U12940 ( .A(n9846), .B(n9847), .Z(n9844) );
  NAND U12941 ( .A(ereg[22]), .B(n9759), .Z(n9847) );
  NANDN U12942 ( .A(n9754), .B(ereg[23]), .Z(n9846) );
  NAND U12943 ( .A(n9848), .B(n9849), .Z(n7674) );
  NANDN U12944 ( .A(init), .B(e[24]), .Z(n9849) );
  AND U12945 ( .A(n9850), .B(n9851), .Z(n9848) );
  NAND U12946 ( .A(ereg[23]), .B(n9759), .Z(n9851) );
  NANDN U12947 ( .A(n9754), .B(ereg[24]), .Z(n9850) );
  NAND U12948 ( .A(n9852), .B(n9853), .Z(n7673) );
  NANDN U12949 ( .A(init), .B(e[25]), .Z(n9853) );
  AND U12950 ( .A(n9854), .B(n9855), .Z(n9852) );
  NAND U12951 ( .A(ereg[24]), .B(n9759), .Z(n9855) );
  NANDN U12952 ( .A(n9754), .B(ereg[25]), .Z(n9854) );
  NAND U12953 ( .A(n9856), .B(n9857), .Z(n7672) );
  NANDN U12954 ( .A(init), .B(e[26]), .Z(n9857) );
  AND U12955 ( .A(n9858), .B(n9859), .Z(n9856) );
  NAND U12956 ( .A(ereg[25]), .B(n9759), .Z(n9859) );
  NANDN U12957 ( .A(n9754), .B(ereg[26]), .Z(n9858) );
  NAND U12958 ( .A(n9860), .B(n9861), .Z(n7671) );
  NANDN U12959 ( .A(init), .B(e[27]), .Z(n9861) );
  AND U12960 ( .A(n9862), .B(n9863), .Z(n9860) );
  NAND U12961 ( .A(ereg[26]), .B(n9759), .Z(n9863) );
  NANDN U12962 ( .A(n9754), .B(ereg[27]), .Z(n9862) );
  NAND U12963 ( .A(n9864), .B(n9865), .Z(n7670) );
  NANDN U12964 ( .A(init), .B(e[28]), .Z(n9865) );
  AND U12965 ( .A(n9866), .B(n9867), .Z(n9864) );
  NAND U12966 ( .A(ereg[27]), .B(n9759), .Z(n9867) );
  NANDN U12967 ( .A(n9754), .B(ereg[28]), .Z(n9866) );
  NAND U12968 ( .A(n9868), .B(n9869), .Z(n7669) );
  NANDN U12969 ( .A(init), .B(e[29]), .Z(n9869) );
  AND U12970 ( .A(n9870), .B(n9871), .Z(n9868) );
  NAND U12971 ( .A(ereg[28]), .B(n9759), .Z(n9871) );
  NANDN U12972 ( .A(n9754), .B(ereg[29]), .Z(n9870) );
  NAND U12973 ( .A(n9872), .B(n9873), .Z(n7668) );
  NANDN U12974 ( .A(init), .B(e[30]), .Z(n9873) );
  AND U12975 ( .A(n9874), .B(n9875), .Z(n9872) );
  NAND U12976 ( .A(ereg[29]), .B(n9759), .Z(n9875) );
  NANDN U12977 ( .A(n9754), .B(ereg[30]), .Z(n9874) );
  NAND U12978 ( .A(n9876), .B(n9877), .Z(n7667) );
  NANDN U12979 ( .A(init), .B(e[31]), .Z(n9877) );
  AND U12980 ( .A(n9878), .B(n9879), .Z(n9876) );
  NAND U12981 ( .A(ereg[30]), .B(n9759), .Z(n9879) );
  NANDN U12982 ( .A(n9754), .B(ereg[31]), .Z(n9878) );
  NAND U12983 ( .A(n9880), .B(n9881), .Z(n7666) );
  NANDN U12984 ( .A(init), .B(e[32]), .Z(n9881) );
  AND U12985 ( .A(n9882), .B(n9883), .Z(n9880) );
  NAND U12986 ( .A(ereg[31]), .B(n9759), .Z(n9883) );
  NANDN U12987 ( .A(n9754), .B(ereg[32]), .Z(n9882) );
  NAND U12988 ( .A(n9884), .B(n9885), .Z(n7665) );
  NANDN U12989 ( .A(init), .B(e[33]), .Z(n9885) );
  AND U12990 ( .A(n9886), .B(n9887), .Z(n9884) );
  NAND U12991 ( .A(ereg[32]), .B(n9759), .Z(n9887) );
  NANDN U12992 ( .A(n9754), .B(ereg[33]), .Z(n9886) );
  NAND U12993 ( .A(n9888), .B(n9889), .Z(n7664) );
  NANDN U12994 ( .A(init), .B(e[34]), .Z(n9889) );
  AND U12995 ( .A(n9890), .B(n9891), .Z(n9888) );
  NAND U12996 ( .A(ereg[33]), .B(n9759), .Z(n9891) );
  NANDN U12997 ( .A(n9754), .B(ereg[34]), .Z(n9890) );
  NAND U12998 ( .A(n9892), .B(n9893), .Z(n7663) );
  NANDN U12999 ( .A(init), .B(e[35]), .Z(n9893) );
  AND U13000 ( .A(n9894), .B(n9895), .Z(n9892) );
  NAND U13001 ( .A(ereg[34]), .B(n9759), .Z(n9895) );
  NANDN U13002 ( .A(n9754), .B(ereg[35]), .Z(n9894) );
  NAND U13003 ( .A(n9896), .B(n9897), .Z(n7662) );
  NANDN U13004 ( .A(init), .B(e[36]), .Z(n9897) );
  AND U13005 ( .A(n9898), .B(n9899), .Z(n9896) );
  NAND U13006 ( .A(ereg[35]), .B(n9759), .Z(n9899) );
  NANDN U13007 ( .A(n9754), .B(ereg[36]), .Z(n9898) );
  NAND U13008 ( .A(n9900), .B(n9901), .Z(n7661) );
  NANDN U13009 ( .A(init), .B(e[37]), .Z(n9901) );
  AND U13010 ( .A(n9902), .B(n9903), .Z(n9900) );
  NAND U13011 ( .A(ereg[36]), .B(n9759), .Z(n9903) );
  NANDN U13012 ( .A(n9754), .B(ereg[37]), .Z(n9902) );
  NAND U13013 ( .A(n9904), .B(n9905), .Z(n7660) );
  NANDN U13014 ( .A(init), .B(e[38]), .Z(n9905) );
  AND U13015 ( .A(n9906), .B(n9907), .Z(n9904) );
  NAND U13016 ( .A(ereg[37]), .B(n9759), .Z(n9907) );
  NANDN U13017 ( .A(n9754), .B(ereg[38]), .Z(n9906) );
  NAND U13018 ( .A(n9908), .B(n9909), .Z(n7659) );
  NANDN U13019 ( .A(init), .B(e[39]), .Z(n9909) );
  AND U13020 ( .A(n9910), .B(n9911), .Z(n9908) );
  NAND U13021 ( .A(ereg[38]), .B(n9759), .Z(n9911) );
  NANDN U13022 ( .A(n9754), .B(ereg[39]), .Z(n9910) );
  NAND U13023 ( .A(n9912), .B(n9913), .Z(n7658) );
  NANDN U13024 ( .A(init), .B(e[40]), .Z(n9913) );
  AND U13025 ( .A(n9914), .B(n9915), .Z(n9912) );
  NAND U13026 ( .A(ereg[39]), .B(n9759), .Z(n9915) );
  NANDN U13027 ( .A(n9754), .B(ereg[40]), .Z(n9914) );
  NAND U13028 ( .A(n9916), .B(n9917), .Z(n7657) );
  NANDN U13029 ( .A(init), .B(e[41]), .Z(n9917) );
  AND U13030 ( .A(n9918), .B(n9919), .Z(n9916) );
  NAND U13031 ( .A(ereg[40]), .B(n9759), .Z(n9919) );
  NANDN U13032 ( .A(n9754), .B(ereg[41]), .Z(n9918) );
  NAND U13033 ( .A(n9920), .B(n9921), .Z(n7656) );
  NANDN U13034 ( .A(init), .B(e[42]), .Z(n9921) );
  AND U13035 ( .A(n9922), .B(n9923), .Z(n9920) );
  NAND U13036 ( .A(ereg[41]), .B(n9759), .Z(n9923) );
  NANDN U13037 ( .A(n9754), .B(ereg[42]), .Z(n9922) );
  NAND U13038 ( .A(n9924), .B(n9925), .Z(n7655) );
  NANDN U13039 ( .A(init), .B(e[43]), .Z(n9925) );
  AND U13040 ( .A(n9926), .B(n9927), .Z(n9924) );
  NAND U13041 ( .A(ereg[42]), .B(n9759), .Z(n9927) );
  NANDN U13042 ( .A(n9754), .B(ereg[43]), .Z(n9926) );
  NAND U13043 ( .A(n9928), .B(n9929), .Z(n7654) );
  NANDN U13044 ( .A(init), .B(e[44]), .Z(n9929) );
  AND U13045 ( .A(n9930), .B(n9931), .Z(n9928) );
  NAND U13046 ( .A(ereg[43]), .B(n9759), .Z(n9931) );
  NANDN U13047 ( .A(n9754), .B(ereg[44]), .Z(n9930) );
  NAND U13048 ( .A(n9932), .B(n9933), .Z(n7653) );
  NANDN U13049 ( .A(init), .B(e[45]), .Z(n9933) );
  AND U13050 ( .A(n9934), .B(n9935), .Z(n9932) );
  NAND U13051 ( .A(ereg[44]), .B(n9759), .Z(n9935) );
  NANDN U13052 ( .A(n9754), .B(ereg[45]), .Z(n9934) );
  NAND U13053 ( .A(n9936), .B(n9937), .Z(n7652) );
  NANDN U13054 ( .A(init), .B(e[46]), .Z(n9937) );
  AND U13055 ( .A(n9938), .B(n9939), .Z(n9936) );
  NAND U13056 ( .A(ereg[45]), .B(n9759), .Z(n9939) );
  NANDN U13057 ( .A(n9754), .B(ereg[46]), .Z(n9938) );
  NAND U13058 ( .A(n9940), .B(n9941), .Z(n7651) );
  NANDN U13059 ( .A(init), .B(e[47]), .Z(n9941) );
  AND U13060 ( .A(n9942), .B(n9943), .Z(n9940) );
  NAND U13061 ( .A(ereg[46]), .B(n9759), .Z(n9943) );
  NANDN U13062 ( .A(n9754), .B(ereg[47]), .Z(n9942) );
  NAND U13063 ( .A(n9944), .B(n9945), .Z(n7650) );
  NANDN U13064 ( .A(init), .B(e[48]), .Z(n9945) );
  AND U13065 ( .A(n9946), .B(n9947), .Z(n9944) );
  NAND U13066 ( .A(ereg[47]), .B(n9759), .Z(n9947) );
  NANDN U13067 ( .A(n9754), .B(ereg[48]), .Z(n9946) );
  NAND U13068 ( .A(n9948), .B(n9949), .Z(n7649) );
  NANDN U13069 ( .A(init), .B(e[49]), .Z(n9949) );
  AND U13070 ( .A(n9950), .B(n9951), .Z(n9948) );
  NAND U13071 ( .A(ereg[48]), .B(n9759), .Z(n9951) );
  NANDN U13072 ( .A(n9754), .B(ereg[49]), .Z(n9950) );
  NAND U13073 ( .A(n9952), .B(n9953), .Z(n7648) );
  NANDN U13074 ( .A(init), .B(e[50]), .Z(n9953) );
  AND U13075 ( .A(n9954), .B(n9955), .Z(n9952) );
  NAND U13076 ( .A(ereg[49]), .B(n9759), .Z(n9955) );
  NANDN U13077 ( .A(n9754), .B(ereg[50]), .Z(n9954) );
  NAND U13078 ( .A(n9956), .B(n9957), .Z(n7647) );
  NANDN U13079 ( .A(init), .B(e[51]), .Z(n9957) );
  AND U13080 ( .A(n9958), .B(n9959), .Z(n9956) );
  NAND U13081 ( .A(ereg[50]), .B(n9759), .Z(n9959) );
  NANDN U13082 ( .A(n9754), .B(ereg[51]), .Z(n9958) );
  NAND U13083 ( .A(n9960), .B(n9961), .Z(n7646) );
  NANDN U13084 ( .A(init), .B(e[52]), .Z(n9961) );
  AND U13085 ( .A(n9962), .B(n9963), .Z(n9960) );
  NAND U13086 ( .A(ereg[51]), .B(n9759), .Z(n9963) );
  NANDN U13087 ( .A(n9754), .B(ereg[52]), .Z(n9962) );
  NAND U13088 ( .A(n9964), .B(n9965), .Z(n7645) );
  NANDN U13089 ( .A(init), .B(e[53]), .Z(n9965) );
  AND U13090 ( .A(n9966), .B(n9967), .Z(n9964) );
  NAND U13091 ( .A(ereg[52]), .B(n9759), .Z(n9967) );
  NANDN U13092 ( .A(n9754), .B(ereg[53]), .Z(n9966) );
  NAND U13093 ( .A(n9968), .B(n9969), .Z(n7644) );
  NANDN U13094 ( .A(init), .B(e[54]), .Z(n9969) );
  AND U13095 ( .A(n9970), .B(n9971), .Z(n9968) );
  NAND U13096 ( .A(ereg[53]), .B(n9759), .Z(n9971) );
  NANDN U13097 ( .A(n9754), .B(ereg[54]), .Z(n9970) );
  NAND U13098 ( .A(n9972), .B(n9973), .Z(n7643) );
  NANDN U13099 ( .A(init), .B(e[55]), .Z(n9973) );
  AND U13100 ( .A(n9974), .B(n9975), .Z(n9972) );
  NAND U13101 ( .A(ereg[54]), .B(n9759), .Z(n9975) );
  NANDN U13102 ( .A(n9754), .B(ereg[55]), .Z(n9974) );
  NAND U13103 ( .A(n9976), .B(n9977), .Z(n7642) );
  NANDN U13104 ( .A(init), .B(e[56]), .Z(n9977) );
  AND U13105 ( .A(n9978), .B(n9979), .Z(n9976) );
  NAND U13106 ( .A(ereg[55]), .B(n9759), .Z(n9979) );
  NANDN U13107 ( .A(n9754), .B(ereg[56]), .Z(n9978) );
  NAND U13108 ( .A(n9980), .B(n9981), .Z(n7641) );
  NANDN U13109 ( .A(init), .B(e[57]), .Z(n9981) );
  AND U13110 ( .A(n9982), .B(n9983), .Z(n9980) );
  NAND U13111 ( .A(ereg[56]), .B(n9759), .Z(n9983) );
  NANDN U13112 ( .A(n9754), .B(ereg[57]), .Z(n9982) );
  NAND U13113 ( .A(n9984), .B(n9985), .Z(n7640) );
  NANDN U13114 ( .A(init), .B(e[58]), .Z(n9985) );
  AND U13115 ( .A(n9986), .B(n9987), .Z(n9984) );
  NAND U13116 ( .A(ereg[57]), .B(n9759), .Z(n9987) );
  NANDN U13117 ( .A(n9754), .B(ereg[58]), .Z(n9986) );
  NAND U13118 ( .A(n9988), .B(n9989), .Z(n7639) );
  NANDN U13119 ( .A(init), .B(e[59]), .Z(n9989) );
  AND U13120 ( .A(n9990), .B(n9991), .Z(n9988) );
  NAND U13121 ( .A(ereg[58]), .B(n9759), .Z(n9991) );
  NANDN U13122 ( .A(n9754), .B(ereg[59]), .Z(n9990) );
  NAND U13123 ( .A(n9992), .B(n9993), .Z(n7638) );
  NANDN U13124 ( .A(init), .B(e[60]), .Z(n9993) );
  AND U13125 ( .A(n9994), .B(n9995), .Z(n9992) );
  NAND U13126 ( .A(ereg[59]), .B(n9759), .Z(n9995) );
  NANDN U13127 ( .A(n9754), .B(ereg[60]), .Z(n9994) );
  NAND U13128 ( .A(n9996), .B(n9997), .Z(n7637) );
  NANDN U13129 ( .A(init), .B(e[61]), .Z(n9997) );
  AND U13130 ( .A(n9998), .B(n9999), .Z(n9996) );
  NAND U13131 ( .A(ereg[60]), .B(n9759), .Z(n9999) );
  NANDN U13132 ( .A(n9754), .B(ereg[61]), .Z(n9998) );
  NAND U13133 ( .A(n10000), .B(n10001), .Z(n7636) );
  NANDN U13134 ( .A(init), .B(e[62]), .Z(n10001) );
  AND U13135 ( .A(n10002), .B(n10003), .Z(n10000) );
  NAND U13136 ( .A(ereg[61]), .B(n9759), .Z(n10003) );
  NANDN U13137 ( .A(n9754), .B(ereg[62]), .Z(n10002) );
  NAND U13138 ( .A(n10004), .B(n10005), .Z(n7635) );
  NANDN U13139 ( .A(init), .B(e[63]), .Z(n10005) );
  AND U13140 ( .A(n10006), .B(n10007), .Z(n10004) );
  NAND U13141 ( .A(ereg[62]), .B(n9759), .Z(n10007) );
  NANDN U13142 ( .A(n9754), .B(ereg[63]), .Z(n10006) );
  NAND U13143 ( .A(n10008), .B(n10009), .Z(n7634) );
  NANDN U13144 ( .A(init), .B(e[64]), .Z(n10009) );
  AND U13145 ( .A(n10010), .B(n10011), .Z(n10008) );
  NAND U13146 ( .A(ereg[63]), .B(n9759), .Z(n10011) );
  NANDN U13147 ( .A(n9754), .B(ereg[64]), .Z(n10010) );
  NAND U13148 ( .A(n10012), .B(n10013), .Z(n7633) );
  NANDN U13149 ( .A(init), .B(e[65]), .Z(n10013) );
  AND U13150 ( .A(n10014), .B(n10015), .Z(n10012) );
  NAND U13151 ( .A(ereg[64]), .B(n9759), .Z(n10015) );
  NANDN U13152 ( .A(n9754), .B(ereg[65]), .Z(n10014) );
  NAND U13153 ( .A(n10016), .B(n10017), .Z(n7632) );
  NANDN U13154 ( .A(init), .B(e[66]), .Z(n10017) );
  AND U13155 ( .A(n10018), .B(n10019), .Z(n10016) );
  NAND U13156 ( .A(ereg[65]), .B(n9759), .Z(n10019) );
  NANDN U13157 ( .A(n9754), .B(ereg[66]), .Z(n10018) );
  NAND U13158 ( .A(n10020), .B(n10021), .Z(n7631) );
  NANDN U13159 ( .A(init), .B(e[67]), .Z(n10021) );
  AND U13160 ( .A(n10022), .B(n10023), .Z(n10020) );
  NAND U13161 ( .A(ereg[66]), .B(n9759), .Z(n10023) );
  NANDN U13162 ( .A(n9754), .B(ereg[67]), .Z(n10022) );
  NAND U13163 ( .A(n10024), .B(n10025), .Z(n7630) );
  NANDN U13164 ( .A(init), .B(e[68]), .Z(n10025) );
  AND U13165 ( .A(n10026), .B(n10027), .Z(n10024) );
  NAND U13166 ( .A(ereg[67]), .B(n9759), .Z(n10027) );
  NANDN U13167 ( .A(n9754), .B(ereg[68]), .Z(n10026) );
  NAND U13168 ( .A(n10028), .B(n10029), .Z(n7629) );
  NANDN U13169 ( .A(init), .B(e[69]), .Z(n10029) );
  AND U13170 ( .A(n10030), .B(n10031), .Z(n10028) );
  NAND U13171 ( .A(ereg[68]), .B(n9759), .Z(n10031) );
  NANDN U13172 ( .A(n9754), .B(ereg[69]), .Z(n10030) );
  NAND U13173 ( .A(n10032), .B(n10033), .Z(n7628) );
  NANDN U13174 ( .A(init), .B(e[70]), .Z(n10033) );
  AND U13175 ( .A(n10034), .B(n10035), .Z(n10032) );
  NAND U13176 ( .A(ereg[69]), .B(n9759), .Z(n10035) );
  NANDN U13177 ( .A(n9754), .B(ereg[70]), .Z(n10034) );
  NAND U13178 ( .A(n10036), .B(n10037), .Z(n7627) );
  NANDN U13179 ( .A(init), .B(e[71]), .Z(n10037) );
  AND U13180 ( .A(n10038), .B(n10039), .Z(n10036) );
  NAND U13181 ( .A(ereg[70]), .B(n9759), .Z(n10039) );
  NANDN U13182 ( .A(n9754), .B(ereg[71]), .Z(n10038) );
  NAND U13183 ( .A(n10040), .B(n10041), .Z(n7626) );
  NANDN U13184 ( .A(init), .B(e[72]), .Z(n10041) );
  AND U13185 ( .A(n10042), .B(n10043), .Z(n10040) );
  NAND U13186 ( .A(ereg[71]), .B(n9759), .Z(n10043) );
  NANDN U13187 ( .A(n9754), .B(ereg[72]), .Z(n10042) );
  NAND U13188 ( .A(n10044), .B(n10045), .Z(n7625) );
  NANDN U13189 ( .A(init), .B(e[73]), .Z(n10045) );
  AND U13190 ( .A(n10046), .B(n10047), .Z(n10044) );
  NAND U13191 ( .A(ereg[72]), .B(n9759), .Z(n10047) );
  NANDN U13192 ( .A(n9754), .B(ereg[73]), .Z(n10046) );
  NAND U13193 ( .A(n10048), .B(n10049), .Z(n7624) );
  NANDN U13194 ( .A(init), .B(e[74]), .Z(n10049) );
  AND U13195 ( .A(n10050), .B(n10051), .Z(n10048) );
  NAND U13196 ( .A(ereg[73]), .B(n9759), .Z(n10051) );
  NANDN U13197 ( .A(n9754), .B(ereg[74]), .Z(n10050) );
  NAND U13198 ( .A(n10052), .B(n10053), .Z(n7623) );
  NANDN U13199 ( .A(init), .B(e[75]), .Z(n10053) );
  AND U13200 ( .A(n10054), .B(n10055), .Z(n10052) );
  NAND U13201 ( .A(ereg[74]), .B(n9759), .Z(n10055) );
  NANDN U13202 ( .A(n9754), .B(ereg[75]), .Z(n10054) );
  NAND U13203 ( .A(n10056), .B(n10057), .Z(n7622) );
  NANDN U13204 ( .A(init), .B(e[76]), .Z(n10057) );
  AND U13205 ( .A(n10058), .B(n10059), .Z(n10056) );
  NAND U13206 ( .A(ereg[75]), .B(n9759), .Z(n10059) );
  NANDN U13207 ( .A(n9754), .B(ereg[76]), .Z(n10058) );
  NAND U13208 ( .A(n10060), .B(n10061), .Z(n7621) );
  NANDN U13209 ( .A(init), .B(e[77]), .Z(n10061) );
  AND U13210 ( .A(n10062), .B(n10063), .Z(n10060) );
  NAND U13211 ( .A(ereg[76]), .B(n9759), .Z(n10063) );
  NANDN U13212 ( .A(n9754), .B(ereg[77]), .Z(n10062) );
  NAND U13213 ( .A(n10064), .B(n10065), .Z(n7620) );
  NANDN U13214 ( .A(init), .B(e[78]), .Z(n10065) );
  AND U13215 ( .A(n10066), .B(n10067), .Z(n10064) );
  NAND U13216 ( .A(ereg[77]), .B(n9759), .Z(n10067) );
  NANDN U13217 ( .A(n9754), .B(ereg[78]), .Z(n10066) );
  NAND U13218 ( .A(n10068), .B(n10069), .Z(n7619) );
  NANDN U13219 ( .A(init), .B(e[79]), .Z(n10069) );
  AND U13220 ( .A(n10070), .B(n10071), .Z(n10068) );
  NAND U13221 ( .A(ereg[78]), .B(n9759), .Z(n10071) );
  NANDN U13222 ( .A(n9754), .B(ereg[79]), .Z(n10070) );
  NAND U13223 ( .A(n10072), .B(n10073), .Z(n7618) );
  NANDN U13224 ( .A(init), .B(e[80]), .Z(n10073) );
  AND U13225 ( .A(n10074), .B(n10075), .Z(n10072) );
  NAND U13226 ( .A(ereg[79]), .B(n9759), .Z(n10075) );
  NANDN U13227 ( .A(n9754), .B(ereg[80]), .Z(n10074) );
  NAND U13228 ( .A(n10076), .B(n10077), .Z(n7617) );
  NANDN U13229 ( .A(init), .B(e[81]), .Z(n10077) );
  AND U13230 ( .A(n10078), .B(n10079), .Z(n10076) );
  NAND U13231 ( .A(ereg[80]), .B(n9759), .Z(n10079) );
  NANDN U13232 ( .A(n9754), .B(ereg[81]), .Z(n10078) );
  NAND U13233 ( .A(n10080), .B(n10081), .Z(n7616) );
  NANDN U13234 ( .A(init), .B(e[82]), .Z(n10081) );
  AND U13235 ( .A(n10082), .B(n10083), .Z(n10080) );
  NAND U13236 ( .A(ereg[81]), .B(n9759), .Z(n10083) );
  NANDN U13237 ( .A(n9754), .B(ereg[82]), .Z(n10082) );
  NAND U13238 ( .A(n10084), .B(n10085), .Z(n7615) );
  NANDN U13239 ( .A(init), .B(e[83]), .Z(n10085) );
  AND U13240 ( .A(n10086), .B(n10087), .Z(n10084) );
  NAND U13241 ( .A(ereg[82]), .B(n9759), .Z(n10087) );
  NANDN U13242 ( .A(n9754), .B(ereg[83]), .Z(n10086) );
  NAND U13243 ( .A(n10088), .B(n10089), .Z(n7614) );
  NANDN U13244 ( .A(init), .B(e[84]), .Z(n10089) );
  AND U13245 ( .A(n10090), .B(n10091), .Z(n10088) );
  NAND U13246 ( .A(ereg[83]), .B(n9759), .Z(n10091) );
  NANDN U13247 ( .A(n9754), .B(ereg[84]), .Z(n10090) );
  NAND U13248 ( .A(n10092), .B(n10093), .Z(n7613) );
  NANDN U13249 ( .A(init), .B(e[85]), .Z(n10093) );
  AND U13250 ( .A(n10094), .B(n10095), .Z(n10092) );
  NAND U13251 ( .A(ereg[84]), .B(n9759), .Z(n10095) );
  NANDN U13252 ( .A(n9754), .B(ereg[85]), .Z(n10094) );
  NAND U13253 ( .A(n10096), .B(n10097), .Z(n7612) );
  NANDN U13254 ( .A(init), .B(e[86]), .Z(n10097) );
  AND U13255 ( .A(n10098), .B(n10099), .Z(n10096) );
  NAND U13256 ( .A(ereg[85]), .B(n9759), .Z(n10099) );
  NANDN U13257 ( .A(n9754), .B(ereg[86]), .Z(n10098) );
  NAND U13258 ( .A(n10100), .B(n10101), .Z(n7611) );
  NANDN U13259 ( .A(init), .B(e[87]), .Z(n10101) );
  AND U13260 ( .A(n10102), .B(n10103), .Z(n10100) );
  NAND U13261 ( .A(ereg[86]), .B(n9759), .Z(n10103) );
  NANDN U13262 ( .A(n9754), .B(ereg[87]), .Z(n10102) );
  NAND U13263 ( .A(n10104), .B(n10105), .Z(n7610) );
  NANDN U13264 ( .A(init), .B(e[88]), .Z(n10105) );
  AND U13265 ( .A(n10106), .B(n10107), .Z(n10104) );
  NAND U13266 ( .A(ereg[87]), .B(n9759), .Z(n10107) );
  NANDN U13267 ( .A(n9754), .B(ereg[88]), .Z(n10106) );
  NAND U13268 ( .A(n10108), .B(n10109), .Z(n7609) );
  NANDN U13269 ( .A(init), .B(e[89]), .Z(n10109) );
  AND U13270 ( .A(n10110), .B(n10111), .Z(n10108) );
  NAND U13271 ( .A(ereg[88]), .B(n9759), .Z(n10111) );
  NANDN U13272 ( .A(n9754), .B(ereg[89]), .Z(n10110) );
  NAND U13273 ( .A(n10112), .B(n10113), .Z(n7608) );
  NANDN U13274 ( .A(init), .B(e[90]), .Z(n10113) );
  AND U13275 ( .A(n10114), .B(n10115), .Z(n10112) );
  NAND U13276 ( .A(ereg[89]), .B(n9759), .Z(n10115) );
  NANDN U13277 ( .A(n9754), .B(ereg[90]), .Z(n10114) );
  NAND U13278 ( .A(n10116), .B(n10117), .Z(n7607) );
  NANDN U13279 ( .A(init), .B(e[91]), .Z(n10117) );
  AND U13280 ( .A(n10118), .B(n10119), .Z(n10116) );
  NAND U13281 ( .A(ereg[90]), .B(n9759), .Z(n10119) );
  NANDN U13282 ( .A(n9754), .B(ereg[91]), .Z(n10118) );
  NAND U13283 ( .A(n10120), .B(n10121), .Z(n7606) );
  NANDN U13284 ( .A(init), .B(e[92]), .Z(n10121) );
  AND U13285 ( .A(n10122), .B(n10123), .Z(n10120) );
  NAND U13286 ( .A(ereg[91]), .B(n9759), .Z(n10123) );
  NANDN U13287 ( .A(n9754), .B(ereg[92]), .Z(n10122) );
  NAND U13288 ( .A(n10124), .B(n10125), .Z(n7605) );
  NANDN U13289 ( .A(init), .B(e[93]), .Z(n10125) );
  AND U13290 ( .A(n10126), .B(n10127), .Z(n10124) );
  NAND U13291 ( .A(ereg[92]), .B(n9759), .Z(n10127) );
  NANDN U13292 ( .A(n9754), .B(ereg[93]), .Z(n10126) );
  NAND U13293 ( .A(n10128), .B(n10129), .Z(n7604) );
  NANDN U13294 ( .A(init), .B(e[94]), .Z(n10129) );
  AND U13295 ( .A(n10130), .B(n10131), .Z(n10128) );
  NAND U13296 ( .A(ereg[93]), .B(n9759), .Z(n10131) );
  NANDN U13297 ( .A(n9754), .B(ereg[94]), .Z(n10130) );
  NAND U13298 ( .A(n10132), .B(n10133), .Z(n7603) );
  NANDN U13299 ( .A(init), .B(e[95]), .Z(n10133) );
  AND U13300 ( .A(n10134), .B(n10135), .Z(n10132) );
  NAND U13301 ( .A(ereg[94]), .B(n9759), .Z(n10135) );
  NANDN U13302 ( .A(n9754), .B(ereg[95]), .Z(n10134) );
  NAND U13303 ( .A(n10136), .B(n10137), .Z(n7602) );
  NANDN U13304 ( .A(init), .B(e[96]), .Z(n10137) );
  AND U13305 ( .A(n10138), .B(n10139), .Z(n10136) );
  NAND U13306 ( .A(ereg[95]), .B(n9759), .Z(n10139) );
  NANDN U13307 ( .A(n9754), .B(ereg[96]), .Z(n10138) );
  NAND U13308 ( .A(n10140), .B(n10141), .Z(n7601) );
  NANDN U13309 ( .A(init), .B(e[97]), .Z(n10141) );
  AND U13310 ( .A(n10142), .B(n10143), .Z(n10140) );
  NAND U13311 ( .A(ereg[96]), .B(n9759), .Z(n10143) );
  NANDN U13312 ( .A(n9754), .B(ereg[97]), .Z(n10142) );
  NAND U13313 ( .A(n10144), .B(n10145), .Z(n7600) );
  NANDN U13314 ( .A(init), .B(e[98]), .Z(n10145) );
  AND U13315 ( .A(n10146), .B(n10147), .Z(n10144) );
  NAND U13316 ( .A(ereg[97]), .B(n9759), .Z(n10147) );
  NANDN U13317 ( .A(n9754), .B(ereg[98]), .Z(n10146) );
  NAND U13318 ( .A(n10148), .B(n10149), .Z(n7599) );
  NANDN U13319 ( .A(init), .B(e[99]), .Z(n10149) );
  AND U13320 ( .A(n10150), .B(n10151), .Z(n10148) );
  NAND U13321 ( .A(ereg[98]), .B(n9759), .Z(n10151) );
  NANDN U13322 ( .A(n9754), .B(ereg[99]), .Z(n10150) );
  NAND U13323 ( .A(n10152), .B(n10153), .Z(n7598) );
  NANDN U13324 ( .A(init), .B(e[100]), .Z(n10153) );
  AND U13325 ( .A(n10154), .B(n10155), .Z(n10152) );
  NAND U13326 ( .A(ereg[99]), .B(n9759), .Z(n10155) );
  NANDN U13327 ( .A(n9754), .B(ereg[100]), .Z(n10154) );
  NAND U13328 ( .A(n10156), .B(n10157), .Z(n7597) );
  NANDN U13329 ( .A(init), .B(e[101]), .Z(n10157) );
  AND U13330 ( .A(n10158), .B(n10159), .Z(n10156) );
  NAND U13331 ( .A(ereg[100]), .B(n9759), .Z(n10159) );
  NANDN U13332 ( .A(n9754), .B(ereg[101]), .Z(n10158) );
  NAND U13333 ( .A(n10160), .B(n10161), .Z(n7596) );
  NANDN U13334 ( .A(init), .B(e[102]), .Z(n10161) );
  AND U13335 ( .A(n10162), .B(n10163), .Z(n10160) );
  NAND U13336 ( .A(ereg[101]), .B(n9759), .Z(n10163) );
  NANDN U13337 ( .A(n9754), .B(ereg[102]), .Z(n10162) );
  NAND U13338 ( .A(n10164), .B(n10165), .Z(n7595) );
  NANDN U13339 ( .A(init), .B(e[103]), .Z(n10165) );
  AND U13340 ( .A(n10166), .B(n10167), .Z(n10164) );
  NAND U13341 ( .A(ereg[102]), .B(n9759), .Z(n10167) );
  NANDN U13342 ( .A(n9754), .B(ereg[103]), .Z(n10166) );
  NAND U13343 ( .A(n10168), .B(n10169), .Z(n7594) );
  NANDN U13344 ( .A(init), .B(e[104]), .Z(n10169) );
  AND U13345 ( .A(n10170), .B(n10171), .Z(n10168) );
  NAND U13346 ( .A(ereg[103]), .B(n9759), .Z(n10171) );
  NANDN U13347 ( .A(n9754), .B(ereg[104]), .Z(n10170) );
  NAND U13348 ( .A(n10172), .B(n10173), .Z(n7593) );
  NANDN U13349 ( .A(init), .B(e[105]), .Z(n10173) );
  AND U13350 ( .A(n10174), .B(n10175), .Z(n10172) );
  NAND U13351 ( .A(ereg[104]), .B(n9759), .Z(n10175) );
  NANDN U13352 ( .A(n9754), .B(ereg[105]), .Z(n10174) );
  NAND U13353 ( .A(n10176), .B(n10177), .Z(n7592) );
  NANDN U13354 ( .A(init), .B(e[106]), .Z(n10177) );
  AND U13355 ( .A(n10178), .B(n10179), .Z(n10176) );
  NAND U13356 ( .A(ereg[105]), .B(n9759), .Z(n10179) );
  NANDN U13357 ( .A(n9754), .B(ereg[106]), .Z(n10178) );
  NAND U13358 ( .A(n10180), .B(n10181), .Z(n7591) );
  NANDN U13359 ( .A(init), .B(e[107]), .Z(n10181) );
  AND U13360 ( .A(n10182), .B(n10183), .Z(n10180) );
  NAND U13361 ( .A(ereg[106]), .B(n9759), .Z(n10183) );
  NANDN U13362 ( .A(n9754), .B(ereg[107]), .Z(n10182) );
  NAND U13363 ( .A(n10184), .B(n10185), .Z(n7590) );
  NANDN U13364 ( .A(init), .B(e[108]), .Z(n10185) );
  AND U13365 ( .A(n10186), .B(n10187), .Z(n10184) );
  NAND U13366 ( .A(ereg[107]), .B(n9759), .Z(n10187) );
  NANDN U13367 ( .A(n9754), .B(ereg[108]), .Z(n10186) );
  NAND U13368 ( .A(n10188), .B(n10189), .Z(n7589) );
  NANDN U13369 ( .A(init), .B(e[109]), .Z(n10189) );
  AND U13370 ( .A(n10190), .B(n10191), .Z(n10188) );
  NAND U13371 ( .A(ereg[108]), .B(n9759), .Z(n10191) );
  NANDN U13372 ( .A(n9754), .B(ereg[109]), .Z(n10190) );
  NAND U13373 ( .A(n10192), .B(n10193), .Z(n7588) );
  NANDN U13374 ( .A(init), .B(e[110]), .Z(n10193) );
  AND U13375 ( .A(n10194), .B(n10195), .Z(n10192) );
  NAND U13376 ( .A(ereg[109]), .B(n9759), .Z(n10195) );
  NANDN U13377 ( .A(n9754), .B(ereg[110]), .Z(n10194) );
  NAND U13378 ( .A(n10196), .B(n10197), .Z(n7587) );
  NANDN U13379 ( .A(init), .B(e[111]), .Z(n10197) );
  AND U13380 ( .A(n10198), .B(n10199), .Z(n10196) );
  NAND U13381 ( .A(ereg[110]), .B(n9759), .Z(n10199) );
  NANDN U13382 ( .A(n9754), .B(ereg[111]), .Z(n10198) );
  NAND U13383 ( .A(n10200), .B(n10201), .Z(n7586) );
  NANDN U13384 ( .A(init), .B(e[112]), .Z(n10201) );
  AND U13385 ( .A(n10202), .B(n10203), .Z(n10200) );
  NAND U13386 ( .A(ereg[111]), .B(n9759), .Z(n10203) );
  NANDN U13387 ( .A(n9754), .B(ereg[112]), .Z(n10202) );
  NAND U13388 ( .A(n10204), .B(n10205), .Z(n7585) );
  NANDN U13389 ( .A(init), .B(e[113]), .Z(n10205) );
  AND U13390 ( .A(n10206), .B(n10207), .Z(n10204) );
  NAND U13391 ( .A(ereg[112]), .B(n9759), .Z(n10207) );
  NANDN U13392 ( .A(n9754), .B(ereg[113]), .Z(n10206) );
  NAND U13393 ( .A(n10208), .B(n10209), .Z(n7584) );
  NANDN U13394 ( .A(init), .B(e[114]), .Z(n10209) );
  AND U13395 ( .A(n10210), .B(n10211), .Z(n10208) );
  NAND U13396 ( .A(ereg[113]), .B(n9759), .Z(n10211) );
  NANDN U13397 ( .A(n9754), .B(ereg[114]), .Z(n10210) );
  NAND U13398 ( .A(n10212), .B(n10213), .Z(n7583) );
  NANDN U13399 ( .A(init), .B(e[115]), .Z(n10213) );
  AND U13400 ( .A(n10214), .B(n10215), .Z(n10212) );
  NAND U13401 ( .A(ereg[114]), .B(n9759), .Z(n10215) );
  NANDN U13402 ( .A(n9754), .B(ereg[115]), .Z(n10214) );
  NAND U13403 ( .A(n10216), .B(n10217), .Z(n7582) );
  NANDN U13404 ( .A(init), .B(e[116]), .Z(n10217) );
  AND U13405 ( .A(n10218), .B(n10219), .Z(n10216) );
  NAND U13406 ( .A(ereg[115]), .B(n9759), .Z(n10219) );
  NANDN U13407 ( .A(n9754), .B(ereg[116]), .Z(n10218) );
  NAND U13408 ( .A(n10220), .B(n10221), .Z(n7581) );
  NANDN U13409 ( .A(init), .B(e[117]), .Z(n10221) );
  AND U13410 ( .A(n10222), .B(n10223), .Z(n10220) );
  NAND U13411 ( .A(ereg[116]), .B(n9759), .Z(n10223) );
  NANDN U13412 ( .A(n9754), .B(ereg[117]), .Z(n10222) );
  NAND U13413 ( .A(n10224), .B(n10225), .Z(n7580) );
  NANDN U13414 ( .A(init), .B(e[118]), .Z(n10225) );
  AND U13415 ( .A(n10226), .B(n10227), .Z(n10224) );
  NAND U13416 ( .A(ereg[117]), .B(n9759), .Z(n10227) );
  NANDN U13417 ( .A(n9754), .B(ereg[118]), .Z(n10226) );
  NAND U13418 ( .A(n10228), .B(n10229), .Z(n7579) );
  NANDN U13419 ( .A(init), .B(e[119]), .Z(n10229) );
  AND U13420 ( .A(n10230), .B(n10231), .Z(n10228) );
  NAND U13421 ( .A(ereg[118]), .B(n9759), .Z(n10231) );
  NANDN U13422 ( .A(n9754), .B(ereg[119]), .Z(n10230) );
  NAND U13423 ( .A(n10232), .B(n10233), .Z(n7578) );
  NANDN U13424 ( .A(init), .B(e[120]), .Z(n10233) );
  AND U13425 ( .A(n10234), .B(n10235), .Z(n10232) );
  NAND U13426 ( .A(ereg[119]), .B(n9759), .Z(n10235) );
  NANDN U13427 ( .A(n9754), .B(ereg[120]), .Z(n10234) );
  NAND U13428 ( .A(n10236), .B(n10237), .Z(n7577) );
  NANDN U13429 ( .A(init), .B(e[121]), .Z(n10237) );
  AND U13430 ( .A(n10238), .B(n10239), .Z(n10236) );
  NAND U13431 ( .A(ereg[120]), .B(n9759), .Z(n10239) );
  NANDN U13432 ( .A(n9754), .B(ereg[121]), .Z(n10238) );
  NAND U13433 ( .A(n10240), .B(n10241), .Z(n7576) );
  NANDN U13434 ( .A(init), .B(e[122]), .Z(n10241) );
  AND U13435 ( .A(n10242), .B(n10243), .Z(n10240) );
  NAND U13436 ( .A(ereg[121]), .B(n9759), .Z(n10243) );
  NANDN U13437 ( .A(n9754), .B(ereg[122]), .Z(n10242) );
  NAND U13438 ( .A(n10244), .B(n10245), .Z(n7575) );
  NANDN U13439 ( .A(init), .B(e[123]), .Z(n10245) );
  AND U13440 ( .A(n10246), .B(n10247), .Z(n10244) );
  NAND U13441 ( .A(ereg[122]), .B(n9759), .Z(n10247) );
  NANDN U13442 ( .A(n9754), .B(ereg[123]), .Z(n10246) );
  NAND U13443 ( .A(n10248), .B(n10249), .Z(n7574) );
  NANDN U13444 ( .A(init), .B(e[124]), .Z(n10249) );
  AND U13445 ( .A(n10250), .B(n10251), .Z(n10248) );
  NAND U13446 ( .A(ereg[123]), .B(n9759), .Z(n10251) );
  NANDN U13447 ( .A(n9754), .B(ereg[124]), .Z(n10250) );
  NAND U13448 ( .A(n10252), .B(n10253), .Z(n7573) );
  NANDN U13449 ( .A(init), .B(e[125]), .Z(n10253) );
  AND U13450 ( .A(n10254), .B(n10255), .Z(n10252) );
  NAND U13451 ( .A(ereg[124]), .B(n9759), .Z(n10255) );
  NANDN U13452 ( .A(n9754), .B(ereg[125]), .Z(n10254) );
  NAND U13453 ( .A(n10256), .B(n10257), .Z(n7572) );
  NANDN U13454 ( .A(init), .B(e[126]), .Z(n10257) );
  AND U13455 ( .A(n10258), .B(n10259), .Z(n10256) );
  NAND U13456 ( .A(ereg[125]), .B(n9759), .Z(n10259) );
  NANDN U13457 ( .A(n9754), .B(ereg[126]), .Z(n10258) );
  NAND U13458 ( .A(n10260), .B(n10261), .Z(n7571) );
  NANDN U13459 ( .A(init), .B(e[127]), .Z(n10261) );
  AND U13460 ( .A(n10262), .B(n10263), .Z(n10260) );
  NAND U13461 ( .A(ereg[126]), .B(n9759), .Z(n10263) );
  NANDN U13462 ( .A(n9754), .B(ereg[127]), .Z(n10262) );
  NAND U13463 ( .A(n10264), .B(n10265), .Z(n7570) );
  NANDN U13464 ( .A(init), .B(e[128]), .Z(n10265) );
  AND U13465 ( .A(n10266), .B(n10267), .Z(n10264) );
  NAND U13466 ( .A(ereg[127]), .B(n9759), .Z(n10267) );
  NANDN U13467 ( .A(n9754), .B(ereg[128]), .Z(n10266) );
  NAND U13468 ( .A(n10268), .B(n10269), .Z(n7569) );
  NANDN U13469 ( .A(init), .B(e[129]), .Z(n10269) );
  AND U13470 ( .A(n10270), .B(n10271), .Z(n10268) );
  NAND U13471 ( .A(ereg[128]), .B(n9759), .Z(n10271) );
  NANDN U13472 ( .A(n9754), .B(ereg[129]), .Z(n10270) );
  NAND U13473 ( .A(n10272), .B(n10273), .Z(n7568) );
  NANDN U13474 ( .A(init), .B(e[130]), .Z(n10273) );
  AND U13475 ( .A(n10274), .B(n10275), .Z(n10272) );
  NAND U13476 ( .A(ereg[129]), .B(n9759), .Z(n10275) );
  NANDN U13477 ( .A(n9754), .B(ereg[130]), .Z(n10274) );
  NAND U13478 ( .A(n10276), .B(n10277), .Z(n7567) );
  NANDN U13479 ( .A(init), .B(e[131]), .Z(n10277) );
  AND U13480 ( .A(n10278), .B(n10279), .Z(n10276) );
  NAND U13481 ( .A(ereg[130]), .B(n9759), .Z(n10279) );
  NANDN U13482 ( .A(n9754), .B(ereg[131]), .Z(n10278) );
  NAND U13483 ( .A(n10280), .B(n10281), .Z(n7566) );
  NANDN U13484 ( .A(init), .B(e[132]), .Z(n10281) );
  AND U13485 ( .A(n10282), .B(n10283), .Z(n10280) );
  NAND U13486 ( .A(ereg[131]), .B(n9759), .Z(n10283) );
  NANDN U13487 ( .A(n9754), .B(ereg[132]), .Z(n10282) );
  NAND U13488 ( .A(n10284), .B(n10285), .Z(n7565) );
  NANDN U13489 ( .A(init), .B(e[133]), .Z(n10285) );
  AND U13490 ( .A(n10286), .B(n10287), .Z(n10284) );
  NAND U13491 ( .A(ereg[132]), .B(n9759), .Z(n10287) );
  NANDN U13492 ( .A(n9754), .B(ereg[133]), .Z(n10286) );
  NAND U13493 ( .A(n10288), .B(n10289), .Z(n7564) );
  NANDN U13494 ( .A(init), .B(e[134]), .Z(n10289) );
  AND U13495 ( .A(n10290), .B(n10291), .Z(n10288) );
  NAND U13496 ( .A(ereg[133]), .B(n9759), .Z(n10291) );
  NANDN U13497 ( .A(n9754), .B(ereg[134]), .Z(n10290) );
  NAND U13498 ( .A(n10292), .B(n10293), .Z(n7563) );
  NANDN U13499 ( .A(init), .B(e[135]), .Z(n10293) );
  AND U13500 ( .A(n10294), .B(n10295), .Z(n10292) );
  NAND U13501 ( .A(ereg[134]), .B(n9759), .Z(n10295) );
  NANDN U13502 ( .A(n9754), .B(ereg[135]), .Z(n10294) );
  NAND U13503 ( .A(n10296), .B(n10297), .Z(n7562) );
  NANDN U13504 ( .A(init), .B(e[136]), .Z(n10297) );
  AND U13505 ( .A(n10298), .B(n10299), .Z(n10296) );
  NAND U13506 ( .A(ereg[135]), .B(n9759), .Z(n10299) );
  NANDN U13507 ( .A(n9754), .B(ereg[136]), .Z(n10298) );
  NAND U13508 ( .A(n10300), .B(n10301), .Z(n7561) );
  NANDN U13509 ( .A(init), .B(e[137]), .Z(n10301) );
  AND U13510 ( .A(n10302), .B(n10303), .Z(n10300) );
  NAND U13511 ( .A(ereg[136]), .B(n9759), .Z(n10303) );
  NANDN U13512 ( .A(n9754), .B(ereg[137]), .Z(n10302) );
  NAND U13513 ( .A(n10304), .B(n10305), .Z(n7560) );
  NANDN U13514 ( .A(init), .B(e[138]), .Z(n10305) );
  AND U13515 ( .A(n10306), .B(n10307), .Z(n10304) );
  NAND U13516 ( .A(ereg[137]), .B(n9759), .Z(n10307) );
  NANDN U13517 ( .A(n9754), .B(ereg[138]), .Z(n10306) );
  NAND U13518 ( .A(n10308), .B(n10309), .Z(n7559) );
  NANDN U13519 ( .A(init), .B(e[139]), .Z(n10309) );
  AND U13520 ( .A(n10310), .B(n10311), .Z(n10308) );
  NAND U13521 ( .A(ereg[138]), .B(n9759), .Z(n10311) );
  NANDN U13522 ( .A(n9754), .B(ereg[139]), .Z(n10310) );
  NAND U13523 ( .A(n10312), .B(n10313), .Z(n7558) );
  NANDN U13524 ( .A(init), .B(e[140]), .Z(n10313) );
  AND U13525 ( .A(n10314), .B(n10315), .Z(n10312) );
  NAND U13526 ( .A(ereg[139]), .B(n9759), .Z(n10315) );
  NANDN U13527 ( .A(n9754), .B(ereg[140]), .Z(n10314) );
  NAND U13528 ( .A(n10316), .B(n10317), .Z(n7557) );
  NANDN U13529 ( .A(init), .B(e[141]), .Z(n10317) );
  AND U13530 ( .A(n10318), .B(n10319), .Z(n10316) );
  NAND U13531 ( .A(ereg[140]), .B(n9759), .Z(n10319) );
  NANDN U13532 ( .A(n9754), .B(ereg[141]), .Z(n10318) );
  NAND U13533 ( .A(n10320), .B(n10321), .Z(n7556) );
  NANDN U13534 ( .A(init), .B(e[142]), .Z(n10321) );
  AND U13535 ( .A(n10322), .B(n10323), .Z(n10320) );
  NAND U13536 ( .A(ereg[141]), .B(n9759), .Z(n10323) );
  NANDN U13537 ( .A(n9754), .B(ereg[142]), .Z(n10322) );
  NAND U13538 ( .A(n10324), .B(n10325), .Z(n7555) );
  NANDN U13539 ( .A(init), .B(e[143]), .Z(n10325) );
  AND U13540 ( .A(n10326), .B(n10327), .Z(n10324) );
  NAND U13541 ( .A(ereg[142]), .B(n9759), .Z(n10327) );
  NANDN U13542 ( .A(n9754), .B(ereg[143]), .Z(n10326) );
  NAND U13543 ( .A(n10328), .B(n10329), .Z(n7554) );
  NANDN U13544 ( .A(init), .B(e[144]), .Z(n10329) );
  AND U13545 ( .A(n10330), .B(n10331), .Z(n10328) );
  NAND U13546 ( .A(ereg[143]), .B(n9759), .Z(n10331) );
  NANDN U13547 ( .A(n9754), .B(ereg[144]), .Z(n10330) );
  NAND U13548 ( .A(n10332), .B(n10333), .Z(n7553) );
  NANDN U13549 ( .A(init), .B(e[145]), .Z(n10333) );
  AND U13550 ( .A(n10334), .B(n10335), .Z(n10332) );
  NAND U13551 ( .A(ereg[144]), .B(n9759), .Z(n10335) );
  NANDN U13552 ( .A(n9754), .B(ereg[145]), .Z(n10334) );
  NAND U13553 ( .A(n10336), .B(n10337), .Z(n7552) );
  NANDN U13554 ( .A(init), .B(e[146]), .Z(n10337) );
  AND U13555 ( .A(n10338), .B(n10339), .Z(n10336) );
  NAND U13556 ( .A(ereg[145]), .B(n9759), .Z(n10339) );
  NANDN U13557 ( .A(n9754), .B(ereg[146]), .Z(n10338) );
  NAND U13558 ( .A(n10340), .B(n10341), .Z(n7551) );
  NANDN U13559 ( .A(init), .B(e[147]), .Z(n10341) );
  AND U13560 ( .A(n10342), .B(n10343), .Z(n10340) );
  NAND U13561 ( .A(ereg[146]), .B(n9759), .Z(n10343) );
  NANDN U13562 ( .A(n9754), .B(ereg[147]), .Z(n10342) );
  NAND U13563 ( .A(n10344), .B(n10345), .Z(n7550) );
  NANDN U13564 ( .A(init), .B(e[148]), .Z(n10345) );
  AND U13565 ( .A(n10346), .B(n10347), .Z(n10344) );
  NAND U13566 ( .A(ereg[147]), .B(n9759), .Z(n10347) );
  NANDN U13567 ( .A(n9754), .B(ereg[148]), .Z(n10346) );
  NAND U13568 ( .A(n10348), .B(n10349), .Z(n7549) );
  NANDN U13569 ( .A(init), .B(e[149]), .Z(n10349) );
  AND U13570 ( .A(n10350), .B(n10351), .Z(n10348) );
  NAND U13571 ( .A(ereg[148]), .B(n9759), .Z(n10351) );
  NANDN U13572 ( .A(n9754), .B(ereg[149]), .Z(n10350) );
  NAND U13573 ( .A(n10352), .B(n10353), .Z(n7548) );
  NANDN U13574 ( .A(init), .B(e[150]), .Z(n10353) );
  AND U13575 ( .A(n10354), .B(n10355), .Z(n10352) );
  NAND U13576 ( .A(ereg[149]), .B(n9759), .Z(n10355) );
  NANDN U13577 ( .A(n9754), .B(ereg[150]), .Z(n10354) );
  NAND U13578 ( .A(n10356), .B(n10357), .Z(n7547) );
  NANDN U13579 ( .A(init), .B(e[151]), .Z(n10357) );
  AND U13580 ( .A(n10358), .B(n10359), .Z(n10356) );
  NAND U13581 ( .A(ereg[150]), .B(n9759), .Z(n10359) );
  NANDN U13582 ( .A(n9754), .B(ereg[151]), .Z(n10358) );
  NAND U13583 ( .A(n10360), .B(n10361), .Z(n7546) );
  NANDN U13584 ( .A(init), .B(e[152]), .Z(n10361) );
  AND U13585 ( .A(n10362), .B(n10363), .Z(n10360) );
  NAND U13586 ( .A(ereg[151]), .B(n9759), .Z(n10363) );
  NANDN U13587 ( .A(n9754), .B(ereg[152]), .Z(n10362) );
  NAND U13588 ( .A(n10364), .B(n10365), .Z(n7545) );
  NANDN U13589 ( .A(init), .B(e[153]), .Z(n10365) );
  AND U13590 ( .A(n10366), .B(n10367), .Z(n10364) );
  NAND U13591 ( .A(ereg[152]), .B(n9759), .Z(n10367) );
  NANDN U13592 ( .A(n9754), .B(ereg[153]), .Z(n10366) );
  NAND U13593 ( .A(n10368), .B(n10369), .Z(n7544) );
  NANDN U13594 ( .A(init), .B(e[154]), .Z(n10369) );
  AND U13595 ( .A(n10370), .B(n10371), .Z(n10368) );
  NAND U13596 ( .A(ereg[153]), .B(n9759), .Z(n10371) );
  NANDN U13597 ( .A(n9754), .B(ereg[154]), .Z(n10370) );
  NAND U13598 ( .A(n10372), .B(n10373), .Z(n7543) );
  NANDN U13599 ( .A(init), .B(e[155]), .Z(n10373) );
  AND U13600 ( .A(n10374), .B(n10375), .Z(n10372) );
  NAND U13601 ( .A(ereg[154]), .B(n9759), .Z(n10375) );
  NANDN U13602 ( .A(n9754), .B(ereg[155]), .Z(n10374) );
  NAND U13603 ( .A(n10376), .B(n10377), .Z(n7542) );
  NANDN U13604 ( .A(init), .B(e[156]), .Z(n10377) );
  AND U13605 ( .A(n10378), .B(n10379), .Z(n10376) );
  NAND U13606 ( .A(ereg[155]), .B(n9759), .Z(n10379) );
  NANDN U13607 ( .A(n9754), .B(ereg[156]), .Z(n10378) );
  NAND U13608 ( .A(n10380), .B(n10381), .Z(n7541) );
  NANDN U13609 ( .A(init), .B(e[157]), .Z(n10381) );
  AND U13610 ( .A(n10382), .B(n10383), .Z(n10380) );
  NAND U13611 ( .A(ereg[156]), .B(n9759), .Z(n10383) );
  NANDN U13612 ( .A(n9754), .B(ereg[157]), .Z(n10382) );
  NAND U13613 ( .A(n10384), .B(n10385), .Z(n7540) );
  NANDN U13614 ( .A(init), .B(e[158]), .Z(n10385) );
  AND U13615 ( .A(n10386), .B(n10387), .Z(n10384) );
  NAND U13616 ( .A(ereg[157]), .B(n9759), .Z(n10387) );
  NANDN U13617 ( .A(n9754), .B(ereg[158]), .Z(n10386) );
  NAND U13618 ( .A(n10388), .B(n10389), .Z(n7539) );
  NANDN U13619 ( .A(init), .B(e[159]), .Z(n10389) );
  AND U13620 ( .A(n10390), .B(n10391), .Z(n10388) );
  NAND U13621 ( .A(ereg[158]), .B(n9759), .Z(n10391) );
  NANDN U13622 ( .A(n9754), .B(ereg[159]), .Z(n10390) );
  NAND U13623 ( .A(n10392), .B(n10393), .Z(n7538) );
  NANDN U13624 ( .A(init), .B(e[160]), .Z(n10393) );
  AND U13625 ( .A(n10394), .B(n10395), .Z(n10392) );
  NAND U13626 ( .A(ereg[159]), .B(n9759), .Z(n10395) );
  NANDN U13627 ( .A(n9754), .B(ereg[160]), .Z(n10394) );
  NAND U13628 ( .A(n10396), .B(n10397), .Z(n7537) );
  NANDN U13629 ( .A(init), .B(e[161]), .Z(n10397) );
  AND U13630 ( .A(n10398), .B(n10399), .Z(n10396) );
  NAND U13631 ( .A(ereg[160]), .B(n9759), .Z(n10399) );
  NANDN U13632 ( .A(n9754), .B(ereg[161]), .Z(n10398) );
  NAND U13633 ( .A(n10400), .B(n10401), .Z(n7536) );
  NANDN U13634 ( .A(init), .B(e[162]), .Z(n10401) );
  AND U13635 ( .A(n10402), .B(n10403), .Z(n10400) );
  NAND U13636 ( .A(ereg[161]), .B(n9759), .Z(n10403) );
  NANDN U13637 ( .A(n9754), .B(ereg[162]), .Z(n10402) );
  NAND U13638 ( .A(n10404), .B(n10405), .Z(n7535) );
  NANDN U13639 ( .A(init), .B(e[163]), .Z(n10405) );
  AND U13640 ( .A(n10406), .B(n10407), .Z(n10404) );
  NAND U13641 ( .A(ereg[162]), .B(n9759), .Z(n10407) );
  NANDN U13642 ( .A(n9754), .B(ereg[163]), .Z(n10406) );
  NAND U13643 ( .A(n10408), .B(n10409), .Z(n7534) );
  NANDN U13644 ( .A(init), .B(e[164]), .Z(n10409) );
  AND U13645 ( .A(n10410), .B(n10411), .Z(n10408) );
  NAND U13646 ( .A(ereg[163]), .B(n9759), .Z(n10411) );
  NANDN U13647 ( .A(n9754), .B(ereg[164]), .Z(n10410) );
  NAND U13648 ( .A(n10412), .B(n10413), .Z(n7533) );
  NANDN U13649 ( .A(init), .B(e[165]), .Z(n10413) );
  AND U13650 ( .A(n10414), .B(n10415), .Z(n10412) );
  NAND U13651 ( .A(ereg[164]), .B(n9759), .Z(n10415) );
  NANDN U13652 ( .A(n9754), .B(ereg[165]), .Z(n10414) );
  NAND U13653 ( .A(n10416), .B(n10417), .Z(n7532) );
  NANDN U13654 ( .A(init), .B(e[166]), .Z(n10417) );
  AND U13655 ( .A(n10418), .B(n10419), .Z(n10416) );
  NAND U13656 ( .A(ereg[165]), .B(n9759), .Z(n10419) );
  NANDN U13657 ( .A(n9754), .B(ereg[166]), .Z(n10418) );
  NAND U13658 ( .A(n10420), .B(n10421), .Z(n7531) );
  NANDN U13659 ( .A(init), .B(e[167]), .Z(n10421) );
  AND U13660 ( .A(n10422), .B(n10423), .Z(n10420) );
  NAND U13661 ( .A(ereg[166]), .B(n9759), .Z(n10423) );
  NANDN U13662 ( .A(n9754), .B(ereg[167]), .Z(n10422) );
  NAND U13663 ( .A(n10424), .B(n10425), .Z(n7530) );
  NANDN U13664 ( .A(init), .B(e[168]), .Z(n10425) );
  AND U13665 ( .A(n10426), .B(n10427), .Z(n10424) );
  NAND U13666 ( .A(ereg[167]), .B(n9759), .Z(n10427) );
  NANDN U13667 ( .A(n9754), .B(ereg[168]), .Z(n10426) );
  NAND U13668 ( .A(n10428), .B(n10429), .Z(n7529) );
  NANDN U13669 ( .A(init), .B(e[169]), .Z(n10429) );
  AND U13670 ( .A(n10430), .B(n10431), .Z(n10428) );
  NAND U13671 ( .A(ereg[168]), .B(n9759), .Z(n10431) );
  NANDN U13672 ( .A(n9754), .B(ereg[169]), .Z(n10430) );
  NAND U13673 ( .A(n10432), .B(n10433), .Z(n7528) );
  NANDN U13674 ( .A(init), .B(e[170]), .Z(n10433) );
  AND U13675 ( .A(n10434), .B(n10435), .Z(n10432) );
  NAND U13676 ( .A(ereg[169]), .B(n9759), .Z(n10435) );
  NANDN U13677 ( .A(n9754), .B(ereg[170]), .Z(n10434) );
  NAND U13678 ( .A(n10436), .B(n10437), .Z(n7527) );
  NANDN U13679 ( .A(init), .B(e[171]), .Z(n10437) );
  AND U13680 ( .A(n10438), .B(n10439), .Z(n10436) );
  NAND U13681 ( .A(ereg[170]), .B(n9759), .Z(n10439) );
  NANDN U13682 ( .A(n9754), .B(ereg[171]), .Z(n10438) );
  NAND U13683 ( .A(n10440), .B(n10441), .Z(n7526) );
  NANDN U13684 ( .A(init), .B(e[172]), .Z(n10441) );
  AND U13685 ( .A(n10442), .B(n10443), .Z(n10440) );
  NAND U13686 ( .A(ereg[171]), .B(n9759), .Z(n10443) );
  NANDN U13687 ( .A(n9754), .B(ereg[172]), .Z(n10442) );
  NAND U13688 ( .A(n10444), .B(n10445), .Z(n7525) );
  NANDN U13689 ( .A(init), .B(e[173]), .Z(n10445) );
  AND U13690 ( .A(n10446), .B(n10447), .Z(n10444) );
  NAND U13691 ( .A(ereg[172]), .B(n9759), .Z(n10447) );
  NANDN U13692 ( .A(n9754), .B(ereg[173]), .Z(n10446) );
  NAND U13693 ( .A(n10448), .B(n10449), .Z(n7524) );
  NANDN U13694 ( .A(init), .B(e[174]), .Z(n10449) );
  AND U13695 ( .A(n10450), .B(n10451), .Z(n10448) );
  NAND U13696 ( .A(ereg[173]), .B(n9759), .Z(n10451) );
  NANDN U13697 ( .A(n9754), .B(ereg[174]), .Z(n10450) );
  NAND U13698 ( .A(n10452), .B(n10453), .Z(n7523) );
  NANDN U13699 ( .A(init), .B(e[175]), .Z(n10453) );
  AND U13700 ( .A(n10454), .B(n10455), .Z(n10452) );
  NAND U13701 ( .A(ereg[174]), .B(n9759), .Z(n10455) );
  NANDN U13702 ( .A(n9754), .B(ereg[175]), .Z(n10454) );
  NAND U13703 ( .A(n10456), .B(n10457), .Z(n7522) );
  NANDN U13704 ( .A(init), .B(e[176]), .Z(n10457) );
  AND U13705 ( .A(n10458), .B(n10459), .Z(n10456) );
  NAND U13706 ( .A(ereg[175]), .B(n9759), .Z(n10459) );
  NANDN U13707 ( .A(n9754), .B(ereg[176]), .Z(n10458) );
  NAND U13708 ( .A(n10460), .B(n10461), .Z(n7521) );
  NANDN U13709 ( .A(init), .B(e[177]), .Z(n10461) );
  AND U13710 ( .A(n10462), .B(n10463), .Z(n10460) );
  NAND U13711 ( .A(ereg[176]), .B(n9759), .Z(n10463) );
  NANDN U13712 ( .A(n9754), .B(ereg[177]), .Z(n10462) );
  NAND U13713 ( .A(n10464), .B(n10465), .Z(n7520) );
  NANDN U13714 ( .A(init), .B(e[178]), .Z(n10465) );
  AND U13715 ( .A(n10466), .B(n10467), .Z(n10464) );
  NAND U13716 ( .A(ereg[177]), .B(n9759), .Z(n10467) );
  NANDN U13717 ( .A(n9754), .B(ereg[178]), .Z(n10466) );
  NAND U13718 ( .A(n10468), .B(n10469), .Z(n7519) );
  NANDN U13719 ( .A(init), .B(e[179]), .Z(n10469) );
  AND U13720 ( .A(n10470), .B(n10471), .Z(n10468) );
  NAND U13721 ( .A(ereg[178]), .B(n9759), .Z(n10471) );
  NANDN U13722 ( .A(n9754), .B(ereg[179]), .Z(n10470) );
  NAND U13723 ( .A(n10472), .B(n10473), .Z(n7518) );
  NANDN U13724 ( .A(init), .B(e[180]), .Z(n10473) );
  AND U13725 ( .A(n10474), .B(n10475), .Z(n10472) );
  NAND U13726 ( .A(ereg[179]), .B(n9759), .Z(n10475) );
  NANDN U13727 ( .A(n9754), .B(ereg[180]), .Z(n10474) );
  NAND U13728 ( .A(n10476), .B(n10477), .Z(n7517) );
  NANDN U13729 ( .A(init), .B(e[181]), .Z(n10477) );
  AND U13730 ( .A(n10478), .B(n10479), .Z(n10476) );
  NAND U13731 ( .A(ereg[180]), .B(n9759), .Z(n10479) );
  NANDN U13732 ( .A(n9754), .B(ereg[181]), .Z(n10478) );
  NAND U13733 ( .A(n10480), .B(n10481), .Z(n7516) );
  NANDN U13734 ( .A(init), .B(e[182]), .Z(n10481) );
  AND U13735 ( .A(n10482), .B(n10483), .Z(n10480) );
  NAND U13736 ( .A(ereg[181]), .B(n9759), .Z(n10483) );
  NANDN U13737 ( .A(n9754), .B(ereg[182]), .Z(n10482) );
  NAND U13738 ( .A(n10484), .B(n10485), .Z(n7515) );
  NANDN U13739 ( .A(init), .B(e[183]), .Z(n10485) );
  AND U13740 ( .A(n10486), .B(n10487), .Z(n10484) );
  NAND U13741 ( .A(ereg[182]), .B(n9759), .Z(n10487) );
  NANDN U13742 ( .A(n9754), .B(ereg[183]), .Z(n10486) );
  NAND U13743 ( .A(n10488), .B(n10489), .Z(n7514) );
  NANDN U13744 ( .A(init), .B(e[184]), .Z(n10489) );
  AND U13745 ( .A(n10490), .B(n10491), .Z(n10488) );
  NAND U13746 ( .A(ereg[183]), .B(n9759), .Z(n10491) );
  NANDN U13747 ( .A(n9754), .B(ereg[184]), .Z(n10490) );
  NAND U13748 ( .A(n10492), .B(n10493), .Z(n7513) );
  NANDN U13749 ( .A(init), .B(e[185]), .Z(n10493) );
  AND U13750 ( .A(n10494), .B(n10495), .Z(n10492) );
  NAND U13751 ( .A(ereg[184]), .B(n9759), .Z(n10495) );
  NANDN U13752 ( .A(n9754), .B(ereg[185]), .Z(n10494) );
  NAND U13753 ( .A(n10496), .B(n10497), .Z(n7512) );
  NANDN U13754 ( .A(init), .B(e[186]), .Z(n10497) );
  AND U13755 ( .A(n10498), .B(n10499), .Z(n10496) );
  NAND U13756 ( .A(ereg[185]), .B(n9759), .Z(n10499) );
  NANDN U13757 ( .A(n9754), .B(ereg[186]), .Z(n10498) );
  NAND U13758 ( .A(n10500), .B(n10501), .Z(n7511) );
  NANDN U13759 ( .A(init), .B(e[187]), .Z(n10501) );
  AND U13760 ( .A(n10502), .B(n10503), .Z(n10500) );
  NAND U13761 ( .A(ereg[186]), .B(n9759), .Z(n10503) );
  NANDN U13762 ( .A(n9754), .B(ereg[187]), .Z(n10502) );
  NAND U13763 ( .A(n10504), .B(n10505), .Z(n7510) );
  NANDN U13764 ( .A(init), .B(e[188]), .Z(n10505) );
  AND U13765 ( .A(n10506), .B(n10507), .Z(n10504) );
  NAND U13766 ( .A(ereg[187]), .B(n9759), .Z(n10507) );
  NANDN U13767 ( .A(n9754), .B(ereg[188]), .Z(n10506) );
  NAND U13768 ( .A(n10508), .B(n10509), .Z(n7509) );
  NANDN U13769 ( .A(init), .B(e[189]), .Z(n10509) );
  AND U13770 ( .A(n10510), .B(n10511), .Z(n10508) );
  NAND U13771 ( .A(ereg[188]), .B(n9759), .Z(n10511) );
  NANDN U13772 ( .A(n9754), .B(ereg[189]), .Z(n10510) );
  NAND U13773 ( .A(n10512), .B(n10513), .Z(n7508) );
  NANDN U13774 ( .A(init), .B(e[190]), .Z(n10513) );
  AND U13775 ( .A(n10514), .B(n10515), .Z(n10512) );
  NAND U13776 ( .A(ereg[189]), .B(n9759), .Z(n10515) );
  NANDN U13777 ( .A(n9754), .B(ereg[190]), .Z(n10514) );
  NAND U13778 ( .A(n10516), .B(n10517), .Z(n7507) );
  NANDN U13779 ( .A(init), .B(e[191]), .Z(n10517) );
  AND U13780 ( .A(n10518), .B(n10519), .Z(n10516) );
  NAND U13781 ( .A(ereg[190]), .B(n9759), .Z(n10519) );
  NANDN U13782 ( .A(n9754), .B(ereg[191]), .Z(n10518) );
  NAND U13783 ( .A(n10520), .B(n10521), .Z(n7506) );
  NANDN U13784 ( .A(init), .B(e[192]), .Z(n10521) );
  AND U13785 ( .A(n10522), .B(n10523), .Z(n10520) );
  NAND U13786 ( .A(ereg[191]), .B(n9759), .Z(n10523) );
  NANDN U13787 ( .A(n9754), .B(ereg[192]), .Z(n10522) );
  NAND U13788 ( .A(n10524), .B(n10525), .Z(n7505) );
  NANDN U13789 ( .A(init), .B(e[193]), .Z(n10525) );
  AND U13790 ( .A(n10526), .B(n10527), .Z(n10524) );
  NAND U13791 ( .A(ereg[192]), .B(n9759), .Z(n10527) );
  NANDN U13792 ( .A(n9754), .B(ereg[193]), .Z(n10526) );
  NAND U13793 ( .A(n10528), .B(n10529), .Z(n7504) );
  NANDN U13794 ( .A(init), .B(e[194]), .Z(n10529) );
  AND U13795 ( .A(n10530), .B(n10531), .Z(n10528) );
  NAND U13796 ( .A(ereg[193]), .B(n9759), .Z(n10531) );
  NANDN U13797 ( .A(n9754), .B(ereg[194]), .Z(n10530) );
  NAND U13798 ( .A(n10532), .B(n10533), .Z(n7503) );
  NANDN U13799 ( .A(init), .B(e[195]), .Z(n10533) );
  AND U13800 ( .A(n10534), .B(n10535), .Z(n10532) );
  NAND U13801 ( .A(ereg[194]), .B(n9759), .Z(n10535) );
  NANDN U13802 ( .A(n9754), .B(ereg[195]), .Z(n10534) );
  NAND U13803 ( .A(n10536), .B(n10537), .Z(n7502) );
  NANDN U13804 ( .A(init), .B(e[196]), .Z(n10537) );
  AND U13805 ( .A(n10538), .B(n10539), .Z(n10536) );
  NAND U13806 ( .A(ereg[195]), .B(n9759), .Z(n10539) );
  NANDN U13807 ( .A(n9754), .B(ereg[196]), .Z(n10538) );
  NAND U13808 ( .A(n10540), .B(n10541), .Z(n7501) );
  NANDN U13809 ( .A(init), .B(e[197]), .Z(n10541) );
  AND U13810 ( .A(n10542), .B(n10543), .Z(n10540) );
  NAND U13811 ( .A(ereg[196]), .B(n9759), .Z(n10543) );
  NANDN U13812 ( .A(n9754), .B(ereg[197]), .Z(n10542) );
  NAND U13813 ( .A(n10544), .B(n10545), .Z(n7500) );
  NANDN U13814 ( .A(init), .B(e[198]), .Z(n10545) );
  AND U13815 ( .A(n10546), .B(n10547), .Z(n10544) );
  NAND U13816 ( .A(ereg[197]), .B(n9759), .Z(n10547) );
  NANDN U13817 ( .A(n9754), .B(ereg[198]), .Z(n10546) );
  NAND U13818 ( .A(n10548), .B(n10549), .Z(n7499) );
  NANDN U13819 ( .A(init), .B(e[199]), .Z(n10549) );
  AND U13820 ( .A(n10550), .B(n10551), .Z(n10548) );
  NAND U13821 ( .A(ereg[198]), .B(n9759), .Z(n10551) );
  NANDN U13822 ( .A(n9754), .B(ereg[199]), .Z(n10550) );
  NAND U13823 ( .A(n10552), .B(n10553), .Z(n7498) );
  NANDN U13824 ( .A(init), .B(e[200]), .Z(n10553) );
  AND U13825 ( .A(n10554), .B(n10555), .Z(n10552) );
  NAND U13826 ( .A(ereg[199]), .B(n9759), .Z(n10555) );
  NANDN U13827 ( .A(n9754), .B(ereg[200]), .Z(n10554) );
  NAND U13828 ( .A(n10556), .B(n10557), .Z(n7497) );
  NANDN U13829 ( .A(init), .B(e[201]), .Z(n10557) );
  AND U13830 ( .A(n10558), .B(n10559), .Z(n10556) );
  NAND U13831 ( .A(ereg[200]), .B(n9759), .Z(n10559) );
  NANDN U13832 ( .A(n9754), .B(ereg[201]), .Z(n10558) );
  NAND U13833 ( .A(n10560), .B(n10561), .Z(n7496) );
  NANDN U13834 ( .A(init), .B(e[202]), .Z(n10561) );
  AND U13835 ( .A(n10562), .B(n10563), .Z(n10560) );
  NAND U13836 ( .A(ereg[201]), .B(n9759), .Z(n10563) );
  NANDN U13837 ( .A(n9754), .B(ereg[202]), .Z(n10562) );
  NAND U13838 ( .A(n10564), .B(n10565), .Z(n7495) );
  NANDN U13839 ( .A(init), .B(e[203]), .Z(n10565) );
  AND U13840 ( .A(n10566), .B(n10567), .Z(n10564) );
  NAND U13841 ( .A(ereg[202]), .B(n9759), .Z(n10567) );
  NANDN U13842 ( .A(n9754), .B(ereg[203]), .Z(n10566) );
  NAND U13843 ( .A(n10568), .B(n10569), .Z(n7494) );
  NANDN U13844 ( .A(init), .B(e[204]), .Z(n10569) );
  AND U13845 ( .A(n10570), .B(n10571), .Z(n10568) );
  NAND U13846 ( .A(ereg[203]), .B(n9759), .Z(n10571) );
  NANDN U13847 ( .A(n9754), .B(ereg[204]), .Z(n10570) );
  NAND U13848 ( .A(n10572), .B(n10573), .Z(n7493) );
  NANDN U13849 ( .A(init), .B(e[205]), .Z(n10573) );
  AND U13850 ( .A(n10574), .B(n10575), .Z(n10572) );
  NAND U13851 ( .A(ereg[204]), .B(n9759), .Z(n10575) );
  NANDN U13852 ( .A(n9754), .B(ereg[205]), .Z(n10574) );
  NAND U13853 ( .A(n10576), .B(n10577), .Z(n7492) );
  NANDN U13854 ( .A(init), .B(e[206]), .Z(n10577) );
  AND U13855 ( .A(n10578), .B(n10579), .Z(n10576) );
  NAND U13856 ( .A(ereg[205]), .B(n9759), .Z(n10579) );
  NANDN U13857 ( .A(n9754), .B(ereg[206]), .Z(n10578) );
  NAND U13858 ( .A(n10580), .B(n10581), .Z(n7491) );
  NANDN U13859 ( .A(init), .B(e[207]), .Z(n10581) );
  AND U13860 ( .A(n10582), .B(n10583), .Z(n10580) );
  NAND U13861 ( .A(ereg[206]), .B(n9759), .Z(n10583) );
  NANDN U13862 ( .A(n9754), .B(ereg[207]), .Z(n10582) );
  NAND U13863 ( .A(n10584), .B(n10585), .Z(n7490) );
  NANDN U13864 ( .A(init), .B(e[208]), .Z(n10585) );
  AND U13865 ( .A(n10586), .B(n10587), .Z(n10584) );
  NAND U13866 ( .A(ereg[207]), .B(n9759), .Z(n10587) );
  NANDN U13867 ( .A(n9754), .B(ereg[208]), .Z(n10586) );
  NAND U13868 ( .A(n10588), .B(n10589), .Z(n7489) );
  NANDN U13869 ( .A(init), .B(e[209]), .Z(n10589) );
  AND U13870 ( .A(n10590), .B(n10591), .Z(n10588) );
  NAND U13871 ( .A(ereg[208]), .B(n9759), .Z(n10591) );
  NANDN U13872 ( .A(n9754), .B(ereg[209]), .Z(n10590) );
  NAND U13873 ( .A(n10592), .B(n10593), .Z(n7488) );
  NANDN U13874 ( .A(init), .B(e[210]), .Z(n10593) );
  AND U13875 ( .A(n10594), .B(n10595), .Z(n10592) );
  NAND U13876 ( .A(ereg[209]), .B(n9759), .Z(n10595) );
  NANDN U13877 ( .A(n9754), .B(ereg[210]), .Z(n10594) );
  NAND U13878 ( .A(n10596), .B(n10597), .Z(n7487) );
  NANDN U13879 ( .A(init), .B(e[211]), .Z(n10597) );
  AND U13880 ( .A(n10598), .B(n10599), .Z(n10596) );
  NAND U13881 ( .A(ereg[210]), .B(n9759), .Z(n10599) );
  NANDN U13882 ( .A(n9754), .B(ereg[211]), .Z(n10598) );
  NAND U13883 ( .A(n10600), .B(n10601), .Z(n7486) );
  NANDN U13884 ( .A(init), .B(e[212]), .Z(n10601) );
  AND U13885 ( .A(n10602), .B(n10603), .Z(n10600) );
  NAND U13886 ( .A(ereg[211]), .B(n9759), .Z(n10603) );
  NANDN U13887 ( .A(n9754), .B(ereg[212]), .Z(n10602) );
  NAND U13888 ( .A(n10604), .B(n10605), .Z(n7485) );
  NANDN U13889 ( .A(init), .B(e[213]), .Z(n10605) );
  AND U13890 ( .A(n10606), .B(n10607), .Z(n10604) );
  NAND U13891 ( .A(ereg[212]), .B(n9759), .Z(n10607) );
  NANDN U13892 ( .A(n9754), .B(ereg[213]), .Z(n10606) );
  NAND U13893 ( .A(n10608), .B(n10609), .Z(n7484) );
  NANDN U13894 ( .A(init), .B(e[214]), .Z(n10609) );
  AND U13895 ( .A(n10610), .B(n10611), .Z(n10608) );
  NAND U13896 ( .A(ereg[213]), .B(n9759), .Z(n10611) );
  NANDN U13897 ( .A(n9754), .B(ereg[214]), .Z(n10610) );
  NAND U13898 ( .A(n10612), .B(n10613), .Z(n7483) );
  NANDN U13899 ( .A(init), .B(e[215]), .Z(n10613) );
  AND U13900 ( .A(n10614), .B(n10615), .Z(n10612) );
  NAND U13901 ( .A(ereg[214]), .B(n9759), .Z(n10615) );
  NANDN U13902 ( .A(n9754), .B(ereg[215]), .Z(n10614) );
  NAND U13903 ( .A(n10616), .B(n10617), .Z(n7482) );
  NANDN U13904 ( .A(init), .B(e[216]), .Z(n10617) );
  AND U13905 ( .A(n10618), .B(n10619), .Z(n10616) );
  NAND U13906 ( .A(ereg[215]), .B(n9759), .Z(n10619) );
  NANDN U13907 ( .A(n9754), .B(ereg[216]), .Z(n10618) );
  NAND U13908 ( .A(n10620), .B(n10621), .Z(n7481) );
  NANDN U13909 ( .A(init), .B(e[217]), .Z(n10621) );
  AND U13910 ( .A(n10622), .B(n10623), .Z(n10620) );
  NAND U13911 ( .A(ereg[216]), .B(n9759), .Z(n10623) );
  NANDN U13912 ( .A(n9754), .B(ereg[217]), .Z(n10622) );
  NAND U13913 ( .A(n10624), .B(n10625), .Z(n7480) );
  NANDN U13914 ( .A(init), .B(e[218]), .Z(n10625) );
  AND U13915 ( .A(n10626), .B(n10627), .Z(n10624) );
  NAND U13916 ( .A(ereg[217]), .B(n9759), .Z(n10627) );
  NANDN U13917 ( .A(n9754), .B(ereg[218]), .Z(n10626) );
  NAND U13918 ( .A(n10628), .B(n10629), .Z(n7479) );
  NANDN U13919 ( .A(init), .B(e[219]), .Z(n10629) );
  AND U13920 ( .A(n10630), .B(n10631), .Z(n10628) );
  NAND U13921 ( .A(ereg[218]), .B(n9759), .Z(n10631) );
  NANDN U13922 ( .A(n9754), .B(ereg[219]), .Z(n10630) );
  NAND U13923 ( .A(n10632), .B(n10633), .Z(n7478) );
  NANDN U13924 ( .A(init), .B(e[220]), .Z(n10633) );
  AND U13925 ( .A(n10634), .B(n10635), .Z(n10632) );
  NAND U13926 ( .A(ereg[219]), .B(n9759), .Z(n10635) );
  NANDN U13927 ( .A(n9754), .B(ereg[220]), .Z(n10634) );
  NAND U13928 ( .A(n10636), .B(n10637), .Z(n7477) );
  NANDN U13929 ( .A(init), .B(e[221]), .Z(n10637) );
  AND U13930 ( .A(n10638), .B(n10639), .Z(n10636) );
  NAND U13931 ( .A(ereg[220]), .B(n9759), .Z(n10639) );
  NANDN U13932 ( .A(n9754), .B(ereg[221]), .Z(n10638) );
  NAND U13933 ( .A(n10640), .B(n10641), .Z(n7476) );
  NANDN U13934 ( .A(init), .B(e[222]), .Z(n10641) );
  AND U13935 ( .A(n10642), .B(n10643), .Z(n10640) );
  NAND U13936 ( .A(ereg[221]), .B(n9759), .Z(n10643) );
  NANDN U13937 ( .A(n9754), .B(ereg[222]), .Z(n10642) );
  NAND U13938 ( .A(n10644), .B(n10645), .Z(n7475) );
  NANDN U13939 ( .A(init), .B(e[223]), .Z(n10645) );
  AND U13940 ( .A(n10646), .B(n10647), .Z(n10644) );
  NAND U13941 ( .A(ereg[222]), .B(n9759), .Z(n10647) );
  NANDN U13942 ( .A(n9754), .B(ereg[223]), .Z(n10646) );
  NAND U13943 ( .A(n10648), .B(n10649), .Z(n7474) );
  NANDN U13944 ( .A(init), .B(e[224]), .Z(n10649) );
  AND U13945 ( .A(n10650), .B(n10651), .Z(n10648) );
  NAND U13946 ( .A(ereg[223]), .B(n9759), .Z(n10651) );
  NANDN U13947 ( .A(n9754), .B(ereg[224]), .Z(n10650) );
  NAND U13948 ( .A(n10652), .B(n10653), .Z(n7473) );
  NANDN U13949 ( .A(init), .B(e[225]), .Z(n10653) );
  AND U13950 ( .A(n10654), .B(n10655), .Z(n10652) );
  NAND U13951 ( .A(ereg[224]), .B(n9759), .Z(n10655) );
  NANDN U13952 ( .A(n9754), .B(ereg[225]), .Z(n10654) );
  NAND U13953 ( .A(n10656), .B(n10657), .Z(n7472) );
  NANDN U13954 ( .A(init), .B(e[226]), .Z(n10657) );
  AND U13955 ( .A(n10658), .B(n10659), .Z(n10656) );
  NAND U13956 ( .A(ereg[225]), .B(n9759), .Z(n10659) );
  NANDN U13957 ( .A(n9754), .B(ereg[226]), .Z(n10658) );
  NAND U13958 ( .A(n10660), .B(n10661), .Z(n7471) );
  NANDN U13959 ( .A(init), .B(e[227]), .Z(n10661) );
  AND U13960 ( .A(n10662), .B(n10663), .Z(n10660) );
  NAND U13961 ( .A(ereg[226]), .B(n9759), .Z(n10663) );
  NANDN U13962 ( .A(n9754), .B(ereg[227]), .Z(n10662) );
  NAND U13963 ( .A(n10664), .B(n10665), .Z(n7470) );
  NANDN U13964 ( .A(init), .B(e[228]), .Z(n10665) );
  AND U13965 ( .A(n10666), .B(n10667), .Z(n10664) );
  NAND U13966 ( .A(ereg[227]), .B(n9759), .Z(n10667) );
  NANDN U13967 ( .A(n9754), .B(ereg[228]), .Z(n10666) );
  NAND U13968 ( .A(n10668), .B(n10669), .Z(n7469) );
  NANDN U13969 ( .A(init), .B(e[229]), .Z(n10669) );
  AND U13970 ( .A(n10670), .B(n10671), .Z(n10668) );
  NAND U13971 ( .A(ereg[228]), .B(n9759), .Z(n10671) );
  NANDN U13972 ( .A(n9754), .B(ereg[229]), .Z(n10670) );
  NAND U13973 ( .A(n10672), .B(n10673), .Z(n7468) );
  NANDN U13974 ( .A(init), .B(e[230]), .Z(n10673) );
  AND U13975 ( .A(n10674), .B(n10675), .Z(n10672) );
  NAND U13976 ( .A(ereg[229]), .B(n9759), .Z(n10675) );
  NANDN U13977 ( .A(n9754), .B(ereg[230]), .Z(n10674) );
  NAND U13978 ( .A(n10676), .B(n10677), .Z(n7467) );
  NANDN U13979 ( .A(init), .B(e[231]), .Z(n10677) );
  AND U13980 ( .A(n10678), .B(n10679), .Z(n10676) );
  NAND U13981 ( .A(ereg[230]), .B(n9759), .Z(n10679) );
  NANDN U13982 ( .A(n9754), .B(ereg[231]), .Z(n10678) );
  NAND U13983 ( .A(n10680), .B(n10681), .Z(n7466) );
  NANDN U13984 ( .A(init), .B(e[232]), .Z(n10681) );
  AND U13985 ( .A(n10682), .B(n10683), .Z(n10680) );
  NAND U13986 ( .A(ereg[231]), .B(n9759), .Z(n10683) );
  NANDN U13987 ( .A(n9754), .B(ereg[232]), .Z(n10682) );
  NAND U13988 ( .A(n10684), .B(n10685), .Z(n7465) );
  NANDN U13989 ( .A(init), .B(e[233]), .Z(n10685) );
  AND U13990 ( .A(n10686), .B(n10687), .Z(n10684) );
  NAND U13991 ( .A(ereg[232]), .B(n9759), .Z(n10687) );
  NANDN U13992 ( .A(n9754), .B(ereg[233]), .Z(n10686) );
  NAND U13993 ( .A(n10688), .B(n10689), .Z(n7464) );
  NANDN U13994 ( .A(init), .B(e[234]), .Z(n10689) );
  AND U13995 ( .A(n10690), .B(n10691), .Z(n10688) );
  NAND U13996 ( .A(ereg[233]), .B(n9759), .Z(n10691) );
  NANDN U13997 ( .A(n9754), .B(ereg[234]), .Z(n10690) );
  NAND U13998 ( .A(n10692), .B(n10693), .Z(n7463) );
  NANDN U13999 ( .A(init), .B(e[235]), .Z(n10693) );
  AND U14000 ( .A(n10694), .B(n10695), .Z(n10692) );
  NAND U14001 ( .A(ereg[234]), .B(n9759), .Z(n10695) );
  NANDN U14002 ( .A(n9754), .B(ereg[235]), .Z(n10694) );
  NAND U14003 ( .A(n10696), .B(n10697), .Z(n7462) );
  NANDN U14004 ( .A(init), .B(e[236]), .Z(n10697) );
  AND U14005 ( .A(n10698), .B(n10699), .Z(n10696) );
  NAND U14006 ( .A(ereg[235]), .B(n9759), .Z(n10699) );
  NANDN U14007 ( .A(n9754), .B(ereg[236]), .Z(n10698) );
  NAND U14008 ( .A(n10700), .B(n10701), .Z(n7461) );
  NANDN U14009 ( .A(init), .B(e[237]), .Z(n10701) );
  AND U14010 ( .A(n10702), .B(n10703), .Z(n10700) );
  NAND U14011 ( .A(ereg[236]), .B(n9759), .Z(n10703) );
  NANDN U14012 ( .A(n9754), .B(ereg[237]), .Z(n10702) );
  NAND U14013 ( .A(n10704), .B(n10705), .Z(n7460) );
  NANDN U14014 ( .A(init), .B(e[238]), .Z(n10705) );
  AND U14015 ( .A(n10706), .B(n10707), .Z(n10704) );
  NAND U14016 ( .A(ereg[237]), .B(n9759), .Z(n10707) );
  NANDN U14017 ( .A(n9754), .B(ereg[238]), .Z(n10706) );
  NAND U14018 ( .A(n10708), .B(n10709), .Z(n7459) );
  NANDN U14019 ( .A(init), .B(e[239]), .Z(n10709) );
  AND U14020 ( .A(n10710), .B(n10711), .Z(n10708) );
  NAND U14021 ( .A(ereg[238]), .B(n9759), .Z(n10711) );
  NANDN U14022 ( .A(n9754), .B(ereg[239]), .Z(n10710) );
  NAND U14023 ( .A(n10712), .B(n10713), .Z(n7458) );
  NANDN U14024 ( .A(init), .B(e[240]), .Z(n10713) );
  AND U14025 ( .A(n10714), .B(n10715), .Z(n10712) );
  NAND U14026 ( .A(ereg[239]), .B(n9759), .Z(n10715) );
  NANDN U14027 ( .A(n9754), .B(ereg[240]), .Z(n10714) );
  NAND U14028 ( .A(n10716), .B(n10717), .Z(n7457) );
  NANDN U14029 ( .A(init), .B(e[241]), .Z(n10717) );
  AND U14030 ( .A(n10718), .B(n10719), .Z(n10716) );
  NAND U14031 ( .A(ereg[240]), .B(n9759), .Z(n10719) );
  NANDN U14032 ( .A(n9754), .B(ereg[241]), .Z(n10718) );
  NAND U14033 ( .A(n10720), .B(n10721), .Z(n7456) );
  NANDN U14034 ( .A(init), .B(e[242]), .Z(n10721) );
  AND U14035 ( .A(n10722), .B(n10723), .Z(n10720) );
  NAND U14036 ( .A(ereg[241]), .B(n9759), .Z(n10723) );
  NANDN U14037 ( .A(n9754), .B(ereg[242]), .Z(n10722) );
  NAND U14038 ( .A(n10724), .B(n10725), .Z(n7455) );
  NANDN U14039 ( .A(init), .B(e[243]), .Z(n10725) );
  AND U14040 ( .A(n10726), .B(n10727), .Z(n10724) );
  NAND U14041 ( .A(ereg[242]), .B(n9759), .Z(n10727) );
  NANDN U14042 ( .A(n9754), .B(ereg[243]), .Z(n10726) );
  NAND U14043 ( .A(n10728), .B(n10729), .Z(n7454) );
  NANDN U14044 ( .A(init), .B(e[244]), .Z(n10729) );
  AND U14045 ( .A(n10730), .B(n10731), .Z(n10728) );
  NAND U14046 ( .A(ereg[243]), .B(n9759), .Z(n10731) );
  NANDN U14047 ( .A(n9754), .B(ereg[244]), .Z(n10730) );
  NAND U14048 ( .A(n10732), .B(n10733), .Z(n7453) );
  NANDN U14049 ( .A(init), .B(e[245]), .Z(n10733) );
  AND U14050 ( .A(n10734), .B(n10735), .Z(n10732) );
  NAND U14051 ( .A(ereg[244]), .B(n9759), .Z(n10735) );
  NANDN U14052 ( .A(n9754), .B(ereg[245]), .Z(n10734) );
  NAND U14053 ( .A(n10736), .B(n10737), .Z(n7452) );
  NANDN U14054 ( .A(init), .B(e[246]), .Z(n10737) );
  AND U14055 ( .A(n10738), .B(n10739), .Z(n10736) );
  NAND U14056 ( .A(ereg[245]), .B(n9759), .Z(n10739) );
  NANDN U14057 ( .A(n9754), .B(ereg[246]), .Z(n10738) );
  NAND U14058 ( .A(n10740), .B(n10741), .Z(n7451) );
  NANDN U14059 ( .A(init), .B(e[247]), .Z(n10741) );
  AND U14060 ( .A(n10742), .B(n10743), .Z(n10740) );
  NAND U14061 ( .A(ereg[246]), .B(n9759), .Z(n10743) );
  NANDN U14062 ( .A(n9754), .B(ereg[247]), .Z(n10742) );
  NAND U14063 ( .A(n10744), .B(n10745), .Z(n7450) );
  NANDN U14064 ( .A(init), .B(e[248]), .Z(n10745) );
  AND U14065 ( .A(n10746), .B(n10747), .Z(n10744) );
  NAND U14066 ( .A(ereg[247]), .B(n9759), .Z(n10747) );
  NANDN U14067 ( .A(n9754), .B(ereg[248]), .Z(n10746) );
  NAND U14068 ( .A(n10748), .B(n10749), .Z(n7449) );
  NANDN U14069 ( .A(init), .B(e[249]), .Z(n10749) );
  AND U14070 ( .A(n10750), .B(n10751), .Z(n10748) );
  NAND U14071 ( .A(ereg[248]), .B(n9759), .Z(n10751) );
  NANDN U14072 ( .A(n9754), .B(ereg[249]), .Z(n10750) );
  NAND U14073 ( .A(n10752), .B(n10753), .Z(n7448) );
  NANDN U14074 ( .A(init), .B(e[250]), .Z(n10753) );
  AND U14075 ( .A(n10754), .B(n10755), .Z(n10752) );
  NAND U14076 ( .A(ereg[249]), .B(n9759), .Z(n10755) );
  NANDN U14077 ( .A(n9754), .B(ereg[250]), .Z(n10754) );
  NAND U14078 ( .A(n10756), .B(n10757), .Z(n7447) );
  NANDN U14079 ( .A(init), .B(e[251]), .Z(n10757) );
  AND U14080 ( .A(n10758), .B(n10759), .Z(n10756) );
  NAND U14081 ( .A(ereg[250]), .B(n9759), .Z(n10759) );
  NANDN U14082 ( .A(n9754), .B(ereg[251]), .Z(n10758) );
  NAND U14083 ( .A(n10760), .B(n10761), .Z(n7446) );
  NANDN U14084 ( .A(init), .B(e[252]), .Z(n10761) );
  AND U14085 ( .A(n10762), .B(n10763), .Z(n10760) );
  NAND U14086 ( .A(ereg[251]), .B(n9759), .Z(n10763) );
  NANDN U14087 ( .A(n9754), .B(ereg[252]), .Z(n10762) );
  NAND U14088 ( .A(n10764), .B(n10765), .Z(n7445) );
  NANDN U14089 ( .A(init), .B(e[253]), .Z(n10765) );
  AND U14090 ( .A(n10766), .B(n10767), .Z(n10764) );
  NAND U14091 ( .A(ereg[252]), .B(n9759), .Z(n10767) );
  NANDN U14092 ( .A(n9754), .B(ereg[253]), .Z(n10766) );
  NAND U14093 ( .A(n10768), .B(n10769), .Z(n7444) );
  NANDN U14094 ( .A(init), .B(e[254]), .Z(n10769) );
  AND U14095 ( .A(n10770), .B(n10771), .Z(n10768) );
  NAND U14096 ( .A(ereg[253]), .B(n9759), .Z(n10771) );
  NANDN U14097 ( .A(n9754), .B(ereg[254]), .Z(n10770) );
  NAND U14098 ( .A(n10772), .B(n10773), .Z(n7443) );
  NANDN U14099 ( .A(init), .B(e[255]), .Z(n10773) );
  AND U14100 ( .A(n10774), .B(n10775), .Z(n10772) );
  NAND U14101 ( .A(ereg[254]), .B(n9759), .Z(n10775) );
  NANDN U14102 ( .A(n9754), .B(ereg[255]), .Z(n10774) );
  NAND U14103 ( .A(n10776), .B(n10777), .Z(n7442) );
  NANDN U14104 ( .A(init), .B(e[256]), .Z(n10777) );
  AND U14105 ( .A(n10778), .B(n10779), .Z(n10776) );
  NAND U14106 ( .A(ereg[255]), .B(n9759), .Z(n10779) );
  NANDN U14107 ( .A(n9754), .B(ereg[256]), .Z(n10778) );
  NAND U14108 ( .A(n10780), .B(n10781), .Z(n7441) );
  NANDN U14109 ( .A(init), .B(e[257]), .Z(n10781) );
  AND U14110 ( .A(n10782), .B(n10783), .Z(n10780) );
  NAND U14111 ( .A(ereg[256]), .B(n9759), .Z(n10783) );
  NANDN U14112 ( .A(n9754), .B(ereg[257]), .Z(n10782) );
  NAND U14113 ( .A(n10784), .B(n10785), .Z(n7440) );
  NANDN U14114 ( .A(init), .B(e[258]), .Z(n10785) );
  AND U14115 ( .A(n10786), .B(n10787), .Z(n10784) );
  NAND U14116 ( .A(ereg[257]), .B(n9759), .Z(n10787) );
  NANDN U14117 ( .A(n9754), .B(ereg[258]), .Z(n10786) );
  NAND U14118 ( .A(n10788), .B(n10789), .Z(n7439) );
  NANDN U14119 ( .A(init), .B(e[259]), .Z(n10789) );
  AND U14120 ( .A(n10790), .B(n10791), .Z(n10788) );
  NAND U14121 ( .A(ereg[258]), .B(n9759), .Z(n10791) );
  NANDN U14122 ( .A(n9754), .B(ereg[259]), .Z(n10790) );
  NAND U14123 ( .A(n10792), .B(n10793), .Z(n7438) );
  NANDN U14124 ( .A(init), .B(e[260]), .Z(n10793) );
  AND U14125 ( .A(n10794), .B(n10795), .Z(n10792) );
  NAND U14126 ( .A(ereg[259]), .B(n9759), .Z(n10795) );
  NANDN U14127 ( .A(n9754), .B(ereg[260]), .Z(n10794) );
  NAND U14128 ( .A(n10796), .B(n10797), .Z(n7437) );
  NANDN U14129 ( .A(init), .B(e[261]), .Z(n10797) );
  AND U14130 ( .A(n10798), .B(n10799), .Z(n10796) );
  NAND U14131 ( .A(ereg[260]), .B(n9759), .Z(n10799) );
  NANDN U14132 ( .A(n9754), .B(ereg[261]), .Z(n10798) );
  NAND U14133 ( .A(n10800), .B(n10801), .Z(n7436) );
  NANDN U14134 ( .A(init), .B(e[262]), .Z(n10801) );
  AND U14135 ( .A(n10802), .B(n10803), .Z(n10800) );
  NAND U14136 ( .A(ereg[261]), .B(n9759), .Z(n10803) );
  NANDN U14137 ( .A(n9754), .B(ereg[262]), .Z(n10802) );
  NAND U14138 ( .A(n10804), .B(n10805), .Z(n7435) );
  NANDN U14139 ( .A(init), .B(e[263]), .Z(n10805) );
  AND U14140 ( .A(n10806), .B(n10807), .Z(n10804) );
  NAND U14141 ( .A(ereg[262]), .B(n9759), .Z(n10807) );
  NANDN U14142 ( .A(n9754), .B(ereg[263]), .Z(n10806) );
  NAND U14143 ( .A(n10808), .B(n10809), .Z(n7434) );
  NANDN U14144 ( .A(init), .B(e[264]), .Z(n10809) );
  AND U14145 ( .A(n10810), .B(n10811), .Z(n10808) );
  NAND U14146 ( .A(ereg[263]), .B(n9759), .Z(n10811) );
  NANDN U14147 ( .A(n9754), .B(ereg[264]), .Z(n10810) );
  NAND U14148 ( .A(n10812), .B(n10813), .Z(n7433) );
  NANDN U14149 ( .A(init), .B(e[265]), .Z(n10813) );
  AND U14150 ( .A(n10814), .B(n10815), .Z(n10812) );
  NAND U14151 ( .A(ereg[264]), .B(n9759), .Z(n10815) );
  NANDN U14152 ( .A(n9754), .B(ereg[265]), .Z(n10814) );
  NAND U14153 ( .A(n10816), .B(n10817), .Z(n7432) );
  NANDN U14154 ( .A(init), .B(e[266]), .Z(n10817) );
  AND U14155 ( .A(n10818), .B(n10819), .Z(n10816) );
  NAND U14156 ( .A(ereg[265]), .B(n9759), .Z(n10819) );
  NANDN U14157 ( .A(n9754), .B(ereg[266]), .Z(n10818) );
  NAND U14158 ( .A(n10820), .B(n10821), .Z(n7431) );
  NANDN U14159 ( .A(init), .B(e[267]), .Z(n10821) );
  AND U14160 ( .A(n10822), .B(n10823), .Z(n10820) );
  NAND U14161 ( .A(ereg[266]), .B(n9759), .Z(n10823) );
  NANDN U14162 ( .A(n9754), .B(ereg[267]), .Z(n10822) );
  NAND U14163 ( .A(n10824), .B(n10825), .Z(n7430) );
  NANDN U14164 ( .A(init), .B(e[268]), .Z(n10825) );
  AND U14165 ( .A(n10826), .B(n10827), .Z(n10824) );
  NAND U14166 ( .A(ereg[267]), .B(n9759), .Z(n10827) );
  NANDN U14167 ( .A(n9754), .B(ereg[268]), .Z(n10826) );
  NAND U14168 ( .A(n10828), .B(n10829), .Z(n7429) );
  NANDN U14169 ( .A(init), .B(e[269]), .Z(n10829) );
  AND U14170 ( .A(n10830), .B(n10831), .Z(n10828) );
  NAND U14171 ( .A(ereg[268]), .B(n9759), .Z(n10831) );
  NANDN U14172 ( .A(n9754), .B(ereg[269]), .Z(n10830) );
  NAND U14173 ( .A(n10832), .B(n10833), .Z(n7428) );
  NANDN U14174 ( .A(init), .B(e[270]), .Z(n10833) );
  AND U14175 ( .A(n10834), .B(n10835), .Z(n10832) );
  NAND U14176 ( .A(ereg[269]), .B(n9759), .Z(n10835) );
  NANDN U14177 ( .A(n9754), .B(ereg[270]), .Z(n10834) );
  NAND U14178 ( .A(n10836), .B(n10837), .Z(n7427) );
  NANDN U14179 ( .A(init), .B(e[271]), .Z(n10837) );
  AND U14180 ( .A(n10838), .B(n10839), .Z(n10836) );
  NAND U14181 ( .A(ereg[270]), .B(n9759), .Z(n10839) );
  NANDN U14182 ( .A(n9754), .B(ereg[271]), .Z(n10838) );
  NAND U14183 ( .A(n10840), .B(n10841), .Z(n7426) );
  NANDN U14184 ( .A(init), .B(e[272]), .Z(n10841) );
  AND U14185 ( .A(n10842), .B(n10843), .Z(n10840) );
  NAND U14186 ( .A(ereg[271]), .B(n9759), .Z(n10843) );
  NANDN U14187 ( .A(n9754), .B(ereg[272]), .Z(n10842) );
  NAND U14188 ( .A(n10844), .B(n10845), .Z(n7425) );
  NANDN U14189 ( .A(init), .B(e[273]), .Z(n10845) );
  AND U14190 ( .A(n10846), .B(n10847), .Z(n10844) );
  NAND U14191 ( .A(ereg[272]), .B(n9759), .Z(n10847) );
  NANDN U14192 ( .A(n9754), .B(ereg[273]), .Z(n10846) );
  NAND U14193 ( .A(n10848), .B(n10849), .Z(n7424) );
  NANDN U14194 ( .A(init), .B(e[274]), .Z(n10849) );
  AND U14195 ( .A(n10850), .B(n10851), .Z(n10848) );
  NAND U14196 ( .A(ereg[273]), .B(n9759), .Z(n10851) );
  NANDN U14197 ( .A(n9754), .B(ereg[274]), .Z(n10850) );
  NAND U14198 ( .A(n10852), .B(n10853), .Z(n7423) );
  NANDN U14199 ( .A(init), .B(e[275]), .Z(n10853) );
  AND U14200 ( .A(n10854), .B(n10855), .Z(n10852) );
  NAND U14201 ( .A(ereg[274]), .B(n9759), .Z(n10855) );
  NANDN U14202 ( .A(n9754), .B(ereg[275]), .Z(n10854) );
  NAND U14203 ( .A(n10856), .B(n10857), .Z(n7422) );
  NANDN U14204 ( .A(init), .B(e[276]), .Z(n10857) );
  AND U14205 ( .A(n10858), .B(n10859), .Z(n10856) );
  NAND U14206 ( .A(ereg[275]), .B(n9759), .Z(n10859) );
  NANDN U14207 ( .A(n9754), .B(ereg[276]), .Z(n10858) );
  NAND U14208 ( .A(n10860), .B(n10861), .Z(n7421) );
  NANDN U14209 ( .A(init), .B(e[277]), .Z(n10861) );
  AND U14210 ( .A(n10862), .B(n10863), .Z(n10860) );
  NAND U14211 ( .A(ereg[276]), .B(n9759), .Z(n10863) );
  NANDN U14212 ( .A(n9754), .B(ereg[277]), .Z(n10862) );
  NAND U14213 ( .A(n10864), .B(n10865), .Z(n7420) );
  NANDN U14214 ( .A(init), .B(e[278]), .Z(n10865) );
  AND U14215 ( .A(n10866), .B(n10867), .Z(n10864) );
  NAND U14216 ( .A(ereg[277]), .B(n9759), .Z(n10867) );
  NANDN U14217 ( .A(n9754), .B(ereg[278]), .Z(n10866) );
  NAND U14218 ( .A(n10868), .B(n10869), .Z(n7419) );
  NANDN U14219 ( .A(init), .B(e[279]), .Z(n10869) );
  AND U14220 ( .A(n10870), .B(n10871), .Z(n10868) );
  NAND U14221 ( .A(ereg[278]), .B(n9759), .Z(n10871) );
  NANDN U14222 ( .A(n9754), .B(ereg[279]), .Z(n10870) );
  NAND U14223 ( .A(n10872), .B(n10873), .Z(n7418) );
  NANDN U14224 ( .A(init), .B(e[280]), .Z(n10873) );
  AND U14225 ( .A(n10874), .B(n10875), .Z(n10872) );
  NAND U14226 ( .A(ereg[279]), .B(n9759), .Z(n10875) );
  NANDN U14227 ( .A(n9754), .B(ereg[280]), .Z(n10874) );
  NAND U14228 ( .A(n10876), .B(n10877), .Z(n7417) );
  NANDN U14229 ( .A(init), .B(e[281]), .Z(n10877) );
  AND U14230 ( .A(n10878), .B(n10879), .Z(n10876) );
  NAND U14231 ( .A(ereg[280]), .B(n9759), .Z(n10879) );
  NANDN U14232 ( .A(n9754), .B(ereg[281]), .Z(n10878) );
  NAND U14233 ( .A(n10880), .B(n10881), .Z(n7416) );
  NANDN U14234 ( .A(init), .B(e[282]), .Z(n10881) );
  AND U14235 ( .A(n10882), .B(n10883), .Z(n10880) );
  NAND U14236 ( .A(ereg[281]), .B(n9759), .Z(n10883) );
  NANDN U14237 ( .A(n9754), .B(ereg[282]), .Z(n10882) );
  NAND U14238 ( .A(n10884), .B(n10885), .Z(n7415) );
  NANDN U14239 ( .A(init), .B(e[283]), .Z(n10885) );
  AND U14240 ( .A(n10886), .B(n10887), .Z(n10884) );
  NAND U14241 ( .A(ereg[282]), .B(n9759), .Z(n10887) );
  NANDN U14242 ( .A(n9754), .B(ereg[283]), .Z(n10886) );
  NAND U14243 ( .A(n10888), .B(n10889), .Z(n7414) );
  NANDN U14244 ( .A(init), .B(e[284]), .Z(n10889) );
  AND U14245 ( .A(n10890), .B(n10891), .Z(n10888) );
  NAND U14246 ( .A(ereg[283]), .B(n9759), .Z(n10891) );
  NANDN U14247 ( .A(n9754), .B(ereg[284]), .Z(n10890) );
  NAND U14248 ( .A(n10892), .B(n10893), .Z(n7413) );
  NANDN U14249 ( .A(init), .B(e[285]), .Z(n10893) );
  AND U14250 ( .A(n10894), .B(n10895), .Z(n10892) );
  NAND U14251 ( .A(ereg[284]), .B(n9759), .Z(n10895) );
  NANDN U14252 ( .A(n9754), .B(ereg[285]), .Z(n10894) );
  NAND U14253 ( .A(n10896), .B(n10897), .Z(n7412) );
  NANDN U14254 ( .A(init), .B(e[286]), .Z(n10897) );
  AND U14255 ( .A(n10898), .B(n10899), .Z(n10896) );
  NAND U14256 ( .A(ereg[285]), .B(n9759), .Z(n10899) );
  NANDN U14257 ( .A(n9754), .B(ereg[286]), .Z(n10898) );
  NAND U14258 ( .A(n10900), .B(n10901), .Z(n7411) );
  NANDN U14259 ( .A(init), .B(e[287]), .Z(n10901) );
  AND U14260 ( .A(n10902), .B(n10903), .Z(n10900) );
  NAND U14261 ( .A(ereg[286]), .B(n9759), .Z(n10903) );
  NANDN U14262 ( .A(n9754), .B(ereg[287]), .Z(n10902) );
  NAND U14263 ( .A(n10904), .B(n10905), .Z(n7410) );
  NANDN U14264 ( .A(init), .B(e[288]), .Z(n10905) );
  AND U14265 ( .A(n10906), .B(n10907), .Z(n10904) );
  NAND U14266 ( .A(ereg[287]), .B(n9759), .Z(n10907) );
  NANDN U14267 ( .A(n9754), .B(ereg[288]), .Z(n10906) );
  NAND U14268 ( .A(n10908), .B(n10909), .Z(n7409) );
  NANDN U14269 ( .A(init), .B(e[289]), .Z(n10909) );
  AND U14270 ( .A(n10910), .B(n10911), .Z(n10908) );
  NAND U14271 ( .A(ereg[288]), .B(n9759), .Z(n10911) );
  NANDN U14272 ( .A(n9754), .B(ereg[289]), .Z(n10910) );
  NAND U14273 ( .A(n10912), .B(n10913), .Z(n7408) );
  NANDN U14274 ( .A(init), .B(e[290]), .Z(n10913) );
  AND U14275 ( .A(n10914), .B(n10915), .Z(n10912) );
  NAND U14276 ( .A(ereg[289]), .B(n9759), .Z(n10915) );
  NANDN U14277 ( .A(n9754), .B(ereg[290]), .Z(n10914) );
  NAND U14278 ( .A(n10916), .B(n10917), .Z(n7407) );
  NANDN U14279 ( .A(init), .B(e[291]), .Z(n10917) );
  AND U14280 ( .A(n10918), .B(n10919), .Z(n10916) );
  NAND U14281 ( .A(ereg[290]), .B(n9759), .Z(n10919) );
  NANDN U14282 ( .A(n9754), .B(ereg[291]), .Z(n10918) );
  NAND U14283 ( .A(n10920), .B(n10921), .Z(n7406) );
  NANDN U14284 ( .A(init), .B(e[292]), .Z(n10921) );
  AND U14285 ( .A(n10922), .B(n10923), .Z(n10920) );
  NAND U14286 ( .A(ereg[291]), .B(n9759), .Z(n10923) );
  NANDN U14287 ( .A(n9754), .B(ereg[292]), .Z(n10922) );
  NAND U14288 ( .A(n10924), .B(n10925), .Z(n7405) );
  NANDN U14289 ( .A(init), .B(e[293]), .Z(n10925) );
  AND U14290 ( .A(n10926), .B(n10927), .Z(n10924) );
  NAND U14291 ( .A(ereg[292]), .B(n9759), .Z(n10927) );
  NANDN U14292 ( .A(n9754), .B(ereg[293]), .Z(n10926) );
  NAND U14293 ( .A(n10928), .B(n10929), .Z(n7404) );
  NANDN U14294 ( .A(init), .B(e[294]), .Z(n10929) );
  AND U14295 ( .A(n10930), .B(n10931), .Z(n10928) );
  NAND U14296 ( .A(ereg[293]), .B(n9759), .Z(n10931) );
  NANDN U14297 ( .A(n9754), .B(ereg[294]), .Z(n10930) );
  NAND U14298 ( .A(n10932), .B(n10933), .Z(n7403) );
  NANDN U14299 ( .A(init), .B(e[295]), .Z(n10933) );
  AND U14300 ( .A(n10934), .B(n10935), .Z(n10932) );
  NAND U14301 ( .A(ereg[294]), .B(n9759), .Z(n10935) );
  NANDN U14302 ( .A(n9754), .B(ereg[295]), .Z(n10934) );
  NAND U14303 ( .A(n10936), .B(n10937), .Z(n7402) );
  NANDN U14304 ( .A(init), .B(e[296]), .Z(n10937) );
  AND U14305 ( .A(n10938), .B(n10939), .Z(n10936) );
  NAND U14306 ( .A(ereg[295]), .B(n9759), .Z(n10939) );
  NANDN U14307 ( .A(n9754), .B(ereg[296]), .Z(n10938) );
  NAND U14308 ( .A(n10940), .B(n10941), .Z(n7401) );
  NANDN U14309 ( .A(init), .B(e[297]), .Z(n10941) );
  AND U14310 ( .A(n10942), .B(n10943), .Z(n10940) );
  NAND U14311 ( .A(ereg[296]), .B(n9759), .Z(n10943) );
  NANDN U14312 ( .A(n9754), .B(ereg[297]), .Z(n10942) );
  NAND U14313 ( .A(n10944), .B(n10945), .Z(n7400) );
  NANDN U14314 ( .A(init), .B(e[298]), .Z(n10945) );
  AND U14315 ( .A(n10946), .B(n10947), .Z(n10944) );
  NAND U14316 ( .A(ereg[297]), .B(n9759), .Z(n10947) );
  NANDN U14317 ( .A(n9754), .B(ereg[298]), .Z(n10946) );
  NAND U14318 ( .A(n10948), .B(n10949), .Z(n7399) );
  NANDN U14319 ( .A(init), .B(e[299]), .Z(n10949) );
  AND U14320 ( .A(n10950), .B(n10951), .Z(n10948) );
  NAND U14321 ( .A(ereg[298]), .B(n9759), .Z(n10951) );
  NANDN U14322 ( .A(n9754), .B(ereg[299]), .Z(n10950) );
  NAND U14323 ( .A(n10952), .B(n10953), .Z(n7398) );
  NANDN U14324 ( .A(init), .B(e[300]), .Z(n10953) );
  AND U14325 ( .A(n10954), .B(n10955), .Z(n10952) );
  NAND U14326 ( .A(ereg[299]), .B(n9759), .Z(n10955) );
  NANDN U14327 ( .A(n9754), .B(ereg[300]), .Z(n10954) );
  NAND U14328 ( .A(n10956), .B(n10957), .Z(n7397) );
  NANDN U14329 ( .A(init), .B(e[301]), .Z(n10957) );
  AND U14330 ( .A(n10958), .B(n10959), .Z(n10956) );
  NAND U14331 ( .A(ereg[300]), .B(n9759), .Z(n10959) );
  NANDN U14332 ( .A(n9754), .B(ereg[301]), .Z(n10958) );
  NAND U14333 ( .A(n10960), .B(n10961), .Z(n7396) );
  NANDN U14334 ( .A(init), .B(e[302]), .Z(n10961) );
  AND U14335 ( .A(n10962), .B(n10963), .Z(n10960) );
  NAND U14336 ( .A(ereg[301]), .B(n9759), .Z(n10963) );
  NANDN U14337 ( .A(n9754), .B(ereg[302]), .Z(n10962) );
  NAND U14338 ( .A(n10964), .B(n10965), .Z(n7395) );
  NANDN U14339 ( .A(init), .B(e[303]), .Z(n10965) );
  AND U14340 ( .A(n10966), .B(n10967), .Z(n10964) );
  NAND U14341 ( .A(ereg[302]), .B(n9759), .Z(n10967) );
  NANDN U14342 ( .A(n9754), .B(ereg[303]), .Z(n10966) );
  NAND U14343 ( .A(n10968), .B(n10969), .Z(n7394) );
  NANDN U14344 ( .A(init), .B(e[304]), .Z(n10969) );
  AND U14345 ( .A(n10970), .B(n10971), .Z(n10968) );
  NAND U14346 ( .A(ereg[303]), .B(n9759), .Z(n10971) );
  NANDN U14347 ( .A(n9754), .B(ereg[304]), .Z(n10970) );
  NAND U14348 ( .A(n10972), .B(n10973), .Z(n7393) );
  NANDN U14349 ( .A(init), .B(e[305]), .Z(n10973) );
  AND U14350 ( .A(n10974), .B(n10975), .Z(n10972) );
  NAND U14351 ( .A(ereg[304]), .B(n9759), .Z(n10975) );
  NANDN U14352 ( .A(n9754), .B(ereg[305]), .Z(n10974) );
  NAND U14353 ( .A(n10976), .B(n10977), .Z(n7392) );
  NANDN U14354 ( .A(init), .B(e[306]), .Z(n10977) );
  AND U14355 ( .A(n10978), .B(n10979), .Z(n10976) );
  NAND U14356 ( .A(ereg[305]), .B(n9759), .Z(n10979) );
  NANDN U14357 ( .A(n9754), .B(ereg[306]), .Z(n10978) );
  NAND U14358 ( .A(n10980), .B(n10981), .Z(n7391) );
  NANDN U14359 ( .A(init), .B(e[307]), .Z(n10981) );
  AND U14360 ( .A(n10982), .B(n10983), .Z(n10980) );
  NAND U14361 ( .A(ereg[306]), .B(n9759), .Z(n10983) );
  NANDN U14362 ( .A(n9754), .B(ereg[307]), .Z(n10982) );
  NAND U14363 ( .A(n10984), .B(n10985), .Z(n7390) );
  NANDN U14364 ( .A(init), .B(e[308]), .Z(n10985) );
  AND U14365 ( .A(n10986), .B(n10987), .Z(n10984) );
  NAND U14366 ( .A(ereg[307]), .B(n9759), .Z(n10987) );
  NANDN U14367 ( .A(n9754), .B(ereg[308]), .Z(n10986) );
  NAND U14368 ( .A(n10988), .B(n10989), .Z(n7389) );
  NANDN U14369 ( .A(init), .B(e[309]), .Z(n10989) );
  AND U14370 ( .A(n10990), .B(n10991), .Z(n10988) );
  NAND U14371 ( .A(ereg[308]), .B(n9759), .Z(n10991) );
  NANDN U14372 ( .A(n9754), .B(ereg[309]), .Z(n10990) );
  NAND U14373 ( .A(n10992), .B(n10993), .Z(n7388) );
  NANDN U14374 ( .A(init), .B(e[310]), .Z(n10993) );
  AND U14375 ( .A(n10994), .B(n10995), .Z(n10992) );
  NAND U14376 ( .A(ereg[309]), .B(n9759), .Z(n10995) );
  NANDN U14377 ( .A(n9754), .B(ereg[310]), .Z(n10994) );
  NAND U14378 ( .A(n10996), .B(n10997), .Z(n7387) );
  NANDN U14379 ( .A(init), .B(e[311]), .Z(n10997) );
  AND U14380 ( .A(n10998), .B(n10999), .Z(n10996) );
  NAND U14381 ( .A(ereg[310]), .B(n9759), .Z(n10999) );
  NANDN U14382 ( .A(n9754), .B(ereg[311]), .Z(n10998) );
  NAND U14383 ( .A(n11000), .B(n11001), .Z(n7386) );
  NANDN U14384 ( .A(init), .B(e[312]), .Z(n11001) );
  AND U14385 ( .A(n11002), .B(n11003), .Z(n11000) );
  NAND U14386 ( .A(ereg[311]), .B(n9759), .Z(n11003) );
  NANDN U14387 ( .A(n9754), .B(ereg[312]), .Z(n11002) );
  NAND U14388 ( .A(n11004), .B(n11005), .Z(n7385) );
  NANDN U14389 ( .A(init), .B(e[313]), .Z(n11005) );
  AND U14390 ( .A(n11006), .B(n11007), .Z(n11004) );
  NAND U14391 ( .A(ereg[312]), .B(n9759), .Z(n11007) );
  NANDN U14392 ( .A(n9754), .B(ereg[313]), .Z(n11006) );
  NAND U14393 ( .A(n11008), .B(n11009), .Z(n7384) );
  NANDN U14394 ( .A(init), .B(e[314]), .Z(n11009) );
  AND U14395 ( .A(n11010), .B(n11011), .Z(n11008) );
  NAND U14396 ( .A(ereg[313]), .B(n9759), .Z(n11011) );
  NANDN U14397 ( .A(n9754), .B(ereg[314]), .Z(n11010) );
  NAND U14398 ( .A(n11012), .B(n11013), .Z(n7383) );
  NANDN U14399 ( .A(init), .B(e[315]), .Z(n11013) );
  AND U14400 ( .A(n11014), .B(n11015), .Z(n11012) );
  NAND U14401 ( .A(ereg[314]), .B(n9759), .Z(n11015) );
  NANDN U14402 ( .A(n9754), .B(ereg[315]), .Z(n11014) );
  NAND U14403 ( .A(n11016), .B(n11017), .Z(n7382) );
  NANDN U14404 ( .A(init), .B(e[316]), .Z(n11017) );
  AND U14405 ( .A(n11018), .B(n11019), .Z(n11016) );
  NAND U14406 ( .A(ereg[315]), .B(n9759), .Z(n11019) );
  NANDN U14407 ( .A(n9754), .B(ereg[316]), .Z(n11018) );
  NAND U14408 ( .A(n11020), .B(n11021), .Z(n7381) );
  NANDN U14409 ( .A(init), .B(e[317]), .Z(n11021) );
  AND U14410 ( .A(n11022), .B(n11023), .Z(n11020) );
  NAND U14411 ( .A(ereg[316]), .B(n9759), .Z(n11023) );
  NANDN U14412 ( .A(n9754), .B(ereg[317]), .Z(n11022) );
  NAND U14413 ( .A(n11024), .B(n11025), .Z(n7380) );
  NANDN U14414 ( .A(init), .B(e[318]), .Z(n11025) );
  AND U14415 ( .A(n11026), .B(n11027), .Z(n11024) );
  NAND U14416 ( .A(ereg[317]), .B(n9759), .Z(n11027) );
  NANDN U14417 ( .A(n9754), .B(ereg[318]), .Z(n11026) );
  NAND U14418 ( .A(n11028), .B(n11029), .Z(n7379) );
  NANDN U14419 ( .A(init), .B(e[319]), .Z(n11029) );
  AND U14420 ( .A(n11030), .B(n11031), .Z(n11028) );
  NAND U14421 ( .A(ereg[318]), .B(n9759), .Z(n11031) );
  NANDN U14422 ( .A(n9754), .B(ereg[319]), .Z(n11030) );
  NAND U14423 ( .A(n11032), .B(n11033), .Z(n7378) );
  NANDN U14424 ( .A(init), .B(e[320]), .Z(n11033) );
  AND U14425 ( .A(n11034), .B(n11035), .Z(n11032) );
  NAND U14426 ( .A(ereg[319]), .B(n9759), .Z(n11035) );
  NANDN U14427 ( .A(n9754), .B(ereg[320]), .Z(n11034) );
  NAND U14428 ( .A(n11036), .B(n11037), .Z(n7377) );
  NANDN U14429 ( .A(init), .B(e[321]), .Z(n11037) );
  AND U14430 ( .A(n11038), .B(n11039), .Z(n11036) );
  NAND U14431 ( .A(ereg[320]), .B(n9759), .Z(n11039) );
  NANDN U14432 ( .A(n9754), .B(ereg[321]), .Z(n11038) );
  NAND U14433 ( .A(n11040), .B(n11041), .Z(n7376) );
  NANDN U14434 ( .A(init), .B(e[322]), .Z(n11041) );
  AND U14435 ( .A(n11042), .B(n11043), .Z(n11040) );
  NAND U14436 ( .A(ereg[321]), .B(n9759), .Z(n11043) );
  NANDN U14437 ( .A(n9754), .B(ereg[322]), .Z(n11042) );
  NAND U14438 ( .A(n11044), .B(n11045), .Z(n7375) );
  NANDN U14439 ( .A(init), .B(e[323]), .Z(n11045) );
  AND U14440 ( .A(n11046), .B(n11047), .Z(n11044) );
  NAND U14441 ( .A(ereg[322]), .B(n9759), .Z(n11047) );
  NANDN U14442 ( .A(n9754), .B(ereg[323]), .Z(n11046) );
  NAND U14443 ( .A(n11048), .B(n11049), .Z(n7374) );
  NANDN U14444 ( .A(init), .B(e[324]), .Z(n11049) );
  AND U14445 ( .A(n11050), .B(n11051), .Z(n11048) );
  NAND U14446 ( .A(ereg[323]), .B(n9759), .Z(n11051) );
  NANDN U14447 ( .A(n9754), .B(ereg[324]), .Z(n11050) );
  NAND U14448 ( .A(n11052), .B(n11053), .Z(n7373) );
  NANDN U14449 ( .A(init), .B(e[325]), .Z(n11053) );
  AND U14450 ( .A(n11054), .B(n11055), .Z(n11052) );
  NAND U14451 ( .A(ereg[324]), .B(n9759), .Z(n11055) );
  NANDN U14452 ( .A(n9754), .B(ereg[325]), .Z(n11054) );
  NAND U14453 ( .A(n11056), .B(n11057), .Z(n7372) );
  NANDN U14454 ( .A(init), .B(e[326]), .Z(n11057) );
  AND U14455 ( .A(n11058), .B(n11059), .Z(n11056) );
  NAND U14456 ( .A(ereg[325]), .B(n9759), .Z(n11059) );
  NANDN U14457 ( .A(n9754), .B(ereg[326]), .Z(n11058) );
  NAND U14458 ( .A(n11060), .B(n11061), .Z(n7371) );
  NANDN U14459 ( .A(init), .B(e[327]), .Z(n11061) );
  AND U14460 ( .A(n11062), .B(n11063), .Z(n11060) );
  NAND U14461 ( .A(ereg[326]), .B(n9759), .Z(n11063) );
  NANDN U14462 ( .A(n9754), .B(ereg[327]), .Z(n11062) );
  NAND U14463 ( .A(n11064), .B(n11065), .Z(n7370) );
  NANDN U14464 ( .A(init), .B(e[328]), .Z(n11065) );
  AND U14465 ( .A(n11066), .B(n11067), .Z(n11064) );
  NAND U14466 ( .A(ereg[327]), .B(n9759), .Z(n11067) );
  NANDN U14467 ( .A(n9754), .B(ereg[328]), .Z(n11066) );
  NAND U14468 ( .A(n11068), .B(n11069), .Z(n7369) );
  NANDN U14469 ( .A(init), .B(e[329]), .Z(n11069) );
  AND U14470 ( .A(n11070), .B(n11071), .Z(n11068) );
  NAND U14471 ( .A(ereg[328]), .B(n9759), .Z(n11071) );
  NANDN U14472 ( .A(n9754), .B(ereg[329]), .Z(n11070) );
  NAND U14473 ( .A(n11072), .B(n11073), .Z(n7368) );
  NANDN U14474 ( .A(init), .B(e[330]), .Z(n11073) );
  AND U14475 ( .A(n11074), .B(n11075), .Z(n11072) );
  NAND U14476 ( .A(ereg[329]), .B(n9759), .Z(n11075) );
  NANDN U14477 ( .A(n9754), .B(ereg[330]), .Z(n11074) );
  NAND U14478 ( .A(n11076), .B(n11077), .Z(n7367) );
  NANDN U14479 ( .A(init), .B(e[331]), .Z(n11077) );
  AND U14480 ( .A(n11078), .B(n11079), .Z(n11076) );
  NAND U14481 ( .A(ereg[330]), .B(n9759), .Z(n11079) );
  NANDN U14482 ( .A(n9754), .B(ereg[331]), .Z(n11078) );
  NAND U14483 ( .A(n11080), .B(n11081), .Z(n7366) );
  NANDN U14484 ( .A(init), .B(e[332]), .Z(n11081) );
  AND U14485 ( .A(n11082), .B(n11083), .Z(n11080) );
  NAND U14486 ( .A(ereg[331]), .B(n9759), .Z(n11083) );
  NANDN U14487 ( .A(n9754), .B(ereg[332]), .Z(n11082) );
  NAND U14488 ( .A(n11084), .B(n11085), .Z(n7365) );
  NANDN U14489 ( .A(init), .B(e[333]), .Z(n11085) );
  AND U14490 ( .A(n11086), .B(n11087), .Z(n11084) );
  NAND U14491 ( .A(ereg[332]), .B(n9759), .Z(n11087) );
  NANDN U14492 ( .A(n9754), .B(ereg[333]), .Z(n11086) );
  NAND U14493 ( .A(n11088), .B(n11089), .Z(n7364) );
  NANDN U14494 ( .A(init), .B(e[334]), .Z(n11089) );
  AND U14495 ( .A(n11090), .B(n11091), .Z(n11088) );
  NAND U14496 ( .A(ereg[333]), .B(n9759), .Z(n11091) );
  NANDN U14497 ( .A(n9754), .B(ereg[334]), .Z(n11090) );
  NAND U14498 ( .A(n11092), .B(n11093), .Z(n7363) );
  NANDN U14499 ( .A(init), .B(e[335]), .Z(n11093) );
  AND U14500 ( .A(n11094), .B(n11095), .Z(n11092) );
  NAND U14501 ( .A(ereg[334]), .B(n9759), .Z(n11095) );
  NANDN U14502 ( .A(n9754), .B(ereg[335]), .Z(n11094) );
  NAND U14503 ( .A(n11096), .B(n11097), .Z(n7362) );
  NANDN U14504 ( .A(init), .B(e[336]), .Z(n11097) );
  AND U14505 ( .A(n11098), .B(n11099), .Z(n11096) );
  NAND U14506 ( .A(ereg[335]), .B(n9759), .Z(n11099) );
  NANDN U14507 ( .A(n9754), .B(ereg[336]), .Z(n11098) );
  NAND U14508 ( .A(n11100), .B(n11101), .Z(n7361) );
  NANDN U14509 ( .A(init), .B(e[337]), .Z(n11101) );
  AND U14510 ( .A(n11102), .B(n11103), .Z(n11100) );
  NAND U14511 ( .A(ereg[336]), .B(n9759), .Z(n11103) );
  NANDN U14512 ( .A(n9754), .B(ereg[337]), .Z(n11102) );
  NAND U14513 ( .A(n11104), .B(n11105), .Z(n7360) );
  NANDN U14514 ( .A(init), .B(e[338]), .Z(n11105) );
  AND U14515 ( .A(n11106), .B(n11107), .Z(n11104) );
  NAND U14516 ( .A(ereg[337]), .B(n9759), .Z(n11107) );
  NANDN U14517 ( .A(n9754), .B(ereg[338]), .Z(n11106) );
  NAND U14518 ( .A(n11108), .B(n11109), .Z(n7359) );
  NANDN U14519 ( .A(init), .B(e[339]), .Z(n11109) );
  AND U14520 ( .A(n11110), .B(n11111), .Z(n11108) );
  NAND U14521 ( .A(ereg[338]), .B(n9759), .Z(n11111) );
  NANDN U14522 ( .A(n9754), .B(ereg[339]), .Z(n11110) );
  NAND U14523 ( .A(n11112), .B(n11113), .Z(n7358) );
  NANDN U14524 ( .A(init), .B(e[340]), .Z(n11113) );
  AND U14525 ( .A(n11114), .B(n11115), .Z(n11112) );
  NAND U14526 ( .A(ereg[339]), .B(n9759), .Z(n11115) );
  NANDN U14527 ( .A(n9754), .B(ereg[340]), .Z(n11114) );
  NAND U14528 ( .A(n11116), .B(n11117), .Z(n7357) );
  NANDN U14529 ( .A(init), .B(e[341]), .Z(n11117) );
  AND U14530 ( .A(n11118), .B(n11119), .Z(n11116) );
  NAND U14531 ( .A(ereg[340]), .B(n9759), .Z(n11119) );
  NANDN U14532 ( .A(n9754), .B(ereg[341]), .Z(n11118) );
  NAND U14533 ( .A(n11120), .B(n11121), .Z(n7356) );
  NANDN U14534 ( .A(init), .B(e[342]), .Z(n11121) );
  AND U14535 ( .A(n11122), .B(n11123), .Z(n11120) );
  NAND U14536 ( .A(ereg[341]), .B(n9759), .Z(n11123) );
  NANDN U14537 ( .A(n9754), .B(ereg[342]), .Z(n11122) );
  NAND U14538 ( .A(n11124), .B(n11125), .Z(n7355) );
  NANDN U14539 ( .A(init), .B(e[343]), .Z(n11125) );
  AND U14540 ( .A(n11126), .B(n11127), .Z(n11124) );
  NAND U14541 ( .A(ereg[342]), .B(n9759), .Z(n11127) );
  NANDN U14542 ( .A(n9754), .B(ereg[343]), .Z(n11126) );
  NAND U14543 ( .A(n11128), .B(n11129), .Z(n7354) );
  NANDN U14544 ( .A(init), .B(e[344]), .Z(n11129) );
  AND U14545 ( .A(n11130), .B(n11131), .Z(n11128) );
  NAND U14546 ( .A(ereg[343]), .B(n9759), .Z(n11131) );
  NANDN U14547 ( .A(n9754), .B(ereg[344]), .Z(n11130) );
  NAND U14548 ( .A(n11132), .B(n11133), .Z(n7353) );
  NANDN U14549 ( .A(init), .B(e[345]), .Z(n11133) );
  AND U14550 ( .A(n11134), .B(n11135), .Z(n11132) );
  NAND U14551 ( .A(ereg[344]), .B(n9759), .Z(n11135) );
  NANDN U14552 ( .A(n9754), .B(ereg[345]), .Z(n11134) );
  NAND U14553 ( .A(n11136), .B(n11137), .Z(n7352) );
  NANDN U14554 ( .A(init), .B(e[346]), .Z(n11137) );
  AND U14555 ( .A(n11138), .B(n11139), .Z(n11136) );
  NAND U14556 ( .A(ereg[345]), .B(n9759), .Z(n11139) );
  NANDN U14557 ( .A(n9754), .B(ereg[346]), .Z(n11138) );
  NAND U14558 ( .A(n11140), .B(n11141), .Z(n7351) );
  NANDN U14559 ( .A(init), .B(e[347]), .Z(n11141) );
  AND U14560 ( .A(n11142), .B(n11143), .Z(n11140) );
  NAND U14561 ( .A(ereg[346]), .B(n9759), .Z(n11143) );
  NANDN U14562 ( .A(n9754), .B(ereg[347]), .Z(n11142) );
  NAND U14563 ( .A(n11144), .B(n11145), .Z(n7350) );
  NANDN U14564 ( .A(init), .B(e[348]), .Z(n11145) );
  AND U14565 ( .A(n11146), .B(n11147), .Z(n11144) );
  NAND U14566 ( .A(ereg[347]), .B(n9759), .Z(n11147) );
  NANDN U14567 ( .A(n9754), .B(ereg[348]), .Z(n11146) );
  NAND U14568 ( .A(n11148), .B(n11149), .Z(n7349) );
  NANDN U14569 ( .A(init), .B(e[349]), .Z(n11149) );
  AND U14570 ( .A(n11150), .B(n11151), .Z(n11148) );
  NAND U14571 ( .A(ereg[348]), .B(n9759), .Z(n11151) );
  NANDN U14572 ( .A(n9754), .B(ereg[349]), .Z(n11150) );
  NAND U14573 ( .A(n11152), .B(n11153), .Z(n7348) );
  NANDN U14574 ( .A(init), .B(e[350]), .Z(n11153) );
  AND U14575 ( .A(n11154), .B(n11155), .Z(n11152) );
  NAND U14576 ( .A(ereg[349]), .B(n9759), .Z(n11155) );
  NANDN U14577 ( .A(n9754), .B(ereg[350]), .Z(n11154) );
  NAND U14578 ( .A(n11156), .B(n11157), .Z(n7347) );
  NANDN U14579 ( .A(init), .B(e[351]), .Z(n11157) );
  AND U14580 ( .A(n11158), .B(n11159), .Z(n11156) );
  NAND U14581 ( .A(ereg[350]), .B(n9759), .Z(n11159) );
  NANDN U14582 ( .A(n9754), .B(ereg[351]), .Z(n11158) );
  NAND U14583 ( .A(n11160), .B(n11161), .Z(n7346) );
  NANDN U14584 ( .A(init), .B(e[352]), .Z(n11161) );
  AND U14585 ( .A(n11162), .B(n11163), .Z(n11160) );
  NAND U14586 ( .A(ereg[351]), .B(n9759), .Z(n11163) );
  NANDN U14587 ( .A(n9754), .B(ereg[352]), .Z(n11162) );
  NAND U14588 ( .A(n11164), .B(n11165), .Z(n7345) );
  NANDN U14589 ( .A(init), .B(e[353]), .Z(n11165) );
  AND U14590 ( .A(n11166), .B(n11167), .Z(n11164) );
  NAND U14591 ( .A(ereg[352]), .B(n9759), .Z(n11167) );
  NANDN U14592 ( .A(n9754), .B(ereg[353]), .Z(n11166) );
  NAND U14593 ( .A(n11168), .B(n11169), .Z(n7344) );
  NANDN U14594 ( .A(init), .B(e[354]), .Z(n11169) );
  AND U14595 ( .A(n11170), .B(n11171), .Z(n11168) );
  NAND U14596 ( .A(ereg[353]), .B(n9759), .Z(n11171) );
  NANDN U14597 ( .A(n9754), .B(ereg[354]), .Z(n11170) );
  NAND U14598 ( .A(n11172), .B(n11173), .Z(n7343) );
  NANDN U14599 ( .A(init), .B(e[355]), .Z(n11173) );
  AND U14600 ( .A(n11174), .B(n11175), .Z(n11172) );
  NAND U14601 ( .A(ereg[354]), .B(n9759), .Z(n11175) );
  NANDN U14602 ( .A(n9754), .B(ereg[355]), .Z(n11174) );
  NAND U14603 ( .A(n11176), .B(n11177), .Z(n7342) );
  NANDN U14604 ( .A(init), .B(e[356]), .Z(n11177) );
  AND U14605 ( .A(n11178), .B(n11179), .Z(n11176) );
  NAND U14606 ( .A(ereg[355]), .B(n9759), .Z(n11179) );
  NANDN U14607 ( .A(n9754), .B(ereg[356]), .Z(n11178) );
  NAND U14608 ( .A(n11180), .B(n11181), .Z(n7341) );
  NANDN U14609 ( .A(init), .B(e[357]), .Z(n11181) );
  AND U14610 ( .A(n11182), .B(n11183), .Z(n11180) );
  NAND U14611 ( .A(ereg[356]), .B(n9759), .Z(n11183) );
  NANDN U14612 ( .A(n9754), .B(ereg[357]), .Z(n11182) );
  NAND U14613 ( .A(n11184), .B(n11185), .Z(n7340) );
  NANDN U14614 ( .A(init), .B(e[358]), .Z(n11185) );
  AND U14615 ( .A(n11186), .B(n11187), .Z(n11184) );
  NAND U14616 ( .A(ereg[357]), .B(n9759), .Z(n11187) );
  NANDN U14617 ( .A(n9754), .B(ereg[358]), .Z(n11186) );
  NAND U14618 ( .A(n11188), .B(n11189), .Z(n7339) );
  NANDN U14619 ( .A(init), .B(e[359]), .Z(n11189) );
  AND U14620 ( .A(n11190), .B(n11191), .Z(n11188) );
  NAND U14621 ( .A(ereg[358]), .B(n9759), .Z(n11191) );
  NANDN U14622 ( .A(n9754), .B(ereg[359]), .Z(n11190) );
  NAND U14623 ( .A(n11192), .B(n11193), .Z(n7338) );
  NANDN U14624 ( .A(init), .B(e[360]), .Z(n11193) );
  AND U14625 ( .A(n11194), .B(n11195), .Z(n11192) );
  NAND U14626 ( .A(ereg[359]), .B(n9759), .Z(n11195) );
  NANDN U14627 ( .A(n9754), .B(ereg[360]), .Z(n11194) );
  NAND U14628 ( .A(n11196), .B(n11197), .Z(n7337) );
  NANDN U14629 ( .A(init), .B(e[361]), .Z(n11197) );
  AND U14630 ( .A(n11198), .B(n11199), .Z(n11196) );
  NAND U14631 ( .A(ereg[360]), .B(n9759), .Z(n11199) );
  NANDN U14632 ( .A(n9754), .B(ereg[361]), .Z(n11198) );
  NAND U14633 ( .A(n11200), .B(n11201), .Z(n7336) );
  NANDN U14634 ( .A(init), .B(e[362]), .Z(n11201) );
  AND U14635 ( .A(n11202), .B(n11203), .Z(n11200) );
  NAND U14636 ( .A(ereg[361]), .B(n9759), .Z(n11203) );
  NANDN U14637 ( .A(n9754), .B(ereg[362]), .Z(n11202) );
  NAND U14638 ( .A(n11204), .B(n11205), .Z(n7335) );
  NANDN U14639 ( .A(init), .B(e[363]), .Z(n11205) );
  AND U14640 ( .A(n11206), .B(n11207), .Z(n11204) );
  NAND U14641 ( .A(ereg[362]), .B(n9759), .Z(n11207) );
  NANDN U14642 ( .A(n9754), .B(ereg[363]), .Z(n11206) );
  NAND U14643 ( .A(n11208), .B(n11209), .Z(n7334) );
  NANDN U14644 ( .A(init), .B(e[364]), .Z(n11209) );
  AND U14645 ( .A(n11210), .B(n11211), .Z(n11208) );
  NAND U14646 ( .A(ereg[363]), .B(n9759), .Z(n11211) );
  NANDN U14647 ( .A(n9754), .B(ereg[364]), .Z(n11210) );
  NAND U14648 ( .A(n11212), .B(n11213), .Z(n7333) );
  NANDN U14649 ( .A(init), .B(e[365]), .Z(n11213) );
  AND U14650 ( .A(n11214), .B(n11215), .Z(n11212) );
  NAND U14651 ( .A(ereg[364]), .B(n9759), .Z(n11215) );
  NANDN U14652 ( .A(n9754), .B(ereg[365]), .Z(n11214) );
  NAND U14653 ( .A(n11216), .B(n11217), .Z(n7332) );
  NANDN U14654 ( .A(init), .B(e[366]), .Z(n11217) );
  AND U14655 ( .A(n11218), .B(n11219), .Z(n11216) );
  NAND U14656 ( .A(ereg[365]), .B(n9759), .Z(n11219) );
  NANDN U14657 ( .A(n9754), .B(ereg[366]), .Z(n11218) );
  NAND U14658 ( .A(n11220), .B(n11221), .Z(n7331) );
  NANDN U14659 ( .A(init), .B(e[367]), .Z(n11221) );
  AND U14660 ( .A(n11222), .B(n11223), .Z(n11220) );
  NAND U14661 ( .A(ereg[366]), .B(n9759), .Z(n11223) );
  NANDN U14662 ( .A(n9754), .B(ereg[367]), .Z(n11222) );
  NAND U14663 ( .A(n11224), .B(n11225), .Z(n7330) );
  NANDN U14664 ( .A(init), .B(e[368]), .Z(n11225) );
  AND U14665 ( .A(n11226), .B(n11227), .Z(n11224) );
  NAND U14666 ( .A(ereg[367]), .B(n9759), .Z(n11227) );
  NANDN U14667 ( .A(n9754), .B(ereg[368]), .Z(n11226) );
  NAND U14668 ( .A(n11228), .B(n11229), .Z(n7329) );
  NANDN U14669 ( .A(init), .B(e[369]), .Z(n11229) );
  AND U14670 ( .A(n11230), .B(n11231), .Z(n11228) );
  NAND U14671 ( .A(ereg[368]), .B(n9759), .Z(n11231) );
  NANDN U14672 ( .A(n9754), .B(ereg[369]), .Z(n11230) );
  NAND U14673 ( .A(n11232), .B(n11233), .Z(n7328) );
  NANDN U14674 ( .A(init), .B(e[370]), .Z(n11233) );
  AND U14675 ( .A(n11234), .B(n11235), .Z(n11232) );
  NAND U14676 ( .A(ereg[369]), .B(n9759), .Z(n11235) );
  NANDN U14677 ( .A(n9754), .B(ereg[370]), .Z(n11234) );
  NAND U14678 ( .A(n11236), .B(n11237), .Z(n7327) );
  NANDN U14679 ( .A(init), .B(e[371]), .Z(n11237) );
  AND U14680 ( .A(n11238), .B(n11239), .Z(n11236) );
  NAND U14681 ( .A(ereg[370]), .B(n9759), .Z(n11239) );
  NANDN U14682 ( .A(n9754), .B(ereg[371]), .Z(n11238) );
  NAND U14683 ( .A(n11240), .B(n11241), .Z(n7326) );
  NANDN U14684 ( .A(init), .B(e[372]), .Z(n11241) );
  AND U14685 ( .A(n11242), .B(n11243), .Z(n11240) );
  NAND U14686 ( .A(ereg[371]), .B(n9759), .Z(n11243) );
  NANDN U14687 ( .A(n9754), .B(ereg[372]), .Z(n11242) );
  NAND U14688 ( .A(n11244), .B(n11245), .Z(n7325) );
  NANDN U14689 ( .A(init), .B(e[373]), .Z(n11245) );
  AND U14690 ( .A(n11246), .B(n11247), .Z(n11244) );
  NAND U14691 ( .A(ereg[372]), .B(n9759), .Z(n11247) );
  NANDN U14692 ( .A(n9754), .B(ereg[373]), .Z(n11246) );
  NAND U14693 ( .A(n11248), .B(n11249), .Z(n7324) );
  NANDN U14694 ( .A(init), .B(e[374]), .Z(n11249) );
  AND U14695 ( .A(n11250), .B(n11251), .Z(n11248) );
  NAND U14696 ( .A(ereg[373]), .B(n9759), .Z(n11251) );
  NANDN U14697 ( .A(n9754), .B(ereg[374]), .Z(n11250) );
  NAND U14698 ( .A(n11252), .B(n11253), .Z(n7323) );
  NANDN U14699 ( .A(init), .B(e[375]), .Z(n11253) );
  AND U14700 ( .A(n11254), .B(n11255), .Z(n11252) );
  NAND U14701 ( .A(ereg[374]), .B(n9759), .Z(n11255) );
  NANDN U14702 ( .A(n9754), .B(ereg[375]), .Z(n11254) );
  NAND U14703 ( .A(n11256), .B(n11257), .Z(n7322) );
  NANDN U14704 ( .A(init), .B(e[376]), .Z(n11257) );
  AND U14705 ( .A(n11258), .B(n11259), .Z(n11256) );
  NAND U14706 ( .A(ereg[375]), .B(n9759), .Z(n11259) );
  NANDN U14707 ( .A(n9754), .B(ereg[376]), .Z(n11258) );
  NAND U14708 ( .A(n11260), .B(n11261), .Z(n7321) );
  NANDN U14709 ( .A(init), .B(e[377]), .Z(n11261) );
  AND U14710 ( .A(n11262), .B(n11263), .Z(n11260) );
  NAND U14711 ( .A(ereg[376]), .B(n9759), .Z(n11263) );
  NANDN U14712 ( .A(n9754), .B(ereg[377]), .Z(n11262) );
  NAND U14713 ( .A(n11264), .B(n11265), .Z(n7320) );
  NANDN U14714 ( .A(init), .B(e[378]), .Z(n11265) );
  AND U14715 ( .A(n11266), .B(n11267), .Z(n11264) );
  NAND U14716 ( .A(ereg[377]), .B(n9759), .Z(n11267) );
  NANDN U14717 ( .A(n9754), .B(ereg[378]), .Z(n11266) );
  NAND U14718 ( .A(n11268), .B(n11269), .Z(n7319) );
  NANDN U14719 ( .A(init), .B(e[379]), .Z(n11269) );
  AND U14720 ( .A(n11270), .B(n11271), .Z(n11268) );
  NAND U14721 ( .A(ereg[378]), .B(n9759), .Z(n11271) );
  NANDN U14722 ( .A(n9754), .B(ereg[379]), .Z(n11270) );
  NAND U14723 ( .A(n11272), .B(n11273), .Z(n7318) );
  NANDN U14724 ( .A(init), .B(e[380]), .Z(n11273) );
  AND U14725 ( .A(n11274), .B(n11275), .Z(n11272) );
  NAND U14726 ( .A(ereg[379]), .B(n9759), .Z(n11275) );
  NANDN U14727 ( .A(n9754), .B(ereg[380]), .Z(n11274) );
  NAND U14728 ( .A(n11276), .B(n11277), .Z(n7317) );
  NANDN U14729 ( .A(init), .B(e[381]), .Z(n11277) );
  AND U14730 ( .A(n11278), .B(n11279), .Z(n11276) );
  NAND U14731 ( .A(ereg[380]), .B(n9759), .Z(n11279) );
  NANDN U14732 ( .A(n9754), .B(ereg[381]), .Z(n11278) );
  NAND U14733 ( .A(n11280), .B(n11281), .Z(n7316) );
  NANDN U14734 ( .A(init), .B(e[382]), .Z(n11281) );
  AND U14735 ( .A(n11282), .B(n11283), .Z(n11280) );
  NAND U14736 ( .A(ereg[381]), .B(n9759), .Z(n11283) );
  NANDN U14737 ( .A(n9754), .B(ereg[382]), .Z(n11282) );
  NAND U14738 ( .A(n11284), .B(n11285), .Z(n7315) );
  NANDN U14739 ( .A(init), .B(e[383]), .Z(n11285) );
  AND U14740 ( .A(n11286), .B(n11287), .Z(n11284) );
  NAND U14741 ( .A(ereg[382]), .B(n9759), .Z(n11287) );
  NANDN U14742 ( .A(n9754), .B(ereg[383]), .Z(n11286) );
  NAND U14743 ( .A(n11288), .B(n11289), .Z(n7314) );
  NANDN U14744 ( .A(init), .B(e[384]), .Z(n11289) );
  AND U14745 ( .A(n11290), .B(n11291), .Z(n11288) );
  NAND U14746 ( .A(ereg[383]), .B(n9759), .Z(n11291) );
  NANDN U14747 ( .A(n9754), .B(ereg[384]), .Z(n11290) );
  NAND U14748 ( .A(n11292), .B(n11293), .Z(n7313) );
  NANDN U14749 ( .A(init), .B(e[385]), .Z(n11293) );
  AND U14750 ( .A(n11294), .B(n11295), .Z(n11292) );
  NAND U14751 ( .A(ereg[384]), .B(n9759), .Z(n11295) );
  NANDN U14752 ( .A(n9754), .B(ereg[385]), .Z(n11294) );
  NAND U14753 ( .A(n11296), .B(n11297), .Z(n7312) );
  NANDN U14754 ( .A(init), .B(e[386]), .Z(n11297) );
  AND U14755 ( .A(n11298), .B(n11299), .Z(n11296) );
  NAND U14756 ( .A(ereg[385]), .B(n9759), .Z(n11299) );
  NANDN U14757 ( .A(n9754), .B(ereg[386]), .Z(n11298) );
  NAND U14758 ( .A(n11300), .B(n11301), .Z(n7311) );
  NANDN U14759 ( .A(init), .B(e[387]), .Z(n11301) );
  AND U14760 ( .A(n11302), .B(n11303), .Z(n11300) );
  NAND U14761 ( .A(ereg[386]), .B(n9759), .Z(n11303) );
  NANDN U14762 ( .A(n9754), .B(ereg[387]), .Z(n11302) );
  NAND U14763 ( .A(n11304), .B(n11305), .Z(n7310) );
  NANDN U14764 ( .A(init), .B(e[388]), .Z(n11305) );
  AND U14765 ( .A(n11306), .B(n11307), .Z(n11304) );
  NAND U14766 ( .A(ereg[387]), .B(n9759), .Z(n11307) );
  NANDN U14767 ( .A(n9754), .B(ereg[388]), .Z(n11306) );
  NAND U14768 ( .A(n11308), .B(n11309), .Z(n7309) );
  NANDN U14769 ( .A(init), .B(e[389]), .Z(n11309) );
  AND U14770 ( .A(n11310), .B(n11311), .Z(n11308) );
  NAND U14771 ( .A(ereg[388]), .B(n9759), .Z(n11311) );
  NANDN U14772 ( .A(n9754), .B(ereg[389]), .Z(n11310) );
  NAND U14773 ( .A(n11312), .B(n11313), .Z(n7308) );
  NANDN U14774 ( .A(init), .B(e[390]), .Z(n11313) );
  AND U14775 ( .A(n11314), .B(n11315), .Z(n11312) );
  NAND U14776 ( .A(ereg[389]), .B(n9759), .Z(n11315) );
  NANDN U14777 ( .A(n9754), .B(ereg[390]), .Z(n11314) );
  NAND U14778 ( .A(n11316), .B(n11317), .Z(n7307) );
  NANDN U14779 ( .A(init), .B(e[391]), .Z(n11317) );
  AND U14780 ( .A(n11318), .B(n11319), .Z(n11316) );
  NAND U14781 ( .A(ereg[390]), .B(n9759), .Z(n11319) );
  NANDN U14782 ( .A(n9754), .B(ereg[391]), .Z(n11318) );
  NAND U14783 ( .A(n11320), .B(n11321), .Z(n7306) );
  NANDN U14784 ( .A(init), .B(e[392]), .Z(n11321) );
  AND U14785 ( .A(n11322), .B(n11323), .Z(n11320) );
  NAND U14786 ( .A(ereg[391]), .B(n9759), .Z(n11323) );
  NANDN U14787 ( .A(n9754), .B(ereg[392]), .Z(n11322) );
  NAND U14788 ( .A(n11324), .B(n11325), .Z(n7305) );
  NANDN U14789 ( .A(init), .B(e[393]), .Z(n11325) );
  AND U14790 ( .A(n11326), .B(n11327), .Z(n11324) );
  NAND U14791 ( .A(ereg[392]), .B(n9759), .Z(n11327) );
  NANDN U14792 ( .A(n9754), .B(ereg[393]), .Z(n11326) );
  NAND U14793 ( .A(n11328), .B(n11329), .Z(n7304) );
  NANDN U14794 ( .A(init), .B(e[394]), .Z(n11329) );
  AND U14795 ( .A(n11330), .B(n11331), .Z(n11328) );
  NAND U14796 ( .A(ereg[393]), .B(n9759), .Z(n11331) );
  NANDN U14797 ( .A(n9754), .B(ereg[394]), .Z(n11330) );
  NAND U14798 ( .A(n11332), .B(n11333), .Z(n7303) );
  NANDN U14799 ( .A(init), .B(e[395]), .Z(n11333) );
  AND U14800 ( .A(n11334), .B(n11335), .Z(n11332) );
  NAND U14801 ( .A(ereg[394]), .B(n9759), .Z(n11335) );
  NANDN U14802 ( .A(n9754), .B(ereg[395]), .Z(n11334) );
  NAND U14803 ( .A(n11336), .B(n11337), .Z(n7302) );
  NANDN U14804 ( .A(init), .B(e[396]), .Z(n11337) );
  AND U14805 ( .A(n11338), .B(n11339), .Z(n11336) );
  NAND U14806 ( .A(ereg[395]), .B(n9759), .Z(n11339) );
  NANDN U14807 ( .A(n9754), .B(ereg[396]), .Z(n11338) );
  NAND U14808 ( .A(n11340), .B(n11341), .Z(n7301) );
  NANDN U14809 ( .A(init), .B(e[397]), .Z(n11341) );
  AND U14810 ( .A(n11342), .B(n11343), .Z(n11340) );
  NAND U14811 ( .A(ereg[396]), .B(n9759), .Z(n11343) );
  NANDN U14812 ( .A(n9754), .B(ereg[397]), .Z(n11342) );
  NAND U14813 ( .A(n11344), .B(n11345), .Z(n7300) );
  NANDN U14814 ( .A(init), .B(e[398]), .Z(n11345) );
  AND U14815 ( .A(n11346), .B(n11347), .Z(n11344) );
  NAND U14816 ( .A(ereg[397]), .B(n9759), .Z(n11347) );
  NANDN U14817 ( .A(n9754), .B(ereg[398]), .Z(n11346) );
  NAND U14818 ( .A(n11348), .B(n11349), .Z(n7299) );
  NANDN U14819 ( .A(init), .B(e[399]), .Z(n11349) );
  AND U14820 ( .A(n11350), .B(n11351), .Z(n11348) );
  NAND U14821 ( .A(ereg[398]), .B(n9759), .Z(n11351) );
  NANDN U14822 ( .A(n9754), .B(ereg[399]), .Z(n11350) );
  NAND U14823 ( .A(n11352), .B(n11353), .Z(n7298) );
  NANDN U14824 ( .A(init), .B(e[400]), .Z(n11353) );
  AND U14825 ( .A(n11354), .B(n11355), .Z(n11352) );
  NAND U14826 ( .A(ereg[399]), .B(n9759), .Z(n11355) );
  NANDN U14827 ( .A(n9754), .B(ereg[400]), .Z(n11354) );
  NAND U14828 ( .A(n11356), .B(n11357), .Z(n7297) );
  NANDN U14829 ( .A(init), .B(e[401]), .Z(n11357) );
  AND U14830 ( .A(n11358), .B(n11359), .Z(n11356) );
  NAND U14831 ( .A(ereg[400]), .B(n9759), .Z(n11359) );
  NANDN U14832 ( .A(n9754), .B(ereg[401]), .Z(n11358) );
  NAND U14833 ( .A(n11360), .B(n11361), .Z(n7296) );
  NANDN U14834 ( .A(init), .B(e[402]), .Z(n11361) );
  AND U14835 ( .A(n11362), .B(n11363), .Z(n11360) );
  NAND U14836 ( .A(ereg[401]), .B(n9759), .Z(n11363) );
  NANDN U14837 ( .A(n9754), .B(ereg[402]), .Z(n11362) );
  NAND U14838 ( .A(n11364), .B(n11365), .Z(n7295) );
  NANDN U14839 ( .A(init), .B(e[403]), .Z(n11365) );
  AND U14840 ( .A(n11366), .B(n11367), .Z(n11364) );
  NAND U14841 ( .A(ereg[402]), .B(n9759), .Z(n11367) );
  NANDN U14842 ( .A(n9754), .B(ereg[403]), .Z(n11366) );
  NAND U14843 ( .A(n11368), .B(n11369), .Z(n7294) );
  NANDN U14844 ( .A(init), .B(e[404]), .Z(n11369) );
  AND U14845 ( .A(n11370), .B(n11371), .Z(n11368) );
  NAND U14846 ( .A(ereg[403]), .B(n9759), .Z(n11371) );
  NANDN U14847 ( .A(n9754), .B(ereg[404]), .Z(n11370) );
  NAND U14848 ( .A(n11372), .B(n11373), .Z(n7293) );
  NANDN U14849 ( .A(init), .B(e[405]), .Z(n11373) );
  AND U14850 ( .A(n11374), .B(n11375), .Z(n11372) );
  NAND U14851 ( .A(ereg[404]), .B(n9759), .Z(n11375) );
  NANDN U14852 ( .A(n9754), .B(ereg[405]), .Z(n11374) );
  NAND U14853 ( .A(n11376), .B(n11377), .Z(n7292) );
  NANDN U14854 ( .A(init), .B(e[406]), .Z(n11377) );
  AND U14855 ( .A(n11378), .B(n11379), .Z(n11376) );
  NAND U14856 ( .A(ereg[405]), .B(n9759), .Z(n11379) );
  NANDN U14857 ( .A(n9754), .B(ereg[406]), .Z(n11378) );
  NAND U14858 ( .A(n11380), .B(n11381), .Z(n7291) );
  NANDN U14859 ( .A(init), .B(e[407]), .Z(n11381) );
  AND U14860 ( .A(n11382), .B(n11383), .Z(n11380) );
  NAND U14861 ( .A(ereg[406]), .B(n9759), .Z(n11383) );
  NANDN U14862 ( .A(n9754), .B(ereg[407]), .Z(n11382) );
  NAND U14863 ( .A(n11384), .B(n11385), .Z(n7290) );
  NANDN U14864 ( .A(init), .B(e[408]), .Z(n11385) );
  AND U14865 ( .A(n11386), .B(n11387), .Z(n11384) );
  NAND U14866 ( .A(ereg[407]), .B(n9759), .Z(n11387) );
  NANDN U14867 ( .A(n9754), .B(ereg[408]), .Z(n11386) );
  NAND U14868 ( .A(n11388), .B(n11389), .Z(n7289) );
  NANDN U14869 ( .A(init), .B(e[409]), .Z(n11389) );
  AND U14870 ( .A(n11390), .B(n11391), .Z(n11388) );
  NAND U14871 ( .A(ereg[408]), .B(n9759), .Z(n11391) );
  NANDN U14872 ( .A(n9754), .B(ereg[409]), .Z(n11390) );
  NAND U14873 ( .A(n11392), .B(n11393), .Z(n7288) );
  NANDN U14874 ( .A(init), .B(e[410]), .Z(n11393) );
  AND U14875 ( .A(n11394), .B(n11395), .Z(n11392) );
  NAND U14876 ( .A(ereg[409]), .B(n9759), .Z(n11395) );
  NANDN U14877 ( .A(n9754), .B(ereg[410]), .Z(n11394) );
  NAND U14878 ( .A(n11396), .B(n11397), .Z(n7287) );
  NANDN U14879 ( .A(init), .B(e[411]), .Z(n11397) );
  AND U14880 ( .A(n11398), .B(n11399), .Z(n11396) );
  NAND U14881 ( .A(ereg[410]), .B(n9759), .Z(n11399) );
  NANDN U14882 ( .A(n9754), .B(ereg[411]), .Z(n11398) );
  NAND U14883 ( .A(n11400), .B(n11401), .Z(n7286) );
  NANDN U14884 ( .A(init), .B(e[412]), .Z(n11401) );
  AND U14885 ( .A(n11402), .B(n11403), .Z(n11400) );
  NAND U14886 ( .A(ereg[411]), .B(n9759), .Z(n11403) );
  NANDN U14887 ( .A(n9754), .B(ereg[412]), .Z(n11402) );
  NAND U14888 ( .A(n11404), .B(n11405), .Z(n7285) );
  NANDN U14889 ( .A(init), .B(e[413]), .Z(n11405) );
  AND U14890 ( .A(n11406), .B(n11407), .Z(n11404) );
  NAND U14891 ( .A(ereg[412]), .B(n9759), .Z(n11407) );
  NANDN U14892 ( .A(n9754), .B(ereg[413]), .Z(n11406) );
  NAND U14893 ( .A(n11408), .B(n11409), .Z(n7284) );
  NANDN U14894 ( .A(init), .B(e[414]), .Z(n11409) );
  AND U14895 ( .A(n11410), .B(n11411), .Z(n11408) );
  NAND U14896 ( .A(ereg[413]), .B(n9759), .Z(n11411) );
  NANDN U14897 ( .A(n9754), .B(ereg[414]), .Z(n11410) );
  NAND U14898 ( .A(n11412), .B(n11413), .Z(n7283) );
  NANDN U14899 ( .A(init), .B(e[415]), .Z(n11413) );
  AND U14900 ( .A(n11414), .B(n11415), .Z(n11412) );
  NAND U14901 ( .A(ereg[414]), .B(n9759), .Z(n11415) );
  NANDN U14902 ( .A(n9754), .B(ereg[415]), .Z(n11414) );
  NAND U14903 ( .A(n11416), .B(n11417), .Z(n7282) );
  NANDN U14904 ( .A(init), .B(e[416]), .Z(n11417) );
  AND U14905 ( .A(n11418), .B(n11419), .Z(n11416) );
  NAND U14906 ( .A(ereg[415]), .B(n9759), .Z(n11419) );
  NANDN U14907 ( .A(n9754), .B(ereg[416]), .Z(n11418) );
  NAND U14908 ( .A(n11420), .B(n11421), .Z(n7281) );
  NANDN U14909 ( .A(init), .B(e[417]), .Z(n11421) );
  AND U14910 ( .A(n11422), .B(n11423), .Z(n11420) );
  NAND U14911 ( .A(ereg[416]), .B(n9759), .Z(n11423) );
  NANDN U14912 ( .A(n9754), .B(ereg[417]), .Z(n11422) );
  NAND U14913 ( .A(n11424), .B(n11425), .Z(n7280) );
  NANDN U14914 ( .A(init), .B(e[418]), .Z(n11425) );
  AND U14915 ( .A(n11426), .B(n11427), .Z(n11424) );
  NAND U14916 ( .A(ereg[417]), .B(n9759), .Z(n11427) );
  NANDN U14917 ( .A(n9754), .B(ereg[418]), .Z(n11426) );
  NAND U14918 ( .A(n11428), .B(n11429), .Z(n7279) );
  NANDN U14919 ( .A(init), .B(e[419]), .Z(n11429) );
  AND U14920 ( .A(n11430), .B(n11431), .Z(n11428) );
  NAND U14921 ( .A(ereg[418]), .B(n9759), .Z(n11431) );
  NANDN U14922 ( .A(n9754), .B(ereg[419]), .Z(n11430) );
  NAND U14923 ( .A(n11432), .B(n11433), .Z(n7278) );
  NANDN U14924 ( .A(init), .B(e[420]), .Z(n11433) );
  AND U14925 ( .A(n11434), .B(n11435), .Z(n11432) );
  NAND U14926 ( .A(ereg[419]), .B(n9759), .Z(n11435) );
  NANDN U14927 ( .A(n9754), .B(ereg[420]), .Z(n11434) );
  NAND U14928 ( .A(n11436), .B(n11437), .Z(n7277) );
  NANDN U14929 ( .A(init), .B(e[421]), .Z(n11437) );
  AND U14930 ( .A(n11438), .B(n11439), .Z(n11436) );
  NAND U14931 ( .A(ereg[420]), .B(n9759), .Z(n11439) );
  NANDN U14932 ( .A(n9754), .B(ereg[421]), .Z(n11438) );
  NAND U14933 ( .A(n11440), .B(n11441), .Z(n7276) );
  NANDN U14934 ( .A(init), .B(e[422]), .Z(n11441) );
  AND U14935 ( .A(n11442), .B(n11443), .Z(n11440) );
  NAND U14936 ( .A(ereg[421]), .B(n9759), .Z(n11443) );
  NANDN U14937 ( .A(n9754), .B(ereg[422]), .Z(n11442) );
  NAND U14938 ( .A(n11444), .B(n11445), .Z(n7275) );
  NANDN U14939 ( .A(init), .B(e[423]), .Z(n11445) );
  AND U14940 ( .A(n11446), .B(n11447), .Z(n11444) );
  NAND U14941 ( .A(ereg[422]), .B(n9759), .Z(n11447) );
  NANDN U14942 ( .A(n9754), .B(ereg[423]), .Z(n11446) );
  NAND U14943 ( .A(n11448), .B(n11449), .Z(n7274) );
  NANDN U14944 ( .A(init), .B(e[424]), .Z(n11449) );
  AND U14945 ( .A(n11450), .B(n11451), .Z(n11448) );
  NAND U14946 ( .A(ereg[423]), .B(n9759), .Z(n11451) );
  NANDN U14947 ( .A(n9754), .B(ereg[424]), .Z(n11450) );
  NAND U14948 ( .A(n11452), .B(n11453), .Z(n7273) );
  NANDN U14949 ( .A(init), .B(e[425]), .Z(n11453) );
  AND U14950 ( .A(n11454), .B(n11455), .Z(n11452) );
  NAND U14951 ( .A(ereg[424]), .B(n9759), .Z(n11455) );
  NANDN U14952 ( .A(n9754), .B(ereg[425]), .Z(n11454) );
  NAND U14953 ( .A(n11456), .B(n11457), .Z(n7272) );
  NANDN U14954 ( .A(init), .B(e[426]), .Z(n11457) );
  AND U14955 ( .A(n11458), .B(n11459), .Z(n11456) );
  NAND U14956 ( .A(ereg[425]), .B(n9759), .Z(n11459) );
  NANDN U14957 ( .A(n9754), .B(ereg[426]), .Z(n11458) );
  NAND U14958 ( .A(n11460), .B(n11461), .Z(n7271) );
  NANDN U14959 ( .A(init), .B(e[427]), .Z(n11461) );
  AND U14960 ( .A(n11462), .B(n11463), .Z(n11460) );
  NAND U14961 ( .A(ereg[426]), .B(n9759), .Z(n11463) );
  NANDN U14962 ( .A(n9754), .B(ereg[427]), .Z(n11462) );
  NAND U14963 ( .A(n11464), .B(n11465), .Z(n7270) );
  NANDN U14964 ( .A(init), .B(e[428]), .Z(n11465) );
  AND U14965 ( .A(n11466), .B(n11467), .Z(n11464) );
  NAND U14966 ( .A(ereg[427]), .B(n9759), .Z(n11467) );
  NANDN U14967 ( .A(n9754), .B(ereg[428]), .Z(n11466) );
  NAND U14968 ( .A(n11468), .B(n11469), .Z(n7269) );
  NANDN U14969 ( .A(init), .B(e[429]), .Z(n11469) );
  AND U14970 ( .A(n11470), .B(n11471), .Z(n11468) );
  NAND U14971 ( .A(ereg[428]), .B(n9759), .Z(n11471) );
  NANDN U14972 ( .A(n9754), .B(ereg[429]), .Z(n11470) );
  NAND U14973 ( .A(n11472), .B(n11473), .Z(n7268) );
  NANDN U14974 ( .A(init), .B(e[430]), .Z(n11473) );
  AND U14975 ( .A(n11474), .B(n11475), .Z(n11472) );
  NAND U14976 ( .A(ereg[429]), .B(n9759), .Z(n11475) );
  NANDN U14977 ( .A(n9754), .B(ereg[430]), .Z(n11474) );
  NAND U14978 ( .A(n11476), .B(n11477), .Z(n7267) );
  NANDN U14979 ( .A(init), .B(e[431]), .Z(n11477) );
  AND U14980 ( .A(n11478), .B(n11479), .Z(n11476) );
  NAND U14981 ( .A(ereg[430]), .B(n9759), .Z(n11479) );
  NANDN U14982 ( .A(n9754), .B(ereg[431]), .Z(n11478) );
  NAND U14983 ( .A(n11480), .B(n11481), .Z(n7266) );
  NANDN U14984 ( .A(init), .B(e[432]), .Z(n11481) );
  AND U14985 ( .A(n11482), .B(n11483), .Z(n11480) );
  NAND U14986 ( .A(ereg[431]), .B(n9759), .Z(n11483) );
  NANDN U14987 ( .A(n9754), .B(ereg[432]), .Z(n11482) );
  NAND U14988 ( .A(n11484), .B(n11485), .Z(n7265) );
  NANDN U14989 ( .A(init), .B(e[433]), .Z(n11485) );
  AND U14990 ( .A(n11486), .B(n11487), .Z(n11484) );
  NAND U14991 ( .A(ereg[432]), .B(n9759), .Z(n11487) );
  NANDN U14992 ( .A(n9754), .B(ereg[433]), .Z(n11486) );
  NAND U14993 ( .A(n11488), .B(n11489), .Z(n7264) );
  NANDN U14994 ( .A(init), .B(e[434]), .Z(n11489) );
  AND U14995 ( .A(n11490), .B(n11491), .Z(n11488) );
  NAND U14996 ( .A(ereg[433]), .B(n9759), .Z(n11491) );
  NANDN U14997 ( .A(n9754), .B(ereg[434]), .Z(n11490) );
  NAND U14998 ( .A(n11492), .B(n11493), .Z(n7263) );
  NANDN U14999 ( .A(init), .B(e[435]), .Z(n11493) );
  AND U15000 ( .A(n11494), .B(n11495), .Z(n11492) );
  NAND U15001 ( .A(ereg[434]), .B(n9759), .Z(n11495) );
  NANDN U15002 ( .A(n9754), .B(ereg[435]), .Z(n11494) );
  NAND U15003 ( .A(n11496), .B(n11497), .Z(n7262) );
  NANDN U15004 ( .A(init), .B(e[436]), .Z(n11497) );
  AND U15005 ( .A(n11498), .B(n11499), .Z(n11496) );
  NAND U15006 ( .A(ereg[435]), .B(n9759), .Z(n11499) );
  NANDN U15007 ( .A(n9754), .B(ereg[436]), .Z(n11498) );
  NAND U15008 ( .A(n11500), .B(n11501), .Z(n7261) );
  NANDN U15009 ( .A(init), .B(e[437]), .Z(n11501) );
  AND U15010 ( .A(n11502), .B(n11503), .Z(n11500) );
  NAND U15011 ( .A(ereg[436]), .B(n9759), .Z(n11503) );
  NANDN U15012 ( .A(n9754), .B(ereg[437]), .Z(n11502) );
  NAND U15013 ( .A(n11504), .B(n11505), .Z(n7260) );
  NANDN U15014 ( .A(init), .B(e[438]), .Z(n11505) );
  AND U15015 ( .A(n11506), .B(n11507), .Z(n11504) );
  NAND U15016 ( .A(ereg[437]), .B(n9759), .Z(n11507) );
  NANDN U15017 ( .A(n9754), .B(ereg[438]), .Z(n11506) );
  NAND U15018 ( .A(n11508), .B(n11509), .Z(n7259) );
  NANDN U15019 ( .A(init), .B(e[439]), .Z(n11509) );
  AND U15020 ( .A(n11510), .B(n11511), .Z(n11508) );
  NAND U15021 ( .A(ereg[438]), .B(n9759), .Z(n11511) );
  NANDN U15022 ( .A(n9754), .B(ereg[439]), .Z(n11510) );
  NAND U15023 ( .A(n11512), .B(n11513), .Z(n7258) );
  NANDN U15024 ( .A(init), .B(e[440]), .Z(n11513) );
  AND U15025 ( .A(n11514), .B(n11515), .Z(n11512) );
  NAND U15026 ( .A(ereg[439]), .B(n9759), .Z(n11515) );
  NANDN U15027 ( .A(n9754), .B(ereg[440]), .Z(n11514) );
  NAND U15028 ( .A(n11516), .B(n11517), .Z(n7257) );
  NANDN U15029 ( .A(init), .B(e[441]), .Z(n11517) );
  AND U15030 ( .A(n11518), .B(n11519), .Z(n11516) );
  NAND U15031 ( .A(ereg[440]), .B(n9759), .Z(n11519) );
  NANDN U15032 ( .A(n9754), .B(ereg[441]), .Z(n11518) );
  NAND U15033 ( .A(n11520), .B(n11521), .Z(n7256) );
  NANDN U15034 ( .A(init), .B(e[442]), .Z(n11521) );
  AND U15035 ( .A(n11522), .B(n11523), .Z(n11520) );
  NAND U15036 ( .A(ereg[441]), .B(n9759), .Z(n11523) );
  NANDN U15037 ( .A(n9754), .B(ereg[442]), .Z(n11522) );
  NAND U15038 ( .A(n11524), .B(n11525), .Z(n7255) );
  NANDN U15039 ( .A(init), .B(e[443]), .Z(n11525) );
  AND U15040 ( .A(n11526), .B(n11527), .Z(n11524) );
  NAND U15041 ( .A(ereg[442]), .B(n9759), .Z(n11527) );
  NANDN U15042 ( .A(n9754), .B(ereg[443]), .Z(n11526) );
  NAND U15043 ( .A(n11528), .B(n11529), .Z(n7254) );
  NANDN U15044 ( .A(init), .B(e[444]), .Z(n11529) );
  AND U15045 ( .A(n11530), .B(n11531), .Z(n11528) );
  NAND U15046 ( .A(ereg[443]), .B(n9759), .Z(n11531) );
  NANDN U15047 ( .A(n9754), .B(ereg[444]), .Z(n11530) );
  NAND U15048 ( .A(n11532), .B(n11533), .Z(n7253) );
  NANDN U15049 ( .A(init), .B(e[445]), .Z(n11533) );
  AND U15050 ( .A(n11534), .B(n11535), .Z(n11532) );
  NAND U15051 ( .A(ereg[444]), .B(n9759), .Z(n11535) );
  NANDN U15052 ( .A(n9754), .B(ereg[445]), .Z(n11534) );
  NAND U15053 ( .A(n11536), .B(n11537), .Z(n7252) );
  NANDN U15054 ( .A(init), .B(e[446]), .Z(n11537) );
  AND U15055 ( .A(n11538), .B(n11539), .Z(n11536) );
  NAND U15056 ( .A(ereg[445]), .B(n9759), .Z(n11539) );
  NANDN U15057 ( .A(n9754), .B(ereg[446]), .Z(n11538) );
  NAND U15058 ( .A(n11540), .B(n11541), .Z(n7251) );
  NANDN U15059 ( .A(init), .B(e[447]), .Z(n11541) );
  AND U15060 ( .A(n11542), .B(n11543), .Z(n11540) );
  NAND U15061 ( .A(ereg[446]), .B(n9759), .Z(n11543) );
  NANDN U15062 ( .A(n9754), .B(ereg[447]), .Z(n11542) );
  NAND U15063 ( .A(n11544), .B(n11545), .Z(n7250) );
  NANDN U15064 ( .A(init), .B(e[448]), .Z(n11545) );
  AND U15065 ( .A(n11546), .B(n11547), .Z(n11544) );
  NAND U15066 ( .A(ereg[447]), .B(n9759), .Z(n11547) );
  NANDN U15067 ( .A(n9754), .B(ereg[448]), .Z(n11546) );
  NAND U15068 ( .A(n11548), .B(n11549), .Z(n7249) );
  NANDN U15069 ( .A(init), .B(e[449]), .Z(n11549) );
  AND U15070 ( .A(n11550), .B(n11551), .Z(n11548) );
  NAND U15071 ( .A(ereg[448]), .B(n9759), .Z(n11551) );
  NANDN U15072 ( .A(n9754), .B(ereg[449]), .Z(n11550) );
  NAND U15073 ( .A(n11552), .B(n11553), .Z(n7248) );
  NANDN U15074 ( .A(init), .B(e[450]), .Z(n11553) );
  AND U15075 ( .A(n11554), .B(n11555), .Z(n11552) );
  NAND U15076 ( .A(ereg[449]), .B(n9759), .Z(n11555) );
  NANDN U15077 ( .A(n9754), .B(ereg[450]), .Z(n11554) );
  NAND U15078 ( .A(n11556), .B(n11557), .Z(n7247) );
  NANDN U15079 ( .A(init), .B(e[451]), .Z(n11557) );
  AND U15080 ( .A(n11558), .B(n11559), .Z(n11556) );
  NAND U15081 ( .A(ereg[450]), .B(n9759), .Z(n11559) );
  NANDN U15082 ( .A(n9754), .B(ereg[451]), .Z(n11558) );
  NAND U15083 ( .A(n11560), .B(n11561), .Z(n7246) );
  NANDN U15084 ( .A(init), .B(e[452]), .Z(n11561) );
  AND U15085 ( .A(n11562), .B(n11563), .Z(n11560) );
  NAND U15086 ( .A(ereg[451]), .B(n9759), .Z(n11563) );
  NANDN U15087 ( .A(n9754), .B(ereg[452]), .Z(n11562) );
  NAND U15088 ( .A(n11564), .B(n11565), .Z(n7245) );
  NANDN U15089 ( .A(init), .B(e[453]), .Z(n11565) );
  AND U15090 ( .A(n11566), .B(n11567), .Z(n11564) );
  NAND U15091 ( .A(ereg[452]), .B(n9759), .Z(n11567) );
  NANDN U15092 ( .A(n9754), .B(ereg[453]), .Z(n11566) );
  NAND U15093 ( .A(n11568), .B(n11569), .Z(n7244) );
  NANDN U15094 ( .A(init), .B(e[454]), .Z(n11569) );
  AND U15095 ( .A(n11570), .B(n11571), .Z(n11568) );
  NAND U15096 ( .A(ereg[453]), .B(n9759), .Z(n11571) );
  NANDN U15097 ( .A(n9754), .B(ereg[454]), .Z(n11570) );
  NAND U15098 ( .A(n11572), .B(n11573), .Z(n7243) );
  NANDN U15099 ( .A(init), .B(e[455]), .Z(n11573) );
  AND U15100 ( .A(n11574), .B(n11575), .Z(n11572) );
  NAND U15101 ( .A(ereg[454]), .B(n9759), .Z(n11575) );
  NANDN U15102 ( .A(n9754), .B(ereg[455]), .Z(n11574) );
  NAND U15103 ( .A(n11576), .B(n11577), .Z(n7242) );
  NANDN U15104 ( .A(init), .B(e[456]), .Z(n11577) );
  AND U15105 ( .A(n11578), .B(n11579), .Z(n11576) );
  NAND U15106 ( .A(ereg[455]), .B(n9759), .Z(n11579) );
  NANDN U15107 ( .A(n9754), .B(ereg[456]), .Z(n11578) );
  NAND U15108 ( .A(n11580), .B(n11581), .Z(n7241) );
  NANDN U15109 ( .A(init), .B(e[457]), .Z(n11581) );
  AND U15110 ( .A(n11582), .B(n11583), .Z(n11580) );
  NAND U15111 ( .A(ereg[456]), .B(n9759), .Z(n11583) );
  NANDN U15112 ( .A(n9754), .B(ereg[457]), .Z(n11582) );
  NAND U15113 ( .A(n11584), .B(n11585), .Z(n7240) );
  NANDN U15114 ( .A(init), .B(e[458]), .Z(n11585) );
  AND U15115 ( .A(n11586), .B(n11587), .Z(n11584) );
  NAND U15116 ( .A(ereg[457]), .B(n9759), .Z(n11587) );
  NANDN U15117 ( .A(n9754), .B(ereg[458]), .Z(n11586) );
  NAND U15118 ( .A(n11588), .B(n11589), .Z(n7239) );
  NANDN U15119 ( .A(init), .B(e[459]), .Z(n11589) );
  AND U15120 ( .A(n11590), .B(n11591), .Z(n11588) );
  NAND U15121 ( .A(ereg[458]), .B(n9759), .Z(n11591) );
  NANDN U15122 ( .A(n9754), .B(ereg[459]), .Z(n11590) );
  NAND U15123 ( .A(n11592), .B(n11593), .Z(n7238) );
  NANDN U15124 ( .A(init), .B(e[460]), .Z(n11593) );
  AND U15125 ( .A(n11594), .B(n11595), .Z(n11592) );
  NAND U15126 ( .A(ereg[459]), .B(n9759), .Z(n11595) );
  NANDN U15127 ( .A(n9754), .B(ereg[460]), .Z(n11594) );
  NAND U15128 ( .A(n11596), .B(n11597), .Z(n7237) );
  NANDN U15129 ( .A(init), .B(e[461]), .Z(n11597) );
  AND U15130 ( .A(n11598), .B(n11599), .Z(n11596) );
  NAND U15131 ( .A(ereg[460]), .B(n9759), .Z(n11599) );
  NANDN U15132 ( .A(n9754), .B(ereg[461]), .Z(n11598) );
  NAND U15133 ( .A(n11600), .B(n11601), .Z(n7236) );
  NANDN U15134 ( .A(init), .B(e[462]), .Z(n11601) );
  AND U15135 ( .A(n11602), .B(n11603), .Z(n11600) );
  NAND U15136 ( .A(ereg[461]), .B(n9759), .Z(n11603) );
  NANDN U15137 ( .A(n9754), .B(ereg[462]), .Z(n11602) );
  NAND U15138 ( .A(n11604), .B(n11605), .Z(n7235) );
  NANDN U15139 ( .A(init), .B(e[463]), .Z(n11605) );
  AND U15140 ( .A(n11606), .B(n11607), .Z(n11604) );
  NAND U15141 ( .A(ereg[462]), .B(n9759), .Z(n11607) );
  NANDN U15142 ( .A(n9754), .B(ereg[463]), .Z(n11606) );
  NAND U15143 ( .A(n11608), .B(n11609), .Z(n7234) );
  NANDN U15144 ( .A(init), .B(e[464]), .Z(n11609) );
  AND U15145 ( .A(n11610), .B(n11611), .Z(n11608) );
  NAND U15146 ( .A(ereg[463]), .B(n9759), .Z(n11611) );
  NANDN U15147 ( .A(n9754), .B(ereg[464]), .Z(n11610) );
  NAND U15148 ( .A(n11612), .B(n11613), .Z(n7233) );
  NANDN U15149 ( .A(init), .B(e[465]), .Z(n11613) );
  AND U15150 ( .A(n11614), .B(n11615), .Z(n11612) );
  NAND U15151 ( .A(ereg[464]), .B(n9759), .Z(n11615) );
  NANDN U15152 ( .A(n9754), .B(ereg[465]), .Z(n11614) );
  NAND U15153 ( .A(n11616), .B(n11617), .Z(n7232) );
  NANDN U15154 ( .A(init), .B(e[466]), .Z(n11617) );
  AND U15155 ( .A(n11618), .B(n11619), .Z(n11616) );
  NAND U15156 ( .A(ereg[465]), .B(n9759), .Z(n11619) );
  NANDN U15157 ( .A(n9754), .B(ereg[466]), .Z(n11618) );
  NAND U15158 ( .A(n11620), .B(n11621), .Z(n7231) );
  NANDN U15159 ( .A(init), .B(e[467]), .Z(n11621) );
  AND U15160 ( .A(n11622), .B(n11623), .Z(n11620) );
  NAND U15161 ( .A(ereg[466]), .B(n9759), .Z(n11623) );
  NANDN U15162 ( .A(n9754), .B(ereg[467]), .Z(n11622) );
  NAND U15163 ( .A(n11624), .B(n11625), .Z(n7230) );
  NANDN U15164 ( .A(init), .B(e[468]), .Z(n11625) );
  AND U15165 ( .A(n11626), .B(n11627), .Z(n11624) );
  NAND U15166 ( .A(ereg[467]), .B(n9759), .Z(n11627) );
  NANDN U15167 ( .A(n9754), .B(ereg[468]), .Z(n11626) );
  NAND U15168 ( .A(n11628), .B(n11629), .Z(n7229) );
  NANDN U15169 ( .A(init), .B(e[469]), .Z(n11629) );
  AND U15170 ( .A(n11630), .B(n11631), .Z(n11628) );
  NAND U15171 ( .A(ereg[468]), .B(n9759), .Z(n11631) );
  NANDN U15172 ( .A(n9754), .B(ereg[469]), .Z(n11630) );
  NAND U15173 ( .A(n11632), .B(n11633), .Z(n7228) );
  NANDN U15174 ( .A(init), .B(e[470]), .Z(n11633) );
  AND U15175 ( .A(n11634), .B(n11635), .Z(n11632) );
  NAND U15176 ( .A(ereg[469]), .B(n9759), .Z(n11635) );
  NANDN U15177 ( .A(n9754), .B(ereg[470]), .Z(n11634) );
  NAND U15178 ( .A(n11636), .B(n11637), .Z(n7227) );
  NANDN U15179 ( .A(init), .B(e[471]), .Z(n11637) );
  AND U15180 ( .A(n11638), .B(n11639), .Z(n11636) );
  NAND U15181 ( .A(ereg[470]), .B(n9759), .Z(n11639) );
  NANDN U15182 ( .A(n9754), .B(ereg[471]), .Z(n11638) );
  NAND U15183 ( .A(n11640), .B(n11641), .Z(n7226) );
  NANDN U15184 ( .A(init), .B(e[472]), .Z(n11641) );
  AND U15185 ( .A(n11642), .B(n11643), .Z(n11640) );
  NAND U15186 ( .A(ereg[471]), .B(n9759), .Z(n11643) );
  NANDN U15187 ( .A(n9754), .B(ereg[472]), .Z(n11642) );
  NAND U15188 ( .A(n11644), .B(n11645), .Z(n7225) );
  NANDN U15189 ( .A(init), .B(e[473]), .Z(n11645) );
  AND U15190 ( .A(n11646), .B(n11647), .Z(n11644) );
  NAND U15191 ( .A(ereg[472]), .B(n9759), .Z(n11647) );
  NANDN U15192 ( .A(n9754), .B(ereg[473]), .Z(n11646) );
  NAND U15193 ( .A(n11648), .B(n11649), .Z(n7224) );
  NANDN U15194 ( .A(init), .B(e[474]), .Z(n11649) );
  AND U15195 ( .A(n11650), .B(n11651), .Z(n11648) );
  NAND U15196 ( .A(ereg[473]), .B(n9759), .Z(n11651) );
  NANDN U15197 ( .A(n9754), .B(ereg[474]), .Z(n11650) );
  NAND U15198 ( .A(n11652), .B(n11653), .Z(n7223) );
  NANDN U15199 ( .A(init), .B(e[475]), .Z(n11653) );
  AND U15200 ( .A(n11654), .B(n11655), .Z(n11652) );
  NAND U15201 ( .A(ereg[474]), .B(n9759), .Z(n11655) );
  NANDN U15202 ( .A(n9754), .B(ereg[475]), .Z(n11654) );
  NAND U15203 ( .A(n11656), .B(n11657), .Z(n7222) );
  NANDN U15204 ( .A(init), .B(e[476]), .Z(n11657) );
  AND U15205 ( .A(n11658), .B(n11659), .Z(n11656) );
  NAND U15206 ( .A(ereg[475]), .B(n9759), .Z(n11659) );
  NANDN U15207 ( .A(n9754), .B(ereg[476]), .Z(n11658) );
  NAND U15208 ( .A(n11660), .B(n11661), .Z(n7221) );
  NANDN U15209 ( .A(init), .B(e[477]), .Z(n11661) );
  AND U15210 ( .A(n11662), .B(n11663), .Z(n11660) );
  NAND U15211 ( .A(ereg[476]), .B(n9759), .Z(n11663) );
  NANDN U15212 ( .A(n9754), .B(ereg[477]), .Z(n11662) );
  NAND U15213 ( .A(n11664), .B(n11665), .Z(n7220) );
  NANDN U15214 ( .A(init), .B(e[478]), .Z(n11665) );
  AND U15215 ( .A(n11666), .B(n11667), .Z(n11664) );
  NAND U15216 ( .A(ereg[477]), .B(n9759), .Z(n11667) );
  NANDN U15217 ( .A(n9754), .B(ereg[478]), .Z(n11666) );
  NAND U15218 ( .A(n11668), .B(n11669), .Z(n7219) );
  NANDN U15219 ( .A(init), .B(e[479]), .Z(n11669) );
  AND U15220 ( .A(n11670), .B(n11671), .Z(n11668) );
  NAND U15221 ( .A(ereg[478]), .B(n9759), .Z(n11671) );
  NANDN U15222 ( .A(n9754), .B(ereg[479]), .Z(n11670) );
  NAND U15223 ( .A(n11672), .B(n11673), .Z(n7218) );
  NANDN U15224 ( .A(init), .B(e[480]), .Z(n11673) );
  AND U15225 ( .A(n11674), .B(n11675), .Z(n11672) );
  NAND U15226 ( .A(ereg[479]), .B(n9759), .Z(n11675) );
  NANDN U15227 ( .A(n9754), .B(ereg[480]), .Z(n11674) );
  NAND U15228 ( .A(n11676), .B(n11677), .Z(n7217) );
  NANDN U15229 ( .A(init), .B(e[481]), .Z(n11677) );
  AND U15230 ( .A(n11678), .B(n11679), .Z(n11676) );
  NAND U15231 ( .A(ereg[480]), .B(n9759), .Z(n11679) );
  NANDN U15232 ( .A(n9754), .B(ereg[481]), .Z(n11678) );
  NAND U15233 ( .A(n11680), .B(n11681), .Z(n7216) );
  NANDN U15234 ( .A(init), .B(e[482]), .Z(n11681) );
  AND U15235 ( .A(n11682), .B(n11683), .Z(n11680) );
  NAND U15236 ( .A(ereg[481]), .B(n9759), .Z(n11683) );
  NANDN U15237 ( .A(n9754), .B(ereg[482]), .Z(n11682) );
  NAND U15238 ( .A(n11684), .B(n11685), .Z(n7215) );
  NANDN U15239 ( .A(init), .B(e[483]), .Z(n11685) );
  AND U15240 ( .A(n11686), .B(n11687), .Z(n11684) );
  NAND U15241 ( .A(ereg[482]), .B(n9759), .Z(n11687) );
  NANDN U15242 ( .A(n9754), .B(ereg[483]), .Z(n11686) );
  NAND U15243 ( .A(n11688), .B(n11689), .Z(n7214) );
  NANDN U15244 ( .A(init), .B(e[484]), .Z(n11689) );
  AND U15245 ( .A(n11690), .B(n11691), .Z(n11688) );
  NAND U15246 ( .A(ereg[483]), .B(n9759), .Z(n11691) );
  NANDN U15247 ( .A(n9754), .B(ereg[484]), .Z(n11690) );
  NAND U15248 ( .A(n11692), .B(n11693), .Z(n7213) );
  NANDN U15249 ( .A(init), .B(e[485]), .Z(n11693) );
  AND U15250 ( .A(n11694), .B(n11695), .Z(n11692) );
  NAND U15251 ( .A(ereg[484]), .B(n9759), .Z(n11695) );
  NANDN U15252 ( .A(n9754), .B(ereg[485]), .Z(n11694) );
  NAND U15253 ( .A(n11696), .B(n11697), .Z(n7212) );
  NANDN U15254 ( .A(init), .B(e[486]), .Z(n11697) );
  AND U15255 ( .A(n11698), .B(n11699), .Z(n11696) );
  NAND U15256 ( .A(ereg[485]), .B(n9759), .Z(n11699) );
  NANDN U15257 ( .A(n9754), .B(ereg[486]), .Z(n11698) );
  NAND U15258 ( .A(n11700), .B(n11701), .Z(n7211) );
  NANDN U15259 ( .A(init), .B(e[487]), .Z(n11701) );
  AND U15260 ( .A(n11702), .B(n11703), .Z(n11700) );
  NAND U15261 ( .A(ereg[486]), .B(n9759), .Z(n11703) );
  NANDN U15262 ( .A(n9754), .B(ereg[487]), .Z(n11702) );
  NAND U15263 ( .A(n11704), .B(n11705), .Z(n7210) );
  NANDN U15264 ( .A(init), .B(e[488]), .Z(n11705) );
  AND U15265 ( .A(n11706), .B(n11707), .Z(n11704) );
  NAND U15266 ( .A(ereg[487]), .B(n9759), .Z(n11707) );
  NANDN U15267 ( .A(n9754), .B(ereg[488]), .Z(n11706) );
  NAND U15268 ( .A(n11708), .B(n11709), .Z(n7209) );
  NANDN U15269 ( .A(init), .B(e[489]), .Z(n11709) );
  AND U15270 ( .A(n11710), .B(n11711), .Z(n11708) );
  NAND U15271 ( .A(ereg[488]), .B(n9759), .Z(n11711) );
  NANDN U15272 ( .A(n9754), .B(ereg[489]), .Z(n11710) );
  NAND U15273 ( .A(n11712), .B(n11713), .Z(n7208) );
  NANDN U15274 ( .A(init), .B(e[490]), .Z(n11713) );
  AND U15275 ( .A(n11714), .B(n11715), .Z(n11712) );
  NAND U15276 ( .A(ereg[489]), .B(n9759), .Z(n11715) );
  NANDN U15277 ( .A(n9754), .B(ereg[490]), .Z(n11714) );
  NAND U15278 ( .A(n11716), .B(n11717), .Z(n7207) );
  NANDN U15279 ( .A(init), .B(e[491]), .Z(n11717) );
  AND U15280 ( .A(n11718), .B(n11719), .Z(n11716) );
  NAND U15281 ( .A(ereg[490]), .B(n9759), .Z(n11719) );
  NANDN U15282 ( .A(n9754), .B(ereg[491]), .Z(n11718) );
  NAND U15283 ( .A(n11720), .B(n11721), .Z(n7206) );
  NANDN U15284 ( .A(init), .B(e[492]), .Z(n11721) );
  AND U15285 ( .A(n11722), .B(n11723), .Z(n11720) );
  NAND U15286 ( .A(ereg[491]), .B(n9759), .Z(n11723) );
  NANDN U15287 ( .A(n9754), .B(ereg[492]), .Z(n11722) );
  NAND U15288 ( .A(n11724), .B(n11725), .Z(n7205) );
  NANDN U15289 ( .A(init), .B(e[493]), .Z(n11725) );
  AND U15290 ( .A(n11726), .B(n11727), .Z(n11724) );
  NAND U15291 ( .A(ereg[492]), .B(n9759), .Z(n11727) );
  NANDN U15292 ( .A(n9754), .B(ereg[493]), .Z(n11726) );
  NAND U15293 ( .A(n11728), .B(n11729), .Z(n7204) );
  NANDN U15294 ( .A(init), .B(e[494]), .Z(n11729) );
  AND U15295 ( .A(n11730), .B(n11731), .Z(n11728) );
  NAND U15296 ( .A(ereg[493]), .B(n9759), .Z(n11731) );
  NANDN U15297 ( .A(n9754), .B(ereg[494]), .Z(n11730) );
  NAND U15298 ( .A(n11732), .B(n11733), .Z(n7203) );
  NANDN U15299 ( .A(init), .B(e[495]), .Z(n11733) );
  AND U15300 ( .A(n11734), .B(n11735), .Z(n11732) );
  NAND U15301 ( .A(ereg[494]), .B(n9759), .Z(n11735) );
  NANDN U15302 ( .A(n9754), .B(ereg[495]), .Z(n11734) );
  NAND U15303 ( .A(n11736), .B(n11737), .Z(n7202) );
  NANDN U15304 ( .A(init), .B(e[496]), .Z(n11737) );
  AND U15305 ( .A(n11738), .B(n11739), .Z(n11736) );
  NAND U15306 ( .A(ereg[495]), .B(n9759), .Z(n11739) );
  NANDN U15307 ( .A(n9754), .B(ereg[496]), .Z(n11738) );
  NAND U15308 ( .A(n11740), .B(n11741), .Z(n7201) );
  NANDN U15309 ( .A(init), .B(e[497]), .Z(n11741) );
  AND U15310 ( .A(n11742), .B(n11743), .Z(n11740) );
  NAND U15311 ( .A(ereg[496]), .B(n9759), .Z(n11743) );
  NANDN U15312 ( .A(n9754), .B(ereg[497]), .Z(n11742) );
  NAND U15313 ( .A(n11744), .B(n11745), .Z(n7200) );
  NANDN U15314 ( .A(init), .B(e[498]), .Z(n11745) );
  AND U15315 ( .A(n11746), .B(n11747), .Z(n11744) );
  NAND U15316 ( .A(ereg[497]), .B(n9759), .Z(n11747) );
  NANDN U15317 ( .A(n9754), .B(ereg[498]), .Z(n11746) );
  NAND U15318 ( .A(n11748), .B(n11749), .Z(n7199) );
  NANDN U15319 ( .A(init), .B(e[499]), .Z(n11749) );
  AND U15320 ( .A(n11750), .B(n11751), .Z(n11748) );
  NAND U15321 ( .A(ereg[498]), .B(n9759), .Z(n11751) );
  NANDN U15322 ( .A(n9754), .B(ereg[499]), .Z(n11750) );
  NAND U15323 ( .A(n11752), .B(n11753), .Z(n7198) );
  NANDN U15324 ( .A(init), .B(e[500]), .Z(n11753) );
  AND U15325 ( .A(n11754), .B(n11755), .Z(n11752) );
  NAND U15326 ( .A(ereg[499]), .B(n9759), .Z(n11755) );
  NANDN U15327 ( .A(n9754), .B(ereg[500]), .Z(n11754) );
  NAND U15328 ( .A(n11756), .B(n11757), .Z(n7197) );
  NANDN U15329 ( .A(init), .B(e[501]), .Z(n11757) );
  AND U15330 ( .A(n11758), .B(n11759), .Z(n11756) );
  NAND U15331 ( .A(ereg[500]), .B(n9759), .Z(n11759) );
  NANDN U15332 ( .A(n9754), .B(ereg[501]), .Z(n11758) );
  NAND U15333 ( .A(n11760), .B(n11761), .Z(n7196) );
  NANDN U15334 ( .A(init), .B(e[502]), .Z(n11761) );
  AND U15335 ( .A(n11762), .B(n11763), .Z(n11760) );
  NAND U15336 ( .A(ereg[501]), .B(n9759), .Z(n11763) );
  NANDN U15337 ( .A(n9754), .B(ereg[502]), .Z(n11762) );
  NAND U15338 ( .A(n11764), .B(n11765), .Z(n7195) );
  NANDN U15339 ( .A(init), .B(e[503]), .Z(n11765) );
  AND U15340 ( .A(n11766), .B(n11767), .Z(n11764) );
  NAND U15341 ( .A(ereg[502]), .B(n9759), .Z(n11767) );
  NANDN U15342 ( .A(n9754), .B(ereg[503]), .Z(n11766) );
  NAND U15343 ( .A(n11768), .B(n11769), .Z(n7194) );
  NANDN U15344 ( .A(init), .B(e[504]), .Z(n11769) );
  AND U15345 ( .A(n11770), .B(n11771), .Z(n11768) );
  NAND U15346 ( .A(ereg[503]), .B(n9759), .Z(n11771) );
  NANDN U15347 ( .A(n9754), .B(ereg[504]), .Z(n11770) );
  NAND U15348 ( .A(n11772), .B(n11773), .Z(n7193) );
  NANDN U15349 ( .A(init), .B(e[505]), .Z(n11773) );
  AND U15350 ( .A(n11774), .B(n11775), .Z(n11772) );
  NAND U15351 ( .A(ereg[504]), .B(n9759), .Z(n11775) );
  NANDN U15352 ( .A(n9754), .B(ereg[505]), .Z(n11774) );
  NAND U15353 ( .A(n11776), .B(n11777), .Z(n7192) );
  NANDN U15354 ( .A(init), .B(e[506]), .Z(n11777) );
  AND U15355 ( .A(n11778), .B(n11779), .Z(n11776) );
  NAND U15356 ( .A(ereg[505]), .B(n9759), .Z(n11779) );
  NANDN U15357 ( .A(n9754), .B(ereg[506]), .Z(n11778) );
  NAND U15358 ( .A(n11780), .B(n11781), .Z(n7191) );
  NANDN U15359 ( .A(init), .B(e[507]), .Z(n11781) );
  AND U15360 ( .A(n11782), .B(n11783), .Z(n11780) );
  NAND U15361 ( .A(ereg[506]), .B(n9759), .Z(n11783) );
  NANDN U15362 ( .A(n9754), .B(ereg[507]), .Z(n11782) );
  NAND U15363 ( .A(n11784), .B(n11785), .Z(n7190) );
  NANDN U15364 ( .A(init), .B(e[508]), .Z(n11785) );
  AND U15365 ( .A(n11786), .B(n11787), .Z(n11784) );
  NAND U15366 ( .A(ereg[507]), .B(n9759), .Z(n11787) );
  NANDN U15367 ( .A(n9754), .B(ereg[508]), .Z(n11786) );
  NAND U15368 ( .A(n11788), .B(n11789), .Z(n7189) );
  NANDN U15369 ( .A(init), .B(e[509]), .Z(n11789) );
  AND U15370 ( .A(n11790), .B(n11791), .Z(n11788) );
  NAND U15371 ( .A(ereg[508]), .B(n9759), .Z(n11791) );
  NANDN U15372 ( .A(n9754), .B(ereg[509]), .Z(n11790) );
  NAND U15373 ( .A(n11792), .B(n11793), .Z(n7188) );
  NANDN U15374 ( .A(init), .B(e[510]), .Z(n11793) );
  AND U15375 ( .A(n11794), .B(n11795), .Z(n11792) );
  NAND U15376 ( .A(ereg[509]), .B(n9759), .Z(n11795) );
  NANDN U15377 ( .A(n9754), .B(ereg[510]), .Z(n11794) );
  NAND U15378 ( .A(n11796), .B(n11797), .Z(n7187) );
  NANDN U15379 ( .A(init), .B(e[511]), .Z(n11797) );
  AND U15380 ( .A(n11798), .B(n11799), .Z(n11796) );
  NAND U15381 ( .A(ereg[510]), .B(n9759), .Z(n11799) );
  AND U15382 ( .A(n9754), .B(n14372), .Z(n9759) );
  NANDN U15383 ( .A(n9754), .B(ereg[511]), .Z(n11798) );
  AND U15384 ( .A(n11800), .B(n7702), .Z(n9754) );
  NANDN U15385 ( .A(mul_pow), .B(init), .Z(n7702) );
  NANDN U15386 ( .A(start_reg[511]), .B(init), .Z(n11800) );
  NAND U15387 ( .A(n11801), .B(n8835), .Z(n7186) );
  NANDN U15388 ( .A(init), .B(m[511]), .Z(n8835) );
  AND U15389 ( .A(n11802), .B(n11803), .Z(n11801) );
  NAND U15390 ( .A(o[511]), .B(n11804), .Z(n11803) );
  NANDN U15391 ( .A(n11805), .B(creg[511]), .Z(n11802) );
  NAND U15392 ( .A(n11806), .B(n9749), .Z(n7185) );
  NANDN U15393 ( .A(init), .B(m[0]), .Z(n9749) );
  AND U15394 ( .A(n11807), .B(n11808), .Z(n11806) );
  NAND U15395 ( .A(o[0]), .B(n11804), .Z(n11808) );
  NANDN U15396 ( .A(n11805), .B(creg[0]), .Z(n11807) );
  NAND U15397 ( .A(n11809), .B(n9527), .Z(n7184) );
  NANDN U15398 ( .A(init), .B(m[1]), .Z(n9527) );
  AND U15399 ( .A(n11810), .B(n11811), .Z(n11809) );
  NAND U15400 ( .A(o[1]), .B(n11804), .Z(n11811) );
  NANDN U15401 ( .A(n11805), .B(creg[1]), .Z(n11810) );
  NAND U15402 ( .A(n11812), .B(n9305), .Z(n7183) );
  NANDN U15403 ( .A(init), .B(m[2]), .Z(n9305) );
  AND U15404 ( .A(n11813), .B(n11814), .Z(n11812) );
  NAND U15405 ( .A(o[2]), .B(n11804), .Z(n11814) );
  NANDN U15406 ( .A(n11805), .B(creg[2]), .Z(n11813) );
  NAND U15407 ( .A(n11815), .B(n9083), .Z(n7182) );
  NANDN U15408 ( .A(init), .B(m[3]), .Z(n9083) );
  AND U15409 ( .A(n11816), .B(n11817), .Z(n11815) );
  NAND U15410 ( .A(o[3]), .B(n11804), .Z(n11817) );
  NANDN U15411 ( .A(n11805), .B(creg[3]), .Z(n11816) );
  NAND U15412 ( .A(n11818), .B(n8861), .Z(n7181) );
  NANDN U15413 ( .A(init), .B(m[4]), .Z(n8861) );
  AND U15414 ( .A(n11819), .B(n11820), .Z(n11818) );
  NAND U15415 ( .A(o[4]), .B(n11804), .Z(n11820) );
  NANDN U15416 ( .A(n11805), .B(creg[4]), .Z(n11819) );
  NAND U15417 ( .A(n11821), .B(n8815), .Z(n7180) );
  NANDN U15418 ( .A(init), .B(m[5]), .Z(n8815) );
  AND U15419 ( .A(n11822), .B(n11823), .Z(n11821) );
  NAND U15420 ( .A(o[5]), .B(n11804), .Z(n11823) );
  NANDN U15421 ( .A(n11805), .B(creg[5]), .Z(n11822) );
  NAND U15422 ( .A(n11824), .B(n8793), .Z(n7179) );
  NANDN U15423 ( .A(init), .B(m[6]), .Z(n8793) );
  AND U15424 ( .A(n11825), .B(n11826), .Z(n11824) );
  NAND U15425 ( .A(o[6]), .B(n11804), .Z(n11826) );
  NANDN U15426 ( .A(n11805), .B(creg[6]), .Z(n11825) );
  NAND U15427 ( .A(n11827), .B(n8771), .Z(n7178) );
  NANDN U15428 ( .A(init), .B(m[7]), .Z(n8771) );
  AND U15429 ( .A(n11828), .B(n11829), .Z(n11827) );
  NAND U15430 ( .A(o[7]), .B(n11804), .Z(n11829) );
  NANDN U15431 ( .A(n11805), .B(creg[7]), .Z(n11828) );
  NAND U15432 ( .A(n11830), .B(n8749), .Z(n7177) );
  NANDN U15433 ( .A(init), .B(m[8]), .Z(n8749) );
  AND U15434 ( .A(n11831), .B(n11832), .Z(n11830) );
  NAND U15435 ( .A(o[8]), .B(n11804), .Z(n11832) );
  NANDN U15436 ( .A(n11805), .B(creg[8]), .Z(n11831) );
  NAND U15437 ( .A(n11833), .B(n8727), .Z(n7176) );
  NANDN U15438 ( .A(init), .B(m[9]), .Z(n8727) );
  AND U15439 ( .A(n11834), .B(n11835), .Z(n11833) );
  NAND U15440 ( .A(o[9]), .B(n11804), .Z(n11835) );
  NANDN U15441 ( .A(n11805), .B(creg[9]), .Z(n11834) );
  NAND U15442 ( .A(n11836), .B(n9727), .Z(n7175) );
  NANDN U15443 ( .A(init), .B(m[10]), .Z(n9727) );
  AND U15444 ( .A(n11837), .B(n11838), .Z(n11836) );
  NAND U15445 ( .A(o[10]), .B(n11804), .Z(n11838) );
  NANDN U15446 ( .A(n11805), .B(creg[10]), .Z(n11837) );
  NAND U15447 ( .A(n11839), .B(n9705), .Z(n7174) );
  NANDN U15448 ( .A(init), .B(m[11]), .Z(n9705) );
  AND U15449 ( .A(n11840), .B(n11841), .Z(n11839) );
  NAND U15450 ( .A(o[11]), .B(n11804), .Z(n11841) );
  NANDN U15451 ( .A(n11805), .B(creg[11]), .Z(n11840) );
  NAND U15452 ( .A(n11842), .B(n9683), .Z(n7173) );
  NANDN U15453 ( .A(init), .B(m[12]), .Z(n9683) );
  AND U15454 ( .A(n11843), .B(n11844), .Z(n11842) );
  NAND U15455 ( .A(o[12]), .B(n11804), .Z(n11844) );
  NANDN U15456 ( .A(n11805), .B(creg[12]), .Z(n11843) );
  NAND U15457 ( .A(n11845), .B(n9661), .Z(n7172) );
  NANDN U15458 ( .A(init), .B(m[13]), .Z(n9661) );
  AND U15459 ( .A(n11846), .B(n11847), .Z(n11845) );
  NAND U15460 ( .A(o[13]), .B(n11804), .Z(n11847) );
  NANDN U15461 ( .A(n11805), .B(creg[13]), .Z(n11846) );
  NAND U15462 ( .A(n11848), .B(n9639), .Z(n7171) );
  NANDN U15463 ( .A(init), .B(m[14]), .Z(n9639) );
  AND U15464 ( .A(n11849), .B(n11850), .Z(n11848) );
  NAND U15465 ( .A(o[14]), .B(n11804), .Z(n11850) );
  NANDN U15466 ( .A(n11805), .B(creg[14]), .Z(n11849) );
  NAND U15467 ( .A(n11851), .B(n9617), .Z(n7170) );
  NANDN U15468 ( .A(init), .B(m[15]), .Z(n9617) );
  AND U15469 ( .A(n11852), .B(n11853), .Z(n11851) );
  NAND U15470 ( .A(o[15]), .B(n11804), .Z(n11853) );
  NANDN U15471 ( .A(n11805), .B(creg[15]), .Z(n11852) );
  NAND U15472 ( .A(n11854), .B(n9595), .Z(n7169) );
  NANDN U15473 ( .A(init), .B(m[16]), .Z(n9595) );
  AND U15474 ( .A(n11855), .B(n11856), .Z(n11854) );
  NAND U15475 ( .A(o[16]), .B(n11804), .Z(n11856) );
  NANDN U15476 ( .A(n11805), .B(creg[16]), .Z(n11855) );
  NAND U15477 ( .A(n11857), .B(n9573), .Z(n7168) );
  NANDN U15478 ( .A(init), .B(m[17]), .Z(n9573) );
  AND U15479 ( .A(n11858), .B(n11859), .Z(n11857) );
  NAND U15480 ( .A(o[17]), .B(n11804), .Z(n11859) );
  NANDN U15481 ( .A(n11805), .B(creg[17]), .Z(n11858) );
  NAND U15482 ( .A(n11860), .B(n9551), .Z(n7167) );
  NANDN U15483 ( .A(init), .B(m[18]), .Z(n9551) );
  AND U15484 ( .A(n11861), .B(n11862), .Z(n11860) );
  NAND U15485 ( .A(o[18]), .B(n11804), .Z(n11862) );
  NANDN U15486 ( .A(n11805), .B(creg[18]), .Z(n11861) );
  NAND U15487 ( .A(n11863), .B(n9529), .Z(n7166) );
  NANDN U15488 ( .A(init), .B(m[19]), .Z(n9529) );
  AND U15489 ( .A(n11864), .B(n11865), .Z(n11863) );
  NAND U15490 ( .A(o[19]), .B(n11804), .Z(n11865) );
  NANDN U15491 ( .A(n11805), .B(creg[19]), .Z(n11864) );
  NAND U15492 ( .A(n11866), .B(n9505), .Z(n7165) );
  NANDN U15493 ( .A(init), .B(m[20]), .Z(n9505) );
  AND U15494 ( .A(n11867), .B(n11868), .Z(n11866) );
  NAND U15495 ( .A(o[20]), .B(n11804), .Z(n11868) );
  NANDN U15496 ( .A(n11805), .B(creg[20]), .Z(n11867) );
  NAND U15497 ( .A(n11869), .B(n9483), .Z(n7164) );
  NANDN U15498 ( .A(init), .B(m[21]), .Z(n9483) );
  AND U15499 ( .A(n11870), .B(n11871), .Z(n11869) );
  NAND U15500 ( .A(o[21]), .B(n11804), .Z(n11871) );
  NANDN U15501 ( .A(n11805), .B(creg[21]), .Z(n11870) );
  NAND U15502 ( .A(n11872), .B(n9461), .Z(n7163) );
  NANDN U15503 ( .A(init), .B(m[22]), .Z(n9461) );
  AND U15504 ( .A(n11873), .B(n11874), .Z(n11872) );
  NAND U15505 ( .A(o[22]), .B(n11804), .Z(n11874) );
  NANDN U15506 ( .A(n11805), .B(creg[22]), .Z(n11873) );
  NAND U15507 ( .A(n11875), .B(n9439), .Z(n7162) );
  NANDN U15508 ( .A(init), .B(m[23]), .Z(n9439) );
  AND U15509 ( .A(n11876), .B(n11877), .Z(n11875) );
  NAND U15510 ( .A(o[23]), .B(n11804), .Z(n11877) );
  NANDN U15511 ( .A(n11805), .B(creg[23]), .Z(n11876) );
  NAND U15512 ( .A(n11878), .B(n9417), .Z(n7161) );
  NANDN U15513 ( .A(init), .B(m[24]), .Z(n9417) );
  AND U15514 ( .A(n11879), .B(n11880), .Z(n11878) );
  NAND U15515 ( .A(o[24]), .B(n11804), .Z(n11880) );
  NANDN U15516 ( .A(n11805), .B(creg[24]), .Z(n11879) );
  NAND U15517 ( .A(n11881), .B(n9395), .Z(n7160) );
  NANDN U15518 ( .A(init), .B(m[25]), .Z(n9395) );
  AND U15519 ( .A(n11882), .B(n11883), .Z(n11881) );
  NAND U15520 ( .A(o[25]), .B(n11804), .Z(n11883) );
  NANDN U15521 ( .A(n11805), .B(creg[25]), .Z(n11882) );
  NAND U15522 ( .A(n11884), .B(n9373), .Z(n7159) );
  NANDN U15523 ( .A(init), .B(m[26]), .Z(n9373) );
  AND U15524 ( .A(n11885), .B(n11886), .Z(n11884) );
  NAND U15525 ( .A(o[26]), .B(n11804), .Z(n11886) );
  NANDN U15526 ( .A(n11805), .B(creg[26]), .Z(n11885) );
  NAND U15527 ( .A(n11887), .B(n9351), .Z(n7158) );
  NANDN U15528 ( .A(init), .B(m[27]), .Z(n9351) );
  AND U15529 ( .A(n11888), .B(n11889), .Z(n11887) );
  NAND U15530 ( .A(o[27]), .B(n11804), .Z(n11889) );
  NANDN U15531 ( .A(n11805), .B(creg[27]), .Z(n11888) );
  NAND U15532 ( .A(n11890), .B(n9329), .Z(n7157) );
  NANDN U15533 ( .A(init), .B(m[28]), .Z(n9329) );
  AND U15534 ( .A(n11891), .B(n11892), .Z(n11890) );
  NAND U15535 ( .A(o[28]), .B(n11804), .Z(n11892) );
  NANDN U15536 ( .A(n11805), .B(creg[28]), .Z(n11891) );
  NAND U15537 ( .A(n11893), .B(n9307), .Z(n7156) );
  NANDN U15538 ( .A(init), .B(m[29]), .Z(n9307) );
  AND U15539 ( .A(n11894), .B(n11895), .Z(n11893) );
  NAND U15540 ( .A(o[29]), .B(n11804), .Z(n11895) );
  NANDN U15541 ( .A(n11805), .B(creg[29]), .Z(n11894) );
  NAND U15542 ( .A(n11896), .B(n9283), .Z(n7155) );
  NANDN U15543 ( .A(init), .B(m[30]), .Z(n9283) );
  AND U15544 ( .A(n11897), .B(n11898), .Z(n11896) );
  NAND U15545 ( .A(o[30]), .B(n11804), .Z(n11898) );
  NANDN U15546 ( .A(n11805), .B(creg[30]), .Z(n11897) );
  NAND U15547 ( .A(n11899), .B(n9261), .Z(n7154) );
  NANDN U15548 ( .A(init), .B(m[31]), .Z(n9261) );
  AND U15549 ( .A(n11900), .B(n11901), .Z(n11899) );
  NAND U15550 ( .A(o[31]), .B(n11804), .Z(n11901) );
  NANDN U15551 ( .A(n11805), .B(creg[31]), .Z(n11900) );
  NAND U15552 ( .A(n11902), .B(n9239), .Z(n7153) );
  NANDN U15553 ( .A(init), .B(m[32]), .Z(n9239) );
  AND U15554 ( .A(n11903), .B(n11904), .Z(n11902) );
  NAND U15555 ( .A(o[32]), .B(n11804), .Z(n11904) );
  NANDN U15556 ( .A(n11805), .B(creg[32]), .Z(n11903) );
  NAND U15557 ( .A(n11905), .B(n9217), .Z(n7152) );
  NANDN U15558 ( .A(init), .B(m[33]), .Z(n9217) );
  AND U15559 ( .A(n11906), .B(n11907), .Z(n11905) );
  NAND U15560 ( .A(o[33]), .B(n11804), .Z(n11907) );
  NANDN U15561 ( .A(n11805), .B(creg[33]), .Z(n11906) );
  NAND U15562 ( .A(n11908), .B(n9195), .Z(n7151) );
  NANDN U15563 ( .A(init), .B(m[34]), .Z(n9195) );
  AND U15564 ( .A(n11909), .B(n11910), .Z(n11908) );
  NAND U15565 ( .A(o[34]), .B(n11804), .Z(n11910) );
  NANDN U15566 ( .A(n11805), .B(creg[34]), .Z(n11909) );
  NAND U15567 ( .A(n11911), .B(n9173), .Z(n7150) );
  NANDN U15568 ( .A(init), .B(m[35]), .Z(n9173) );
  AND U15569 ( .A(n11912), .B(n11913), .Z(n11911) );
  NAND U15570 ( .A(o[35]), .B(n11804), .Z(n11913) );
  NANDN U15571 ( .A(n11805), .B(creg[35]), .Z(n11912) );
  NAND U15572 ( .A(n11914), .B(n9151), .Z(n7149) );
  NANDN U15573 ( .A(init), .B(m[36]), .Z(n9151) );
  AND U15574 ( .A(n11915), .B(n11916), .Z(n11914) );
  NAND U15575 ( .A(o[36]), .B(n11804), .Z(n11916) );
  NANDN U15576 ( .A(n11805), .B(creg[36]), .Z(n11915) );
  NAND U15577 ( .A(n11917), .B(n9129), .Z(n7148) );
  NANDN U15578 ( .A(init), .B(m[37]), .Z(n9129) );
  AND U15579 ( .A(n11918), .B(n11919), .Z(n11917) );
  NAND U15580 ( .A(o[37]), .B(n11804), .Z(n11919) );
  NANDN U15581 ( .A(n11805), .B(creg[37]), .Z(n11918) );
  NAND U15582 ( .A(n11920), .B(n9107), .Z(n7147) );
  NANDN U15583 ( .A(init), .B(m[38]), .Z(n9107) );
  AND U15584 ( .A(n11921), .B(n11922), .Z(n11920) );
  NAND U15585 ( .A(o[38]), .B(n11804), .Z(n11922) );
  NANDN U15586 ( .A(n11805), .B(creg[38]), .Z(n11921) );
  NAND U15587 ( .A(n11923), .B(n9085), .Z(n7146) );
  NANDN U15588 ( .A(init), .B(m[39]), .Z(n9085) );
  AND U15589 ( .A(n11924), .B(n11925), .Z(n11923) );
  NAND U15590 ( .A(o[39]), .B(n11804), .Z(n11925) );
  NANDN U15591 ( .A(n11805), .B(creg[39]), .Z(n11924) );
  NAND U15592 ( .A(n11926), .B(n9061), .Z(n7145) );
  NANDN U15593 ( .A(init), .B(m[40]), .Z(n9061) );
  AND U15594 ( .A(n11927), .B(n11928), .Z(n11926) );
  NAND U15595 ( .A(o[40]), .B(n11804), .Z(n11928) );
  NANDN U15596 ( .A(n11805), .B(creg[40]), .Z(n11927) );
  NAND U15597 ( .A(n11929), .B(n9039), .Z(n7144) );
  NANDN U15598 ( .A(init), .B(m[41]), .Z(n9039) );
  AND U15599 ( .A(n11930), .B(n11931), .Z(n11929) );
  NAND U15600 ( .A(o[41]), .B(n11804), .Z(n11931) );
  NANDN U15601 ( .A(n11805), .B(creg[41]), .Z(n11930) );
  NAND U15602 ( .A(n11932), .B(n9017), .Z(n7143) );
  NANDN U15603 ( .A(init), .B(m[42]), .Z(n9017) );
  AND U15604 ( .A(n11933), .B(n11934), .Z(n11932) );
  NAND U15605 ( .A(o[42]), .B(n11804), .Z(n11934) );
  NANDN U15606 ( .A(n11805), .B(creg[42]), .Z(n11933) );
  NAND U15607 ( .A(n11935), .B(n8995), .Z(n7142) );
  NANDN U15608 ( .A(init), .B(m[43]), .Z(n8995) );
  AND U15609 ( .A(n11936), .B(n11937), .Z(n11935) );
  NAND U15610 ( .A(o[43]), .B(n11804), .Z(n11937) );
  NANDN U15611 ( .A(n11805), .B(creg[43]), .Z(n11936) );
  NAND U15612 ( .A(n11938), .B(n8973), .Z(n7141) );
  NANDN U15613 ( .A(init), .B(m[44]), .Z(n8973) );
  AND U15614 ( .A(n11939), .B(n11940), .Z(n11938) );
  NAND U15615 ( .A(o[44]), .B(n11804), .Z(n11940) );
  NANDN U15616 ( .A(n11805), .B(creg[44]), .Z(n11939) );
  NAND U15617 ( .A(n11941), .B(n8951), .Z(n7140) );
  NANDN U15618 ( .A(init), .B(m[45]), .Z(n8951) );
  AND U15619 ( .A(n11942), .B(n11943), .Z(n11941) );
  NAND U15620 ( .A(o[45]), .B(n11804), .Z(n11943) );
  NANDN U15621 ( .A(n11805), .B(creg[45]), .Z(n11942) );
  NAND U15622 ( .A(n11944), .B(n8929), .Z(n7139) );
  NANDN U15623 ( .A(init), .B(m[46]), .Z(n8929) );
  AND U15624 ( .A(n11945), .B(n11946), .Z(n11944) );
  NAND U15625 ( .A(o[46]), .B(n11804), .Z(n11946) );
  NANDN U15626 ( .A(n11805), .B(creg[46]), .Z(n11945) );
  NAND U15627 ( .A(n11947), .B(n8907), .Z(n7138) );
  NANDN U15628 ( .A(init), .B(m[47]), .Z(n8907) );
  AND U15629 ( .A(n11948), .B(n11949), .Z(n11947) );
  NAND U15630 ( .A(o[47]), .B(n11804), .Z(n11949) );
  NANDN U15631 ( .A(n11805), .B(creg[47]), .Z(n11948) );
  NAND U15632 ( .A(n11950), .B(n8885), .Z(n7137) );
  NANDN U15633 ( .A(init), .B(m[48]), .Z(n8885) );
  AND U15634 ( .A(n11951), .B(n11952), .Z(n11950) );
  NAND U15635 ( .A(o[48]), .B(n11804), .Z(n11952) );
  NANDN U15636 ( .A(n11805), .B(creg[48]), .Z(n11951) );
  NAND U15637 ( .A(n11953), .B(n8863), .Z(n7136) );
  NANDN U15638 ( .A(init), .B(m[49]), .Z(n8863) );
  AND U15639 ( .A(n11954), .B(n11955), .Z(n11953) );
  NAND U15640 ( .A(o[49]), .B(n11804), .Z(n11955) );
  NANDN U15641 ( .A(n11805), .B(creg[49]), .Z(n11954) );
  NAND U15642 ( .A(n11956), .B(n8839), .Z(n7135) );
  NANDN U15643 ( .A(init), .B(m[50]), .Z(n8839) );
  AND U15644 ( .A(n11957), .B(n11958), .Z(n11956) );
  NAND U15645 ( .A(o[50]), .B(n11804), .Z(n11958) );
  NANDN U15646 ( .A(n11805), .B(creg[50]), .Z(n11957) );
  NAND U15647 ( .A(n11959), .B(n8833), .Z(n7134) );
  NANDN U15648 ( .A(init), .B(m[51]), .Z(n8833) );
  AND U15649 ( .A(n11960), .B(n11961), .Z(n11959) );
  NAND U15650 ( .A(o[51]), .B(n11804), .Z(n11961) );
  NANDN U15651 ( .A(n11805), .B(creg[51]), .Z(n11960) );
  NAND U15652 ( .A(n11962), .B(n8831), .Z(n7133) );
  NANDN U15653 ( .A(init), .B(m[52]), .Z(n8831) );
  AND U15654 ( .A(n11963), .B(n11964), .Z(n11962) );
  NAND U15655 ( .A(o[52]), .B(n11804), .Z(n11964) );
  NANDN U15656 ( .A(n11805), .B(creg[52]), .Z(n11963) );
  NAND U15657 ( .A(n11965), .B(n8829), .Z(n7132) );
  NANDN U15658 ( .A(init), .B(m[53]), .Z(n8829) );
  AND U15659 ( .A(n11966), .B(n11967), .Z(n11965) );
  NAND U15660 ( .A(o[53]), .B(n11804), .Z(n11967) );
  NANDN U15661 ( .A(n11805), .B(creg[53]), .Z(n11966) );
  NAND U15662 ( .A(n11968), .B(n8827), .Z(n7131) );
  NANDN U15663 ( .A(init), .B(m[54]), .Z(n8827) );
  AND U15664 ( .A(n11969), .B(n11970), .Z(n11968) );
  NAND U15665 ( .A(o[54]), .B(n11804), .Z(n11970) );
  NANDN U15666 ( .A(n11805), .B(creg[54]), .Z(n11969) );
  NAND U15667 ( .A(n11971), .B(n8825), .Z(n7130) );
  NANDN U15668 ( .A(init), .B(m[55]), .Z(n8825) );
  AND U15669 ( .A(n11972), .B(n11973), .Z(n11971) );
  NAND U15670 ( .A(o[55]), .B(n11804), .Z(n11973) );
  NANDN U15671 ( .A(n11805), .B(creg[55]), .Z(n11972) );
  NAND U15672 ( .A(n11974), .B(n8823), .Z(n7129) );
  NANDN U15673 ( .A(init), .B(m[56]), .Z(n8823) );
  AND U15674 ( .A(n11975), .B(n11976), .Z(n11974) );
  NAND U15675 ( .A(o[56]), .B(n11804), .Z(n11976) );
  NANDN U15676 ( .A(n11805), .B(creg[56]), .Z(n11975) );
  NAND U15677 ( .A(n11977), .B(n8821), .Z(n7128) );
  NANDN U15678 ( .A(init), .B(m[57]), .Z(n8821) );
  AND U15679 ( .A(n11978), .B(n11979), .Z(n11977) );
  NAND U15680 ( .A(o[57]), .B(n11804), .Z(n11979) );
  NANDN U15681 ( .A(n11805), .B(creg[57]), .Z(n11978) );
  NAND U15682 ( .A(n11980), .B(n8819), .Z(n7127) );
  NANDN U15683 ( .A(init), .B(m[58]), .Z(n8819) );
  AND U15684 ( .A(n11981), .B(n11982), .Z(n11980) );
  NAND U15685 ( .A(o[58]), .B(n11804), .Z(n11982) );
  NANDN U15686 ( .A(n11805), .B(creg[58]), .Z(n11981) );
  NAND U15687 ( .A(n11983), .B(n8817), .Z(n7126) );
  NANDN U15688 ( .A(init), .B(m[59]), .Z(n8817) );
  AND U15689 ( .A(n11984), .B(n11985), .Z(n11983) );
  NAND U15690 ( .A(o[59]), .B(n11804), .Z(n11985) );
  NANDN U15691 ( .A(n11805), .B(creg[59]), .Z(n11984) );
  NAND U15692 ( .A(n11986), .B(n8813), .Z(n7125) );
  NANDN U15693 ( .A(init), .B(m[60]), .Z(n8813) );
  AND U15694 ( .A(n11987), .B(n11988), .Z(n11986) );
  NAND U15695 ( .A(o[60]), .B(n11804), .Z(n11988) );
  NANDN U15696 ( .A(n11805), .B(creg[60]), .Z(n11987) );
  NAND U15697 ( .A(n11989), .B(n8811), .Z(n7124) );
  NANDN U15698 ( .A(init), .B(m[61]), .Z(n8811) );
  AND U15699 ( .A(n11990), .B(n11991), .Z(n11989) );
  NAND U15700 ( .A(o[61]), .B(n11804), .Z(n11991) );
  NANDN U15701 ( .A(n11805), .B(creg[61]), .Z(n11990) );
  NAND U15702 ( .A(n11992), .B(n8809), .Z(n7123) );
  NANDN U15703 ( .A(init), .B(m[62]), .Z(n8809) );
  AND U15704 ( .A(n11993), .B(n11994), .Z(n11992) );
  NAND U15705 ( .A(o[62]), .B(n11804), .Z(n11994) );
  NANDN U15706 ( .A(n11805), .B(creg[62]), .Z(n11993) );
  NAND U15707 ( .A(n11995), .B(n8807), .Z(n7122) );
  NANDN U15708 ( .A(init), .B(m[63]), .Z(n8807) );
  AND U15709 ( .A(n11996), .B(n11997), .Z(n11995) );
  NAND U15710 ( .A(o[63]), .B(n11804), .Z(n11997) );
  NANDN U15711 ( .A(n11805), .B(creg[63]), .Z(n11996) );
  NAND U15712 ( .A(n11998), .B(n8805), .Z(n7121) );
  NANDN U15713 ( .A(init), .B(m[64]), .Z(n8805) );
  AND U15714 ( .A(n11999), .B(n12000), .Z(n11998) );
  NAND U15715 ( .A(o[64]), .B(n11804), .Z(n12000) );
  NANDN U15716 ( .A(n11805), .B(creg[64]), .Z(n11999) );
  NAND U15717 ( .A(n12001), .B(n8803), .Z(n7120) );
  NANDN U15718 ( .A(init), .B(m[65]), .Z(n8803) );
  AND U15719 ( .A(n12002), .B(n12003), .Z(n12001) );
  NAND U15720 ( .A(o[65]), .B(n11804), .Z(n12003) );
  NANDN U15721 ( .A(n11805), .B(creg[65]), .Z(n12002) );
  NAND U15722 ( .A(n12004), .B(n8801), .Z(n7119) );
  NANDN U15723 ( .A(init), .B(m[66]), .Z(n8801) );
  AND U15724 ( .A(n12005), .B(n12006), .Z(n12004) );
  NAND U15725 ( .A(o[66]), .B(n11804), .Z(n12006) );
  NANDN U15726 ( .A(n11805), .B(creg[66]), .Z(n12005) );
  NAND U15727 ( .A(n12007), .B(n8799), .Z(n7118) );
  NANDN U15728 ( .A(init), .B(m[67]), .Z(n8799) );
  AND U15729 ( .A(n12008), .B(n12009), .Z(n12007) );
  NAND U15730 ( .A(o[67]), .B(n11804), .Z(n12009) );
  NANDN U15731 ( .A(n11805), .B(creg[67]), .Z(n12008) );
  NAND U15732 ( .A(n12010), .B(n8797), .Z(n7117) );
  NANDN U15733 ( .A(init), .B(m[68]), .Z(n8797) );
  AND U15734 ( .A(n12011), .B(n12012), .Z(n12010) );
  NAND U15735 ( .A(o[68]), .B(n11804), .Z(n12012) );
  NANDN U15736 ( .A(n11805), .B(creg[68]), .Z(n12011) );
  NAND U15737 ( .A(n12013), .B(n8795), .Z(n7116) );
  NANDN U15738 ( .A(init), .B(m[69]), .Z(n8795) );
  AND U15739 ( .A(n12014), .B(n12015), .Z(n12013) );
  NAND U15740 ( .A(o[69]), .B(n11804), .Z(n12015) );
  NANDN U15741 ( .A(n11805), .B(creg[69]), .Z(n12014) );
  NAND U15742 ( .A(n12016), .B(n8791), .Z(n7115) );
  NANDN U15743 ( .A(init), .B(m[70]), .Z(n8791) );
  AND U15744 ( .A(n12017), .B(n12018), .Z(n12016) );
  NAND U15745 ( .A(o[70]), .B(n11804), .Z(n12018) );
  NANDN U15746 ( .A(n11805), .B(creg[70]), .Z(n12017) );
  NAND U15747 ( .A(n12019), .B(n8789), .Z(n7114) );
  NANDN U15748 ( .A(init), .B(m[71]), .Z(n8789) );
  AND U15749 ( .A(n12020), .B(n12021), .Z(n12019) );
  NAND U15750 ( .A(o[71]), .B(n11804), .Z(n12021) );
  NANDN U15751 ( .A(n11805), .B(creg[71]), .Z(n12020) );
  NAND U15752 ( .A(n12022), .B(n8787), .Z(n7113) );
  NANDN U15753 ( .A(init), .B(m[72]), .Z(n8787) );
  AND U15754 ( .A(n12023), .B(n12024), .Z(n12022) );
  NAND U15755 ( .A(o[72]), .B(n11804), .Z(n12024) );
  NANDN U15756 ( .A(n11805), .B(creg[72]), .Z(n12023) );
  NAND U15757 ( .A(n12025), .B(n8785), .Z(n7112) );
  NANDN U15758 ( .A(init), .B(m[73]), .Z(n8785) );
  AND U15759 ( .A(n12026), .B(n12027), .Z(n12025) );
  NAND U15760 ( .A(o[73]), .B(n11804), .Z(n12027) );
  NANDN U15761 ( .A(n11805), .B(creg[73]), .Z(n12026) );
  NAND U15762 ( .A(n12028), .B(n8783), .Z(n7111) );
  NANDN U15763 ( .A(init), .B(m[74]), .Z(n8783) );
  AND U15764 ( .A(n12029), .B(n12030), .Z(n12028) );
  NAND U15765 ( .A(o[74]), .B(n11804), .Z(n12030) );
  NANDN U15766 ( .A(n11805), .B(creg[74]), .Z(n12029) );
  NAND U15767 ( .A(n12031), .B(n8781), .Z(n7110) );
  NANDN U15768 ( .A(init), .B(m[75]), .Z(n8781) );
  AND U15769 ( .A(n12032), .B(n12033), .Z(n12031) );
  NAND U15770 ( .A(o[75]), .B(n11804), .Z(n12033) );
  NANDN U15771 ( .A(n11805), .B(creg[75]), .Z(n12032) );
  NAND U15772 ( .A(n12034), .B(n8779), .Z(n7109) );
  NANDN U15773 ( .A(init), .B(m[76]), .Z(n8779) );
  AND U15774 ( .A(n12035), .B(n12036), .Z(n12034) );
  NAND U15775 ( .A(o[76]), .B(n11804), .Z(n12036) );
  NANDN U15776 ( .A(n11805), .B(creg[76]), .Z(n12035) );
  NAND U15777 ( .A(n12037), .B(n8777), .Z(n7108) );
  NANDN U15778 ( .A(init), .B(m[77]), .Z(n8777) );
  AND U15779 ( .A(n12038), .B(n12039), .Z(n12037) );
  NAND U15780 ( .A(o[77]), .B(n11804), .Z(n12039) );
  NANDN U15781 ( .A(n11805), .B(creg[77]), .Z(n12038) );
  NAND U15782 ( .A(n12040), .B(n8775), .Z(n7107) );
  NANDN U15783 ( .A(init), .B(m[78]), .Z(n8775) );
  AND U15784 ( .A(n12041), .B(n12042), .Z(n12040) );
  NAND U15785 ( .A(o[78]), .B(n11804), .Z(n12042) );
  NANDN U15786 ( .A(n11805), .B(creg[78]), .Z(n12041) );
  NAND U15787 ( .A(n12043), .B(n8773), .Z(n7106) );
  NANDN U15788 ( .A(init), .B(m[79]), .Z(n8773) );
  AND U15789 ( .A(n12044), .B(n12045), .Z(n12043) );
  NAND U15790 ( .A(o[79]), .B(n11804), .Z(n12045) );
  NANDN U15791 ( .A(n11805), .B(creg[79]), .Z(n12044) );
  NAND U15792 ( .A(n12046), .B(n8769), .Z(n7105) );
  NANDN U15793 ( .A(init), .B(m[80]), .Z(n8769) );
  AND U15794 ( .A(n12047), .B(n12048), .Z(n12046) );
  NAND U15795 ( .A(o[80]), .B(n11804), .Z(n12048) );
  NANDN U15796 ( .A(n11805), .B(creg[80]), .Z(n12047) );
  NAND U15797 ( .A(n12049), .B(n8767), .Z(n7104) );
  NANDN U15798 ( .A(init), .B(m[81]), .Z(n8767) );
  AND U15799 ( .A(n12050), .B(n12051), .Z(n12049) );
  NAND U15800 ( .A(o[81]), .B(n11804), .Z(n12051) );
  NANDN U15801 ( .A(n11805), .B(creg[81]), .Z(n12050) );
  NAND U15802 ( .A(n12052), .B(n8765), .Z(n7103) );
  NANDN U15803 ( .A(init), .B(m[82]), .Z(n8765) );
  AND U15804 ( .A(n12053), .B(n12054), .Z(n12052) );
  NAND U15805 ( .A(o[82]), .B(n11804), .Z(n12054) );
  NANDN U15806 ( .A(n11805), .B(creg[82]), .Z(n12053) );
  NAND U15807 ( .A(n12055), .B(n8763), .Z(n7102) );
  NANDN U15808 ( .A(init), .B(m[83]), .Z(n8763) );
  AND U15809 ( .A(n12056), .B(n12057), .Z(n12055) );
  NAND U15810 ( .A(o[83]), .B(n11804), .Z(n12057) );
  NANDN U15811 ( .A(n11805), .B(creg[83]), .Z(n12056) );
  NAND U15812 ( .A(n12058), .B(n8761), .Z(n7101) );
  NANDN U15813 ( .A(init), .B(m[84]), .Z(n8761) );
  AND U15814 ( .A(n12059), .B(n12060), .Z(n12058) );
  NAND U15815 ( .A(o[84]), .B(n11804), .Z(n12060) );
  NANDN U15816 ( .A(n11805), .B(creg[84]), .Z(n12059) );
  NAND U15817 ( .A(n12061), .B(n8759), .Z(n7100) );
  NANDN U15818 ( .A(init), .B(m[85]), .Z(n8759) );
  AND U15819 ( .A(n12062), .B(n12063), .Z(n12061) );
  NAND U15820 ( .A(o[85]), .B(n11804), .Z(n12063) );
  NANDN U15821 ( .A(n11805), .B(creg[85]), .Z(n12062) );
  NAND U15822 ( .A(n12064), .B(n8757), .Z(n7099) );
  NANDN U15823 ( .A(init), .B(m[86]), .Z(n8757) );
  AND U15824 ( .A(n12065), .B(n12066), .Z(n12064) );
  NAND U15825 ( .A(o[86]), .B(n11804), .Z(n12066) );
  NANDN U15826 ( .A(n11805), .B(creg[86]), .Z(n12065) );
  NAND U15827 ( .A(n12067), .B(n8755), .Z(n7098) );
  NANDN U15828 ( .A(init), .B(m[87]), .Z(n8755) );
  AND U15829 ( .A(n12068), .B(n12069), .Z(n12067) );
  NAND U15830 ( .A(o[87]), .B(n11804), .Z(n12069) );
  NANDN U15831 ( .A(n11805), .B(creg[87]), .Z(n12068) );
  NAND U15832 ( .A(n12070), .B(n8753), .Z(n7097) );
  NANDN U15833 ( .A(init), .B(m[88]), .Z(n8753) );
  AND U15834 ( .A(n12071), .B(n12072), .Z(n12070) );
  NAND U15835 ( .A(o[88]), .B(n11804), .Z(n12072) );
  NANDN U15836 ( .A(n11805), .B(creg[88]), .Z(n12071) );
  NAND U15837 ( .A(n12073), .B(n8751), .Z(n7096) );
  NANDN U15838 ( .A(init), .B(m[89]), .Z(n8751) );
  AND U15839 ( .A(n12074), .B(n12075), .Z(n12073) );
  NAND U15840 ( .A(o[89]), .B(n11804), .Z(n12075) );
  NANDN U15841 ( .A(n11805), .B(creg[89]), .Z(n12074) );
  NAND U15842 ( .A(n12076), .B(n8747), .Z(n7095) );
  NANDN U15843 ( .A(init), .B(m[90]), .Z(n8747) );
  AND U15844 ( .A(n12077), .B(n12078), .Z(n12076) );
  NAND U15845 ( .A(o[90]), .B(n11804), .Z(n12078) );
  NANDN U15846 ( .A(n11805), .B(creg[90]), .Z(n12077) );
  NAND U15847 ( .A(n12079), .B(n8745), .Z(n7094) );
  NANDN U15848 ( .A(init), .B(m[91]), .Z(n8745) );
  AND U15849 ( .A(n12080), .B(n12081), .Z(n12079) );
  NAND U15850 ( .A(o[91]), .B(n11804), .Z(n12081) );
  NANDN U15851 ( .A(n11805), .B(creg[91]), .Z(n12080) );
  NAND U15852 ( .A(n12082), .B(n8743), .Z(n7093) );
  NANDN U15853 ( .A(init), .B(m[92]), .Z(n8743) );
  AND U15854 ( .A(n12083), .B(n12084), .Z(n12082) );
  NAND U15855 ( .A(o[92]), .B(n11804), .Z(n12084) );
  NANDN U15856 ( .A(n11805), .B(creg[92]), .Z(n12083) );
  NAND U15857 ( .A(n12085), .B(n8741), .Z(n7092) );
  NANDN U15858 ( .A(init), .B(m[93]), .Z(n8741) );
  AND U15859 ( .A(n12086), .B(n12087), .Z(n12085) );
  NAND U15860 ( .A(o[93]), .B(n11804), .Z(n12087) );
  NANDN U15861 ( .A(n11805), .B(creg[93]), .Z(n12086) );
  NAND U15862 ( .A(n12088), .B(n8739), .Z(n7091) );
  NANDN U15863 ( .A(init), .B(m[94]), .Z(n8739) );
  AND U15864 ( .A(n12089), .B(n12090), .Z(n12088) );
  NAND U15865 ( .A(o[94]), .B(n11804), .Z(n12090) );
  NANDN U15866 ( .A(n11805), .B(creg[94]), .Z(n12089) );
  NAND U15867 ( .A(n12091), .B(n8737), .Z(n7090) );
  NANDN U15868 ( .A(init), .B(m[95]), .Z(n8737) );
  AND U15869 ( .A(n12092), .B(n12093), .Z(n12091) );
  NAND U15870 ( .A(o[95]), .B(n11804), .Z(n12093) );
  NANDN U15871 ( .A(n11805), .B(creg[95]), .Z(n12092) );
  NAND U15872 ( .A(n12094), .B(n8735), .Z(n7089) );
  NANDN U15873 ( .A(init), .B(m[96]), .Z(n8735) );
  AND U15874 ( .A(n12095), .B(n12096), .Z(n12094) );
  NAND U15875 ( .A(o[96]), .B(n11804), .Z(n12096) );
  NANDN U15876 ( .A(n11805), .B(creg[96]), .Z(n12095) );
  NAND U15877 ( .A(n12097), .B(n8733), .Z(n7088) );
  NANDN U15878 ( .A(init), .B(m[97]), .Z(n8733) );
  AND U15879 ( .A(n12098), .B(n12099), .Z(n12097) );
  NAND U15880 ( .A(o[97]), .B(n11804), .Z(n12099) );
  NANDN U15881 ( .A(n11805), .B(creg[97]), .Z(n12098) );
  NAND U15882 ( .A(n12100), .B(n8731), .Z(n7087) );
  NANDN U15883 ( .A(init), .B(m[98]), .Z(n8731) );
  AND U15884 ( .A(n12101), .B(n12102), .Z(n12100) );
  NAND U15885 ( .A(o[98]), .B(n11804), .Z(n12102) );
  NANDN U15886 ( .A(n11805), .B(creg[98]), .Z(n12101) );
  NAND U15887 ( .A(n12103), .B(n8729), .Z(n7086) );
  NANDN U15888 ( .A(init), .B(m[99]), .Z(n8729) );
  AND U15889 ( .A(n12104), .B(n12105), .Z(n12103) );
  NAND U15890 ( .A(o[99]), .B(n11804), .Z(n12105) );
  NANDN U15891 ( .A(n11805), .B(creg[99]), .Z(n12104) );
  NAND U15892 ( .A(n12106), .B(n9747), .Z(n7085) );
  NANDN U15893 ( .A(init), .B(m[100]), .Z(n9747) );
  AND U15894 ( .A(n12107), .B(n12108), .Z(n12106) );
  NAND U15895 ( .A(o[100]), .B(n11804), .Z(n12108) );
  NANDN U15896 ( .A(n11805), .B(creg[100]), .Z(n12107) );
  NAND U15897 ( .A(n12109), .B(n9745), .Z(n7084) );
  NANDN U15898 ( .A(init), .B(m[101]), .Z(n9745) );
  AND U15899 ( .A(n12110), .B(n12111), .Z(n12109) );
  NAND U15900 ( .A(o[101]), .B(n11804), .Z(n12111) );
  NANDN U15901 ( .A(n11805), .B(creg[101]), .Z(n12110) );
  NAND U15902 ( .A(n12112), .B(n9743), .Z(n7083) );
  NANDN U15903 ( .A(init), .B(m[102]), .Z(n9743) );
  AND U15904 ( .A(n12113), .B(n12114), .Z(n12112) );
  NAND U15905 ( .A(o[102]), .B(n11804), .Z(n12114) );
  NANDN U15906 ( .A(n11805), .B(creg[102]), .Z(n12113) );
  NAND U15907 ( .A(n12115), .B(n9741), .Z(n7082) );
  NANDN U15908 ( .A(init), .B(m[103]), .Z(n9741) );
  AND U15909 ( .A(n12116), .B(n12117), .Z(n12115) );
  NAND U15910 ( .A(o[103]), .B(n11804), .Z(n12117) );
  NANDN U15911 ( .A(n11805), .B(creg[103]), .Z(n12116) );
  NAND U15912 ( .A(n12118), .B(n9739), .Z(n7081) );
  NANDN U15913 ( .A(init), .B(m[104]), .Z(n9739) );
  AND U15914 ( .A(n12119), .B(n12120), .Z(n12118) );
  NAND U15915 ( .A(o[104]), .B(n11804), .Z(n12120) );
  NANDN U15916 ( .A(n11805), .B(creg[104]), .Z(n12119) );
  NAND U15917 ( .A(n12121), .B(n9737), .Z(n7080) );
  NANDN U15918 ( .A(init), .B(m[105]), .Z(n9737) );
  AND U15919 ( .A(n12122), .B(n12123), .Z(n12121) );
  NAND U15920 ( .A(o[105]), .B(n11804), .Z(n12123) );
  NANDN U15921 ( .A(n11805), .B(creg[105]), .Z(n12122) );
  NAND U15922 ( .A(n12124), .B(n9735), .Z(n7079) );
  NANDN U15923 ( .A(init), .B(m[106]), .Z(n9735) );
  AND U15924 ( .A(n12125), .B(n12126), .Z(n12124) );
  NAND U15925 ( .A(o[106]), .B(n11804), .Z(n12126) );
  NANDN U15926 ( .A(n11805), .B(creg[106]), .Z(n12125) );
  NAND U15927 ( .A(n12127), .B(n9733), .Z(n7078) );
  NANDN U15928 ( .A(init), .B(m[107]), .Z(n9733) );
  AND U15929 ( .A(n12128), .B(n12129), .Z(n12127) );
  NAND U15930 ( .A(o[107]), .B(n11804), .Z(n12129) );
  NANDN U15931 ( .A(n11805), .B(creg[107]), .Z(n12128) );
  NAND U15932 ( .A(n12130), .B(n9731), .Z(n7077) );
  NANDN U15933 ( .A(init), .B(m[108]), .Z(n9731) );
  AND U15934 ( .A(n12131), .B(n12132), .Z(n12130) );
  NAND U15935 ( .A(o[108]), .B(n11804), .Z(n12132) );
  NANDN U15936 ( .A(n11805), .B(creg[108]), .Z(n12131) );
  NAND U15937 ( .A(n12133), .B(n9729), .Z(n7076) );
  NANDN U15938 ( .A(init), .B(m[109]), .Z(n9729) );
  AND U15939 ( .A(n12134), .B(n12135), .Z(n12133) );
  NAND U15940 ( .A(o[109]), .B(n11804), .Z(n12135) );
  NANDN U15941 ( .A(n11805), .B(creg[109]), .Z(n12134) );
  NAND U15942 ( .A(n12136), .B(n9725), .Z(n7075) );
  NANDN U15943 ( .A(init), .B(m[110]), .Z(n9725) );
  AND U15944 ( .A(n12137), .B(n12138), .Z(n12136) );
  NAND U15945 ( .A(o[110]), .B(n11804), .Z(n12138) );
  NANDN U15946 ( .A(n11805), .B(creg[110]), .Z(n12137) );
  NAND U15947 ( .A(n12139), .B(n9723), .Z(n7074) );
  NANDN U15948 ( .A(init), .B(m[111]), .Z(n9723) );
  AND U15949 ( .A(n12140), .B(n12141), .Z(n12139) );
  NAND U15950 ( .A(o[111]), .B(n11804), .Z(n12141) );
  NANDN U15951 ( .A(n11805), .B(creg[111]), .Z(n12140) );
  NAND U15952 ( .A(n12142), .B(n9721), .Z(n7073) );
  NANDN U15953 ( .A(init), .B(m[112]), .Z(n9721) );
  AND U15954 ( .A(n12143), .B(n12144), .Z(n12142) );
  NAND U15955 ( .A(o[112]), .B(n11804), .Z(n12144) );
  NANDN U15956 ( .A(n11805), .B(creg[112]), .Z(n12143) );
  NAND U15957 ( .A(n12145), .B(n9719), .Z(n7072) );
  NANDN U15958 ( .A(init), .B(m[113]), .Z(n9719) );
  AND U15959 ( .A(n12146), .B(n12147), .Z(n12145) );
  NAND U15960 ( .A(o[113]), .B(n11804), .Z(n12147) );
  NANDN U15961 ( .A(n11805), .B(creg[113]), .Z(n12146) );
  NAND U15962 ( .A(n12148), .B(n9717), .Z(n7071) );
  NANDN U15963 ( .A(init), .B(m[114]), .Z(n9717) );
  AND U15964 ( .A(n12149), .B(n12150), .Z(n12148) );
  NAND U15965 ( .A(o[114]), .B(n11804), .Z(n12150) );
  NANDN U15966 ( .A(n11805), .B(creg[114]), .Z(n12149) );
  NAND U15967 ( .A(n12151), .B(n9715), .Z(n7070) );
  NANDN U15968 ( .A(init), .B(m[115]), .Z(n9715) );
  AND U15969 ( .A(n12152), .B(n12153), .Z(n12151) );
  NAND U15970 ( .A(o[115]), .B(n11804), .Z(n12153) );
  NANDN U15971 ( .A(n11805), .B(creg[115]), .Z(n12152) );
  NAND U15972 ( .A(n12154), .B(n9713), .Z(n7069) );
  NANDN U15973 ( .A(init), .B(m[116]), .Z(n9713) );
  AND U15974 ( .A(n12155), .B(n12156), .Z(n12154) );
  NAND U15975 ( .A(o[116]), .B(n11804), .Z(n12156) );
  NANDN U15976 ( .A(n11805), .B(creg[116]), .Z(n12155) );
  NAND U15977 ( .A(n12157), .B(n9711), .Z(n7068) );
  NANDN U15978 ( .A(init), .B(m[117]), .Z(n9711) );
  AND U15979 ( .A(n12158), .B(n12159), .Z(n12157) );
  NAND U15980 ( .A(o[117]), .B(n11804), .Z(n12159) );
  NANDN U15981 ( .A(n11805), .B(creg[117]), .Z(n12158) );
  NAND U15982 ( .A(n12160), .B(n9709), .Z(n7067) );
  NANDN U15983 ( .A(init), .B(m[118]), .Z(n9709) );
  AND U15984 ( .A(n12161), .B(n12162), .Z(n12160) );
  NAND U15985 ( .A(o[118]), .B(n11804), .Z(n12162) );
  NANDN U15986 ( .A(n11805), .B(creg[118]), .Z(n12161) );
  NAND U15987 ( .A(n12163), .B(n9707), .Z(n7066) );
  NANDN U15988 ( .A(init), .B(m[119]), .Z(n9707) );
  AND U15989 ( .A(n12164), .B(n12165), .Z(n12163) );
  NAND U15990 ( .A(o[119]), .B(n11804), .Z(n12165) );
  NANDN U15991 ( .A(n11805), .B(creg[119]), .Z(n12164) );
  NAND U15992 ( .A(n12166), .B(n9703), .Z(n7065) );
  NANDN U15993 ( .A(init), .B(m[120]), .Z(n9703) );
  AND U15994 ( .A(n12167), .B(n12168), .Z(n12166) );
  NAND U15995 ( .A(o[120]), .B(n11804), .Z(n12168) );
  NANDN U15996 ( .A(n11805), .B(creg[120]), .Z(n12167) );
  NAND U15997 ( .A(n12169), .B(n9701), .Z(n7064) );
  NANDN U15998 ( .A(init), .B(m[121]), .Z(n9701) );
  AND U15999 ( .A(n12170), .B(n12171), .Z(n12169) );
  NAND U16000 ( .A(o[121]), .B(n11804), .Z(n12171) );
  NANDN U16001 ( .A(n11805), .B(creg[121]), .Z(n12170) );
  NAND U16002 ( .A(n12172), .B(n9699), .Z(n7063) );
  NANDN U16003 ( .A(init), .B(m[122]), .Z(n9699) );
  AND U16004 ( .A(n12173), .B(n12174), .Z(n12172) );
  NAND U16005 ( .A(o[122]), .B(n11804), .Z(n12174) );
  NANDN U16006 ( .A(n11805), .B(creg[122]), .Z(n12173) );
  NAND U16007 ( .A(n12175), .B(n9697), .Z(n7062) );
  NANDN U16008 ( .A(init), .B(m[123]), .Z(n9697) );
  AND U16009 ( .A(n12176), .B(n12177), .Z(n12175) );
  NAND U16010 ( .A(o[123]), .B(n11804), .Z(n12177) );
  NANDN U16011 ( .A(n11805), .B(creg[123]), .Z(n12176) );
  NAND U16012 ( .A(n12178), .B(n9695), .Z(n7061) );
  NANDN U16013 ( .A(init), .B(m[124]), .Z(n9695) );
  AND U16014 ( .A(n12179), .B(n12180), .Z(n12178) );
  NAND U16015 ( .A(o[124]), .B(n11804), .Z(n12180) );
  NANDN U16016 ( .A(n11805), .B(creg[124]), .Z(n12179) );
  NAND U16017 ( .A(n12181), .B(n9693), .Z(n7060) );
  NANDN U16018 ( .A(init), .B(m[125]), .Z(n9693) );
  AND U16019 ( .A(n12182), .B(n12183), .Z(n12181) );
  NAND U16020 ( .A(o[125]), .B(n11804), .Z(n12183) );
  NANDN U16021 ( .A(n11805), .B(creg[125]), .Z(n12182) );
  NAND U16022 ( .A(n12184), .B(n9691), .Z(n7059) );
  NANDN U16023 ( .A(init), .B(m[126]), .Z(n9691) );
  AND U16024 ( .A(n12185), .B(n12186), .Z(n12184) );
  NAND U16025 ( .A(o[126]), .B(n11804), .Z(n12186) );
  NANDN U16026 ( .A(n11805), .B(creg[126]), .Z(n12185) );
  NAND U16027 ( .A(n12187), .B(n9689), .Z(n7058) );
  NANDN U16028 ( .A(init), .B(m[127]), .Z(n9689) );
  AND U16029 ( .A(n12188), .B(n12189), .Z(n12187) );
  NAND U16030 ( .A(o[127]), .B(n11804), .Z(n12189) );
  NANDN U16031 ( .A(n11805), .B(creg[127]), .Z(n12188) );
  NAND U16032 ( .A(n12190), .B(n9687), .Z(n7057) );
  NANDN U16033 ( .A(init), .B(m[128]), .Z(n9687) );
  AND U16034 ( .A(n12191), .B(n12192), .Z(n12190) );
  NAND U16035 ( .A(o[128]), .B(n11804), .Z(n12192) );
  NANDN U16036 ( .A(n11805), .B(creg[128]), .Z(n12191) );
  NAND U16037 ( .A(n12193), .B(n9685), .Z(n7056) );
  NANDN U16038 ( .A(init), .B(m[129]), .Z(n9685) );
  AND U16039 ( .A(n12194), .B(n12195), .Z(n12193) );
  NAND U16040 ( .A(o[129]), .B(n11804), .Z(n12195) );
  NANDN U16041 ( .A(n11805), .B(creg[129]), .Z(n12194) );
  NAND U16042 ( .A(n12196), .B(n9681), .Z(n7055) );
  NANDN U16043 ( .A(init), .B(m[130]), .Z(n9681) );
  AND U16044 ( .A(n12197), .B(n12198), .Z(n12196) );
  NAND U16045 ( .A(o[130]), .B(n11804), .Z(n12198) );
  NANDN U16046 ( .A(n11805), .B(creg[130]), .Z(n12197) );
  NAND U16047 ( .A(n12199), .B(n9679), .Z(n7054) );
  NANDN U16048 ( .A(init), .B(m[131]), .Z(n9679) );
  AND U16049 ( .A(n12200), .B(n12201), .Z(n12199) );
  NAND U16050 ( .A(o[131]), .B(n11804), .Z(n12201) );
  NANDN U16051 ( .A(n11805), .B(creg[131]), .Z(n12200) );
  NAND U16052 ( .A(n12202), .B(n9677), .Z(n7053) );
  NANDN U16053 ( .A(init), .B(m[132]), .Z(n9677) );
  AND U16054 ( .A(n12203), .B(n12204), .Z(n12202) );
  NAND U16055 ( .A(o[132]), .B(n11804), .Z(n12204) );
  NANDN U16056 ( .A(n11805), .B(creg[132]), .Z(n12203) );
  NAND U16057 ( .A(n12205), .B(n9675), .Z(n7052) );
  NANDN U16058 ( .A(init), .B(m[133]), .Z(n9675) );
  AND U16059 ( .A(n12206), .B(n12207), .Z(n12205) );
  NAND U16060 ( .A(o[133]), .B(n11804), .Z(n12207) );
  NANDN U16061 ( .A(n11805), .B(creg[133]), .Z(n12206) );
  NAND U16062 ( .A(n12208), .B(n9673), .Z(n7051) );
  NANDN U16063 ( .A(init), .B(m[134]), .Z(n9673) );
  AND U16064 ( .A(n12209), .B(n12210), .Z(n12208) );
  NAND U16065 ( .A(o[134]), .B(n11804), .Z(n12210) );
  NANDN U16066 ( .A(n11805), .B(creg[134]), .Z(n12209) );
  NAND U16067 ( .A(n12211), .B(n9671), .Z(n7050) );
  NANDN U16068 ( .A(init), .B(m[135]), .Z(n9671) );
  AND U16069 ( .A(n12212), .B(n12213), .Z(n12211) );
  NAND U16070 ( .A(o[135]), .B(n11804), .Z(n12213) );
  NANDN U16071 ( .A(n11805), .B(creg[135]), .Z(n12212) );
  NAND U16072 ( .A(n12214), .B(n9669), .Z(n7049) );
  NANDN U16073 ( .A(init), .B(m[136]), .Z(n9669) );
  AND U16074 ( .A(n12215), .B(n12216), .Z(n12214) );
  NAND U16075 ( .A(o[136]), .B(n11804), .Z(n12216) );
  NANDN U16076 ( .A(n11805), .B(creg[136]), .Z(n12215) );
  NAND U16077 ( .A(n12217), .B(n9667), .Z(n7048) );
  NANDN U16078 ( .A(init), .B(m[137]), .Z(n9667) );
  AND U16079 ( .A(n12218), .B(n12219), .Z(n12217) );
  NAND U16080 ( .A(o[137]), .B(n11804), .Z(n12219) );
  NANDN U16081 ( .A(n11805), .B(creg[137]), .Z(n12218) );
  NAND U16082 ( .A(n12220), .B(n9665), .Z(n7047) );
  NANDN U16083 ( .A(init), .B(m[138]), .Z(n9665) );
  AND U16084 ( .A(n12221), .B(n12222), .Z(n12220) );
  NAND U16085 ( .A(o[138]), .B(n11804), .Z(n12222) );
  NANDN U16086 ( .A(n11805), .B(creg[138]), .Z(n12221) );
  NAND U16087 ( .A(n12223), .B(n9663), .Z(n7046) );
  NANDN U16088 ( .A(init), .B(m[139]), .Z(n9663) );
  AND U16089 ( .A(n12224), .B(n12225), .Z(n12223) );
  NAND U16090 ( .A(o[139]), .B(n11804), .Z(n12225) );
  NANDN U16091 ( .A(n11805), .B(creg[139]), .Z(n12224) );
  NAND U16092 ( .A(n12226), .B(n9659), .Z(n7045) );
  NANDN U16093 ( .A(init), .B(m[140]), .Z(n9659) );
  AND U16094 ( .A(n12227), .B(n12228), .Z(n12226) );
  NAND U16095 ( .A(o[140]), .B(n11804), .Z(n12228) );
  NANDN U16096 ( .A(n11805), .B(creg[140]), .Z(n12227) );
  NAND U16097 ( .A(n12229), .B(n9657), .Z(n7044) );
  NANDN U16098 ( .A(init), .B(m[141]), .Z(n9657) );
  AND U16099 ( .A(n12230), .B(n12231), .Z(n12229) );
  NAND U16100 ( .A(o[141]), .B(n11804), .Z(n12231) );
  NANDN U16101 ( .A(n11805), .B(creg[141]), .Z(n12230) );
  NAND U16102 ( .A(n12232), .B(n9655), .Z(n7043) );
  NANDN U16103 ( .A(init), .B(m[142]), .Z(n9655) );
  AND U16104 ( .A(n12233), .B(n12234), .Z(n12232) );
  NAND U16105 ( .A(o[142]), .B(n11804), .Z(n12234) );
  NANDN U16106 ( .A(n11805), .B(creg[142]), .Z(n12233) );
  NAND U16107 ( .A(n12235), .B(n9653), .Z(n7042) );
  NANDN U16108 ( .A(init), .B(m[143]), .Z(n9653) );
  AND U16109 ( .A(n12236), .B(n12237), .Z(n12235) );
  NAND U16110 ( .A(o[143]), .B(n11804), .Z(n12237) );
  NANDN U16111 ( .A(n11805), .B(creg[143]), .Z(n12236) );
  NAND U16112 ( .A(n12238), .B(n9651), .Z(n7041) );
  NANDN U16113 ( .A(init), .B(m[144]), .Z(n9651) );
  AND U16114 ( .A(n12239), .B(n12240), .Z(n12238) );
  NAND U16115 ( .A(o[144]), .B(n11804), .Z(n12240) );
  NANDN U16116 ( .A(n11805), .B(creg[144]), .Z(n12239) );
  NAND U16117 ( .A(n12241), .B(n9649), .Z(n7040) );
  NANDN U16118 ( .A(init), .B(m[145]), .Z(n9649) );
  AND U16119 ( .A(n12242), .B(n12243), .Z(n12241) );
  NAND U16120 ( .A(o[145]), .B(n11804), .Z(n12243) );
  NANDN U16121 ( .A(n11805), .B(creg[145]), .Z(n12242) );
  NAND U16122 ( .A(n12244), .B(n9647), .Z(n7039) );
  NANDN U16123 ( .A(init), .B(m[146]), .Z(n9647) );
  AND U16124 ( .A(n12245), .B(n12246), .Z(n12244) );
  NAND U16125 ( .A(o[146]), .B(n11804), .Z(n12246) );
  NANDN U16126 ( .A(n11805), .B(creg[146]), .Z(n12245) );
  NAND U16127 ( .A(n12247), .B(n9645), .Z(n7038) );
  NANDN U16128 ( .A(init), .B(m[147]), .Z(n9645) );
  AND U16129 ( .A(n12248), .B(n12249), .Z(n12247) );
  NAND U16130 ( .A(o[147]), .B(n11804), .Z(n12249) );
  NANDN U16131 ( .A(n11805), .B(creg[147]), .Z(n12248) );
  NAND U16132 ( .A(n12250), .B(n9643), .Z(n7037) );
  NANDN U16133 ( .A(init), .B(m[148]), .Z(n9643) );
  AND U16134 ( .A(n12251), .B(n12252), .Z(n12250) );
  NAND U16135 ( .A(o[148]), .B(n11804), .Z(n12252) );
  NANDN U16136 ( .A(n11805), .B(creg[148]), .Z(n12251) );
  NAND U16137 ( .A(n12253), .B(n9641), .Z(n7036) );
  NANDN U16138 ( .A(init), .B(m[149]), .Z(n9641) );
  AND U16139 ( .A(n12254), .B(n12255), .Z(n12253) );
  NAND U16140 ( .A(o[149]), .B(n11804), .Z(n12255) );
  NANDN U16141 ( .A(n11805), .B(creg[149]), .Z(n12254) );
  NAND U16142 ( .A(n12256), .B(n9637), .Z(n7035) );
  NANDN U16143 ( .A(init), .B(m[150]), .Z(n9637) );
  AND U16144 ( .A(n12257), .B(n12258), .Z(n12256) );
  NAND U16145 ( .A(o[150]), .B(n11804), .Z(n12258) );
  NANDN U16146 ( .A(n11805), .B(creg[150]), .Z(n12257) );
  NAND U16147 ( .A(n12259), .B(n9635), .Z(n7034) );
  NANDN U16148 ( .A(init), .B(m[151]), .Z(n9635) );
  AND U16149 ( .A(n12260), .B(n12261), .Z(n12259) );
  NAND U16150 ( .A(o[151]), .B(n11804), .Z(n12261) );
  NANDN U16151 ( .A(n11805), .B(creg[151]), .Z(n12260) );
  NAND U16152 ( .A(n12262), .B(n9633), .Z(n7033) );
  NANDN U16153 ( .A(init), .B(m[152]), .Z(n9633) );
  AND U16154 ( .A(n12263), .B(n12264), .Z(n12262) );
  NAND U16155 ( .A(o[152]), .B(n11804), .Z(n12264) );
  NANDN U16156 ( .A(n11805), .B(creg[152]), .Z(n12263) );
  NAND U16157 ( .A(n12265), .B(n9631), .Z(n7032) );
  NANDN U16158 ( .A(init), .B(m[153]), .Z(n9631) );
  AND U16159 ( .A(n12266), .B(n12267), .Z(n12265) );
  NAND U16160 ( .A(o[153]), .B(n11804), .Z(n12267) );
  NANDN U16161 ( .A(n11805), .B(creg[153]), .Z(n12266) );
  NAND U16162 ( .A(n12268), .B(n9629), .Z(n7031) );
  NANDN U16163 ( .A(init), .B(m[154]), .Z(n9629) );
  AND U16164 ( .A(n12269), .B(n12270), .Z(n12268) );
  NAND U16165 ( .A(o[154]), .B(n11804), .Z(n12270) );
  NANDN U16166 ( .A(n11805), .B(creg[154]), .Z(n12269) );
  NAND U16167 ( .A(n12271), .B(n9627), .Z(n7030) );
  NANDN U16168 ( .A(init), .B(m[155]), .Z(n9627) );
  AND U16169 ( .A(n12272), .B(n12273), .Z(n12271) );
  NAND U16170 ( .A(o[155]), .B(n11804), .Z(n12273) );
  NANDN U16171 ( .A(n11805), .B(creg[155]), .Z(n12272) );
  NAND U16172 ( .A(n12274), .B(n9625), .Z(n7029) );
  NANDN U16173 ( .A(init), .B(m[156]), .Z(n9625) );
  AND U16174 ( .A(n12275), .B(n12276), .Z(n12274) );
  NAND U16175 ( .A(o[156]), .B(n11804), .Z(n12276) );
  NANDN U16176 ( .A(n11805), .B(creg[156]), .Z(n12275) );
  NAND U16177 ( .A(n12277), .B(n9623), .Z(n7028) );
  NANDN U16178 ( .A(init), .B(m[157]), .Z(n9623) );
  AND U16179 ( .A(n12278), .B(n12279), .Z(n12277) );
  NAND U16180 ( .A(o[157]), .B(n11804), .Z(n12279) );
  NANDN U16181 ( .A(n11805), .B(creg[157]), .Z(n12278) );
  NAND U16182 ( .A(n12280), .B(n9621), .Z(n7027) );
  NANDN U16183 ( .A(init), .B(m[158]), .Z(n9621) );
  AND U16184 ( .A(n12281), .B(n12282), .Z(n12280) );
  NAND U16185 ( .A(o[158]), .B(n11804), .Z(n12282) );
  NANDN U16186 ( .A(n11805), .B(creg[158]), .Z(n12281) );
  NAND U16187 ( .A(n12283), .B(n9619), .Z(n7026) );
  NANDN U16188 ( .A(init), .B(m[159]), .Z(n9619) );
  AND U16189 ( .A(n12284), .B(n12285), .Z(n12283) );
  NAND U16190 ( .A(o[159]), .B(n11804), .Z(n12285) );
  NANDN U16191 ( .A(n11805), .B(creg[159]), .Z(n12284) );
  NAND U16192 ( .A(n12286), .B(n9615), .Z(n7025) );
  NANDN U16193 ( .A(init), .B(m[160]), .Z(n9615) );
  AND U16194 ( .A(n12287), .B(n12288), .Z(n12286) );
  NAND U16195 ( .A(o[160]), .B(n11804), .Z(n12288) );
  NANDN U16196 ( .A(n11805), .B(creg[160]), .Z(n12287) );
  NAND U16197 ( .A(n12289), .B(n9613), .Z(n7024) );
  NANDN U16198 ( .A(init), .B(m[161]), .Z(n9613) );
  AND U16199 ( .A(n12290), .B(n12291), .Z(n12289) );
  NAND U16200 ( .A(o[161]), .B(n11804), .Z(n12291) );
  NANDN U16201 ( .A(n11805), .B(creg[161]), .Z(n12290) );
  NAND U16202 ( .A(n12292), .B(n9611), .Z(n7023) );
  NANDN U16203 ( .A(init), .B(m[162]), .Z(n9611) );
  AND U16204 ( .A(n12293), .B(n12294), .Z(n12292) );
  NAND U16205 ( .A(o[162]), .B(n11804), .Z(n12294) );
  NANDN U16206 ( .A(n11805), .B(creg[162]), .Z(n12293) );
  NAND U16207 ( .A(n12295), .B(n9609), .Z(n7022) );
  NANDN U16208 ( .A(init), .B(m[163]), .Z(n9609) );
  AND U16209 ( .A(n12296), .B(n12297), .Z(n12295) );
  NAND U16210 ( .A(o[163]), .B(n11804), .Z(n12297) );
  NANDN U16211 ( .A(n11805), .B(creg[163]), .Z(n12296) );
  NAND U16212 ( .A(n12298), .B(n9607), .Z(n7021) );
  NANDN U16213 ( .A(init), .B(m[164]), .Z(n9607) );
  AND U16214 ( .A(n12299), .B(n12300), .Z(n12298) );
  NAND U16215 ( .A(o[164]), .B(n11804), .Z(n12300) );
  NANDN U16216 ( .A(n11805), .B(creg[164]), .Z(n12299) );
  NAND U16217 ( .A(n12301), .B(n9605), .Z(n7020) );
  NANDN U16218 ( .A(init), .B(m[165]), .Z(n9605) );
  AND U16219 ( .A(n12302), .B(n12303), .Z(n12301) );
  NAND U16220 ( .A(o[165]), .B(n11804), .Z(n12303) );
  NANDN U16221 ( .A(n11805), .B(creg[165]), .Z(n12302) );
  NAND U16222 ( .A(n12304), .B(n9603), .Z(n7019) );
  NANDN U16223 ( .A(init), .B(m[166]), .Z(n9603) );
  AND U16224 ( .A(n12305), .B(n12306), .Z(n12304) );
  NAND U16225 ( .A(o[166]), .B(n11804), .Z(n12306) );
  NANDN U16226 ( .A(n11805), .B(creg[166]), .Z(n12305) );
  NAND U16227 ( .A(n12307), .B(n9601), .Z(n7018) );
  NANDN U16228 ( .A(init), .B(m[167]), .Z(n9601) );
  AND U16229 ( .A(n12308), .B(n12309), .Z(n12307) );
  NAND U16230 ( .A(o[167]), .B(n11804), .Z(n12309) );
  NANDN U16231 ( .A(n11805), .B(creg[167]), .Z(n12308) );
  NAND U16232 ( .A(n12310), .B(n9599), .Z(n7017) );
  NANDN U16233 ( .A(init), .B(m[168]), .Z(n9599) );
  AND U16234 ( .A(n12311), .B(n12312), .Z(n12310) );
  NAND U16235 ( .A(o[168]), .B(n11804), .Z(n12312) );
  NANDN U16236 ( .A(n11805), .B(creg[168]), .Z(n12311) );
  NAND U16237 ( .A(n12313), .B(n9597), .Z(n7016) );
  NANDN U16238 ( .A(init), .B(m[169]), .Z(n9597) );
  AND U16239 ( .A(n12314), .B(n12315), .Z(n12313) );
  NAND U16240 ( .A(o[169]), .B(n11804), .Z(n12315) );
  NANDN U16241 ( .A(n11805), .B(creg[169]), .Z(n12314) );
  NAND U16242 ( .A(n12316), .B(n9593), .Z(n7015) );
  NANDN U16243 ( .A(init), .B(m[170]), .Z(n9593) );
  AND U16244 ( .A(n12317), .B(n12318), .Z(n12316) );
  NAND U16245 ( .A(o[170]), .B(n11804), .Z(n12318) );
  NANDN U16246 ( .A(n11805), .B(creg[170]), .Z(n12317) );
  NAND U16247 ( .A(n12319), .B(n9591), .Z(n7014) );
  NANDN U16248 ( .A(init), .B(m[171]), .Z(n9591) );
  AND U16249 ( .A(n12320), .B(n12321), .Z(n12319) );
  NAND U16250 ( .A(o[171]), .B(n11804), .Z(n12321) );
  NANDN U16251 ( .A(n11805), .B(creg[171]), .Z(n12320) );
  NAND U16252 ( .A(n12322), .B(n9589), .Z(n7013) );
  NANDN U16253 ( .A(init), .B(m[172]), .Z(n9589) );
  AND U16254 ( .A(n12323), .B(n12324), .Z(n12322) );
  NAND U16255 ( .A(o[172]), .B(n11804), .Z(n12324) );
  NANDN U16256 ( .A(n11805), .B(creg[172]), .Z(n12323) );
  NAND U16257 ( .A(n12325), .B(n9587), .Z(n7012) );
  NANDN U16258 ( .A(init), .B(m[173]), .Z(n9587) );
  AND U16259 ( .A(n12326), .B(n12327), .Z(n12325) );
  NAND U16260 ( .A(o[173]), .B(n11804), .Z(n12327) );
  NANDN U16261 ( .A(n11805), .B(creg[173]), .Z(n12326) );
  NAND U16262 ( .A(n12328), .B(n9585), .Z(n7011) );
  NANDN U16263 ( .A(init), .B(m[174]), .Z(n9585) );
  AND U16264 ( .A(n12329), .B(n12330), .Z(n12328) );
  NAND U16265 ( .A(o[174]), .B(n11804), .Z(n12330) );
  NANDN U16266 ( .A(n11805), .B(creg[174]), .Z(n12329) );
  NAND U16267 ( .A(n12331), .B(n9583), .Z(n7010) );
  NANDN U16268 ( .A(init), .B(m[175]), .Z(n9583) );
  AND U16269 ( .A(n12332), .B(n12333), .Z(n12331) );
  NAND U16270 ( .A(o[175]), .B(n11804), .Z(n12333) );
  NANDN U16271 ( .A(n11805), .B(creg[175]), .Z(n12332) );
  NAND U16272 ( .A(n12334), .B(n9581), .Z(n7009) );
  NANDN U16273 ( .A(init), .B(m[176]), .Z(n9581) );
  AND U16274 ( .A(n12335), .B(n12336), .Z(n12334) );
  NAND U16275 ( .A(o[176]), .B(n11804), .Z(n12336) );
  NANDN U16276 ( .A(n11805), .B(creg[176]), .Z(n12335) );
  NAND U16277 ( .A(n12337), .B(n9579), .Z(n7008) );
  NANDN U16278 ( .A(init), .B(m[177]), .Z(n9579) );
  AND U16279 ( .A(n12338), .B(n12339), .Z(n12337) );
  NAND U16280 ( .A(o[177]), .B(n11804), .Z(n12339) );
  NANDN U16281 ( .A(n11805), .B(creg[177]), .Z(n12338) );
  NAND U16282 ( .A(n12340), .B(n9577), .Z(n7007) );
  NANDN U16283 ( .A(init), .B(m[178]), .Z(n9577) );
  AND U16284 ( .A(n12341), .B(n12342), .Z(n12340) );
  NAND U16285 ( .A(o[178]), .B(n11804), .Z(n12342) );
  NANDN U16286 ( .A(n11805), .B(creg[178]), .Z(n12341) );
  NAND U16287 ( .A(n12343), .B(n9575), .Z(n7006) );
  NANDN U16288 ( .A(init), .B(m[179]), .Z(n9575) );
  AND U16289 ( .A(n12344), .B(n12345), .Z(n12343) );
  NAND U16290 ( .A(o[179]), .B(n11804), .Z(n12345) );
  NANDN U16291 ( .A(n11805), .B(creg[179]), .Z(n12344) );
  NAND U16292 ( .A(n12346), .B(n9571), .Z(n7005) );
  NANDN U16293 ( .A(init), .B(m[180]), .Z(n9571) );
  AND U16294 ( .A(n12347), .B(n12348), .Z(n12346) );
  NAND U16295 ( .A(o[180]), .B(n11804), .Z(n12348) );
  NANDN U16296 ( .A(n11805), .B(creg[180]), .Z(n12347) );
  NAND U16297 ( .A(n12349), .B(n9569), .Z(n7004) );
  NANDN U16298 ( .A(init), .B(m[181]), .Z(n9569) );
  AND U16299 ( .A(n12350), .B(n12351), .Z(n12349) );
  NAND U16300 ( .A(o[181]), .B(n11804), .Z(n12351) );
  NANDN U16301 ( .A(n11805), .B(creg[181]), .Z(n12350) );
  NAND U16302 ( .A(n12352), .B(n9567), .Z(n7003) );
  NANDN U16303 ( .A(init), .B(m[182]), .Z(n9567) );
  AND U16304 ( .A(n12353), .B(n12354), .Z(n12352) );
  NAND U16305 ( .A(o[182]), .B(n11804), .Z(n12354) );
  NANDN U16306 ( .A(n11805), .B(creg[182]), .Z(n12353) );
  NAND U16307 ( .A(n12355), .B(n9565), .Z(n7002) );
  NANDN U16308 ( .A(init), .B(m[183]), .Z(n9565) );
  AND U16309 ( .A(n12356), .B(n12357), .Z(n12355) );
  NAND U16310 ( .A(o[183]), .B(n11804), .Z(n12357) );
  NANDN U16311 ( .A(n11805), .B(creg[183]), .Z(n12356) );
  NAND U16312 ( .A(n12358), .B(n9563), .Z(n7001) );
  NANDN U16313 ( .A(init), .B(m[184]), .Z(n9563) );
  AND U16314 ( .A(n12359), .B(n12360), .Z(n12358) );
  NAND U16315 ( .A(o[184]), .B(n11804), .Z(n12360) );
  NANDN U16316 ( .A(n11805), .B(creg[184]), .Z(n12359) );
  NAND U16317 ( .A(n12361), .B(n9561), .Z(n7000) );
  NANDN U16318 ( .A(init), .B(m[185]), .Z(n9561) );
  AND U16319 ( .A(n12362), .B(n12363), .Z(n12361) );
  NAND U16320 ( .A(o[185]), .B(n11804), .Z(n12363) );
  NANDN U16321 ( .A(n11805), .B(creg[185]), .Z(n12362) );
  NAND U16322 ( .A(n12364), .B(n9559), .Z(n6999) );
  NANDN U16323 ( .A(init), .B(m[186]), .Z(n9559) );
  AND U16324 ( .A(n12365), .B(n12366), .Z(n12364) );
  NAND U16325 ( .A(o[186]), .B(n11804), .Z(n12366) );
  NANDN U16326 ( .A(n11805), .B(creg[186]), .Z(n12365) );
  NAND U16327 ( .A(n12367), .B(n9557), .Z(n6998) );
  NANDN U16328 ( .A(init), .B(m[187]), .Z(n9557) );
  AND U16329 ( .A(n12368), .B(n12369), .Z(n12367) );
  NAND U16330 ( .A(o[187]), .B(n11804), .Z(n12369) );
  NANDN U16331 ( .A(n11805), .B(creg[187]), .Z(n12368) );
  NAND U16332 ( .A(n12370), .B(n9555), .Z(n6997) );
  NANDN U16333 ( .A(init), .B(m[188]), .Z(n9555) );
  AND U16334 ( .A(n12371), .B(n12372), .Z(n12370) );
  NAND U16335 ( .A(o[188]), .B(n11804), .Z(n12372) );
  NANDN U16336 ( .A(n11805), .B(creg[188]), .Z(n12371) );
  NAND U16337 ( .A(n12373), .B(n9553), .Z(n6996) );
  NANDN U16338 ( .A(init), .B(m[189]), .Z(n9553) );
  AND U16339 ( .A(n12374), .B(n12375), .Z(n12373) );
  NAND U16340 ( .A(o[189]), .B(n11804), .Z(n12375) );
  NANDN U16341 ( .A(n11805), .B(creg[189]), .Z(n12374) );
  NAND U16342 ( .A(n12376), .B(n9549), .Z(n6995) );
  NANDN U16343 ( .A(init), .B(m[190]), .Z(n9549) );
  AND U16344 ( .A(n12377), .B(n12378), .Z(n12376) );
  NAND U16345 ( .A(o[190]), .B(n11804), .Z(n12378) );
  NANDN U16346 ( .A(n11805), .B(creg[190]), .Z(n12377) );
  NAND U16347 ( .A(n12379), .B(n9547), .Z(n6994) );
  NANDN U16348 ( .A(init), .B(m[191]), .Z(n9547) );
  AND U16349 ( .A(n12380), .B(n12381), .Z(n12379) );
  NAND U16350 ( .A(o[191]), .B(n11804), .Z(n12381) );
  NANDN U16351 ( .A(n11805), .B(creg[191]), .Z(n12380) );
  NAND U16352 ( .A(n12382), .B(n9545), .Z(n6993) );
  NANDN U16353 ( .A(init), .B(m[192]), .Z(n9545) );
  AND U16354 ( .A(n12383), .B(n12384), .Z(n12382) );
  NAND U16355 ( .A(o[192]), .B(n11804), .Z(n12384) );
  NANDN U16356 ( .A(n11805), .B(creg[192]), .Z(n12383) );
  NAND U16357 ( .A(n12385), .B(n9543), .Z(n6992) );
  NANDN U16358 ( .A(init), .B(m[193]), .Z(n9543) );
  AND U16359 ( .A(n12386), .B(n12387), .Z(n12385) );
  NAND U16360 ( .A(o[193]), .B(n11804), .Z(n12387) );
  NANDN U16361 ( .A(n11805), .B(creg[193]), .Z(n12386) );
  NAND U16362 ( .A(n12388), .B(n9541), .Z(n6991) );
  NANDN U16363 ( .A(init), .B(m[194]), .Z(n9541) );
  AND U16364 ( .A(n12389), .B(n12390), .Z(n12388) );
  NAND U16365 ( .A(o[194]), .B(n11804), .Z(n12390) );
  NANDN U16366 ( .A(n11805), .B(creg[194]), .Z(n12389) );
  NAND U16367 ( .A(n12391), .B(n9539), .Z(n6990) );
  NANDN U16368 ( .A(init), .B(m[195]), .Z(n9539) );
  AND U16369 ( .A(n12392), .B(n12393), .Z(n12391) );
  NAND U16370 ( .A(o[195]), .B(n11804), .Z(n12393) );
  NANDN U16371 ( .A(n11805), .B(creg[195]), .Z(n12392) );
  NAND U16372 ( .A(n12394), .B(n9537), .Z(n6989) );
  NANDN U16373 ( .A(init), .B(m[196]), .Z(n9537) );
  AND U16374 ( .A(n12395), .B(n12396), .Z(n12394) );
  NAND U16375 ( .A(o[196]), .B(n11804), .Z(n12396) );
  NANDN U16376 ( .A(n11805), .B(creg[196]), .Z(n12395) );
  NAND U16377 ( .A(n12397), .B(n9535), .Z(n6988) );
  NANDN U16378 ( .A(init), .B(m[197]), .Z(n9535) );
  AND U16379 ( .A(n12398), .B(n12399), .Z(n12397) );
  NAND U16380 ( .A(o[197]), .B(n11804), .Z(n12399) );
  NANDN U16381 ( .A(n11805), .B(creg[197]), .Z(n12398) );
  NAND U16382 ( .A(n12400), .B(n9533), .Z(n6987) );
  NANDN U16383 ( .A(init), .B(m[198]), .Z(n9533) );
  AND U16384 ( .A(n12401), .B(n12402), .Z(n12400) );
  NAND U16385 ( .A(o[198]), .B(n11804), .Z(n12402) );
  NANDN U16386 ( .A(n11805), .B(creg[198]), .Z(n12401) );
  NAND U16387 ( .A(n12403), .B(n9531), .Z(n6986) );
  NANDN U16388 ( .A(init), .B(m[199]), .Z(n9531) );
  AND U16389 ( .A(n12404), .B(n12405), .Z(n12403) );
  NAND U16390 ( .A(o[199]), .B(n11804), .Z(n12405) );
  NANDN U16391 ( .A(n11805), .B(creg[199]), .Z(n12404) );
  NAND U16392 ( .A(n12406), .B(n9525), .Z(n6985) );
  NANDN U16393 ( .A(init), .B(m[200]), .Z(n9525) );
  AND U16394 ( .A(n12407), .B(n12408), .Z(n12406) );
  NAND U16395 ( .A(o[200]), .B(n11804), .Z(n12408) );
  NANDN U16396 ( .A(n11805), .B(creg[200]), .Z(n12407) );
  NAND U16397 ( .A(n12409), .B(n9523), .Z(n6984) );
  NANDN U16398 ( .A(init), .B(m[201]), .Z(n9523) );
  AND U16399 ( .A(n12410), .B(n12411), .Z(n12409) );
  NAND U16400 ( .A(o[201]), .B(n11804), .Z(n12411) );
  NANDN U16401 ( .A(n11805), .B(creg[201]), .Z(n12410) );
  NAND U16402 ( .A(n12412), .B(n9521), .Z(n6983) );
  NANDN U16403 ( .A(init), .B(m[202]), .Z(n9521) );
  AND U16404 ( .A(n12413), .B(n12414), .Z(n12412) );
  NAND U16405 ( .A(o[202]), .B(n11804), .Z(n12414) );
  NANDN U16406 ( .A(n11805), .B(creg[202]), .Z(n12413) );
  NAND U16407 ( .A(n12415), .B(n9519), .Z(n6982) );
  NANDN U16408 ( .A(init), .B(m[203]), .Z(n9519) );
  AND U16409 ( .A(n12416), .B(n12417), .Z(n12415) );
  NAND U16410 ( .A(o[203]), .B(n11804), .Z(n12417) );
  NANDN U16411 ( .A(n11805), .B(creg[203]), .Z(n12416) );
  NAND U16412 ( .A(n12418), .B(n9517), .Z(n6981) );
  NANDN U16413 ( .A(init), .B(m[204]), .Z(n9517) );
  AND U16414 ( .A(n12419), .B(n12420), .Z(n12418) );
  NAND U16415 ( .A(o[204]), .B(n11804), .Z(n12420) );
  NANDN U16416 ( .A(n11805), .B(creg[204]), .Z(n12419) );
  NAND U16417 ( .A(n12421), .B(n9515), .Z(n6980) );
  NANDN U16418 ( .A(init), .B(m[205]), .Z(n9515) );
  AND U16419 ( .A(n12422), .B(n12423), .Z(n12421) );
  NAND U16420 ( .A(o[205]), .B(n11804), .Z(n12423) );
  NANDN U16421 ( .A(n11805), .B(creg[205]), .Z(n12422) );
  NAND U16422 ( .A(n12424), .B(n9513), .Z(n6979) );
  NANDN U16423 ( .A(init), .B(m[206]), .Z(n9513) );
  AND U16424 ( .A(n12425), .B(n12426), .Z(n12424) );
  NAND U16425 ( .A(o[206]), .B(n11804), .Z(n12426) );
  NANDN U16426 ( .A(n11805), .B(creg[206]), .Z(n12425) );
  NAND U16427 ( .A(n12427), .B(n9511), .Z(n6978) );
  NANDN U16428 ( .A(init), .B(m[207]), .Z(n9511) );
  AND U16429 ( .A(n12428), .B(n12429), .Z(n12427) );
  NAND U16430 ( .A(o[207]), .B(n11804), .Z(n12429) );
  NANDN U16431 ( .A(n11805), .B(creg[207]), .Z(n12428) );
  NAND U16432 ( .A(n12430), .B(n9509), .Z(n6977) );
  NANDN U16433 ( .A(init), .B(m[208]), .Z(n9509) );
  AND U16434 ( .A(n12431), .B(n12432), .Z(n12430) );
  NAND U16435 ( .A(o[208]), .B(n11804), .Z(n12432) );
  NANDN U16436 ( .A(n11805), .B(creg[208]), .Z(n12431) );
  NAND U16437 ( .A(n12433), .B(n9507), .Z(n6976) );
  NANDN U16438 ( .A(init), .B(m[209]), .Z(n9507) );
  AND U16439 ( .A(n12434), .B(n12435), .Z(n12433) );
  NAND U16440 ( .A(o[209]), .B(n11804), .Z(n12435) );
  NANDN U16441 ( .A(n11805), .B(creg[209]), .Z(n12434) );
  NAND U16442 ( .A(n12436), .B(n9503), .Z(n6975) );
  NANDN U16443 ( .A(init), .B(m[210]), .Z(n9503) );
  AND U16444 ( .A(n12437), .B(n12438), .Z(n12436) );
  NAND U16445 ( .A(o[210]), .B(n11804), .Z(n12438) );
  NANDN U16446 ( .A(n11805), .B(creg[210]), .Z(n12437) );
  NAND U16447 ( .A(n12439), .B(n9501), .Z(n6974) );
  NANDN U16448 ( .A(init), .B(m[211]), .Z(n9501) );
  AND U16449 ( .A(n12440), .B(n12441), .Z(n12439) );
  NAND U16450 ( .A(o[211]), .B(n11804), .Z(n12441) );
  NANDN U16451 ( .A(n11805), .B(creg[211]), .Z(n12440) );
  NAND U16452 ( .A(n12442), .B(n9499), .Z(n6973) );
  NANDN U16453 ( .A(init), .B(m[212]), .Z(n9499) );
  AND U16454 ( .A(n12443), .B(n12444), .Z(n12442) );
  NAND U16455 ( .A(o[212]), .B(n11804), .Z(n12444) );
  NANDN U16456 ( .A(n11805), .B(creg[212]), .Z(n12443) );
  NAND U16457 ( .A(n12445), .B(n9497), .Z(n6972) );
  NANDN U16458 ( .A(init), .B(m[213]), .Z(n9497) );
  AND U16459 ( .A(n12446), .B(n12447), .Z(n12445) );
  NAND U16460 ( .A(o[213]), .B(n11804), .Z(n12447) );
  NANDN U16461 ( .A(n11805), .B(creg[213]), .Z(n12446) );
  NAND U16462 ( .A(n12448), .B(n9495), .Z(n6971) );
  NANDN U16463 ( .A(init), .B(m[214]), .Z(n9495) );
  AND U16464 ( .A(n12449), .B(n12450), .Z(n12448) );
  NAND U16465 ( .A(o[214]), .B(n11804), .Z(n12450) );
  NANDN U16466 ( .A(n11805), .B(creg[214]), .Z(n12449) );
  NAND U16467 ( .A(n12451), .B(n9493), .Z(n6970) );
  NANDN U16468 ( .A(init), .B(m[215]), .Z(n9493) );
  AND U16469 ( .A(n12452), .B(n12453), .Z(n12451) );
  NAND U16470 ( .A(o[215]), .B(n11804), .Z(n12453) );
  NANDN U16471 ( .A(n11805), .B(creg[215]), .Z(n12452) );
  NAND U16472 ( .A(n12454), .B(n9491), .Z(n6969) );
  NANDN U16473 ( .A(init), .B(m[216]), .Z(n9491) );
  AND U16474 ( .A(n12455), .B(n12456), .Z(n12454) );
  NAND U16475 ( .A(o[216]), .B(n11804), .Z(n12456) );
  NANDN U16476 ( .A(n11805), .B(creg[216]), .Z(n12455) );
  NAND U16477 ( .A(n12457), .B(n9489), .Z(n6968) );
  NANDN U16478 ( .A(init), .B(m[217]), .Z(n9489) );
  AND U16479 ( .A(n12458), .B(n12459), .Z(n12457) );
  NAND U16480 ( .A(o[217]), .B(n11804), .Z(n12459) );
  NANDN U16481 ( .A(n11805), .B(creg[217]), .Z(n12458) );
  NAND U16482 ( .A(n12460), .B(n9487), .Z(n6967) );
  NANDN U16483 ( .A(init), .B(m[218]), .Z(n9487) );
  AND U16484 ( .A(n12461), .B(n12462), .Z(n12460) );
  NAND U16485 ( .A(o[218]), .B(n11804), .Z(n12462) );
  NANDN U16486 ( .A(n11805), .B(creg[218]), .Z(n12461) );
  NAND U16487 ( .A(n12463), .B(n9485), .Z(n6966) );
  NANDN U16488 ( .A(init), .B(m[219]), .Z(n9485) );
  AND U16489 ( .A(n12464), .B(n12465), .Z(n12463) );
  NAND U16490 ( .A(o[219]), .B(n11804), .Z(n12465) );
  NANDN U16491 ( .A(n11805), .B(creg[219]), .Z(n12464) );
  NAND U16492 ( .A(n12466), .B(n9481), .Z(n6965) );
  NANDN U16493 ( .A(init), .B(m[220]), .Z(n9481) );
  AND U16494 ( .A(n12467), .B(n12468), .Z(n12466) );
  NAND U16495 ( .A(o[220]), .B(n11804), .Z(n12468) );
  NANDN U16496 ( .A(n11805), .B(creg[220]), .Z(n12467) );
  NAND U16497 ( .A(n12469), .B(n9479), .Z(n6964) );
  NANDN U16498 ( .A(init), .B(m[221]), .Z(n9479) );
  AND U16499 ( .A(n12470), .B(n12471), .Z(n12469) );
  NAND U16500 ( .A(o[221]), .B(n11804), .Z(n12471) );
  NANDN U16501 ( .A(n11805), .B(creg[221]), .Z(n12470) );
  NAND U16502 ( .A(n12472), .B(n9477), .Z(n6963) );
  NANDN U16503 ( .A(init), .B(m[222]), .Z(n9477) );
  AND U16504 ( .A(n12473), .B(n12474), .Z(n12472) );
  NAND U16505 ( .A(o[222]), .B(n11804), .Z(n12474) );
  NANDN U16506 ( .A(n11805), .B(creg[222]), .Z(n12473) );
  NAND U16507 ( .A(n12475), .B(n9475), .Z(n6962) );
  NANDN U16508 ( .A(init), .B(m[223]), .Z(n9475) );
  AND U16509 ( .A(n12476), .B(n12477), .Z(n12475) );
  NAND U16510 ( .A(o[223]), .B(n11804), .Z(n12477) );
  NANDN U16511 ( .A(n11805), .B(creg[223]), .Z(n12476) );
  NAND U16512 ( .A(n12478), .B(n9473), .Z(n6961) );
  NANDN U16513 ( .A(init), .B(m[224]), .Z(n9473) );
  AND U16514 ( .A(n12479), .B(n12480), .Z(n12478) );
  NAND U16515 ( .A(o[224]), .B(n11804), .Z(n12480) );
  NANDN U16516 ( .A(n11805), .B(creg[224]), .Z(n12479) );
  NAND U16517 ( .A(n12481), .B(n9471), .Z(n6960) );
  NANDN U16518 ( .A(init), .B(m[225]), .Z(n9471) );
  AND U16519 ( .A(n12482), .B(n12483), .Z(n12481) );
  NAND U16520 ( .A(o[225]), .B(n11804), .Z(n12483) );
  NANDN U16521 ( .A(n11805), .B(creg[225]), .Z(n12482) );
  NAND U16522 ( .A(n12484), .B(n9469), .Z(n6959) );
  NANDN U16523 ( .A(init), .B(m[226]), .Z(n9469) );
  AND U16524 ( .A(n12485), .B(n12486), .Z(n12484) );
  NAND U16525 ( .A(o[226]), .B(n11804), .Z(n12486) );
  NANDN U16526 ( .A(n11805), .B(creg[226]), .Z(n12485) );
  NAND U16527 ( .A(n12487), .B(n9467), .Z(n6958) );
  NANDN U16528 ( .A(init), .B(m[227]), .Z(n9467) );
  AND U16529 ( .A(n12488), .B(n12489), .Z(n12487) );
  NAND U16530 ( .A(o[227]), .B(n11804), .Z(n12489) );
  NANDN U16531 ( .A(n11805), .B(creg[227]), .Z(n12488) );
  NAND U16532 ( .A(n12490), .B(n9465), .Z(n6957) );
  NANDN U16533 ( .A(init), .B(m[228]), .Z(n9465) );
  AND U16534 ( .A(n12491), .B(n12492), .Z(n12490) );
  NAND U16535 ( .A(o[228]), .B(n11804), .Z(n12492) );
  NANDN U16536 ( .A(n11805), .B(creg[228]), .Z(n12491) );
  NAND U16537 ( .A(n12493), .B(n9463), .Z(n6956) );
  NANDN U16538 ( .A(init), .B(m[229]), .Z(n9463) );
  AND U16539 ( .A(n12494), .B(n12495), .Z(n12493) );
  NAND U16540 ( .A(o[229]), .B(n11804), .Z(n12495) );
  NANDN U16541 ( .A(n11805), .B(creg[229]), .Z(n12494) );
  NAND U16542 ( .A(n12496), .B(n9459), .Z(n6955) );
  NANDN U16543 ( .A(init), .B(m[230]), .Z(n9459) );
  AND U16544 ( .A(n12497), .B(n12498), .Z(n12496) );
  NAND U16545 ( .A(o[230]), .B(n11804), .Z(n12498) );
  NANDN U16546 ( .A(n11805), .B(creg[230]), .Z(n12497) );
  NAND U16547 ( .A(n12499), .B(n9457), .Z(n6954) );
  NANDN U16548 ( .A(init), .B(m[231]), .Z(n9457) );
  AND U16549 ( .A(n12500), .B(n12501), .Z(n12499) );
  NAND U16550 ( .A(o[231]), .B(n11804), .Z(n12501) );
  NANDN U16551 ( .A(n11805), .B(creg[231]), .Z(n12500) );
  NAND U16552 ( .A(n12502), .B(n9455), .Z(n6953) );
  NANDN U16553 ( .A(init), .B(m[232]), .Z(n9455) );
  AND U16554 ( .A(n12503), .B(n12504), .Z(n12502) );
  NAND U16555 ( .A(o[232]), .B(n11804), .Z(n12504) );
  NANDN U16556 ( .A(n11805), .B(creg[232]), .Z(n12503) );
  NAND U16557 ( .A(n12505), .B(n9453), .Z(n6952) );
  NANDN U16558 ( .A(init), .B(m[233]), .Z(n9453) );
  AND U16559 ( .A(n12506), .B(n12507), .Z(n12505) );
  NAND U16560 ( .A(o[233]), .B(n11804), .Z(n12507) );
  NANDN U16561 ( .A(n11805), .B(creg[233]), .Z(n12506) );
  NAND U16562 ( .A(n12508), .B(n9451), .Z(n6951) );
  NANDN U16563 ( .A(init), .B(m[234]), .Z(n9451) );
  AND U16564 ( .A(n12509), .B(n12510), .Z(n12508) );
  NAND U16565 ( .A(o[234]), .B(n11804), .Z(n12510) );
  NANDN U16566 ( .A(n11805), .B(creg[234]), .Z(n12509) );
  NAND U16567 ( .A(n12511), .B(n9449), .Z(n6950) );
  NANDN U16568 ( .A(init), .B(m[235]), .Z(n9449) );
  AND U16569 ( .A(n12512), .B(n12513), .Z(n12511) );
  NAND U16570 ( .A(o[235]), .B(n11804), .Z(n12513) );
  NANDN U16571 ( .A(n11805), .B(creg[235]), .Z(n12512) );
  NAND U16572 ( .A(n12514), .B(n9447), .Z(n6949) );
  NANDN U16573 ( .A(init), .B(m[236]), .Z(n9447) );
  AND U16574 ( .A(n12515), .B(n12516), .Z(n12514) );
  NAND U16575 ( .A(o[236]), .B(n11804), .Z(n12516) );
  NANDN U16576 ( .A(n11805), .B(creg[236]), .Z(n12515) );
  NAND U16577 ( .A(n12517), .B(n9445), .Z(n6948) );
  NANDN U16578 ( .A(init), .B(m[237]), .Z(n9445) );
  AND U16579 ( .A(n12518), .B(n12519), .Z(n12517) );
  NAND U16580 ( .A(o[237]), .B(n11804), .Z(n12519) );
  NANDN U16581 ( .A(n11805), .B(creg[237]), .Z(n12518) );
  NAND U16582 ( .A(n12520), .B(n9443), .Z(n6947) );
  NANDN U16583 ( .A(init), .B(m[238]), .Z(n9443) );
  AND U16584 ( .A(n12521), .B(n12522), .Z(n12520) );
  NAND U16585 ( .A(o[238]), .B(n11804), .Z(n12522) );
  NANDN U16586 ( .A(n11805), .B(creg[238]), .Z(n12521) );
  NAND U16587 ( .A(n12523), .B(n9441), .Z(n6946) );
  NANDN U16588 ( .A(init), .B(m[239]), .Z(n9441) );
  AND U16589 ( .A(n12524), .B(n12525), .Z(n12523) );
  NAND U16590 ( .A(o[239]), .B(n11804), .Z(n12525) );
  NANDN U16591 ( .A(n11805), .B(creg[239]), .Z(n12524) );
  NAND U16592 ( .A(n12526), .B(n9437), .Z(n6945) );
  NANDN U16593 ( .A(init), .B(m[240]), .Z(n9437) );
  AND U16594 ( .A(n12527), .B(n12528), .Z(n12526) );
  NAND U16595 ( .A(o[240]), .B(n11804), .Z(n12528) );
  NANDN U16596 ( .A(n11805), .B(creg[240]), .Z(n12527) );
  NAND U16597 ( .A(n12529), .B(n9435), .Z(n6944) );
  NANDN U16598 ( .A(init), .B(m[241]), .Z(n9435) );
  AND U16599 ( .A(n12530), .B(n12531), .Z(n12529) );
  NAND U16600 ( .A(o[241]), .B(n11804), .Z(n12531) );
  NANDN U16601 ( .A(n11805), .B(creg[241]), .Z(n12530) );
  NAND U16602 ( .A(n12532), .B(n9433), .Z(n6943) );
  NANDN U16603 ( .A(init), .B(m[242]), .Z(n9433) );
  AND U16604 ( .A(n12533), .B(n12534), .Z(n12532) );
  NAND U16605 ( .A(o[242]), .B(n11804), .Z(n12534) );
  NANDN U16606 ( .A(n11805), .B(creg[242]), .Z(n12533) );
  NAND U16607 ( .A(n12535), .B(n9431), .Z(n6942) );
  NANDN U16608 ( .A(init), .B(m[243]), .Z(n9431) );
  AND U16609 ( .A(n12536), .B(n12537), .Z(n12535) );
  NAND U16610 ( .A(o[243]), .B(n11804), .Z(n12537) );
  NANDN U16611 ( .A(n11805), .B(creg[243]), .Z(n12536) );
  NAND U16612 ( .A(n12538), .B(n9429), .Z(n6941) );
  NANDN U16613 ( .A(init), .B(m[244]), .Z(n9429) );
  AND U16614 ( .A(n12539), .B(n12540), .Z(n12538) );
  NAND U16615 ( .A(o[244]), .B(n11804), .Z(n12540) );
  NANDN U16616 ( .A(n11805), .B(creg[244]), .Z(n12539) );
  NAND U16617 ( .A(n12541), .B(n9427), .Z(n6940) );
  NANDN U16618 ( .A(init), .B(m[245]), .Z(n9427) );
  AND U16619 ( .A(n12542), .B(n12543), .Z(n12541) );
  NAND U16620 ( .A(o[245]), .B(n11804), .Z(n12543) );
  NANDN U16621 ( .A(n11805), .B(creg[245]), .Z(n12542) );
  NAND U16622 ( .A(n12544), .B(n9425), .Z(n6939) );
  NANDN U16623 ( .A(init), .B(m[246]), .Z(n9425) );
  AND U16624 ( .A(n12545), .B(n12546), .Z(n12544) );
  NAND U16625 ( .A(o[246]), .B(n11804), .Z(n12546) );
  NANDN U16626 ( .A(n11805), .B(creg[246]), .Z(n12545) );
  NAND U16627 ( .A(n12547), .B(n9423), .Z(n6938) );
  NANDN U16628 ( .A(init), .B(m[247]), .Z(n9423) );
  AND U16629 ( .A(n12548), .B(n12549), .Z(n12547) );
  NAND U16630 ( .A(o[247]), .B(n11804), .Z(n12549) );
  NANDN U16631 ( .A(n11805), .B(creg[247]), .Z(n12548) );
  NAND U16632 ( .A(n12550), .B(n9421), .Z(n6937) );
  NANDN U16633 ( .A(init), .B(m[248]), .Z(n9421) );
  AND U16634 ( .A(n12551), .B(n12552), .Z(n12550) );
  NAND U16635 ( .A(o[248]), .B(n11804), .Z(n12552) );
  NANDN U16636 ( .A(n11805), .B(creg[248]), .Z(n12551) );
  NAND U16637 ( .A(n12553), .B(n9419), .Z(n6936) );
  NANDN U16638 ( .A(init), .B(m[249]), .Z(n9419) );
  AND U16639 ( .A(n12554), .B(n12555), .Z(n12553) );
  NAND U16640 ( .A(o[249]), .B(n11804), .Z(n12555) );
  NANDN U16641 ( .A(n11805), .B(creg[249]), .Z(n12554) );
  NAND U16642 ( .A(n12556), .B(n9415), .Z(n6935) );
  NANDN U16643 ( .A(init), .B(m[250]), .Z(n9415) );
  AND U16644 ( .A(n12557), .B(n12558), .Z(n12556) );
  NAND U16645 ( .A(o[250]), .B(n11804), .Z(n12558) );
  NANDN U16646 ( .A(n11805), .B(creg[250]), .Z(n12557) );
  NAND U16647 ( .A(n12559), .B(n9413), .Z(n6934) );
  NANDN U16648 ( .A(init), .B(m[251]), .Z(n9413) );
  AND U16649 ( .A(n12560), .B(n12561), .Z(n12559) );
  NAND U16650 ( .A(o[251]), .B(n11804), .Z(n12561) );
  NANDN U16651 ( .A(n11805), .B(creg[251]), .Z(n12560) );
  NAND U16652 ( .A(n12562), .B(n9411), .Z(n6933) );
  NANDN U16653 ( .A(init), .B(m[252]), .Z(n9411) );
  AND U16654 ( .A(n12563), .B(n12564), .Z(n12562) );
  NAND U16655 ( .A(o[252]), .B(n11804), .Z(n12564) );
  NANDN U16656 ( .A(n11805), .B(creg[252]), .Z(n12563) );
  NAND U16657 ( .A(n12565), .B(n9409), .Z(n6932) );
  NANDN U16658 ( .A(init), .B(m[253]), .Z(n9409) );
  AND U16659 ( .A(n12566), .B(n12567), .Z(n12565) );
  NAND U16660 ( .A(o[253]), .B(n11804), .Z(n12567) );
  NANDN U16661 ( .A(n11805), .B(creg[253]), .Z(n12566) );
  NAND U16662 ( .A(n12568), .B(n9407), .Z(n6931) );
  NANDN U16663 ( .A(init), .B(m[254]), .Z(n9407) );
  AND U16664 ( .A(n12569), .B(n12570), .Z(n12568) );
  NAND U16665 ( .A(o[254]), .B(n11804), .Z(n12570) );
  NANDN U16666 ( .A(n11805), .B(creg[254]), .Z(n12569) );
  NAND U16667 ( .A(n12571), .B(n9405), .Z(n6930) );
  NANDN U16668 ( .A(init), .B(m[255]), .Z(n9405) );
  AND U16669 ( .A(n12572), .B(n12573), .Z(n12571) );
  NAND U16670 ( .A(o[255]), .B(n11804), .Z(n12573) );
  NANDN U16671 ( .A(n11805), .B(creg[255]), .Z(n12572) );
  NAND U16672 ( .A(n12574), .B(n9403), .Z(n6929) );
  NANDN U16673 ( .A(init), .B(m[256]), .Z(n9403) );
  AND U16674 ( .A(n12575), .B(n12576), .Z(n12574) );
  NAND U16675 ( .A(o[256]), .B(n11804), .Z(n12576) );
  NANDN U16676 ( .A(n11805), .B(creg[256]), .Z(n12575) );
  NAND U16677 ( .A(n12577), .B(n9401), .Z(n6928) );
  NANDN U16678 ( .A(init), .B(m[257]), .Z(n9401) );
  AND U16679 ( .A(n12578), .B(n12579), .Z(n12577) );
  NAND U16680 ( .A(o[257]), .B(n11804), .Z(n12579) );
  NANDN U16681 ( .A(n11805), .B(creg[257]), .Z(n12578) );
  NAND U16682 ( .A(n12580), .B(n9399), .Z(n6927) );
  NANDN U16683 ( .A(init), .B(m[258]), .Z(n9399) );
  AND U16684 ( .A(n12581), .B(n12582), .Z(n12580) );
  NAND U16685 ( .A(o[258]), .B(n11804), .Z(n12582) );
  NANDN U16686 ( .A(n11805), .B(creg[258]), .Z(n12581) );
  NAND U16687 ( .A(n12583), .B(n9397), .Z(n6926) );
  NANDN U16688 ( .A(init), .B(m[259]), .Z(n9397) );
  AND U16689 ( .A(n12584), .B(n12585), .Z(n12583) );
  NAND U16690 ( .A(o[259]), .B(n11804), .Z(n12585) );
  NANDN U16691 ( .A(n11805), .B(creg[259]), .Z(n12584) );
  NAND U16692 ( .A(n12586), .B(n9393), .Z(n6925) );
  NANDN U16693 ( .A(init), .B(m[260]), .Z(n9393) );
  AND U16694 ( .A(n12587), .B(n12588), .Z(n12586) );
  NAND U16695 ( .A(o[260]), .B(n11804), .Z(n12588) );
  NANDN U16696 ( .A(n11805), .B(creg[260]), .Z(n12587) );
  NAND U16697 ( .A(n12589), .B(n9391), .Z(n6924) );
  NANDN U16698 ( .A(init), .B(m[261]), .Z(n9391) );
  AND U16699 ( .A(n12590), .B(n12591), .Z(n12589) );
  NAND U16700 ( .A(o[261]), .B(n11804), .Z(n12591) );
  NANDN U16701 ( .A(n11805), .B(creg[261]), .Z(n12590) );
  NAND U16702 ( .A(n12592), .B(n9389), .Z(n6923) );
  NANDN U16703 ( .A(init), .B(m[262]), .Z(n9389) );
  AND U16704 ( .A(n12593), .B(n12594), .Z(n12592) );
  NAND U16705 ( .A(o[262]), .B(n11804), .Z(n12594) );
  NANDN U16706 ( .A(n11805), .B(creg[262]), .Z(n12593) );
  NAND U16707 ( .A(n12595), .B(n9387), .Z(n6922) );
  NANDN U16708 ( .A(init), .B(m[263]), .Z(n9387) );
  AND U16709 ( .A(n12596), .B(n12597), .Z(n12595) );
  NAND U16710 ( .A(o[263]), .B(n11804), .Z(n12597) );
  NANDN U16711 ( .A(n11805), .B(creg[263]), .Z(n12596) );
  NAND U16712 ( .A(n12598), .B(n9385), .Z(n6921) );
  NANDN U16713 ( .A(init), .B(m[264]), .Z(n9385) );
  AND U16714 ( .A(n12599), .B(n12600), .Z(n12598) );
  NAND U16715 ( .A(o[264]), .B(n11804), .Z(n12600) );
  NANDN U16716 ( .A(n11805), .B(creg[264]), .Z(n12599) );
  NAND U16717 ( .A(n12601), .B(n9383), .Z(n6920) );
  NANDN U16718 ( .A(init), .B(m[265]), .Z(n9383) );
  AND U16719 ( .A(n12602), .B(n12603), .Z(n12601) );
  NAND U16720 ( .A(o[265]), .B(n11804), .Z(n12603) );
  NANDN U16721 ( .A(n11805), .B(creg[265]), .Z(n12602) );
  NAND U16722 ( .A(n12604), .B(n9381), .Z(n6919) );
  NANDN U16723 ( .A(init), .B(m[266]), .Z(n9381) );
  AND U16724 ( .A(n12605), .B(n12606), .Z(n12604) );
  NAND U16725 ( .A(o[266]), .B(n11804), .Z(n12606) );
  NANDN U16726 ( .A(n11805), .B(creg[266]), .Z(n12605) );
  NAND U16727 ( .A(n12607), .B(n9379), .Z(n6918) );
  NANDN U16728 ( .A(init), .B(m[267]), .Z(n9379) );
  AND U16729 ( .A(n12608), .B(n12609), .Z(n12607) );
  NAND U16730 ( .A(o[267]), .B(n11804), .Z(n12609) );
  NANDN U16731 ( .A(n11805), .B(creg[267]), .Z(n12608) );
  NAND U16732 ( .A(n12610), .B(n9377), .Z(n6917) );
  NANDN U16733 ( .A(init), .B(m[268]), .Z(n9377) );
  AND U16734 ( .A(n12611), .B(n12612), .Z(n12610) );
  NAND U16735 ( .A(o[268]), .B(n11804), .Z(n12612) );
  NANDN U16736 ( .A(n11805), .B(creg[268]), .Z(n12611) );
  NAND U16737 ( .A(n12613), .B(n9375), .Z(n6916) );
  NANDN U16738 ( .A(init), .B(m[269]), .Z(n9375) );
  AND U16739 ( .A(n12614), .B(n12615), .Z(n12613) );
  NAND U16740 ( .A(o[269]), .B(n11804), .Z(n12615) );
  NANDN U16741 ( .A(n11805), .B(creg[269]), .Z(n12614) );
  NAND U16742 ( .A(n12616), .B(n9371), .Z(n6915) );
  NANDN U16743 ( .A(init), .B(m[270]), .Z(n9371) );
  AND U16744 ( .A(n12617), .B(n12618), .Z(n12616) );
  NAND U16745 ( .A(o[270]), .B(n11804), .Z(n12618) );
  NANDN U16746 ( .A(n11805), .B(creg[270]), .Z(n12617) );
  NAND U16747 ( .A(n12619), .B(n9369), .Z(n6914) );
  NANDN U16748 ( .A(init), .B(m[271]), .Z(n9369) );
  AND U16749 ( .A(n12620), .B(n12621), .Z(n12619) );
  NAND U16750 ( .A(o[271]), .B(n11804), .Z(n12621) );
  NANDN U16751 ( .A(n11805), .B(creg[271]), .Z(n12620) );
  NAND U16752 ( .A(n12622), .B(n9367), .Z(n6913) );
  NANDN U16753 ( .A(init), .B(m[272]), .Z(n9367) );
  AND U16754 ( .A(n12623), .B(n12624), .Z(n12622) );
  NAND U16755 ( .A(o[272]), .B(n11804), .Z(n12624) );
  NANDN U16756 ( .A(n11805), .B(creg[272]), .Z(n12623) );
  NAND U16757 ( .A(n12625), .B(n9365), .Z(n6912) );
  NANDN U16758 ( .A(init), .B(m[273]), .Z(n9365) );
  AND U16759 ( .A(n12626), .B(n12627), .Z(n12625) );
  NAND U16760 ( .A(o[273]), .B(n11804), .Z(n12627) );
  NANDN U16761 ( .A(n11805), .B(creg[273]), .Z(n12626) );
  NAND U16762 ( .A(n12628), .B(n9363), .Z(n6911) );
  NANDN U16763 ( .A(init), .B(m[274]), .Z(n9363) );
  AND U16764 ( .A(n12629), .B(n12630), .Z(n12628) );
  NAND U16765 ( .A(o[274]), .B(n11804), .Z(n12630) );
  NANDN U16766 ( .A(n11805), .B(creg[274]), .Z(n12629) );
  NAND U16767 ( .A(n12631), .B(n9361), .Z(n6910) );
  NANDN U16768 ( .A(init), .B(m[275]), .Z(n9361) );
  AND U16769 ( .A(n12632), .B(n12633), .Z(n12631) );
  NAND U16770 ( .A(o[275]), .B(n11804), .Z(n12633) );
  NANDN U16771 ( .A(n11805), .B(creg[275]), .Z(n12632) );
  NAND U16772 ( .A(n12634), .B(n9359), .Z(n6909) );
  NANDN U16773 ( .A(init), .B(m[276]), .Z(n9359) );
  AND U16774 ( .A(n12635), .B(n12636), .Z(n12634) );
  NAND U16775 ( .A(o[276]), .B(n11804), .Z(n12636) );
  NANDN U16776 ( .A(n11805), .B(creg[276]), .Z(n12635) );
  NAND U16777 ( .A(n12637), .B(n9357), .Z(n6908) );
  NANDN U16778 ( .A(init), .B(m[277]), .Z(n9357) );
  AND U16779 ( .A(n12638), .B(n12639), .Z(n12637) );
  NAND U16780 ( .A(o[277]), .B(n11804), .Z(n12639) );
  NANDN U16781 ( .A(n11805), .B(creg[277]), .Z(n12638) );
  NAND U16782 ( .A(n12640), .B(n9355), .Z(n6907) );
  NANDN U16783 ( .A(init), .B(m[278]), .Z(n9355) );
  AND U16784 ( .A(n12641), .B(n12642), .Z(n12640) );
  NAND U16785 ( .A(o[278]), .B(n11804), .Z(n12642) );
  NANDN U16786 ( .A(n11805), .B(creg[278]), .Z(n12641) );
  NAND U16787 ( .A(n12643), .B(n9353), .Z(n6906) );
  NANDN U16788 ( .A(init), .B(m[279]), .Z(n9353) );
  AND U16789 ( .A(n12644), .B(n12645), .Z(n12643) );
  NAND U16790 ( .A(o[279]), .B(n11804), .Z(n12645) );
  NANDN U16791 ( .A(n11805), .B(creg[279]), .Z(n12644) );
  NAND U16792 ( .A(n12646), .B(n9349), .Z(n6905) );
  NANDN U16793 ( .A(init), .B(m[280]), .Z(n9349) );
  AND U16794 ( .A(n12647), .B(n12648), .Z(n12646) );
  NAND U16795 ( .A(o[280]), .B(n11804), .Z(n12648) );
  NANDN U16796 ( .A(n11805), .B(creg[280]), .Z(n12647) );
  NAND U16797 ( .A(n12649), .B(n9347), .Z(n6904) );
  NANDN U16798 ( .A(init), .B(m[281]), .Z(n9347) );
  AND U16799 ( .A(n12650), .B(n12651), .Z(n12649) );
  NAND U16800 ( .A(o[281]), .B(n11804), .Z(n12651) );
  NANDN U16801 ( .A(n11805), .B(creg[281]), .Z(n12650) );
  NAND U16802 ( .A(n12652), .B(n9345), .Z(n6903) );
  NANDN U16803 ( .A(init), .B(m[282]), .Z(n9345) );
  AND U16804 ( .A(n12653), .B(n12654), .Z(n12652) );
  NAND U16805 ( .A(o[282]), .B(n11804), .Z(n12654) );
  NANDN U16806 ( .A(n11805), .B(creg[282]), .Z(n12653) );
  NAND U16807 ( .A(n12655), .B(n9343), .Z(n6902) );
  NANDN U16808 ( .A(init), .B(m[283]), .Z(n9343) );
  AND U16809 ( .A(n12656), .B(n12657), .Z(n12655) );
  NAND U16810 ( .A(o[283]), .B(n11804), .Z(n12657) );
  NANDN U16811 ( .A(n11805), .B(creg[283]), .Z(n12656) );
  NAND U16812 ( .A(n12658), .B(n9341), .Z(n6901) );
  NANDN U16813 ( .A(init), .B(m[284]), .Z(n9341) );
  AND U16814 ( .A(n12659), .B(n12660), .Z(n12658) );
  NAND U16815 ( .A(o[284]), .B(n11804), .Z(n12660) );
  NANDN U16816 ( .A(n11805), .B(creg[284]), .Z(n12659) );
  NAND U16817 ( .A(n12661), .B(n9339), .Z(n6900) );
  NANDN U16818 ( .A(init), .B(m[285]), .Z(n9339) );
  AND U16819 ( .A(n12662), .B(n12663), .Z(n12661) );
  NAND U16820 ( .A(o[285]), .B(n11804), .Z(n12663) );
  NANDN U16821 ( .A(n11805), .B(creg[285]), .Z(n12662) );
  NAND U16822 ( .A(n12664), .B(n9337), .Z(n6899) );
  NANDN U16823 ( .A(init), .B(m[286]), .Z(n9337) );
  AND U16824 ( .A(n12665), .B(n12666), .Z(n12664) );
  NAND U16825 ( .A(o[286]), .B(n11804), .Z(n12666) );
  NANDN U16826 ( .A(n11805), .B(creg[286]), .Z(n12665) );
  NAND U16827 ( .A(n12667), .B(n9335), .Z(n6898) );
  NANDN U16828 ( .A(init), .B(m[287]), .Z(n9335) );
  AND U16829 ( .A(n12668), .B(n12669), .Z(n12667) );
  NAND U16830 ( .A(o[287]), .B(n11804), .Z(n12669) );
  NANDN U16831 ( .A(n11805), .B(creg[287]), .Z(n12668) );
  NAND U16832 ( .A(n12670), .B(n9333), .Z(n6897) );
  NANDN U16833 ( .A(init), .B(m[288]), .Z(n9333) );
  AND U16834 ( .A(n12671), .B(n12672), .Z(n12670) );
  NAND U16835 ( .A(o[288]), .B(n11804), .Z(n12672) );
  NANDN U16836 ( .A(n11805), .B(creg[288]), .Z(n12671) );
  NAND U16837 ( .A(n12673), .B(n9331), .Z(n6896) );
  NANDN U16838 ( .A(init), .B(m[289]), .Z(n9331) );
  AND U16839 ( .A(n12674), .B(n12675), .Z(n12673) );
  NAND U16840 ( .A(o[289]), .B(n11804), .Z(n12675) );
  NANDN U16841 ( .A(n11805), .B(creg[289]), .Z(n12674) );
  NAND U16842 ( .A(n12676), .B(n9327), .Z(n6895) );
  NANDN U16843 ( .A(init), .B(m[290]), .Z(n9327) );
  AND U16844 ( .A(n12677), .B(n12678), .Z(n12676) );
  NAND U16845 ( .A(o[290]), .B(n11804), .Z(n12678) );
  NANDN U16846 ( .A(n11805), .B(creg[290]), .Z(n12677) );
  NAND U16847 ( .A(n12679), .B(n9325), .Z(n6894) );
  NANDN U16848 ( .A(init), .B(m[291]), .Z(n9325) );
  AND U16849 ( .A(n12680), .B(n12681), .Z(n12679) );
  NAND U16850 ( .A(o[291]), .B(n11804), .Z(n12681) );
  NANDN U16851 ( .A(n11805), .B(creg[291]), .Z(n12680) );
  NAND U16852 ( .A(n12682), .B(n9323), .Z(n6893) );
  NANDN U16853 ( .A(init), .B(m[292]), .Z(n9323) );
  AND U16854 ( .A(n12683), .B(n12684), .Z(n12682) );
  NAND U16855 ( .A(o[292]), .B(n11804), .Z(n12684) );
  NANDN U16856 ( .A(n11805), .B(creg[292]), .Z(n12683) );
  NAND U16857 ( .A(n12685), .B(n9321), .Z(n6892) );
  NANDN U16858 ( .A(init), .B(m[293]), .Z(n9321) );
  AND U16859 ( .A(n12686), .B(n12687), .Z(n12685) );
  NAND U16860 ( .A(o[293]), .B(n11804), .Z(n12687) );
  NANDN U16861 ( .A(n11805), .B(creg[293]), .Z(n12686) );
  NAND U16862 ( .A(n12688), .B(n9319), .Z(n6891) );
  NANDN U16863 ( .A(init), .B(m[294]), .Z(n9319) );
  AND U16864 ( .A(n12689), .B(n12690), .Z(n12688) );
  NAND U16865 ( .A(o[294]), .B(n11804), .Z(n12690) );
  NANDN U16866 ( .A(n11805), .B(creg[294]), .Z(n12689) );
  NAND U16867 ( .A(n12691), .B(n9317), .Z(n6890) );
  NANDN U16868 ( .A(init), .B(m[295]), .Z(n9317) );
  AND U16869 ( .A(n12692), .B(n12693), .Z(n12691) );
  NAND U16870 ( .A(o[295]), .B(n11804), .Z(n12693) );
  NANDN U16871 ( .A(n11805), .B(creg[295]), .Z(n12692) );
  NAND U16872 ( .A(n12694), .B(n9315), .Z(n6889) );
  NANDN U16873 ( .A(init), .B(m[296]), .Z(n9315) );
  AND U16874 ( .A(n12695), .B(n12696), .Z(n12694) );
  NAND U16875 ( .A(o[296]), .B(n11804), .Z(n12696) );
  NANDN U16876 ( .A(n11805), .B(creg[296]), .Z(n12695) );
  NAND U16877 ( .A(n12697), .B(n9313), .Z(n6888) );
  NANDN U16878 ( .A(init), .B(m[297]), .Z(n9313) );
  AND U16879 ( .A(n12698), .B(n12699), .Z(n12697) );
  NAND U16880 ( .A(o[297]), .B(n11804), .Z(n12699) );
  NANDN U16881 ( .A(n11805), .B(creg[297]), .Z(n12698) );
  NAND U16882 ( .A(n12700), .B(n9311), .Z(n6887) );
  NANDN U16883 ( .A(init), .B(m[298]), .Z(n9311) );
  AND U16884 ( .A(n12701), .B(n12702), .Z(n12700) );
  NAND U16885 ( .A(o[298]), .B(n11804), .Z(n12702) );
  NANDN U16886 ( .A(n11805), .B(creg[298]), .Z(n12701) );
  NAND U16887 ( .A(n12703), .B(n9309), .Z(n6886) );
  NANDN U16888 ( .A(init), .B(m[299]), .Z(n9309) );
  AND U16889 ( .A(n12704), .B(n12705), .Z(n12703) );
  NAND U16890 ( .A(o[299]), .B(n11804), .Z(n12705) );
  NANDN U16891 ( .A(n11805), .B(creg[299]), .Z(n12704) );
  NAND U16892 ( .A(n12706), .B(n9303), .Z(n6885) );
  NANDN U16893 ( .A(init), .B(m[300]), .Z(n9303) );
  AND U16894 ( .A(n12707), .B(n12708), .Z(n12706) );
  NAND U16895 ( .A(o[300]), .B(n11804), .Z(n12708) );
  NANDN U16896 ( .A(n11805), .B(creg[300]), .Z(n12707) );
  NAND U16897 ( .A(n12709), .B(n9301), .Z(n6884) );
  NANDN U16898 ( .A(init), .B(m[301]), .Z(n9301) );
  AND U16899 ( .A(n12710), .B(n12711), .Z(n12709) );
  NAND U16900 ( .A(o[301]), .B(n11804), .Z(n12711) );
  NANDN U16901 ( .A(n11805), .B(creg[301]), .Z(n12710) );
  NAND U16902 ( .A(n12712), .B(n9299), .Z(n6883) );
  NANDN U16903 ( .A(init), .B(m[302]), .Z(n9299) );
  AND U16904 ( .A(n12713), .B(n12714), .Z(n12712) );
  NAND U16905 ( .A(o[302]), .B(n11804), .Z(n12714) );
  NANDN U16906 ( .A(n11805), .B(creg[302]), .Z(n12713) );
  NAND U16907 ( .A(n12715), .B(n9297), .Z(n6882) );
  NANDN U16908 ( .A(init), .B(m[303]), .Z(n9297) );
  AND U16909 ( .A(n12716), .B(n12717), .Z(n12715) );
  NAND U16910 ( .A(o[303]), .B(n11804), .Z(n12717) );
  NANDN U16911 ( .A(n11805), .B(creg[303]), .Z(n12716) );
  NAND U16912 ( .A(n12718), .B(n9295), .Z(n6881) );
  NANDN U16913 ( .A(init), .B(m[304]), .Z(n9295) );
  AND U16914 ( .A(n12719), .B(n12720), .Z(n12718) );
  NAND U16915 ( .A(o[304]), .B(n11804), .Z(n12720) );
  NANDN U16916 ( .A(n11805), .B(creg[304]), .Z(n12719) );
  NAND U16917 ( .A(n12721), .B(n9293), .Z(n6880) );
  NANDN U16918 ( .A(init), .B(m[305]), .Z(n9293) );
  AND U16919 ( .A(n12722), .B(n12723), .Z(n12721) );
  NAND U16920 ( .A(o[305]), .B(n11804), .Z(n12723) );
  NANDN U16921 ( .A(n11805), .B(creg[305]), .Z(n12722) );
  NAND U16922 ( .A(n12724), .B(n9291), .Z(n6879) );
  NANDN U16923 ( .A(init), .B(m[306]), .Z(n9291) );
  AND U16924 ( .A(n12725), .B(n12726), .Z(n12724) );
  NAND U16925 ( .A(o[306]), .B(n11804), .Z(n12726) );
  NANDN U16926 ( .A(n11805), .B(creg[306]), .Z(n12725) );
  NAND U16927 ( .A(n12727), .B(n9289), .Z(n6878) );
  NANDN U16928 ( .A(init), .B(m[307]), .Z(n9289) );
  AND U16929 ( .A(n12728), .B(n12729), .Z(n12727) );
  NAND U16930 ( .A(o[307]), .B(n11804), .Z(n12729) );
  NANDN U16931 ( .A(n11805), .B(creg[307]), .Z(n12728) );
  NAND U16932 ( .A(n12730), .B(n9287), .Z(n6877) );
  NANDN U16933 ( .A(init), .B(m[308]), .Z(n9287) );
  AND U16934 ( .A(n12731), .B(n12732), .Z(n12730) );
  NAND U16935 ( .A(o[308]), .B(n11804), .Z(n12732) );
  NANDN U16936 ( .A(n11805), .B(creg[308]), .Z(n12731) );
  NAND U16937 ( .A(n12733), .B(n9285), .Z(n6876) );
  NANDN U16938 ( .A(init), .B(m[309]), .Z(n9285) );
  AND U16939 ( .A(n12734), .B(n12735), .Z(n12733) );
  NAND U16940 ( .A(o[309]), .B(n11804), .Z(n12735) );
  NANDN U16941 ( .A(n11805), .B(creg[309]), .Z(n12734) );
  NAND U16942 ( .A(n12736), .B(n9281), .Z(n6875) );
  NANDN U16943 ( .A(init), .B(m[310]), .Z(n9281) );
  AND U16944 ( .A(n12737), .B(n12738), .Z(n12736) );
  NAND U16945 ( .A(o[310]), .B(n11804), .Z(n12738) );
  NANDN U16946 ( .A(n11805), .B(creg[310]), .Z(n12737) );
  NAND U16947 ( .A(n12739), .B(n9279), .Z(n6874) );
  NANDN U16948 ( .A(init), .B(m[311]), .Z(n9279) );
  AND U16949 ( .A(n12740), .B(n12741), .Z(n12739) );
  NAND U16950 ( .A(o[311]), .B(n11804), .Z(n12741) );
  NANDN U16951 ( .A(n11805), .B(creg[311]), .Z(n12740) );
  NAND U16952 ( .A(n12742), .B(n9277), .Z(n6873) );
  NANDN U16953 ( .A(init), .B(m[312]), .Z(n9277) );
  AND U16954 ( .A(n12743), .B(n12744), .Z(n12742) );
  NAND U16955 ( .A(o[312]), .B(n11804), .Z(n12744) );
  NANDN U16956 ( .A(n11805), .B(creg[312]), .Z(n12743) );
  NAND U16957 ( .A(n12745), .B(n9275), .Z(n6872) );
  NANDN U16958 ( .A(init), .B(m[313]), .Z(n9275) );
  AND U16959 ( .A(n12746), .B(n12747), .Z(n12745) );
  NAND U16960 ( .A(o[313]), .B(n11804), .Z(n12747) );
  NANDN U16961 ( .A(n11805), .B(creg[313]), .Z(n12746) );
  NAND U16962 ( .A(n12748), .B(n9273), .Z(n6871) );
  NANDN U16963 ( .A(init), .B(m[314]), .Z(n9273) );
  AND U16964 ( .A(n12749), .B(n12750), .Z(n12748) );
  NAND U16965 ( .A(o[314]), .B(n11804), .Z(n12750) );
  NANDN U16966 ( .A(n11805), .B(creg[314]), .Z(n12749) );
  NAND U16967 ( .A(n12751), .B(n9271), .Z(n6870) );
  NANDN U16968 ( .A(init), .B(m[315]), .Z(n9271) );
  AND U16969 ( .A(n12752), .B(n12753), .Z(n12751) );
  NAND U16970 ( .A(o[315]), .B(n11804), .Z(n12753) );
  NANDN U16971 ( .A(n11805), .B(creg[315]), .Z(n12752) );
  NAND U16972 ( .A(n12754), .B(n9269), .Z(n6869) );
  NANDN U16973 ( .A(init), .B(m[316]), .Z(n9269) );
  AND U16974 ( .A(n12755), .B(n12756), .Z(n12754) );
  NAND U16975 ( .A(o[316]), .B(n11804), .Z(n12756) );
  NANDN U16976 ( .A(n11805), .B(creg[316]), .Z(n12755) );
  NAND U16977 ( .A(n12757), .B(n9267), .Z(n6868) );
  NANDN U16978 ( .A(init), .B(m[317]), .Z(n9267) );
  AND U16979 ( .A(n12758), .B(n12759), .Z(n12757) );
  NAND U16980 ( .A(o[317]), .B(n11804), .Z(n12759) );
  NANDN U16981 ( .A(n11805), .B(creg[317]), .Z(n12758) );
  NAND U16982 ( .A(n12760), .B(n9265), .Z(n6867) );
  NANDN U16983 ( .A(init), .B(m[318]), .Z(n9265) );
  AND U16984 ( .A(n12761), .B(n12762), .Z(n12760) );
  NAND U16985 ( .A(o[318]), .B(n11804), .Z(n12762) );
  NANDN U16986 ( .A(n11805), .B(creg[318]), .Z(n12761) );
  NAND U16987 ( .A(n12763), .B(n9263), .Z(n6866) );
  NANDN U16988 ( .A(init), .B(m[319]), .Z(n9263) );
  AND U16989 ( .A(n12764), .B(n12765), .Z(n12763) );
  NAND U16990 ( .A(o[319]), .B(n11804), .Z(n12765) );
  NANDN U16991 ( .A(n11805), .B(creg[319]), .Z(n12764) );
  NAND U16992 ( .A(n12766), .B(n9259), .Z(n6865) );
  NANDN U16993 ( .A(init), .B(m[320]), .Z(n9259) );
  AND U16994 ( .A(n12767), .B(n12768), .Z(n12766) );
  NAND U16995 ( .A(o[320]), .B(n11804), .Z(n12768) );
  NANDN U16996 ( .A(n11805), .B(creg[320]), .Z(n12767) );
  NAND U16997 ( .A(n12769), .B(n9257), .Z(n6864) );
  NANDN U16998 ( .A(init), .B(m[321]), .Z(n9257) );
  AND U16999 ( .A(n12770), .B(n12771), .Z(n12769) );
  NAND U17000 ( .A(o[321]), .B(n11804), .Z(n12771) );
  NANDN U17001 ( .A(n11805), .B(creg[321]), .Z(n12770) );
  NAND U17002 ( .A(n12772), .B(n9255), .Z(n6863) );
  NANDN U17003 ( .A(init), .B(m[322]), .Z(n9255) );
  AND U17004 ( .A(n12773), .B(n12774), .Z(n12772) );
  NAND U17005 ( .A(o[322]), .B(n11804), .Z(n12774) );
  NANDN U17006 ( .A(n11805), .B(creg[322]), .Z(n12773) );
  NAND U17007 ( .A(n12775), .B(n9253), .Z(n6862) );
  NANDN U17008 ( .A(init), .B(m[323]), .Z(n9253) );
  AND U17009 ( .A(n12776), .B(n12777), .Z(n12775) );
  NAND U17010 ( .A(o[323]), .B(n11804), .Z(n12777) );
  NANDN U17011 ( .A(n11805), .B(creg[323]), .Z(n12776) );
  NAND U17012 ( .A(n12778), .B(n9251), .Z(n6861) );
  NANDN U17013 ( .A(init), .B(m[324]), .Z(n9251) );
  AND U17014 ( .A(n12779), .B(n12780), .Z(n12778) );
  NAND U17015 ( .A(o[324]), .B(n11804), .Z(n12780) );
  NANDN U17016 ( .A(n11805), .B(creg[324]), .Z(n12779) );
  NAND U17017 ( .A(n12781), .B(n9249), .Z(n6860) );
  NANDN U17018 ( .A(init), .B(m[325]), .Z(n9249) );
  AND U17019 ( .A(n12782), .B(n12783), .Z(n12781) );
  NAND U17020 ( .A(o[325]), .B(n11804), .Z(n12783) );
  NANDN U17021 ( .A(n11805), .B(creg[325]), .Z(n12782) );
  NAND U17022 ( .A(n12784), .B(n9247), .Z(n6859) );
  NANDN U17023 ( .A(init), .B(m[326]), .Z(n9247) );
  AND U17024 ( .A(n12785), .B(n12786), .Z(n12784) );
  NAND U17025 ( .A(o[326]), .B(n11804), .Z(n12786) );
  NANDN U17026 ( .A(n11805), .B(creg[326]), .Z(n12785) );
  NAND U17027 ( .A(n12787), .B(n9245), .Z(n6858) );
  NANDN U17028 ( .A(init), .B(m[327]), .Z(n9245) );
  AND U17029 ( .A(n12788), .B(n12789), .Z(n12787) );
  NAND U17030 ( .A(o[327]), .B(n11804), .Z(n12789) );
  NANDN U17031 ( .A(n11805), .B(creg[327]), .Z(n12788) );
  NAND U17032 ( .A(n12790), .B(n9243), .Z(n6857) );
  NANDN U17033 ( .A(init), .B(m[328]), .Z(n9243) );
  AND U17034 ( .A(n12791), .B(n12792), .Z(n12790) );
  NAND U17035 ( .A(o[328]), .B(n11804), .Z(n12792) );
  NANDN U17036 ( .A(n11805), .B(creg[328]), .Z(n12791) );
  NAND U17037 ( .A(n12793), .B(n9241), .Z(n6856) );
  NANDN U17038 ( .A(init), .B(m[329]), .Z(n9241) );
  AND U17039 ( .A(n12794), .B(n12795), .Z(n12793) );
  NAND U17040 ( .A(o[329]), .B(n11804), .Z(n12795) );
  NANDN U17041 ( .A(n11805), .B(creg[329]), .Z(n12794) );
  NAND U17042 ( .A(n12796), .B(n9237), .Z(n6855) );
  NANDN U17043 ( .A(init), .B(m[330]), .Z(n9237) );
  AND U17044 ( .A(n12797), .B(n12798), .Z(n12796) );
  NAND U17045 ( .A(o[330]), .B(n11804), .Z(n12798) );
  NANDN U17046 ( .A(n11805), .B(creg[330]), .Z(n12797) );
  NAND U17047 ( .A(n12799), .B(n9235), .Z(n6854) );
  NANDN U17048 ( .A(init), .B(m[331]), .Z(n9235) );
  AND U17049 ( .A(n12800), .B(n12801), .Z(n12799) );
  NAND U17050 ( .A(o[331]), .B(n11804), .Z(n12801) );
  NANDN U17051 ( .A(n11805), .B(creg[331]), .Z(n12800) );
  NAND U17052 ( .A(n12802), .B(n9233), .Z(n6853) );
  NANDN U17053 ( .A(init), .B(m[332]), .Z(n9233) );
  AND U17054 ( .A(n12803), .B(n12804), .Z(n12802) );
  NAND U17055 ( .A(o[332]), .B(n11804), .Z(n12804) );
  NANDN U17056 ( .A(n11805), .B(creg[332]), .Z(n12803) );
  NAND U17057 ( .A(n12805), .B(n9231), .Z(n6852) );
  NANDN U17058 ( .A(init), .B(m[333]), .Z(n9231) );
  AND U17059 ( .A(n12806), .B(n12807), .Z(n12805) );
  NAND U17060 ( .A(o[333]), .B(n11804), .Z(n12807) );
  NANDN U17061 ( .A(n11805), .B(creg[333]), .Z(n12806) );
  NAND U17062 ( .A(n12808), .B(n9229), .Z(n6851) );
  NANDN U17063 ( .A(init), .B(m[334]), .Z(n9229) );
  AND U17064 ( .A(n12809), .B(n12810), .Z(n12808) );
  NAND U17065 ( .A(o[334]), .B(n11804), .Z(n12810) );
  NANDN U17066 ( .A(n11805), .B(creg[334]), .Z(n12809) );
  NAND U17067 ( .A(n12811), .B(n9227), .Z(n6850) );
  NANDN U17068 ( .A(init), .B(m[335]), .Z(n9227) );
  AND U17069 ( .A(n12812), .B(n12813), .Z(n12811) );
  NAND U17070 ( .A(o[335]), .B(n11804), .Z(n12813) );
  NANDN U17071 ( .A(n11805), .B(creg[335]), .Z(n12812) );
  NAND U17072 ( .A(n12814), .B(n9225), .Z(n6849) );
  NANDN U17073 ( .A(init), .B(m[336]), .Z(n9225) );
  AND U17074 ( .A(n12815), .B(n12816), .Z(n12814) );
  NAND U17075 ( .A(o[336]), .B(n11804), .Z(n12816) );
  NANDN U17076 ( .A(n11805), .B(creg[336]), .Z(n12815) );
  NAND U17077 ( .A(n12817), .B(n9223), .Z(n6848) );
  NANDN U17078 ( .A(init), .B(m[337]), .Z(n9223) );
  AND U17079 ( .A(n12818), .B(n12819), .Z(n12817) );
  NAND U17080 ( .A(o[337]), .B(n11804), .Z(n12819) );
  NANDN U17081 ( .A(n11805), .B(creg[337]), .Z(n12818) );
  NAND U17082 ( .A(n12820), .B(n9221), .Z(n6847) );
  NANDN U17083 ( .A(init), .B(m[338]), .Z(n9221) );
  AND U17084 ( .A(n12821), .B(n12822), .Z(n12820) );
  NAND U17085 ( .A(o[338]), .B(n11804), .Z(n12822) );
  NANDN U17086 ( .A(n11805), .B(creg[338]), .Z(n12821) );
  NAND U17087 ( .A(n12823), .B(n9219), .Z(n6846) );
  NANDN U17088 ( .A(init), .B(m[339]), .Z(n9219) );
  AND U17089 ( .A(n12824), .B(n12825), .Z(n12823) );
  NAND U17090 ( .A(o[339]), .B(n11804), .Z(n12825) );
  NANDN U17091 ( .A(n11805), .B(creg[339]), .Z(n12824) );
  NAND U17092 ( .A(n12826), .B(n9215), .Z(n6845) );
  NANDN U17093 ( .A(init), .B(m[340]), .Z(n9215) );
  AND U17094 ( .A(n12827), .B(n12828), .Z(n12826) );
  NAND U17095 ( .A(o[340]), .B(n11804), .Z(n12828) );
  NANDN U17096 ( .A(n11805), .B(creg[340]), .Z(n12827) );
  NAND U17097 ( .A(n12829), .B(n9213), .Z(n6844) );
  NANDN U17098 ( .A(init), .B(m[341]), .Z(n9213) );
  AND U17099 ( .A(n12830), .B(n12831), .Z(n12829) );
  NAND U17100 ( .A(o[341]), .B(n11804), .Z(n12831) );
  NANDN U17101 ( .A(n11805), .B(creg[341]), .Z(n12830) );
  NAND U17102 ( .A(n12832), .B(n9211), .Z(n6843) );
  NANDN U17103 ( .A(init), .B(m[342]), .Z(n9211) );
  AND U17104 ( .A(n12833), .B(n12834), .Z(n12832) );
  NAND U17105 ( .A(o[342]), .B(n11804), .Z(n12834) );
  NANDN U17106 ( .A(n11805), .B(creg[342]), .Z(n12833) );
  NAND U17107 ( .A(n12835), .B(n9209), .Z(n6842) );
  NANDN U17108 ( .A(init), .B(m[343]), .Z(n9209) );
  AND U17109 ( .A(n12836), .B(n12837), .Z(n12835) );
  NAND U17110 ( .A(o[343]), .B(n11804), .Z(n12837) );
  NANDN U17111 ( .A(n11805), .B(creg[343]), .Z(n12836) );
  NAND U17112 ( .A(n12838), .B(n9207), .Z(n6841) );
  NANDN U17113 ( .A(init), .B(m[344]), .Z(n9207) );
  AND U17114 ( .A(n12839), .B(n12840), .Z(n12838) );
  NAND U17115 ( .A(o[344]), .B(n11804), .Z(n12840) );
  NANDN U17116 ( .A(n11805), .B(creg[344]), .Z(n12839) );
  NAND U17117 ( .A(n12841), .B(n9205), .Z(n6840) );
  NANDN U17118 ( .A(init), .B(m[345]), .Z(n9205) );
  AND U17119 ( .A(n12842), .B(n12843), .Z(n12841) );
  NAND U17120 ( .A(o[345]), .B(n11804), .Z(n12843) );
  NANDN U17121 ( .A(n11805), .B(creg[345]), .Z(n12842) );
  NAND U17122 ( .A(n12844), .B(n9203), .Z(n6839) );
  NANDN U17123 ( .A(init), .B(m[346]), .Z(n9203) );
  AND U17124 ( .A(n12845), .B(n12846), .Z(n12844) );
  NAND U17125 ( .A(o[346]), .B(n11804), .Z(n12846) );
  NANDN U17126 ( .A(n11805), .B(creg[346]), .Z(n12845) );
  NAND U17127 ( .A(n12847), .B(n9201), .Z(n6838) );
  NANDN U17128 ( .A(init), .B(m[347]), .Z(n9201) );
  AND U17129 ( .A(n12848), .B(n12849), .Z(n12847) );
  NAND U17130 ( .A(o[347]), .B(n11804), .Z(n12849) );
  NANDN U17131 ( .A(n11805), .B(creg[347]), .Z(n12848) );
  NAND U17132 ( .A(n12850), .B(n9199), .Z(n6837) );
  NANDN U17133 ( .A(init), .B(m[348]), .Z(n9199) );
  AND U17134 ( .A(n12851), .B(n12852), .Z(n12850) );
  NAND U17135 ( .A(o[348]), .B(n11804), .Z(n12852) );
  NANDN U17136 ( .A(n11805), .B(creg[348]), .Z(n12851) );
  NAND U17137 ( .A(n12853), .B(n9197), .Z(n6836) );
  NANDN U17138 ( .A(init), .B(m[349]), .Z(n9197) );
  AND U17139 ( .A(n12854), .B(n12855), .Z(n12853) );
  NAND U17140 ( .A(o[349]), .B(n11804), .Z(n12855) );
  NANDN U17141 ( .A(n11805), .B(creg[349]), .Z(n12854) );
  NAND U17142 ( .A(n12856), .B(n9193), .Z(n6835) );
  NANDN U17143 ( .A(init), .B(m[350]), .Z(n9193) );
  AND U17144 ( .A(n12857), .B(n12858), .Z(n12856) );
  NAND U17145 ( .A(o[350]), .B(n11804), .Z(n12858) );
  NANDN U17146 ( .A(n11805), .B(creg[350]), .Z(n12857) );
  NAND U17147 ( .A(n12859), .B(n9191), .Z(n6834) );
  NANDN U17148 ( .A(init), .B(m[351]), .Z(n9191) );
  AND U17149 ( .A(n12860), .B(n12861), .Z(n12859) );
  NAND U17150 ( .A(o[351]), .B(n11804), .Z(n12861) );
  NANDN U17151 ( .A(n11805), .B(creg[351]), .Z(n12860) );
  NAND U17152 ( .A(n12862), .B(n9189), .Z(n6833) );
  NANDN U17153 ( .A(init), .B(m[352]), .Z(n9189) );
  AND U17154 ( .A(n12863), .B(n12864), .Z(n12862) );
  NAND U17155 ( .A(o[352]), .B(n11804), .Z(n12864) );
  NANDN U17156 ( .A(n11805), .B(creg[352]), .Z(n12863) );
  NAND U17157 ( .A(n12865), .B(n9187), .Z(n6832) );
  NANDN U17158 ( .A(init), .B(m[353]), .Z(n9187) );
  AND U17159 ( .A(n12866), .B(n12867), .Z(n12865) );
  NAND U17160 ( .A(o[353]), .B(n11804), .Z(n12867) );
  NANDN U17161 ( .A(n11805), .B(creg[353]), .Z(n12866) );
  NAND U17162 ( .A(n12868), .B(n9185), .Z(n6831) );
  NANDN U17163 ( .A(init), .B(m[354]), .Z(n9185) );
  AND U17164 ( .A(n12869), .B(n12870), .Z(n12868) );
  NAND U17165 ( .A(o[354]), .B(n11804), .Z(n12870) );
  NANDN U17166 ( .A(n11805), .B(creg[354]), .Z(n12869) );
  NAND U17167 ( .A(n12871), .B(n9183), .Z(n6830) );
  NANDN U17168 ( .A(init), .B(m[355]), .Z(n9183) );
  AND U17169 ( .A(n12872), .B(n12873), .Z(n12871) );
  NAND U17170 ( .A(o[355]), .B(n11804), .Z(n12873) );
  NANDN U17171 ( .A(n11805), .B(creg[355]), .Z(n12872) );
  NAND U17172 ( .A(n12874), .B(n9181), .Z(n6829) );
  NANDN U17173 ( .A(init), .B(m[356]), .Z(n9181) );
  AND U17174 ( .A(n12875), .B(n12876), .Z(n12874) );
  NAND U17175 ( .A(o[356]), .B(n11804), .Z(n12876) );
  NANDN U17176 ( .A(n11805), .B(creg[356]), .Z(n12875) );
  NAND U17177 ( .A(n12877), .B(n9179), .Z(n6828) );
  NANDN U17178 ( .A(init), .B(m[357]), .Z(n9179) );
  AND U17179 ( .A(n12878), .B(n12879), .Z(n12877) );
  NAND U17180 ( .A(o[357]), .B(n11804), .Z(n12879) );
  NANDN U17181 ( .A(n11805), .B(creg[357]), .Z(n12878) );
  NAND U17182 ( .A(n12880), .B(n9177), .Z(n6827) );
  NANDN U17183 ( .A(init), .B(m[358]), .Z(n9177) );
  AND U17184 ( .A(n12881), .B(n12882), .Z(n12880) );
  NAND U17185 ( .A(o[358]), .B(n11804), .Z(n12882) );
  NANDN U17186 ( .A(n11805), .B(creg[358]), .Z(n12881) );
  NAND U17187 ( .A(n12883), .B(n9175), .Z(n6826) );
  NANDN U17188 ( .A(init), .B(m[359]), .Z(n9175) );
  AND U17189 ( .A(n12884), .B(n12885), .Z(n12883) );
  NAND U17190 ( .A(o[359]), .B(n11804), .Z(n12885) );
  NANDN U17191 ( .A(n11805), .B(creg[359]), .Z(n12884) );
  NAND U17192 ( .A(n12886), .B(n9171), .Z(n6825) );
  NANDN U17193 ( .A(init), .B(m[360]), .Z(n9171) );
  AND U17194 ( .A(n12887), .B(n12888), .Z(n12886) );
  NAND U17195 ( .A(o[360]), .B(n11804), .Z(n12888) );
  NANDN U17196 ( .A(n11805), .B(creg[360]), .Z(n12887) );
  NAND U17197 ( .A(n12889), .B(n9169), .Z(n6824) );
  NANDN U17198 ( .A(init), .B(m[361]), .Z(n9169) );
  AND U17199 ( .A(n12890), .B(n12891), .Z(n12889) );
  NAND U17200 ( .A(o[361]), .B(n11804), .Z(n12891) );
  NANDN U17201 ( .A(n11805), .B(creg[361]), .Z(n12890) );
  NAND U17202 ( .A(n12892), .B(n9167), .Z(n6823) );
  NANDN U17203 ( .A(init), .B(m[362]), .Z(n9167) );
  AND U17204 ( .A(n12893), .B(n12894), .Z(n12892) );
  NAND U17205 ( .A(o[362]), .B(n11804), .Z(n12894) );
  NANDN U17206 ( .A(n11805), .B(creg[362]), .Z(n12893) );
  NAND U17207 ( .A(n12895), .B(n9165), .Z(n6822) );
  NANDN U17208 ( .A(init), .B(m[363]), .Z(n9165) );
  AND U17209 ( .A(n12896), .B(n12897), .Z(n12895) );
  NAND U17210 ( .A(o[363]), .B(n11804), .Z(n12897) );
  NANDN U17211 ( .A(n11805), .B(creg[363]), .Z(n12896) );
  NAND U17212 ( .A(n12898), .B(n9163), .Z(n6821) );
  NANDN U17213 ( .A(init), .B(m[364]), .Z(n9163) );
  AND U17214 ( .A(n12899), .B(n12900), .Z(n12898) );
  NAND U17215 ( .A(o[364]), .B(n11804), .Z(n12900) );
  NANDN U17216 ( .A(n11805), .B(creg[364]), .Z(n12899) );
  NAND U17217 ( .A(n12901), .B(n9161), .Z(n6820) );
  NANDN U17218 ( .A(init), .B(m[365]), .Z(n9161) );
  AND U17219 ( .A(n12902), .B(n12903), .Z(n12901) );
  NAND U17220 ( .A(o[365]), .B(n11804), .Z(n12903) );
  NANDN U17221 ( .A(n11805), .B(creg[365]), .Z(n12902) );
  NAND U17222 ( .A(n12904), .B(n9159), .Z(n6819) );
  NANDN U17223 ( .A(init), .B(m[366]), .Z(n9159) );
  AND U17224 ( .A(n12905), .B(n12906), .Z(n12904) );
  NAND U17225 ( .A(o[366]), .B(n11804), .Z(n12906) );
  NANDN U17226 ( .A(n11805), .B(creg[366]), .Z(n12905) );
  NAND U17227 ( .A(n12907), .B(n9157), .Z(n6818) );
  NANDN U17228 ( .A(init), .B(m[367]), .Z(n9157) );
  AND U17229 ( .A(n12908), .B(n12909), .Z(n12907) );
  NAND U17230 ( .A(o[367]), .B(n11804), .Z(n12909) );
  NANDN U17231 ( .A(n11805), .B(creg[367]), .Z(n12908) );
  NAND U17232 ( .A(n12910), .B(n9155), .Z(n6817) );
  NANDN U17233 ( .A(init), .B(m[368]), .Z(n9155) );
  AND U17234 ( .A(n12911), .B(n12912), .Z(n12910) );
  NAND U17235 ( .A(o[368]), .B(n11804), .Z(n12912) );
  NANDN U17236 ( .A(n11805), .B(creg[368]), .Z(n12911) );
  NAND U17237 ( .A(n12913), .B(n9153), .Z(n6816) );
  NANDN U17238 ( .A(init), .B(m[369]), .Z(n9153) );
  AND U17239 ( .A(n12914), .B(n12915), .Z(n12913) );
  NAND U17240 ( .A(o[369]), .B(n11804), .Z(n12915) );
  NANDN U17241 ( .A(n11805), .B(creg[369]), .Z(n12914) );
  NAND U17242 ( .A(n12916), .B(n9149), .Z(n6815) );
  NANDN U17243 ( .A(init), .B(m[370]), .Z(n9149) );
  AND U17244 ( .A(n12917), .B(n12918), .Z(n12916) );
  NAND U17245 ( .A(o[370]), .B(n11804), .Z(n12918) );
  NANDN U17246 ( .A(n11805), .B(creg[370]), .Z(n12917) );
  NAND U17247 ( .A(n12919), .B(n9147), .Z(n6814) );
  NANDN U17248 ( .A(init), .B(m[371]), .Z(n9147) );
  AND U17249 ( .A(n12920), .B(n12921), .Z(n12919) );
  NAND U17250 ( .A(o[371]), .B(n11804), .Z(n12921) );
  NANDN U17251 ( .A(n11805), .B(creg[371]), .Z(n12920) );
  NAND U17252 ( .A(n12922), .B(n9145), .Z(n6813) );
  NANDN U17253 ( .A(init), .B(m[372]), .Z(n9145) );
  AND U17254 ( .A(n12923), .B(n12924), .Z(n12922) );
  NAND U17255 ( .A(o[372]), .B(n11804), .Z(n12924) );
  NANDN U17256 ( .A(n11805), .B(creg[372]), .Z(n12923) );
  NAND U17257 ( .A(n12925), .B(n9143), .Z(n6812) );
  NANDN U17258 ( .A(init), .B(m[373]), .Z(n9143) );
  AND U17259 ( .A(n12926), .B(n12927), .Z(n12925) );
  NAND U17260 ( .A(o[373]), .B(n11804), .Z(n12927) );
  NANDN U17261 ( .A(n11805), .B(creg[373]), .Z(n12926) );
  NAND U17262 ( .A(n12928), .B(n9141), .Z(n6811) );
  NANDN U17263 ( .A(init), .B(m[374]), .Z(n9141) );
  AND U17264 ( .A(n12929), .B(n12930), .Z(n12928) );
  NAND U17265 ( .A(o[374]), .B(n11804), .Z(n12930) );
  NANDN U17266 ( .A(n11805), .B(creg[374]), .Z(n12929) );
  NAND U17267 ( .A(n12931), .B(n9139), .Z(n6810) );
  NANDN U17268 ( .A(init), .B(m[375]), .Z(n9139) );
  AND U17269 ( .A(n12932), .B(n12933), .Z(n12931) );
  NAND U17270 ( .A(o[375]), .B(n11804), .Z(n12933) );
  NANDN U17271 ( .A(n11805), .B(creg[375]), .Z(n12932) );
  NAND U17272 ( .A(n12934), .B(n9137), .Z(n6809) );
  NANDN U17273 ( .A(init), .B(m[376]), .Z(n9137) );
  AND U17274 ( .A(n12935), .B(n12936), .Z(n12934) );
  NAND U17275 ( .A(o[376]), .B(n11804), .Z(n12936) );
  NANDN U17276 ( .A(n11805), .B(creg[376]), .Z(n12935) );
  NAND U17277 ( .A(n12937), .B(n9135), .Z(n6808) );
  NANDN U17278 ( .A(init), .B(m[377]), .Z(n9135) );
  AND U17279 ( .A(n12938), .B(n12939), .Z(n12937) );
  NAND U17280 ( .A(o[377]), .B(n11804), .Z(n12939) );
  NANDN U17281 ( .A(n11805), .B(creg[377]), .Z(n12938) );
  NAND U17282 ( .A(n12940), .B(n9133), .Z(n6807) );
  NANDN U17283 ( .A(init), .B(m[378]), .Z(n9133) );
  AND U17284 ( .A(n12941), .B(n12942), .Z(n12940) );
  NAND U17285 ( .A(o[378]), .B(n11804), .Z(n12942) );
  NANDN U17286 ( .A(n11805), .B(creg[378]), .Z(n12941) );
  NAND U17287 ( .A(n12943), .B(n9131), .Z(n6806) );
  NANDN U17288 ( .A(init), .B(m[379]), .Z(n9131) );
  AND U17289 ( .A(n12944), .B(n12945), .Z(n12943) );
  NAND U17290 ( .A(o[379]), .B(n11804), .Z(n12945) );
  NANDN U17291 ( .A(n11805), .B(creg[379]), .Z(n12944) );
  NAND U17292 ( .A(n12946), .B(n9127), .Z(n6805) );
  NANDN U17293 ( .A(init), .B(m[380]), .Z(n9127) );
  AND U17294 ( .A(n12947), .B(n12948), .Z(n12946) );
  NAND U17295 ( .A(o[380]), .B(n11804), .Z(n12948) );
  NANDN U17296 ( .A(n11805), .B(creg[380]), .Z(n12947) );
  NAND U17297 ( .A(n12949), .B(n9125), .Z(n6804) );
  NANDN U17298 ( .A(init), .B(m[381]), .Z(n9125) );
  AND U17299 ( .A(n12950), .B(n12951), .Z(n12949) );
  NAND U17300 ( .A(o[381]), .B(n11804), .Z(n12951) );
  NANDN U17301 ( .A(n11805), .B(creg[381]), .Z(n12950) );
  NAND U17302 ( .A(n12952), .B(n9123), .Z(n6803) );
  NANDN U17303 ( .A(init), .B(m[382]), .Z(n9123) );
  AND U17304 ( .A(n12953), .B(n12954), .Z(n12952) );
  NAND U17305 ( .A(o[382]), .B(n11804), .Z(n12954) );
  NANDN U17306 ( .A(n11805), .B(creg[382]), .Z(n12953) );
  NAND U17307 ( .A(n12955), .B(n9121), .Z(n6802) );
  NANDN U17308 ( .A(init), .B(m[383]), .Z(n9121) );
  AND U17309 ( .A(n12956), .B(n12957), .Z(n12955) );
  NAND U17310 ( .A(o[383]), .B(n11804), .Z(n12957) );
  NANDN U17311 ( .A(n11805), .B(creg[383]), .Z(n12956) );
  NAND U17312 ( .A(n12958), .B(n9119), .Z(n6801) );
  NANDN U17313 ( .A(init), .B(m[384]), .Z(n9119) );
  AND U17314 ( .A(n12959), .B(n12960), .Z(n12958) );
  NAND U17315 ( .A(o[384]), .B(n11804), .Z(n12960) );
  NANDN U17316 ( .A(n11805), .B(creg[384]), .Z(n12959) );
  NAND U17317 ( .A(n12961), .B(n9117), .Z(n6800) );
  NANDN U17318 ( .A(init), .B(m[385]), .Z(n9117) );
  AND U17319 ( .A(n12962), .B(n12963), .Z(n12961) );
  NAND U17320 ( .A(o[385]), .B(n11804), .Z(n12963) );
  NANDN U17321 ( .A(n11805), .B(creg[385]), .Z(n12962) );
  NAND U17322 ( .A(n12964), .B(n9115), .Z(n6799) );
  NANDN U17323 ( .A(init), .B(m[386]), .Z(n9115) );
  AND U17324 ( .A(n12965), .B(n12966), .Z(n12964) );
  NAND U17325 ( .A(o[386]), .B(n11804), .Z(n12966) );
  NANDN U17326 ( .A(n11805), .B(creg[386]), .Z(n12965) );
  NAND U17327 ( .A(n12967), .B(n9113), .Z(n6798) );
  NANDN U17328 ( .A(init), .B(m[387]), .Z(n9113) );
  AND U17329 ( .A(n12968), .B(n12969), .Z(n12967) );
  NAND U17330 ( .A(o[387]), .B(n11804), .Z(n12969) );
  NANDN U17331 ( .A(n11805), .B(creg[387]), .Z(n12968) );
  NAND U17332 ( .A(n12970), .B(n9111), .Z(n6797) );
  NANDN U17333 ( .A(init), .B(m[388]), .Z(n9111) );
  AND U17334 ( .A(n12971), .B(n12972), .Z(n12970) );
  NAND U17335 ( .A(o[388]), .B(n11804), .Z(n12972) );
  NANDN U17336 ( .A(n11805), .B(creg[388]), .Z(n12971) );
  NAND U17337 ( .A(n12973), .B(n9109), .Z(n6796) );
  NANDN U17338 ( .A(init), .B(m[389]), .Z(n9109) );
  AND U17339 ( .A(n12974), .B(n12975), .Z(n12973) );
  NAND U17340 ( .A(o[389]), .B(n11804), .Z(n12975) );
  NANDN U17341 ( .A(n11805), .B(creg[389]), .Z(n12974) );
  NAND U17342 ( .A(n12976), .B(n9105), .Z(n6795) );
  NANDN U17343 ( .A(init), .B(m[390]), .Z(n9105) );
  AND U17344 ( .A(n12977), .B(n12978), .Z(n12976) );
  NAND U17345 ( .A(o[390]), .B(n11804), .Z(n12978) );
  NANDN U17346 ( .A(n11805), .B(creg[390]), .Z(n12977) );
  NAND U17347 ( .A(n12979), .B(n9103), .Z(n6794) );
  NANDN U17348 ( .A(init), .B(m[391]), .Z(n9103) );
  AND U17349 ( .A(n12980), .B(n12981), .Z(n12979) );
  NAND U17350 ( .A(o[391]), .B(n11804), .Z(n12981) );
  NANDN U17351 ( .A(n11805), .B(creg[391]), .Z(n12980) );
  NAND U17352 ( .A(n12982), .B(n9101), .Z(n6793) );
  NANDN U17353 ( .A(init), .B(m[392]), .Z(n9101) );
  AND U17354 ( .A(n12983), .B(n12984), .Z(n12982) );
  NAND U17355 ( .A(o[392]), .B(n11804), .Z(n12984) );
  NANDN U17356 ( .A(n11805), .B(creg[392]), .Z(n12983) );
  NAND U17357 ( .A(n12985), .B(n9099), .Z(n6792) );
  NANDN U17358 ( .A(init), .B(m[393]), .Z(n9099) );
  AND U17359 ( .A(n12986), .B(n12987), .Z(n12985) );
  NAND U17360 ( .A(o[393]), .B(n11804), .Z(n12987) );
  NANDN U17361 ( .A(n11805), .B(creg[393]), .Z(n12986) );
  NAND U17362 ( .A(n12988), .B(n9097), .Z(n6791) );
  NANDN U17363 ( .A(init), .B(m[394]), .Z(n9097) );
  AND U17364 ( .A(n12989), .B(n12990), .Z(n12988) );
  NAND U17365 ( .A(o[394]), .B(n11804), .Z(n12990) );
  NANDN U17366 ( .A(n11805), .B(creg[394]), .Z(n12989) );
  NAND U17367 ( .A(n12991), .B(n9095), .Z(n6790) );
  NANDN U17368 ( .A(init), .B(m[395]), .Z(n9095) );
  AND U17369 ( .A(n12992), .B(n12993), .Z(n12991) );
  NAND U17370 ( .A(o[395]), .B(n11804), .Z(n12993) );
  NANDN U17371 ( .A(n11805), .B(creg[395]), .Z(n12992) );
  NAND U17372 ( .A(n12994), .B(n9093), .Z(n6789) );
  NANDN U17373 ( .A(init), .B(m[396]), .Z(n9093) );
  AND U17374 ( .A(n12995), .B(n12996), .Z(n12994) );
  NAND U17375 ( .A(o[396]), .B(n11804), .Z(n12996) );
  NANDN U17376 ( .A(n11805), .B(creg[396]), .Z(n12995) );
  NAND U17377 ( .A(n12997), .B(n9091), .Z(n6788) );
  NANDN U17378 ( .A(init), .B(m[397]), .Z(n9091) );
  AND U17379 ( .A(n12998), .B(n12999), .Z(n12997) );
  NAND U17380 ( .A(o[397]), .B(n11804), .Z(n12999) );
  NANDN U17381 ( .A(n11805), .B(creg[397]), .Z(n12998) );
  NAND U17382 ( .A(n13000), .B(n9089), .Z(n6787) );
  NANDN U17383 ( .A(init), .B(m[398]), .Z(n9089) );
  AND U17384 ( .A(n13001), .B(n13002), .Z(n13000) );
  NAND U17385 ( .A(o[398]), .B(n11804), .Z(n13002) );
  NANDN U17386 ( .A(n11805), .B(creg[398]), .Z(n13001) );
  NAND U17387 ( .A(n13003), .B(n9087), .Z(n6786) );
  NANDN U17388 ( .A(init), .B(m[399]), .Z(n9087) );
  AND U17389 ( .A(n13004), .B(n13005), .Z(n13003) );
  NAND U17390 ( .A(o[399]), .B(n11804), .Z(n13005) );
  NANDN U17391 ( .A(n11805), .B(creg[399]), .Z(n13004) );
  NAND U17392 ( .A(n13006), .B(n9081), .Z(n6785) );
  NANDN U17393 ( .A(init), .B(m[400]), .Z(n9081) );
  AND U17394 ( .A(n13007), .B(n13008), .Z(n13006) );
  NAND U17395 ( .A(o[400]), .B(n11804), .Z(n13008) );
  NANDN U17396 ( .A(n11805), .B(creg[400]), .Z(n13007) );
  NAND U17397 ( .A(n13009), .B(n9079), .Z(n6784) );
  NANDN U17398 ( .A(init), .B(m[401]), .Z(n9079) );
  AND U17399 ( .A(n13010), .B(n13011), .Z(n13009) );
  NAND U17400 ( .A(o[401]), .B(n11804), .Z(n13011) );
  NANDN U17401 ( .A(n11805), .B(creg[401]), .Z(n13010) );
  NAND U17402 ( .A(n13012), .B(n9077), .Z(n6783) );
  NANDN U17403 ( .A(init), .B(m[402]), .Z(n9077) );
  AND U17404 ( .A(n13013), .B(n13014), .Z(n13012) );
  NAND U17405 ( .A(o[402]), .B(n11804), .Z(n13014) );
  NANDN U17406 ( .A(n11805), .B(creg[402]), .Z(n13013) );
  NAND U17407 ( .A(n13015), .B(n9075), .Z(n6782) );
  NANDN U17408 ( .A(init), .B(m[403]), .Z(n9075) );
  AND U17409 ( .A(n13016), .B(n13017), .Z(n13015) );
  NAND U17410 ( .A(o[403]), .B(n11804), .Z(n13017) );
  NANDN U17411 ( .A(n11805), .B(creg[403]), .Z(n13016) );
  NAND U17412 ( .A(n13018), .B(n9073), .Z(n6781) );
  NANDN U17413 ( .A(init), .B(m[404]), .Z(n9073) );
  AND U17414 ( .A(n13019), .B(n13020), .Z(n13018) );
  NAND U17415 ( .A(o[404]), .B(n11804), .Z(n13020) );
  NANDN U17416 ( .A(n11805), .B(creg[404]), .Z(n13019) );
  NAND U17417 ( .A(n13021), .B(n9071), .Z(n6780) );
  NANDN U17418 ( .A(init), .B(m[405]), .Z(n9071) );
  AND U17419 ( .A(n13022), .B(n13023), .Z(n13021) );
  NAND U17420 ( .A(o[405]), .B(n11804), .Z(n13023) );
  NANDN U17421 ( .A(n11805), .B(creg[405]), .Z(n13022) );
  NAND U17422 ( .A(n13024), .B(n9069), .Z(n6779) );
  NANDN U17423 ( .A(init), .B(m[406]), .Z(n9069) );
  AND U17424 ( .A(n13025), .B(n13026), .Z(n13024) );
  NAND U17425 ( .A(o[406]), .B(n11804), .Z(n13026) );
  NANDN U17426 ( .A(n11805), .B(creg[406]), .Z(n13025) );
  NAND U17427 ( .A(n13027), .B(n9067), .Z(n6778) );
  NANDN U17428 ( .A(init), .B(m[407]), .Z(n9067) );
  AND U17429 ( .A(n13028), .B(n13029), .Z(n13027) );
  NAND U17430 ( .A(o[407]), .B(n11804), .Z(n13029) );
  NANDN U17431 ( .A(n11805), .B(creg[407]), .Z(n13028) );
  NAND U17432 ( .A(n13030), .B(n9065), .Z(n6777) );
  NANDN U17433 ( .A(init), .B(m[408]), .Z(n9065) );
  AND U17434 ( .A(n13031), .B(n13032), .Z(n13030) );
  NAND U17435 ( .A(o[408]), .B(n11804), .Z(n13032) );
  NANDN U17436 ( .A(n11805), .B(creg[408]), .Z(n13031) );
  NAND U17437 ( .A(n13033), .B(n9063), .Z(n6776) );
  NANDN U17438 ( .A(init), .B(m[409]), .Z(n9063) );
  AND U17439 ( .A(n13034), .B(n13035), .Z(n13033) );
  NAND U17440 ( .A(o[409]), .B(n11804), .Z(n13035) );
  NANDN U17441 ( .A(n11805), .B(creg[409]), .Z(n13034) );
  NAND U17442 ( .A(n13036), .B(n9059), .Z(n6775) );
  NANDN U17443 ( .A(init), .B(m[410]), .Z(n9059) );
  AND U17444 ( .A(n13037), .B(n13038), .Z(n13036) );
  NAND U17445 ( .A(o[410]), .B(n11804), .Z(n13038) );
  NANDN U17446 ( .A(n11805), .B(creg[410]), .Z(n13037) );
  NAND U17447 ( .A(n13039), .B(n9057), .Z(n6774) );
  NANDN U17448 ( .A(init), .B(m[411]), .Z(n9057) );
  AND U17449 ( .A(n13040), .B(n13041), .Z(n13039) );
  NAND U17450 ( .A(o[411]), .B(n11804), .Z(n13041) );
  NANDN U17451 ( .A(n11805), .B(creg[411]), .Z(n13040) );
  NAND U17452 ( .A(n13042), .B(n9055), .Z(n6773) );
  NANDN U17453 ( .A(init), .B(m[412]), .Z(n9055) );
  AND U17454 ( .A(n13043), .B(n13044), .Z(n13042) );
  NAND U17455 ( .A(o[412]), .B(n11804), .Z(n13044) );
  NANDN U17456 ( .A(n11805), .B(creg[412]), .Z(n13043) );
  NAND U17457 ( .A(n13045), .B(n9053), .Z(n6772) );
  NANDN U17458 ( .A(init), .B(m[413]), .Z(n9053) );
  AND U17459 ( .A(n13046), .B(n13047), .Z(n13045) );
  NAND U17460 ( .A(o[413]), .B(n11804), .Z(n13047) );
  NANDN U17461 ( .A(n11805), .B(creg[413]), .Z(n13046) );
  NAND U17462 ( .A(n13048), .B(n9051), .Z(n6771) );
  NANDN U17463 ( .A(init), .B(m[414]), .Z(n9051) );
  AND U17464 ( .A(n13049), .B(n13050), .Z(n13048) );
  NAND U17465 ( .A(o[414]), .B(n11804), .Z(n13050) );
  NANDN U17466 ( .A(n11805), .B(creg[414]), .Z(n13049) );
  NAND U17467 ( .A(n13051), .B(n9049), .Z(n6770) );
  NANDN U17468 ( .A(init), .B(m[415]), .Z(n9049) );
  AND U17469 ( .A(n13052), .B(n13053), .Z(n13051) );
  NAND U17470 ( .A(o[415]), .B(n11804), .Z(n13053) );
  NANDN U17471 ( .A(n11805), .B(creg[415]), .Z(n13052) );
  NAND U17472 ( .A(n13054), .B(n9047), .Z(n6769) );
  NANDN U17473 ( .A(init), .B(m[416]), .Z(n9047) );
  AND U17474 ( .A(n13055), .B(n13056), .Z(n13054) );
  NAND U17475 ( .A(o[416]), .B(n11804), .Z(n13056) );
  NANDN U17476 ( .A(n11805), .B(creg[416]), .Z(n13055) );
  NAND U17477 ( .A(n13057), .B(n9045), .Z(n6768) );
  NANDN U17478 ( .A(init), .B(m[417]), .Z(n9045) );
  AND U17479 ( .A(n13058), .B(n13059), .Z(n13057) );
  NAND U17480 ( .A(o[417]), .B(n11804), .Z(n13059) );
  NANDN U17481 ( .A(n11805), .B(creg[417]), .Z(n13058) );
  NAND U17482 ( .A(n13060), .B(n9043), .Z(n6767) );
  NANDN U17483 ( .A(init), .B(m[418]), .Z(n9043) );
  AND U17484 ( .A(n13061), .B(n13062), .Z(n13060) );
  NAND U17485 ( .A(o[418]), .B(n11804), .Z(n13062) );
  NANDN U17486 ( .A(n11805), .B(creg[418]), .Z(n13061) );
  NAND U17487 ( .A(n13063), .B(n9041), .Z(n6766) );
  NANDN U17488 ( .A(init), .B(m[419]), .Z(n9041) );
  AND U17489 ( .A(n13064), .B(n13065), .Z(n13063) );
  NAND U17490 ( .A(o[419]), .B(n11804), .Z(n13065) );
  NANDN U17491 ( .A(n11805), .B(creg[419]), .Z(n13064) );
  NAND U17492 ( .A(n13066), .B(n9037), .Z(n6765) );
  NANDN U17493 ( .A(init), .B(m[420]), .Z(n9037) );
  AND U17494 ( .A(n13067), .B(n13068), .Z(n13066) );
  NAND U17495 ( .A(o[420]), .B(n11804), .Z(n13068) );
  NANDN U17496 ( .A(n11805), .B(creg[420]), .Z(n13067) );
  NAND U17497 ( .A(n13069), .B(n9035), .Z(n6764) );
  NANDN U17498 ( .A(init), .B(m[421]), .Z(n9035) );
  AND U17499 ( .A(n13070), .B(n13071), .Z(n13069) );
  NAND U17500 ( .A(o[421]), .B(n11804), .Z(n13071) );
  NANDN U17501 ( .A(n11805), .B(creg[421]), .Z(n13070) );
  NAND U17502 ( .A(n13072), .B(n9033), .Z(n6763) );
  NANDN U17503 ( .A(init), .B(m[422]), .Z(n9033) );
  AND U17504 ( .A(n13073), .B(n13074), .Z(n13072) );
  NAND U17505 ( .A(o[422]), .B(n11804), .Z(n13074) );
  NANDN U17506 ( .A(n11805), .B(creg[422]), .Z(n13073) );
  NAND U17507 ( .A(n13075), .B(n9031), .Z(n6762) );
  NANDN U17508 ( .A(init), .B(m[423]), .Z(n9031) );
  AND U17509 ( .A(n13076), .B(n13077), .Z(n13075) );
  NAND U17510 ( .A(o[423]), .B(n11804), .Z(n13077) );
  NANDN U17511 ( .A(n11805), .B(creg[423]), .Z(n13076) );
  NAND U17512 ( .A(n13078), .B(n9029), .Z(n6761) );
  NANDN U17513 ( .A(init), .B(m[424]), .Z(n9029) );
  AND U17514 ( .A(n13079), .B(n13080), .Z(n13078) );
  NAND U17515 ( .A(o[424]), .B(n11804), .Z(n13080) );
  NANDN U17516 ( .A(n11805), .B(creg[424]), .Z(n13079) );
  NAND U17517 ( .A(n13081), .B(n9027), .Z(n6760) );
  NANDN U17518 ( .A(init), .B(m[425]), .Z(n9027) );
  AND U17519 ( .A(n13082), .B(n13083), .Z(n13081) );
  NAND U17520 ( .A(o[425]), .B(n11804), .Z(n13083) );
  NANDN U17521 ( .A(n11805), .B(creg[425]), .Z(n13082) );
  NAND U17522 ( .A(n13084), .B(n9025), .Z(n6759) );
  NANDN U17523 ( .A(init), .B(m[426]), .Z(n9025) );
  AND U17524 ( .A(n13085), .B(n13086), .Z(n13084) );
  NAND U17525 ( .A(o[426]), .B(n11804), .Z(n13086) );
  NANDN U17526 ( .A(n11805), .B(creg[426]), .Z(n13085) );
  NAND U17527 ( .A(n13087), .B(n9023), .Z(n6758) );
  NANDN U17528 ( .A(init), .B(m[427]), .Z(n9023) );
  AND U17529 ( .A(n13088), .B(n13089), .Z(n13087) );
  NAND U17530 ( .A(o[427]), .B(n11804), .Z(n13089) );
  NANDN U17531 ( .A(n11805), .B(creg[427]), .Z(n13088) );
  NAND U17532 ( .A(n13090), .B(n9021), .Z(n6757) );
  NANDN U17533 ( .A(init), .B(m[428]), .Z(n9021) );
  AND U17534 ( .A(n13091), .B(n13092), .Z(n13090) );
  NAND U17535 ( .A(o[428]), .B(n11804), .Z(n13092) );
  NANDN U17536 ( .A(n11805), .B(creg[428]), .Z(n13091) );
  NAND U17537 ( .A(n13093), .B(n9019), .Z(n6756) );
  NANDN U17538 ( .A(init), .B(m[429]), .Z(n9019) );
  AND U17539 ( .A(n13094), .B(n13095), .Z(n13093) );
  NAND U17540 ( .A(o[429]), .B(n11804), .Z(n13095) );
  NANDN U17541 ( .A(n11805), .B(creg[429]), .Z(n13094) );
  NAND U17542 ( .A(n13096), .B(n9015), .Z(n6755) );
  NANDN U17543 ( .A(init), .B(m[430]), .Z(n9015) );
  AND U17544 ( .A(n13097), .B(n13098), .Z(n13096) );
  NAND U17545 ( .A(o[430]), .B(n11804), .Z(n13098) );
  NANDN U17546 ( .A(n11805), .B(creg[430]), .Z(n13097) );
  NAND U17547 ( .A(n13099), .B(n9013), .Z(n6754) );
  NANDN U17548 ( .A(init), .B(m[431]), .Z(n9013) );
  AND U17549 ( .A(n13100), .B(n13101), .Z(n13099) );
  NAND U17550 ( .A(o[431]), .B(n11804), .Z(n13101) );
  NANDN U17551 ( .A(n11805), .B(creg[431]), .Z(n13100) );
  NAND U17552 ( .A(n13102), .B(n9011), .Z(n6753) );
  NANDN U17553 ( .A(init), .B(m[432]), .Z(n9011) );
  AND U17554 ( .A(n13103), .B(n13104), .Z(n13102) );
  NAND U17555 ( .A(o[432]), .B(n11804), .Z(n13104) );
  NANDN U17556 ( .A(n11805), .B(creg[432]), .Z(n13103) );
  NAND U17557 ( .A(n13105), .B(n9009), .Z(n6752) );
  NANDN U17558 ( .A(init), .B(m[433]), .Z(n9009) );
  AND U17559 ( .A(n13106), .B(n13107), .Z(n13105) );
  NAND U17560 ( .A(o[433]), .B(n11804), .Z(n13107) );
  NANDN U17561 ( .A(n11805), .B(creg[433]), .Z(n13106) );
  NAND U17562 ( .A(n13108), .B(n9007), .Z(n6751) );
  NANDN U17563 ( .A(init), .B(m[434]), .Z(n9007) );
  AND U17564 ( .A(n13109), .B(n13110), .Z(n13108) );
  NAND U17565 ( .A(o[434]), .B(n11804), .Z(n13110) );
  NANDN U17566 ( .A(n11805), .B(creg[434]), .Z(n13109) );
  NAND U17567 ( .A(n13111), .B(n9005), .Z(n6750) );
  NANDN U17568 ( .A(init), .B(m[435]), .Z(n9005) );
  AND U17569 ( .A(n13112), .B(n13113), .Z(n13111) );
  NAND U17570 ( .A(o[435]), .B(n11804), .Z(n13113) );
  NANDN U17571 ( .A(n11805), .B(creg[435]), .Z(n13112) );
  NAND U17572 ( .A(n13114), .B(n9003), .Z(n6749) );
  NANDN U17573 ( .A(init), .B(m[436]), .Z(n9003) );
  AND U17574 ( .A(n13115), .B(n13116), .Z(n13114) );
  NAND U17575 ( .A(o[436]), .B(n11804), .Z(n13116) );
  NANDN U17576 ( .A(n11805), .B(creg[436]), .Z(n13115) );
  NAND U17577 ( .A(n13117), .B(n9001), .Z(n6748) );
  NANDN U17578 ( .A(init), .B(m[437]), .Z(n9001) );
  AND U17579 ( .A(n13118), .B(n13119), .Z(n13117) );
  NAND U17580 ( .A(o[437]), .B(n11804), .Z(n13119) );
  NANDN U17581 ( .A(n11805), .B(creg[437]), .Z(n13118) );
  NAND U17582 ( .A(n13120), .B(n8999), .Z(n6747) );
  NANDN U17583 ( .A(init), .B(m[438]), .Z(n8999) );
  AND U17584 ( .A(n13121), .B(n13122), .Z(n13120) );
  NAND U17585 ( .A(o[438]), .B(n11804), .Z(n13122) );
  NANDN U17586 ( .A(n11805), .B(creg[438]), .Z(n13121) );
  NAND U17587 ( .A(n13123), .B(n8997), .Z(n6746) );
  NANDN U17588 ( .A(init), .B(m[439]), .Z(n8997) );
  AND U17589 ( .A(n13124), .B(n13125), .Z(n13123) );
  NAND U17590 ( .A(o[439]), .B(n11804), .Z(n13125) );
  NANDN U17591 ( .A(n11805), .B(creg[439]), .Z(n13124) );
  NAND U17592 ( .A(n13126), .B(n8993), .Z(n6745) );
  NANDN U17593 ( .A(init), .B(m[440]), .Z(n8993) );
  AND U17594 ( .A(n13127), .B(n13128), .Z(n13126) );
  NAND U17595 ( .A(o[440]), .B(n11804), .Z(n13128) );
  NANDN U17596 ( .A(n11805), .B(creg[440]), .Z(n13127) );
  NAND U17597 ( .A(n13129), .B(n8991), .Z(n6744) );
  NANDN U17598 ( .A(init), .B(m[441]), .Z(n8991) );
  AND U17599 ( .A(n13130), .B(n13131), .Z(n13129) );
  NAND U17600 ( .A(o[441]), .B(n11804), .Z(n13131) );
  NANDN U17601 ( .A(n11805), .B(creg[441]), .Z(n13130) );
  NAND U17602 ( .A(n13132), .B(n8989), .Z(n6743) );
  NANDN U17603 ( .A(init), .B(m[442]), .Z(n8989) );
  AND U17604 ( .A(n13133), .B(n13134), .Z(n13132) );
  NAND U17605 ( .A(o[442]), .B(n11804), .Z(n13134) );
  NANDN U17606 ( .A(n11805), .B(creg[442]), .Z(n13133) );
  NAND U17607 ( .A(n13135), .B(n8987), .Z(n6742) );
  NANDN U17608 ( .A(init), .B(m[443]), .Z(n8987) );
  AND U17609 ( .A(n13136), .B(n13137), .Z(n13135) );
  NAND U17610 ( .A(o[443]), .B(n11804), .Z(n13137) );
  NANDN U17611 ( .A(n11805), .B(creg[443]), .Z(n13136) );
  NAND U17612 ( .A(n13138), .B(n8985), .Z(n6741) );
  NANDN U17613 ( .A(init), .B(m[444]), .Z(n8985) );
  AND U17614 ( .A(n13139), .B(n13140), .Z(n13138) );
  NAND U17615 ( .A(o[444]), .B(n11804), .Z(n13140) );
  NANDN U17616 ( .A(n11805), .B(creg[444]), .Z(n13139) );
  NAND U17617 ( .A(n13141), .B(n8983), .Z(n6740) );
  NANDN U17618 ( .A(init), .B(m[445]), .Z(n8983) );
  AND U17619 ( .A(n13142), .B(n13143), .Z(n13141) );
  NAND U17620 ( .A(o[445]), .B(n11804), .Z(n13143) );
  NANDN U17621 ( .A(n11805), .B(creg[445]), .Z(n13142) );
  NAND U17622 ( .A(n13144), .B(n8981), .Z(n6739) );
  NANDN U17623 ( .A(init), .B(m[446]), .Z(n8981) );
  AND U17624 ( .A(n13145), .B(n13146), .Z(n13144) );
  NAND U17625 ( .A(o[446]), .B(n11804), .Z(n13146) );
  NANDN U17626 ( .A(n11805), .B(creg[446]), .Z(n13145) );
  NAND U17627 ( .A(n13147), .B(n8979), .Z(n6738) );
  NANDN U17628 ( .A(init), .B(m[447]), .Z(n8979) );
  AND U17629 ( .A(n13148), .B(n13149), .Z(n13147) );
  NAND U17630 ( .A(o[447]), .B(n11804), .Z(n13149) );
  NANDN U17631 ( .A(n11805), .B(creg[447]), .Z(n13148) );
  NAND U17632 ( .A(n13150), .B(n8977), .Z(n6737) );
  NANDN U17633 ( .A(init), .B(m[448]), .Z(n8977) );
  AND U17634 ( .A(n13151), .B(n13152), .Z(n13150) );
  NAND U17635 ( .A(o[448]), .B(n11804), .Z(n13152) );
  NANDN U17636 ( .A(n11805), .B(creg[448]), .Z(n13151) );
  NAND U17637 ( .A(n13153), .B(n8975), .Z(n6736) );
  NANDN U17638 ( .A(init), .B(m[449]), .Z(n8975) );
  AND U17639 ( .A(n13154), .B(n13155), .Z(n13153) );
  NAND U17640 ( .A(o[449]), .B(n11804), .Z(n13155) );
  NANDN U17641 ( .A(n11805), .B(creg[449]), .Z(n13154) );
  NAND U17642 ( .A(n13156), .B(n8971), .Z(n6735) );
  NANDN U17643 ( .A(init), .B(m[450]), .Z(n8971) );
  AND U17644 ( .A(n13157), .B(n13158), .Z(n13156) );
  NAND U17645 ( .A(o[450]), .B(n11804), .Z(n13158) );
  NANDN U17646 ( .A(n11805), .B(creg[450]), .Z(n13157) );
  NAND U17647 ( .A(n13159), .B(n8969), .Z(n6734) );
  NANDN U17648 ( .A(init), .B(m[451]), .Z(n8969) );
  AND U17649 ( .A(n13160), .B(n13161), .Z(n13159) );
  NAND U17650 ( .A(o[451]), .B(n11804), .Z(n13161) );
  NANDN U17651 ( .A(n11805), .B(creg[451]), .Z(n13160) );
  NAND U17652 ( .A(n13162), .B(n8967), .Z(n6733) );
  NANDN U17653 ( .A(init), .B(m[452]), .Z(n8967) );
  AND U17654 ( .A(n13163), .B(n13164), .Z(n13162) );
  NAND U17655 ( .A(o[452]), .B(n11804), .Z(n13164) );
  NANDN U17656 ( .A(n11805), .B(creg[452]), .Z(n13163) );
  NAND U17657 ( .A(n13165), .B(n8965), .Z(n6732) );
  NANDN U17658 ( .A(init), .B(m[453]), .Z(n8965) );
  AND U17659 ( .A(n13166), .B(n13167), .Z(n13165) );
  NAND U17660 ( .A(o[453]), .B(n11804), .Z(n13167) );
  NANDN U17661 ( .A(n11805), .B(creg[453]), .Z(n13166) );
  NAND U17662 ( .A(n13168), .B(n8963), .Z(n6731) );
  NANDN U17663 ( .A(init), .B(m[454]), .Z(n8963) );
  AND U17664 ( .A(n13169), .B(n13170), .Z(n13168) );
  NAND U17665 ( .A(o[454]), .B(n11804), .Z(n13170) );
  NANDN U17666 ( .A(n11805), .B(creg[454]), .Z(n13169) );
  NAND U17667 ( .A(n13171), .B(n8961), .Z(n6730) );
  NANDN U17668 ( .A(init), .B(m[455]), .Z(n8961) );
  AND U17669 ( .A(n13172), .B(n13173), .Z(n13171) );
  NAND U17670 ( .A(o[455]), .B(n11804), .Z(n13173) );
  NANDN U17671 ( .A(n11805), .B(creg[455]), .Z(n13172) );
  NAND U17672 ( .A(n13174), .B(n8959), .Z(n6729) );
  NANDN U17673 ( .A(init), .B(m[456]), .Z(n8959) );
  AND U17674 ( .A(n13175), .B(n13176), .Z(n13174) );
  NAND U17675 ( .A(o[456]), .B(n11804), .Z(n13176) );
  NANDN U17676 ( .A(n11805), .B(creg[456]), .Z(n13175) );
  NAND U17677 ( .A(n13177), .B(n8957), .Z(n6728) );
  NANDN U17678 ( .A(init), .B(m[457]), .Z(n8957) );
  AND U17679 ( .A(n13178), .B(n13179), .Z(n13177) );
  NAND U17680 ( .A(o[457]), .B(n11804), .Z(n13179) );
  NANDN U17681 ( .A(n11805), .B(creg[457]), .Z(n13178) );
  NAND U17682 ( .A(n13180), .B(n8955), .Z(n6727) );
  NANDN U17683 ( .A(init), .B(m[458]), .Z(n8955) );
  AND U17684 ( .A(n13181), .B(n13182), .Z(n13180) );
  NAND U17685 ( .A(o[458]), .B(n11804), .Z(n13182) );
  NANDN U17686 ( .A(n11805), .B(creg[458]), .Z(n13181) );
  NAND U17687 ( .A(n13183), .B(n8953), .Z(n6726) );
  NANDN U17688 ( .A(init), .B(m[459]), .Z(n8953) );
  AND U17689 ( .A(n13184), .B(n13185), .Z(n13183) );
  NAND U17690 ( .A(o[459]), .B(n11804), .Z(n13185) );
  NANDN U17691 ( .A(n11805), .B(creg[459]), .Z(n13184) );
  NAND U17692 ( .A(n13186), .B(n8949), .Z(n6725) );
  NANDN U17693 ( .A(init), .B(m[460]), .Z(n8949) );
  AND U17694 ( .A(n13187), .B(n13188), .Z(n13186) );
  NAND U17695 ( .A(o[460]), .B(n11804), .Z(n13188) );
  NANDN U17696 ( .A(n11805), .B(creg[460]), .Z(n13187) );
  NAND U17697 ( .A(n13189), .B(n8947), .Z(n6724) );
  NANDN U17698 ( .A(init), .B(m[461]), .Z(n8947) );
  AND U17699 ( .A(n13190), .B(n13191), .Z(n13189) );
  NAND U17700 ( .A(o[461]), .B(n11804), .Z(n13191) );
  NANDN U17701 ( .A(n11805), .B(creg[461]), .Z(n13190) );
  NAND U17702 ( .A(n13192), .B(n8945), .Z(n6723) );
  NANDN U17703 ( .A(init), .B(m[462]), .Z(n8945) );
  AND U17704 ( .A(n13193), .B(n13194), .Z(n13192) );
  NAND U17705 ( .A(o[462]), .B(n11804), .Z(n13194) );
  NANDN U17706 ( .A(n11805), .B(creg[462]), .Z(n13193) );
  NAND U17707 ( .A(n13195), .B(n8943), .Z(n6722) );
  NANDN U17708 ( .A(init), .B(m[463]), .Z(n8943) );
  AND U17709 ( .A(n13196), .B(n13197), .Z(n13195) );
  NAND U17710 ( .A(o[463]), .B(n11804), .Z(n13197) );
  NANDN U17711 ( .A(n11805), .B(creg[463]), .Z(n13196) );
  NAND U17712 ( .A(n13198), .B(n8941), .Z(n6721) );
  NANDN U17713 ( .A(init), .B(m[464]), .Z(n8941) );
  AND U17714 ( .A(n13199), .B(n13200), .Z(n13198) );
  NAND U17715 ( .A(o[464]), .B(n11804), .Z(n13200) );
  NANDN U17716 ( .A(n11805), .B(creg[464]), .Z(n13199) );
  NAND U17717 ( .A(n13201), .B(n8939), .Z(n6720) );
  NANDN U17718 ( .A(init), .B(m[465]), .Z(n8939) );
  AND U17719 ( .A(n13202), .B(n13203), .Z(n13201) );
  NAND U17720 ( .A(o[465]), .B(n11804), .Z(n13203) );
  NANDN U17721 ( .A(n11805), .B(creg[465]), .Z(n13202) );
  NAND U17722 ( .A(n13204), .B(n8937), .Z(n6719) );
  NANDN U17723 ( .A(init), .B(m[466]), .Z(n8937) );
  AND U17724 ( .A(n13205), .B(n13206), .Z(n13204) );
  NAND U17725 ( .A(o[466]), .B(n11804), .Z(n13206) );
  NANDN U17726 ( .A(n11805), .B(creg[466]), .Z(n13205) );
  NAND U17727 ( .A(n13207), .B(n8935), .Z(n6718) );
  NANDN U17728 ( .A(init), .B(m[467]), .Z(n8935) );
  AND U17729 ( .A(n13208), .B(n13209), .Z(n13207) );
  NAND U17730 ( .A(o[467]), .B(n11804), .Z(n13209) );
  NANDN U17731 ( .A(n11805), .B(creg[467]), .Z(n13208) );
  NAND U17732 ( .A(n13210), .B(n8933), .Z(n6717) );
  NANDN U17733 ( .A(init), .B(m[468]), .Z(n8933) );
  AND U17734 ( .A(n13211), .B(n13212), .Z(n13210) );
  NAND U17735 ( .A(o[468]), .B(n11804), .Z(n13212) );
  NANDN U17736 ( .A(n11805), .B(creg[468]), .Z(n13211) );
  NAND U17737 ( .A(n13213), .B(n8931), .Z(n6716) );
  NANDN U17738 ( .A(init), .B(m[469]), .Z(n8931) );
  AND U17739 ( .A(n13214), .B(n13215), .Z(n13213) );
  NAND U17740 ( .A(o[469]), .B(n11804), .Z(n13215) );
  NANDN U17741 ( .A(n11805), .B(creg[469]), .Z(n13214) );
  NAND U17742 ( .A(n13216), .B(n8927), .Z(n6715) );
  NANDN U17743 ( .A(init), .B(m[470]), .Z(n8927) );
  AND U17744 ( .A(n13217), .B(n13218), .Z(n13216) );
  NAND U17745 ( .A(o[470]), .B(n11804), .Z(n13218) );
  NANDN U17746 ( .A(n11805), .B(creg[470]), .Z(n13217) );
  NAND U17747 ( .A(n13219), .B(n8925), .Z(n6714) );
  NANDN U17748 ( .A(init), .B(m[471]), .Z(n8925) );
  AND U17749 ( .A(n13220), .B(n13221), .Z(n13219) );
  NAND U17750 ( .A(o[471]), .B(n11804), .Z(n13221) );
  NANDN U17751 ( .A(n11805), .B(creg[471]), .Z(n13220) );
  NAND U17752 ( .A(n13222), .B(n8923), .Z(n6713) );
  NANDN U17753 ( .A(init), .B(m[472]), .Z(n8923) );
  AND U17754 ( .A(n13223), .B(n13224), .Z(n13222) );
  NAND U17755 ( .A(o[472]), .B(n11804), .Z(n13224) );
  NANDN U17756 ( .A(n11805), .B(creg[472]), .Z(n13223) );
  NAND U17757 ( .A(n13225), .B(n8921), .Z(n6712) );
  NANDN U17758 ( .A(init), .B(m[473]), .Z(n8921) );
  AND U17759 ( .A(n13226), .B(n13227), .Z(n13225) );
  NAND U17760 ( .A(o[473]), .B(n11804), .Z(n13227) );
  NANDN U17761 ( .A(n11805), .B(creg[473]), .Z(n13226) );
  NAND U17762 ( .A(n13228), .B(n8919), .Z(n6711) );
  NANDN U17763 ( .A(init), .B(m[474]), .Z(n8919) );
  AND U17764 ( .A(n13229), .B(n13230), .Z(n13228) );
  NAND U17765 ( .A(o[474]), .B(n11804), .Z(n13230) );
  NANDN U17766 ( .A(n11805), .B(creg[474]), .Z(n13229) );
  NAND U17767 ( .A(n13231), .B(n8917), .Z(n6710) );
  NANDN U17768 ( .A(init), .B(m[475]), .Z(n8917) );
  AND U17769 ( .A(n13232), .B(n13233), .Z(n13231) );
  NAND U17770 ( .A(o[475]), .B(n11804), .Z(n13233) );
  NANDN U17771 ( .A(n11805), .B(creg[475]), .Z(n13232) );
  NAND U17772 ( .A(n13234), .B(n8915), .Z(n6709) );
  NANDN U17773 ( .A(init), .B(m[476]), .Z(n8915) );
  AND U17774 ( .A(n13235), .B(n13236), .Z(n13234) );
  NAND U17775 ( .A(o[476]), .B(n11804), .Z(n13236) );
  NANDN U17776 ( .A(n11805), .B(creg[476]), .Z(n13235) );
  NAND U17777 ( .A(n13237), .B(n8913), .Z(n6708) );
  NANDN U17778 ( .A(init), .B(m[477]), .Z(n8913) );
  AND U17779 ( .A(n13238), .B(n13239), .Z(n13237) );
  NAND U17780 ( .A(o[477]), .B(n11804), .Z(n13239) );
  NANDN U17781 ( .A(n11805), .B(creg[477]), .Z(n13238) );
  NAND U17782 ( .A(n13240), .B(n8911), .Z(n6707) );
  NANDN U17783 ( .A(init), .B(m[478]), .Z(n8911) );
  AND U17784 ( .A(n13241), .B(n13242), .Z(n13240) );
  NAND U17785 ( .A(o[478]), .B(n11804), .Z(n13242) );
  NANDN U17786 ( .A(n11805), .B(creg[478]), .Z(n13241) );
  NAND U17787 ( .A(n13243), .B(n8909), .Z(n6706) );
  NANDN U17788 ( .A(init), .B(m[479]), .Z(n8909) );
  AND U17789 ( .A(n13244), .B(n13245), .Z(n13243) );
  NAND U17790 ( .A(o[479]), .B(n11804), .Z(n13245) );
  NANDN U17791 ( .A(n11805), .B(creg[479]), .Z(n13244) );
  NAND U17792 ( .A(n13246), .B(n8905), .Z(n6705) );
  NANDN U17793 ( .A(init), .B(m[480]), .Z(n8905) );
  AND U17794 ( .A(n13247), .B(n13248), .Z(n13246) );
  NAND U17795 ( .A(o[480]), .B(n11804), .Z(n13248) );
  NANDN U17796 ( .A(n11805), .B(creg[480]), .Z(n13247) );
  NAND U17797 ( .A(n13249), .B(n8903), .Z(n6704) );
  NANDN U17798 ( .A(init), .B(m[481]), .Z(n8903) );
  AND U17799 ( .A(n13250), .B(n13251), .Z(n13249) );
  NAND U17800 ( .A(o[481]), .B(n11804), .Z(n13251) );
  NANDN U17801 ( .A(n11805), .B(creg[481]), .Z(n13250) );
  NAND U17802 ( .A(n13252), .B(n8901), .Z(n6703) );
  NANDN U17803 ( .A(init), .B(m[482]), .Z(n8901) );
  AND U17804 ( .A(n13253), .B(n13254), .Z(n13252) );
  NAND U17805 ( .A(o[482]), .B(n11804), .Z(n13254) );
  NANDN U17806 ( .A(n11805), .B(creg[482]), .Z(n13253) );
  NAND U17807 ( .A(n13255), .B(n8899), .Z(n6702) );
  NANDN U17808 ( .A(init), .B(m[483]), .Z(n8899) );
  AND U17809 ( .A(n13256), .B(n13257), .Z(n13255) );
  NAND U17810 ( .A(o[483]), .B(n11804), .Z(n13257) );
  NANDN U17811 ( .A(n11805), .B(creg[483]), .Z(n13256) );
  NAND U17812 ( .A(n13258), .B(n8897), .Z(n6701) );
  NANDN U17813 ( .A(init), .B(m[484]), .Z(n8897) );
  AND U17814 ( .A(n13259), .B(n13260), .Z(n13258) );
  NAND U17815 ( .A(o[484]), .B(n11804), .Z(n13260) );
  NANDN U17816 ( .A(n11805), .B(creg[484]), .Z(n13259) );
  NAND U17817 ( .A(n13261), .B(n8895), .Z(n6700) );
  NANDN U17818 ( .A(init), .B(m[485]), .Z(n8895) );
  AND U17819 ( .A(n13262), .B(n13263), .Z(n13261) );
  NAND U17820 ( .A(o[485]), .B(n11804), .Z(n13263) );
  NANDN U17821 ( .A(n11805), .B(creg[485]), .Z(n13262) );
  NAND U17822 ( .A(n13264), .B(n8893), .Z(n6699) );
  NANDN U17823 ( .A(init), .B(m[486]), .Z(n8893) );
  AND U17824 ( .A(n13265), .B(n13266), .Z(n13264) );
  NAND U17825 ( .A(o[486]), .B(n11804), .Z(n13266) );
  NANDN U17826 ( .A(n11805), .B(creg[486]), .Z(n13265) );
  NAND U17827 ( .A(n13267), .B(n8891), .Z(n6698) );
  NANDN U17828 ( .A(init), .B(m[487]), .Z(n8891) );
  AND U17829 ( .A(n13268), .B(n13269), .Z(n13267) );
  NAND U17830 ( .A(o[487]), .B(n11804), .Z(n13269) );
  NANDN U17831 ( .A(n11805), .B(creg[487]), .Z(n13268) );
  NAND U17832 ( .A(n13270), .B(n8889), .Z(n6697) );
  NANDN U17833 ( .A(init), .B(m[488]), .Z(n8889) );
  AND U17834 ( .A(n13271), .B(n13272), .Z(n13270) );
  NAND U17835 ( .A(o[488]), .B(n11804), .Z(n13272) );
  NANDN U17836 ( .A(n11805), .B(creg[488]), .Z(n13271) );
  NAND U17837 ( .A(n13273), .B(n8887), .Z(n6696) );
  NANDN U17838 ( .A(init), .B(m[489]), .Z(n8887) );
  AND U17839 ( .A(n13274), .B(n13275), .Z(n13273) );
  NAND U17840 ( .A(o[489]), .B(n11804), .Z(n13275) );
  NANDN U17841 ( .A(n11805), .B(creg[489]), .Z(n13274) );
  NAND U17842 ( .A(n13276), .B(n8883), .Z(n6695) );
  NANDN U17843 ( .A(init), .B(m[490]), .Z(n8883) );
  AND U17844 ( .A(n13277), .B(n13278), .Z(n13276) );
  NAND U17845 ( .A(o[490]), .B(n11804), .Z(n13278) );
  NANDN U17846 ( .A(n11805), .B(creg[490]), .Z(n13277) );
  NAND U17847 ( .A(n13279), .B(n8881), .Z(n6694) );
  NANDN U17848 ( .A(init), .B(m[491]), .Z(n8881) );
  AND U17849 ( .A(n13280), .B(n13281), .Z(n13279) );
  NAND U17850 ( .A(o[491]), .B(n11804), .Z(n13281) );
  NANDN U17851 ( .A(n11805), .B(creg[491]), .Z(n13280) );
  NAND U17852 ( .A(n13282), .B(n8879), .Z(n6693) );
  NANDN U17853 ( .A(init), .B(m[492]), .Z(n8879) );
  AND U17854 ( .A(n13283), .B(n13284), .Z(n13282) );
  NAND U17855 ( .A(o[492]), .B(n11804), .Z(n13284) );
  NANDN U17856 ( .A(n11805), .B(creg[492]), .Z(n13283) );
  NAND U17857 ( .A(n13285), .B(n8877), .Z(n6692) );
  NANDN U17858 ( .A(init), .B(m[493]), .Z(n8877) );
  AND U17859 ( .A(n13286), .B(n13287), .Z(n13285) );
  NAND U17860 ( .A(o[493]), .B(n11804), .Z(n13287) );
  NANDN U17861 ( .A(n11805), .B(creg[493]), .Z(n13286) );
  NAND U17862 ( .A(n13288), .B(n8875), .Z(n6691) );
  NANDN U17863 ( .A(init), .B(m[494]), .Z(n8875) );
  AND U17864 ( .A(n13289), .B(n13290), .Z(n13288) );
  NAND U17865 ( .A(o[494]), .B(n11804), .Z(n13290) );
  NANDN U17866 ( .A(n11805), .B(creg[494]), .Z(n13289) );
  NAND U17867 ( .A(n13291), .B(n8873), .Z(n6690) );
  NANDN U17868 ( .A(init), .B(m[495]), .Z(n8873) );
  AND U17869 ( .A(n13292), .B(n13293), .Z(n13291) );
  NAND U17870 ( .A(o[495]), .B(n11804), .Z(n13293) );
  NANDN U17871 ( .A(n11805), .B(creg[495]), .Z(n13292) );
  NAND U17872 ( .A(n13294), .B(n8871), .Z(n6689) );
  NANDN U17873 ( .A(init), .B(m[496]), .Z(n8871) );
  AND U17874 ( .A(n13295), .B(n13296), .Z(n13294) );
  NAND U17875 ( .A(o[496]), .B(n11804), .Z(n13296) );
  NANDN U17876 ( .A(n11805), .B(creg[496]), .Z(n13295) );
  NAND U17877 ( .A(n13297), .B(n8869), .Z(n6688) );
  NANDN U17878 ( .A(init), .B(m[497]), .Z(n8869) );
  AND U17879 ( .A(n13298), .B(n13299), .Z(n13297) );
  NAND U17880 ( .A(o[497]), .B(n11804), .Z(n13299) );
  NANDN U17881 ( .A(n11805), .B(creg[497]), .Z(n13298) );
  NAND U17882 ( .A(n13300), .B(n8867), .Z(n6687) );
  NANDN U17883 ( .A(init), .B(m[498]), .Z(n8867) );
  AND U17884 ( .A(n13301), .B(n13302), .Z(n13300) );
  NAND U17885 ( .A(o[498]), .B(n11804), .Z(n13302) );
  NANDN U17886 ( .A(n11805), .B(creg[498]), .Z(n13301) );
  NAND U17887 ( .A(n13303), .B(n8865), .Z(n6686) );
  NANDN U17888 ( .A(init), .B(m[499]), .Z(n8865) );
  AND U17889 ( .A(n13304), .B(n13305), .Z(n13303) );
  NAND U17890 ( .A(o[499]), .B(n11804), .Z(n13305) );
  NANDN U17891 ( .A(n11805), .B(creg[499]), .Z(n13304) );
  NAND U17892 ( .A(n13306), .B(n8859), .Z(n6685) );
  NANDN U17893 ( .A(init), .B(m[500]), .Z(n8859) );
  AND U17894 ( .A(n13307), .B(n13308), .Z(n13306) );
  NAND U17895 ( .A(o[500]), .B(n11804), .Z(n13308) );
  NANDN U17896 ( .A(n11805), .B(creg[500]), .Z(n13307) );
  NAND U17897 ( .A(n13309), .B(n8857), .Z(n6684) );
  NANDN U17898 ( .A(init), .B(m[501]), .Z(n8857) );
  AND U17899 ( .A(n13310), .B(n13311), .Z(n13309) );
  NAND U17900 ( .A(o[501]), .B(n11804), .Z(n13311) );
  NANDN U17901 ( .A(n11805), .B(creg[501]), .Z(n13310) );
  NAND U17902 ( .A(n13312), .B(n8855), .Z(n6683) );
  NANDN U17903 ( .A(init), .B(m[502]), .Z(n8855) );
  AND U17904 ( .A(n13313), .B(n13314), .Z(n13312) );
  NAND U17905 ( .A(o[502]), .B(n11804), .Z(n13314) );
  NANDN U17906 ( .A(n11805), .B(creg[502]), .Z(n13313) );
  NAND U17907 ( .A(n13315), .B(n8853), .Z(n6682) );
  NANDN U17908 ( .A(init), .B(m[503]), .Z(n8853) );
  AND U17909 ( .A(n13316), .B(n13317), .Z(n13315) );
  NAND U17910 ( .A(o[503]), .B(n11804), .Z(n13317) );
  NANDN U17911 ( .A(n11805), .B(creg[503]), .Z(n13316) );
  NAND U17912 ( .A(n13318), .B(n8851), .Z(n6681) );
  NANDN U17913 ( .A(init), .B(m[504]), .Z(n8851) );
  AND U17914 ( .A(n13319), .B(n13320), .Z(n13318) );
  NAND U17915 ( .A(o[504]), .B(n11804), .Z(n13320) );
  NANDN U17916 ( .A(n11805), .B(creg[504]), .Z(n13319) );
  NAND U17917 ( .A(n13321), .B(n8849), .Z(n6680) );
  NANDN U17918 ( .A(init), .B(m[505]), .Z(n8849) );
  AND U17919 ( .A(n13322), .B(n13323), .Z(n13321) );
  NAND U17920 ( .A(o[505]), .B(n11804), .Z(n13323) );
  NANDN U17921 ( .A(n11805), .B(creg[505]), .Z(n13322) );
  NAND U17922 ( .A(n13324), .B(n8847), .Z(n6679) );
  NANDN U17923 ( .A(init), .B(m[506]), .Z(n8847) );
  AND U17924 ( .A(n13325), .B(n13326), .Z(n13324) );
  NAND U17925 ( .A(o[506]), .B(n11804), .Z(n13326) );
  NANDN U17926 ( .A(n11805), .B(creg[506]), .Z(n13325) );
  NAND U17927 ( .A(n13327), .B(n8845), .Z(n6678) );
  NANDN U17928 ( .A(init), .B(m[507]), .Z(n8845) );
  AND U17929 ( .A(n13328), .B(n13329), .Z(n13327) );
  NAND U17930 ( .A(o[507]), .B(n11804), .Z(n13329) );
  NANDN U17931 ( .A(n11805), .B(creg[507]), .Z(n13328) );
  NAND U17932 ( .A(n13330), .B(n8843), .Z(n6677) );
  NANDN U17933 ( .A(init), .B(m[508]), .Z(n8843) );
  AND U17934 ( .A(n13331), .B(n13332), .Z(n13330) );
  NAND U17935 ( .A(o[508]), .B(n11804), .Z(n13332) );
  NANDN U17936 ( .A(n11805), .B(creg[508]), .Z(n13331) );
  NAND U17937 ( .A(n13333), .B(n8841), .Z(n6676) );
  NANDN U17938 ( .A(init), .B(m[509]), .Z(n8841) );
  AND U17939 ( .A(n13334), .B(n13335), .Z(n13333) );
  NAND U17940 ( .A(o[509]), .B(n11804), .Z(n13335) );
  NANDN U17941 ( .A(n11805), .B(creg[509]), .Z(n13334) );
  NAND U17942 ( .A(n13336), .B(n8837), .Z(n6675) );
  NANDN U17943 ( .A(init), .B(m[510]), .Z(n8837) );
  AND U17944 ( .A(n13337), .B(n13338), .Z(n13336) );
  NAND U17945 ( .A(o[510]), .B(n11804), .Z(n13338) );
  AND U17946 ( .A(n14372), .B(n11805), .Z(n11804) );
  NANDN U17947 ( .A(n11805), .B(creg[510]), .Z(n13337) );
  NAND U17948 ( .A(init), .B(n13339), .Z(n11805) );
  NAND U17949 ( .A(first_one), .B(n13340), .Z(n13339) );
  AND U17950 ( .A(start_reg[511]), .B(n13341), .Z(n13340) );
  NAND U17951 ( .A(n13342), .B(mul_pow), .Z(n13341) );
  NANDN U17952 ( .A(first_one), .B(n13343), .Z(n6674) );
  NAND U17953 ( .A(n13344), .B(ereg[511]), .Z(n13343) );
  AND U17954 ( .A(n14372), .B(mul_pow), .Z(n13344) );
  AND U17955 ( .A(start_reg[511]), .B(init), .Z(n14372) );
  NAND U17956 ( .A(n13345), .B(n13346), .Z(c[9]) );
  NAND U17957 ( .A(n13347), .B(o[9]), .Z(n13346) );
  NAND U17958 ( .A(n13342), .B(creg[9]), .Z(n13345) );
  NAND U17959 ( .A(n13348), .B(n13349), .Z(c[99]) );
  NAND U17960 ( .A(n13347), .B(o[99]), .Z(n13349) );
  NAND U17961 ( .A(n13342), .B(creg[99]), .Z(n13348) );
  NAND U17962 ( .A(n13350), .B(n13351), .Z(c[98]) );
  NAND U17963 ( .A(n13347), .B(o[98]), .Z(n13351) );
  NAND U17964 ( .A(n13342), .B(creg[98]), .Z(n13350) );
  NAND U17965 ( .A(n13352), .B(n13353), .Z(c[97]) );
  NAND U17966 ( .A(n13347), .B(o[97]), .Z(n13353) );
  NAND U17967 ( .A(n13342), .B(creg[97]), .Z(n13352) );
  NAND U17968 ( .A(n13354), .B(n13355), .Z(c[96]) );
  NAND U17969 ( .A(n13347), .B(o[96]), .Z(n13355) );
  NAND U17970 ( .A(n13342), .B(creg[96]), .Z(n13354) );
  NAND U17971 ( .A(n13356), .B(n13357), .Z(c[95]) );
  NAND U17972 ( .A(n13347), .B(o[95]), .Z(n13357) );
  NAND U17973 ( .A(n13342), .B(creg[95]), .Z(n13356) );
  NAND U17974 ( .A(n13358), .B(n13359), .Z(c[94]) );
  NAND U17975 ( .A(n13347), .B(o[94]), .Z(n13359) );
  NAND U17976 ( .A(n13342), .B(creg[94]), .Z(n13358) );
  NAND U17977 ( .A(n13360), .B(n13361), .Z(c[93]) );
  NAND U17978 ( .A(n13347), .B(o[93]), .Z(n13361) );
  NAND U17979 ( .A(n13342), .B(creg[93]), .Z(n13360) );
  NAND U17980 ( .A(n13362), .B(n13363), .Z(c[92]) );
  NAND U17981 ( .A(n13347), .B(o[92]), .Z(n13363) );
  NAND U17982 ( .A(n13342), .B(creg[92]), .Z(n13362) );
  NAND U17983 ( .A(n13364), .B(n13365), .Z(c[91]) );
  NAND U17984 ( .A(n13347), .B(o[91]), .Z(n13365) );
  NAND U17985 ( .A(n13342), .B(creg[91]), .Z(n13364) );
  NAND U17986 ( .A(n13366), .B(n13367), .Z(c[90]) );
  NAND U17987 ( .A(n13347), .B(o[90]), .Z(n13367) );
  NAND U17988 ( .A(n13342), .B(creg[90]), .Z(n13366) );
  NAND U17989 ( .A(n13368), .B(n13369), .Z(c[8]) );
  NAND U17990 ( .A(n13347), .B(o[8]), .Z(n13369) );
  NAND U17991 ( .A(n13342), .B(creg[8]), .Z(n13368) );
  NAND U17992 ( .A(n13370), .B(n13371), .Z(c[89]) );
  NAND U17993 ( .A(n13347), .B(o[89]), .Z(n13371) );
  NAND U17994 ( .A(n13342), .B(creg[89]), .Z(n13370) );
  NAND U17995 ( .A(n13372), .B(n13373), .Z(c[88]) );
  NAND U17996 ( .A(n13347), .B(o[88]), .Z(n13373) );
  NAND U17997 ( .A(n13342), .B(creg[88]), .Z(n13372) );
  NAND U17998 ( .A(n13374), .B(n13375), .Z(c[87]) );
  NAND U17999 ( .A(n13347), .B(o[87]), .Z(n13375) );
  NAND U18000 ( .A(n13342), .B(creg[87]), .Z(n13374) );
  NAND U18001 ( .A(n13376), .B(n13377), .Z(c[86]) );
  NAND U18002 ( .A(n13347), .B(o[86]), .Z(n13377) );
  NAND U18003 ( .A(n13342), .B(creg[86]), .Z(n13376) );
  NAND U18004 ( .A(n13378), .B(n13379), .Z(c[85]) );
  NAND U18005 ( .A(n13347), .B(o[85]), .Z(n13379) );
  NAND U18006 ( .A(n13342), .B(creg[85]), .Z(n13378) );
  NAND U18007 ( .A(n13380), .B(n13381), .Z(c[84]) );
  NAND U18008 ( .A(n13347), .B(o[84]), .Z(n13381) );
  NAND U18009 ( .A(n13342), .B(creg[84]), .Z(n13380) );
  NAND U18010 ( .A(n13382), .B(n13383), .Z(c[83]) );
  NAND U18011 ( .A(n13347), .B(o[83]), .Z(n13383) );
  NAND U18012 ( .A(n13342), .B(creg[83]), .Z(n13382) );
  NAND U18013 ( .A(n13384), .B(n13385), .Z(c[82]) );
  NAND U18014 ( .A(n13347), .B(o[82]), .Z(n13385) );
  NAND U18015 ( .A(n13342), .B(creg[82]), .Z(n13384) );
  NAND U18016 ( .A(n13386), .B(n13387), .Z(c[81]) );
  NAND U18017 ( .A(n13347), .B(o[81]), .Z(n13387) );
  NAND U18018 ( .A(n13342), .B(creg[81]), .Z(n13386) );
  NAND U18019 ( .A(n13388), .B(n13389), .Z(c[80]) );
  NAND U18020 ( .A(n13347), .B(o[80]), .Z(n13389) );
  NAND U18021 ( .A(n13342), .B(creg[80]), .Z(n13388) );
  NAND U18022 ( .A(n13390), .B(n13391), .Z(c[7]) );
  NAND U18023 ( .A(n13347), .B(o[7]), .Z(n13391) );
  NAND U18024 ( .A(n13342), .B(creg[7]), .Z(n13390) );
  NAND U18025 ( .A(n13392), .B(n13393), .Z(c[79]) );
  NAND U18026 ( .A(n13347), .B(o[79]), .Z(n13393) );
  NAND U18027 ( .A(n13342), .B(creg[79]), .Z(n13392) );
  NAND U18028 ( .A(n13394), .B(n13395), .Z(c[78]) );
  NAND U18029 ( .A(n13347), .B(o[78]), .Z(n13395) );
  NAND U18030 ( .A(n13342), .B(creg[78]), .Z(n13394) );
  NAND U18031 ( .A(n13396), .B(n13397), .Z(c[77]) );
  NAND U18032 ( .A(n13347), .B(o[77]), .Z(n13397) );
  NAND U18033 ( .A(n13342), .B(creg[77]), .Z(n13396) );
  NAND U18034 ( .A(n13398), .B(n13399), .Z(c[76]) );
  NAND U18035 ( .A(n13347), .B(o[76]), .Z(n13399) );
  NAND U18036 ( .A(n13342), .B(creg[76]), .Z(n13398) );
  NAND U18037 ( .A(n13400), .B(n13401), .Z(c[75]) );
  NAND U18038 ( .A(n13347), .B(o[75]), .Z(n13401) );
  NAND U18039 ( .A(n13342), .B(creg[75]), .Z(n13400) );
  NAND U18040 ( .A(n13402), .B(n13403), .Z(c[74]) );
  NAND U18041 ( .A(n13347), .B(o[74]), .Z(n13403) );
  NAND U18042 ( .A(n13342), .B(creg[74]), .Z(n13402) );
  NAND U18043 ( .A(n13404), .B(n13405), .Z(c[73]) );
  NAND U18044 ( .A(n13347), .B(o[73]), .Z(n13405) );
  NAND U18045 ( .A(n13342), .B(creg[73]), .Z(n13404) );
  NAND U18046 ( .A(n13406), .B(n13407), .Z(c[72]) );
  NAND U18047 ( .A(n13347), .B(o[72]), .Z(n13407) );
  NAND U18048 ( .A(n13342), .B(creg[72]), .Z(n13406) );
  NAND U18049 ( .A(n13408), .B(n13409), .Z(c[71]) );
  NAND U18050 ( .A(n13347), .B(o[71]), .Z(n13409) );
  NAND U18051 ( .A(n13342), .B(creg[71]), .Z(n13408) );
  NAND U18052 ( .A(n13410), .B(n13411), .Z(c[70]) );
  NAND U18053 ( .A(n13347), .B(o[70]), .Z(n13411) );
  NAND U18054 ( .A(n13342), .B(creg[70]), .Z(n13410) );
  NAND U18055 ( .A(n13412), .B(n13413), .Z(c[6]) );
  NAND U18056 ( .A(n13347), .B(o[6]), .Z(n13413) );
  NAND U18057 ( .A(n13342), .B(creg[6]), .Z(n13412) );
  NAND U18058 ( .A(n13414), .B(n13415), .Z(c[69]) );
  NAND U18059 ( .A(n13347), .B(o[69]), .Z(n13415) );
  NAND U18060 ( .A(n13342), .B(creg[69]), .Z(n13414) );
  NAND U18061 ( .A(n13416), .B(n13417), .Z(c[68]) );
  NAND U18062 ( .A(n13347), .B(o[68]), .Z(n13417) );
  NAND U18063 ( .A(n13342), .B(creg[68]), .Z(n13416) );
  NAND U18064 ( .A(n13418), .B(n13419), .Z(c[67]) );
  NAND U18065 ( .A(n13347), .B(o[67]), .Z(n13419) );
  NAND U18066 ( .A(n13342), .B(creg[67]), .Z(n13418) );
  NAND U18067 ( .A(n13420), .B(n13421), .Z(c[66]) );
  NAND U18068 ( .A(n13347), .B(o[66]), .Z(n13421) );
  NAND U18069 ( .A(n13342), .B(creg[66]), .Z(n13420) );
  NAND U18070 ( .A(n13422), .B(n13423), .Z(c[65]) );
  NAND U18071 ( .A(n13347), .B(o[65]), .Z(n13423) );
  NAND U18072 ( .A(n13342), .B(creg[65]), .Z(n13422) );
  NAND U18073 ( .A(n13424), .B(n13425), .Z(c[64]) );
  NAND U18074 ( .A(n13347), .B(o[64]), .Z(n13425) );
  NAND U18075 ( .A(n13342), .B(creg[64]), .Z(n13424) );
  NAND U18076 ( .A(n13426), .B(n13427), .Z(c[63]) );
  NAND U18077 ( .A(n13347), .B(o[63]), .Z(n13427) );
  NAND U18078 ( .A(n13342), .B(creg[63]), .Z(n13426) );
  NAND U18079 ( .A(n13428), .B(n13429), .Z(c[62]) );
  NAND U18080 ( .A(n13347), .B(o[62]), .Z(n13429) );
  NAND U18081 ( .A(n13342), .B(creg[62]), .Z(n13428) );
  NAND U18082 ( .A(n13430), .B(n13431), .Z(c[61]) );
  NAND U18083 ( .A(n13347), .B(o[61]), .Z(n13431) );
  NAND U18084 ( .A(n13342), .B(creg[61]), .Z(n13430) );
  NAND U18085 ( .A(n13432), .B(n13433), .Z(c[60]) );
  NAND U18086 ( .A(n13347), .B(o[60]), .Z(n13433) );
  NAND U18087 ( .A(n13342), .B(creg[60]), .Z(n13432) );
  NAND U18088 ( .A(n13434), .B(n13435), .Z(c[5]) );
  NAND U18089 ( .A(n13347), .B(o[5]), .Z(n13435) );
  NAND U18090 ( .A(n13342), .B(creg[5]), .Z(n13434) );
  NAND U18091 ( .A(n13436), .B(n13437), .Z(c[59]) );
  NAND U18092 ( .A(n13347), .B(o[59]), .Z(n13437) );
  NAND U18093 ( .A(n13342), .B(creg[59]), .Z(n13436) );
  NAND U18094 ( .A(n13438), .B(n13439), .Z(c[58]) );
  NAND U18095 ( .A(n13347), .B(o[58]), .Z(n13439) );
  NAND U18096 ( .A(n13342), .B(creg[58]), .Z(n13438) );
  NAND U18097 ( .A(n13440), .B(n13441), .Z(c[57]) );
  NAND U18098 ( .A(n13347), .B(o[57]), .Z(n13441) );
  NAND U18099 ( .A(n13342), .B(creg[57]), .Z(n13440) );
  NAND U18100 ( .A(n13442), .B(n13443), .Z(c[56]) );
  NAND U18101 ( .A(n13347), .B(o[56]), .Z(n13443) );
  NAND U18102 ( .A(n13342), .B(creg[56]), .Z(n13442) );
  NAND U18103 ( .A(n13444), .B(n13445), .Z(c[55]) );
  NAND U18104 ( .A(n13347), .B(o[55]), .Z(n13445) );
  NAND U18105 ( .A(n13342), .B(creg[55]), .Z(n13444) );
  NAND U18106 ( .A(n13446), .B(n13447), .Z(c[54]) );
  NAND U18107 ( .A(n13347), .B(o[54]), .Z(n13447) );
  NAND U18108 ( .A(n13342), .B(creg[54]), .Z(n13446) );
  NAND U18109 ( .A(n13448), .B(n13449), .Z(c[53]) );
  NAND U18110 ( .A(n13347), .B(o[53]), .Z(n13449) );
  NAND U18111 ( .A(n13342), .B(creg[53]), .Z(n13448) );
  NAND U18112 ( .A(n13450), .B(n13451), .Z(c[52]) );
  NAND U18113 ( .A(n13347), .B(o[52]), .Z(n13451) );
  NAND U18114 ( .A(n13342), .B(creg[52]), .Z(n13450) );
  NAND U18115 ( .A(n13452), .B(n13453), .Z(c[51]) );
  NAND U18116 ( .A(n13347), .B(o[51]), .Z(n13453) );
  NAND U18117 ( .A(n13342), .B(creg[51]), .Z(n13452) );
  NAND U18118 ( .A(n13454), .B(n13455), .Z(c[511]) );
  NAND U18119 ( .A(n13347), .B(o[511]), .Z(n13455) );
  NAND U18120 ( .A(n13342), .B(creg[511]), .Z(n13454) );
  NAND U18121 ( .A(n13456), .B(n13457), .Z(c[510]) );
  NAND U18122 ( .A(n13347), .B(o[510]), .Z(n13457) );
  NAND U18123 ( .A(n13342), .B(creg[510]), .Z(n13456) );
  NAND U18124 ( .A(n13458), .B(n13459), .Z(c[50]) );
  NAND U18125 ( .A(n13347), .B(o[50]), .Z(n13459) );
  NAND U18126 ( .A(n13342), .B(creg[50]), .Z(n13458) );
  NAND U18127 ( .A(n13460), .B(n13461), .Z(c[509]) );
  NAND U18128 ( .A(n13347), .B(o[509]), .Z(n13461) );
  NAND U18129 ( .A(n13342), .B(creg[509]), .Z(n13460) );
  NAND U18130 ( .A(n13462), .B(n13463), .Z(c[508]) );
  NAND U18131 ( .A(n13347), .B(o[508]), .Z(n13463) );
  NAND U18132 ( .A(n13342), .B(creg[508]), .Z(n13462) );
  NAND U18133 ( .A(n13464), .B(n13465), .Z(c[507]) );
  NAND U18134 ( .A(n13347), .B(o[507]), .Z(n13465) );
  NAND U18135 ( .A(n13342), .B(creg[507]), .Z(n13464) );
  NAND U18136 ( .A(n13466), .B(n13467), .Z(c[506]) );
  NAND U18137 ( .A(n13347), .B(o[506]), .Z(n13467) );
  NAND U18138 ( .A(n13342), .B(creg[506]), .Z(n13466) );
  NAND U18139 ( .A(n13468), .B(n13469), .Z(c[505]) );
  NAND U18140 ( .A(n13347), .B(o[505]), .Z(n13469) );
  NAND U18141 ( .A(n13342), .B(creg[505]), .Z(n13468) );
  NAND U18142 ( .A(n13470), .B(n13471), .Z(c[504]) );
  NAND U18143 ( .A(n13347), .B(o[504]), .Z(n13471) );
  NAND U18144 ( .A(n13342), .B(creg[504]), .Z(n13470) );
  NAND U18145 ( .A(n13472), .B(n13473), .Z(c[503]) );
  NAND U18146 ( .A(n13347), .B(o[503]), .Z(n13473) );
  NAND U18147 ( .A(n13342), .B(creg[503]), .Z(n13472) );
  NAND U18148 ( .A(n13474), .B(n13475), .Z(c[502]) );
  NAND U18149 ( .A(n13347), .B(o[502]), .Z(n13475) );
  NAND U18150 ( .A(n13342), .B(creg[502]), .Z(n13474) );
  NAND U18151 ( .A(n13476), .B(n13477), .Z(c[501]) );
  NAND U18152 ( .A(n13347), .B(o[501]), .Z(n13477) );
  NAND U18153 ( .A(n13342), .B(creg[501]), .Z(n13476) );
  NAND U18154 ( .A(n13478), .B(n13479), .Z(c[500]) );
  NAND U18155 ( .A(n13347), .B(o[500]), .Z(n13479) );
  NAND U18156 ( .A(n13342), .B(creg[500]), .Z(n13478) );
  NAND U18157 ( .A(n13480), .B(n13481), .Z(c[4]) );
  NAND U18158 ( .A(n13347), .B(o[4]), .Z(n13481) );
  NAND U18159 ( .A(n13342), .B(creg[4]), .Z(n13480) );
  NAND U18160 ( .A(n13482), .B(n13483), .Z(c[49]) );
  NAND U18161 ( .A(n13347), .B(o[49]), .Z(n13483) );
  NAND U18162 ( .A(n13342), .B(creg[49]), .Z(n13482) );
  NAND U18163 ( .A(n13484), .B(n13485), .Z(c[499]) );
  NAND U18164 ( .A(n13347), .B(o[499]), .Z(n13485) );
  NAND U18165 ( .A(n13342), .B(creg[499]), .Z(n13484) );
  NAND U18166 ( .A(n13486), .B(n13487), .Z(c[498]) );
  NAND U18167 ( .A(n13347), .B(o[498]), .Z(n13487) );
  NAND U18168 ( .A(n13342), .B(creg[498]), .Z(n13486) );
  NAND U18169 ( .A(n13488), .B(n13489), .Z(c[497]) );
  NAND U18170 ( .A(n13347), .B(o[497]), .Z(n13489) );
  NAND U18171 ( .A(n13342), .B(creg[497]), .Z(n13488) );
  NAND U18172 ( .A(n13490), .B(n13491), .Z(c[496]) );
  NAND U18173 ( .A(n13347), .B(o[496]), .Z(n13491) );
  NAND U18174 ( .A(n13342), .B(creg[496]), .Z(n13490) );
  NAND U18175 ( .A(n13492), .B(n13493), .Z(c[495]) );
  NAND U18176 ( .A(n13347), .B(o[495]), .Z(n13493) );
  NAND U18177 ( .A(n13342), .B(creg[495]), .Z(n13492) );
  NAND U18178 ( .A(n13494), .B(n13495), .Z(c[494]) );
  NAND U18179 ( .A(n13347), .B(o[494]), .Z(n13495) );
  NAND U18180 ( .A(n13342), .B(creg[494]), .Z(n13494) );
  NAND U18181 ( .A(n13496), .B(n13497), .Z(c[493]) );
  NAND U18182 ( .A(n13347), .B(o[493]), .Z(n13497) );
  NAND U18183 ( .A(n13342), .B(creg[493]), .Z(n13496) );
  NAND U18184 ( .A(n13498), .B(n13499), .Z(c[492]) );
  NAND U18185 ( .A(n13347), .B(o[492]), .Z(n13499) );
  NAND U18186 ( .A(n13342), .B(creg[492]), .Z(n13498) );
  NAND U18187 ( .A(n13500), .B(n13501), .Z(c[491]) );
  NAND U18188 ( .A(n13347), .B(o[491]), .Z(n13501) );
  NAND U18189 ( .A(n13342), .B(creg[491]), .Z(n13500) );
  NAND U18190 ( .A(n13502), .B(n13503), .Z(c[490]) );
  NAND U18191 ( .A(n13347), .B(o[490]), .Z(n13503) );
  NAND U18192 ( .A(n13342), .B(creg[490]), .Z(n13502) );
  NAND U18193 ( .A(n13504), .B(n13505), .Z(c[48]) );
  NAND U18194 ( .A(n13347), .B(o[48]), .Z(n13505) );
  NAND U18195 ( .A(n13342), .B(creg[48]), .Z(n13504) );
  NAND U18196 ( .A(n13506), .B(n13507), .Z(c[489]) );
  NAND U18197 ( .A(n13347), .B(o[489]), .Z(n13507) );
  NAND U18198 ( .A(n13342), .B(creg[489]), .Z(n13506) );
  NAND U18199 ( .A(n13508), .B(n13509), .Z(c[488]) );
  NAND U18200 ( .A(n13347), .B(o[488]), .Z(n13509) );
  NAND U18201 ( .A(n13342), .B(creg[488]), .Z(n13508) );
  NAND U18202 ( .A(n13510), .B(n13511), .Z(c[487]) );
  NAND U18203 ( .A(n13347), .B(o[487]), .Z(n13511) );
  NAND U18204 ( .A(n13342), .B(creg[487]), .Z(n13510) );
  NAND U18205 ( .A(n13512), .B(n13513), .Z(c[486]) );
  NAND U18206 ( .A(n13347), .B(o[486]), .Z(n13513) );
  NAND U18207 ( .A(n13342), .B(creg[486]), .Z(n13512) );
  NAND U18208 ( .A(n13514), .B(n13515), .Z(c[485]) );
  NAND U18209 ( .A(n13347), .B(o[485]), .Z(n13515) );
  NAND U18210 ( .A(n13342), .B(creg[485]), .Z(n13514) );
  NAND U18211 ( .A(n13516), .B(n13517), .Z(c[484]) );
  NAND U18212 ( .A(n13347), .B(o[484]), .Z(n13517) );
  NAND U18213 ( .A(n13342), .B(creg[484]), .Z(n13516) );
  NAND U18214 ( .A(n13518), .B(n13519), .Z(c[483]) );
  NAND U18215 ( .A(n13347), .B(o[483]), .Z(n13519) );
  NAND U18216 ( .A(n13342), .B(creg[483]), .Z(n13518) );
  NAND U18217 ( .A(n13520), .B(n13521), .Z(c[482]) );
  NAND U18218 ( .A(n13347), .B(o[482]), .Z(n13521) );
  NAND U18219 ( .A(n13342), .B(creg[482]), .Z(n13520) );
  NAND U18220 ( .A(n13522), .B(n13523), .Z(c[481]) );
  NAND U18221 ( .A(n13347), .B(o[481]), .Z(n13523) );
  NAND U18222 ( .A(n13342), .B(creg[481]), .Z(n13522) );
  NAND U18223 ( .A(n13524), .B(n13525), .Z(c[480]) );
  NAND U18224 ( .A(n13347), .B(o[480]), .Z(n13525) );
  NAND U18225 ( .A(n13342), .B(creg[480]), .Z(n13524) );
  NAND U18226 ( .A(n13526), .B(n13527), .Z(c[47]) );
  NAND U18227 ( .A(n13347), .B(o[47]), .Z(n13527) );
  NAND U18228 ( .A(n13342), .B(creg[47]), .Z(n13526) );
  NAND U18229 ( .A(n13528), .B(n13529), .Z(c[479]) );
  NAND U18230 ( .A(n13347), .B(o[479]), .Z(n13529) );
  NAND U18231 ( .A(n13342), .B(creg[479]), .Z(n13528) );
  NAND U18232 ( .A(n13530), .B(n13531), .Z(c[478]) );
  NAND U18233 ( .A(n13347), .B(o[478]), .Z(n13531) );
  NAND U18234 ( .A(n13342), .B(creg[478]), .Z(n13530) );
  NAND U18235 ( .A(n13532), .B(n13533), .Z(c[477]) );
  NAND U18236 ( .A(n13347), .B(o[477]), .Z(n13533) );
  NAND U18237 ( .A(n13342), .B(creg[477]), .Z(n13532) );
  NAND U18238 ( .A(n13534), .B(n13535), .Z(c[476]) );
  NAND U18239 ( .A(n13347), .B(o[476]), .Z(n13535) );
  NAND U18240 ( .A(n13342), .B(creg[476]), .Z(n13534) );
  NAND U18241 ( .A(n13536), .B(n13537), .Z(c[475]) );
  NAND U18242 ( .A(n13347), .B(o[475]), .Z(n13537) );
  NAND U18243 ( .A(n13342), .B(creg[475]), .Z(n13536) );
  NAND U18244 ( .A(n13538), .B(n13539), .Z(c[474]) );
  NAND U18245 ( .A(n13347), .B(o[474]), .Z(n13539) );
  NAND U18246 ( .A(n13342), .B(creg[474]), .Z(n13538) );
  NAND U18247 ( .A(n13540), .B(n13541), .Z(c[473]) );
  NAND U18248 ( .A(n13347), .B(o[473]), .Z(n13541) );
  NAND U18249 ( .A(n13342), .B(creg[473]), .Z(n13540) );
  NAND U18250 ( .A(n13542), .B(n13543), .Z(c[472]) );
  NAND U18251 ( .A(n13347), .B(o[472]), .Z(n13543) );
  NAND U18252 ( .A(n13342), .B(creg[472]), .Z(n13542) );
  NAND U18253 ( .A(n13544), .B(n13545), .Z(c[471]) );
  NAND U18254 ( .A(n13347), .B(o[471]), .Z(n13545) );
  NAND U18255 ( .A(n13342), .B(creg[471]), .Z(n13544) );
  NAND U18256 ( .A(n13546), .B(n13547), .Z(c[470]) );
  NAND U18257 ( .A(n13347), .B(o[470]), .Z(n13547) );
  NAND U18258 ( .A(n13342), .B(creg[470]), .Z(n13546) );
  NAND U18259 ( .A(n13548), .B(n13549), .Z(c[46]) );
  NAND U18260 ( .A(n13347), .B(o[46]), .Z(n13549) );
  NAND U18261 ( .A(n13342), .B(creg[46]), .Z(n13548) );
  NAND U18262 ( .A(n13550), .B(n13551), .Z(c[469]) );
  NAND U18263 ( .A(n13347), .B(o[469]), .Z(n13551) );
  NAND U18264 ( .A(n13342), .B(creg[469]), .Z(n13550) );
  NAND U18265 ( .A(n13552), .B(n13553), .Z(c[468]) );
  NAND U18266 ( .A(n13347), .B(o[468]), .Z(n13553) );
  NAND U18267 ( .A(n13342), .B(creg[468]), .Z(n13552) );
  NAND U18268 ( .A(n13554), .B(n13555), .Z(c[467]) );
  NAND U18269 ( .A(n13347), .B(o[467]), .Z(n13555) );
  NAND U18270 ( .A(n13342), .B(creg[467]), .Z(n13554) );
  NAND U18271 ( .A(n13556), .B(n13557), .Z(c[466]) );
  NAND U18272 ( .A(n13347), .B(o[466]), .Z(n13557) );
  NAND U18273 ( .A(n13342), .B(creg[466]), .Z(n13556) );
  NAND U18274 ( .A(n13558), .B(n13559), .Z(c[465]) );
  NAND U18275 ( .A(n13347), .B(o[465]), .Z(n13559) );
  NAND U18276 ( .A(n13342), .B(creg[465]), .Z(n13558) );
  NAND U18277 ( .A(n13560), .B(n13561), .Z(c[464]) );
  NAND U18278 ( .A(n13347), .B(o[464]), .Z(n13561) );
  NAND U18279 ( .A(n13342), .B(creg[464]), .Z(n13560) );
  NAND U18280 ( .A(n13562), .B(n13563), .Z(c[463]) );
  NAND U18281 ( .A(n13347), .B(o[463]), .Z(n13563) );
  NAND U18282 ( .A(n13342), .B(creg[463]), .Z(n13562) );
  NAND U18283 ( .A(n13564), .B(n13565), .Z(c[462]) );
  NAND U18284 ( .A(n13347), .B(o[462]), .Z(n13565) );
  NAND U18285 ( .A(n13342), .B(creg[462]), .Z(n13564) );
  NAND U18286 ( .A(n13566), .B(n13567), .Z(c[461]) );
  NAND U18287 ( .A(n13347), .B(o[461]), .Z(n13567) );
  NAND U18288 ( .A(n13342), .B(creg[461]), .Z(n13566) );
  NAND U18289 ( .A(n13568), .B(n13569), .Z(c[460]) );
  NAND U18290 ( .A(n13347), .B(o[460]), .Z(n13569) );
  NAND U18291 ( .A(n13342), .B(creg[460]), .Z(n13568) );
  NAND U18292 ( .A(n13570), .B(n13571), .Z(c[45]) );
  NAND U18293 ( .A(n13347), .B(o[45]), .Z(n13571) );
  NAND U18294 ( .A(n13342), .B(creg[45]), .Z(n13570) );
  NAND U18295 ( .A(n13572), .B(n13573), .Z(c[459]) );
  NAND U18296 ( .A(n13347), .B(o[459]), .Z(n13573) );
  NAND U18297 ( .A(n13342), .B(creg[459]), .Z(n13572) );
  NAND U18298 ( .A(n13574), .B(n13575), .Z(c[458]) );
  NAND U18299 ( .A(n13347), .B(o[458]), .Z(n13575) );
  NAND U18300 ( .A(n13342), .B(creg[458]), .Z(n13574) );
  NAND U18301 ( .A(n13576), .B(n13577), .Z(c[457]) );
  NAND U18302 ( .A(n13347), .B(o[457]), .Z(n13577) );
  NAND U18303 ( .A(n13342), .B(creg[457]), .Z(n13576) );
  NAND U18304 ( .A(n13578), .B(n13579), .Z(c[456]) );
  NAND U18305 ( .A(n13347), .B(o[456]), .Z(n13579) );
  NAND U18306 ( .A(n13342), .B(creg[456]), .Z(n13578) );
  NAND U18307 ( .A(n13580), .B(n13581), .Z(c[455]) );
  NAND U18308 ( .A(n13347), .B(o[455]), .Z(n13581) );
  NAND U18309 ( .A(n13342), .B(creg[455]), .Z(n13580) );
  NAND U18310 ( .A(n13582), .B(n13583), .Z(c[454]) );
  NAND U18311 ( .A(n13347), .B(o[454]), .Z(n13583) );
  NAND U18312 ( .A(n13342), .B(creg[454]), .Z(n13582) );
  NAND U18313 ( .A(n13584), .B(n13585), .Z(c[453]) );
  NAND U18314 ( .A(n13347), .B(o[453]), .Z(n13585) );
  NAND U18315 ( .A(n13342), .B(creg[453]), .Z(n13584) );
  NAND U18316 ( .A(n13586), .B(n13587), .Z(c[452]) );
  NAND U18317 ( .A(n13347), .B(o[452]), .Z(n13587) );
  NAND U18318 ( .A(n13342), .B(creg[452]), .Z(n13586) );
  NAND U18319 ( .A(n13588), .B(n13589), .Z(c[451]) );
  NAND U18320 ( .A(n13347), .B(o[451]), .Z(n13589) );
  NAND U18321 ( .A(n13342), .B(creg[451]), .Z(n13588) );
  NAND U18322 ( .A(n13590), .B(n13591), .Z(c[450]) );
  NAND U18323 ( .A(n13347), .B(o[450]), .Z(n13591) );
  NAND U18324 ( .A(n13342), .B(creg[450]), .Z(n13590) );
  NAND U18325 ( .A(n13592), .B(n13593), .Z(c[44]) );
  NAND U18326 ( .A(n13347), .B(o[44]), .Z(n13593) );
  NAND U18327 ( .A(n13342), .B(creg[44]), .Z(n13592) );
  NAND U18328 ( .A(n13594), .B(n13595), .Z(c[449]) );
  NAND U18329 ( .A(n13347), .B(o[449]), .Z(n13595) );
  NAND U18330 ( .A(n13342), .B(creg[449]), .Z(n13594) );
  NAND U18331 ( .A(n13596), .B(n13597), .Z(c[448]) );
  NAND U18332 ( .A(n13347), .B(o[448]), .Z(n13597) );
  NAND U18333 ( .A(n13342), .B(creg[448]), .Z(n13596) );
  NAND U18334 ( .A(n13598), .B(n13599), .Z(c[447]) );
  NAND U18335 ( .A(n13347), .B(o[447]), .Z(n13599) );
  NAND U18336 ( .A(n13342), .B(creg[447]), .Z(n13598) );
  NAND U18337 ( .A(n13600), .B(n13601), .Z(c[446]) );
  NAND U18338 ( .A(n13347), .B(o[446]), .Z(n13601) );
  NAND U18339 ( .A(n13342), .B(creg[446]), .Z(n13600) );
  NAND U18340 ( .A(n13602), .B(n13603), .Z(c[445]) );
  NAND U18341 ( .A(n13347), .B(o[445]), .Z(n13603) );
  NAND U18342 ( .A(n13342), .B(creg[445]), .Z(n13602) );
  NAND U18343 ( .A(n13604), .B(n13605), .Z(c[444]) );
  NAND U18344 ( .A(n13347), .B(o[444]), .Z(n13605) );
  NAND U18345 ( .A(n13342), .B(creg[444]), .Z(n13604) );
  NAND U18346 ( .A(n13606), .B(n13607), .Z(c[443]) );
  NAND U18347 ( .A(n13347), .B(o[443]), .Z(n13607) );
  NAND U18348 ( .A(n13342), .B(creg[443]), .Z(n13606) );
  NAND U18349 ( .A(n13608), .B(n13609), .Z(c[442]) );
  NAND U18350 ( .A(n13347), .B(o[442]), .Z(n13609) );
  NAND U18351 ( .A(n13342), .B(creg[442]), .Z(n13608) );
  NAND U18352 ( .A(n13610), .B(n13611), .Z(c[441]) );
  NAND U18353 ( .A(n13347), .B(o[441]), .Z(n13611) );
  NAND U18354 ( .A(n13342), .B(creg[441]), .Z(n13610) );
  NAND U18355 ( .A(n13612), .B(n13613), .Z(c[440]) );
  NAND U18356 ( .A(n13347), .B(o[440]), .Z(n13613) );
  NAND U18357 ( .A(n13342), .B(creg[440]), .Z(n13612) );
  NAND U18358 ( .A(n13614), .B(n13615), .Z(c[43]) );
  NAND U18359 ( .A(n13347), .B(o[43]), .Z(n13615) );
  NAND U18360 ( .A(n13342), .B(creg[43]), .Z(n13614) );
  NAND U18361 ( .A(n13616), .B(n13617), .Z(c[439]) );
  NAND U18362 ( .A(n13347), .B(o[439]), .Z(n13617) );
  NAND U18363 ( .A(n13342), .B(creg[439]), .Z(n13616) );
  NAND U18364 ( .A(n13618), .B(n13619), .Z(c[438]) );
  NAND U18365 ( .A(n13347), .B(o[438]), .Z(n13619) );
  NAND U18366 ( .A(n13342), .B(creg[438]), .Z(n13618) );
  NAND U18367 ( .A(n13620), .B(n13621), .Z(c[437]) );
  NAND U18368 ( .A(n13347), .B(o[437]), .Z(n13621) );
  NAND U18369 ( .A(n13342), .B(creg[437]), .Z(n13620) );
  NAND U18370 ( .A(n13622), .B(n13623), .Z(c[436]) );
  NAND U18371 ( .A(n13347), .B(o[436]), .Z(n13623) );
  NAND U18372 ( .A(n13342), .B(creg[436]), .Z(n13622) );
  NAND U18373 ( .A(n13624), .B(n13625), .Z(c[435]) );
  NAND U18374 ( .A(n13347), .B(o[435]), .Z(n13625) );
  NAND U18375 ( .A(n13342), .B(creg[435]), .Z(n13624) );
  NAND U18376 ( .A(n13626), .B(n13627), .Z(c[434]) );
  NAND U18377 ( .A(n13347), .B(o[434]), .Z(n13627) );
  NAND U18378 ( .A(n13342), .B(creg[434]), .Z(n13626) );
  NAND U18379 ( .A(n13628), .B(n13629), .Z(c[433]) );
  NAND U18380 ( .A(n13347), .B(o[433]), .Z(n13629) );
  NAND U18381 ( .A(n13342), .B(creg[433]), .Z(n13628) );
  NAND U18382 ( .A(n13630), .B(n13631), .Z(c[432]) );
  NAND U18383 ( .A(n13347), .B(o[432]), .Z(n13631) );
  NAND U18384 ( .A(n13342), .B(creg[432]), .Z(n13630) );
  NAND U18385 ( .A(n13632), .B(n13633), .Z(c[431]) );
  NAND U18386 ( .A(n13347), .B(o[431]), .Z(n13633) );
  NAND U18387 ( .A(n13342), .B(creg[431]), .Z(n13632) );
  NAND U18388 ( .A(n13634), .B(n13635), .Z(c[430]) );
  NAND U18389 ( .A(n13347), .B(o[430]), .Z(n13635) );
  NAND U18390 ( .A(n13342), .B(creg[430]), .Z(n13634) );
  NAND U18391 ( .A(n13636), .B(n13637), .Z(c[42]) );
  NAND U18392 ( .A(n13347), .B(o[42]), .Z(n13637) );
  NAND U18393 ( .A(n13342), .B(creg[42]), .Z(n13636) );
  NAND U18394 ( .A(n13638), .B(n13639), .Z(c[429]) );
  NAND U18395 ( .A(n13347), .B(o[429]), .Z(n13639) );
  NAND U18396 ( .A(n13342), .B(creg[429]), .Z(n13638) );
  NAND U18397 ( .A(n13640), .B(n13641), .Z(c[428]) );
  NAND U18398 ( .A(n13347), .B(o[428]), .Z(n13641) );
  NAND U18399 ( .A(n13342), .B(creg[428]), .Z(n13640) );
  NAND U18400 ( .A(n13642), .B(n13643), .Z(c[427]) );
  NAND U18401 ( .A(n13347), .B(o[427]), .Z(n13643) );
  NAND U18402 ( .A(n13342), .B(creg[427]), .Z(n13642) );
  NAND U18403 ( .A(n13644), .B(n13645), .Z(c[426]) );
  NAND U18404 ( .A(n13347), .B(o[426]), .Z(n13645) );
  NAND U18405 ( .A(n13342), .B(creg[426]), .Z(n13644) );
  NAND U18406 ( .A(n13646), .B(n13647), .Z(c[425]) );
  NAND U18407 ( .A(n13347), .B(o[425]), .Z(n13647) );
  NAND U18408 ( .A(n13342), .B(creg[425]), .Z(n13646) );
  NAND U18409 ( .A(n13648), .B(n13649), .Z(c[424]) );
  NAND U18410 ( .A(n13347), .B(o[424]), .Z(n13649) );
  NAND U18411 ( .A(n13342), .B(creg[424]), .Z(n13648) );
  NAND U18412 ( .A(n13650), .B(n13651), .Z(c[423]) );
  NAND U18413 ( .A(n13347), .B(o[423]), .Z(n13651) );
  NAND U18414 ( .A(n13342), .B(creg[423]), .Z(n13650) );
  NAND U18415 ( .A(n13652), .B(n13653), .Z(c[422]) );
  NAND U18416 ( .A(n13347), .B(o[422]), .Z(n13653) );
  NAND U18417 ( .A(n13342), .B(creg[422]), .Z(n13652) );
  NAND U18418 ( .A(n13654), .B(n13655), .Z(c[421]) );
  NAND U18419 ( .A(n13347), .B(o[421]), .Z(n13655) );
  NAND U18420 ( .A(n13342), .B(creg[421]), .Z(n13654) );
  NAND U18421 ( .A(n13656), .B(n13657), .Z(c[420]) );
  NAND U18422 ( .A(n13347), .B(o[420]), .Z(n13657) );
  NAND U18423 ( .A(n13342), .B(creg[420]), .Z(n13656) );
  NAND U18424 ( .A(n13658), .B(n13659), .Z(c[41]) );
  NAND U18425 ( .A(n13347), .B(o[41]), .Z(n13659) );
  NAND U18426 ( .A(n13342), .B(creg[41]), .Z(n13658) );
  NAND U18427 ( .A(n13660), .B(n13661), .Z(c[419]) );
  NAND U18428 ( .A(n13347), .B(o[419]), .Z(n13661) );
  NAND U18429 ( .A(n13342), .B(creg[419]), .Z(n13660) );
  NAND U18430 ( .A(n13662), .B(n13663), .Z(c[418]) );
  NAND U18431 ( .A(n13347), .B(o[418]), .Z(n13663) );
  NAND U18432 ( .A(n13342), .B(creg[418]), .Z(n13662) );
  NAND U18433 ( .A(n13664), .B(n13665), .Z(c[417]) );
  NAND U18434 ( .A(n13347), .B(o[417]), .Z(n13665) );
  NAND U18435 ( .A(n13342), .B(creg[417]), .Z(n13664) );
  NAND U18436 ( .A(n13666), .B(n13667), .Z(c[416]) );
  NAND U18437 ( .A(n13347), .B(o[416]), .Z(n13667) );
  NAND U18438 ( .A(n13342), .B(creg[416]), .Z(n13666) );
  NAND U18439 ( .A(n13668), .B(n13669), .Z(c[415]) );
  NAND U18440 ( .A(n13347), .B(o[415]), .Z(n13669) );
  NAND U18441 ( .A(n13342), .B(creg[415]), .Z(n13668) );
  NAND U18442 ( .A(n13670), .B(n13671), .Z(c[414]) );
  NAND U18443 ( .A(n13347), .B(o[414]), .Z(n13671) );
  NAND U18444 ( .A(n13342), .B(creg[414]), .Z(n13670) );
  NAND U18445 ( .A(n13672), .B(n13673), .Z(c[413]) );
  NAND U18446 ( .A(n13347), .B(o[413]), .Z(n13673) );
  NAND U18447 ( .A(n13342), .B(creg[413]), .Z(n13672) );
  NAND U18448 ( .A(n13674), .B(n13675), .Z(c[412]) );
  NAND U18449 ( .A(n13347), .B(o[412]), .Z(n13675) );
  NAND U18450 ( .A(n13342), .B(creg[412]), .Z(n13674) );
  NAND U18451 ( .A(n13676), .B(n13677), .Z(c[411]) );
  NAND U18452 ( .A(n13347), .B(o[411]), .Z(n13677) );
  NAND U18453 ( .A(n13342), .B(creg[411]), .Z(n13676) );
  NAND U18454 ( .A(n13678), .B(n13679), .Z(c[410]) );
  NAND U18455 ( .A(n13347), .B(o[410]), .Z(n13679) );
  NAND U18456 ( .A(n13342), .B(creg[410]), .Z(n13678) );
  NAND U18457 ( .A(n13680), .B(n13681), .Z(c[40]) );
  NAND U18458 ( .A(n13347), .B(o[40]), .Z(n13681) );
  NAND U18459 ( .A(n13342), .B(creg[40]), .Z(n13680) );
  NAND U18460 ( .A(n13682), .B(n13683), .Z(c[409]) );
  NAND U18461 ( .A(n13347), .B(o[409]), .Z(n13683) );
  NAND U18462 ( .A(n13342), .B(creg[409]), .Z(n13682) );
  NAND U18463 ( .A(n13684), .B(n13685), .Z(c[408]) );
  NAND U18464 ( .A(n13347), .B(o[408]), .Z(n13685) );
  NAND U18465 ( .A(n13342), .B(creg[408]), .Z(n13684) );
  NAND U18466 ( .A(n13686), .B(n13687), .Z(c[407]) );
  NAND U18467 ( .A(n13347), .B(o[407]), .Z(n13687) );
  NAND U18468 ( .A(n13342), .B(creg[407]), .Z(n13686) );
  NAND U18469 ( .A(n13688), .B(n13689), .Z(c[406]) );
  NAND U18470 ( .A(n13347), .B(o[406]), .Z(n13689) );
  NAND U18471 ( .A(n13342), .B(creg[406]), .Z(n13688) );
  NAND U18472 ( .A(n13690), .B(n13691), .Z(c[405]) );
  NAND U18473 ( .A(n13347), .B(o[405]), .Z(n13691) );
  NAND U18474 ( .A(n13342), .B(creg[405]), .Z(n13690) );
  NAND U18475 ( .A(n13692), .B(n13693), .Z(c[404]) );
  NAND U18476 ( .A(n13347), .B(o[404]), .Z(n13693) );
  NAND U18477 ( .A(n13342), .B(creg[404]), .Z(n13692) );
  NAND U18478 ( .A(n13694), .B(n13695), .Z(c[403]) );
  NAND U18479 ( .A(n13347), .B(o[403]), .Z(n13695) );
  NAND U18480 ( .A(n13342), .B(creg[403]), .Z(n13694) );
  NAND U18481 ( .A(n13696), .B(n13697), .Z(c[402]) );
  NAND U18482 ( .A(n13347), .B(o[402]), .Z(n13697) );
  NAND U18483 ( .A(n13342), .B(creg[402]), .Z(n13696) );
  NAND U18484 ( .A(n13698), .B(n13699), .Z(c[401]) );
  NAND U18485 ( .A(n13347), .B(o[401]), .Z(n13699) );
  NAND U18486 ( .A(n13342), .B(creg[401]), .Z(n13698) );
  NAND U18487 ( .A(n13700), .B(n13701), .Z(c[400]) );
  NAND U18488 ( .A(n13347), .B(o[400]), .Z(n13701) );
  NAND U18489 ( .A(n13342), .B(creg[400]), .Z(n13700) );
  NAND U18490 ( .A(n13702), .B(n13703), .Z(c[3]) );
  NAND U18491 ( .A(n13347), .B(o[3]), .Z(n13703) );
  NAND U18492 ( .A(n13342), .B(creg[3]), .Z(n13702) );
  NAND U18493 ( .A(n13704), .B(n13705), .Z(c[39]) );
  NAND U18494 ( .A(n13347), .B(o[39]), .Z(n13705) );
  NAND U18495 ( .A(n13342), .B(creg[39]), .Z(n13704) );
  NAND U18496 ( .A(n13706), .B(n13707), .Z(c[399]) );
  NAND U18497 ( .A(n13347), .B(o[399]), .Z(n13707) );
  NAND U18498 ( .A(n13342), .B(creg[399]), .Z(n13706) );
  NAND U18499 ( .A(n13708), .B(n13709), .Z(c[398]) );
  NAND U18500 ( .A(n13347), .B(o[398]), .Z(n13709) );
  NAND U18501 ( .A(n13342), .B(creg[398]), .Z(n13708) );
  NAND U18502 ( .A(n13710), .B(n13711), .Z(c[397]) );
  NAND U18503 ( .A(n13347), .B(o[397]), .Z(n13711) );
  NAND U18504 ( .A(n13342), .B(creg[397]), .Z(n13710) );
  NAND U18505 ( .A(n13712), .B(n13713), .Z(c[396]) );
  NAND U18506 ( .A(n13347), .B(o[396]), .Z(n13713) );
  NAND U18507 ( .A(n13342), .B(creg[396]), .Z(n13712) );
  NAND U18508 ( .A(n13714), .B(n13715), .Z(c[395]) );
  NAND U18509 ( .A(n13347), .B(o[395]), .Z(n13715) );
  NAND U18510 ( .A(n13342), .B(creg[395]), .Z(n13714) );
  NAND U18511 ( .A(n13716), .B(n13717), .Z(c[394]) );
  NAND U18512 ( .A(n13347), .B(o[394]), .Z(n13717) );
  NAND U18513 ( .A(n13342), .B(creg[394]), .Z(n13716) );
  NAND U18514 ( .A(n13718), .B(n13719), .Z(c[393]) );
  NAND U18515 ( .A(n13347), .B(o[393]), .Z(n13719) );
  NAND U18516 ( .A(n13342), .B(creg[393]), .Z(n13718) );
  NAND U18517 ( .A(n13720), .B(n13721), .Z(c[392]) );
  NAND U18518 ( .A(n13347), .B(o[392]), .Z(n13721) );
  NAND U18519 ( .A(n13342), .B(creg[392]), .Z(n13720) );
  NAND U18520 ( .A(n13722), .B(n13723), .Z(c[391]) );
  NAND U18521 ( .A(n13347), .B(o[391]), .Z(n13723) );
  NAND U18522 ( .A(n13342), .B(creg[391]), .Z(n13722) );
  NAND U18523 ( .A(n13724), .B(n13725), .Z(c[390]) );
  NAND U18524 ( .A(n13347), .B(o[390]), .Z(n13725) );
  NAND U18525 ( .A(n13342), .B(creg[390]), .Z(n13724) );
  NAND U18526 ( .A(n13726), .B(n13727), .Z(c[38]) );
  NAND U18527 ( .A(n13347), .B(o[38]), .Z(n13727) );
  NAND U18528 ( .A(n13342), .B(creg[38]), .Z(n13726) );
  NAND U18529 ( .A(n13728), .B(n13729), .Z(c[389]) );
  NAND U18530 ( .A(n13347), .B(o[389]), .Z(n13729) );
  NAND U18531 ( .A(n13342), .B(creg[389]), .Z(n13728) );
  NAND U18532 ( .A(n13730), .B(n13731), .Z(c[388]) );
  NAND U18533 ( .A(n13347), .B(o[388]), .Z(n13731) );
  NAND U18534 ( .A(n13342), .B(creg[388]), .Z(n13730) );
  NAND U18535 ( .A(n13732), .B(n13733), .Z(c[387]) );
  NAND U18536 ( .A(n13347), .B(o[387]), .Z(n13733) );
  NAND U18537 ( .A(n13342), .B(creg[387]), .Z(n13732) );
  NAND U18538 ( .A(n13734), .B(n13735), .Z(c[386]) );
  NAND U18539 ( .A(n13347), .B(o[386]), .Z(n13735) );
  NAND U18540 ( .A(n13342), .B(creg[386]), .Z(n13734) );
  NAND U18541 ( .A(n13736), .B(n13737), .Z(c[385]) );
  NAND U18542 ( .A(n13347), .B(o[385]), .Z(n13737) );
  NAND U18543 ( .A(n13342), .B(creg[385]), .Z(n13736) );
  NAND U18544 ( .A(n13738), .B(n13739), .Z(c[384]) );
  NAND U18545 ( .A(n13347), .B(o[384]), .Z(n13739) );
  NAND U18546 ( .A(n13342), .B(creg[384]), .Z(n13738) );
  NAND U18547 ( .A(n13740), .B(n13741), .Z(c[383]) );
  NAND U18548 ( .A(n13347), .B(o[383]), .Z(n13741) );
  NAND U18549 ( .A(n13342), .B(creg[383]), .Z(n13740) );
  NAND U18550 ( .A(n13742), .B(n13743), .Z(c[382]) );
  NAND U18551 ( .A(n13347), .B(o[382]), .Z(n13743) );
  NAND U18552 ( .A(n13342), .B(creg[382]), .Z(n13742) );
  NAND U18553 ( .A(n13744), .B(n13745), .Z(c[381]) );
  NAND U18554 ( .A(n13347), .B(o[381]), .Z(n13745) );
  NAND U18555 ( .A(n13342), .B(creg[381]), .Z(n13744) );
  NAND U18556 ( .A(n13746), .B(n13747), .Z(c[380]) );
  NAND U18557 ( .A(n13347), .B(o[380]), .Z(n13747) );
  NAND U18558 ( .A(n13342), .B(creg[380]), .Z(n13746) );
  NAND U18559 ( .A(n13748), .B(n13749), .Z(c[37]) );
  NAND U18560 ( .A(n13347), .B(o[37]), .Z(n13749) );
  NAND U18561 ( .A(n13342), .B(creg[37]), .Z(n13748) );
  NAND U18562 ( .A(n13750), .B(n13751), .Z(c[379]) );
  NAND U18563 ( .A(n13347), .B(o[379]), .Z(n13751) );
  NAND U18564 ( .A(n13342), .B(creg[379]), .Z(n13750) );
  NAND U18565 ( .A(n13752), .B(n13753), .Z(c[378]) );
  NAND U18566 ( .A(n13347), .B(o[378]), .Z(n13753) );
  NAND U18567 ( .A(n13342), .B(creg[378]), .Z(n13752) );
  NAND U18568 ( .A(n13754), .B(n13755), .Z(c[377]) );
  NAND U18569 ( .A(n13347), .B(o[377]), .Z(n13755) );
  NAND U18570 ( .A(n13342), .B(creg[377]), .Z(n13754) );
  NAND U18571 ( .A(n13756), .B(n13757), .Z(c[376]) );
  NAND U18572 ( .A(n13347), .B(o[376]), .Z(n13757) );
  NAND U18573 ( .A(n13342), .B(creg[376]), .Z(n13756) );
  NAND U18574 ( .A(n13758), .B(n13759), .Z(c[375]) );
  NAND U18575 ( .A(n13347), .B(o[375]), .Z(n13759) );
  NAND U18576 ( .A(n13342), .B(creg[375]), .Z(n13758) );
  NAND U18577 ( .A(n13760), .B(n13761), .Z(c[374]) );
  NAND U18578 ( .A(n13347), .B(o[374]), .Z(n13761) );
  NAND U18579 ( .A(n13342), .B(creg[374]), .Z(n13760) );
  NAND U18580 ( .A(n13762), .B(n13763), .Z(c[373]) );
  NAND U18581 ( .A(n13347), .B(o[373]), .Z(n13763) );
  NAND U18582 ( .A(n13342), .B(creg[373]), .Z(n13762) );
  NAND U18583 ( .A(n13764), .B(n13765), .Z(c[372]) );
  NAND U18584 ( .A(n13347), .B(o[372]), .Z(n13765) );
  NAND U18585 ( .A(n13342), .B(creg[372]), .Z(n13764) );
  NAND U18586 ( .A(n13766), .B(n13767), .Z(c[371]) );
  NAND U18587 ( .A(n13347), .B(o[371]), .Z(n13767) );
  NAND U18588 ( .A(n13342), .B(creg[371]), .Z(n13766) );
  NAND U18589 ( .A(n13768), .B(n13769), .Z(c[370]) );
  NAND U18590 ( .A(n13347), .B(o[370]), .Z(n13769) );
  NAND U18591 ( .A(n13342), .B(creg[370]), .Z(n13768) );
  NAND U18592 ( .A(n13770), .B(n13771), .Z(c[36]) );
  NAND U18593 ( .A(n13347), .B(o[36]), .Z(n13771) );
  NAND U18594 ( .A(n13342), .B(creg[36]), .Z(n13770) );
  NAND U18595 ( .A(n13772), .B(n13773), .Z(c[369]) );
  NAND U18596 ( .A(n13347), .B(o[369]), .Z(n13773) );
  NAND U18597 ( .A(n13342), .B(creg[369]), .Z(n13772) );
  NAND U18598 ( .A(n13774), .B(n13775), .Z(c[368]) );
  NAND U18599 ( .A(n13347), .B(o[368]), .Z(n13775) );
  NAND U18600 ( .A(n13342), .B(creg[368]), .Z(n13774) );
  NAND U18601 ( .A(n13776), .B(n13777), .Z(c[367]) );
  NAND U18602 ( .A(n13347), .B(o[367]), .Z(n13777) );
  NAND U18603 ( .A(n13342), .B(creg[367]), .Z(n13776) );
  NAND U18604 ( .A(n13778), .B(n13779), .Z(c[366]) );
  NAND U18605 ( .A(n13347), .B(o[366]), .Z(n13779) );
  NAND U18606 ( .A(n13342), .B(creg[366]), .Z(n13778) );
  NAND U18607 ( .A(n13780), .B(n13781), .Z(c[365]) );
  NAND U18608 ( .A(n13347), .B(o[365]), .Z(n13781) );
  NAND U18609 ( .A(n13342), .B(creg[365]), .Z(n13780) );
  NAND U18610 ( .A(n13782), .B(n13783), .Z(c[364]) );
  NAND U18611 ( .A(n13347), .B(o[364]), .Z(n13783) );
  NAND U18612 ( .A(n13342), .B(creg[364]), .Z(n13782) );
  NAND U18613 ( .A(n13784), .B(n13785), .Z(c[363]) );
  NAND U18614 ( .A(n13347), .B(o[363]), .Z(n13785) );
  NAND U18615 ( .A(n13342), .B(creg[363]), .Z(n13784) );
  NAND U18616 ( .A(n13786), .B(n13787), .Z(c[362]) );
  NAND U18617 ( .A(n13347), .B(o[362]), .Z(n13787) );
  NAND U18618 ( .A(n13342), .B(creg[362]), .Z(n13786) );
  NAND U18619 ( .A(n13788), .B(n13789), .Z(c[361]) );
  NAND U18620 ( .A(n13347), .B(o[361]), .Z(n13789) );
  NAND U18621 ( .A(n13342), .B(creg[361]), .Z(n13788) );
  NAND U18622 ( .A(n13790), .B(n13791), .Z(c[360]) );
  NAND U18623 ( .A(n13347), .B(o[360]), .Z(n13791) );
  NAND U18624 ( .A(n13342), .B(creg[360]), .Z(n13790) );
  NAND U18625 ( .A(n13792), .B(n13793), .Z(c[35]) );
  NAND U18626 ( .A(n13347), .B(o[35]), .Z(n13793) );
  NAND U18627 ( .A(n13342), .B(creg[35]), .Z(n13792) );
  NAND U18628 ( .A(n13794), .B(n13795), .Z(c[359]) );
  NAND U18629 ( .A(n13347), .B(o[359]), .Z(n13795) );
  NAND U18630 ( .A(n13342), .B(creg[359]), .Z(n13794) );
  NAND U18631 ( .A(n13796), .B(n13797), .Z(c[358]) );
  NAND U18632 ( .A(n13347), .B(o[358]), .Z(n13797) );
  NAND U18633 ( .A(n13342), .B(creg[358]), .Z(n13796) );
  NAND U18634 ( .A(n13798), .B(n13799), .Z(c[357]) );
  NAND U18635 ( .A(n13347), .B(o[357]), .Z(n13799) );
  NAND U18636 ( .A(n13342), .B(creg[357]), .Z(n13798) );
  NAND U18637 ( .A(n13800), .B(n13801), .Z(c[356]) );
  NAND U18638 ( .A(n13347), .B(o[356]), .Z(n13801) );
  NAND U18639 ( .A(n13342), .B(creg[356]), .Z(n13800) );
  NAND U18640 ( .A(n13802), .B(n13803), .Z(c[355]) );
  NAND U18641 ( .A(n13347), .B(o[355]), .Z(n13803) );
  NAND U18642 ( .A(n13342), .B(creg[355]), .Z(n13802) );
  NAND U18643 ( .A(n13804), .B(n13805), .Z(c[354]) );
  NAND U18644 ( .A(n13347), .B(o[354]), .Z(n13805) );
  NAND U18645 ( .A(n13342), .B(creg[354]), .Z(n13804) );
  NAND U18646 ( .A(n13806), .B(n13807), .Z(c[353]) );
  NAND U18647 ( .A(n13347), .B(o[353]), .Z(n13807) );
  NAND U18648 ( .A(n13342), .B(creg[353]), .Z(n13806) );
  NAND U18649 ( .A(n13808), .B(n13809), .Z(c[352]) );
  NAND U18650 ( .A(n13347), .B(o[352]), .Z(n13809) );
  NAND U18651 ( .A(n13342), .B(creg[352]), .Z(n13808) );
  NAND U18652 ( .A(n13810), .B(n13811), .Z(c[351]) );
  NAND U18653 ( .A(n13347), .B(o[351]), .Z(n13811) );
  NAND U18654 ( .A(n13342), .B(creg[351]), .Z(n13810) );
  NAND U18655 ( .A(n13812), .B(n13813), .Z(c[350]) );
  NAND U18656 ( .A(n13347), .B(o[350]), .Z(n13813) );
  NAND U18657 ( .A(n13342), .B(creg[350]), .Z(n13812) );
  NAND U18658 ( .A(n13814), .B(n13815), .Z(c[34]) );
  NAND U18659 ( .A(n13347), .B(o[34]), .Z(n13815) );
  NAND U18660 ( .A(n13342), .B(creg[34]), .Z(n13814) );
  NAND U18661 ( .A(n13816), .B(n13817), .Z(c[349]) );
  NAND U18662 ( .A(n13347), .B(o[349]), .Z(n13817) );
  NAND U18663 ( .A(n13342), .B(creg[349]), .Z(n13816) );
  NAND U18664 ( .A(n13818), .B(n13819), .Z(c[348]) );
  NAND U18665 ( .A(n13347), .B(o[348]), .Z(n13819) );
  NAND U18666 ( .A(n13342), .B(creg[348]), .Z(n13818) );
  NAND U18667 ( .A(n13820), .B(n13821), .Z(c[347]) );
  NAND U18668 ( .A(n13347), .B(o[347]), .Z(n13821) );
  NAND U18669 ( .A(n13342), .B(creg[347]), .Z(n13820) );
  NAND U18670 ( .A(n13822), .B(n13823), .Z(c[346]) );
  NAND U18671 ( .A(n13347), .B(o[346]), .Z(n13823) );
  NAND U18672 ( .A(n13342), .B(creg[346]), .Z(n13822) );
  NAND U18673 ( .A(n13824), .B(n13825), .Z(c[345]) );
  NAND U18674 ( .A(n13347), .B(o[345]), .Z(n13825) );
  NAND U18675 ( .A(n13342), .B(creg[345]), .Z(n13824) );
  NAND U18676 ( .A(n13826), .B(n13827), .Z(c[344]) );
  NAND U18677 ( .A(n13347), .B(o[344]), .Z(n13827) );
  NAND U18678 ( .A(n13342), .B(creg[344]), .Z(n13826) );
  NAND U18679 ( .A(n13828), .B(n13829), .Z(c[343]) );
  NAND U18680 ( .A(n13347), .B(o[343]), .Z(n13829) );
  NAND U18681 ( .A(n13342), .B(creg[343]), .Z(n13828) );
  NAND U18682 ( .A(n13830), .B(n13831), .Z(c[342]) );
  NAND U18683 ( .A(n13347), .B(o[342]), .Z(n13831) );
  NAND U18684 ( .A(n13342), .B(creg[342]), .Z(n13830) );
  NAND U18685 ( .A(n13832), .B(n13833), .Z(c[341]) );
  NAND U18686 ( .A(n13347), .B(o[341]), .Z(n13833) );
  NAND U18687 ( .A(n13342), .B(creg[341]), .Z(n13832) );
  NAND U18688 ( .A(n13834), .B(n13835), .Z(c[340]) );
  NAND U18689 ( .A(n13347), .B(o[340]), .Z(n13835) );
  NAND U18690 ( .A(n13342), .B(creg[340]), .Z(n13834) );
  NAND U18691 ( .A(n13836), .B(n13837), .Z(c[33]) );
  NAND U18692 ( .A(n13347), .B(o[33]), .Z(n13837) );
  NAND U18693 ( .A(n13342), .B(creg[33]), .Z(n13836) );
  NAND U18694 ( .A(n13838), .B(n13839), .Z(c[339]) );
  NAND U18695 ( .A(n13347), .B(o[339]), .Z(n13839) );
  NAND U18696 ( .A(n13342), .B(creg[339]), .Z(n13838) );
  NAND U18697 ( .A(n13840), .B(n13841), .Z(c[338]) );
  NAND U18698 ( .A(n13347), .B(o[338]), .Z(n13841) );
  NAND U18699 ( .A(n13342), .B(creg[338]), .Z(n13840) );
  NAND U18700 ( .A(n13842), .B(n13843), .Z(c[337]) );
  NAND U18701 ( .A(n13347), .B(o[337]), .Z(n13843) );
  NAND U18702 ( .A(n13342), .B(creg[337]), .Z(n13842) );
  NAND U18703 ( .A(n13844), .B(n13845), .Z(c[336]) );
  NAND U18704 ( .A(n13347), .B(o[336]), .Z(n13845) );
  NAND U18705 ( .A(n13342), .B(creg[336]), .Z(n13844) );
  NAND U18706 ( .A(n13846), .B(n13847), .Z(c[335]) );
  NAND U18707 ( .A(n13347), .B(o[335]), .Z(n13847) );
  NAND U18708 ( .A(n13342), .B(creg[335]), .Z(n13846) );
  NAND U18709 ( .A(n13848), .B(n13849), .Z(c[334]) );
  NAND U18710 ( .A(n13347), .B(o[334]), .Z(n13849) );
  NAND U18711 ( .A(n13342), .B(creg[334]), .Z(n13848) );
  NAND U18712 ( .A(n13850), .B(n13851), .Z(c[333]) );
  NAND U18713 ( .A(n13347), .B(o[333]), .Z(n13851) );
  NAND U18714 ( .A(n13342), .B(creg[333]), .Z(n13850) );
  NAND U18715 ( .A(n13852), .B(n13853), .Z(c[332]) );
  NAND U18716 ( .A(n13347), .B(o[332]), .Z(n13853) );
  NAND U18717 ( .A(n13342), .B(creg[332]), .Z(n13852) );
  NAND U18718 ( .A(n13854), .B(n13855), .Z(c[331]) );
  NAND U18719 ( .A(n13347), .B(o[331]), .Z(n13855) );
  NAND U18720 ( .A(n13342), .B(creg[331]), .Z(n13854) );
  NAND U18721 ( .A(n13856), .B(n13857), .Z(c[330]) );
  NAND U18722 ( .A(n13347), .B(o[330]), .Z(n13857) );
  NAND U18723 ( .A(n13342), .B(creg[330]), .Z(n13856) );
  NAND U18724 ( .A(n13858), .B(n13859), .Z(c[32]) );
  NAND U18725 ( .A(n13347), .B(o[32]), .Z(n13859) );
  NAND U18726 ( .A(n13342), .B(creg[32]), .Z(n13858) );
  NAND U18727 ( .A(n13860), .B(n13861), .Z(c[329]) );
  NAND U18728 ( .A(n13347), .B(o[329]), .Z(n13861) );
  NAND U18729 ( .A(n13342), .B(creg[329]), .Z(n13860) );
  NAND U18730 ( .A(n13862), .B(n13863), .Z(c[328]) );
  NAND U18731 ( .A(n13347), .B(o[328]), .Z(n13863) );
  NAND U18732 ( .A(n13342), .B(creg[328]), .Z(n13862) );
  NAND U18733 ( .A(n13864), .B(n13865), .Z(c[327]) );
  NAND U18734 ( .A(n13347), .B(o[327]), .Z(n13865) );
  NAND U18735 ( .A(n13342), .B(creg[327]), .Z(n13864) );
  NAND U18736 ( .A(n13866), .B(n13867), .Z(c[326]) );
  NAND U18737 ( .A(n13347), .B(o[326]), .Z(n13867) );
  NAND U18738 ( .A(n13342), .B(creg[326]), .Z(n13866) );
  NAND U18739 ( .A(n13868), .B(n13869), .Z(c[325]) );
  NAND U18740 ( .A(n13347), .B(o[325]), .Z(n13869) );
  NAND U18741 ( .A(n13342), .B(creg[325]), .Z(n13868) );
  NAND U18742 ( .A(n13870), .B(n13871), .Z(c[324]) );
  NAND U18743 ( .A(n13347), .B(o[324]), .Z(n13871) );
  NAND U18744 ( .A(n13342), .B(creg[324]), .Z(n13870) );
  NAND U18745 ( .A(n13872), .B(n13873), .Z(c[323]) );
  NAND U18746 ( .A(n13347), .B(o[323]), .Z(n13873) );
  NAND U18747 ( .A(n13342), .B(creg[323]), .Z(n13872) );
  NAND U18748 ( .A(n13874), .B(n13875), .Z(c[322]) );
  NAND U18749 ( .A(n13347), .B(o[322]), .Z(n13875) );
  NAND U18750 ( .A(n13342), .B(creg[322]), .Z(n13874) );
  NAND U18751 ( .A(n13876), .B(n13877), .Z(c[321]) );
  NAND U18752 ( .A(n13347), .B(o[321]), .Z(n13877) );
  NAND U18753 ( .A(n13342), .B(creg[321]), .Z(n13876) );
  NAND U18754 ( .A(n13878), .B(n13879), .Z(c[320]) );
  NAND U18755 ( .A(n13347), .B(o[320]), .Z(n13879) );
  NAND U18756 ( .A(n13342), .B(creg[320]), .Z(n13878) );
  NAND U18757 ( .A(n13880), .B(n13881), .Z(c[31]) );
  NAND U18758 ( .A(n13347), .B(o[31]), .Z(n13881) );
  NAND U18759 ( .A(n13342), .B(creg[31]), .Z(n13880) );
  NAND U18760 ( .A(n13882), .B(n13883), .Z(c[319]) );
  NAND U18761 ( .A(n13347), .B(o[319]), .Z(n13883) );
  NAND U18762 ( .A(n13342), .B(creg[319]), .Z(n13882) );
  NAND U18763 ( .A(n13884), .B(n13885), .Z(c[318]) );
  NAND U18764 ( .A(n13347), .B(o[318]), .Z(n13885) );
  NAND U18765 ( .A(n13342), .B(creg[318]), .Z(n13884) );
  NAND U18766 ( .A(n13886), .B(n13887), .Z(c[317]) );
  NAND U18767 ( .A(n13347), .B(o[317]), .Z(n13887) );
  NAND U18768 ( .A(n13342), .B(creg[317]), .Z(n13886) );
  NAND U18769 ( .A(n13888), .B(n13889), .Z(c[316]) );
  NAND U18770 ( .A(n13347), .B(o[316]), .Z(n13889) );
  NAND U18771 ( .A(n13342), .B(creg[316]), .Z(n13888) );
  NAND U18772 ( .A(n13890), .B(n13891), .Z(c[315]) );
  NAND U18773 ( .A(n13347), .B(o[315]), .Z(n13891) );
  NAND U18774 ( .A(n13342), .B(creg[315]), .Z(n13890) );
  NAND U18775 ( .A(n13892), .B(n13893), .Z(c[314]) );
  NAND U18776 ( .A(n13347), .B(o[314]), .Z(n13893) );
  NAND U18777 ( .A(n13342), .B(creg[314]), .Z(n13892) );
  NAND U18778 ( .A(n13894), .B(n13895), .Z(c[313]) );
  NAND U18779 ( .A(n13347), .B(o[313]), .Z(n13895) );
  NAND U18780 ( .A(n13342), .B(creg[313]), .Z(n13894) );
  NAND U18781 ( .A(n13896), .B(n13897), .Z(c[312]) );
  NAND U18782 ( .A(n13347), .B(o[312]), .Z(n13897) );
  NAND U18783 ( .A(n13342), .B(creg[312]), .Z(n13896) );
  NAND U18784 ( .A(n13898), .B(n13899), .Z(c[311]) );
  NAND U18785 ( .A(n13347), .B(o[311]), .Z(n13899) );
  NAND U18786 ( .A(n13342), .B(creg[311]), .Z(n13898) );
  NAND U18787 ( .A(n13900), .B(n13901), .Z(c[310]) );
  NAND U18788 ( .A(n13347), .B(o[310]), .Z(n13901) );
  NAND U18789 ( .A(n13342), .B(creg[310]), .Z(n13900) );
  NAND U18790 ( .A(n13902), .B(n13903), .Z(c[30]) );
  NAND U18791 ( .A(n13347), .B(o[30]), .Z(n13903) );
  NAND U18792 ( .A(n13342), .B(creg[30]), .Z(n13902) );
  NAND U18793 ( .A(n13904), .B(n13905), .Z(c[309]) );
  NAND U18794 ( .A(n13347), .B(o[309]), .Z(n13905) );
  NAND U18795 ( .A(n13342), .B(creg[309]), .Z(n13904) );
  NAND U18796 ( .A(n13906), .B(n13907), .Z(c[308]) );
  NAND U18797 ( .A(n13347), .B(o[308]), .Z(n13907) );
  NAND U18798 ( .A(n13342), .B(creg[308]), .Z(n13906) );
  NAND U18799 ( .A(n13908), .B(n13909), .Z(c[307]) );
  NAND U18800 ( .A(n13347), .B(o[307]), .Z(n13909) );
  NAND U18801 ( .A(n13342), .B(creg[307]), .Z(n13908) );
  NAND U18802 ( .A(n13910), .B(n13911), .Z(c[306]) );
  NAND U18803 ( .A(n13347), .B(o[306]), .Z(n13911) );
  NAND U18804 ( .A(n13342), .B(creg[306]), .Z(n13910) );
  NAND U18805 ( .A(n13912), .B(n13913), .Z(c[305]) );
  NAND U18806 ( .A(n13347), .B(o[305]), .Z(n13913) );
  NAND U18807 ( .A(n13342), .B(creg[305]), .Z(n13912) );
  NAND U18808 ( .A(n13914), .B(n13915), .Z(c[304]) );
  NAND U18809 ( .A(n13347), .B(o[304]), .Z(n13915) );
  NAND U18810 ( .A(n13342), .B(creg[304]), .Z(n13914) );
  NAND U18811 ( .A(n13916), .B(n13917), .Z(c[303]) );
  NAND U18812 ( .A(n13347), .B(o[303]), .Z(n13917) );
  NAND U18813 ( .A(n13342), .B(creg[303]), .Z(n13916) );
  NAND U18814 ( .A(n13918), .B(n13919), .Z(c[302]) );
  NAND U18815 ( .A(n13347), .B(o[302]), .Z(n13919) );
  NAND U18816 ( .A(n13342), .B(creg[302]), .Z(n13918) );
  NAND U18817 ( .A(n13920), .B(n13921), .Z(c[301]) );
  NAND U18818 ( .A(n13347), .B(o[301]), .Z(n13921) );
  NAND U18819 ( .A(n13342), .B(creg[301]), .Z(n13920) );
  NAND U18820 ( .A(n13922), .B(n13923), .Z(c[300]) );
  NAND U18821 ( .A(n13347), .B(o[300]), .Z(n13923) );
  NAND U18822 ( .A(n13342), .B(creg[300]), .Z(n13922) );
  NAND U18823 ( .A(n13924), .B(n13925), .Z(c[2]) );
  NAND U18824 ( .A(n13347), .B(o[2]), .Z(n13925) );
  NAND U18825 ( .A(n13342), .B(creg[2]), .Z(n13924) );
  NAND U18826 ( .A(n13926), .B(n13927), .Z(c[29]) );
  NAND U18827 ( .A(n13347), .B(o[29]), .Z(n13927) );
  NAND U18828 ( .A(n13342), .B(creg[29]), .Z(n13926) );
  NAND U18829 ( .A(n13928), .B(n13929), .Z(c[299]) );
  NAND U18830 ( .A(n13347), .B(o[299]), .Z(n13929) );
  NAND U18831 ( .A(n13342), .B(creg[299]), .Z(n13928) );
  NAND U18832 ( .A(n13930), .B(n13931), .Z(c[298]) );
  NAND U18833 ( .A(n13347), .B(o[298]), .Z(n13931) );
  NAND U18834 ( .A(n13342), .B(creg[298]), .Z(n13930) );
  NAND U18835 ( .A(n13932), .B(n13933), .Z(c[297]) );
  NAND U18836 ( .A(n13347), .B(o[297]), .Z(n13933) );
  NAND U18837 ( .A(n13342), .B(creg[297]), .Z(n13932) );
  NAND U18838 ( .A(n13934), .B(n13935), .Z(c[296]) );
  NAND U18839 ( .A(n13347), .B(o[296]), .Z(n13935) );
  NAND U18840 ( .A(n13342), .B(creg[296]), .Z(n13934) );
  NAND U18841 ( .A(n13936), .B(n13937), .Z(c[295]) );
  NAND U18842 ( .A(n13347), .B(o[295]), .Z(n13937) );
  NAND U18843 ( .A(n13342), .B(creg[295]), .Z(n13936) );
  NAND U18844 ( .A(n13938), .B(n13939), .Z(c[294]) );
  NAND U18845 ( .A(n13347), .B(o[294]), .Z(n13939) );
  NAND U18846 ( .A(n13342), .B(creg[294]), .Z(n13938) );
  NAND U18847 ( .A(n13940), .B(n13941), .Z(c[293]) );
  NAND U18848 ( .A(n13347), .B(o[293]), .Z(n13941) );
  NAND U18849 ( .A(n13342), .B(creg[293]), .Z(n13940) );
  NAND U18850 ( .A(n13942), .B(n13943), .Z(c[292]) );
  NAND U18851 ( .A(n13347), .B(o[292]), .Z(n13943) );
  NAND U18852 ( .A(n13342), .B(creg[292]), .Z(n13942) );
  NAND U18853 ( .A(n13944), .B(n13945), .Z(c[291]) );
  NAND U18854 ( .A(n13347), .B(o[291]), .Z(n13945) );
  NAND U18855 ( .A(n13342), .B(creg[291]), .Z(n13944) );
  NAND U18856 ( .A(n13946), .B(n13947), .Z(c[290]) );
  NAND U18857 ( .A(n13347), .B(o[290]), .Z(n13947) );
  NAND U18858 ( .A(n13342), .B(creg[290]), .Z(n13946) );
  NAND U18859 ( .A(n13948), .B(n13949), .Z(c[28]) );
  NAND U18860 ( .A(n13347), .B(o[28]), .Z(n13949) );
  NAND U18861 ( .A(n13342), .B(creg[28]), .Z(n13948) );
  NAND U18862 ( .A(n13950), .B(n13951), .Z(c[289]) );
  NAND U18863 ( .A(n13347), .B(o[289]), .Z(n13951) );
  NAND U18864 ( .A(n13342), .B(creg[289]), .Z(n13950) );
  NAND U18865 ( .A(n13952), .B(n13953), .Z(c[288]) );
  NAND U18866 ( .A(n13347), .B(o[288]), .Z(n13953) );
  NAND U18867 ( .A(n13342), .B(creg[288]), .Z(n13952) );
  NAND U18868 ( .A(n13954), .B(n13955), .Z(c[287]) );
  NAND U18869 ( .A(n13347), .B(o[287]), .Z(n13955) );
  NAND U18870 ( .A(n13342), .B(creg[287]), .Z(n13954) );
  NAND U18871 ( .A(n13956), .B(n13957), .Z(c[286]) );
  NAND U18872 ( .A(n13347), .B(o[286]), .Z(n13957) );
  NAND U18873 ( .A(n13342), .B(creg[286]), .Z(n13956) );
  NAND U18874 ( .A(n13958), .B(n13959), .Z(c[285]) );
  NAND U18875 ( .A(n13347), .B(o[285]), .Z(n13959) );
  NAND U18876 ( .A(n13342), .B(creg[285]), .Z(n13958) );
  NAND U18877 ( .A(n13960), .B(n13961), .Z(c[284]) );
  NAND U18878 ( .A(n13347), .B(o[284]), .Z(n13961) );
  NAND U18879 ( .A(n13342), .B(creg[284]), .Z(n13960) );
  NAND U18880 ( .A(n13962), .B(n13963), .Z(c[283]) );
  NAND U18881 ( .A(n13347), .B(o[283]), .Z(n13963) );
  NAND U18882 ( .A(n13342), .B(creg[283]), .Z(n13962) );
  NAND U18883 ( .A(n13964), .B(n13965), .Z(c[282]) );
  NAND U18884 ( .A(n13347), .B(o[282]), .Z(n13965) );
  NAND U18885 ( .A(n13342), .B(creg[282]), .Z(n13964) );
  NAND U18886 ( .A(n13966), .B(n13967), .Z(c[281]) );
  NAND U18887 ( .A(n13347), .B(o[281]), .Z(n13967) );
  NAND U18888 ( .A(n13342), .B(creg[281]), .Z(n13966) );
  NAND U18889 ( .A(n13968), .B(n13969), .Z(c[280]) );
  NAND U18890 ( .A(n13347), .B(o[280]), .Z(n13969) );
  NAND U18891 ( .A(n13342), .B(creg[280]), .Z(n13968) );
  NAND U18892 ( .A(n13970), .B(n13971), .Z(c[27]) );
  NAND U18893 ( .A(n13347), .B(o[27]), .Z(n13971) );
  NAND U18894 ( .A(n13342), .B(creg[27]), .Z(n13970) );
  NAND U18895 ( .A(n13972), .B(n13973), .Z(c[279]) );
  NAND U18896 ( .A(n13347), .B(o[279]), .Z(n13973) );
  NAND U18897 ( .A(n13342), .B(creg[279]), .Z(n13972) );
  NAND U18898 ( .A(n13974), .B(n13975), .Z(c[278]) );
  NAND U18899 ( .A(n13347), .B(o[278]), .Z(n13975) );
  NAND U18900 ( .A(n13342), .B(creg[278]), .Z(n13974) );
  NAND U18901 ( .A(n13976), .B(n13977), .Z(c[277]) );
  NAND U18902 ( .A(n13347), .B(o[277]), .Z(n13977) );
  NAND U18903 ( .A(n13342), .B(creg[277]), .Z(n13976) );
  NAND U18904 ( .A(n13978), .B(n13979), .Z(c[276]) );
  NAND U18905 ( .A(n13347), .B(o[276]), .Z(n13979) );
  NAND U18906 ( .A(n13342), .B(creg[276]), .Z(n13978) );
  NAND U18907 ( .A(n13980), .B(n13981), .Z(c[275]) );
  NAND U18908 ( .A(n13347), .B(o[275]), .Z(n13981) );
  NAND U18909 ( .A(n13342), .B(creg[275]), .Z(n13980) );
  NAND U18910 ( .A(n13982), .B(n13983), .Z(c[274]) );
  NAND U18911 ( .A(n13347), .B(o[274]), .Z(n13983) );
  NAND U18912 ( .A(n13342), .B(creg[274]), .Z(n13982) );
  NAND U18913 ( .A(n13984), .B(n13985), .Z(c[273]) );
  NAND U18914 ( .A(n13347), .B(o[273]), .Z(n13985) );
  NAND U18915 ( .A(n13342), .B(creg[273]), .Z(n13984) );
  NAND U18916 ( .A(n13986), .B(n13987), .Z(c[272]) );
  NAND U18917 ( .A(n13347), .B(o[272]), .Z(n13987) );
  NAND U18918 ( .A(n13342), .B(creg[272]), .Z(n13986) );
  NAND U18919 ( .A(n13988), .B(n13989), .Z(c[271]) );
  NAND U18920 ( .A(n13347), .B(o[271]), .Z(n13989) );
  NAND U18921 ( .A(n13342), .B(creg[271]), .Z(n13988) );
  NAND U18922 ( .A(n13990), .B(n13991), .Z(c[270]) );
  NAND U18923 ( .A(n13347), .B(o[270]), .Z(n13991) );
  NAND U18924 ( .A(n13342), .B(creg[270]), .Z(n13990) );
  NAND U18925 ( .A(n13992), .B(n13993), .Z(c[26]) );
  NAND U18926 ( .A(n13347), .B(o[26]), .Z(n13993) );
  NAND U18927 ( .A(n13342), .B(creg[26]), .Z(n13992) );
  NAND U18928 ( .A(n13994), .B(n13995), .Z(c[269]) );
  NAND U18929 ( .A(n13347), .B(o[269]), .Z(n13995) );
  NAND U18930 ( .A(n13342), .B(creg[269]), .Z(n13994) );
  NAND U18931 ( .A(n13996), .B(n13997), .Z(c[268]) );
  NAND U18932 ( .A(n13347), .B(o[268]), .Z(n13997) );
  NAND U18933 ( .A(n13342), .B(creg[268]), .Z(n13996) );
  NAND U18934 ( .A(n13998), .B(n13999), .Z(c[267]) );
  NAND U18935 ( .A(n13347), .B(o[267]), .Z(n13999) );
  NAND U18936 ( .A(n13342), .B(creg[267]), .Z(n13998) );
  NAND U18937 ( .A(n14000), .B(n14001), .Z(c[266]) );
  NAND U18938 ( .A(n13347), .B(o[266]), .Z(n14001) );
  NAND U18939 ( .A(n13342), .B(creg[266]), .Z(n14000) );
  NAND U18940 ( .A(n14002), .B(n14003), .Z(c[265]) );
  NAND U18941 ( .A(n13347), .B(o[265]), .Z(n14003) );
  NAND U18942 ( .A(n13342), .B(creg[265]), .Z(n14002) );
  NAND U18943 ( .A(n14004), .B(n14005), .Z(c[264]) );
  NAND U18944 ( .A(n13347), .B(o[264]), .Z(n14005) );
  NAND U18945 ( .A(n13342), .B(creg[264]), .Z(n14004) );
  NAND U18946 ( .A(n14006), .B(n14007), .Z(c[263]) );
  NAND U18947 ( .A(n13347), .B(o[263]), .Z(n14007) );
  NAND U18948 ( .A(n13342), .B(creg[263]), .Z(n14006) );
  NAND U18949 ( .A(n14008), .B(n14009), .Z(c[262]) );
  NAND U18950 ( .A(n13347), .B(o[262]), .Z(n14009) );
  NAND U18951 ( .A(n13342), .B(creg[262]), .Z(n14008) );
  NAND U18952 ( .A(n14010), .B(n14011), .Z(c[261]) );
  NAND U18953 ( .A(n13347), .B(o[261]), .Z(n14011) );
  NAND U18954 ( .A(n13342), .B(creg[261]), .Z(n14010) );
  NAND U18955 ( .A(n14012), .B(n14013), .Z(c[260]) );
  NAND U18956 ( .A(n13347), .B(o[260]), .Z(n14013) );
  NAND U18957 ( .A(n13342), .B(creg[260]), .Z(n14012) );
  NAND U18958 ( .A(n14014), .B(n14015), .Z(c[25]) );
  NAND U18959 ( .A(n13347), .B(o[25]), .Z(n14015) );
  NAND U18960 ( .A(n13342), .B(creg[25]), .Z(n14014) );
  NAND U18961 ( .A(n14016), .B(n14017), .Z(c[259]) );
  NAND U18962 ( .A(n13347), .B(o[259]), .Z(n14017) );
  NAND U18963 ( .A(n13342), .B(creg[259]), .Z(n14016) );
  NAND U18964 ( .A(n14018), .B(n14019), .Z(c[258]) );
  NAND U18965 ( .A(n13347), .B(o[258]), .Z(n14019) );
  NAND U18966 ( .A(n13342), .B(creg[258]), .Z(n14018) );
  NAND U18967 ( .A(n14020), .B(n14021), .Z(c[257]) );
  NAND U18968 ( .A(n13347), .B(o[257]), .Z(n14021) );
  NAND U18969 ( .A(n13342), .B(creg[257]), .Z(n14020) );
  NAND U18970 ( .A(n14022), .B(n14023), .Z(c[256]) );
  NAND U18971 ( .A(n13347), .B(o[256]), .Z(n14023) );
  NAND U18972 ( .A(n13342), .B(creg[256]), .Z(n14022) );
  NAND U18973 ( .A(n14024), .B(n14025), .Z(c[255]) );
  NAND U18974 ( .A(n13347), .B(o[255]), .Z(n14025) );
  NAND U18975 ( .A(n13342), .B(creg[255]), .Z(n14024) );
  NAND U18976 ( .A(n14026), .B(n14027), .Z(c[254]) );
  NAND U18977 ( .A(n13347), .B(o[254]), .Z(n14027) );
  NAND U18978 ( .A(n13342), .B(creg[254]), .Z(n14026) );
  NAND U18979 ( .A(n14028), .B(n14029), .Z(c[253]) );
  NAND U18980 ( .A(n13347), .B(o[253]), .Z(n14029) );
  NAND U18981 ( .A(n13342), .B(creg[253]), .Z(n14028) );
  NAND U18982 ( .A(n14030), .B(n14031), .Z(c[252]) );
  NAND U18983 ( .A(n13347), .B(o[252]), .Z(n14031) );
  NAND U18984 ( .A(n13342), .B(creg[252]), .Z(n14030) );
  NAND U18985 ( .A(n14032), .B(n14033), .Z(c[251]) );
  NAND U18986 ( .A(n13347), .B(o[251]), .Z(n14033) );
  NAND U18987 ( .A(n13342), .B(creg[251]), .Z(n14032) );
  NAND U18988 ( .A(n14034), .B(n14035), .Z(c[250]) );
  NAND U18989 ( .A(n13347), .B(o[250]), .Z(n14035) );
  NAND U18990 ( .A(n13342), .B(creg[250]), .Z(n14034) );
  NAND U18991 ( .A(n14036), .B(n14037), .Z(c[24]) );
  NAND U18992 ( .A(n13347), .B(o[24]), .Z(n14037) );
  NAND U18993 ( .A(n13342), .B(creg[24]), .Z(n14036) );
  NAND U18994 ( .A(n14038), .B(n14039), .Z(c[249]) );
  NAND U18995 ( .A(n13347), .B(o[249]), .Z(n14039) );
  NAND U18996 ( .A(n13342), .B(creg[249]), .Z(n14038) );
  NAND U18997 ( .A(n14040), .B(n14041), .Z(c[248]) );
  NAND U18998 ( .A(n13347), .B(o[248]), .Z(n14041) );
  NAND U18999 ( .A(n13342), .B(creg[248]), .Z(n14040) );
  NAND U19000 ( .A(n14042), .B(n14043), .Z(c[247]) );
  NAND U19001 ( .A(n13347), .B(o[247]), .Z(n14043) );
  NAND U19002 ( .A(n13342), .B(creg[247]), .Z(n14042) );
  NAND U19003 ( .A(n14044), .B(n14045), .Z(c[246]) );
  NAND U19004 ( .A(n13347), .B(o[246]), .Z(n14045) );
  NAND U19005 ( .A(n13342), .B(creg[246]), .Z(n14044) );
  NAND U19006 ( .A(n14046), .B(n14047), .Z(c[245]) );
  NAND U19007 ( .A(n13347), .B(o[245]), .Z(n14047) );
  NAND U19008 ( .A(n13342), .B(creg[245]), .Z(n14046) );
  NAND U19009 ( .A(n14048), .B(n14049), .Z(c[244]) );
  NAND U19010 ( .A(n13347), .B(o[244]), .Z(n14049) );
  NAND U19011 ( .A(n13342), .B(creg[244]), .Z(n14048) );
  NAND U19012 ( .A(n14050), .B(n14051), .Z(c[243]) );
  NAND U19013 ( .A(n13347), .B(o[243]), .Z(n14051) );
  NAND U19014 ( .A(n13342), .B(creg[243]), .Z(n14050) );
  NAND U19015 ( .A(n14052), .B(n14053), .Z(c[242]) );
  NAND U19016 ( .A(n13347), .B(o[242]), .Z(n14053) );
  NAND U19017 ( .A(n13342), .B(creg[242]), .Z(n14052) );
  NAND U19018 ( .A(n14054), .B(n14055), .Z(c[241]) );
  NAND U19019 ( .A(n13347), .B(o[241]), .Z(n14055) );
  NAND U19020 ( .A(n13342), .B(creg[241]), .Z(n14054) );
  NAND U19021 ( .A(n14056), .B(n14057), .Z(c[240]) );
  NAND U19022 ( .A(n13347), .B(o[240]), .Z(n14057) );
  NAND U19023 ( .A(n13342), .B(creg[240]), .Z(n14056) );
  NAND U19024 ( .A(n14058), .B(n14059), .Z(c[23]) );
  NAND U19025 ( .A(n13347), .B(o[23]), .Z(n14059) );
  NAND U19026 ( .A(n13342), .B(creg[23]), .Z(n14058) );
  NAND U19027 ( .A(n14060), .B(n14061), .Z(c[239]) );
  NAND U19028 ( .A(n13347), .B(o[239]), .Z(n14061) );
  NAND U19029 ( .A(n13342), .B(creg[239]), .Z(n14060) );
  NAND U19030 ( .A(n14062), .B(n14063), .Z(c[238]) );
  NAND U19031 ( .A(n13347), .B(o[238]), .Z(n14063) );
  NAND U19032 ( .A(n13342), .B(creg[238]), .Z(n14062) );
  NAND U19033 ( .A(n14064), .B(n14065), .Z(c[237]) );
  NAND U19034 ( .A(n13347), .B(o[237]), .Z(n14065) );
  NAND U19035 ( .A(n13342), .B(creg[237]), .Z(n14064) );
  NAND U19036 ( .A(n14066), .B(n14067), .Z(c[236]) );
  NAND U19037 ( .A(n13347), .B(o[236]), .Z(n14067) );
  NAND U19038 ( .A(n13342), .B(creg[236]), .Z(n14066) );
  NAND U19039 ( .A(n14068), .B(n14069), .Z(c[235]) );
  NAND U19040 ( .A(n13347), .B(o[235]), .Z(n14069) );
  NAND U19041 ( .A(n13342), .B(creg[235]), .Z(n14068) );
  NAND U19042 ( .A(n14070), .B(n14071), .Z(c[234]) );
  NAND U19043 ( .A(n13347), .B(o[234]), .Z(n14071) );
  NAND U19044 ( .A(n13342), .B(creg[234]), .Z(n14070) );
  NAND U19045 ( .A(n14072), .B(n14073), .Z(c[233]) );
  NAND U19046 ( .A(n13347), .B(o[233]), .Z(n14073) );
  NAND U19047 ( .A(n13342), .B(creg[233]), .Z(n14072) );
  NAND U19048 ( .A(n14074), .B(n14075), .Z(c[232]) );
  NAND U19049 ( .A(n13347), .B(o[232]), .Z(n14075) );
  NAND U19050 ( .A(n13342), .B(creg[232]), .Z(n14074) );
  NAND U19051 ( .A(n14076), .B(n14077), .Z(c[231]) );
  NAND U19052 ( .A(n13347), .B(o[231]), .Z(n14077) );
  NAND U19053 ( .A(n13342), .B(creg[231]), .Z(n14076) );
  NAND U19054 ( .A(n14078), .B(n14079), .Z(c[230]) );
  NAND U19055 ( .A(n13347), .B(o[230]), .Z(n14079) );
  NAND U19056 ( .A(n13342), .B(creg[230]), .Z(n14078) );
  NAND U19057 ( .A(n14080), .B(n14081), .Z(c[22]) );
  NAND U19058 ( .A(n13347), .B(o[22]), .Z(n14081) );
  NAND U19059 ( .A(n13342), .B(creg[22]), .Z(n14080) );
  NAND U19060 ( .A(n14082), .B(n14083), .Z(c[229]) );
  NAND U19061 ( .A(n13347), .B(o[229]), .Z(n14083) );
  NAND U19062 ( .A(n13342), .B(creg[229]), .Z(n14082) );
  NAND U19063 ( .A(n14084), .B(n14085), .Z(c[228]) );
  NAND U19064 ( .A(n13347), .B(o[228]), .Z(n14085) );
  NAND U19065 ( .A(n13342), .B(creg[228]), .Z(n14084) );
  NAND U19066 ( .A(n14086), .B(n14087), .Z(c[227]) );
  NAND U19067 ( .A(n13347), .B(o[227]), .Z(n14087) );
  NAND U19068 ( .A(n13342), .B(creg[227]), .Z(n14086) );
  NAND U19069 ( .A(n14088), .B(n14089), .Z(c[226]) );
  NAND U19070 ( .A(n13347), .B(o[226]), .Z(n14089) );
  NAND U19071 ( .A(n13342), .B(creg[226]), .Z(n14088) );
  NAND U19072 ( .A(n14090), .B(n14091), .Z(c[225]) );
  NAND U19073 ( .A(n13347), .B(o[225]), .Z(n14091) );
  NAND U19074 ( .A(n13342), .B(creg[225]), .Z(n14090) );
  NAND U19075 ( .A(n14092), .B(n14093), .Z(c[224]) );
  NAND U19076 ( .A(n13347), .B(o[224]), .Z(n14093) );
  NAND U19077 ( .A(n13342), .B(creg[224]), .Z(n14092) );
  NAND U19078 ( .A(n14094), .B(n14095), .Z(c[223]) );
  NAND U19079 ( .A(n13347), .B(o[223]), .Z(n14095) );
  NAND U19080 ( .A(n13342), .B(creg[223]), .Z(n14094) );
  NAND U19081 ( .A(n14096), .B(n14097), .Z(c[222]) );
  NAND U19082 ( .A(n13347), .B(o[222]), .Z(n14097) );
  NAND U19083 ( .A(n13342), .B(creg[222]), .Z(n14096) );
  NAND U19084 ( .A(n14098), .B(n14099), .Z(c[221]) );
  NAND U19085 ( .A(n13347), .B(o[221]), .Z(n14099) );
  NAND U19086 ( .A(n13342), .B(creg[221]), .Z(n14098) );
  NAND U19087 ( .A(n14100), .B(n14101), .Z(c[220]) );
  NAND U19088 ( .A(n13347), .B(o[220]), .Z(n14101) );
  NAND U19089 ( .A(n13342), .B(creg[220]), .Z(n14100) );
  NAND U19090 ( .A(n14102), .B(n14103), .Z(c[21]) );
  NAND U19091 ( .A(n13347), .B(o[21]), .Z(n14103) );
  NAND U19092 ( .A(n13342), .B(creg[21]), .Z(n14102) );
  NAND U19093 ( .A(n14104), .B(n14105), .Z(c[219]) );
  NAND U19094 ( .A(n13347), .B(o[219]), .Z(n14105) );
  NAND U19095 ( .A(n13342), .B(creg[219]), .Z(n14104) );
  NAND U19096 ( .A(n14106), .B(n14107), .Z(c[218]) );
  NAND U19097 ( .A(n13347), .B(o[218]), .Z(n14107) );
  NAND U19098 ( .A(n13342), .B(creg[218]), .Z(n14106) );
  NAND U19099 ( .A(n14108), .B(n14109), .Z(c[217]) );
  NAND U19100 ( .A(n13347), .B(o[217]), .Z(n14109) );
  NAND U19101 ( .A(n13342), .B(creg[217]), .Z(n14108) );
  NAND U19102 ( .A(n14110), .B(n14111), .Z(c[216]) );
  NAND U19103 ( .A(n13347), .B(o[216]), .Z(n14111) );
  NAND U19104 ( .A(n13342), .B(creg[216]), .Z(n14110) );
  NAND U19105 ( .A(n14112), .B(n14113), .Z(c[215]) );
  NAND U19106 ( .A(n13347), .B(o[215]), .Z(n14113) );
  NAND U19107 ( .A(n13342), .B(creg[215]), .Z(n14112) );
  NAND U19108 ( .A(n14114), .B(n14115), .Z(c[214]) );
  NAND U19109 ( .A(n13347), .B(o[214]), .Z(n14115) );
  NAND U19110 ( .A(n13342), .B(creg[214]), .Z(n14114) );
  NAND U19111 ( .A(n14116), .B(n14117), .Z(c[213]) );
  NAND U19112 ( .A(n13347), .B(o[213]), .Z(n14117) );
  NAND U19113 ( .A(n13342), .B(creg[213]), .Z(n14116) );
  NAND U19114 ( .A(n14118), .B(n14119), .Z(c[212]) );
  NAND U19115 ( .A(n13347), .B(o[212]), .Z(n14119) );
  NAND U19116 ( .A(n13342), .B(creg[212]), .Z(n14118) );
  NAND U19117 ( .A(n14120), .B(n14121), .Z(c[211]) );
  NAND U19118 ( .A(n13347), .B(o[211]), .Z(n14121) );
  NAND U19119 ( .A(n13342), .B(creg[211]), .Z(n14120) );
  NAND U19120 ( .A(n14122), .B(n14123), .Z(c[210]) );
  NAND U19121 ( .A(n13347), .B(o[210]), .Z(n14123) );
  NAND U19122 ( .A(n13342), .B(creg[210]), .Z(n14122) );
  NAND U19123 ( .A(n14124), .B(n14125), .Z(c[20]) );
  NAND U19124 ( .A(n13347), .B(o[20]), .Z(n14125) );
  NAND U19125 ( .A(n13342), .B(creg[20]), .Z(n14124) );
  NAND U19126 ( .A(n14126), .B(n14127), .Z(c[209]) );
  NAND U19127 ( .A(n13347), .B(o[209]), .Z(n14127) );
  NAND U19128 ( .A(n13342), .B(creg[209]), .Z(n14126) );
  NAND U19129 ( .A(n14128), .B(n14129), .Z(c[208]) );
  NAND U19130 ( .A(n13347), .B(o[208]), .Z(n14129) );
  NAND U19131 ( .A(n13342), .B(creg[208]), .Z(n14128) );
  NAND U19132 ( .A(n14130), .B(n14131), .Z(c[207]) );
  NAND U19133 ( .A(n13347), .B(o[207]), .Z(n14131) );
  NAND U19134 ( .A(n13342), .B(creg[207]), .Z(n14130) );
  NAND U19135 ( .A(n14132), .B(n14133), .Z(c[206]) );
  NAND U19136 ( .A(n13347), .B(o[206]), .Z(n14133) );
  NAND U19137 ( .A(n13342), .B(creg[206]), .Z(n14132) );
  NAND U19138 ( .A(n14134), .B(n14135), .Z(c[205]) );
  NAND U19139 ( .A(n13347), .B(o[205]), .Z(n14135) );
  NAND U19140 ( .A(n13342), .B(creg[205]), .Z(n14134) );
  NAND U19141 ( .A(n14136), .B(n14137), .Z(c[204]) );
  NAND U19142 ( .A(n13347), .B(o[204]), .Z(n14137) );
  NAND U19143 ( .A(n13342), .B(creg[204]), .Z(n14136) );
  NAND U19144 ( .A(n14138), .B(n14139), .Z(c[203]) );
  NAND U19145 ( .A(n13347), .B(o[203]), .Z(n14139) );
  NAND U19146 ( .A(n13342), .B(creg[203]), .Z(n14138) );
  NAND U19147 ( .A(n14140), .B(n14141), .Z(c[202]) );
  NAND U19148 ( .A(n13347), .B(o[202]), .Z(n14141) );
  NAND U19149 ( .A(n13342), .B(creg[202]), .Z(n14140) );
  NAND U19150 ( .A(n14142), .B(n14143), .Z(c[201]) );
  NAND U19151 ( .A(n13347), .B(o[201]), .Z(n14143) );
  NAND U19152 ( .A(n13342), .B(creg[201]), .Z(n14142) );
  NAND U19153 ( .A(n14144), .B(n14145), .Z(c[200]) );
  NAND U19154 ( .A(n13347), .B(o[200]), .Z(n14145) );
  NAND U19155 ( .A(n13342), .B(creg[200]), .Z(n14144) );
  NAND U19156 ( .A(n14146), .B(n14147), .Z(c[1]) );
  NAND U19157 ( .A(n13347), .B(o[1]), .Z(n14147) );
  NAND U19158 ( .A(n13342), .B(creg[1]), .Z(n14146) );
  NAND U19159 ( .A(n14148), .B(n14149), .Z(c[19]) );
  NAND U19160 ( .A(n13347), .B(o[19]), .Z(n14149) );
  NAND U19161 ( .A(n13342), .B(creg[19]), .Z(n14148) );
  NAND U19162 ( .A(n14150), .B(n14151), .Z(c[199]) );
  NAND U19163 ( .A(n13347), .B(o[199]), .Z(n14151) );
  NAND U19164 ( .A(n13342), .B(creg[199]), .Z(n14150) );
  NAND U19165 ( .A(n14152), .B(n14153), .Z(c[198]) );
  NAND U19166 ( .A(n13347), .B(o[198]), .Z(n14153) );
  NAND U19167 ( .A(n13342), .B(creg[198]), .Z(n14152) );
  NAND U19168 ( .A(n14154), .B(n14155), .Z(c[197]) );
  NAND U19169 ( .A(n13347), .B(o[197]), .Z(n14155) );
  NAND U19170 ( .A(n13342), .B(creg[197]), .Z(n14154) );
  NAND U19171 ( .A(n14156), .B(n14157), .Z(c[196]) );
  NAND U19172 ( .A(n13347), .B(o[196]), .Z(n14157) );
  NAND U19173 ( .A(n13342), .B(creg[196]), .Z(n14156) );
  NAND U19174 ( .A(n14158), .B(n14159), .Z(c[195]) );
  NAND U19175 ( .A(n13347), .B(o[195]), .Z(n14159) );
  NAND U19176 ( .A(n13342), .B(creg[195]), .Z(n14158) );
  NAND U19177 ( .A(n14160), .B(n14161), .Z(c[194]) );
  NAND U19178 ( .A(n13347), .B(o[194]), .Z(n14161) );
  NAND U19179 ( .A(n13342), .B(creg[194]), .Z(n14160) );
  NAND U19180 ( .A(n14162), .B(n14163), .Z(c[193]) );
  NAND U19181 ( .A(n13347), .B(o[193]), .Z(n14163) );
  NAND U19182 ( .A(n13342), .B(creg[193]), .Z(n14162) );
  NAND U19183 ( .A(n14164), .B(n14165), .Z(c[192]) );
  NAND U19184 ( .A(n13347), .B(o[192]), .Z(n14165) );
  NAND U19185 ( .A(n13342), .B(creg[192]), .Z(n14164) );
  NAND U19186 ( .A(n14166), .B(n14167), .Z(c[191]) );
  NAND U19187 ( .A(n13347), .B(o[191]), .Z(n14167) );
  NAND U19188 ( .A(n13342), .B(creg[191]), .Z(n14166) );
  NAND U19189 ( .A(n14168), .B(n14169), .Z(c[190]) );
  NAND U19190 ( .A(n13347), .B(o[190]), .Z(n14169) );
  NAND U19191 ( .A(n13342), .B(creg[190]), .Z(n14168) );
  NAND U19192 ( .A(n14170), .B(n14171), .Z(c[18]) );
  NAND U19193 ( .A(n13347), .B(o[18]), .Z(n14171) );
  NAND U19194 ( .A(n13342), .B(creg[18]), .Z(n14170) );
  NAND U19195 ( .A(n14172), .B(n14173), .Z(c[189]) );
  NAND U19196 ( .A(n13347), .B(o[189]), .Z(n14173) );
  NAND U19197 ( .A(n13342), .B(creg[189]), .Z(n14172) );
  NAND U19198 ( .A(n14174), .B(n14175), .Z(c[188]) );
  NAND U19199 ( .A(n13347), .B(o[188]), .Z(n14175) );
  NAND U19200 ( .A(n13342), .B(creg[188]), .Z(n14174) );
  NAND U19201 ( .A(n14176), .B(n14177), .Z(c[187]) );
  NAND U19202 ( .A(n13347), .B(o[187]), .Z(n14177) );
  NAND U19203 ( .A(n13342), .B(creg[187]), .Z(n14176) );
  NAND U19204 ( .A(n14178), .B(n14179), .Z(c[186]) );
  NAND U19205 ( .A(n13347), .B(o[186]), .Z(n14179) );
  NAND U19206 ( .A(n13342), .B(creg[186]), .Z(n14178) );
  NAND U19207 ( .A(n14180), .B(n14181), .Z(c[185]) );
  NAND U19208 ( .A(n13347), .B(o[185]), .Z(n14181) );
  NAND U19209 ( .A(n13342), .B(creg[185]), .Z(n14180) );
  NAND U19210 ( .A(n14182), .B(n14183), .Z(c[184]) );
  NAND U19211 ( .A(n13347), .B(o[184]), .Z(n14183) );
  NAND U19212 ( .A(n13342), .B(creg[184]), .Z(n14182) );
  NAND U19213 ( .A(n14184), .B(n14185), .Z(c[183]) );
  NAND U19214 ( .A(n13347), .B(o[183]), .Z(n14185) );
  NAND U19215 ( .A(n13342), .B(creg[183]), .Z(n14184) );
  NAND U19216 ( .A(n14186), .B(n14187), .Z(c[182]) );
  NAND U19217 ( .A(n13347), .B(o[182]), .Z(n14187) );
  NAND U19218 ( .A(n13342), .B(creg[182]), .Z(n14186) );
  NAND U19219 ( .A(n14188), .B(n14189), .Z(c[181]) );
  NAND U19220 ( .A(n13347), .B(o[181]), .Z(n14189) );
  NAND U19221 ( .A(n13342), .B(creg[181]), .Z(n14188) );
  NAND U19222 ( .A(n14190), .B(n14191), .Z(c[180]) );
  NAND U19223 ( .A(n13347), .B(o[180]), .Z(n14191) );
  NAND U19224 ( .A(n13342), .B(creg[180]), .Z(n14190) );
  NAND U19225 ( .A(n14192), .B(n14193), .Z(c[17]) );
  NAND U19226 ( .A(n13347), .B(o[17]), .Z(n14193) );
  NAND U19227 ( .A(n13342), .B(creg[17]), .Z(n14192) );
  NAND U19228 ( .A(n14194), .B(n14195), .Z(c[179]) );
  NAND U19229 ( .A(n13347), .B(o[179]), .Z(n14195) );
  NAND U19230 ( .A(n13342), .B(creg[179]), .Z(n14194) );
  NAND U19231 ( .A(n14196), .B(n14197), .Z(c[178]) );
  NAND U19232 ( .A(n13347), .B(o[178]), .Z(n14197) );
  NAND U19233 ( .A(n13342), .B(creg[178]), .Z(n14196) );
  NAND U19234 ( .A(n14198), .B(n14199), .Z(c[177]) );
  NAND U19235 ( .A(n13347), .B(o[177]), .Z(n14199) );
  NAND U19236 ( .A(n13342), .B(creg[177]), .Z(n14198) );
  NAND U19237 ( .A(n14200), .B(n14201), .Z(c[176]) );
  NAND U19238 ( .A(n13347), .B(o[176]), .Z(n14201) );
  NAND U19239 ( .A(n13342), .B(creg[176]), .Z(n14200) );
  NAND U19240 ( .A(n14202), .B(n14203), .Z(c[175]) );
  NAND U19241 ( .A(n13347), .B(o[175]), .Z(n14203) );
  NAND U19242 ( .A(n13342), .B(creg[175]), .Z(n14202) );
  NAND U19243 ( .A(n14204), .B(n14205), .Z(c[174]) );
  NAND U19244 ( .A(n13347), .B(o[174]), .Z(n14205) );
  NAND U19245 ( .A(n13342), .B(creg[174]), .Z(n14204) );
  NAND U19246 ( .A(n14206), .B(n14207), .Z(c[173]) );
  NAND U19247 ( .A(n13347), .B(o[173]), .Z(n14207) );
  NAND U19248 ( .A(n13342), .B(creg[173]), .Z(n14206) );
  NAND U19249 ( .A(n14208), .B(n14209), .Z(c[172]) );
  NAND U19250 ( .A(n13347), .B(o[172]), .Z(n14209) );
  NAND U19251 ( .A(n13342), .B(creg[172]), .Z(n14208) );
  NAND U19252 ( .A(n14210), .B(n14211), .Z(c[171]) );
  NAND U19253 ( .A(n13347), .B(o[171]), .Z(n14211) );
  NAND U19254 ( .A(n13342), .B(creg[171]), .Z(n14210) );
  NAND U19255 ( .A(n14212), .B(n14213), .Z(c[170]) );
  NAND U19256 ( .A(n13347), .B(o[170]), .Z(n14213) );
  NAND U19257 ( .A(n13342), .B(creg[170]), .Z(n14212) );
  NAND U19258 ( .A(n14214), .B(n14215), .Z(c[16]) );
  NAND U19259 ( .A(n13347), .B(o[16]), .Z(n14215) );
  NAND U19260 ( .A(n13342), .B(creg[16]), .Z(n14214) );
  NAND U19261 ( .A(n14216), .B(n14217), .Z(c[169]) );
  NAND U19262 ( .A(n13347), .B(o[169]), .Z(n14217) );
  NAND U19263 ( .A(n13342), .B(creg[169]), .Z(n14216) );
  NAND U19264 ( .A(n14218), .B(n14219), .Z(c[168]) );
  NAND U19265 ( .A(n13347), .B(o[168]), .Z(n14219) );
  NAND U19266 ( .A(n13342), .B(creg[168]), .Z(n14218) );
  NAND U19267 ( .A(n14220), .B(n14221), .Z(c[167]) );
  NAND U19268 ( .A(n13347), .B(o[167]), .Z(n14221) );
  NAND U19269 ( .A(n13342), .B(creg[167]), .Z(n14220) );
  NAND U19270 ( .A(n14222), .B(n14223), .Z(c[166]) );
  NAND U19271 ( .A(n13347), .B(o[166]), .Z(n14223) );
  NAND U19272 ( .A(n13342), .B(creg[166]), .Z(n14222) );
  NAND U19273 ( .A(n14224), .B(n14225), .Z(c[165]) );
  NAND U19274 ( .A(n13347), .B(o[165]), .Z(n14225) );
  NAND U19275 ( .A(n13342), .B(creg[165]), .Z(n14224) );
  NAND U19276 ( .A(n14226), .B(n14227), .Z(c[164]) );
  NAND U19277 ( .A(n13347), .B(o[164]), .Z(n14227) );
  NAND U19278 ( .A(n13342), .B(creg[164]), .Z(n14226) );
  NAND U19279 ( .A(n14228), .B(n14229), .Z(c[163]) );
  NAND U19280 ( .A(n13347), .B(o[163]), .Z(n14229) );
  NAND U19281 ( .A(n13342), .B(creg[163]), .Z(n14228) );
  NAND U19282 ( .A(n14230), .B(n14231), .Z(c[162]) );
  NAND U19283 ( .A(n13347), .B(o[162]), .Z(n14231) );
  NAND U19284 ( .A(n13342), .B(creg[162]), .Z(n14230) );
  NAND U19285 ( .A(n14232), .B(n14233), .Z(c[161]) );
  NAND U19286 ( .A(n13347), .B(o[161]), .Z(n14233) );
  NAND U19287 ( .A(n13342), .B(creg[161]), .Z(n14232) );
  NAND U19288 ( .A(n14234), .B(n14235), .Z(c[160]) );
  NAND U19289 ( .A(n13347), .B(o[160]), .Z(n14235) );
  NAND U19290 ( .A(n13342), .B(creg[160]), .Z(n14234) );
  NAND U19291 ( .A(n14236), .B(n14237), .Z(c[15]) );
  NAND U19292 ( .A(n13347), .B(o[15]), .Z(n14237) );
  NAND U19293 ( .A(n13342), .B(creg[15]), .Z(n14236) );
  NAND U19294 ( .A(n14238), .B(n14239), .Z(c[159]) );
  NAND U19295 ( .A(n13347), .B(o[159]), .Z(n14239) );
  NAND U19296 ( .A(n13342), .B(creg[159]), .Z(n14238) );
  NAND U19297 ( .A(n14240), .B(n14241), .Z(c[158]) );
  NAND U19298 ( .A(n13347), .B(o[158]), .Z(n14241) );
  NAND U19299 ( .A(n13342), .B(creg[158]), .Z(n14240) );
  NAND U19300 ( .A(n14242), .B(n14243), .Z(c[157]) );
  NAND U19301 ( .A(n13347), .B(o[157]), .Z(n14243) );
  NAND U19302 ( .A(n13342), .B(creg[157]), .Z(n14242) );
  NAND U19303 ( .A(n14244), .B(n14245), .Z(c[156]) );
  NAND U19304 ( .A(n13347), .B(o[156]), .Z(n14245) );
  NAND U19305 ( .A(n13342), .B(creg[156]), .Z(n14244) );
  NAND U19306 ( .A(n14246), .B(n14247), .Z(c[155]) );
  NAND U19307 ( .A(n13347), .B(o[155]), .Z(n14247) );
  NAND U19308 ( .A(n13342), .B(creg[155]), .Z(n14246) );
  NAND U19309 ( .A(n14248), .B(n14249), .Z(c[154]) );
  NAND U19310 ( .A(n13347), .B(o[154]), .Z(n14249) );
  NAND U19311 ( .A(n13342), .B(creg[154]), .Z(n14248) );
  NAND U19312 ( .A(n14250), .B(n14251), .Z(c[153]) );
  NAND U19313 ( .A(n13347), .B(o[153]), .Z(n14251) );
  NAND U19314 ( .A(n13342), .B(creg[153]), .Z(n14250) );
  NAND U19315 ( .A(n14252), .B(n14253), .Z(c[152]) );
  NAND U19316 ( .A(n13347), .B(o[152]), .Z(n14253) );
  NAND U19317 ( .A(n13342), .B(creg[152]), .Z(n14252) );
  NAND U19318 ( .A(n14254), .B(n14255), .Z(c[151]) );
  NAND U19319 ( .A(n13347), .B(o[151]), .Z(n14255) );
  NAND U19320 ( .A(n13342), .B(creg[151]), .Z(n14254) );
  NAND U19321 ( .A(n14256), .B(n14257), .Z(c[150]) );
  NAND U19322 ( .A(n13347), .B(o[150]), .Z(n14257) );
  NAND U19323 ( .A(n13342), .B(creg[150]), .Z(n14256) );
  NAND U19324 ( .A(n14258), .B(n14259), .Z(c[14]) );
  NAND U19325 ( .A(n13347), .B(o[14]), .Z(n14259) );
  NAND U19326 ( .A(n13342), .B(creg[14]), .Z(n14258) );
  NAND U19327 ( .A(n14260), .B(n14261), .Z(c[149]) );
  NAND U19328 ( .A(n13347), .B(o[149]), .Z(n14261) );
  NAND U19329 ( .A(n13342), .B(creg[149]), .Z(n14260) );
  NAND U19330 ( .A(n14262), .B(n14263), .Z(c[148]) );
  NAND U19331 ( .A(n13347), .B(o[148]), .Z(n14263) );
  NAND U19332 ( .A(n13342), .B(creg[148]), .Z(n14262) );
  NAND U19333 ( .A(n14264), .B(n14265), .Z(c[147]) );
  NAND U19334 ( .A(n13347), .B(o[147]), .Z(n14265) );
  NAND U19335 ( .A(n13342), .B(creg[147]), .Z(n14264) );
  NAND U19336 ( .A(n14266), .B(n14267), .Z(c[146]) );
  NAND U19337 ( .A(n13347), .B(o[146]), .Z(n14267) );
  NAND U19338 ( .A(n13342), .B(creg[146]), .Z(n14266) );
  NAND U19339 ( .A(n14268), .B(n14269), .Z(c[145]) );
  NAND U19340 ( .A(n13347), .B(o[145]), .Z(n14269) );
  NAND U19341 ( .A(n13342), .B(creg[145]), .Z(n14268) );
  NAND U19342 ( .A(n14270), .B(n14271), .Z(c[144]) );
  NAND U19343 ( .A(n13347), .B(o[144]), .Z(n14271) );
  NAND U19344 ( .A(n13342), .B(creg[144]), .Z(n14270) );
  NAND U19345 ( .A(n14272), .B(n14273), .Z(c[143]) );
  NAND U19346 ( .A(n13347), .B(o[143]), .Z(n14273) );
  NAND U19347 ( .A(n13342), .B(creg[143]), .Z(n14272) );
  NAND U19348 ( .A(n14274), .B(n14275), .Z(c[142]) );
  NAND U19349 ( .A(n13347), .B(o[142]), .Z(n14275) );
  NAND U19350 ( .A(n13342), .B(creg[142]), .Z(n14274) );
  NAND U19351 ( .A(n14276), .B(n14277), .Z(c[141]) );
  NAND U19352 ( .A(n13347), .B(o[141]), .Z(n14277) );
  NAND U19353 ( .A(n13342), .B(creg[141]), .Z(n14276) );
  NAND U19354 ( .A(n14278), .B(n14279), .Z(c[140]) );
  NAND U19355 ( .A(n13347), .B(o[140]), .Z(n14279) );
  NAND U19356 ( .A(n13342), .B(creg[140]), .Z(n14278) );
  NAND U19357 ( .A(n14280), .B(n14281), .Z(c[13]) );
  NAND U19358 ( .A(n13347), .B(o[13]), .Z(n14281) );
  NAND U19359 ( .A(n13342), .B(creg[13]), .Z(n14280) );
  NAND U19360 ( .A(n14282), .B(n14283), .Z(c[139]) );
  NAND U19361 ( .A(n13347), .B(o[139]), .Z(n14283) );
  NAND U19362 ( .A(n13342), .B(creg[139]), .Z(n14282) );
  NAND U19363 ( .A(n14284), .B(n14285), .Z(c[138]) );
  NAND U19364 ( .A(n13347), .B(o[138]), .Z(n14285) );
  NAND U19365 ( .A(n13342), .B(creg[138]), .Z(n14284) );
  NAND U19366 ( .A(n14286), .B(n14287), .Z(c[137]) );
  NAND U19367 ( .A(n13347), .B(o[137]), .Z(n14287) );
  NAND U19368 ( .A(n13342), .B(creg[137]), .Z(n14286) );
  NAND U19369 ( .A(n14288), .B(n14289), .Z(c[136]) );
  NAND U19370 ( .A(n13347), .B(o[136]), .Z(n14289) );
  NAND U19371 ( .A(n13342), .B(creg[136]), .Z(n14288) );
  NAND U19372 ( .A(n14290), .B(n14291), .Z(c[135]) );
  NAND U19373 ( .A(n13347), .B(o[135]), .Z(n14291) );
  NAND U19374 ( .A(n13342), .B(creg[135]), .Z(n14290) );
  NAND U19375 ( .A(n14292), .B(n14293), .Z(c[134]) );
  NAND U19376 ( .A(n13347), .B(o[134]), .Z(n14293) );
  NAND U19377 ( .A(n13342), .B(creg[134]), .Z(n14292) );
  NAND U19378 ( .A(n14294), .B(n14295), .Z(c[133]) );
  NAND U19379 ( .A(n13347), .B(o[133]), .Z(n14295) );
  NAND U19380 ( .A(n13342), .B(creg[133]), .Z(n14294) );
  NAND U19381 ( .A(n14296), .B(n14297), .Z(c[132]) );
  NAND U19382 ( .A(n13347), .B(o[132]), .Z(n14297) );
  NAND U19383 ( .A(n13342), .B(creg[132]), .Z(n14296) );
  NAND U19384 ( .A(n14298), .B(n14299), .Z(c[131]) );
  NAND U19385 ( .A(n13347), .B(o[131]), .Z(n14299) );
  NAND U19386 ( .A(n13342), .B(creg[131]), .Z(n14298) );
  NAND U19387 ( .A(n14300), .B(n14301), .Z(c[130]) );
  NAND U19388 ( .A(n13347), .B(o[130]), .Z(n14301) );
  NAND U19389 ( .A(n13342), .B(creg[130]), .Z(n14300) );
  NAND U19390 ( .A(n14302), .B(n14303), .Z(c[12]) );
  NAND U19391 ( .A(n13347), .B(o[12]), .Z(n14303) );
  NAND U19392 ( .A(n13342), .B(creg[12]), .Z(n14302) );
  NAND U19393 ( .A(n14304), .B(n14305), .Z(c[129]) );
  NAND U19394 ( .A(n13347), .B(o[129]), .Z(n14305) );
  NAND U19395 ( .A(n13342), .B(creg[129]), .Z(n14304) );
  NAND U19396 ( .A(n14306), .B(n14307), .Z(c[128]) );
  NAND U19397 ( .A(n13347), .B(o[128]), .Z(n14307) );
  NAND U19398 ( .A(n13342), .B(creg[128]), .Z(n14306) );
  NAND U19399 ( .A(n14308), .B(n14309), .Z(c[127]) );
  NAND U19400 ( .A(n13347), .B(o[127]), .Z(n14309) );
  NAND U19401 ( .A(n13342), .B(creg[127]), .Z(n14308) );
  NAND U19402 ( .A(n14310), .B(n14311), .Z(c[126]) );
  NAND U19403 ( .A(n13347), .B(o[126]), .Z(n14311) );
  NAND U19404 ( .A(n13342), .B(creg[126]), .Z(n14310) );
  NAND U19405 ( .A(n14312), .B(n14313), .Z(c[125]) );
  NAND U19406 ( .A(n13347), .B(o[125]), .Z(n14313) );
  NAND U19407 ( .A(n13342), .B(creg[125]), .Z(n14312) );
  NAND U19408 ( .A(n14314), .B(n14315), .Z(c[124]) );
  NAND U19409 ( .A(n13347), .B(o[124]), .Z(n14315) );
  NAND U19410 ( .A(n13342), .B(creg[124]), .Z(n14314) );
  NAND U19411 ( .A(n14316), .B(n14317), .Z(c[123]) );
  NAND U19412 ( .A(n13347), .B(o[123]), .Z(n14317) );
  NAND U19413 ( .A(n13342), .B(creg[123]), .Z(n14316) );
  NAND U19414 ( .A(n14318), .B(n14319), .Z(c[122]) );
  NAND U19415 ( .A(n13347), .B(o[122]), .Z(n14319) );
  NAND U19416 ( .A(n13342), .B(creg[122]), .Z(n14318) );
  NAND U19417 ( .A(n14320), .B(n14321), .Z(c[121]) );
  NAND U19418 ( .A(n13347), .B(o[121]), .Z(n14321) );
  NAND U19419 ( .A(n13342), .B(creg[121]), .Z(n14320) );
  NAND U19420 ( .A(n14322), .B(n14323), .Z(c[120]) );
  NAND U19421 ( .A(n13347), .B(o[120]), .Z(n14323) );
  NAND U19422 ( .A(n13342), .B(creg[120]), .Z(n14322) );
  NAND U19423 ( .A(n14324), .B(n14325), .Z(c[11]) );
  NAND U19424 ( .A(n13347), .B(o[11]), .Z(n14325) );
  NAND U19425 ( .A(n13342), .B(creg[11]), .Z(n14324) );
  NAND U19426 ( .A(n14326), .B(n14327), .Z(c[119]) );
  NAND U19427 ( .A(n13347), .B(o[119]), .Z(n14327) );
  NAND U19428 ( .A(n13342), .B(creg[119]), .Z(n14326) );
  NAND U19429 ( .A(n14328), .B(n14329), .Z(c[118]) );
  NAND U19430 ( .A(n13347), .B(o[118]), .Z(n14329) );
  NAND U19431 ( .A(n13342), .B(creg[118]), .Z(n14328) );
  NAND U19432 ( .A(n14330), .B(n14331), .Z(c[117]) );
  NAND U19433 ( .A(n13347), .B(o[117]), .Z(n14331) );
  NAND U19434 ( .A(n13342), .B(creg[117]), .Z(n14330) );
  NAND U19435 ( .A(n14332), .B(n14333), .Z(c[116]) );
  NAND U19436 ( .A(n13347), .B(o[116]), .Z(n14333) );
  NAND U19437 ( .A(n13342), .B(creg[116]), .Z(n14332) );
  NAND U19438 ( .A(n14334), .B(n14335), .Z(c[115]) );
  NAND U19439 ( .A(n13347), .B(o[115]), .Z(n14335) );
  NAND U19440 ( .A(n13342), .B(creg[115]), .Z(n14334) );
  NAND U19441 ( .A(n14336), .B(n14337), .Z(c[114]) );
  NAND U19442 ( .A(n13347), .B(o[114]), .Z(n14337) );
  NAND U19443 ( .A(n13342), .B(creg[114]), .Z(n14336) );
  NAND U19444 ( .A(n14338), .B(n14339), .Z(c[113]) );
  NAND U19445 ( .A(n13347), .B(o[113]), .Z(n14339) );
  NAND U19446 ( .A(n13342), .B(creg[113]), .Z(n14338) );
  NAND U19447 ( .A(n14340), .B(n14341), .Z(c[112]) );
  NAND U19448 ( .A(n13347), .B(o[112]), .Z(n14341) );
  NAND U19449 ( .A(n13342), .B(creg[112]), .Z(n14340) );
  NAND U19450 ( .A(n14342), .B(n14343), .Z(c[111]) );
  NAND U19451 ( .A(n13347), .B(o[111]), .Z(n14343) );
  NAND U19452 ( .A(n13342), .B(creg[111]), .Z(n14342) );
  NAND U19453 ( .A(n14344), .B(n14345), .Z(c[110]) );
  NAND U19454 ( .A(n13347), .B(o[110]), .Z(n14345) );
  NAND U19455 ( .A(n13342), .B(creg[110]), .Z(n14344) );
  NAND U19456 ( .A(n14346), .B(n14347), .Z(c[10]) );
  NAND U19457 ( .A(n13347), .B(o[10]), .Z(n14347) );
  NAND U19458 ( .A(n13342), .B(creg[10]), .Z(n14346) );
  NAND U19459 ( .A(n14348), .B(n14349), .Z(c[109]) );
  NAND U19460 ( .A(n13347), .B(o[109]), .Z(n14349) );
  NAND U19461 ( .A(n13342), .B(creg[109]), .Z(n14348) );
  NAND U19462 ( .A(n14350), .B(n14351), .Z(c[108]) );
  NAND U19463 ( .A(n13347), .B(o[108]), .Z(n14351) );
  NAND U19464 ( .A(n13342), .B(creg[108]), .Z(n14350) );
  NAND U19465 ( .A(n14352), .B(n14353), .Z(c[107]) );
  NAND U19466 ( .A(n13347), .B(o[107]), .Z(n14353) );
  NAND U19467 ( .A(n13342), .B(creg[107]), .Z(n14352) );
  NAND U19468 ( .A(n14354), .B(n14355), .Z(c[106]) );
  NAND U19469 ( .A(n13347), .B(o[106]), .Z(n14355) );
  NAND U19470 ( .A(n13342), .B(creg[106]), .Z(n14354) );
  NAND U19471 ( .A(n14356), .B(n14357), .Z(c[105]) );
  NAND U19472 ( .A(n13347), .B(o[105]), .Z(n14357) );
  NAND U19473 ( .A(n13342), .B(creg[105]), .Z(n14356) );
  NAND U19474 ( .A(n14358), .B(n14359), .Z(c[104]) );
  NAND U19475 ( .A(n13347), .B(o[104]), .Z(n14359) );
  NAND U19476 ( .A(n13342), .B(creg[104]), .Z(n14358) );
  NAND U19477 ( .A(n14360), .B(n14361), .Z(c[103]) );
  NAND U19478 ( .A(n13347), .B(o[103]), .Z(n14361) );
  NAND U19479 ( .A(n13342), .B(creg[103]), .Z(n14360) );
  NAND U19480 ( .A(n14362), .B(n14363), .Z(c[102]) );
  NAND U19481 ( .A(n13347), .B(o[102]), .Z(n14363) );
  NAND U19482 ( .A(n13342), .B(creg[102]), .Z(n14362) );
  NAND U19483 ( .A(n14364), .B(n14365), .Z(c[101]) );
  NAND U19484 ( .A(n13347), .B(o[101]), .Z(n14365) );
  NAND U19485 ( .A(n13342), .B(creg[101]), .Z(n14364) );
  NAND U19486 ( .A(n14366), .B(n14367), .Z(c[100]) );
  NAND U19487 ( .A(n13347), .B(o[100]), .Z(n14367) );
  NAND U19488 ( .A(n13342), .B(creg[100]), .Z(n14366) );
  NAND U19489 ( .A(n14368), .B(n14369), .Z(c[0]) );
  NAND U19490 ( .A(n13347), .B(o[0]), .Z(n14369) );
  IV U19491 ( .A(n13342), .Z(n13347) );
  NAND U19492 ( .A(n13342), .B(creg[0]), .Z(n14368) );
  NAND U19493 ( .A(n14370), .B(n14371), .Z(n13342) );
  NANDN U19494 ( .A(ereg[511]), .B(init), .Z(n14371) );
  OR U19495 ( .A(init), .B(e[511]), .Z(n14370) );
endmodule

