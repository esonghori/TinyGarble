
module k_nns_seq_W31_K4 ( clk, rst, g_input, e_input, o );
  input [30:0] g_input;
  input [30:0] e_input;
  output [123:0] o;
  input clk, rst;
  wire   \min_dist_reg[3][4] , \min_dist_reg[3][3] , \min_dist_reg[3][2] ,
         \min_dist_reg[3][1] , \min_dist_reg[3][0] , \min_dist_reg[2][4] ,
         \min_dist_reg[2][3] , \min_dist_reg[2][2] , \min_dist_reg[2][1] ,
         \min_dist_reg[2][0] , \min_dist_reg[1][4] , \min_dist_reg[1][3] ,
         \min_dist_reg[1][2] , \min_dist_reg[1][1] , \min_dist_reg[1][0] ,
         \min_dist_reg[0][4] , \min_dist_reg[0][3] , \min_dist_reg[0][2] ,
         \min_dist_reg[0][1] , \min_dist_reg[0][0] , \local_min_dist[0][4] ,
         \local_min_dist[0][3] , \local_min_dist[0][2] ,
         \local_min_dist[0][1] , \local_min_dist[0][0] , \min_dist[3][4] ,
         \min_dist[3][3] , \min_dist[3][2] , \min_dist[3][1] ,
         \min_dist[3][0] , \min_dist[2][4] , \min_dist[2][3] ,
         \min_dist[2][2] , \min_dist[2][1] , \min_dist[2][0] ,
         \min_dist[1][4] , \min_dist[1][3] , \min_dist[1][2] ,
         \min_dist[1][1] , \min_dist[1][0] , \min_val_reg[3][30] ,
         \min_val_reg[3][29] , \min_val_reg[3][28] , \min_val_reg[3][27] ,
         \min_val_reg[3][26] , \min_val_reg[3][25] , \min_val_reg[3][24] ,
         \min_val_reg[3][23] , \min_val_reg[3][22] , \min_val_reg[3][21] ,
         \min_val_reg[3][20] , \min_val_reg[3][19] , \min_val_reg[3][18] ,
         \min_val_reg[3][17] , \min_val_reg[3][16] , \min_val_reg[3][15] ,
         \min_val_reg[3][14] , \min_val_reg[3][13] , \min_val_reg[3][12] ,
         \min_val_reg[3][11] , \min_val_reg[3][10] , \min_val_reg[3][9] ,
         \min_val_reg[3][8] , \min_val_reg[3][7] , \min_val_reg[3][6] ,
         \min_val_reg[3][5] , \min_val_reg[3][4] , \min_val_reg[3][3] ,
         \min_val_reg[3][2] , \min_val_reg[3][1] , \min_val_reg[3][0] ,
         \min_val_reg[2][30] , \min_val_reg[2][29] , \min_val_reg[2][28] ,
         \min_val_reg[2][27] , \min_val_reg[2][26] , \min_val_reg[2][25] ,
         \min_val_reg[2][24] , \min_val_reg[2][23] , \min_val_reg[2][22] ,
         \min_val_reg[2][21] , \min_val_reg[2][20] , \min_val_reg[2][19] ,
         \min_val_reg[2][18] , \min_val_reg[2][17] , \min_val_reg[2][16] ,
         \min_val_reg[2][15] , \min_val_reg[2][14] , \min_val_reg[2][13] ,
         \min_val_reg[2][12] , \min_val_reg[2][11] , \min_val_reg[2][10] ,
         \min_val_reg[2][9] , \min_val_reg[2][8] , \min_val_reg[2][7] ,
         \min_val_reg[2][6] , \min_val_reg[2][5] , \min_val_reg[2][4] ,
         \min_val_reg[2][3] , \min_val_reg[2][2] , \min_val_reg[2][1] ,
         \min_val_reg[2][0] , \min_val_reg[1][30] , \min_val_reg[1][29] ,
         \min_val_reg[1][28] , \min_val_reg[1][27] , \min_val_reg[1][26] ,
         \min_val_reg[1][25] , \min_val_reg[1][24] , \min_val_reg[1][23] ,
         \min_val_reg[1][22] , \min_val_reg[1][21] , \min_val_reg[1][20] ,
         \min_val_reg[1][19] , \min_val_reg[1][18] , \min_val_reg[1][17] ,
         \min_val_reg[1][16] , \min_val_reg[1][15] , \min_val_reg[1][14] ,
         \min_val_reg[1][13] , \min_val_reg[1][12] , \min_val_reg[1][11] ,
         \min_val_reg[1][10] , \min_val_reg[1][9] , \min_val_reg[1][8] ,
         \min_val_reg[1][7] , \min_val_reg[1][6] , \min_val_reg[1][5] ,
         \min_val_reg[1][4] , \min_val_reg[1][3] , \min_val_reg[1][2] ,
         \min_val_reg[1][1] , \min_val_reg[1][0] , \min_val_reg[0][30] ,
         \min_val_reg[0][29] , \min_val_reg[0][28] , \min_val_reg[0][27] ,
         \min_val_reg[0][26] , \min_val_reg[0][25] , \min_val_reg[0][24] ,
         \min_val_reg[0][23] , \min_val_reg[0][22] , \min_val_reg[0][21] ,
         \min_val_reg[0][20] , \min_val_reg[0][19] , \min_val_reg[0][18] ,
         \min_val_reg[0][17] , \min_val_reg[0][16] , \min_val_reg[0][15] ,
         \min_val_reg[0][14] , \min_val_reg[0][13] , \min_val_reg[0][12] ,
         \min_val_reg[0][11] , \min_val_reg[0][10] , \min_val_reg[0][9] ,
         \min_val_reg[0][8] , \min_val_reg[0][7] , \min_val_reg[0][6] ,
         \min_val_reg[0][5] , \min_val_reg[0][4] , \min_val_reg[0][3] ,
         \min_val_reg[0][2] , \min_val_reg[0][1] , \min_val_reg[0][0] , n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952;

  DFF \min_dist_reg_reg[0][0]  ( .D(\local_min_dist[0][0] ), .CLK(clk), .RST(
        rst), .I(1'b1), .Q(\min_dist_reg[0][0] ) );
  DFF \min_dist_reg_reg[0][1]  ( .D(\local_min_dist[0][1] ), .CLK(clk), .RST(
        rst), .I(1'b1), .Q(\min_dist_reg[0][1] ) );
  DFF \min_dist_reg_reg[0][2]  ( .D(\local_min_dist[0][2] ), .CLK(clk), .RST(
        rst), .I(1'b1), .Q(\min_dist_reg[0][2] ) );
  DFF \min_dist_reg_reg[0][3]  ( .D(\local_min_dist[0][3] ), .CLK(clk), .RST(
        rst), .I(1'b1), .Q(\min_dist_reg[0][3] ) );
  DFF \min_dist_reg_reg[0][4]  ( .D(\local_min_dist[0][4] ), .CLK(clk), .RST(
        rst), .I(1'b1), .Q(\min_dist_reg[0][4] ) );
  DFF \min_dist_reg_reg[1][0]  ( .D(\min_dist[1][0] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[1][0] ) );
  DFF \min_dist_reg_reg[1][1]  ( .D(\min_dist[1][1] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[1][1] ) );
  DFF \min_dist_reg_reg[1][2]  ( .D(\min_dist[1][2] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[1][2] ) );
  DFF \min_dist_reg_reg[1][3]  ( .D(\min_dist[1][3] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[1][3] ) );
  DFF \min_dist_reg_reg[1][4]  ( .D(\min_dist[1][4] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[1][4] ) );
  DFF \min_dist_reg_reg[2][0]  ( .D(\min_dist[2][0] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[2][0] ) );
  DFF \min_dist_reg_reg[2][1]  ( .D(\min_dist[2][1] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[2][1] ) );
  DFF \min_dist_reg_reg[2][2]  ( .D(\min_dist[2][2] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[2][2] ) );
  DFF \min_dist_reg_reg[2][3]  ( .D(\min_dist[2][3] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[2][3] ) );
  DFF \min_dist_reg_reg[2][4]  ( .D(\min_dist[2][4] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[2][4] ) );
  DFF \min_dist_reg_reg[3][0]  ( .D(\min_dist[3][0] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[3][0] ) );
  DFF \min_dist_reg_reg[3][1]  ( .D(\min_dist[3][1] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[3][1] ) );
  DFF \min_dist_reg_reg[3][2]  ( .D(\min_dist[3][2] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[3][2] ) );
  DFF \min_dist_reg_reg[3][3]  ( .D(\min_dist[3][3] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[3][3] ) );
  DFF \min_dist_reg_reg[3][4]  ( .D(\min_dist[3][4] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[3][4] ) );
  DFF \min_val_reg_reg[0][0]  ( .D(o[0]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \min_val_reg[0][0] ) );
  DFF \min_val_reg_reg[0][1]  ( .D(o[1]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \min_val_reg[0][1] ) );
  DFF \min_val_reg_reg[0][2]  ( .D(o[2]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \min_val_reg[0][2] ) );
  DFF \min_val_reg_reg[0][3]  ( .D(o[3]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \min_val_reg[0][3] ) );
  DFF \min_val_reg_reg[0][4]  ( .D(o[4]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \min_val_reg[0][4] ) );
  DFF \min_val_reg_reg[0][5]  ( .D(o[5]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \min_val_reg[0][5] ) );
  DFF \min_val_reg_reg[0][6]  ( .D(o[6]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \min_val_reg[0][6] ) );
  DFF \min_val_reg_reg[0][7]  ( .D(o[7]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \min_val_reg[0][7] ) );
  DFF \min_val_reg_reg[0][8]  ( .D(o[8]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \min_val_reg[0][8] ) );
  DFF \min_val_reg_reg[0][9]  ( .D(o[9]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \min_val_reg[0][9] ) );
  DFF \min_val_reg_reg[0][10]  ( .D(o[10]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][10] ) );
  DFF \min_val_reg_reg[0][11]  ( .D(o[11]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][11] ) );
  DFF \min_val_reg_reg[0][12]  ( .D(o[12]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][12] ) );
  DFF \min_val_reg_reg[0][13]  ( .D(o[13]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][13] ) );
  DFF \min_val_reg_reg[0][14]  ( .D(o[14]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][14] ) );
  DFF \min_val_reg_reg[0][15]  ( .D(o[15]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][15] ) );
  DFF \min_val_reg_reg[0][16]  ( .D(o[16]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][16] ) );
  DFF \min_val_reg_reg[0][17]  ( .D(o[17]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][17] ) );
  DFF \min_val_reg_reg[0][18]  ( .D(o[18]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][18] ) );
  DFF \min_val_reg_reg[0][19]  ( .D(o[19]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][19] ) );
  DFF \min_val_reg_reg[0][20]  ( .D(o[20]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][20] ) );
  DFF \min_val_reg_reg[0][21]  ( .D(o[21]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][21] ) );
  DFF \min_val_reg_reg[0][22]  ( .D(o[22]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][22] ) );
  DFF \min_val_reg_reg[0][23]  ( .D(o[23]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][23] ) );
  DFF \min_val_reg_reg[0][24]  ( .D(o[24]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][24] ) );
  DFF \min_val_reg_reg[0][25]  ( .D(o[25]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][25] ) );
  DFF \min_val_reg_reg[0][26]  ( .D(o[26]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][26] ) );
  DFF \min_val_reg_reg[0][27]  ( .D(o[27]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][27] ) );
  DFF \min_val_reg_reg[0][28]  ( .D(o[28]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][28] ) );
  DFF \min_val_reg_reg[0][29]  ( .D(o[29]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][29] ) );
  DFF \min_val_reg_reg[0][30]  ( .D(o[30]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[0][30] ) );
  DFF \min_val_reg_reg[1][0]  ( .D(o[31]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \min_val_reg[1][0] ) );
  DFF \min_val_reg_reg[1][1]  ( .D(o[32]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \min_val_reg[1][1] ) );
  DFF \min_val_reg_reg[1][2]  ( .D(o[33]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \min_val_reg[1][2] ) );
  DFF \min_val_reg_reg[1][3]  ( .D(o[34]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \min_val_reg[1][3] ) );
  DFF \min_val_reg_reg[1][4]  ( .D(o[35]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \min_val_reg[1][4] ) );
  DFF \min_val_reg_reg[1][5]  ( .D(o[36]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \min_val_reg[1][5] ) );
  DFF \min_val_reg_reg[1][6]  ( .D(o[37]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \min_val_reg[1][6] ) );
  DFF \min_val_reg_reg[1][7]  ( .D(o[38]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \min_val_reg[1][7] ) );
  DFF \min_val_reg_reg[1][8]  ( .D(o[39]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \min_val_reg[1][8] ) );
  DFF \min_val_reg_reg[1][9]  ( .D(o[40]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \min_val_reg[1][9] ) );
  DFF \min_val_reg_reg[1][10]  ( .D(o[41]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][10] ) );
  DFF \min_val_reg_reg[1][11]  ( .D(o[42]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][11] ) );
  DFF \min_val_reg_reg[1][12]  ( .D(o[43]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][12] ) );
  DFF \min_val_reg_reg[1][13]  ( .D(o[44]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][13] ) );
  DFF \min_val_reg_reg[1][14]  ( .D(o[45]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][14] ) );
  DFF \min_val_reg_reg[1][15]  ( .D(o[46]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][15] ) );
  DFF \min_val_reg_reg[1][16]  ( .D(o[47]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][16] ) );
  DFF \min_val_reg_reg[1][17]  ( .D(o[48]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][17] ) );
  DFF \min_val_reg_reg[1][18]  ( .D(o[49]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][18] ) );
  DFF \min_val_reg_reg[1][19]  ( .D(o[50]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][19] ) );
  DFF \min_val_reg_reg[1][20]  ( .D(o[51]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][20] ) );
  DFF \min_val_reg_reg[1][21]  ( .D(o[52]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][21] ) );
  DFF \min_val_reg_reg[1][22]  ( .D(o[53]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][22] ) );
  DFF \min_val_reg_reg[1][23]  ( .D(o[54]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][23] ) );
  DFF \min_val_reg_reg[1][24]  ( .D(o[55]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][24] ) );
  DFF \min_val_reg_reg[1][25]  ( .D(o[56]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][25] ) );
  DFF \min_val_reg_reg[1][26]  ( .D(o[57]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][26] ) );
  DFF \min_val_reg_reg[1][27]  ( .D(o[58]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][27] ) );
  DFF \min_val_reg_reg[1][28]  ( .D(o[59]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][28] ) );
  DFF \min_val_reg_reg[1][29]  ( .D(o[60]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][29] ) );
  DFF \min_val_reg_reg[1][30]  ( .D(o[61]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[1][30] ) );
  DFF \min_val_reg_reg[2][0]  ( .D(o[62]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \min_val_reg[2][0] ) );
  DFF \min_val_reg_reg[2][1]  ( .D(o[63]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \min_val_reg[2][1] ) );
  DFF \min_val_reg_reg[2][2]  ( .D(o[64]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \min_val_reg[2][2] ) );
  DFF \min_val_reg_reg[2][3]  ( .D(o[65]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \min_val_reg[2][3] ) );
  DFF \min_val_reg_reg[2][4]  ( .D(o[66]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \min_val_reg[2][4] ) );
  DFF \min_val_reg_reg[2][5]  ( .D(o[67]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \min_val_reg[2][5] ) );
  DFF \min_val_reg_reg[2][6]  ( .D(o[68]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \min_val_reg[2][6] ) );
  DFF \min_val_reg_reg[2][7]  ( .D(o[69]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \min_val_reg[2][7] ) );
  DFF \min_val_reg_reg[2][8]  ( .D(o[70]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \min_val_reg[2][8] ) );
  DFF \min_val_reg_reg[2][9]  ( .D(o[71]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \min_val_reg[2][9] ) );
  DFF \min_val_reg_reg[2][10]  ( .D(o[72]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][10] ) );
  DFF \min_val_reg_reg[2][11]  ( .D(o[73]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][11] ) );
  DFF \min_val_reg_reg[2][12]  ( .D(o[74]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][12] ) );
  DFF \min_val_reg_reg[2][13]  ( .D(o[75]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][13] ) );
  DFF \min_val_reg_reg[2][14]  ( .D(o[76]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][14] ) );
  DFF \min_val_reg_reg[2][15]  ( .D(o[77]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][15] ) );
  DFF \min_val_reg_reg[2][16]  ( .D(o[78]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][16] ) );
  DFF \min_val_reg_reg[2][17]  ( .D(o[79]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][17] ) );
  DFF \min_val_reg_reg[2][18]  ( .D(o[80]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][18] ) );
  DFF \min_val_reg_reg[2][19]  ( .D(o[81]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][19] ) );
  DFF \min_val_reg_reg[2][20]  ( .D(o[82]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][20] ) );
  DFF \min_val_reg_reg[2][21]  ( .D(o[83]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][21] ) );
  DFF \min_val_reg_reg[2][22]  ( .D(o[84]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][22] ) );
  DFF \min_val_reg_reg[2][23]  ( .D(o[85]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][23] ) );
  DFF \min_val_reg_reg[2][24]  ( .D(o[86]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][24] ) );
  DFF \min_val_reg_reg[2][25]  ( .D(o[87]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][25] ) );
  DFF \min_val_reg_reg[2][26]  ( .D(o[88]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][26] ) );
  DFF \min_val_reg_reg[2][27]  ( .D(o[89]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][27] ) );
  DFF \min_val_reg_reg[2][28]  ( .D(o[90]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][28] ) );
  DFF \min_val_reg_reg[2][29]  ( .D(o[91]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][29] ) );
  DFF \min_val_reg_reg[2][30]  ( .D(o[92]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[2][30] ) );
  DFF \min_val_reg_reg[3][0]  ( .D(o[93]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \min_val_reg[3][0] ) );
  DFF \min_val_reg_reg[3][1]  ( .D(o[94]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \min_val_reg[3][1] ) );
  DFF \min_val_reg_reg[3][2]  ( .D(o[95]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \min_val_reg[3][2] ) );
  DFF \min_val_reg_reg[3][3]  ( .D(o[96]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \min_val_reg[3][3] ) );
  DFF \min_val_reg_reg[3][4]  ( .D(o[97]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \min_val_reg[3][4] ) );
  DFF \min_val_reg_reg[3][5]  ( .D(o[98]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \min_val_reg[3][5] ) );
  DFF \min_val_reg_reg[3][6]  ( .D(o[99]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \min_val_reg[3][6] ) );
  DFF \min_val_reg_reg[3][7]  ( .D(o[100]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][7] ) );
  DFF \min_val_reg_reg[3][8]  ( .D(o[101]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][8] ) );
  DFF \min_val_reg_reg[3][9]  ( .D(o[102]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][9] ) );
  DFF \min_val_reg_reg[3][10]  ( .D(o[103]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][10] ) );
  DFF \min_val_reg_reg[3][11]  ( .D(o[104]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][11] ) );
  DFF \min_val_reg_reg[3][12]  ( .D(o[105]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][12] ) );
  DFF \min_val_reg_reg[3][13]  ( .D(o[106]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][13] ) );
  DFF \min_val_reg_reg[3][14]  ( .D(o[107]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][14] ) );
  DFF \min_val_reg_reg[3][15]  ( .D(o[108]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][15] ) );
  DFF \min_val_reg_reg[3][16]  ( .D(o[109]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][16] ) );
  DFF \min_val_reg_reg[3][17]  ( .D(o[110]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][17] ) );
  DFF \min_val_reg_reg[3][18]  ( .D(o[111]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][18] ) );
  DFF \min_val_reg_reg[3][19]  ( .D(o[112]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][19] ) );
  DFF \min_val_reg_reg[3][20]  ( .D(o[113]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][20] ) );
  DFF \min_val_reg_reg[3][21]  ( .D(o[114]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][21] ) );
  DFF \min_val_reg_reg[3][22]  ( .D(o[115]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][22] ) );
  DFF \min_val_reg_reg[3][23]  ( .D(o[116]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][23] ) );
  DFF \min_val_reg_reg[3][24]  ( .D(o[117]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][24] ) );
  DFF \min_val_reg_reg[3][25]  ( .D(o[118]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][25] ) );
  DFF \min_val_reg_reg[3][26]  ( .D(o[119]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][26] ) );
  DFF \min_val_reg_reg[3][27]  ( .D(o[120]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][27] ) );
  DFF \min_val_reg_reg[3][28]  ( .D(o[121]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][28] ) );
  DFF \min_val_reg_reg[3][29]  ( .D(o[122]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][29] ) );
  DFF \min_val_reg_reg[3][30]  ( .D(o[123]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(\min_val_reg[3][30] ) );
  XOR U178 ( .A(\min_val_reg[0][9] ), .B(n145), .Z(o[9]) );
  AND U179 ( .A(n146), .B(n147), .Z(n145) );
  XNOR U180 ( .A(n148), .B(n149), .Z(o[99]) );
  AND U181 ( .A(n150), .B(n151), .Z(n148) );
  XNOR U182 ( .A(n152), .B(n153), .Z(o[98]) );
  AND U183 ( .A(n150), .B(n154), .Z(n152) );
  XNOR U184 ( .A(n155), .B(n156), .Z(o[97]) );
  AND U185 ( .A(n150), .B(n157), .Z(n155) );
  XNOR U186 ( .A(n158), .B(n159), .Z(o[96]) );
  AND U187 ( .A(n150), .B(n160), .Z(n158) );
  XNOR U188 ( .A(n161), .B(n162), .Z(o[95]) );
  AND U189 ( .A(n150), .B(n163), .Z(n161) );
  XNOR U190 ( .A(n164), .B(n165), .Z(o[94]) );
  AND U191 ( .A(n150), .B(n166), .Z(n164) );
  XNOR U192 ( .A(n167), .B(n168), .Z(o[93]) );
  AND U193 ( .A(n150), .B(n169), .Z(n167) );
  XOR U194 ( .A(n170), .B(n171), .Z(o[92]) );
  AND U195 ( .A(n172), .B(n173), .Z(n170) );
  XOR U196 ( .A(n174), .B(n175), .Z(o[91]) );
  AND U197 ( .A(n172), .B(n176), .Z(n174) );
  XOR U198 ( .A(n177), .B(n178), .Z(o[90]) );
  AND U199 ( .A(n172), .B(n179), .Z(n177) );
  XOR U200 ( .A(\min_val_reg[0][8] ), .B(n180), .Z(o[8]) );
  AND U201 ( .A(n146), .B(n181), .Z(n180) );
  XOR U202 ( .A(n182), .B(n183), .Z(o[89]) );
  AND U203 ( .A(n172), .B(n184), .Z(n182) );
  XOR U204 ( .A(n185), .B(n186), .Z(o[88]) );
  AND U205 ( .A(n172), .B(n187), .Z(n185) );
  XOR U206 ( .A(n188), .B(n189), .Z(o[87]) );
  AND U207 ( .A(n172), .B(n190), .Z(n188) );
  XOR U208 ( .A(n191), .B(n192), .Z(o[86]) );
  AND U209 ( .A(n172), .B(n193), .Z(n191) );
  XOR U210 ( .A(n194), .B(n195), .Z(o[85]) );
  AND U211 ( .A(n172), .B(n196), .Z(n194) );
  XOR U212 ( .A(n197), .B(n198), .Z(o[84]) );
  AND U213 ( .A(n172), .B(n199), .Z(n197) );
  XOR U214 ( .A(n200), .B(n201), .Z(o[83]) );
  AND U215 ( .A(n172), .B(n202), .Z(n200) );
  XOR U216 ( .A(n203), .B(n204), .Z(o[82]) );
  AND U217 ( .A(n172), .B(n205), .Z(n203) );
  XOR U218 ( .A(n206), .B(n207), .Z(o[81]) );
  AND U219 ( .A(n172), .B(n208), .Z(n206) );
  XOR U220 ( .A(n209), .B(n210), .Z(o[80]) );
  AND U221 ( .A(n172), .B(n211), .Z(n209) );
  XOR U222 ( .A(\min_val_reg[0][7] ), .B(n212), .Z(o[7]) );
  AND U223 ( .A(n146), .B(n213), .Z(n212) );
  XOR U224 ( .A(n214), .B(n215), .Z(o[79]) );
  AND U225 ( .A(n172), .B(n216), .Z(n214) );
  XOR U226 ( .A(n217), .B(n218), .Z(o[78]) );
  AND U227 ( .A(n172), .B(n219), .Z(n217) );
  XOR U228 ( .A(n220), .B(n221), .Z(o[77]) );
  AND U229 ( .A(n172), .B(n222), .Z(n220) );
  XOR U230 ( .A(n223), .B(n224), .Z(o[76]) );
  AND U231 ( .A(n172), .B(n225), .Z(n223) );
  XOR U232 ( .A(n226), .B(n227), .Z(o[75]) );
  AND U233 ( .A(n172), .B(n228), .Z(n226) );
  XOR U234 ( .A(n229), .B(n230), .Z(o[74]) );
  AND U235 ( .A(n172), .B(n231), .Z(n229) );
  XOR U236 ( .A(n232), .B(n233), .Z(o[73]) );
  AND U237 ( .A(n172), .B(n234), .Z(n232) );
  XOR U238 ( .A(n235), .B(n236), .Z(o[72]) );
  AND U239 ( .A(n172), .B(n237), .Z(n235) );
  XOR U240 ( .A(n238), .B(n239), .Z(o[71]) );
  AND U241 ( .A(n172), .B(n240), .Z(n238) );
  XOR U242 ( .A(n241), .B(n242), .Z(o[70]) );
  AND U243 ( .A(n172), .B(n243), .Z(n241) );
  XOR U244 ( .A(\min_val_reg[0][6] ), .B(n244), .Z(o[6]) );
  AND U245 ( .A(n146), .B(n245), .Z(n244) );
  XOR U246 ( .A(n246), .B(n247), .Z(o[69]) );
  AND U247 ( .A(n172), .B(n248), .Z(n246) );
  XNOR U248 ( .A(n249), .B(n250), .Z(o[68]) );
  AND U249 ( .A(n172), .B(n251), .Z(n249) );
  XNOR U250 ( .A(n252), .B(n253), .Z(o[67]) );
  AND U251 ( .A(n172), .B(n254), .Z(n252) );
  XNOR U252 ( .A(n255), .B(n256), .Z(o[66]) );
  AND U253 ( .A(n172), .B(n257), .Z(n255) );
  XNOR U254 ( .A(n258), .B(n259), .Z(o[65]) );
  AND U255 ( .A(n172), .B(n260), .Z(n258) );
  XNOR U256 ( .A(n261), .B(n262), .Z(o[64]) );
  AND U257 ( .A(n172), .B(n263), .Z(n261) );
  XNOR U258 ( .A(n264), .B(n265), .Z(o[63]) );
  AND U259 ( .A(n172), .B(n266), .Z(n264) );
  XNOR U260 ( .A(n267), .B(n268), .Z(o[62]) );
  AND U261 ( .A(n172), .B(n269), .Z(n267) );
  XNOR U262 ( .A(n270), .B(n271), .Z(o[61]) );
  AND U263 ( .A(n272), .B(n273), .Z(n270) );
  XNOR U264 ( .A(n274), .B(n275), .Z(o[60]) );
  AND U265 ( .A(n272), .B(n276), .Z(n274) );
  XOR U266 ( .A(\min_val_reg[0][5] ), .B(n277), .Z(o[5]) );
  AND U267 ( .A(n146), .B(n278), .Z(n277) );
  XNOR U268 ( .A(n279), .B(n280), .Z(o[59]) );
  AND U269 ( .A(n272), .B(n281), .Z(n279) );
  XNOR U270 ( .A(n282), .B(n283), .Z(o[58]) );
  AND U271 ( .A(n272), .B(n284), .Z(n282) );
  XNOR U272 ( .A(n285), .B(n286), .Z(o[57]) );
  AND U273 ( .A(n272), .B(n287), .Z(n285) );
  XNOR U274 ( .A(n288), .B(n289), .Z(o[56]) );
  AND U275 ( .A(n272), .B(n290), .Z(n288) );
  XNOR U276 ( .A(n291), .B(n292), .Z(o[55]) );
  AND U277 ( .A(n272), .B(n293), .Z(n291) );
  XNOR U278 ( .A(n294), .B(n295), .Z(o[54]) );
  AND U279 ( .A(n272), .B(n296), .Z(n294) );
  XNOR U280 ( .A(n297), .B(n298), .Z(o[53]) );
  AND U281 ( .A(n272), .B(n299), .Z(n297) );
  XNOR U282 ( .A(n300), .B(n301), .Z(o[52]) );
  AND U283 ( .A(n272), .B(n302), .Z(n300) );
  XNOR U284 ( .A(n303), .B(n304), .Z(o[51]) );
  AND U285 ( .A(n272), .B(n305), .Z(n303) );
  XNOR U286 ( .A(n306), .B(n307), .Z(o[50]) );
  AND U287 ( .A(n272), .B(n308), .Z(n306) );
  XOR U288 ( .A(\min_val_reg[0][4] ), .B(n309), .Z(o[4]) );
  AND U289 ( .A(n146), .B(n310), .Z(n309) );
  XNOR U290 ( .A(n311), .B(n312), .Z(o[49]) );
  AND U291 ( .A(n272), .B(n313), .Z(n311) );
  XNOR U292 ( .A(n314), .B(n315), .Z(o[48]) );
  AND U293 ( .A(n272), .B(n316), .Z(n314) );
  XNOR U294 ( .A(n317), .B(n318), .Z(o[47]) );
  AND U295 ( .A(n272), .B(n319), .Z(n317) );
  XNOR U296 ( .A(n320), .B(n321), .Z(o[46]) );
  AND U297 ( .A(n272), .B(n322), .Z(n320) );
  XNOR U298 ( .A(n323), .B(n324), .Z(o[45]) );
  AND U299 ( .A(n272), .B(n325), .Z(n323) );
  XNOR U300 ( .A(n326), .B(n327), .Z(o[44]) );
  AND U301 ( .A(n272), .B(n328), .Z(n326) );
  XNOR U302 ( .A(n329), .B(n330), .Z(o[43]) );
  AND U303 ( .A(n272), .B(n331), .Z(n329) );
  XNOR U304 ( .A(n332), .B(n333), .Z(o[42]) );
  AND U305 ( .A(n272), .B(n334), .Z(n332) );
  XNOR U306 ( .A(n335), .B(n336), .Z(o[41]) );
  AND U307 ( .A(n272), .B(n337), .Z(n335) );
  XOR U308 ( .A(n338), .B(n339), .Z(o[40]) );
  AND U309 ( .A(n272), .B(n147), .Z(n338) );
  XOR U310 ( .A(\min_val_reg[0][9] ), .B(n339), .Z(n147) );
  XNOR U311 ( .A(n340), .B(\min_val_reg[1][9] ), .Z(n339) );
  NAND U312 ( .A(n240), .B(n172), .Z(n340) );
  XOR U313 ( .A(\min_val_reg[1][9] ), .B(n239), .Z(n240) );
  XNOR U314 ( .A(n341), .B(\min_val_reg[2][9] ), .Z(n239) );
  NAND U315 ( .A(n342), .B(n343), .Z(n341) );
  XOR U316 ( .A(\min_val_reg[0][3] ), .B(n344), .Z(o[3]) );
  AND U317 ( .A(n146), .B(n345), .Z(n344) );
  XOR U318 ( .A(n346), .B(n347), .Z(o[39]) );
  AND U319 ( .A(n272), .B(n181), .Z(n346) );
  XOR U320 ( .A(\min_val_reg[0][8] ), .B(n347), .Z(n181) );
  XNOR U321 ( .A(n348), .B(\min_val_reg[1][8] ), .Z(n347) );
  NAND U322 ( .A(n243), .B(n172), .Z(n348) );
  XOR U323 ( .A(\min_val_reg[1][8] ), .B(n242), .Z(n243) );
  XNOR U324 ( .A(n349), .B(\min_val_reg[2][8] ), .Z(n242) );
  NAND U325 ( .A(n350), .B(n343), .Z(n349) );
  XOR U326 ( .A(n351), .B(n352), .Z(o[38]) );
  AND U327 ( .A(n272), .B(n213), .Z(n351) );
  XOR U328 ( .A(\min_val_reg[0][7] ), .B(n352), .Z(n213) );
  XNOR U329 ( .A(n353), .B(\min_val_reg[1][7] ), .Z(n352) );
  NAND U330 ( .A(n248), .B(n172), .Z(n353) );
  XOR U331 ( .A(\min_val_reg[1][7] ), .B(n247), .Z(n248) );
  XNOR U332 ( .A(n354), .B(\min_val_reg[2][7] ), .Z(n247) );
  NAND U333 ( .A(n355), .B(n343), .Z(n354) );
  XOR U334 ( .A(n356), .B(n357), .Z(o[37]) );
  AND U335 ( .A(n272), .B(n245), .Z(n356) );
  XOR U336 ( .A(\min_val_reg[0][6] ), .B(n357), .Z(n245) );
  XNOR U337 ( .A(n358), .B(\min_val_reg[1][6] ), .Z(n357) );
  NAND U338 ( .A(n251), .B(n172), .Z(n358) );
  XNOR U339 ( .A(\min_val_reg[1][6] ), .B(n250), .Z(n251) );
  XOR U340 ( .A(n359), .B(\min_val_reg[2][6] ), .Z(n250) );
  NAND U341 ( .A(n151), .B(n343), .Z(n359) );
  XNOR U342 ( .A(\min_val_reg[2][6] ), .B(n149), .Z(n151) );
  XOR U343 ( .A(n360), .B(\min_val_reg[3][6] ), .Z(n149) );
  NAND U344 ( .A(n361), .B(n362), .Z(n360) );
  XOR U345 ( .A(\min_val_reg[3][6] ), .B(e_input[6]), .Z(n361) );
  XNOR U346 ( .A(n363), .B(n364), .Z(o[36]) );
  AND U347 ( .A(n272), .B(n278), .Z(n363) );
  XNOR U348 ( .A(\min_val_reg[0][5] ), .B(n364), .Z(n278) );
  XOR U349 ( .A(n365), .B(\min_val_reg[1][5] ), .Z(n364) );
  NAND U350 ( .A(n254), .B(n172), .Z(n365) );
  XNOR U351 ( .A(\min_val_reg[1][5] ), .B(n253), .Z(n254) );
  XOR U352 ( .A(n366), .B(\min_val_reg[2][5] ), .Z(n253) );
  NAND U353 ( .A(n154), .B(n343), .Z(n366) );
  XNOR U354 ( .A(\min_val_reg[2][5] ), .B(n153), .Z(n154) );
  XOR U355 ( .A(n367), .B(\min_val_reg[3][5] ), .Z(n153) );
  NAND U356 ( .A(n368), .B(n362), .Z(n367) );
  XOR U357 ( .A(\min_val_reg[3][5] ), .B(e_input[5]), .Z(n368) );
  XNOR U358 ( .A(n369), .B(n370), .Z(o[35]) );
  AND U359 ( .A(n272), .B(n310), .Z(n369) );
  XNOR U360 ( .A(\min_val_reg[0][4] ), .B(n370), .Z(n310) );
  XOR U361 ( .A(n371), .B(\min_val_reg[1][4] ), .Z(n370) );
  NAND U362 ( .A(n257), .B(n172), .Z(n371) );
  XNOR U363 ( .A(\min_val_reg[1][4] ), .B(n256), .Z(n257) );
  XOR U364 ( .A(n372), .B(\min_val_reg[2][4] ), .Z(n256) );
  NAND U365 ( .A(n157), .B(n343), .Z(n372) );
  XNOR U366 ( .A(\min_val_reg[2][4] ), .B(n156), .Z(n157) );
  XOR U367 ( .A(n373), .B(\min_val_reg[3][4] ), .Z(n156) );
  NAND U368 ( .A(n374), .B(n362), .Z(n373) );
  XOR U369 ( .A(\min_val_reg[3][4] ), .B(e_input[4]), .Z(n374) );
  XNOR U370 ( .A(n375), .B(n376), .Z(o[34]) );
  AND U371 ( .A(n272), .B(n345), .Z(n375) );
  XNOR U372 ( .A(\min_val_reg[0][3] ), .B(n376), .Z(n345) );
  XOR U373 ( .A(n377), .B(\min_val_reg[1][3] ), .Z(n376) );
  NAND U374 ( .A(n260), .B(n172), .Z(n377) );
  XNOR U375 ( .A(\min_val_reg[1][3] ), .B(n259), .Z(n260) );
  XOR U376 ( .A(n378), .B(\min_val_reg[2][3] ), .Z(n259) );
  NAND U377 ( .A(n160), .B(n343), .Z(n378) );
  XNOR U378 ( .A(\min_val_reg[2][3] ), .B(n159), .Z(n160) );
  XOR U379 ( .A(n379), .B(\min_val_reg[3][3] ), .Z(n159) );
  NAND U380 ( .A(n380), .B(n362), .Z(n379) );
  XOR U381 ( .A(\min_val_reg[3][3] ), .B(e_input[3]), .Z(n380) );
  XNOR U382 ( .A(n381), .B(n382), .Z(o[33]) );
  AND U383 ( .A(n272), .B(n383), .Z(n381) );
  XNOR U384 ( .A(n384), .B(n385), .Z(o[32]) );
  AND U385 ( .A(n272), .B(n386), .Z(n384) );
  XNOR U386 ( .A(n387), .B(n388), .Z(o[31]) );
  AND U387 ( .A(n272), .B(n389), .Z(n387) );
  XOR U388 ( .A(\min_val_reg[0][30] ), .B(n390), .Z(o[30]) );
  AND U389 ( .A(n146), .B(n273), .Z(n390) );
  XNOR U390 ( .A(\min_val_reg[0][30] ), .B(n271), .Z(n273) );
  XOR U391 ( .A(n391), .B(\min_val_reg[1][30] ), .Z(n271) );
  NAND U392 ( .A(n173), .B(n172), .Z(n391) );
  XOR U393 ( .A(\min_val_reg[1][30] ), .B(n171), .Z(n173) );
  XNOR U394 ( .A(n392), .B(\min_val_reg[2][30] ), .Z(n171) );
  NAND U395 ( .A(n393), .B(n343), .Z(n392) );
  XOR U396 ( .A(\min_val_reg[0][2] ), .B(n394), .Z(o[2]) );
  AND U397 ( .A(n146), .B(n383), .Z(n394) );
  XNOR U398 ( .A(\min_val_reg[0][2] ), .B(n382), .Z(n383) );
  XOR U399 ( .A(n395), .B(\min_val_reg[1][2] ), .Z(n382) );
  NAND U400 ( .A(n263), .B(n172), .Z(n395) );
  XNOR U401 ( .A(\min_val_reg[1][2] ), .B(n262), .Z(n263) );
  XOR U402 ( .A(n396), .B(\min_val_reg[2][2] ), .Z(n262) );
  NAND U403 ( .A(n163), .B(n343), .Z(n396) );
  XNOR U404 ( .A(\min_val_reg[2][2] ), .B(n162), .Z(n163) );
  XOR U405 ( .A(n397), .B(\min_val_reg[3][2] ), .Z(n162) );
  NAND U406 ( .A(n398), .B(n362), .Z(n397) );
  XOR U407 ( .A(\min_val_reg[3][2] ), .B(e_input[2]), .Z(n398) );
  XOR U408 ( .A(\min_val_reg[0][29] ), .B(n399), .Z(o[29]) );
  AND U409 ( .A(n146), .B(n276), .Z(n399) );
  XNOR U410 ( .A(\min_val_reg[0][29] ), .B(n275), .Z(n276) );
  XOR U411 ( .A(n400), .B(\min_val_reg[1][29] ), .Z(n275) );
  NAND U412 ( .A(n176), .B(n172), .Z(n400) );
  XOR U413 ( .A(\min_val_reg[1][29] ), .B(n175), .Z(n176) );
  XNOR U414 ( .A(n401), .B(\min_val_reg[2][29] ), .Z(n175) );
  NAND U415 ( .A(n402), .B(n343), .Z(n401) );
  XOR U416 ( .A(\min_val_reg[0][28] ), .B(n403), .Z(o[28]) );
  AND U417 ( .A(n146), .B(n281), .Z(n403) );
  XNOR U418 ( .A(\min_val_reg[0][28] ), .B(n280), .Z(n281) );
  XOR U419 ( .A(n404), .B(\min_val_reg[1][28] ), .Z(n280) );
  NAND U420 ( .A(n179), .B(n172), .Z(n404) );
  XOR U421 ( .A(\min_val_reg[1][28] ), .B(n178), .Z(n179) );
  XNOR U422 ( .A(n405), .B(\min_val_reg[2][28] ), .Z(n178) );
  NAND U423 ( .A(n406), .B(n343), .Z(n405) );
  XOR U424 ( .A(\min_val_reg[0][27] ), .B(n407), .Z(o[27]) );
  AND U425 ( .A(n146), .B(n284), .Z(n407) );
  XNOR U426 ( .A(\min_val_reg[0][27] ), .B(n283), .Z(n284) );
  XOR U427 ( .A(n408), .B(\min_val_reg[1][27] ), .Z(n283) );
  NAND U428 ( .A(n184), .B(n172), .Z(n408) );
  XOR U429 ( .A(\min_val_reg[1][27] ), .B(n183), .Z(n184) );
  XNOR U430 ( .A(n409), .B(\min_val_reg[2][27] ), .Z(n183) );
  NAND U431 ( .A(n410), .B(n343), .Z(n409) );
  XOR U432 ( .A(\min_val_reg[0][26] ), .B(n411), .Z(o[26]) );
  AND U433 ( .A(n146), .B(n287), .Z(n411) );
  XNOR U434 ( .A(\min_val_reg[0][26] ), .B(n286), .Z(n287) );
  XOR U435 ( .A(n412), .B(\min_val_reg[1][26] ), .Z(n286) );
  NAND U436 ( .A(n187), .B(n172), .Z(n412) );
  XOR U437 ( .A(\min_val_reg[1][26] ), .B(n186), .Z(n187) );
  XNOR U438 ( .A(n413), .B(\min_val_reg[2][26] ), .Z(n186) );
  NAND U439 ( .A(n414), .B(n343), .Z(n413) );
  XOR U440 ( .A(\min_val_reg[0][25] ), .B(n415), .Z(o[25]) );
  AND U441 ( .A(n146), .B(n290), .Z(n415) );
  XNOR U442 ( .A(\min_val_reg[0][25] ), .B(n289), .Z(n290) );
  XOR U443 ( .A(n416), .B(\min_val_reg[1][25] ), .Z(n289) );
  NAND U444 ( .A(n190), .B(n172), .Z(n416) );
  XOR U445 ( .A(\min_val_reg[1][25] ), .B(n189), .Z(n190) );
  XNOR U446 ( .A(n417), .B(\min_val_reg[2][25] ), .Z(n189) );
  NAND U447 ( .A(n418), .B(n343), .Z(n417) );
  XOR U448 ( .A(\min_val_reg[0][24] ), .B(n419), .Z(o[24]) );
  AND U449 ( .A(n146), .B(n293), .Z(n419) );
  XNOR U450 ( .A(\min_val_reg[0][24] ), .B(n292), .Z(n293) );
  XOR U451 ( .A(n420), .B(\min_val_reg[1][24] ), .Z(n292) );
  NAND U452 ( .A(n193), .B(n172), .Z(n420) );
  XOR U453 ( .A(\min_val_reg[1][24] ), .B(n192), .Z(n193) );
  XNOR U454 ( .A(n421), .B(\min_val_reg[2][24] ), .Z(n192) );
  NAND U455 ( .A(n422), .B(n343), .Z(n421) );
  XOR U456 ( .A(\min_val_reg[0][23] ), .B(n423), .Z(o[23]) );
  AND U457 ( .A(n146), .B(n296), .Z(n423) );
  XNOR U458 ( .A(\min_val_reg[0][23] ), .B(n295), .Z(n296) );
  XOR U459 ( .A(n424), .B(\min_val_reg[1][23] ), .Z(n295) );
  NAND U460 ( .A(n196), .B(n172), .Z(n424) );
  XOR U461 ( .A(\min_val_reg[1][23] ), .B(n195), .Z(n196) );
  XNOR U462 ( .A(n425), .B(\min_val_reg[2][23] ), .Z(n195) );
  NAND U463 ( .A(n426), .B(n343), .Z(n425) );
  XOR U464 ( .A(\min_val_reg[0][22] ), .B(n427), .Z(o[22]) );
  AND U465 ( .A(n146), .B(n299), .Z(n427) );
  XNOR U466 ( .A(\min_val_reg[0][22] ), .B(n298), .Z(n299) );
  XOR U467 ( .A(n428), .B(\min_val_reg[1][22] ), .Z(n298) );
  NAND U468 ( .A(n199), .B(n172), .Z(n428) );
  XOR U469 ( .A(\min_val_reg[1][22] ), .B(n198), .Z(n199) );
  XNOR U470 ( .A(n429), .B(\min_val_reg[2][22] ), .Z(n198) );
  NAND U471 ( .A(n430), .B(n343), .Z(n429) );
  XOR U472 ( .A(\min_val_reg[0][21] ), .B(n431), .Z(o[21]) );
  AND U473 ( .A(n146), .B(n302), .Z(n431) );
  XNOR U474 ( .A(\min_val_reg[0][21] ), .B(n301), .Z(n302) );
  XOR U475 ( .A(n432), .B(\min_val_reg[1][21] ), .Z(n301) );
  NAND U476 ( .A(n202), .B(n172), .Z(n432) );
  XOR U477 ( .A(\min_val_reg[1][21] ), .B(n201), .Z(n202) );
  XNOR U478 ( .A(n433), .B(\min_val_reg[2][21] ), .Z(n201) );
  NAND U479 ( .A(n434), .B(n343), .Z(n433) );
  XOR U480 ( .A(\min_val_reg[0][20] ), .B(n435), .Z(o[20]) );
  AND U481 ( .A(n146), .B(n305), .Z(n435) );
  XNOR U482 ( .A(\min_val_reg[0][20] ), .B(n304), .Z(n305) );
  XOR U483 ( .A(n436), .B(\min_val_reg[1][20] ), .Z(n304) );
  NAND U484 ( .A(n205), .B(n172), .Z(n436) );
  XOR U485 ( .A(\min_val_reg[1][20] ), .B(n204), .Z(n205) );
  XNOR U486 ( .A(n437), .B(\min_val_reg[2][20] ), .Z(n204) );
  NAND U487 ( .A(n438), .B(n343), .Z(n437) );
  XOR U488 ( .A(\min_val_reg[0][1] ), .B(n439), .Z(o[1]) );
  AND U489 ( .A(n146), .B(n386), .Z(n439) );
  XNOR U490 ( .A(\min_val_reg[0][1] ), .B(n385), .Z(n386) );
  XOR U491 ( .A(n440), .B(\min_val_reg[1][1] ), .Z(n385) );
  NAND U492 ( .A(n266), .B(n172), .Z(n440) );
  XNOR U493 ( .A(\min_val_reg[1][1] ), .B(n265), .Z(n266) );
  XOR U494 ( .A(n441), .B(\min_val_reg[2][1] ), .Z(n265) );
  NAND U495 ( .A(n166), .B(n343), .Z(n441) );
  XNOR U496 ( .A(\min_val_reg[2][1] ), .B(n165), .Z(n166) );
  XOR U497 ( .A(n442), .B(\min_val_reg[3][1] ), .Z(n165) );
  NAND U498 ( .A(n443), .B(n362), .Z(n442) );
  XOR U499 ( .A(\min_val_reg[3][1] ), .B(e_input[1]), .Z(n443) );
  XOR U500 ( .A(\min_val_reg[0][19] ), .B(n444), .Z(o[19]) );
  AND U501 ( .A(n146), .B(n308), .Z(n444) );
  XNOR U502 ( .A(\min_val_reg[0][19] ), .B(n307), .Z(n308) );
  XOR U503 ( .A(n445), .B(\min_val_reg[1][19] ), .Z(n307) );
  NAND U504 ( .A(n208), .B(n172), .Z(n445) );
  XOR U505 ( .A(\min_val_reg[1][19] ), .B(n207), .Z(n208) );
  XNOR U506 ( .A(n446), .B(\min_val_reg[2][19] ), .Z(n207) );
  NAND U507 ( .A(n447), .B(n343), .Z(n446) );
  XOR U508 ( .A(\min_val_reg[0][18] ), .B(n448), .Z(o[18]) );
  AND U509 ( .A(n146), .B(n313), .Z(n448) );
  XNOR U510 ( .A(\min_val_reg[0][18] ), .B(n312), .Z(n313) );
  XOR U511 ( .A(n449), .B(\min_val_reg[1][18] ), .Z(n312) );
  NAND U512 ( .A(n211), .B(n172), .Z(n449) );
  XOR U513 ( .A(\min_val_reg[1][18] ), .B(n210), .Z(n211) );
  XNOR U514 ( .A(n450), .B(\min_val_reg[2][18] ), .Z(n210) );
  NAND U515 ( .A(n451), .B(n343), .Z(n450) );
  XOR U516 ( .A(\min_val_reg[0][17] ), .B(n452), .Z(o[17]) );
  AND U517 ( .A(n146), .B(n316), .Z(n452) );
  XNOR U518 ( .A(\min_val_reg[0][17] ), .B(n315), .Z(n316) );
  XOR U519 ( .A(n453), .B(\min_val_reg[1][17] ), .Z(n315) );
  NAND U520 ( .A(n216), .B(n172), .Z(n453) );
  XOR U521 ( .A(\min_val_reg[1][17] ), .B(n215), .Z(n216) );
  XNOR U522 ( .A(n454), .B(\min_val_reg[2][17] ), .Z(n215) );
  NAND U523 ( .A(n455), .B(n343), .Z(n454) );
  XOR U524 ( .A(\min_val_reg[0][16] ), .B(n456), .Z(o[16]) );
  AND U525 ( .A(n146), .B(n319), .Z(n456) );
  XNOR U526 ( .A(\min_val_reg[0][16] ), .B(n318), .Z(n319) );
  XOR U527 ( .A(n457), .B(\min_val_reg[1][16] ), .Z(n318) );
  NAND U528 ( .A(n219), .B(n172), .Z(n457) );
  XOR U529 ( .A(\min_val_reg[1][16] ), .B(n218), .Z(n219) );
  XNOR U530 ( .A(n458), .B(\min_val_reg[2][16] ), .Z(n218) );
  NAND U531 ( .A(n459), .B(n343), .Z(n458) );
  XOR U532 ( .A(\min_val_reg[0][15] ), .B(n460), .Z(o[15]) );
  AND U533 ( .A(n146), .B(n322), .Z(n460) );
  XNOR U534 ( .A(\min_val_reg[0][15] ), .B(n321), .Z(n322) );
  XOR U535 ( .A(n461), .B(\min_val_reg[1][15] ), .Z(n321) );
  NAND U536 ( .A(n222), .B(n172), .Z(n461) );
  XOR U537 ( .A(\min_val_reg[1][15] ), .B(n221), .Z(n222) );
  XNOR U538 ( .A(n462), .B(\min_val_reg[2][15] ), .Z(n221) );
  NAND U539 ( .A(n463), .B(n343), .Z(n462) );
  XOR U540 ( .A(\min_val_reg[0][14] ), .B(n464), .Z(o[14]) );
  AND U541 ( .A(n146), .B(n325), .Z(n464) );
  XNOR U542 ( .A(\min_val_reg[0][14] ), .B(n324), .Z(n325) );
  XOR U543 ( .A(n465), .B(\min_val_reg[1][14] ), .Z(n324) );
  NAND U544 ( .A(n225), .B(n172), .Z(n465) );
  XOR U545 ( .A(\min_val_reg[1][14] ), .B(n224), .Z(n225) );
  XNOR U546 ( .A(n466), .B(\min_val_reg[2][14] ), .Z(n224) );
  NAND U547 ( .A(n467), .B(n343), .Z(n466) );
  XOR U548 ( .A(\min_val_reg[0][13] ), .B(n468), .Z(o[13]) );
  AND U549 ( .A(n146), .B(n328), .Z(n468) );
  XNOR U550 ( .A(\min_val_reg[0][13] ), .B(n327), .Z(n328) );
  XOR U551 ( .A(n469), .B(\min_val_reg[1][13] ), .Z(n327) );
  NAND U552 ( .A(n228), .B(n172), .Z(n469) );
  XOR U553 ( .A(\min_val_reg[1][13] ), .B(n227), .Z(n228) );
  XNOR U554 ( .A(n470), .B(\min_val_reg[2][13] ), .Z(n227) );
  NAND U555 ( .A(n471), .B(n343), .Z(n470) );
  XOR U556 ( .A(\min_val_reg[0][12] ), .B(n472), .Z(o[12]) );
  AND U557 ( .A(n146), .B(n331), .Z(n472) );
  XNOR U558 ( .A(\min_val_reg[0][12] ), .B(n330), .Z(n331) );
  XOR U559 ( .A(n473), .B(\min_val_reg[1][12] ), .Z(n330) );
  NAND U560 ( .A(n231), .B(n172), .Z(n473) );
  XOR U561 ( .A(\min_val_reg[1][12] ), .B(n230), .Z(n231) );
  XNOR U562 ( .A(n474), .B(\min_val_reg[2][12] ), .Z(n230) );
  NAND U563 ( .A(n475), .B(n343), .Z(n474) );
  XNOR U564 ( .A(n476), .B(n477), .Z(o[123]) );
  AND U565 ( .A(n150), .B(n393), .Z(n476) );
  XNOR U566 ( .A(\min_val_reg[2][30] ), .B(n477), .Z(n393) );
  XOR U567 ( .A(n478), .B(\min_val_reg[3][30] ), .Z(n477) );
  NAND U568 ( .A(n479), .B(n362), .Z(n478) );
  XOR U569 ( .A(\min_val_reg[3][30] ), .B(e_input[30]), .Z(n479) );
  XNOR U570 ( .A(n480), .B(n481), .Z(o[122]) );
  AND U571 ( .A(n150), .B(n402), .Z(n480) );
  XNOR U572 ( .A(\min_val_reg[2][29] ), .B(n481), .Z(n402) );
  XOR U573 ( .A(n482), .B(\min_val_reg[3][29] ), .Z(n481) );
  NAND U574 ( .A(n483), .B(n362), .Z(n482) );
  XOR U575 ( .A(\min_val_reg[3][29] ), .B(e_input[29]), .Z(n483) );
  XNOR U576 ( .A(n484), .B(n485), .Z(o[121]) );
  AND U577 ( .A(n150), .B(n406), .Z(n484) );
  XNOR U578 ( .A(\min_val_reg[2][28] ), .B(n485), .Z(n406) );
  XOR U579 ( .A(n486), .B(\min_val_reg[3][28] ), .Z(n485) );
  NAND U580 ( .A(n487), .B(n362), .Z(n486) );
  XOR U581 ( .A(\min_val_reg[3][28] ), .B(e_input[28]), .Z(n487) );
  XNOR U582 ( .A(n488), .B(n489), .Z(o[120]) );
  AND U583 ( .A(n150), .B(n410), .Z(n488) );
  XNOR U584 ( .A(\min_val_reg[2][27] ), .B(n489), .Z(n410) );
  XOR U585 ( .A(n490), .B(\min_val_reg[3][27] ), .Z(n489) );
  NAND U586 ( .A(n491), .B(n362), .Z(n490) );
  XOR U587 ( .A(\min_val_reg[3][27] ), .B(e_input[27]), .Z(n491) );
  XOR U588 ( .A(\min_val_reg[0][11] ), .B(n492), .Z(o[11]) );
  AND U589 ( .A(n146), .B(n334), .Z(n492) );
  XNOR U590 ( .A(\min_val_reg[0][11] ), .B(n333), .Z(n334) );
  XOR U591 ( .A(n493), .B(\min_val_reg[1][11] ), .Z(n333) );
  NAND U592 ( .A(n234), .B(n172), .Z(n493) );
  XOR U593 ( .A(\min_val_reg[1][11] ), .B(n233), .Z(n234) );
  XNOR U594 ( .A(n494), .B(\min_val_reg[2][11] ), .Z(n233) );
  NAND U595 ( .A(n495), .B(n343), .Z(n494) );
  XNOR U596 ( .A(n496), .B(n497), .Z(o[119]) );
  AND U597 ( .A(n150), .B(n414), .Z(n496) );
  XNOR U598 ( .A(\min_val_reg[2][26] ), .B(n497), .Z(n414) );
  XOR U599 ( .A(n498), .B(\min_val_reg[3][26] ), .Z(n497) );
  NAND U600 ( .A(n499), .B(n362), .Z(n498) );
  XOR U601 ( .A(\min_val_reg[3][26] ), .B(e_input[26]), .Z(n499) );
  XNOR U602 ( .A(n500), .B(n501), .Z(o[118]) );
  AND U603 ( .A(n150), .B(n418), .Z(n500) );
  XNOR U604 ( .A(\min_val_reg[2][25] ), .B(n501), .Z(n418) );
  XOR U605 ( .A(n502), .B(\min_val_reg[3][25] ), .Z(n501) );
  NAND U606 ( .A(n503), .B(n362), .Z(n502) );
  XOR U607 ( .A(\min_val_reg[3][25] ), .B(e_input[25]), .Z(n503) );
  XNOR U608 ( .A(n504), .B(n505), .Z(o[117]) );
  AND U609 ( .A(n150), .B(n422), .Z(n504) );
  XNOR U610 ( .A(\min_val_reg[2][24] ), .B(n505), .Z(n422) );
  XOR U611 ( .A(n506), .B(\min_val_reg[3][24] ), .Z(n505) );
  NAND U612 ( .A(n507), .B(n362), .Z(n506) );
  XOR U613 ( .A(\min_val_reg[3][24] ), .B(e_input[24]), .Z(n507) );
  XNOR U614 ( .A(n508), .B(n509), .Z(o[116]) );
  AND U615 ( .A(n150), .B(n426), .Z(n508) );
  XNOR U616 ( .A(\min_val_reg[2][23] ), .B(n509), .Z(n426) );
  XOR U617 ( .A(n510), .B(\min_val_reg[3][23] ), .Z(n509) );
  NAND U618 ( .A(n511), .B(n362), .Z(n510) );
  XOR U619 ( .A(\min_val_reg[3][23] ), .B(e_input[23]), .Z(n511) );
  XNOR U620 ( .A(n512), .B(n513), .Z(o[115]) );
  AND U621 ( .A(n150), .B(n430), .Z(n512) );
  XNOR U622 ( .A(\min_val_reg[2][22] ), .B(n513), .Z(n430) );
  XOR U623 ( .A(n514), .B(\min_val_reg[3][22] ), .Z(n513) );
  NAND U624 ( .A(n515), .B(n362), .Z(n514) );
  XOR U625 ( .A(\min_val_reg[3][22] ), .B(e_input[22]), .Z(n515) );
  XNOR U626 ( .A(n516), .B(n517), .Z(o[114]) );
  AND U627 ( .A(n150), .B(n434), .Z(n516) );
  XNOR U628 ( .A(\min_val_reg[2][21] ), .B(n517), .Z(n434) );
  XOR U629 ( .A(n518), .B(\min_val_reg[3][21] ), .Z(n517) );
  NAND U630 ( .A(n519), .B(n362), .Z(n518) );
  XOR U631 ( .A(\min_val_reg[3][21] ), .B(e_input[21]), .Z(n519) );
  XNOR U632 ( .A(n520), .B(n521), .Z(o[113]) );
  AND U633 ( .A(n150), .B(n438), .Z(n520) );
  XNOR U634 ( .A(\min_val_reg[2][20] ), .B(n521), .Z(n438) );
  XOR U635 ( .A(n522), .B(\min_val_reg[3][20] ), .Z(n521) );
  NAND U636 ( .A(n523), .B(n362), .Z(n522) );
  XOR U637 ( .A(\min_val_reg[3][20] ), .B(e_input[20]), .Z(n523) );
  XNOR U638 ( .A(n524), .B(n525), .Z(o[112]) );
  AND U639 ( .A(n150), .B(n447), .Z(n524) );
  XNOR U640 ( .A(\min_val_reg[2][19] ), .B(n525), .Z(n447) );
  XOR U641 ( .A(n526), .B(\min_val_reg[3][19] ), .Z(n525) );
  NAND U642 ( .A(n527), .B(n362), .Z(n526) );
  XOR U643 ( .A(\min_val_reg[3][19] ), .B(e_input[19]), .Z(n527) );
  XNOR U644 ( .A(n528), .B(n529), .Z(o[111]) );
  AND U645 ( .A(n150), .B(n451), .Z(n528) );
  XNOR U646 ( .A(\min_val_reg[2][18] ), .B(n529), .Z(n451) );
  XOR U647 ( .A(n530), .B(\min_val_reg[3][18] ), .Z(n529) );
  NAND U648 ( .A(n531), .B(n362), .Z(n530) );
  XOR U649 ( .A(\min_val_reg[3][18] ), .B(e_input[18]), .Z(n531) );
  XNOR U650 ( .A(n532), .B(n533), .Z(o[110]) );
  AND U651 ( .A(n150), .B(n455), .Z(n532) );
  XNOR U652 ( .A(\min_val_reg[2][17] ), .B(n533), .Z(n455) );
  XOR U653 ( .A(n534), .B(\min_val_reg[3][17] ), .Z(n533) );
  NAND U654 ( .A(n535), .B(n362), .Z(n534) );
  XOR U655 ( .A(\min_val_reg[3][17] ), .B(e_input[17]), .Z(n535) );
  XOR U656 ( .A(\min_val_reg[0][10] ), .B(n536), .Z(o[10]) );
  AND U657 ( .A(n146), .B(n337), .Z(n536) );
  XNOR U658 ( .A(\min_val_reg[0][10] ), .B(n336), .Z(n337) );
  XOR U659 ( .A(n537), .B(\min_val_reg[1][10] ), .Z(n336) );
  NAND U660 ( .A(n237), .B(n172), .Z(n537) );
  XOR U661 ( .A(\min_val_reg[1][10] ), .B(n236), .Z(n237) );
  XNOR U662 ( .A(n538), .B(\min_val_reg[2][10] ), .Z(n236) );
  NAND U663 ( .A(n539), .B(n343), .Z(n538) );
  XNOR U664 ( .A(n540), .B(n541), .Z(o[109]) );
  AND U665 ( .A(n150), .B(n459), .Z(n540) );
  XNOR U666 ( .A(\min_val_reg[2][16] ), .B(n541), .Z(n459) );
  XOR U667 ( .A(n542), .B(\min_val_reg[3][16] ), .Z(n541) );
  NAND U668 ( .A(n543), .B(n362), .Z(n542) );
  XOR U669 ( .A(\min_val_reg[3][16] ), .B(e_input[16]), .Z(n543) );
  XNOR U670 ( .A(n544), .B(n545), .Z(o[108]) );
  AND U671 ( .A(n150), .B(n463), .Z(n544) );
  XNOR U672 ( .A(\min_val_reg[2][15] ), .B(n545), .Z(n463) );
  XOR U673 ( .A(n546), .B(\min_val_reg[3][15] ), .Z(n545) );
  NAND U674 ( .A(n547), .B(n362), .Z(n546) );
  XOR U675 ( .A(\min_val_reg[3][15] ), .B(e_input[15]), .Z(n547) );
  XNOR U676 ( .A(n548), .B(n549), .Z(o[107]) );
  AND U677 ( .A(n150), .B(n467), .Z(n548) );
  XNOR U678 ( .A(\min_val_reg[2][14] ), .B(n549), .Z(n467) );
  XOR U679 ( .A(n550), .B(\min_val_reg[3][14] ), .Z(n549) );
  NAND U680 ( .A(n551), .B(n362), .Z(n550) );
  XOR U681 ( .A(\min_val_reg[3][14] ), .B(e_input[14]), .Z(n551) );
  XNOR U682 ( .A(n552), .B(n553), .Z(o[106]) );
  AND U683 ( .A(n150), .B(n471), .Z(n552) );
  XNOR U684 ( .A(\min_val_reg[2][13] ), .B(n553), .Z(n471) );
  XOR U685 ( .A(n554), .B(\min_val_reg[3][13] ), .Z(n553) );
  NAND U686 ( .A(n555), .B(n362), .Z(n554) );
  XOR U687 ( .A(\min_val_reg[3][13] ), .B(e_input[13]), .Z(n555) );
  XNOR U688 ( .A(n556), .B(n557), .Z(o[105]) );
  AND U689 ( .A(n150), .B(n475), .Z(n556) );
  XNOR U690 ( .A(\min_val_reg[2][12] ), .B(n557), .Z(n475) );
  XOR U691 ( .A(n558), .B(\min_val_reg[3][12] ), .Z(n557) );
  NAND U692 ( .A(n559), .B(n362), .Z(n558) );
  XOR U693 ( .A(\min_val_reg[3][12] ), .B(e_input[12]), .Z(n559) );
  XNOR U694 ( .A(n560), .B(n561), .Z(o[104]) );
  AND U695 ( .A(n150), .B(n495), .Z(n560) );
  XNOR U696 ( .A(\min_val_reg[2][11] ), .B(n561), .Z(n495) );
  XOR U697 ( .A(n562), .B(\min_val_reg[3][11] ), .Z(n561) );
  NAND U698 ( .A(n563), .B(n362), .Z(n562) );
  XOR U699 ( .A(\min_val_reg[3][11] ), .B(e_input[11]), .Z(n563) );
  XNOR U700 ( .A(n564), .B(n565), .Z(o[103]) );
  AND U701 ( .A(n150), .B(n539), .Z(n564) );
  XNOR U702 ( .A(\min_val_reg[2][10] ), .B(n565), .Z(n539) );
  XOR U703 ( .A(n566), .B(\min_val_reg[3][10] ), .Z(n565) );
  NAND U704 ( .A(n567), .B(n362), .Z(n566) );
  XOR U705 ( .A(\min_val_reg[3][10] ), .B(e_input[10]), .Z(n567) );
  XNOR U706 ( .A(n568), .B(n569), .Z(o[102]) );
  AND U707 ( .A(n150), .B(n342), .Z(n568) );
  XNOR U708 ( .A(\min_val_reg[2][9] ), .B(n569), .Z(n342) );
  XOR U709 ( .A(n570), .B(\min_val_reg[3][9] ), .Z(n569) );
  NAND U710 ( .A(n571), .B(n362), .Z(n570) );
  XOR U711 ( .A(\min_val_reg[3][9] ), .B(e_input[9]), .Z(n571) );
  XNOR U712 ( .A(n572), .B(n573), .Z(o[101]) );
  AND U713 ( .A(n150), .B(n350), .Z(n572) );
  XNOR U714 ( .A(\min_val_reg[2][8] ), .B(n573), .Z(n350) );
  XOR U715 ( .A(n574), .B(\min_val_reg[3][8] ), .Z(n573) );
  NAND U716 ( .A(n575), .B(n362), .Z(n574) );
  XOR U717 ( .A(\min_val_reg[3][8] ), .B(e_input[8]), .Z(n575) );
  XNOR U718 ( .A(n576), .B(n577), .Z(o[100]) );
  AND U719 ( .A(n150), .B(n355), .Z(n576) );
  XNOR U720 ( .A(\min_val_reg[2][7] ), .B(n577), .Z(n355) );
  XOR U721 ( .A(n578), .B(\min_val_reg[3][7] ), .Z(n577) );
  NAND U722 ( .A(n579), .B(n362), .Z(n578) );
  XOR U723 ( .A(\min_val_reg[3][7] ), .B(e_input[7]), .Z(n579) );
  XOR U724 ( .A(\min_val_reg[0][0] ), .B(n580), .Z(o[0]) );
  AND U725 ( .A(n146), .B(n389), .Z(n580) );
  XNOR U726 ( .A(\min_val_reg[0][0] ), .B(n388), .Z(n389) );
  XOR U727 ( .A(n581), .B(\min_val_reg[1][0] ), .Z(n388) );
  NAND U728 ( .A(n269), .B(n172), .Z(n581) );
  XNOR U729 ( .A(\min_val_reg[1][0] ), .B(n268), .Z(n269) );
  XOR U730 ( .A(n582), .B(\min_val_reg[2][0] ), .Z(n268) );
  NAND U731 ( .A(n169), .B(n343), .Z(n582) );
  XNOR U732 ( .A(\min_val_reg[2][0] ), .B(n168), .Z(n169) );
  XOR U733 ( .A(n583), .B(\min_val_reg[3][0] ), .Z(n168) );
  NAND U734 ( .A(n584), .B(n362), .Z(n583) );
  XOR U735 ( .A(\min_val_reg[3][0] ), .B(e_input[0]), .Z(n584) );
  XOR U736 ( .A(n585), .B(n586), .Z(\min_dist[3][4] ) );
  AND U737 ( .A(n150), .B(n587), .Z(n585) );
  XOR U738 ( .A(\min_dist_reg[2][4] ), .B(n586), .Z(n587) );
  XOR U739 ( .A(n588), .B(n589), .Z(\min_dist[3][3] ) );
  AND U740 ( .A(n150), .B(n590), .Z(n588) );
  XOR U741 ( .A(n591), .B(n592), .Z(\min_dist[3][2] ) );
  AND U742 ( .A(n150), .B(n593), .Z(n591) );
  XNOR U743 ( .A(\min_dist_reg[2][2] ), .B(n594), .Z(n593) );
  XOR U744 ( .A(n595), .B(n596), .Z(\min_dist[3][1] ) );
  AND U745 ( .A(n150), .B(n597), .Z(n595) );
  XNOR U746 ( .A(\min_dist_reg[2][1] ), .B(n598), .Z(n597) );
  XOR U747 ( .A(n599), .B(n600), .Z(\min_dist[3][0] ) );
  AND U748 ( .A(n150), .B(n601), .Z(n599) );
  XNOR U749 ( .A(n602), .B(n603), .Z(n150) );
  AND U750 ( .A(n604), .B(n605), .Z(n603) );
  XNOR U751 ( .A(n586), .B(n606), .Z(n605) );
  XNOR U752 ( .A(n602), .B(\min_dist_reg[2][4] ), .Z(n604) );
  IV U753 ( .A(n606), .Z(n602) );
  XOR U754 ( .A(n607), .B(n608), .Z(n606) );
  AND U755 ( .A(n609), .B(n610), .Z(n608) );
  XNOR U756 ( .A(n611), .B(n612), .Z(n610) );
  XOR U757 ( .A(n613), .B(n614), .Z(\min_dist[2][4] ) );
  AND U758 ( .A(n172), .B(n615), .Z(n613) );
  XOR U759 ( .A(\min_dist_reg[1][4] ), .B(n614), .Z(n615) );
  XOR U760 ( .A(n616), .B(n617), .Z(\min_dist[2][3] ) );
  AND U761 ( .A(n172), .B(n618), .Z(n616) );
  XOR U762 ( .A(n619), .B(n620), .Z(\min_dist[2][2] ) );
  AND U763 ( .A(n172), .B(n621), .Z(n619) );
  XOR U764 ( .A(\min_dist_reg[1][2] ), .B(n620), .Z(n621) );
  XOR U765 ( .A(n622), .B(n623), .Z(\min_dist[2][1] ) );
  AND U766 ( .A(n172), .B(n624), .Z(n622) );
  XOR U767 ( .A(\min_dist_reg[1][1] ), .B(n623), .Z(n624) );
  XOR U768 ( .A(n625), .B(n626), .Z(\min_dist[2][0] ) );
  AND U769 ( .A(n172), .B(n627), .Z(n625) );
  XOR U770 ( .A(n628), .B(n629), .Z(\min_dist[1][4] ) );
  AND U771 ( .A(n272), .B(n630), .Z(n628) );
  XNOR U772 ( .A(\min_dist_reg[0][4] ), .B(n631), .Z(n630) );
  XOR U773 ( .A(n632), .B(n633), .Z(\min_dist[1][3] ) );
  AND U774 ( .A(n272), .B(n634), .Z(n632) );
  XOR U775 ( .A(n635), .B(n636), .Z(\min_dist[1][2] ) );
  AND U776 ( .A(n272), .B(n637), .Z(n635) );
  XOR U777 ( .A(n638), .B(n639), .Z(\min_dist[1][1] ) );
  AND U778 ( .A(n272), .B(n640), .Z(n638) );
  XNOR U779 ( .A(n641), .B(n642), .Z(\min_dist[1][0] ) );
  AND U780 ( .A(n272), .B(n643), .Z(n641) );
  XNOR U781 ( .A(\min_dist_reg[0][0] ), .B(n642), .Z(n643) );
  XNOR U782 ( .A(n644), .B(n645), .Z(n272) );
  AND U783 ( .A(n646), .B(n647), .Z(n645) );
  XNOR U784 ( .A(n631), .B(n644), .Z(n647) );
  XNOR U785 ( .A(n644), .B(\min_dist_reg[0][4] ), .Z(n646) );
  XOR U786 ( .A(n648), .B(n649), .Z(n644) );
  AND U787 ( .A(n650), .B(n651), .Z(n649) );
  XNOR U788 ( .A(n633), .B(n652), .Z(n651) );
  XNOR U789 ( .A(n648), .B(\min_dist_reg[0][3] ), .Z(n650) );
  IV U790 ( .A(n652), .Z(n648) );
  XOR U791 ( .A(n653), .B(n654), .Z(n652) );
  AND U792 ( .A(n655), .B(n656), .Z(n654) );
  XNOR U793 ( .A(n636), .B(n653), .Z(n656) );
  XOR U794 ( .A(n653), .B(\min_dist_reg[0][2] ), .Z(n655) );
  XOR U795 ( .A(n657), .B(n658), .Z(n653) );
  NAND U796 ( .A(n659), .B(n660), .Z(n657) );
  XOR U797 ( .A(n658), .B(n639), .Z(n660) );
  XNOR U798 ( .A(n658), .B(\min_dist_reg[0][1] ), .Z(n659) );
  NOR U799 ( .A(n642), .B(\min_dist_reg[0][0] ), .Z(n658) );
  AND U800 ( .A(\min_dist_reg[0][4] ), .B(n661), .Z(\local_min_dist[0][4] ) );
  NANDN U801 ( .B(n629), .A(n146), .Z(n661) );
  XOR U802 ( .A(\min_dist_reg[0][3] ), .B(n662), .Z(\local_min_dist[0][3] ) );
  AND U803 ( .A(n146), .B(n634), .Z(n662) );
  XOR U804 ( .A(\min_dist_reg[0][3] ), .B(n633), .Z(n634) );
  XOR U805 ( .A(\min_dist_reg[0][2] ), .B(n663), .Z(\local_min_dist[0][2] ) );
  AND U806 ( .A(n146), .B(n637), .Z(n663) );
  XOR U807 ( .A(\min_dist_reg[0][2] ), .B(n636), .Z(n637) );
  XOR U808 ( .A(\min_dist_reg[0][1] ), .B(n664), .Z(\local_min_dist[0][1] ) );
  AND U809 ( .A(n146), .B(n640), .Z(n664) );
  XOR U810 ( .A(\min_dist_reg[0][1] ), .B(n639), .Z(n640) );
  XOR U811 ( .A(\min_dist_reg[0][0] ), .B(n665), .Z(\local_min_dist[0][0] ) );
  AND U812 ( .A(n146), .B(n666), .Z(n665) );
  XOR U813 ( .A(\min_dist_reg[0][0] ), .B(n667), .Z(n666) );
  XNOR U814 ( .A(n668), .B(n669), .Z(n146) );
  AND U815 ( .A(n670), .B(n671), .Z(n669) );
  XNOR U816 ( .A(n631), .B(n668), .Z(n671) );
  IV U817 ( .A(n629), .Z(n631) );
  AND U818 ( .A(n672), .B(\min_dist_reg[1][4] ), .Z(n629) );
  NANDN U819 ( .B(n614), .A(n172), .Z(n672) );
  XNOR U820 ( .A(n668), .B(\min_dist_reg[0][4] ), .Z(n670) );
  XOR U821 ( .A(n673), .B(n674), .Z(n668) );
  AND U822 ( .A(n675), .B(n676), .Z(n674) );
  XNOR U823 ( .A(n677), .B(n633), .Z(n676) );
  XNOR U824 ( .A(n678), .B(\min_dist_reg[1][3] ), .Z(n633) );
  NAND U825 ( .A(n618), .B(n172), .Z(n678) );
  XOR U826 ( .A(\min_dist_reg[1][3] ), .B(n617), .Z(n618) );
  XNOR U827 ( .A(n673), .B(\min_dist_reg[0][3] ), .Z(n675) );
  IV U828 ( .A(n677), .Z(n673) );
  XOR U829 ( .A(n679), .B(n680), .Z(n677) );
  AND U830 ( .A(n681), .B(n682), .Z(n680) );
  XNOR U831 ( .A(n679), .B(n636), .Z(n682) );
  XNOR U832 ( .A(n683), .B(\min_dist_reg[1][2] ), .Z(n636) );
  NAND U833 ( .A(n684), .B(n172), .Z(n683) );
  XNOR U834 ( .A(n685), .B(n620), .Z(n684) );
  XOR U835 ( .A(n679), .B(\min_dist_reg[0][2] ), .Z(n681) );
  XOR U836 ( .A(n686), .B(n687), .Z(n679) );
  NAND U837 ( .A(n688), .B(n689), .Z(n686) );
  XOR U838 ( .A(n687), .B(n639), .Z(n689) );
  XNOR U839 ( .A(n690), .B(\min_dist_reg[1][1] ), .Z(n639) );
  NAND U840 ( .A(n691), .B(n172), .Z(n690) );
  XNOR U841 ( .A(n692), .B(n623), .Z(n691) );
  XNOR U842 ( .A(n687), .B(\min_dist_reg[0][1] ), .Z(n688) );
  ANDN U843 ( .A(n667), .B(\min_dist_reg[0][0] ), .Z(n687) );
  IV U844 ( .A(n642), .Z(n667) );
  XOR U845 ( .A(n693), .B(\min_dist_reg[1][0] ), .Z(n642) );
  NAND U846 ( .A(n627), .B(n172), .Z(n693) );
  XNOR U847 ( .A(n694), .B(n695), .Z(n172) );
  AND U848 ( .A(n696), .B(n697), .Z(n695) );
  XNOR U849 ( .A(n614), .B(n698), .Z(n697) );
  AND U850 ( .A(n699), .B(\min_dist_reg[2][4] ), .Z(n614) );
  NANDN U851 ( .B(n586), .A(n343), .Z(n699) );
  XNOR U852 ( .A(n694), .B(\min_dist_reg[1][4] ), .Z(n696) );
  IV U853 ( .A(n698), .Z(n694) );
  XOR U854 ( .A(n700), .B(n701), .Z(n698) );
  AND U855 ( .A(n702), .B(n703), .Z(n701) );
  XNOR U856 ( .A(n617), .B(n700), .Z(n703) );
  XNOR U857 ( .A(n704), .B(\min_dist_reg[2][3] ), .Z(n617) );
  NAND U858 ( .A(n590), .B(n343), .Z(n704) );
  XNOR U859 ( .A(\min_dist_reg[2][3] ), .B(n611), .Z(n590) );
  IV U860 ( .A(n589), .Z(n611) );
  XNOR U861 ( .A(n705), .B(\min_dist_reg[1][3] ), .Z(n702) );
  IV U862 ( .A(n700), .Z(n705) );
  XOR U863 ( .A(n706), .B(n707), .Z(n700) );
  AND U864 ( .A(n708), .B(n709), .Z(n707) );
  XNOR U865 ( .A(n620), .B(n706), .Z(n709) );
  XNOR U866 ( .A(n710), .B(\min_dist_reg[2][2] ), .Z(n620) );
  NAND U867 ( .A(n711), .B(n343), .Z(n710) );
  XNOR U868 ( .A(n712), .B(n592), .Z(n711) );
  XNOR U869 ( .A(n706), .B(n685), .Z(n708) );
  IV U870 ( .A(\min_dist_reg[1][2] ), .Z(n685) );
  XOR U871 ( .A(n713), .B(n714), .Z(n706) );
  NAND U872 ( .A(n715), .B(n716), .Z(n713) );
  XOR U873 ( .A(n714), .B(n623), .Z(n716) );
  XNOR U874 ( .A(n717), .B(\min_dist_reg[2][1] ), .Z(n623) );
  NAND U875 ( .A(n718), .B(n343), .Z(n717) );
  XNOR U876 ( .A(n719), .B(n596), .Z(n718) );
  XOR U877 ( .A(n714), .B(n692), .Z(n715) );
  IV U878 ( .A(\min_dist_reg[1][1] ), .Z(n692) );
  AND U879 ( .A(n626), .B(n720), .Z(n714) );
  XNOR U880 ( .A(n720), .B(n626), .Z(n627) );
  XNOR U881 ( .A(n721), .B(\min_dist_reg[2][0] ), .Z(n626) );
  NAND U882 ( .A(n601), .B(n343), .Z(n721) );
  XNOR U883 ( .A(n722), .B(n723), .Z(n343) );
  AND U884 ( .A(n724), .B(n725), .Z(n723) );
  XNOR U885 ( .A(n726), .B(n586), .Z(n725) );
  XNOR U886 ( .A(n727), .B(\min_dist_reg[3][4] ), .Z(n586) );
  NAND U887 ( .A(n728), .B(n362), .Z(n727) );
  XOR U888 ( .A(\min_dist_reg[3][4] ), .B(n729), .Z(n728) );
  XNOR U889 ( .A(n722), .B(\min_dist_reg[2][4] ), .Z(n724) );
  IV U890 ( .A(n726), .Z(n722) );
  XOR U891 ( .A(n607), .B(n730), .Z(n726) );
  AND U892 ( .A(n609), .B(n731), .Z(n730) );
  XNOR U893 ( .A(n607), .B(n589), .Z(n731) );
  XNOR U894 ( .A(n732), .B(\min_dist_reg[3][3] ), .Z(n589) );
  NAND U895 ( .A(n733), .B(n362), .Z(n732) );
  XNOR U896 ( .A(\min_dist_reg[3][3] ), .B(n734), .Z(n733) );
  XNOR U897 ( .A(n612), .B(\min_dist_reg[2][3] ), .Z(n609) );
  IV U898 ( .A(n607), .Z(n612) );
  XOR U899 ( .A(n735), .B(n736), .Z(n607) );
  AND U900 ( .A(n737), .B(n738), .Z(n736) );
  XOR U901 ( .A(n594), .B(n735), .Z(n738) );
  IV U902 ( .A(n592), .Z(n594) );
  XNOR U903 ( .A(n739), .B(\min_dist_reg[3][2] ), .Z(n592) );
  NAND U904 ( .A(n740), .B(n362), .Z(n739) );
  XNOR U905 ( .A(\min_dist_reg[3][2] ), .B(n741), .Z(n740) );
  XNOR U906 ( .A(n735), .B(n712), .Z(n737) );
  IV U907 ( .A(\min_dist_reg[2][2] ), .Z(n712) );
  XOR U908 ( .A(n742), .B(n743), .Z(n735) );
  NAND U909 ( .A(n744), .B(n745), .Z(n742) );
  XNOR U910 ( .A(n743), .B(n598), .Z(n745) );
  IV U911 ( .A(n596), .Z(n598) );
  XNOR U912 ( .A(n746), .B(\min_dist_reg[3][1] ), .Z(n596) );
  NAND U913 ( .A(n747), .B(n362), .Z(n746) );
  XNOR U914 ( .A(\min_dist_reg[3][1] ), .B(n748), .Z(n747) );
  XOR U915 ( .A(n743), .B(n719), .Z(n744) );
  IV U916 ( .A(\min_dist_reg[2][1] ), .Z(n719) );
  ANDN U917 ( .A(n600), .B(\min_dist_reg[2][0] ), .Z(n743) );
  XOR U918 ( .A(\min_dist_reg[2][0] ), .B(n600), .Z(n601) );
  XOR U919 ( .A(n749), .B(n750), .Z(n600) );
  NAND U920 ( .A(n751), .B(n362), .Z(n749) );
  XNOR U921 ( .A(n752), .B(n753), .Z(n362) );
  AND U922 ( .A(n754), .B(n755), .Z(n753) );
  XNOR U923 ( .A(n756), .B(n729), .Z(n755) );
  XNOR U924 ( .A(n757), .B(n758), .Z(n729) );
  ANDN U925 ( .A(n759), .B(n760), .Z(n758) );
  XOR U926 ( .A(n757), .B(n761), .Z(n759) );
  XNOR U927 ( .A(n752), .B(\min_dist_reg[3][4] ), .Z(n754) );
  IV U928 ( .A(n756), .Z(n752) );
  XOR U929 ( .A(n762), .B(n763), .Z(n756) );
  AND U930 ( .A(n764), .B(n765), .Z(n763) );
  XOR U931 ( .A(n762), .B(n734), .Z(n765) );
  XOR U932 ( .A(n761), .B(n766), .Z(n734) );
  IV U933 ( .A(n760), .Z(n766) );
  XOR U934 ( .A(n767), .B(n768), .Z(n760) );
  IV U935 ( .A(n757), .Z(n768) );
  XNOR U936 ( .A(n769), .B(n770), .Z(n757) );
  ANDN U937 ( .A(n771), .B(n772), .Z(n770) );
  XNOR U938 ( .A(n769), .B(n773), .Z(n771) );
  XNOR U939 ( .A(n774), .B(n775), .Z(n767) );
  AND U940 ( .A(n776), .B(n777), .Z(n775) );
  XOR U941 ( .A(n778), .B(n779), .Z(n777) );
  XNOR U942 ( .A(n780), .B(n781), .Z(n761) );
  ANDN U943 ( .A(n782), .B(n783), .Z(n781) );
  XOR U944 ( .A(n784), .B(n785), .Z(n782) );
  XNOR U945 ( .A(n786), .B(\min_dist_reg[3][3] ), .Z(n764) );
  IV U946 ( .A(n762), .Z(n786) );
  XOR U947 ( .A(n787), .B(n788), .Z(n762) );
  AND U948 ( .A(n789), .B(n790), .Z(n788) );
  XOR U949 ( .A(n787), .B(n741), .Z(n790) );
  XOR U950 ( .A(n773), .B(n791), .Z(n741) );
  IV U951 ( .A(n772), .Z(n791) );
  XNOR U952 ( .A(n792), .B(n779), .Z(n772) );
  XNOR U953 ( .A(n793), .B(n794), .Z(n779) );
  ANDN U954 ( .A(n795), .B(n796), .Z(n794) );
  XOR U955 ( .A(n797), .B(n798), .Z(n795) );
  XNOR U956 ( .A(n776), .B(n769), .Z(n792) );
  XOR U957 ( .A(n799), .B(n800), .Z(n769) );
  ANDN U958 ( .A(n801), .B(n802), .Z(n800) );
  XNOR U959 ( .A(n799), .B(n803), .Z(n801) );
  XNOR U960 ( .A(n804), .B(n774), .Z(n776) );
  IV U961 ( .A(n778), .Z(n774) );
  XNOR U962 ( .A(n805), .B(n806), .Z(n778) );
  AND U963 ( .A(n807), .B(n808), .Z(n806) );
  XNOR U964 ( .A(n805), .B(n809), .Z(n808) );
  XNOR U965 ( .A(n810), .B(n811), .Z(n804) );
  AND U966 ( .A(n812), .B(n813), .Z(n811) );
  XOR U967 ( .A(n814), .B(n815), .Z(n813) );
  XOR U968 ( .A(n785), .B(n816), .Z(n773) );
  IV U969 ( .A(n783), .Z(n816) );
  XOR U970 ( .A(n817), .B(n780), .Z(n783) );
  IV U971 ( .A(n784), .Z(n780) );
  XNOR U972 ( .A(n818), .B(n819), .Z(n784) );
  ANDN U973 ( .A(n820), .B(n821), .Z(n819) );
  XNOR U974 ( .A(n818), .B(n822), .Z(n820) );
  XNOR U975 ( .A(n823), .B(n824), .Z(n817) );
  AND U976 ( .A(n825), .B(n826), .Z(n824) );
  XOR U977 ( .A(n827), .B(n828), .Z(n826) );
  XNOR U978 ( .A(n829), .B(n830), .Z(n785) );
  ANDN U979 ( .A(n831), .B(n832), .Z(n830) );
  XOR U980 ( .A(n833), .B(n834), .Z(n831) );
  XOR U981 ( .A(n787), .B(\min_dist_reg[3][2] ), .Z(n789) );
  XOR U982 ( .A(n835), .B(n836), .Z(n787) );
  NAND U983 ( .A(n837), .B(n838), .Z(n835) );
  XNOR U984 ( .A(n836), .B(n748), .Z(n838) );
  XOR U985 ( .A(n803), .B(n839), .Z(n748) );
  IV U986 ( .A(n802), .Z(n839) );
  XNOR U987 ( .A(n840), .B(n809), .Z(n802) );
  XOR U988 ( .A(n798), .B(n841), .Z(n809) );
  IV U989 ( .A(n796), .Z(n841) );
  XOR U990 ( .A(n842), .B(n793), .Z(n796) );
  IV U991 ( .A(n797), .Z(n793) );
  XNOR U992 ( .A(n843), .B(n844), .Z(n797) );
  ANDN U993 ( .A(n845), .B(n846), .Z(n844) );
  XNOR U994 ( .A(n843), .B(n847), .Z(n845) );
  XNOR U995 ( .A(n848), .B(n849), .Z(n842) );
  AND U996 ( .A(n850), .B(n851), .Z(n849) );
  XOR U997 ( .A(n852), .B(n853), .Z(n851) );
  IV U998 ( .A(n848), .Z(n852) );
  XNOR U999 ( .A(n854), .B(n855), .Z(n798) );
  ANDN U1000 ( .A(n856), .B(n857), .Z(n855) );
  XNOR U1001 ( .A(n854), .B(n858), .Z(n856) );
  XNOR U1002 ( .A(n807), .B(n799), .Z(n840) );
  XOR U1003 ( .A(n859), .B(n860), .Z(n799) );
  ANDN U1004 ( .A(n861), .B(n862), .Z(n860) );
  XNOR U1005 ( .A(n859), .B(n863), .Z(n861) );
  XOR U1006 ( .A(n864), .B(n815), .Z(n807) );
  XNOR U1007 ( .A(n865), .B(n866), .Z(n815) );
  ANDN U1008 ( .A(n867), .B(n868), .Z(n866) );
  XNOR U1009 ( .A(n865), .B(n869), .Z(n867) );
  XNOR U1010 ( .A(n812), .B(n805), .Z(n864) );
  XOR U1011 ( .A(n870), .B(n871), .Z(n805) );
  AND U1012 ( .A(n872), .B(n873), .Z(n871) );
  XNOR U1013 ( .A(n870), .B(n874), .Z(n873) );
  XNOR U1014 ( .A(n875), .B(n810), .Z(n812) );
  IV U1015 ( .A(n814), .Z(n810) );
  XNOR U1016 ( .A(n876), .B(n877), .Z(n814) );
  AND U1017 ( .A(n878), .B(n879), .Z(n877) );
  XNOR U1018 ( .A(n876), .B(n880), .Z(n879) );
  XNOR U1019 ( .A(n881), .B(n882), .Z(n875) );
  AND U1020 ( .A(n883), .B(n884), .Z(n882) );
  XOR U1021 ( .A(n885), .B(n886), .Z(n884) );
  IV U1022 ( .A(n881), .Z(n885) );
  XOR U1023 ( .A(n822), .B(n887), .Z(n803) );
  IV U1024 ( .A(n821), .Z(n887) );
  XNOR U1025 ( .A(n888), .B(n828), .Z(n821) );
  XNOR U1026 ( .A(n889), .B(n890), .Z(n828) );
  ANDN U1027 ( .A(n891), .B(n892), .Z(n890) );
  XNOR U1028 ( .A(n889), .B(n893), .Z(n891) );
  XNOR U1029 ( .A(n825), .B(n818), .Z(n888) );
  XOR U1030 ( .A(n894), .B(n895), .Z(n818) );
  ANDN U1031 ( .A(n896), .B(n897), .Z(n895) );
  XNOR U1032 ( .A(n894), .B(n898), .Z(n896) );
  XNOR U1033 ( .A(n899), .B(n823), .Z(n825) );
  IV U1034 ( .A(n827), .Z(n823) );
  XNOR U1035 ( .A(n900), .B(n901), .Z(n827) );
  AND U1036 ( .A(n902), .B(n903), .Z(n901) );
  XNOR U1037 ( .A(n900), .B(n904), .Z(n903) );
  XNOR U1038 ( .A(n905), .B(n906), .Z(n899) );
  AND U1039 ( .A(n907), .B(n908), .Z(n906) );
  XOR U1040 ( .A(n909), .B(n910), .Z(n908) );
  IV U1041 ( .A(n905), .Z(n909) );
  XOR U1042 ( .A(n834), .B(n911), .Z(n822) );
  IV U1043 ( .A(n832), .Z(n911) );
  XOR U1044 ( .A(n912), .B(n829), .Z(n832) );
  IV U1045 ( .A(n833), .Z(n829) );
  XNOR U1046 ( .A(n913), .B(n914), .Z(n833) );
  ANDN U1047 ( .A(n915), .B(n916), .Z(n914) );
  XNOR U1048 ( .A(n913), .B(n917), .Z(n915) );
  XNOR U1049 ( .A(n918), .B(n919), .Z(n912) );
  AND U1050 ( .A(n920), .B(n921), .Z(n919) );
  XOR U1051 ( .A(n922), .B(n923), .Z(n921) );
  IV U1052 ( .A(n918), .Z(n922) );
  XNOR U1053 ( .A(n924), .B(n925), .Z(n834) );
  ANDN U1054 ( .A(n926), .B(n927), .Z(n925) );
  XNOR U1055 ( .A(n924), .B(n928), .Z(n926) );
  XNOR U1056 ( .A(n836), .B(\min_dist_reg[3][1] ), .Z(n837) );
  NOR U1057 ( .A(\min_dist_reg[3][0] ), .B(n929), .Z(n836) );
  XOR U1058 ( .A(n750), .B(n929), .Z(n751) );
  XOR U1059 ( .A(n863), .B(n930), .Z(n929) );
  IV U1060 ( .A(n862), .Z(n930) );
  XNOR U1061 ( .A(n931), .B(n874), .Z(n862) );
  XOR U1062 ( .A(n847), .B(n932), .Z(n874) );
  IV U1063 ( .A(n846), .Z(n932) );
  XNOR U1064 ( .A(n933), .B(n853), .Z(n846) );
  XNOR U1065 ( .A(e_input[23]), .B(g_input[23]), .Z(n853) );
  XNOR U1066 ( .A(n843), .B(n850), .Z(n933) );
  XNOR U1067 ( .A(n934), .B(n848), .Z(n850) );
  XOR U1068 ( .A(e_input[21]), .B(g_input[21]), .Z(n848) );
  XNOR U1069 ( .A(e_input[22]), .B(g_input[22]), .Z(n934) );
  XOR U1070 ( .A(e_input[17]), .B(g_input[17]), .Z(n843) );
  XOR U1071 ( .A(n858), .B(n935), .Z(n847) );
  IV U1072 ( .A(n857), .Z(n935) );
  XOR U1073 ( .A(n936), .B(n854), .Z(n857) );
  XOR U1074 ( .A(e_input[18]), .B(g_input[18]), .Z(n854) );
  XNOR U1075 ( .A(e_input[19]), .B(g_input[19]), .Z(n936) );
  XNOR U1076 ( .A(e_input[20]), .B(g_input[20]), .Z(n858) );
  XNOR U1077 ( .A(n872), .B(n859), .Z(n931) );
  XOR U1078 ( .A(e_input[0]), .B(g_input[0]), .Z(n859) );
  XOR U1079 ( .A(n937), .B(n880), .Z(n872) );
  XOR U1080 ( .A(n869), .B(n938), .Z(n880) );
  IV U1081 ( .A(n868), .Z(n938) );
  XOR U1082 ( .A(n939), .B(n865), .Z(n868) );
  XOR U1083 ( .A(e_input[25]), .B(g_input[25]), .Z(n865) );
  XNOR U1084 ( .A(e_input[26]), .B(g_input[26]), .Z(n939) );
  XNOR U1085 ( .A(e_input[27]), .B(g_input[27]), .Z(n869) );
  XNOR U1086 ( .A(n878), .B(n870), .Z(n937) );
  XOR U1087 ( .A(e_input[16]), .B(g_input[16]), .Z(n870) );
  XOR U1088 ( .A(n940), .B(n886), .Z(n878) );
  XNOR U1089 ( .A(e_input[30]), .B(g_input[30]), .Z(n886) );
  XNOR U1090 ( .A(n876), .B(n883), .Z(n940) );
  XNOR U1091 ( .A(n941), .B(n881), .Z(n883) );
  XOR U1092 ( .A(e_input[28]), .B(g_input[28]), .Z(n881) );
  XNOR U1093 ( .A(e_input[29]), .B(g_input[29]), .Z(n941) );
  XOR U1094 ( .A(e_input[24]), .B(g_input[24]), .Z(n876) );
  XOR U1095 ( .A(n898), .B(n942), .Z(n863) );
  IV U1096 ( .A(n897), .Z(n942) );
  XNOR U1097 ( .A(n943), .B(n904), .Z(n897) );
  XOR U1098 ( .A(n893), .B(n944), .Z(n904) );
  IV U1099 ( .A(n892), .Z(n944) );
  XOR U1100 ( .A(n945), .B(n889), .Z(n892) );
  XOR U1101 ( .A(e_input[10]), .B(g_input[10]), .Z(n889) );
  XNOR U1102 ( .A(e_input[11]), .B(g_input[11]), .Z(n945) );
  XNOR U1103 ( .A(e_input[12]), .B(g_input[12]), .Z(n893) );
  XNOR U1104 ( .A(n902), .B(n894), .Z(n943) );
  XOR U1105 ( .A(e_input[1]), .B(g_input[1]), .Z(n894) );
  XOR U1106 ( .A(n946), .B(n910), .Z(n902) );
  XNOR U1107 ( .A(e_input[15]), .B(g_input[15]), .Z(n910) );
  XNOR U1108 ( .A(n900), .B(n907), .Z(n946) );
  XNOR U1109 ( .A(n947), .B(n905), .Z(n907) );
  XOR U1110 ( .A(e_input[13]), .B(g_input[13]), .Z(n905) );
  XNOR U1111 ( .A(e_input[14]), .B(g_input[14]), .Z(n947) );
  XOR U1112 ( .A(e_input[9]), .B(g_input[9]), .Z(n900) );
  XOR U1113 ( .A(n917), .B(n948), .Z(n898) );
  IV U1114 ( .A(n916), .Z(n948) );
  XNOR U1115 ( .A(n949), .B(n923), .Z(n916) );
  XNOR U1116 ( .A(e_input[8]), .B(g_input[8]), .Z(n923) );
  XNOR U1117 ( .A(n913), .B(n920), .Z(n949) );
  XNOR U1118 ( .A(n950), .B(n918), .Z(n920) );
  XOR U1119 ( .A(e_input[6]), .B(g_input[6]), .Z(n918) );
  XNOR U1120 ( .A(e_input[7]), .B(g_input[7]), .Z(n950) );
  XOR U1121 ( .A(e_input[2]), .B(g_input[2]), .Z(n913) );
  XOR U1122 ( .A(n928), .B(n951), .Z(n917) );
  IV U1123 ( .A(n927), .Z(n951) );
  XOR U1124 ( .A(n952), .B(n924), .Z(n927) );
  XOR U1125 ( .A(e_input[3]), .B(g_input[3]), .Z(n924) );
  XNOR U1126 ( .A(e_input[4]), .B(g_input[4]), .Z(n952) );
  XNOR U1127 ( .A(e_input[5]), .B(g_input[5]), .Z(n928) );
  IV U1128 ( .A(\min_dist_reg[3][0] ), .Z(n750) );
  IV U1129 ( .A(\min_dist_reg[1][0] ), .Z(n720) );
endmodule

