
module compare_N16384_CC2 ( clk, rst, x, y, g, e );
  input [8191:0] x;
  input [8191:0] y;
  input clk, rst;
  output g, e;
  wire   ebreg, n4, n5, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
         n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
         n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
         n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
         n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
         n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
         n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
         n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
         n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
         n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
         n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
         n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
         n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
         n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
         n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
         n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
         n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
         n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
         n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
         n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
         n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
         n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
         n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
         n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
         n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
         n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
         n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
         n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
         n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
         n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
         n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
         n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
         n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193,
         n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
         n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
         n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
         n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
         n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
         n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
         n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
         n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
         n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
         n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
         n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
         n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
         n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
         n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
         n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
         n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
         n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
         n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
         n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
         n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
         n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
         n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
         n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
         n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373,
         n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383,
         n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393,
         n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403,
         n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413,
         n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423,
         n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433,
         n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
         n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
         n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
         n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
         n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
         n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
         n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
         n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
         n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
         n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
         n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
         n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
         n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
         n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
         n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
         n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
         n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
         n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
         n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
         n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
         n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
         n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
         n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
         n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
         n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
         n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
         n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
         n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
         n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723,
         n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
         n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
         n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753,
         n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763,
         n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773,
         n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783,
         n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793,
         n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803,
         n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813,
         n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823,
         n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
         n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
         n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
         n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863,
         n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873,
         n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883,
         n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893,
         n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903,
         n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913,
         n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923,
         n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933,
         n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943,
         n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
         n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
         n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973,
         n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983,
         n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993,
         n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003,
         n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013,
         n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023,
         n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033,
         n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043,
         n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053,
         n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063,
         n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073,
         n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083,
         n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093,
         n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103,
         n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113,
         n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123,
         n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133,
         n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143,
         n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153,
         n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163,
         n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173,
         n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
         n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
         n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
         n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
         n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223,
         n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233,
         n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243,
         n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253,
         n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263,
         n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273,
         n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283,
         n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293,
         n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303,
         n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313,
         n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323,
         n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333,
         n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343,
         n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353,
         n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363,
         n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373,
         n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383,
         n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393,
         n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403,
         n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413,
         n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423,
         n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433,
         n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443,
         n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453,
         n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463,
         n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473,
         n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483,
         n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493,
         n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503,
         n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513,
         n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523,
         n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533,
         n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543,
         n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553,
         n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563,
         n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573,
         n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583,
         n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593,
         n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603,
         n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613,
         n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623,
         n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633,
         n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643,
         n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653,
         n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663,
         n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673,
         n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683,
         n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693,
         n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703,
         n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713,
         n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723,
         n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733,
         n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743,
         n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753,
         n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763,
         n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773,
         n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783,
         n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793,
         n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803,
         n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813,
         n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823,
         n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833,
         n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843,
         n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853,
         n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863,
         n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873,
         n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883,
         n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893,
         n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903,
         n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913,
         n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923,
         n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933,
         n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943,
         n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953,
         n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963,
         n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973,
         n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983,
         n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993,
         n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003,
         n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013,
         n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023,
         n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033,
         n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043,
         n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053,
         n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063,
         n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073,
         n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083,
         n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093,
         n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103,
         n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113,
         n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123,
         n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133,
         n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143,
         n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153,
         n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163,
         n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173,
         n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183,
         n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193,
         n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203,
         n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213,
         n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223,
         n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233,
         n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243,
         n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253,
         n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263,
         n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273,
         n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283,
         n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293,
         n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303,
         n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313,
         n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323,
         n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333,
         n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343,
         n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353,
         n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363,
         n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373,
         n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383,
         n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393,
         n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403,
         n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413,
         n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
         n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433,
         n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443,
         n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453,
         n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463,
         n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
         n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483,
         n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
         n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
         n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
         n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523,
         n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533,
         n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543,
         n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553,
         n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563,
         n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573,
         n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583,
         n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
         n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603,
         n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613,
         n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623,
         n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633,
         n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643,
         n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653,
         n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
         n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673,
         n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683,
         n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693,
         n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703,
         n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713,
         n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723,
         n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733,
         n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
         n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
         n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
         n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783,
         n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793,
         n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803,
         n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813,
         n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
         n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
         n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
         n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
         n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
         n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
         n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
         n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
         n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
         n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
         n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386,
         n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
         n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
         n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
         n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
         n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,
         n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
         n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
         n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554,
         n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562,
         n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570,
         n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578,
         n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586,
         n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594,
         n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602,
         n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610,
         n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618,
         n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626,
         n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634,
         n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642,
         n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650,
         n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658,
         n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666,
         n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674,
         n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682,
         n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690,
         n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698,
         n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706,
         n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714,
         n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722,
         n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730,
         n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738,
         n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746,
         n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754,
         n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762,
         n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770,
         n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778,
         n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786,
         n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794,
         n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802,
         n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810,
         n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818,
         n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826,
         n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834,
         n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842,
         n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850,
         n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858,
         n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866,
         n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874,
         n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882,
         n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890,
         n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898,
         n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906,
         n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914,
         n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922,
         n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930,
         n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938,
         n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946,
         n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954,
         n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962,
         n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970,
         n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978,
         n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986,
         n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994,
         n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002,
         n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010,
         n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018,
         n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026,
         n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034,
         n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042,
         n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050,
         n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058,
         n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066,
         n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074,
         n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082,
         n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090,
         n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098,
         n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106,
         n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114,
         n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122,
         n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130,
         n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138,
         n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146,
         n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154,
         n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162,
         n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170,
         n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178,
         n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186,
         n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194,
         n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202,
         n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210,
         n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218,
         n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226,
         n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234,
         n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242,
         n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250,
         n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258,
         n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266,
         n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274,
         n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282,
         n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290,
         n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298,
         n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306,
         n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314,
         n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322,
         n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330,
         n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338,
         n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346,
         n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354,
         n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362,
         n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370,
         n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378,
         n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386,
         n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394,
         n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402,
         n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410,
         n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418,
         n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426,
         n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434,
         n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442,
         n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450,
         n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458,
         n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466,
         n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474,
         n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482,
         n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490,
         n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498,
         n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506,
         n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514,
         n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522,
         n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530,
         n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538,
         n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546,
         n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554,
         n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562,
         n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570,
         n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578,
         n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586,
         n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594,
         n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602,
         n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610,
         n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618,
         n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626,
         n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634,
         n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642,
         n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650,
         n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658,
         n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666,
         n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674,
         n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682,
         n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690,
         n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698,
         n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706,
         n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714,
         n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722,
         n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730,
         n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738,
         n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746,
         n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754,
         n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762,
         n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770,
         n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778,
         n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786,
         n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794,
         n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802,
         n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810,
         n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818,
         n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826,
         n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834,
         n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842,
         n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850,
         n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858,
         n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866,
         n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874,
         n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882,
         n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890,
         n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898,
         n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906,
         n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914,
         n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922,
         n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930,
         n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938,
         n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946,
         n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954,
         n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962,
         n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970,
         n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978,
         n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986,
         n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994,
         n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002,
         n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010,
         n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018,
         n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026,
         n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034,
         n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042,
         n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050,
         n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058,
         n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066,
         n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074,
         n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082,
         n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090,
         n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098,
         n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106,
         n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114,
         n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122,
         n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130,
         n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138,
         n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146,
         n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154,
         n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162,
         n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170,
         n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178,
         n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186,
         n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194,
         n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202,
         n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210,
         n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218,
         n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226,
         n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234,
         n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242,
         n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250,
         n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258,
         n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266,
         n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274,
         n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282,
         n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290,
         n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,
         n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306,
         n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314,
         n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322,
         n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330,
         n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338,
         n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346,
         n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354,
         n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362,
         n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370,
         n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378,
         n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386,
         n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394,
         n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402,
         n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410,
         n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418,
         n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426,
         n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434,
         n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442,
         n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450,
         n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458,
         n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466,
         n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474,
         n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482,
         n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490,
         n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498,
         n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506,
         n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514,
         n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522,
         n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530,
         n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538,
         n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546,
         n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554,
         n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562,
         n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570,
         n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578,
         n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586,
         n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594,
         n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602,
         n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610,
         n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618,
         n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626,
         n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634,
         n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642,
         n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650,
         n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658,
         n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666,
         n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674,
         n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682,
         n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690,
         n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698,
         n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706,
         n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714,
         n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722,
         n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730,
         n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738,
         n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746,
         n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754,
         n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762,
         n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770,
         n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778,
         n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786,
         n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794,
         n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802,
         n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810,
         n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818,
         n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826,
         n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834,
         n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842,
         n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850,
         n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858,
         n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866,
         n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874,
         n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882,
         n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890,
         n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898,
         n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906,
         n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914,
         n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922,
         n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930,
         n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938,
         n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946,
         n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954,
         n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962,
         n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970,
         n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978,
         n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986,
         n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994,
         n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002,
         n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010,
         n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018,
         n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026,
         n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034,
         n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042,
         n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050,
         n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058,
         n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066,
         n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074,
         n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082,
         n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090,
         n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098,
         n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106,
         n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114,
         n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122,
         n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130,
         n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138,
         n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146,
         n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154,
         n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162,
         n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170,
         n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178,
         n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186,
         n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194,
         n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202,
         n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210,
         n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218,
         n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226,
         n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234,
         n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242,
         n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250,
         n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258,
         n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266,
         n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274,
         n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282,
         n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290,
         n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298,
         n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306,
         n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314,
         n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322,
         n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330,
         n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338,
         n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346,
         n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354,
         n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362,
         n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370,
         n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378,
         n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386,
         n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394,
         n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402,
         n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410,
         n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418,
         n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426,
         n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434,
         n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,
         n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450,
         n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458,
         n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466,
         n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474,
         n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
         n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490,
         n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498,
         n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506,
         n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,
         n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522,
         n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530,
         n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538,
         n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
         n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
         n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,
         n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,
         n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578,
         n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586,
         n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594,
         n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602,
         n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610,
         n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618,
         n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626,
         n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634,
         n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642,
         n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650,
         n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,
         n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666,
         n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674,
         n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682,
         n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690,
         n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698,
         n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706,
         n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714,
         n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722,
         n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730,
         n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738,
         n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746,
         n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754,
         n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762,
         n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770,
         n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778,
         n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786,
         n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794,
         n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802,
         n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810,
         n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818,
         n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826,
         n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834,
         n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842,
         n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
         n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858,
         n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866,
         n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
         n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882,
         n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890,
         n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898,
         n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906,
         n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914,
         n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,
         n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930,
         n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938,
         n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
         n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,
         n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
         n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970,
         n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
         n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
         n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
         n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
         n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,
         n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
         n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,
         n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034,
         n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042,
         n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,
         n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058,
         n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066,
         n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074,
         n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082,
         n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090,
         n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,
         n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106,
         n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114,
         n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122,
         n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130,
         n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138,
         n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146,
         n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154,
         n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162,
         n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170,
         n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178,
         n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186,
         n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194,
         n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202,
         n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210,
         n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218,
         n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226,
         n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234,
         n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242,
         n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250,
         n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258,
         n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266,
         n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274,
         n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282,
         n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290,
         n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298,
         n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306,
         n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314,
         n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322,
         n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330,
         n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338,
         n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346,
         n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354,
         n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362,
         n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370,
         n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378,
         n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386,
         n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394,
         n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402,
         n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410,
         n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418,
         n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426,
         n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434,
         n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442,
         n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450,
         n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458,
         n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466,
         n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474,
         n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482,
         n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490,
         n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498,
         n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506,
         n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514,
         n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522,
         n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530,
         n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538,
         n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546,
         n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554,
         n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562,
         n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570,
         n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578,
         n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586,
         n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594,
         n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602,
         n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610,
         n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618,
         n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626,
         n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634,
         n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642,
         n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650,
         n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658,
         n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666,
         n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674,
         n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682,
         n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690,
         n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698,
         n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706,
         n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714,
         n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722,
         n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730,
         n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738,
         n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746,
         n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754,
         n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762,
         n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770,
         n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778,
         n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786,
         n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794,
         n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802,
         n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810,
         n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818,
         n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826,
         n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834,
         n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842,
         n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850,
         n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858,
         n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866,
         n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874,
         n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882,
         n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890,
         n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898,
         n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906,
         n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914,
         n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922,
         n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930,
         n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938,
         n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946,
         n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954,
         n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962,
         n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970,
         n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978,
         n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986,
         n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994,
         n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002,
         n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010,
         n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018,
         n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026,
         n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034,
         n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042,
         n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050,
         n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058,
         n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066,
         n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074,
         n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082,
         n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090,
         n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098,
         n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106,
         n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114,
         n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122,
         n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130,
         n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138,
         n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146,
         n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154,
         n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162,
         n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170,
         n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178,
         n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186,
         n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194,
         n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202,
         n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210,
         n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218,
         n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226,
         n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234,
         n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242,
         n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250,
         n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258,
         n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266,
         n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274,
         n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282,
         n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290,
         n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298,
         n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306,
         n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314,
         n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322,
         n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330,
         n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338,
         n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346,
         n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354,
         n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362,
         n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370,
         n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378,
         n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386,
         n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394,
         n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402,
         n15403, n15404, n15405, n15406, n15407, n15408, n15409, n15410,
         n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418,
         n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426,
         n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434,
         n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442,
         n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450,
         n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458,
         n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466,
         n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474,
         n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482,
         n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490,
         n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498,
         n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506,
         n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514,
         n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522,
         n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530,
         n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538,
         n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546,
         n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554,
         n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562,
         n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570,
         n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578,
         n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586,
         n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15594,
         n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602,
         n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610,
         n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618,
         n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626,
         n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634,
         n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642,
         n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650,
         n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658,
         n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666,
         n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674,
         n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682,
         n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690,
         n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698,
         n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706,
         n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714,
         n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722,
         n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730,
         n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738,
         n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746,
         n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754,
         n15755, n15756, n15757, n15758, n15759, n15760, n15761, n15762,
         n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770,
         n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778,
         n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786,
         n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794,
         n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802,
         n15803, n15804, n15805, n15806, n15807, n15808, n15809, n15810,
         n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818,
         n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826,
         n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834,
         n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842,
         n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850,
         n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858,
         n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866,
         n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874,
         n15875, n15876, n15877, n15878, n15879, n15880, n15881, n15882,
         n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890,
         n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898,
         n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906,
         n15907, n15908, n15909, n15910, n15911, n15912, n15913, n15914,
         n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922,
         n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930,
         n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938,
         n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946,
         n15947, n15948, n15949, n15950, n15951, n15952, n15953, n15954,
         n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962,
         n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970,
         n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978,
         n15979, n15980, n15981, n15982, n15983, n15984, n15985, n15986,
         n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994,
         n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002,
         n16003, n16004, n16005, n16006, n16007, n16008, n16009, n16010,
         n16011, n16012, n16013, n16014, n16015, n16016, n16017, n16018,
         n16019, n16020, n16021, n16022, n16023, n16024, n16025, n16026,
         n16027, n16028, n16029, n16030, n16031, n16032, n16033, n16034,
         n16035, n16036, n16037, n16038, n16039, n16040, n16041, n16042,
         n16043, n16044, n16045, n16046, n16047, n16048, n16049, n16050,
         n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058,
         n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066,
         n16067, n16068, n16069, n16070, n16071, n16072, n16073, n16074,
         n16075, n16076, n16077, n16078, n16079, n16080, n16081, n16082,
         n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090,
         n16091, n16092, n16093, n16094, n16095, n16096, n16097, n16098,
         n16099, n16100, n16101, n16102, n16103, n16104, n16105, n16106,
         n16107, n16108, n16109, n16110, n16111, n16112, n16113, n16114,
         n16115, n16116, n16117, n16118, n16119, n16120, n16121, n16122,
         n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130,
         n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138,
         n16139, n16140, n16141, n16142, n16143, n16144, n16145, n16146,
         n16147, n16148, n16149, n16150, n16151, n16152, n16153, n16154,
         n16155, n16156, n16157, n16158, n16159, n16160, n16161, n16162,
         n16163, n16164, n16165, n16166, n16167, n16168, n16169, n16170,
         n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178,
         n16179, n16180, n16181, n16182, n16183, n16184, n16185, n16186,
         n16187, n16188, n16189, n16190, n16191, n16192, n16193, n16194,
         n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202,
         n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210,
         n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218,
         n16219, n16220, n16221, n16222, n16223, n16224, n16225, n16226,
         n16227, n16228, n16229, n16230, n16231, n16232, n16233, n16234,
         n16235, n16236, n16237, n16238, n16239, n16240, n16241, n16242,
         n16243, n16244, n16245, n16246, n16247, n16248, n16249, n16250,
         n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16258,
         n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16266,
         n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16274,
         n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282,
         n16283, n16284, n16285, n16286, n16287, n16288, n16289, n16290,
         n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298,
         n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16306,
         n16307, n16308, n16309, n16310, n16311, n16312, n16313, n16314,
         n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322,
         n16323, n16324, n16325, n16326, n16327, n16328, n16329, n16330,
         n16331, n16332, n16333, n16334, n16335, n16336, n16337, n16338,
         n16339, n16340, n16341, n16342, n16343, n16344, n16345, n16346,
         n16347, n16348, n16349, n16350, n16351, n16352, n16353, n16354,
         n16355, n16356, n16357, n16358, n16359, n16360, n16361, n16362,
         n16363, n16364, n16365, n16366, n16367, n16368, n16369, n16370,
         n16371, n16372, n16373, n16374, n16375, n16376, n16377, n16378,
         n16379, n16380, n16381, n16382, n16383, n16384, n16385, n16386,
         n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394,
         n16395, n16396, n16397, n16398, n16399, n16400, n16401, n16402,
         n16403, n16404, n16405, n16406, n16407, n16408, n16409, n16410,
         n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418,
         n16419, n16420, n16421, n16422, n16423, n16424, n16425, n16426,
         n16427, n16428, n16429, n16430, n16431, n16432, n16433, n16434,
         n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442,
         n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450,
         n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16458,
         n16459, n16460, n16461, n16462, n16463, n16464, n16465, n16466,
         n16467, n16468, n16469, n16470, n16471, n16472, n16473, n16474,
         n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16482,
         n16483, n16484, n16485, n16486, n16487, n16488, n16489, n16490,
         n16491, n16492, n16493, n16494, n16495, n16496, n16497, n16498,
         n16499, n16500, n16501, n16502, n16503, n16504, n16505, n16506,
         n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514,
         n16515, n16516, n16517, n16518, n16519, n16520, n16521, n16522,
         n16523, n16524, n16525, n16526, n16527, n16528, n16529, n16530,
         n16531, n16532, n16533, n16534, n16535, n16536, n16537, n16538,
         n16539, n16540, n16541, n16542, n16543, n16544, n16545, n16546,
         n16547, n16548, n16549, n16550, n16551, n16552, n16553, n16554,
         n16555, n16556, n16557, n16558, n16559, n16560, n16561, n16562,
         n16563, n16564, n16565, n16566, n16567, n16568, n16569, n16570,
         n16571, n16572, n16573, n16574, n16575, n16576, n16577, n16578,
         n16579, n16580, n16581, n16582, n16583, n16584, n16585, n16586,
         n16587, n16588, n16589, n16590, n16591, n16592, n16593, n16594,
         n16595, n16596, n16597, n16598, n16599, n16600, n16601, n16602,
         n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610,
         n16611, n16612, n16613, n16614, n16615, n16616, n16617, n16618,
         n16619, n16620, n16621, n16622, n16623, n16624, n16625, n16626,
         n16627, n16628, n16629, n16630, n16631, n16632, n16633, n16634,
         n16635, n16636, n16637, n16638, n16639, n16640, n16641, n16642,
         n16643, n16644, n16645, n16646, n16647, n16648, n16649, n16650,
         n16651, n16652, n16653, n16654, n16655, n16656, n16657, n16658,
         n16659, n16660, n16661, n16662, n16663, n16664, n16665, n16666,
         n16667, n16668, n16669, n16670, n16671, n16672, n16673, n16674,
         n16675, n16676, n16677, n16678, n16679, n16680, n16681, n16682,
         n16683, n16684, n16685, n16686, n16687, n16688, n16689, n16690,
         n16691, n16692, n16693, n16694, n16695, n16696, n16697, n16698,
         n16699, n16700, n16701, n16702, n16703, n16704, n16705, n16706,
         n16707, n16708, n16709, n16710, n16711, n16712, n16713, n16714,
         n16715, n16716, n16717, n16718, n16719, n16720, n16721, n16722,
         n16723, n16724, n16725, n16726, n16727, n16728, n16729, n16730,
         n16731, n16732, n16733, n16734, n16735, n16736, n16737, n16738,
         n16739, n16740, n16741, n16742, n16743, n16744, n16745, n16746,
         n16747, n16748, n16749, n16750, n16751, n16752, n16753, n16754,
         n16755, n16756, n16757, n16758, n16759, n16760, n16761, n16762,
         n16763, n16764, n16765, n16766, n16767, n16768, n16769, n16770,
         n16771, n16772, n16773, n16774, n16775, n16776, n16777, n16778,
         n16779, n16780, n16781, n16782, n16783, n16784, n16785, n16786,
         n16787, n16788, n16789, n16790, n16791, n16792, n16793, n16794,
         n16795, n16796, n16797, n16798, n16799, n16800, n16801, n16802,
         n16803, n16804, n16805, n16806, n16807, n16808, n16809, n16810,
         n16811, n16812, n16813, n16814, n16815, n16816, n16817, n16818,
         n16819, n16820, n16821, n16822, n16823, n16824, n16825, n16826,
         n16827, n16828, n16829, n16830, n16831, n16832, n16833, n16834,
         n16835, n16836, n16837, n16838, n16839, n16840, n16841, n16842,
         n16843, n16844, n16845, n16846, n16847, n16848, n16849, n16850,
         n16851, n16852, n16853, n16854, n16855, n16856, n16857, n16858,
         n16859, n16860, n16861, n16862, n16863, n16864, n16865, n16866,
         n16867, n16868, n16869, n16870, n16871, n16872, n16873, n16874,
         n16875, n16876, n16877, n16878, n16879, n16880, n16881, n16882,
         n16883, n16884, n16885, n16886, n16887, n16888, n16889, n16890,
         n16891, n16892, n16893, n16894, n16895, n16896, n16897, n16898,
         n16899, n16900, n16901, n16902, n16903, n16904, n16905, n16906,
         n16907, n16908, n16909, n16910, n16911, n16912, n16913, n16914,
         n16915, n16916, n16917, n16918, n16919, n16920, n16921, n16922,
         n16923, n16924, n16925, n16926, n16927, n16928, n16929, n16930,
         n16931, n16932, n16933, n16934, n16935, n16936, n16937, n16938,
         n16939, n16940, n16941, n16942, n16943, n16944, n16945, n16946,
         n16947, n16948, n16949, n16950, n16951, n16952, n16953, n16954,
         n16955, n16956, n16957, n16958, n16959, n16960, n16961, n16962,
         n16963, n16964, n16965, n16966, n16967, n16968, n16969, n16970,
         n16971, n16972, n16973, n16974, n16975, n16976, n16977, n16978,
         n16979, n16980, n16981, n16982, n16983, n16984, n16985, n16986,
         n16987, n16988, n16989, n16990, n16991, n16992, n16993, n16994,
         n16995, n16996, n16997, n16998, n16999, n17000, n17001, n17002,
         n17003, n17004, n17005, n17006, n17007, n17008, n17009, n17010,
         n17011, n17012, n17013, n17014, n17015, n17016, n17017, n17018,
         n17019, n17020, n17021, n17022, n17023, n17024, n17025, n17026,
         n17027, n17028, n17029, n17030, n17031, n17032, n17033, n17034,
         n17035, n17036, n17037, n17038, n17039, n17040, n17041, n17042,
         n17043, n17044, n17045, n17046, n17047, n17048, n17049, n17050,
         n17051, n17052, n17053, n17054, n17055, n17056, n17057, n17058,
         n17059, n17060, n17061, n17062, n17063, n17064, n17065, n17066,
         n17067, n17068, n17069, n17070, n17071, n17072, n17073, n17074,
         n17075, n17076, n17077, n17078, n17079, n17080, n17081, n17082,
         n17083, n17084, n17085, n17086, n17087, n17088, n17089, n17090,
         n17091, n17092, n17093, n17094, n17095, n17096, n17097, n17098,
         n17099, n17100, n17101, n17102, n17103, n17104, n17105, n17106,
         n17107, n17108, n17109, n17110, n17111, n17112, n17113, n17114,
         n17115, n17116, n17117, n17118, n17119, n17120, n17121, n17122,
         n17123, n17124, n17125, n17126, n17127, n17128, n17129, n17130,
         n17131, n17132, n17133, n17134, n17135, n17136, n17137, n17138,
         n17139, n17140, n17141, n17142, n17143, n17144, n17145, n17146,
         n17147, n17148, n17149, n17150, n17151, n17152, n17153, n17154,
         n17155, n17156, n17157, n17158, n17159, n17160, n17161, n17162,
         n17163, n17164, n17165, n17166, n17167, n17168, n17169, n17170,
         n17171, n17172, n17173, n17174, n17175, n17176, n17177, n17178,
         n17179, n17180, n17181, n17182, n17183, n17184, n17185, n17186,
         n17187, n17188, n17189, n17190, n17191, n17192, n17193, n17194,
         n17195, n17196, n17197, n17198, n17199, n17200, n17201, n17202,
         n17203, n17204, n17205, n17206, n17207, n17208, n17209, n17210,
         n17211, n17212, n17213, n17214, n17215, n17216, n17217, n17218,
         n17219, n17220, n17221, n17222, n17223, n17224, n17225, n17226,
         n17227, n17228, n17229, n17230, n17231, n17232, n17233, n17234,
         n17235, n17236, n17237, n17238, n17239, n17240, n17241, n17242,
         n17243, n17244, n17245, n17246, n17247, n17248, n17249, n17250,
         n17251, n17252, n17253, n17254, n17255, n17256, n17257, n17258,
         n17259, n17260, n17261, n17262, n17263, n17264, n17265, n17266,
         n17267, n17268, n17269, n17270, n17271, n17272, n17273, n17274,
         n17275, n17276, n17277, n17278, n17279, n17280, n17281, n17282,
         n17283, n17284, n17285, n17286, n17287, n17288, n17289, n17290,
         n17291, n17292, n17293, n17294, n17295, n17296, n17297, n17298,
         n17299, n17300, n17301, n17302, n17303, n17304, n17305, n17306,
         n17307, n17308, n17309, n17310, n17311, n17312, n17313, n17314,
         n17315, n17316, n17317, n17318, n17319, n17320, n17321, n17322,
         n17323, n17324, n17325, n17326, n17327, n17328, n17329, n17330,
         n17331, n17332, n17333, n17334, n17335, n17336, n17337, n17338,
         n17339, n17340, n17341, n17342, n17343, n17344, n17345, n17346,
         n17347, n17348, n17349, n17350, n17351, n17352, n17353, n17354,
         n17355, n17356, n17357, n17358, n17359, n17360, n17361, n17362,
         n17363, n17364, n17365, n17366, n17367, n17368, n17369, n17370,
         n17371, n17372, n17373, n17374, n17375, n17376, n17377, n17378,
         n17379, n17380, n17381, n17382, n17383, n17384, n17385, n17386,
         n17387, n17388, n17389, n17390, n17391, n17392, n17393, n17394,
         n17395, n17396, n17397, n17398, n17399, n17400, n17401, n17402,
         n17403, n17404, n17405, n17406, n17407, n17408, n17409, n17410,
         n17411, n17412, n17413, n17414, n17415, n17416, n17417, n17418,
         n17419, n17420, n17421, n17422, n17423, n17424, n17425, n17426,
         n17427, n17428, n17429, n17430, n17431, n17432, n17433, n17434,
         n17435, n17436, n17437, n17438, n17439, n17440, n17441, n17442,
         n17443, n17444, n17445, n17446, n17447, n17448, n17449, n17450,
         n17451, n17452, n17453, n17454, n17455, n17456, n17457, n17458,
         n17459, n17460, n17461, n17462, n17463, n17464, n17465, n17466,
         n17467, n17468, n17469, n17470, n17471, n17472, n17473, n17474,
         n17475, n17476, n17477, n17478, n17479, n17480, n17481, n17482,
         n17483, n17484, n17485, n17486, n17487, n17488, n17489, n17490,
         n17491, n17492, n17493, n17494, n17495, n17496, n17497, n17498,
         n17499, n17500, n17501, n17502, n17503, n17504, n17505, n17506,
         n17507, n17508, n17509, n17510, n17511, n17512, n17513, n17514,
         n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522,
         n17523, n17524, n17525, n17526, n17527, n17528, n17529, n17530,
         n17531, n17532, n17533, n17534, n17535, n17536, n17537, n17538,
         n17539, n17540, n17541, n17542, n17543, n17544, n17545, n17546,
         n17547, n17548, n17549, n17550, n17551, n17552, n17553, n17554,
         n17555, n17556, n17557, n17558, n17559, n17560, n17561, n17562,
         n17563, n17564, n17565, n17566, n17567, n17568, n17569, n17570,
         n17571, n17572, n17573, n17574, n17575, n17576, n17577, n17578,
         n17579, n17580, n17581, n17582, n17583, n17584, n17585, n17586,
         n17587, n17588, n17589, n17590, n17591, n17592, n17593, n17594,
         n17595, n17596, n17597, n17598, n17599, n17600, n17601, n17602,
         n17603, n17604, n17605, n17606, n17607, n17608, n17609, n17610,
         n17611, n17612, n17613, n17614, n17615, n17616, n17617, n17618,
         n17619, n17620, n17621, n17622, n17623, n17624, n17625, n17626,
         n17627, n17628, n17629, n17630, n17631, n17632, n17633, n17634,
         n17635, n17636, n17637, n17638, n17639, n17640, n17641, n17642,
         n17643, n17644, n17645, n17646, n17647, n17648, n17649, n17650,
         n17651, n17652, n17653, n17654, n17655, n17656, n17657, n17658,
         n17659, n17660, n17661, n17662, n17663, n17664, n17665, n17666,
         n17667, n17668, n17669, n17670, n17671, n17672, n17673, n17674,
         n17675, n17676, n17677, n17678, n17679, n17680, n17681, n17682,
         n17683, n17684, n17685, n17686, n17687, n17688, n17689, n17690,
         n17691, n17692, n17693, n17694, n17695, n17696, n17697, n17698,
         n17699, n17700, n17701, n17702, n17703, n17704, n17705, n17706,
         n17707, n17708, n17709, n17710, n17711, n17712, n17713, n17714,
         n17715, n17716, n17717, n17718, n17719, n17720, n17721, n17722,
         n17723, n17724, n17725, n17726, n17727, n17728, n17729, n17730,
         n17731, n17732, n17733, n17734, n17735, n17736, n17737, n17738,
         n17739, n17740, n17741, n17742, n17743, n17744, n17745, n17746,
         n17747, n17748, n17749, n17750, n17751, n17752, n17753, n17754,
         n17755, n17756, n17757, n17758, n17759, n17760, n17761, n17762,
         n17763, n17764, n17765, n17766, n17767, n17768, n17769, n17770,
         n17771, n17772, n17773, n17774, n17775, n17776, n17777, n17778,
         n17779, n17780, n17781, n17782, n17783, n17784, n17785, n17786,
         n17787, n17788, n17789, n17790, n17791, n17792, n17793, n17794,
         n17795, n17796, n17797, n17798, n17799, n17800, n17801, n17802,
         n17803, n17804, n17805, n17806, n17807, n17808, n17809, n17810,
         n17811, n17812, n17813, n17814, n17815, n17816, n17817, n17818,
         n17819, n17820, n17821, n17822, n17823, n17824, n17825, n17826,
         n17827, n17828, n17829, n17830, n17831, n17832, n17833, n17834,
         n17835, n17836, n17837, n17838, n17839, n17840, n17841, n17842,
         n17843, n17844, n17845, n17846, n17847, n17848, n17849, n17850,
         n17851, n17852, n17853, n17854, n17855, n17856, n17857, n17858,
         n17859, n17860, n17861, n17862, n17863, n17864, n17865, n17866,
         n17867, n17868, n17869, n17870, n17871, n17872, n17873, n17874,
         n17875, n17876, n17877, n17878, n17879, n17880, n17881, n17882,
         n17883, n17884, n17885, n17886, n17887, n17888, n17889, n17890,
         n17891, n17892, n17893, n17894, n17895, n17896, n17897, n17898,
         n17899, n17900, n17901, n17902, n17903, n17904, n17905, n17906,
         n17907, n17908, n17909, n17910, n17911, n17912, n17913, n17914,
         n17915, n17916, n17917, n17918, n17919, n17920, n17921, n17922,
         n17923, n17924, n17925, n17926, n17927, n17928, n17929, n17930,
         n17931, n17932, n17933, n17934, n17935, n17936, n17937, n17938,
         n17939, n17940, n17941, n17942, n17943, n17944, n17945, n17946,
         n17947, n17948, n17949, n17950, n17951, n17952, n17953, n17954,
         n17955, n17956, n17957, n17958, n17959, n17960, n17961, n17962,
         n17963, n17964, n17965, n17966, n17967, n17968, n17969, n17970,
         n17971, n17972, n17973, n17974, n17975, n17976, n17977, n17978,
         n17979, n17980, n17981, n17982, n17983, n17984, n17985, n17986,
         n17987, n17988, n17989, n17990, n17991, n17992, n17993, n17994,
         n17995, n17996, n17997, n17998, n17999, n18000, n18001, n18002,
         n18003, n18004, n18005, n18006, n18007, n18008, n18009, n18010,
         n18011, n18012, n18013, n18014, n18015, n18016, n18017, n18018,
         n18019, n18020, n18021, n18022, n18023, n18024, n18025, n18026,
         n18027, n18028, n18029, n18030, n18031, n18032, n18033, n18034,
         n18035, n18036, n18037, n18038, n18039, n18040, n18041, n18042,
         n18043, n18044, n18045, n18046, n18047, n18048, n18049, n18050,
         n18051, n18052, n18053, n18054, n18055, n18056, n18057, n18058,
         n18059, n18060, n18061, n18062, n18063, n18064, n18065, n18066,
         n18067, n18068, n18069, n18070, n18071, n18072, n18073, n18074,
         n18075, n18076, n18077, n18078, n18079, n18080, n18081, n18082,
         n18083, n18084, n18085, n18086, n18087, n18088, n18089, n18090,
         n18091, n18092, n18093, n18094, n18095, n18096, n18097, n18098,
         n18099, n18100, n18101, n18102, n18103, n18104, n18105, n18106,
         n18107, n18108, n18109, n18110, n18111, n18112, n18113, n18114,
         n18115, n18116, n18117, n18118, n18119, n18120, n18121, n18122,
         n18123, n18124, n18125, n18126, n18127, n18128, n18129, n18130,
         n18131, n18132, n18133, n18134, n18135, n18136, n18137, n18138,
         n18139, n18140, n18141, n18142, n18143, n18144, n18145, n18146,
         n18147, n18148, n18149, n18150, n18151, n18152, n18153, n18154,
         n18155, n18156, n18157, n18158, n18159, n18160, n18161, n18162,
         n18163, n18164, n18165, n18166, n18167, n18168, n18169, n18170,
         n18171, n18172, n18173, n18174, n18175, n18176, n18177, n18178,
         n18179, n18180, n18181, n18182, n18183, n18184, n18185, n18186,
         n18187, n18188, n18189, n18190, n18191, n18192, n18193, n18194,
         n18195, n18196, n18197, n18198, n18199, n18200, n18201, n18202,
         n18203, n18204, n18205, n18206, n18207, n18208, n18209, n18210,
         n18211, n18212, n18213, n18214, n18215, n18216, n18217, n18218,
         n18219, n18220, n18221, n18222, n18223, n18224, n18225, n18226,
         n18227, n18228, n18229, n18230, n18231, n18232, n18233, n18234,
         n18235, n18236, n18237, n18238, n18239, n18240, n18241, n18242,
         n18243, n18244, n18245, n18246, n18247, n18248, n18249, n18250,
         n18251, n18252, n18253, n18254, n18255, n18256, n18257, n18258,
         n18259, n18260, n18261, n18262, n18263, n18264, n18265, n18266,
         n18267, n18268, n18269, n18270, n18271, n18272, n18273, n18274,
         n18275, n18276, n18277, n18278, n18279, n18280, n18281, n18282,
         n18283, n18284, n18285, n18286, n18287, n18288, n18289, n18290,
         n18291, n18292, n18293, n18294, n18295, n18296, n18297, n18298,
         n18299, n18300, n18301, n18302, n18303, n18304, n18305, n18306,
         n18307, n18308, n18309, n18310, n18311, n18312, n18313, n18314,
         n18315, n18316, n18317, n18318, n18319, n18320, n18321, n18322,
         n18323, n18324, n18325, n18326, n18327, n18328, n18329, n18330,
         n18331, n18332, n18333, n18334, n18335, n18336, n18337, n18338,
         n18339, n18340, n18341, n18342, n18343, n18344, n18345, n18346,
         n18347, n18348, n18349, n18350, n18351, n18352, n18353, n18354,
         n18355, n18356, n18357, n18358, n18359, n18360, n18361, n18362,
         n18363, n18364, n18365, n18366, n18367, n18368, n18369, n18370,
         n18371, n18372, n18373, n18374, n18375, n18376, n18377, n18378,
         n18379, n18380, n18381, n18382, n18383, n18384, n18385, n18386,
         n18387, n18388, n18389, n18390, n18391, n18392, n18393, n18394,
         n18395, n18396, n18397, n18398, n18399, n18400, n18401, n18402,
         n18403, n18404, n18405, n18406, n18407, n18408, n18409, n18410,
         n18411, n18412, n18413, n18414, n18415, n18416, n18417, n18418,
         n18419, n18420, n18421, n18422, n18423, n18424, n18425, n18426,
         n18427, n18428, n18429, n18430, n18431, n18432, n18433, n18434,
         n18435, n18436, n18437, n18438, n18439, n18440, n18441, n18442,
         n18443, n18444, n18445, n18446, n18447, n18448, n18449, n18450,
         n18451, n18452, n18453, n18454, n18455, n18456, n18457, n18458,
         n18459, n18460, n18461, n18462, n18463, n18464, n18465, n18466,
         n18467, n18468, n18469, n18470, n18471, n18472, n18473, n18474,
         n18475, n18476, n18477, n18478, n18479, n18480, n18481, n18482,
         n18483, n18484, n18485, n18486, n18487, n18488, n18489, n18490,
         n18491, n18492, n18493, n18494, n18495, n18496, n18497, n18498,
         n18499, n18500, n18501, n18502, n18503, n18504, n18505, n18506,
         n18507, n18508, n18509, n18510, n18511, n18512, n18513, n18514,
         n18515, n18516, n18517, n18518, n18519, n18520, n18521, n18522,
         n18523, n18524, n18525, n18526, n18527, n18528, n18529, n18530,
         n18531, n18532, n18533, n18534, n18535, n18536, n18537, n18538,
         n18539, n18540, n18541, n18542, n18543, n18544, n18545, n18546,
         n18547, n18548, n18549, n18550, n18551, n18552, n18553, n18554,
         n18555, n18556, n18557, n18558, n18559, n18560, n18561, n18562,
         n18563, n18564, n18565, n18566, n18567, n18568, n18569, n18570,
         n18571, n18572, n18573, n18574, n18575, n18576, n18577, n18578,
         n18579, n18580, n18581, n18582, n18583, n18584, n18585, n18586,
         n18587, n18588, n18589, n18590, n18591, n18592, n18593, n18594,
         n18595, n18596, n18597, n18598, n18599, n18600, n18601, n18602,
         n18603, n18604, n18605, n18606, n18607, n18608, n18609, n18610,
         n18611, n18612, n18613, n18614, n18615, n18616, n18617, n18618,
         n18619, n18620, n18621, n18622, n18623, n18624, n18625, n18626,
         n18627, n18628, n18629, n18630, n18631, n18632, n18633, n18634,
         n18635, n18636, n18637, n18638, n18639, n18640, n18641, n18642,
         n18643, n18644, n18645, n18646, n18647, n18648, n18649, n18650,
         n18651, n18652, n18653, n18654, n18655, n18656, n18657, n18658,
         n18659, n18660, n18661, n18662, n18663, n18664, n18665, n18666,
         n18667, n18668, n18669, n18670, n18671, n18672, n18673, n18674,
         n18675, n18676, n18677, n18678, n18679, n18680, n18681, n18682,
         n18683, n18684, n18685, n18686, n18687, n18688, n18689, n18690,
         n18691, n18692, n18693, n18694, n18695, n18696, n18697, n18698,
         n18699, n18700, n18701, n18702, n18703, n18704, n18705, n18706,
         n18707, n18708, n18709, n18710, n18711, n18712, n18713, n18714,
         n18715, n18716, n18717, n18718, n18719, n18720, n18721, n18722,
         n18723, n18724, n18725, n18726, n18727, n18728, n18729, n18730,
         n18731, n18732, n18733, n18734, n18735, n18736, n18737, n18738,
         n18739, n18740, n18741, n18742, n18743, n18744, n18745, n18746,
         n18747, n18748, n18749, n18750, n18751, n18752, n18753, n18754,
         n18755, n18756, n18757, n18758, n18759, n18760, n18761, n18762,
         n18763, n18764, n18765, n18766, n18767, n18768, n18769, n18770,
         n18771, n18772, n18773, n18774, n18775, n18776, n18777, n18778,
         n18779, n18780, n18781, n18782, n18783, n18784, n18785, n18786,
         n18787, n18788, n18789, n18790, n18791, n18792, n18793, n18794,
         n18795, n18796, n18797, n18798, n18799, n18800, n18801, n18802,
         n18803, n18804, n18805, n18806, n18807, n18808, n18809, n18810,
         n18811, n18812, n18813, n18814, n18815, n18816, n18817, n18818,
         n18819, n18820, n18821, n18822, n18823, n18824, n18825, n18826,
         n18827, n18828, n18829, n18830, n18831, n18832, n18833, n18834,
         n18835, n18836, n18837, n18838, n18839, n18840, n18841, n18842,
         n18843, n18844, n18845, n18846, n18847, n18848, n18849, n18850,
         n18851, n18852, n18853, n18854, n18855, n18856, n18857, n18858,
         n18859, n18860, n18861, n18862, n18863, n18864, n18865, n18866,
         n18867, n18868, n18869, n18870, n18871, n18872, n18873, n18874,
         n18875, n18876, n18877, n18878, n18879, n18880, n18881, n18882,
         n18883, n18884, n18885, n18886, n18887, n18888, n18889, n18890,
         n18891, n18892, n18893, n18894, n18895, n18896, n18897, n18898,
         n18899, n18900, n18901, n18902, n18903, n18904, n18905, n18906,
         n18907, n18908, n18909, n18910, n18911, n18912, n18913, n18914,
         n18915, n18916, n18917, n18918, n18919, n18920, n18921, n18922,
         n18923, n18924, n18925, n18926, n18927, n18928, n18929, n18930,
         n18931, n18932, n18933, n18934, n18935, n18936, n18937, n18938,
         n18939, n18940, n18941, n18942, n18943, n18944, n18945, n18946,
         n18947, n18948, n18949, n18950, n18951, n18952, n18953, n18954,
         n18955, n18956, n18957, n18958, n18959, n18960, n18961, n18962,
         n18963, n18964, n18965, n18966, n18967, n18968, n18969, n18970,
         n18971, n18972, n18973, n18974, n18975, n18976, n18977, n18978,
         n18979, n18980, n18981, n18982, n18983, n18984, n18985, n18986,
         n18987, n18988, n18989, n18990, n18991, n18992, n18993, n18994,
         n18995, n18996, n18997, n18998, n18999, n19000, n19001, n19002,
         n19003, n19004, n19005, n19006, n19007, n19008, n19009, n19010,
         n19011, n19012, n19013, n19014, n19015, n19016, n19017, n19018,
         n19019, n19020, n19021, n19022, n19023, n19024, n19025, n19026,
         n19027, n19028, n19029, n19030, n19031, n19032, n19033, n19034,
         n19035, n19036, n19037, n19038, n19039, n19040, n19041, n19042,
         n19043, n19044, n19045, n19046, n19047, n19048, n19049, n19050,
         n19051, n19052, n19053, n19054, n19055, n19056, n19057, n19058,
         n19059, n19060, n19061, n19062, n19063, n19064, n19065, n19066,
         n19067, n19068, n19069, n19070, n19071, n19072, n19073, n19074,
         n19075, n19076, n19077, n19078, n19079, n19080, n19081, n19082,
         n19083, n19084, n19085, n19086, n19087, n19088, n19089, n19090,
         n19091, n19092, n19093, n19094, n19095, n19096, n19097, n19098,
         n19099, n19100, n19101, n19102, n19103, n19104, n19105, n19106,
         n19107, n19108, n19109, n19110, n19111, n19112, n19113, n19114,
         n19115, n19116, n19117, n19118, n19119, n19120, n19121, n19122,
         n19123, n19124, n19125, n19126, n19127, n19128, n19129, n19130,
         n19131, n19132, n19133, n19134, n19135, n19136, n19137, n19138,
         n19139, n19140, n19141, n19142, n19143, n19144, n19145, n19146,
         n19147, n19148, n19149, n19150, n19151, n19152, n19153, n19154,
         n19155, n19156, n19157, n19158, n19159, n19160, n19161, n19162,
         n19163, n19164, n19165, n19166, n19167, n19168, n19169, n19170,
         n19171, n19172, n19173, n19174, n19175, n19176, n19177, n19178,
         n19179, n19180, n19181, n19182, n19183, n19184, n19185, n19186,
         n19187, n19188, n19189, n19190, n19191, n19192, n19193, n19194,
         n19195, n19196, n19197, n19198, n19199, n19200, n19201, n19202,
         n19203, n19204, n19205, n19206, n19207, n19208, n19209, n19210,
         n19211, n19212, n19213, n19214, n19215, n19216, n19217, n19218,
         n19219, n19220, n19221, n19222, n19223, n19224, n19225, n19226,
         n19227, n19228, n19229, n19230, n19231, n19232, n19233, n19234,
         n19235, n19236, n19237, n19238, n19239, n19240, n19241, n19242,
         n19243, n19244, n19245, n19246, n19247, n19248, n19249, n19250,
         n19251, n19252, n19253, n19254, n19255, n19256, n19257, n19258,
         n19259, n19260, n19261, n19262, n19263, n19264, n19265, n19266,
         n19267, n19268, n19269, n19270, n19271, n19272, n19273, n19274,
         n19275, n19276, n19277, n19278, n19279, n19280, n19281, n19282,
         n19283, n19284, n19285, n19286, n19287, n19288, n19289, n19290,
         n19291, n19292, n19293, n19294, n19295, n19296, n19297, n19298,
         n19299, n19300, n19301, n19302, n19303, n19304, n19305, n19306,
         n19307, n19308, n19309, n19310, n19311, n19312, n19313, n19314,
         n19315, n19316, n19317, n19318, n19319, n19320, n19321, n19322,
         n19323, n19324, n19325, n19326, n19327, n19328, n19329, n19330,
         n19331, n19332, n19333, n19334, n19335, n19336, n19337, n19338,
         n19339, n19340, n19341, n19342, n19343, n19344, n19345, n19346,
         n19347, n19348, n19349, n19350, n19351, n19352, n19353, n19354,
         n19355, n19356, n19357, n19358, n19359, n19360, n19361, n19362,
         n19363, n19364, n19365, n19366, n19367, n19368, n19369, n19370,
         n19371, n19372, n19373, n19374, n19375, n19376, n19377, n19378,
         n19379, n19380, n19381, n19382, n19383, n19384, n19385, n19386,
         n19387, n19388, n19389, n19390, n19391, n19392, n19393, n19394,
         n19395, n19396, n19397, n19398, n19399, n19400, n19401, n19402,
         n19403, n19404, n19405, n19406, n19407, n19408, n19409, n19410,
         n19411, n19412, n19413, n19414, n19415, n19416, n19417, n19418,
         n19419, n19420, n19421, n19422, n19423, n19424, n19425, n19426,
         n19427, n19428, n19429, n19430, n19431, n19432, n19433, n19434,
         n19435, n19436, n19437, n19438, n19439, n19440, n19441, n19442,
         n19443, n19444, n19445, n19446, n19447, n19448, n19449, n19450,
         n19451, n19452, n19453, n19454, n19455, n19456, n19457, n19458,
         n19459, n19460, n19461, n19462, n19463, n19464, n19465, n19466,
         n19467, n19468, n19469, n19470, n19471, n19472, n19473, n19474,
         n19475, n19476, n19477, n19478, n19479, n19480, n19481, n19482,
         n19483, n19484, n19485, n19486, n19487, n19488, n19489, n19490,
         n19491, n19492, n19493, n19494, n19495, n19496, n19497, n19498,
         n19499, n19500, n19501, n19502, n19503, n19504, n19505, n19506,
         n19507, n19508, n19509, n19510, n19511, n19512, n19513, n19514,
         n19515, n19516, n19517, n19518, n19519, n19520, n19521, n19522,
         n19523, n19524, n19525, n19526, n19527, n19528, n19529, n19530,
         n19531, n19532, n19533, n19534, n19535, n19536, n19537, n19538,
         n19539, n19540, n19541, n19542, n19543, n19544, n19545, n19546,
         n19547, n19548, n19549, n19550, n19551, n19552, n19553, n19554,
         n19555, n19556, n19557, n19558, n19559, n19560, n19561, n19562,
         n19563, n19564, n19565, n19566, n19567, n19568, n19569, n19570,
         n19571, n19572, n19573, n19574, n19575, n19576, n19577, n19578,
         n19579, n19580, n19581, n19582, n19583, n19584, n19585, n19586,
         n19587, n19588, n19589, n19590, n19591, n19592, n19593, n19594,
         n19595, n19596, n19597, n19598, n19599, n19600, n19601, n19602,
         n19603, n19604, n19605, n19606, n19607, n19608, n19609, n19610,
         n19611, n19612, n19613, n19614, n19615, n19616, n19617, n19618,
         n19619, n19620, n19621, n19622, n19623, n19624, n19625, n19626,
         n19627, n19628, n19629, n19630, n19631, n19632, n19633, n19634,
         n19635, n19636, n19637, n19638, n19639, n19640, n19641, n19642,
         n19643, n19644, n19645, n19646, n19647, n19648, n19649, n19650,
         n19651, n19652, n19653, n19654, n19655, n19656, n19657, n19658,
         n19659, n19660, n19661, n19662, n19663, n19664, n19665, n19666,
         n19667, n19668, n19669, n19670, n19671, n19672, n19673, n19674,
         n19675, n19676, n19677, n19678, n19679, n19680, n19681, n19682,
         n19683, n19684, n19685, n19686, n19687, n19688, n19689, n19690,
         n19691, n19692, n19693, n19694, n19695, n19696, n19697, n19698,
         n19699, n19700, n19701, n19702, n19703, n19704, n19705, n19706,
         n19707, n19708, n19709, n19710, n19711, n19712, n19713, n19714,
         n19715, n19716, n19717, n19718, n19719, n19720, n19721, n19722,
         n19723, n19724, n19725, n19726, n19727, n19728, n19729, n19730,
         n19731, n19732, n19733, n19734, n19735, n19736, n19737, n19738,
         n19739, n19740, n19741, n19742, n19743, n19744, n19745, n19746,
         n19747, n19748, n19749, n19750, n19751, n19752, n19753, n19754,
         n19755, n19756, n19757, n19758, n19759, n19760, n19761, n19762,
         n19763, n19764, n19765, n19766, n19767, n19768, n19769, n19770,
         n19771, n19772, n19773, n19774, n19775, n19776, n19777, n19778,
         n19779, n19780, n19781, n19782, n19783, n19784, n19785, n19786,
         n19787, n19788, n19789, n19790, n19791, n19792, n19793, n19794,
         n19795, n19796, n19797, n19798, n19799, n19800, n19801, n19802,
         n19803, n19804, n19805, n19806, n19807, n19808, n19809, n19810,
         n19811, n19812, n19813, n19814, n19815, n19816, n19817, n19818,
         n19819, n19820, n19821, n19822, n19823, n19824, n19825, n19826,
         n19827, n19828, n19829, n19830, n19831, n19832, n19833, n19834,
         n19835, n19836, n19837, n19838, n19839, n19840, n19841, n19842,
         n19843, n19844, n19845, n19846, n19847, n19848, n19849, n19850,
         n19851, n19852, n19853, n19854, n19855, n19856, n19857, n19858,
         n19859, n19860, n19861, n19862, n19863, n19864, n19865, n19866,
         n19867, n19868, n19869, n19870, n19871, n19872, n19873, n19874,
         n19875, n19876, n19877, n19878, n19879, n19880, n19881, n19882,
         n19883, n19884, n19885, n19886, n19887, n19888, n19889, n19890,
         n19891, n19892, n19893, n19894, n19895, n19896, n19897, n19898,
         n19899, n19900, n19901, n19902, n19903, n19904, n19905, n19906,
         n19907, n19908, n19909, n19910, n19911, n19912, n19913, n19914,
         n19915, n19916, n19917, n19918, n19919, n19920, n19921, n19922,
         n19923, n19924, n19925, n19926, n19927, n19928, n19929, n19930,
         n19931, n19932, n19933, n19934, n19935, n19936, n19937, n19938,
         n19939, n19940, n19941, n19942, n19943, n19944, n19945, n19946,
         n19947, n19948, n19949, n19950, n19951, n19952, n19953, n19954,
         n19955, n19956, n19957, n19958, n19959, n19960, n19961, n19962,
         n19963, n19964, n19965, n19966, n19967, n19968, n19969, n19970,
         n19971, n19972, n19973, n19974, n19975, n19976, n19977, n19978,
         n19979, n19980, n19981, n19982, n19983, n19984, n19985, n19986,
         n19987, n19988, n19989, n19990, n19991, n19992, n19993, n19994,
         n19995, n19996, n19997, n19998, n19999, n20000, n20001, n20002,
         n20003, n20004, n20005, n20006, n20007, n20008, n20009, n20010,
         n20011, n20012, n20013, n20014, n20015, n20016, n20017, n20018,
         n20019, n20020, n20021, n20022, n20023, n20024, n20025, n20026,
         n20027, n20028, n20029, n20030, n20031, n20032, n20033, n20034,
         n20035, n20036, n20037, n20038, n20039, n20040, n20041, n20042,
         n20043, n20044, n20045, n20046, n20047, n20048, n20049, n20050,
         n20051, n20052, n20053, n20054, n20055, n20056, n20057, n20058,
         n20059, n20060, n20061, n20062, n20063, n20064, n20065, n20066,
         n20067, n20068, n20069, n20070, n20071, n20072, n20073, n20074,
         n20075, n20076, n20077, n20078, n20079, n20080, n20081, n20082,
         n20083, n20084, n20085, n20086, n20087, n20088, n20089, n20090,
         n20091, n20092, n20093, n20094, n20095, n20096, n20097, n20098,
         n20099, n20100, n20101, n20102, n20103, n20104, n20105, n20106,
         n20107, n20108, n20109, n20110, n20111, n20112, n20113, n20114,
         n20115, n20116, n20117, n20118, n20119, n20120, n20121, n20122,
         n20123, n20124, n20125, n20126, n20127, n20128, n20129, n20130,
         n20131, n20132, n20133, n20134, n20135, n20136, n20137, n20138,
         n20139, n20140, n20141, n20142, n20143, n20144, n20145, n20146,
         n20147, n20148, n20149, n20150, n20151, n20152, n20153, n20154,
         n20155, n20156, n20157, n20158, n20159, n20160, n20161, n20162,
         n20163, n20164, n20165, n20166, n20167, n20168, n20169, n20170,
         n20171, n20172, n20173, n20174, n20175, n20176, n20177, n20178,
         n20179, n20180, n20181, n20182, n20183, n20184, n20185, n20186,
         n20187, n20188, n20189, n20190, n20191, n20192, n20193, n20194,
         n20195, n20196, n20197, n20198, n20199, n20200, n20201, n20202,
         n20203, n20204, n20205, n20206, n20207, n20208, n20209, n20210,
         n20211, n20212, n20213, n20214, n20215, n20216, n20217, n20218,
         n20219, n20220, n20221, n20222, n20223, n20224, n20225, n20226,
         n20227, n20228, n20229, n20230, n20231, n20232, n20233, n20234,
         n20235, n20236, n20237, n20238, n20239, n20240, n20241, n20242,
         n20243, n20244, n20245, n20246, n20247, n20248, n20249, n20250,
         n20251, n20252, n20253, n20254, n20255, n20256, n20257, n20258,
         n20259, n20260, n20261, n20262, n20263, n20264, n20265, n20266,
         n20267, n20268, n20269, n20270, n20271, n20272, n20273, n20274,
         n20275, n20276, n20277, n20278, n20279, n20280, n20281, n20282,
         n20283, n20284, n20285, n20286, n20287, n20288, n20289, n20290,
         n20291, n20292, n20293, n20294, n20295, n20296, n20297, n20298,
         n20299, n20300, n20301, n20302, n20303, n20304, n20305, n20306,
         n20307, n20308, n20309, n20310, n20311, n20312, n20313, n20314,
         n20315, n20316, n20317, n20318, n20319, n20320, n20321, n20322,
         n20323, n20324, n20325, n20326, n20327, n20328, n20329, n20330,
         n20331, n20332, n20333, n20334, n20335, n20336, n20337, n20338,
         n20339, n20340, n20341, n20342, n20343, n20344, n20345, n20346,
         n20347, n20348, n20349, n20350, n20351, n20352, n20353, n20354,
         n20355, n20356, n20357, n20358, n20359, n20360, n20361, n20362,
         n20363, n20364, n20365, n20366, n20367, n20368, n20369, n20370,
         n20371, n20372, n20373, n20374, n20375, n20376, n20377, n20378,
         n20379, n20380, n20381, n20382, n20383, n20384, n20385, n20386,
         n20387, n20388, n20389, n20390, n20391, n20392, n20393, n20394,
         n20395, n20396, n20397, n20398, n20399, n20400, n20401, n20402,
         n20403, n20404, n20405, n20406, n20407, n20408, n20409, n20410,
         n20411, n20412, n20413, n20414, n20415, n20416, n20417, n20418,
         n20419, n20420, n20421, n20422, n20423, n20424, n20425, n20426,
         n20427, n20428, n20429, n20430, n20431, n20432, n20433, n20434,
         n20435, n20436, n20437, n20438, n20439, n20440, n20441, n20442,
         n20443, n20444, n20445, n20446, n20447, n20448, n20449, n20450,
         n20451, n20452, n20453, n20454, n20455, n20456, n20457, n20458,
         n20459, n20460, n20461, n20462, n20463, n20464, n20465, n20466,
         n20467, n20468, n20469, n20470, n20471, n20472, n20473, n20474,
         n20475, n20476, n20477, n20478, n20479, n20480, n20481, n20482,
         n20483, n20484, n20485, n20486, n20487, n20488, n20489, n20490,
         n20491, n20492, n20493, n20494, n20495, n20496, n20497, n20498,
         n20499, n20500, n20501, n20502, n20503, n20504, n20505, n20506,
         n20507, n20508, n20509, n20510, n20511, n20512, n20513, n20514,
         n20515, n20516, n20517, n20518, n20519, n20520, n20521, n20522,
         n20523, n20524, n20525, n20526, n20527, n20528, n20529, n20530,
         n20531, n20532, n20533, n20534, n20535, n20536, n20537, n20538,
         n20539, n20540, n20541, n20542, n20543, n20544, n20545, n20546,
         n20547, n20548, n20549, n20550, n20551, n20552, n20553, n20554,
         n20555, n20556, n20557, n20558, n20559, n20560, n20561, n20562,
         n20563, n20564, n20565, n20566, n20567, n20568, n20569, n20570,
         n20571, n20572, n20573, n20574, n20575, n20576, n20577, n20578,
         n20579, n20580, n20581, n20582, n20583, n20584, n20585, n20586,
         n20587, n20588, n20589, n20590, n20591, n20592, n20593, n20594,
         n20595, n20596, n20597, n20598, n20599, n20600, n20601, n20602,
         n20603, n20604, n20605, n20606, n20607, n20608, n20609, n20610,
         n20611, n20612, n20613, n20614, n20615, n20616, n20617, n20618,
         n20619, n20620, n20621, n20622, n20623, n20624, n20625, n20626,
         n20627, n20628, n20629, n20630, n20631, n20632, n20633, n20634,
         n20635, n20636, n20637, n20638, n20639, n20640, n20641, n20642,
         n20643, n20644, n20645, n20646, n20647, n20648, n20649, n20650,
         n20651, n20652, n20653, n20654, n20655, n20656, n20657, n20658,
         n20659, n20660, n20661, n20662, n20663, n20664, n20665, n20666,
         n20667, n20668, n20669, n20670, n20671, n20672, n20673, n20674,
         n20675, n20676, n20677, n20678, n20679, n20680, n20681, n20682,
         n20683, n20684, n20685, n20686, n20687, n20688, n20689, n20690,
         n20691, n20692, n20693, n20694, n20695, n20696, n20697, n20698,
         n20699, n20700, n20701, n20702, n20703, n20704, n20705, n20706,
         n20707, n20708, n20709, n20710, n20711, n20712, n20713, n20714,
         n20715, n20716, n20717, n20718, n20719, n20720, n20721, n20722,
         n20723, n20724, n20725, n20726, n20727, n20728, n20729, n20730,
         n20731, n20732, n20733, n20734, n20735, n20736, n20737, n20738,
         n20739, n20740, n20741, n20742, n20743, n20744, n20745, n20746,
         n20747, n20748, n20749, n20750, n20751, n20752, n20753, n20754,
         n20755, n20756, n20757, n20758, n20759, n20760, n20761, n20762,
         n20763, n20764, n20765, n20766, n20767, n20768, n20769, n20770,
         n20771, n20772, n20773, n20774, n20775, n20776, n20777, n20778,
         n20779, n20780, n20781, n20782, n20783, n20784, n20785, n20786,
         n20787, n20788, n20789, n20790, n20791, n20792, n20793, n20794,
         n20795, n20796, n20797, n20798, n20799, n20800, n20801, n20802,
         n20803, n20804, n20805, n20806, n20807, n20808, n20809, n20810,
         n20811, n20812, n20813, n20814, n20815, n20816, n20817, n20818,
         n20819, n20820, n20821, n20822, n20823, n20824, n20825, n20826,
         n20827, n20828, n20829, n20830, n20831, n20832, n20833, n20834,
         n20835, n20836, n20837, n20838, n20839, n20840, n20841, n20842,
         n20843, n20844, n20845, n20846, n20847, n20848, n20849, n20850,
         n20851, n20852, n20853, n20854, n20855, n20856, n20857, n20858,
         n20859, n20860, n20861, n20862, n20863, n20864, n20865, n20866,
         n20867, n20868, n20869, n20870, n20871, n20872, n20873, n20874,
         n20875, n20876, n20877, n20878, n20879, n20880, n20881, n20882,
         n20883, n20884, n20885, n20886, n20887, n20888, n20889, n20890,
         n20891, n20892, n20893, n20894, n20895, n20896, n20897, n20898,
         n20899, n20900, n20901, n20902, n20903, n20904, n20905, n20906,
         n20907, n20908, n20909, n20910, n20911, n20912, n20913, n20914,
         n20915, n20916, n20917, n20918, n20919, n20920, n20921, n20922,
         n20923, n20924, n20925, n20926, n20927, n20928, n20929, n20930,
         n20931, n20932, n20933, n20934, n20935, n20936, n20937, n20938,
         n20939, n20940, n20941, n20942, n20943, n20944, n20945, n20946,
         n20947, n20948, n20949, n20950, n20951, n20952, n20953, n20954,
         n20955, n20956, n20957, n20958, n20959, n20960, n20961, n20962,
         n20963, n20964, n20965, n20966, n20967, n20968, n20969, n20970,
         n20971, n20972, n20973, n20974, n20975, n20976, n20977, n20978,
         n20979, n20980, n20981, n20982, n20983, n20984, n20985, n20986,
         n20987, n20988, n20989, n20990, n20991, n20992, n20993, n20994,
         n20995, n20996, n20997, n20998, n20999, n21000, n21001, n21002,
         n21003, n21004, n21005, n21006, n21007, n21008, n21009, n21010,
         n21011, n21012, n21013, n21014, n21015, n21016, n21017, n21018,
         n21019, n21020, n21021, n21022, n21023, n21024, n21025, n21026,
         n21027, n21028, n21029, n21030, n21031, n21032, n21033, n21034,
         n21035, n21036, n21037, n21038, n21039, n21040, n21041, n21042,
         n21043, n21044, n21045, n21046, n21047, n21048, n21049, n21050,
         n21051, n21052, n21053, n21054, n21055, n21056, n21057, n21058,
         n21059, n21060, n21061, n21062, n21063, n21064, n21065, n21066,
         n21067, n21068, n21069, n21070, n21071, n21072, n21073, n21074,
         n21075, n21076, n21077, n21078, n21079, n21080, n21081, n21082,
         n21083, n21084, n21085, n21086, n21087, n21088, n21089, n21090,
         n21091, n21092, n21093, n21094, n21095, n21096, n21097, n21098,
         n21099, n21100, n21101, n21102, n21103, n21104, n21105, n21106,
         n21107, n21108, n21109, n21110, n21111, n21112, n21113, n21114,
         n21115, n21116, n21117, n21118, n21119, n21120, n21121, n21122,
         n21123, n21124, n21125, n21126, n21127, n21128, n21129, n21130,
         n21131, n21132, n21133, n21134, n21135, n21136, n21137, n21138,
         n21139, n21140, n21141, n21142, n21143, n21144, n21145, n21146,
         n21147, n21148, n21149, n21150, n21151, n21152, n21153, n21154,
         n21155, n21156, n21157, n21158, n21159, n21160, n21161, n21162,
         n21163, n21164, n21165, n21166, n21167, n21168, n21169, n21170,
         n21171, n21172, n21173, n21174, n21175, n21176, n21177, n21178,
         n21179, n21180, n21181, n21182, n21183, n21184, n21185, n21186,
         n21187, n21188, n21189, n21190, n21191, n21192, n21193, n21194,
         n21195, n21196, n21197, n21198, n21199, n21200, n21201, n21202,
         n21203, n21204, n21205, n21206, n21207, n21208, n21209, n21210,
         n21211, n21212, n21213, n21214, n21215, n21216, n21217, n21218,
         n21219, n21220, n21221, n21222, n21223, n21224, n21225, n21226,
         n21227, n21228, n21229, n21230, n21231, n21232, n21233, n21234,
         n21235, n21236, n21237, n21238, n21239, n21240, n21241, n21242,
         n21243, n21244, n21245, n21246, n21247, n21248, n21249, n21250,
         n21251, n21252, n21253, n21254, n21255, n21256, n21257, n21258,
         n21259, n21260, n21261, n21262, n21263, n21264, n21265, n21266,
         n21267, n21268, n21269, n21270, n21271, n21272, n21273, n21274,
         n21275, n21276, n21277, n21278, n21279, n21280, n21281, n21282,
         n21283, n21284, n21285, n21286, n21287, n21288, n21289, n21290,
         n21291, n21292, n21293, n21294, n21295, n21296, n21297, n21298,
         n21299, n21300, n21301, n21302, n21303, n21304, n21305, n21306,
         n21307, n21308, n21309, n21310, n21311, n21312, n21313, n21314,
         n21315, n21316, n21317, n21318, n21319, n21320, n21321, n21322,
         n21323, n21324, n21325, n21326, n21327, n21328, n21329, n21330,
         n21331, n21332, n21333, n21334, n21335, n21336, n21337, n21338,
         n21339, n21340, n21341, n21342, n21343, n21344, n21345, n21346,
         n21347, n21348, n21349, n21350, n21351, n21352, n21353, n21354,
         n21355, n21356, n21357, n21358, n21359, n21360, n21361, n21362,
         n21363, n21364, n21365, n21366, n21367, n21368, n21369, n21370,
         n21371, n21372, n21373, n21374, n21375, n21376, n21377, n21378,
         n21379, n21380, n21381, n21382, n21383, n21384, n21385, n21386,
         n21387, n21388, n21389, n21390, n21391, n21392, n21393, n21394,
         n21395, n21396, n21397, n21398, n21399, n21400, n21401, n21402,
         n21403, n21404, n21405, n21406, n21407, n21408, n21409, n21410,
         n21411, n21412, n21413, n21414, n21415, n21416, n21417, n21418,
         n21419, n21420, n21421, n21422, n21423, n21424, n21425, n21426,
         n21427, n21428, n21429, n21430, n21431, n21432, n21433, n21434,
         n21435, n21436, n21437, n21438, n21439, n21440, n21441, n21442,
         n21443, n21444, n21445, n21446, n21447, n21448, n21449, n21450,
         n21451, n21452, n21453, n21454, n21455, n21456, n21457, n21458,
         n21459, n21460, n21461, n21462, n21463, n21464, n21465, n21466,
         n21467, n21468, n21469, n21470, n21471, n21472, n21473, n21474,
         n21475, n21476, n21477, n21478, n21479, n21480, n21481, n21482,
         n21483, n21484, n21485, n21486, n21487, n21488, n21489, n21490,
         n21491, n21492, n21493, n21494, n21495, n21496, n21497, n21498,
         n21499, n21500, n21501, n21502, n21503, n21504, n21505, n21506,
         n21507, n21508, n21509, n21510, n21511, n21512, n21513, n21514,
         n21515, n21516, n21517, n21518, n21519, n21520, n21521, n21522,
         n21523, n21524, n21525, n21526, n21527, n21528, n21529, n21530,
         n21531, n21532, n21533, n21534, n21535, n21536, n21537, n21538,
         n21539, n21540, n21541, n21542, n21543, n21544, n21545, n21546,
         n21547, n21548, n21549, n21550, n21551, n21552, n21553, n21554,
         n21555, n21556, n21557, n21558, n21559, n21560, n21561, n21562,
         n21563, n21564, n21565, n21566, n21567, n21568, n21569, n21570,
         n21571, n21572, n21573, n21574, n21575, n21576, n21577, n21578,
         n21579, n21580, n21581, n21582, n21583, n21584, n21585, n21586,
         n21587, n21588, n21589, n21590, n21591, n21592, n21593, n21594,
         n21595, n21596, n21597, n21598, n21599, n21600, n21601, n21602,
         n21603, n21604, n21605, n21606, n21607, n21608, n21609, n21610,
         n21611, n21612, n21613, n21614, n21615, n21616, n21617, n21618,
         n21619, n21620, n21621, n21622, n21623, n21624, n21625, n21626,
         n21627, n21628, n21629, n21630, n21631, n21632, n21633, n21634,
         n21635, n21636, n21637, n21638, n21639, n21640, n21641, n21642,
         n21643, n21644, n21645, n21646, n21647, n21648, n21649, n21650,
         n21651, n21652, n21653, n21654, n21655, n21656, n21657, n21658,
         n21659, n21660, n21661, n21662, n21663, n21664, n21665, n21666,
         n21667, n21668, n21669, n21670, n21671, n21672, n21673, n21674,
         n21675, n21676, n21677, n21678, n21679, n21680, n21681, n21682,
         n21683, n21684, n21685, n21686, n21687, n21688, n21689, n21690,
         n21691, n21692, n21693, n21694, n21695, n21696, n21697, n21698,
         n21699, n21700, n21701, n21702, n21703, n21704, n21705, n21706,
         n21707, n21708, n21709, n21710, n21711, n21712, n21713, n21714,
         n21715, n21716, n21717, n21718, n21719, n21720, n21721, n21722,
         n21723, n21724, n21725, n21726, n21727, n21728, n21729, n21730,
         n21731, n21732, n21733, n21734, n21735, n21736, n21737, n21738,
         n21739, n21740, n21741, n21742, n21743, n21744, n21745, n21746,
         n21747, n21748, n21749, n21750, n21751, n21752, n21753, n21754,
         n21755, n21756, n21757, n21758, n21759, n21760, n21761, n21762,
         n21763, n21764, n21765, n21766, n21767, n21768, n21769, n21770,
         n21771, n21772, n21773, n21774, n21775, n21776, n21777, n21778,
         n21779, n21780, n21781, n21782, n21783, n21784, n21785, n21786,
         n21787, n21788, n21789, n21790, n21791, n21792, n21793, n21794,
         n21795, n21796, n21797, n21798, n21799, n21800, n21801, n21802,
         n21803, n21804, n21805, n21806, n21807, n21808, n21809, n21810,
         n21811, n21812, n21813, n21814, n21815, n21816, n21817, n21818,
         n21819, n21820, n21821, n21822, n21823, n21824, n21825, n21826,
         n21827, n21828, n21829, n21830, n21831, n21832, n21833, n21834,
         n21835, n21836, n21837, n21838, n21839, n21840, n21841, n21842,
         n21843, n21844, n21845, n21846, n21847, n21848, n21849, n21850,
         n21851, n21852, n21853, n21854, n21855, n21856, n21857, n21858,
         n21859, n21860, n21861, n21862, n21863, n21864, n21865, n21866,
         n21867, n21868, n21869, n21870, n21871, n21872, n21873, n21874,
         n21875, n21876, n21877, n21878, n21879, n21880, n21881, n21882,
         n21883, n21884, n21885, n21886, n21887, n21888, n21889, n21890,
         n21891, n21892, n21893, n21894, n21895, n21896, n21897, n21898,
         n21899, n21900, n21901, n21902, n21903, n21904, n21905, n21906,
         n21907, n21908, n21909, n21910, n21911, n21912, n21913, n21914,
         n21915, n21916, n21917, n21918, n21919, n21920, n21921, n21922,
         n21923, n21924, n21925, n21926, n21927, n21928, n21929, n21930,
         n21931, n21932, n21933, n21934, n21935, n21936, n21937, n21938,
         n21939, n21940, n21941, n21942, n21943, n21944, n21945, n21946,
         n21947, n21948, n21949, n21950, n21951, n21952, n21953, n21954,
         n21955, n21956, n21957, n21958, n21959, n21960, n21961, n21962,
         n21963, n21964, n21965, n21966, n21967, n21968, n21969, n21970,
         n21971, n21972, n21973, n21974, n21975, n21976, n21977, n21978,
         n21979, n21980, n21981, n21982, n21983, n21984, n21985, n21986,
         n21987, n21988, n21989, n21990, n21991, n21992, n21993, n21994,
         n21995, n21996, n21997, n21998, n21999, n22000, n22001, n22002,
         n22003, n22004, n22005, n22006, n22007, n22008, n22009, n22010,
         n22011, n22012, n22013, n22014, n22015, n22016, n22017, n22018,
         n22019, n22020, n22021, n22022, n22023, n22024, n22025, n22026,
         n22027, n22028, n22029, n22030, n22031, n22032, n22033, n22034,
         n22035, n22036, n22037, n22038, n22039, n22040, n22041, n22042,
         n22043, n22044, n22045, n22046, n22047, n22048, n22049, n22050,
         n22051, n22052, n22053, n22054, n22055, n22056, n22057, n22058,
         n22059, n22060, n22061, n22062, n22063, n22064, n22065, n22066,
         n22067, n22068, n22069, n22070, n22071, n22072, n22073, n22074,
         n22075, n22076, n22077, n22078, n22079, n22080, n22081, n22082,
         n22083, n22084, n22085, n22086, n22087, n22088, n22089, n22090,
         n22091, n22092, n22093, n22094, n22095, n22096, n22097, n22098,
         n22099, n22100, n22101, n22102, n22103, n22104, n22105, n22106,
         n22107, n22108, n22109, n22110, n22111, n22112, n22113, n22114,
         n22115, n22116, n22117, n22118, n22119, n22120, n22121, n22122,
         n22123, n22124, n22125, n22126, n22127, n22128, n22129, n22130,
         n22131, n22132, n22133, n22134, n22135, n22136, n22137, n22138,
         n22139, n22140, n22141, n22142, n22143, n22144, n22145, n22146,
         n22147, n22148, n22149, n22150, n22151, n22152, n22153, n22154,
         n22155, n22156, n22157, n22158, n22159, n22160, n22161, n22162,
         n22163, n22164, n22165, n22166, n22167, n22168, n22169, n22170,
         n22171, n22172, n22173, n22174, n22175, n22176, n22177, n22178,
         n22179, n22180, n22181, n22182, n22183, n22184, n22185, n22186,
         n22187, n22188, n22189, n22190, n22191, n22192, n22193, n22194,
         n22195, n22196, n22197, n22198, n22199, n22200, n22201, n22202,
         n22203, n22204, n22205, n22206, n22207, n22208, n22209, n22210,
         n22211, n22212, n22213, n22214, n22215, n22216, n22217, n22218,
         n22219, n22220, n22221, n22222, n22223, n22224, n22225, n22226,
         n22227, n22228, n22229, n22230, n22231, n22232, n22233, n22234,
         n22235, n22236, n22237, n22238, n22239, n22240, n22241, n22242,
         n22243, n22244, n22245, n22246, n22247, n22248, n22249, n22250,
         n22251, n22252, n22253, n22254, n22255, n22256, n22257, n22258,
         n22259, n22260, n22261, n22262, n22263, n22264, n22265, n22266,
         n22267, n22268, n22269, n22270, n22271, n22272, n22273, n22274,
         n22275, n22276, n22277, n22278, n22279, n22280, n22281, n22282,
         n22283, n22284, n22285, n22286, n22287, n22288, n22289, n22290,
         n22291, n22292, n22293, n22294, n22295, n22296, n22297, n22298,
         n22299, n22300, n22301, n22302, n22303, n22304, n22305, n22306,
         n22307, n22308, n22309, n22310, n22311, n22312, n22313, n22314,
         n22315, n22316, n22317, n22318, n22319, n22320, n22321, n22322,
         n22323, n22324, n22325, n22326, n22327, n22328, n22329, n22330,
         n22331, n22332, n22333, n22334, n22335, n22336, n22337, n22338,
         n22339, n22340, n22341, n22342, n22343, n22344, n22345, n22346,
         n22347, n22348, n22349, n22350, n22351, n22352, n22353, n22354,
         n22355, n22356, n22357, n22358, n22359, n22360, n22361, n22362,
         n22363, n22364, n22365, n22366, n22367, n22368, n22369, n22370,
         n22371, n22372, n22373, n22374, n22375, n22376, n22377, n22378,
         n22379, n22380, n22381, n22382, n22383, n22384, n22385, n22386,
         n22387, n22388, n22389, n22390, n22391, n22392, n22393, n22394,
         n22395, n22396, n22397, n22398, n22399, n22400, n22401, n22402,
         n22403, n22404, n22405, n22406, n22407, n22408, n22409, n22410,
         n22411, n22412, n22413, n22414, n22415, n22416, n22417, n22418,
         n22419, n22420, n22421, n22422, n22423, n22424, n22425, n22426,
         n22427, n22428, n22429, n22430, n22431, n22432, n22433, n22434,
         n22435, n22436, n22437, n22438, n22439, n22440, n22441, n22442,
         n22443, n22444, n22445, n22446, n22447, n22448, n22449, n22450,
         n22451, n22452, n22453, n22454, n22455, n22456, n22457, n22458,
         n22459, n22460, n22461, n22462, n22463, n22464, n22465, n22466,
         n22467, n22468, n22469, n22470, n22471, n22472, n22473, n22474,
         n22475, n22476, n22477, n22478, n22479, n22480, n22481, n22482,
         n22483, n22484, n22485, n22486, n22487, n22488, n22489, n22490,
         n22491, n22492, n22493, n22494, n22495, n22496, n22497, n22498,
         n22499, n22500, n22501, n22502, n22503, n22504, n22505, n22506,
         n22507, n22508, n22509, n22510, n22511, n22512, n22513, n22514,
         n22515, n22516, n22517, n22518, n22519, n22520, n22521, n22522,
         n22523, n22524, n22525, n22526, n22527, n22528, n22529, n22530,
         n22531, n22532, n22533, n22534, n22535, n22536, n22537, n22538,
         n22539, n22540, n22541, n22542, n22543, n22544, n22545, n22546,
         n22547, n22548, n22549, n22550, n22551, n22552, n22553, n22554,
         n22555, n22556, n22557, n22558, n22559, n22560, n22561, n22562,
         n22563, n22564, n22565, n22566, n22567, n22568, n22569, n22570,
         n22571, n22572, n22573, n22574, n22575, n22576, n22577, n22578,
         n22579, n22580, n22581, n22582, n22583, n22584, n22585, n22586,
         n22587, n22588, n22589, n22590, n22591, n22592, n22593, n22594,
         n22595, n22596, n22597, n22598, n22599, n22600, n22601, n22602,
         n22603, n22604, n22605, n22606, n22607, n22608, n22609, n22610,
         n22611, n22612, n22613, n22614, n22615, n22616, n22617, n22618,
         n22619, n22620, n22621, n22622, n22623, n22624, n22625, n22626,
         n22627, n22628, n22629, n22630, n22631, n22632, n22633, n22634,
         n22635, n22636, n22637, n22638, n22639, n22640, n22641, n22642,
         n22643, n22644, n22645, n22646, n22647, n22648, n22649, n22650,
         n22651, n22652, n22653, n22654, n22655, n22656, n22657, n22658,
         n22659, n22660, n22661, n22662, n22663, n22664, n22665, n22666,
         n22667, n22668, n22669, n22670, n22671, n22672, n22673, n22674,
         n22675, n22676, n22677, n22678, n22679, n22680, n22681, n22682,
         n22683, n22684, n22685, n22686, n22687, n22688, n22689, n22690,
         n22691, n22692, n22693, n22694, n22695, n22696, n22697, n22698,
         n22699, n22700, n22701, n22702, n22703, n22704, n22705, n22706,
         n22707, n22708, n22709, n22710, n22711, n22712, n22713, n22714,
         n22715, n22716, n22717, n22718, n22719, n22720, n22721, n22722,
         n22723, n22724, n22725, n22726, n22727, n22728, n22729, n22730,
         n22731, n22732, n22733, n22734, n22735, n22736, n22737, n22738,
         n22739, n22740, n22741, n22742, n22743, n22744, n22745, n22746,
         n22747, n22748, n22749, n22750, n22751, n22752, n22753, n22754,
         n22755, n22756, n22757, n22758, n22759, n22760, n22761, n22762,
         n22763, n22764, n22765, n22766, n22767, n22768, n22769, n22770,
         n22771, n22772, n22773, n22774, n22775, n22776, n22777, n22778,
         n22779, n22780, n22781, n22782, n22783, n22784, n22785, n22786,
         n22787, n22788, n22789, n22790, n22791, n22792, n22793, n22794,
         n22795, n22796, n22797, n22798, n22799, n22800, n22801, n22802,
         n22803, n22804, n22805, n22806, n22807, n22808, n22809, n22810,
         n22811, n22812, n22813, n22814, n22815, n22816, n22817, n22818,
         n22819, n22820, n22821, n22822, n22823, n22824, n22825, n22826,
         n22827, n22828, n22829, n22830, n22831, n22832, n22833, n22834,
         n22835, n22836, n22837, n22838, n22839, n22840, n22841, n22842,
         n22843, n22844, n22845, n22846, n22847, n22848, n22849, n22850,
         n22851, n22852, n22853, n22854, n22855, n22856, n22857, n22858,
         n22859, n22860, n22861, n22862, n22863, n22864, n22865, n22866,
         n22867, n22868, n22869, n22870, n22871, n22872, n22873, n22874,
         n22875, n22876, n22877, n22878, n22879, n22880, n22881, n22882,
         n22883, n22884, n22885, n22886, n22887, n22888, n22889, n22890,
         n22891, n22892, n22893, n22894, n22895, n22896, n22897, n22898,
         n22899, n22900, n22901, n22902, n22903, n22904, n22905, n22906,
         n22907, n22908, n22909, n22910, n22911, n22912, n22913, n22914,
         n22915, n22916, n22917, n22918, n22919, n22920, n22921, n22922,
         n22923, n22924, n22925, n22926, n22927, n22928, n22929, n22930,
         n22931, n22932, n22933, n22934, n22935, n22936, n22937, n22938,
         n22939, n22940, n22941, n22942, n22943, n22944, n22945, n22946,
         n22947, n22948, n22949, n22950, n22951, n22952, n22953, n22954,
         n22955, n22956, n22957, n22958, n22959, n22960, n22961, n22962,
         n22963, n22964, n22965, n22966, n22967, n22968, n22969, n22970,
         n22971, n22972, n22973, n22974, n22975, n22976, n22977, n22978,
         n22979, n22980, n22981, n22982, n22983, n22984, n22985, n22986,
         n22987, n22988, n22989, n22990, n22991, n22992, n22993, n22994,
         n22995, n22996, n22997, n22998, n22999, n23000, n23001, n23002,
         n23003, n23004, n23005, n23006, n23007, n23008, n23009, n23010,
         n23011, n23012, n23013, n23014, n23015, n23016, n23017, n23018,
         n23019, n23020, n23021, n23022, n23023, n23024, n23025, n23026,
         n23027, n23028, n23029, n23030, n23031, n23032, n23033, n23034,
         n23035, n23036, n23037, n23038, n23039, n23040, n23041, n23042,
         n23043, n23044, n23045, n23046, n23047, n23048, n23049, n23050,
         n23051, n23052, n23053, n23054, n23055, n23056, n23057, n23058,
         n23059, n23060, n23061, n23062, n23063, n23064, n23065, n23066,
         n23067, n23068, n23069, n23070, n23071, n23072, n23073, n23074,
         n23075, n23076, n23077, n23078, n23079, n23080, n23081, n23082,
         n23083, n23084, n23085, n23086, n23087, n23088, n23089, n23090,
         n23091, n23092, n23093, n23094, n23095, n23096, n23097, n23098,
         n23099, n23100, n23101, n23102, n23103, n23104, n23105, n23106,
         n23107, n23108, n23109, n23110, n23111, n23112, n23113, n23114,
         n23115, n23116, n23117, n23118, n23119, n23120, n23121, n23122,
         n23123, n23124, n23125, n23126, n23127, n23128, n23129, n23130,
         n23131, n23132, n23133, n23134, n23135, n23136, n23137, n23138,
         n23139, n23140, n23141, n23142, n23143, n23144, n23145, n23146,
         n23147, n23148, n23149, n23150, n23151, n23152, n23153, n23154,
         n23155, n23156, n23157, n23158, n23159, n23160, n23161, n23162,
         n23163, n23164, n23165, n23166, n23167, n23168, n23169, n23170,
         n23171, n23172, n23173, n23174, n23175, n23176, n23177, n23178,
         n23179, n23180, n23181, n23182, n23183, n23184, n23185, n23186,
         n23187, n23188, n23189, n23190, n23191, n23192, n23193, n23194,
         n23195, n23196, n23197, n23198, n23199, n23200, n23201, n23202,
         n23203, n23204, n23205, n23206, n23207, n23208, n23209, n23210,
         n23211, n23212, n23213, n23214, n23215, n23216, n23217, n23218,
         n23219, n23220, n23221, n23222, n23223, n23224, n23225, n23226,
         n23227, n23228, n23229, n23230, n23231, n23232, n23233, n23234,
         n23235, n23236, n23237, n23238, n23239, n23240, n23241, n23242,
         n23243, n23244, n23245, n23246, n23247, n23248, n23249, n23250,
         n23251, n23252, n23253, n23254, n23255, n23256, n23257, n23258,
         n23259, n23260, n23261, n23262, n23263, n23264, n23265, n23266,
         n23267, n23268, n23269, n23270, n23271, n23272, n23273, n23274,
         n23275, n23276, n23277, n23278, n23279, n23280, n23281, n23282,
         n23283, n23284, n23285, n23286, n23287, n23288, n23289, n23290,
         n23291, n23292, n23293, n23294, n23295, n23296, n23297, n23298,
         n23299, n23300, n23301, n23302, n23303, n23304, n23305, n23306,
         n23307, n23308, n23309, n23310, n23311, n23312, n23313, n23314,
         n23315, n23316, n23317, n23318, n23319, n23320, n23321, n23322,
         n23323, n23324, n23325, n23326, n23327, n23328, n23329, n23330,
         n23331, n23332, n23333, n23334, n23335, n23336, n23337, n23338,
         n23339, n23340, n23341, n23342, n23343, n23344, n23345, n23346,
         n23347, n23348, n23349, n23350, n23351, n23352, n23353, n23354,
         n23355, n23356, n23357, n23358, n23359, n23360, n23361, n23362,
         n23363, n23364, n23365, n23366, n23367, n23368, n23369, n23370,
         n23371, n23372, n23373, n23374, n23375, n23376, n23377, n23378,
         n23379, n23380, n23381, n23382, n23383, n23384, n23385, n23386,
         n23387, n23388, n23389, n23390, n23391, n23392, n23393, n23394,
         n23395, n23396, n23397, n23398, n23399, n23400, n23401, n23402,
         n23403, n23404, n23405, n23406, n23407, n23408, n23409, n23410,
         n23411, n23412, n23413, n23414, n23415, n23416, n23417, n23418,
         n23419, n23420, n23421, n23422, n23423, n23424, n23425, n23426,
         n23427, n23428, n23429, n23430, n23431, n23432, n23433, n23434,
         n23435, n23436, n23437, n23438, n23439, n23440, n23441, n23442,
         n23443, n23444, n23445, n23446, n23447, n23448, n23449, n23450,
         n23451, n23452, n23453, n23454, n23455, n23456, n23457, n23458,
         n23459, n23460, n23461, n23462, n23463, n23464, n23465, n23466,
         n23467, n23468, n23469, n23470, n23471, n23472, n23473, n23474,
         n23475, n23476, n23477, n23478, n23479, n23480, n23481, n23482,
         n23483, n23484, n23485, n23486, n23487, n23488, n23489, n23490,
         n23491, n23492, n23493, n23494, n23495, n23496, n23497, n23498,
         n23499, n23500, n23501, n23502, n23503, n23504, n23505, n23506,
         n23507, n23508, n23509, n23510, n23511, n23512, n23513, n23514,
         n23515, n23516, n23517, n23518, n23519, n23520, n23521, n23522,
         n23523, n23524, n23525, n23526, n23527, n23528, n23529, n23530,
         n23531, n23532, n23533, n23534, n23535, n23536, n23537, n23538,
         n23539, n23540, n23541, n23542, n23543, n23544, n23545, n23546,
         n23547, n23548, n23549, n23550, n23551, n23552, n23553, n23554,
         n23555, n23556, n23557, n23558, n23559, n23560, n23561, n23562,
         n23563, n23564, n23565, n23566, n23567, n23568, n23569, n23570,
         n23571, n23572, n23573, n23574, n23575, n23576, n23577, n23578,
         n23579, n23580, n23581, n23582, n23583, n23584, n23585, n23586,
         n23587, n23588, n23589, n23590, n23591, n23592, n23593, n23594,
         n23595, n23596, n23597, n23598, n23599, n23600, n23601, n23602,
         n23603, n23604, n23605, n23606, n23607, n23608, n23609, n23610,
         n23611, n23612, n23613, n23614, n23615, n23616, n23617, n23618,
         n23619, n23620, n23621, n23622, n23623, n23624, n23625, n23626,
         n23627, n23628, n23629, n23630, n23631, n23632, n23633, n23634,
         n23635, n23636, n23637, n23638, n23639, n23640, n23641, n23642,
         n23643, n23644, n23645, n23646, n23647, n23648, n23649, n23650,
         n23651, n23652, n23653, n23654, n23655, n23656, n23657, n23658,
         n23659, n23660, n23661, n23662, n23663, n23664, n23665, n23666,
         n23667, n23668, n23669, n23670, n23671, n23672, n23673, n23674,
         n23675, n23676, n23677, n23678, n23679, n23680, n23681, n23682,
         n23683, n23684, n23685, n23686, n23687, n23688, n23689, n23690,
         n23691, n23692, n23693, n23694, n23695, n23696, n23697, n23698,
         n23699, n23700, n23701, n23702, n23703, n23704, n23705, n23706,
         n23707, n23708, n23709, n23710, n23711, n23712, n23713, n23714,
         n23715, n23716, n23717, n23718, n23719, n23720, n23721, n23722,
         n23723, n23724, n23725, n23726, n23727, n23728, n23729, n23730,
         n23731, n23732, n23733, n23734, n23735, n23736, n23737, n23738,
         n23739, n23740, n23741, n23742, n23743, n23744, n23745, n23746,
         n23747, n23748, n23749, n23750, n23751, n23752, n23753, n23754,
         n23755, n23756, n23757, n23758, n23759, n23760, n23761, n23762,
         n23763, n23764, n23765, n23766, n23767, n23768, n23769, n23770,
         n23771, n23772, n23773, n23774, n23775, n23776, n23777, n23778,
         n23779, n23780, n23781, n23782, n23783, n23784, n23785, n23786,
         n23787, n23788, n23789, n23790, n23791, n23792, n23793, n23794,
         n23795, n23796, n23797, n23798, n23799, n23800, n23801, n23802,
         n23803, n23804, n23805, n23806, n23807, n23808, n23809, n23810,
         n23811, n23812, n23813, n23814, n23815, n23816, n23817, n23818,
         n23819, n23820, n23821, n23822, n23823, n23824, n23825, n23826,
         n23827, n23828, n23829, n23830, n23831, n23832, n23833, n23834,
         n23835, n23836, n23837, n23838, n23839, n23840, n23841, n23842,
         n23843, n23844, n23845, n23846, n23847, n23848, n23849, n23850,
         n23851, n23852, n23853, n23854, n23855, n23856, n23857, n23858,
         n23859, n23860, n23861, n23862, n23863, n23864, n23865, n23866,
         n23867, n23868, n23869, n23870, n23871, n23872, n23873, n23874,
         n23875, n23876, n23877, n23878, n23879, n23880, n23881, n23882,
         n23883, n23884, n23885, n23886, n23887, n23888, n23889, n23890,
         n23891, n23892, n23893, n23894, n23895, n23896, n23897, n23898,
         n23899, n23900, n23901, n23902, n23903, n23904, n23905, n23906,
         n23907, n23908, n23909, n23910, n23911, n23912, n23913, n23914,
         n23915, n23916, n23917, n23918, n23919, n23920, n23921, n23922,
         n23923, n23924, n23925, n23926, n23927, n23928, n23929, n23930,
         n23931, n23932, n23933, n23934, n23935, n23936, n23937, n23938,
         n23939, n23940, n23941, n23942, n23943, n23944, n23945, n23946,
         n23947, n23948, n23949, n23950, n23951, n23952, n23953, n23954,
         n23955, n23956, n23957, n23958, n23959, n23960, n23961, n23962,
         n23963, n23964, n23965, n23966, n23967, n23968, n23969, n23970,
         n23971, n23972, n23973, n23974, n23975, n23976, n23977, n23978,
         n23979, n23980, n23981, n23982, n23983, n23984, n23985, n23986,
         n23987, n23988, n23989, n23990, n23991, n23992, n23993, n23994,
         n23995, n23996, n23997, n23998, n23999, n24000, n24001, n24002,
         n24003, n24004, n24005, n24006, n24007, n24008, n24009, n24010,
         n24011, n24012, n24013, n24014, n24015, n24016, n24017, n24018,
         n24019, n24020, n24021, n24022, n24023, n24024, n24025, n24026,
         n24027, n24028, n24029, n24030, n24031, n24032, n24033, n24034,
         n24035, n24036, n24037, n24038, n24039, n24040, n24041, n24042,
         n24043, n24044, n24045, n24046, n24047, n24048, n24049, n24050,
         n24051, n24052, n24053, n24054, n24055, n24056, n24057, n24058,
         n24059, n24060, n24061, n24062, n24063, n24064, n24065, n24066,
         n24067, n24068, n24069, n24070, n24071, n24072, n24073, n24074,
         n24075, n24076, n24077, n24078, n24079, n24080, n24081, n24082,
         n24083, n24084, n24085, n24086, n24087, n24088, n24089, n24090,
         n24091, n24092, n24093, n24094, n24095, n24096, n24097, n24098,
         n24099, n24100, n24101, n24102, n24103, n24104, n24105, n24106,
         n24107, n24108, n24109, n24110, n24111, n24112, n24113, n24114,
         n24115, n24116, n24117, n24118, n24119, n24120, n24121, n24122,
         n24123, n24124, n24125, n24126, n24127, n24128, n24129, n24130,
         n24131, n24132, n24133, n24134, n24135, n24136, n24137, n24138,
         n24139, n24140, n24141, n24142, n24143, n24144, n24145, n24146,
         n24147, n24148, n24149, n24150, n24151, n24152, n24153, n24154,
         n24155, n24156, n24157, n24158, n24159, n24160, n24161, n24162,
         n24163, n24164, n24165, n24166, n24167, n24168, n24169, n24170,
         n24171, n24172, n24173, n24174, n24175, n24176, n24177, n24178,
         n24179, n24180, n24181, n24182, n24183, n24184, n24185, n24186,
         n24187, n24188, n24189, n24190, n24191, n24192, n24193, n24194,
         n24195, n24196, n24197, n24198, n24199, n24200, n24201, n24202,
         n24203, n24204, n24205, n24206, n24207, n24208, n24209, n24210,
         n24211, n24212, n24213, n24214, n24215, n24216, n24217, n24218,
         n24219, n24220, n24221, n24222, n24223, n24224, n24225, n24226,
         n24227, n24228, n24229, n24230, n24231, n24232, n24233, n24234,
         n24235, n24236, n24237, n24238, n24239, n24240, n24241, n24242,
         n24243, n24244, n24245, n24246, n24247, n24248, n24249, n24250,
         n24251, n24252, n24253, n24254, n24255, n24256, n24257, n24258,
         n24259, n24260, n24261, n24262, n24263, n24264, n24265, n24266,
         n24267, n24268, n24269, n24270, n24271, n24272, n24273, n24274,
         n24275, n24276, n24277, n24278, n24279, n24280, n24281, n24282,
         n24283, n24284, n24285, n24286, n24287, n24288, n24289, n24290,
         n24291, n24292, n24293, n24294, n24295, n24296, n24297, n24298,
         n24299, n24300, n24301, n24302, n24303, n24304, n24305, n24306,
         n24307, n24308, n24309, n24310, n24311, n24312, n24313, n24314,
         n24315, n24316, n24317, n24318, n24319, n24320, n24321, n24322,
         n24323, n24324, n24325, n24326, n24327, n24328, n24329, n24330,
         n24331, n24332, n24333, n24334, n24335, n24336, n24337, n24338,
         n24339, n24340, n24341, n24342, n24343, n24344, n24345, n24346,
         n24347, n24348, n24349, n24350, n24351, n24352, n24353, n24354,
         n24355, n24356, n24357, n24358, n24359, n24360, n24361, n24362,
         n24363, n24364, n24365, n24366, n24367, n24368, n24369, n24370,
         n24371, n24372, n24373, n24374, n24375, n24376, n24377, n24378,
         n24379, n24380, n24381, n24382, n24383, n24384, n24385, n24386,
         n24387, n24388, n24389, n24390, n24391, n24392, n24393, n24394,
         n24395, n24396, n24397, n24398, n24399, n24400, n24401, n24402,
         n24403, n24404, n24405, n24406, n24407, n24408, n24409, n24410,
         n24411, n24412, n24413, n24414, n24415, n24416, n24417, n24418,
         n24419, n24420, n24421, n24422, n24423, n24424, n24425, n24426,
         n24427, n24428, n24429, n24430, n24431, n24432, n24433, n24434,
         n24435, n24436, n24437, n24438, n24439, n24440, n24441, n24442,
         n24443, n24444, n24445, n24446, n24447, n24448, n24449, n24450,
         n24451, n24452, n24453, n24454, n24455, n24456, n24457, n24458,
         n24459, n24460, n24461, n24462, n24463, n24464, n24465, n24466,
         n24467, n24468, n24469, n24470, n24471, n24472, n24473, n24474,
         n24475, n24476, n24477, n24478, n24479, n24480, n24481, n24482,
         n24483, n24484, n24485, n24486, n24487, n24488, n24489, n24490,
         n24491, n24492, n24493, n24494, n24495, n24496, n24497, n24498,
         n24499, n24500, n24501, n24502, n24503, n24504, n24505, n24506,
         n24507, n24508, n24509, n24510, n24511, n24512, n24513, n24514,
         n24515, n24516, n24517, n24518, n24519, n24520, n24521, n24522,
         n24523, n24524, n24525, n24526, n24527, n24528, n24529, n24530,
         n24531, n24532, n24533, n24534, n24535, n24536, n24537, n24538,
         n24539, n24540, n24541, n24542, n24543, n24544, n24545, n24546,
         n24547, n24548, n24549, n24550, n24551, n24552, n24553, n24554,
         n24555, n24556, n24557, n24558, n24559, n24560, n24561, n24562,
         n24563, n24564, n24565, n24566, n24567, n24568, n24569, n24570,
         n24571, n24572, n24573, n24574, n24575, n24576, n24577, n24578,
         n24579, n24580, n24581, n24582, n24583, n24584, n24585, n24586,
         n24587, n24588, n24589, n24590, n24591, n24592, n24593, n24594,
         n24595, n24596, n24597, n24598, n24599, n24600, n24601, n24602,
         n24603, n24604, n24605, n24606, n24607, n24608, n24609, n24610,
         n24611, n24612, n24613, n24614, n24615, n24616, n24617, n24618,
         n24619, n24620, n24621, n24622, n24623, n24624, n24625, n24626,
         n24627, n24628, n24629, n24630, n24631, n24632, n24633, n24634,
         n24635, n24636, n24637, n24638, n24639, n24640, n24641, n24642,
         n24643, n24644, n24645, n24646, n24647, n24648, n24649, n24650,
         n24651, n24652, n24653, n24654, n24655, n24656, n24657, n24658,
         n24659, n24660, n24661, n24662, n24663, n24664, n24665, n24666,
         n24667, n24668, n24669, n24670, n24671, n24672, n24673, n24674,
         n24675, n24676, n24677, n24678, n24679, n24680, n24681, n24682,
         n24683, n24684, n24685, n24686, n24687, n24688, n24689, n24690,
         n24691, n24692, n24693, n24694, n24695, n24696, n24697, n24698,
         n24699, n24700, n24701, n24702, n24703, n24704, n24705, n24706,
         n24707, n24708, n24709, n24710, n24711, n24712, n24713, n24714,
         n24715, n24716, n24717, n24718, n24719, n24720, n24721, n24722,
         n24723, n24724, n24725, n24726, n24727, n24728, n24729, n24730,
         n24731, n24732, n24733, n24734, n24735, n24736, n24737, n24738,
         n24739, n24740, n24741, n24742, n24743, n24744, n24745, n24746,
         n24747, n24748, n24749, n24750, n24751, n24752, n24753, n24754,
         n24755, n24756, n24757, n24758, n24759, n24760, n24761, n24762,
         n24763, n24764, n24765, n24766, n24767, n24768, n24769, n24770,
         n24771, n24772, n24773, n24774, n24775, n24776, n24777, n24778,
         n24779, n24780, n24781, n24782, n24783, n24784, n24785, n24786,
         n24787, n24788, n24789, n24790, n24791, n24792, n24793, n24794,
         n24795, n24796, n24797, n24798, n24799, n24800, n24801, n24802,
         n24803, n24804, n24805, n24806, n24807, n24808, n24809, n24810,
         n24811, n24812, n24813, n24814, n24815, n24816, n24817, n24818,
         n24819, n24820, n24821, n24822, n24823, n24824, n24825, n24826,
         n24827, n24828, n24829, n24830, n24831, n24832, n24833, n24834,
         n24835, n24836, n24837, n24838, n24839, n24840, n24841, n24842,
         n24843, n24844, n24845, n24846, n24847, n24848, n24849, n24850,
         n24851, n24852, n24853, n24854, n24855, n24856, n24857, n24858,
         n24859, n24860, n24861, n24862, n24863, n24864, n24865, n24866,
         n24867, n24868, n24869, n24870, n24871, n24872, n24873, n24874,
         n24875, n24876, n24877, n24878, n24879, n24880, n24881, n24882,
         n24883, n24884, n24885, n24886, n24887, n24888, n24889, n24890,
         n24891, n24892, n24893, n24894, n24895, n24896, n24897, n24898,
         n24899, n24900, n24901, n24902, n24903, n24904, n24905, n24906,
         n24907, n24908, n24909, n24910, n24911, n24912, n24913, n24914,
         n24915, n24916, n24917, n24918, n24919, n24920, n24921, n24922,
         n24923, n24924, n24925, n24926, n24927, n24928, n24929, n24930,
         n24931, n24932, n24933, n24934, n24935, n24936, n24937, n24938,
         n24939, n24940, n24941, n24942, n24943, n24944, n24945, n24946,
         n24947, n24948, n24949, n24950, n24951, n24952, n24953, n24954,
         n24955, n24956, n24957, n24958, n24959, n24960, n24961, n24962,
         n24963, n24964, n24965, n24966, n24967, n24968, n24969, n24970,
         n24971, n24972, n24973, n24974, n24975, n24976, n24977, n24978,
         n24979, n24980, n24981, n24982, n24983, n24984, n24985, n24986,
         n24987, n24988, n24989, n24990, n24991, n24992, n24993, n24994,
         n24995, n24996, n24997, n24998, n24999, n25000, n25001, n25002,
         n25003, n25004, n25005, n25006, n25007, n25008, n25009, n25010,
         n25011, n25012, n25013, n25014, n25015, n25016, n25017, n25018,
         n25019, n25020, n25021, n25022, n25023, n25024, n25025, n25026,
         n25027, n25028, n25029, n25030, n25031, n25032, n25033, n25034,
         n25035, n25036, n25037, n25038, n25039, n25040, n25041, n25042,
         n25043, n25044, n25045, n25046, n25047, n25048, n25049, n25050,
         n25051, n25052, n25053, n25054, n25055, n25056, n25057, n25058,
         n25059, n25060, n25061, n25062, n25063, n25064, n25065, n25066,
         n25067, n25068, n25069, n25070, n25071, n25072, n25073, n25074,
         n25075, n25076, n25077, n25078, n25079, n25080, n25081, n25082,
         n25083, n25084, n25085, n25086, n25087, n25088, n25089, n25090,
         n25091, n25092, n25093, n25094, n25095, n25096, n25097, n25098,
         n25099, n25100, n25101, n25102, n25103, n25104, n25105, n25106,
         n25107, n25108, n25109, n25110, n25111, n25112, n25113, n25114,
         n25115, n25116, n25117, n25118, n25119, n25120, n25121, n25122,
         n25123, n25124, n25125, n25126, n25127, n25128, n25129, n25130,
         n25131, n25132, n25133, n25134, n25135, n25136, n25137, n25138,
         n25139, n25140, n25141, n25142, n25143, n25144, n25145, n25146,
         n25147, n25148, n25149, n25150, n25151, n25152, n25153, n25154,
         n25155, n25156, n25157, n25158, n25159, n25160, n25161, n25162,
         n25163, n25164, n25165, n25166, n25167, n25168, n25169, n25170,
         n25171, n25172, n25173, n25174, n25175, n25176, n25177, n25178,
         n25179, n25180, n25181, n25182, n25183, n25184, n25185, n25186,
         n25187, n25188, n25189, n25190, n25191, n25192, n25193, n25194,
         n25195, n25196, n25197, n25198, n25199, n25200, n25201, n25202,
         n25203, n25204, n25205, n25206, n25207, n25208, n25209, n25210,
         n25211, n25212, n25213, n25214, n25215, n25216, n25217, n25218,
         n25219, n25220, n25221, n25222, n25223, n25224, n25225, n25226,
         n25227, n25228, n25229, n25230, n25231, n25232, n25233, n25234,
         n25235, n25236, n25237, n25238, n25239, n25240, n25241, n25242,
         n25243, n25244, n25245, n25246, n25247, n25248, n25249, n25250,
         n25251, n25252, n25253, n25254, n25255, n25256, n25257, n25258,
         n25259, n25260, n25261, n25262, n25263, n25264, n25265, n25266,
         n25267, n25268, n25269, n25270, n25271, n25272, n25273, n25274,
         n25275, n25276, n25277, n25278, n25279, n25280, n25281, n25282,
         n25283, n25284, n25285, n25286, n25287, n25288, n25289, n25290,
         n25291, n25292, n25293, n25294, n25295, n25296, n25297, n25298,
         n25299, n25300, n25301, n25302, n25303, n25304, n25305, n25306,
         n25307, n25308, n25309, n25310, n25311, n25312, n25313, n25314,
         n25315, n25316, n25317, n25318, n25319, n25320, n25321, n25322,
         n25323, n25324, n25325, n25326, n25327, n25328, n25329, n25330,
         n25331, n25332, n25333, n25334, n25335, n25336, n25337, n25338,
         n25339, n25340, n25341, n25342, n25343, n25344, n25345, n25346,
         n25347, n25348, n25349, n25350, n25351, n25352, n25353, n25354,
         n25355, n25356, n25357, n25358, n25359, n25360, n25361, n25362,
         n25363, n25364, n25365, n25366, n25367, n25368, n25369, n25370,
         n25371, n25372, n25373, n25374, n25375, n25376, n25377, n25378,
         n25379, n25380, n25381, n25382, n25383, n25384, n25385, n25386,
         n25387, n25388, n25389, n25390, n25391, n25392, n25393, n25394,
         n25395, n25396, n25397, n25398, n25399, n25400, n25401, n25402,
         n25403, n25404, n25405, n25406, n25407, n25408, n25409, n25410,
         n25411, n25412, n25413, n25414, n25415, n25416, n25417, n25418,
         n25419, n25420, n25421, n25422, n25423, n25424, n25425, n25426,
         n25427, n25428, n25429, n25430, n25431, n25432, n25433, n25434,
         n25435, n25436, n25437, n25438, n25439, n25440, n25441, n25442,
         n25443, n25444, n25445, n25446, n25447, n25448, n25449, n25450,
         n25451, n25452, n25453, n25454, n25455, n25456, n25457, n25458,
         n25459, n25460, n25461, n25462, n25463, n25464, n25465, n25466,
         n25467, n25468, n25469, n25470, n25471, n25472, n25473, n25474,
         n25475, n25476, n25477, n25478, n25479, n25480, n25481, n25482,
         n25483, n25484, n25485, n25486, n25487, n25488, n25489, n25490,
         n25491, n25492, n25493, n25494, n25495, n25496, n25497, n25498,
         n25499, n25500, n25501, n25502, n25503, n25504, n25505, n25506,
         n25507, n25508, n25509, n25510, n25511, n25512, n25513, n25514,
         n25515, n25516, n25517, n25518, n25519, n25520, n25521, n25522,
         n25523, n25524, n25525, n25526, n25527, n25528, n25529, n25530,
         n25531, n25532, n25533, n25534, n25535, n25536, n25537, n25538,
         n25539, n25540, n25541, n25542, n25543, n25544, n25545, n25546,
         n25547, n25548, n25549, n25550, n25551, n25552, n25553, n25554,
         n25555, n25556, n25557, n25558, n25559, n25560, n25561, n25562,
         n25563, n25564, n25565, n25566, n25567, n25568, n25569, n25570,
         n25571, n25572, n25573, n25574, n25575, n25576, n25577, n25578,
         n25579, n25580, n25581, n25582, n25583, n25584, n25585, n25586,
         n25587, n25588, n25589, n25590, n25591, n25592, n25593, n25594,
         n25595, n25596, n25597, n25598, n25599, n25600, n25601, n25602,
         n25603, n25604, n25605, n25606, n25607, n25608, n25609, n25610,
         n25611, n25612, n25613, n25614, n25615, n25616, n25617, n25618,
         n25619, n25620, n25621, n25622, n25623, n25624, n25625, n25626,
         n25627, n25628, n25629, n25630, n25631, n25632, n25633, n25634,
         n25635, n25636, n25637, n25638, n25639, n25640, n25641, n25642,
         n25643, n25644, n25645, n25646, n25647, n25648, n25649, n25650,
         n25651, n25652, n25653, n25654, n25655, n25656, n25657, n25658,
         n25659, n25660, n25661, n25662, n25663, n25664, n25665, n25666,
         n25667, n25668, n25669, n25670, n25671, n25672, n25673, n25674,
         n25675, n25676, n25677, n25678, n25679, n25680, n25681, n25682,
         n25683, n25684, n25685, n25686, n25687, n25688, n25689, n25690,
         n25691, n25692, n25693, n25694, n25695, n25696, n25697, n25698,
         n25699, n25700, n25701, n25702, n25703, n25704, n25705, n25706,
         n25707, n25708, n25709, n25710, n25711, n25712, n25713, n25714,
         n25715, n25716, n25717, n25718, n25719, n25720, n25721, n25722,
         n25723, n25724, n25725, n25726, n25727, n25728, n25729, n25730,
         n25731, n25732, n25733, n25734, n25735, n25736, n25737, n25738,
         n25739, n25740, n25741, n25742, n25743, n25744, n25745, n25746,
         n25747, n25748, n25749, n25750, n25751, n25752, n25753, n25754,
         n25755, n25756, n25757, n25758, n25759, n25760, n25761, n25762,
         n25763, n25764, n25765, n25766, n25767, n25768, n25769, n25770,
         n25771, n25772, n25773, n25774, n25775, n25776, n25777, n25778,
         n25779, n25780, n25781, n25782, n25783, n25784, n25785, n25786,
         n25787, n25788, n25789, n25790, n25791, n25792, n25793, n25794,
         n25795, n25796, n25797, n25798, n25799, n25800, n25801, n25802,
         n25803, n25804, n25805, n25806, n25807, n25808, n25809, n25810,
         n25811, n25812, n25813, n25814, n25815, n25816, n25817, n25818,
         n25819, n25820, n25821, n25822, n25823, n25824, n25825, n25826,
         n25827, n25828, n25829, n25830, n25831, n25832, n25833, n25834,
         n25835, n25836, n25837, n25838, n25839, n25840, n25841, n25842,
         n25843, n25844, n25845, n25846, n25847, n25848, n25849, n25850,
         n25851, n25852, n25853, n25854, n25855, n25856, n25857, n25858,
         n25859, n25860, n25861, n25862, n25863, n25864, n25865, n25866,
         n25867, n25868, n25869, n25870, n25871, n25872, n25873, n25874,
         n25875, n25876, n25877, n25878, n25879, n25880, n25881, n25882,
         n25883, n25884, n25885, n25886, n25887, n25888, n25889, n25890,
         n25891, n25892, n25893, n25894, n25895, n25896, n25897, n25898,
         n25899, n25900, n25901, n25902, n25903, n25904, n25905, n25906,
         n25907, n25908, n25909, n25910, n25911, n25912, n25913, n25914,
         n25915, n25916, n25917, n25918, n25919, n25920, n25921, n25922,
         n25923, n25924, n25925, n25926, n25927, n25928, n25929, n25930,
         n25931, n25932, n25933, n25934, n25935, n25936, n25937, n25938,
         n25939, n25940, n25941, n25942, n25943, n25944, n25945, n25946,
         n25947, n25948, n25949, n25950, n25951, n25952, n25953, n25954,
         n25955, n25956, n25957, n25958, n25959, n25960, n25961, n25962,
         n25963, n25964, n25965, n25966, n25967, n25968, n25969, n25970,
         n25971, n25972, n25973, n25974, n25975, n25976, n25977, n25978,
         n25979, n25980, n25981, n25982, n25983, n25984, n25985, n25986,
         n25987, n25988, n25989, n25990, n25991, n25992, n25993, n25994,
         n25995, n25996, n25997, n25998, n25999, n26000, n26001, n26002,
         n26003, n26004, n26005, n26006, n26007, n26008, n26009, n26010,
         n26011, n26012, n26013, n26014, n26015, n26016, n26017, n26018,
         n26019, n26020, n26021, n26022, n26023, n26024, n26025, n26026,
         n26027, n26028, n26029, n26030, n26031, n26032, n26033, n26034,
         n26035, n26036, n26037, n26038, n26039, n26040, n26041, n26042,
         n26043, n26044, n26045, n26046, n26047, n26048, n26049, n26050,
         n26051, n26052, n26053, n26054, n26055, n26056, n26057, n26058,
         n26059, n26060, n26061, n26062, n26063, n26064, n26065, n26066,
         n26067, n26068, n26069, n26070, n26071, n26072, n26073, n26074,
         n26075, n26076, n26077, n26078, n26079, n26080, n26081, n26082,
         n26083, n26084, n26085, n26086, n26087, n26088, n26089, n26090,
         n26091, n26092, n26093, n26094, n26095, n26096, n26097, n26098,
         n26099, n26100, n26101, n26102, n26103, n26104, n26105, n26106,
         n26107, n26108, n26109, n26110, n26111, n26112, n26113, n26114,
         n26115, n26116, n26117, n26118, n26119, n26120, n26121, n26122,
         n26123, n26124, n26125, n26126, n26127, n26128, n26129, n26130,
         n26131, n26132, n26133, n26134, n26135, n26136, n26137, n26138,
         n26139, n26140, n26141, n26142, n26143, n26144, n26145, n26146,
         n26147, n26148, n26149, n26150, n26151, n26152, n26153, n26154,
         n26155, n26156, n26157, n26158, n26159, n26160, n26161, n26162,
         n26163, n26164, n26165, n26166, n26167, n26168, n26169, n26170,
         n26171, n26172, n26173, n26174, n26175, n26176, n26177, n26178,
         n26179, n26180, n26181, n26182, n26183, n26184, n26185, n26186,
         n26187, n26188, n26189, n26190, n26191, n26192, n26193, n26194,
         n26195, n26196, n26197, n26198, n26199, n26200, n26201, n26202,
         n26203, n26204, n26205, n26206, n26207, n26208, n26209, n26210,
         n26211, n26212, n26213, n26214, n26215, n26216, n26217, n26218,
         n26219, n26220, n26221, n26222, n26223, n26224, n26225, n26226,
         n26227, n26228, n26229, n26230, n26231, n26232, n26233, n26234,
         n26235, n26236, n26237, n26238, n26239, n26240, n26241, n26242,
         n26243, n26244, n26245, n26246, n26247, n26248, n26249, n26250,
         n26251, n26252, n26253, n26254, n26255, n26256, n26257, n26258,
         n26259, n26260, n26261, n26262, n26263, n26264, n26265, n26266,
         n26267, n26268, n26269, n26270, n26271, n26272, n26273, n26274,
         n26275, n26276, n26277, n26278, n26279, n26280, n26281, n26282,
         n26283, n26284, n26285, n26286, n26287, n26288, n26289, n26290,
         n26291, n26292, n26293, n26294, n26295, n26296, n26297, n26298,
         n26299, n26300, n26301, n26302, n26303, n26304, n26305, n26306,
         n26307, n26308, n26309, n26310, n26311, n26312, n26313, n26314,
         n26315, n26316, n26317, n26318, n26319, n26320, n26321, n26322,
         n26323, n26324, n26325, n26326, n26327, n26328, n26329, n26330,
         n26331, n26332, n26333, n26334, n26335, n26336, n26337, n26338,
         n26339, n26340, n26341, n26342, n26343, n26344, n26345, n26346,
         n26347, n26348, n26349, n26350, n26351, n26352, n26353, n26354,
         n26355, n26356, n26357, n26358, n26359, n26360, n26361, n26362,
         n26363, n26364, n26365, n26366, n26367, n26368, n26369, n26370,
         n26371, n26372, n26373, n26374, n26375, n26376, n26377, n26378,
         n26379, n26380, n26381, n26382, n26383, n26384, n26385, n26386,
         n26387, n26388, n26389, n26390, n26391, n26392, n26393, n26394,
         n26395, n26396, n26397, n26398, n26399, n26400, n26401, n26402,
         n26403, n26404, n26405, n26406, n26407, n26408, n26409, n26410,
         n26411, n26412, n26413, n26414, n26415, n26416, n26417, n26418,
         n26419, n26420, n26421, n26422, n26423, n26424, n26425, n26426,
         n26427, n26428, n26429, n26430, n26431, n26432, n26433, n26434,
         n26435, n26436, n26437, n26438, n26439, n26440, n26441, n26442,
         n26443, n26444, n26445, n26446, n26447, n26448, n26449, n26450,
         n26451, n26452, n26453, n26454, n26455, n26456, n26457, n26458,
         n26459, n26460, n26461, n26462, n26463, n26464, n26465, n26466,
         n26467, n26468, n26469, n26470, n26471, n26472, n26473, n26474,
         n26475, n26476, n26477, n26478, n26479, n26480, n26481, n26482,
         n26483, n26484, n26485, n26486, n26487, n26488, n26489, n26490,
         n26491, n26492, n26493, n26494, n26495, n26496, n26497, n26498,
         n26499, n26500, n26501, n26502, n26503, n26504, n26505, n26506,
         n26507, n26508, n26509, n26510, n26511, n26512, n26513, n26514,
         n26515, n26516, n26517, n26518, n26519, n26520, n26521, n26522,
         n26523, n26524, n26525, n26526, n26527, n26528, n26529, n26530,
         n26531, n26532, n26533, n26534, n26535, n26536, n26537, n26538,
         n26539, n26540, n26541, n26542, n26543, n26544, n26545, n26546,
         n26547, n26548, n26549, n26550, n26551, n26552, n26553, n26554,
         n26555, n26556, n26557, n26558, n26559, n26560, n26561, n26562,
         n26563, n26564, n26565, n26566, n26567, n26568, n26569, n26570,
         n26571, n26572, n26573, n26574, n26575, n26576, n26577, n26578,
         n26579, n26580, n26581, n26582, n26583, n26584, n26585, n26586,
         n26587, n26588, n26589, n26590, n26591, n26592, n26593, n26594,
         n26595, n26596, n26597, n26598, n26599, n26600, n26601, n26602,
         n26603, n26604, n26605, n26606, n26607, n26608, n26609, n26610,
         n26611, n26612, n26613, n26614, n26615, n26616, n26617, n26618,
         n26619, n26620, n26621, n26622, n26623, n26624, n26625, n26626,
         n26627, n26628, n26629, n26630, n26631, n26632, n26633, n26634,
         n26635, n26636, n26637, n26638, n26639, n26640, n26641, n26642,
         n26643, n26644, n26645, n26646, n26647, n26648, n26649, n26650,
         n26651, n26652, n26653, n26654, n26655, n26656, n26657, n26658,
         n26659, n26660, n26661, n26662, n26663, n26664, n26665, n26666,
         n26667, n26668, n26669, n26670, n26671, n26672, n26673, n26674,
         n26675, n26676, n26677, n26678, n26679, n26680, n26681, n26682,
         n26683, n26684, n26685, n26686, n26687, n26688, n26689, n26690,
         n26691, n26692, n26693, n26694, n26695, n26696, n26697, n26698,
         n26699, n26700, n26701, n26702, n26703, n26704, n26705, n26706,
         n26707, n26708, n26709, n26710, n26711, n26712, n26713, n26714,
         n26715, n26716, n26717, n26718, n26719, n26720, n26721, n26722,
         n26723, n26724, n26725, n26726, n26727, n26728, n26729, n26730,
         n26731, n26732, n26733, n26734, n26735, n26736, n26737, n26738,
         n26739, n26740, n26741, n26742, n26743, n26744, n26745, n26746,
         n26747, n26748, n26749, n26750, n26751, n26752, n26753, n26754,
         n26755, n26756, n26757, n26758, n26759, n26760, n26761, n26762,
         n26763, n26764, n26765, n26766, n26767, n26768, n26769, n26770,
         n26771, n26772, n26773, n26774, n26775, n26776, n26777, n26778,
         n26779, n26780, n26781, n26782, n26783, n26784, n26785, n26786,
         n26787, n26788, n26789, n26790, n26791, n26792, n26793, n26794,
         n26795, n26796, n26797, n26798, n26799, n26800, n26801, n26802,
         n26803, n26804, n26805, n26806, n26807, n26808, n26809, n26810,
         n26811, n26812, n26813, n26814, n26815, n26816, n26817, n26818,
         n26819, n26820, n26821, n26822, n26823, n26824, n26825, n26826,
         n26827, n26828, n26829, n26830, n26831, n26832, n26833, n26834,
         n26835, n26836, n26837, n26838, n26839, n26840, n26841, n26842,
         n26843, n26844, n26845, n26846, n26847, n26848, n26849, n26850,
         n26851, n26852, n26853, n26854, n26855, n26856, n26857, n26858,
         n26859, n26860, n26861, n26862, n26863, n26864, n26865, n26866,
         n26867, n26868, n26869, n26870, n26871, n26872, n26873, n26874,
         n26875, n26876, n26877, n26878, n26879, n26880, n26881, n26882,
         n26883, n26884, n26885, n26886, n26887, n26888, n26889, n26890,
         n26891, n26892, n26893, n26894, n26895, n26896, n26897, n26898,
         n26899, n26900, n26901, n26902, n26903, n26904, n26905, n26906,
         n26907, n26908, n26909, n26910, n26911, n26912, n26913, n26914,
         n26915, n26916, n26917, n26918, n26919, n26920, n26921, n26922,
         n26923, n26924, n26925, n26926, n26927, n26928, n26929, n26930,
         n26931, n26932, n26933, n26934, n26935, n26936, n26937, n26938,
         n26939, n26940, n26941, n26942, n26943, n26944, n26945, n26946,
         n26947, n26948, n26949, n26950, n26951, n26952, n26953, n26954,
         n26955, n26956, n26957, n26958, n26959, n26960, n26961, n26962,
         n26963, n26964, n26965, n26966, n26967, n26968, n26969, n26970,
         n26971, n26972, n26973, n26974, n26975, n26976, n26977, n26978,
         n26979, n26980, n26981, n26982, n26983, n26984, n26985, n26986,
         n26987, n26988, n26989, n26990, n26991, n26992, n26993, n26994,
         n26995, n26996, n26997, n26998, n26999, n27000, n27001, n27002,
         n27003, n27004, n27005, n27006, n27007, n27008, n27009, n27010,
         n27011, n27012, n27013, n27014, n27015, n27016, n27017, n27018,
         n27019, n27020, n27021, n27022, n27023, n27024, n27025, n27026,
         n27027, n27028, n27029, n27030, n27031, n27032, n27033, n27034,
         n27035, n27036, n27037, n27038, n27039, n27040, n27041, n27042,
         n27043, n27044, n27045, n27046, n27047, n27048, n27049, n27050,
         n27051, n27052, n27053, n27054, n27055, n27056, n27057, n27058,
         n27059, n27060, n27061, n27062, n27063, n27064, n27065, n27066,
         n27067, n27068, n27069, n27070, n27071, n27072, n27073, n27074,
         n27075, n27076, n27077, n27078, n27079, n27080, n27081, n27082,
         n27083, n27084, n27085, n27086, n27087, n27088, n27089, n27090,
         n27091, n27092, n27093, n27094, n27095, n27096, n27097, n27098,
         n27099, n27100, n27101, n27102, n27103, n27104, n27105, n27106,
         n27107, n27108, n27109, n27110, n27111, n27112, n27113, n27114,
         n27115, n27116, n27117, n27118, n27119, n27120, n27121, n27122,
         n27123, n27124, n27125, n27126, n27127, n27128, n27129, n27130,
         n27131, n27132, n27133, n27134, n27135, n27136, n27137, n27138,
         n27139, n27140, n27141, n27142, n27143, n27144, n27145, n27146,
         n27147, n27148, n27149, n27150, n27151, n27152, n27153, n27154,
         n27155, n27156, n27157, n27158, n27159, n27160, n27161, n27162,
         n27163, n27164, n27165, n27166, n27167, n27168, n27169, n27170,
         n27171, n27172, n27173, n27174, n27175, n27176, n27177, n27178,
         n27179, n27180, n27181, n27182, n27183, n27184, n27185, n27186,
         n27187, n27188, n27189, n27190, n27191, n27192, n27193, n27194,
         n27195, n27196, n27197, n27198, n27199, n27200, n27201, n27202,
         n27203, n27204, n27205, n27206, n27207, n27208, n27209, n27210,
         n27211, n27212, n27213, n27214, n27215, n27216, n27217, n27218,
         n27219, n27220, n27221, n27222, n27223, n27224, n27225, n27226,
         n27227, n27228, n27229, n27230, n27231, n27232, n27233, n27234,
         n27235, n27236, n27237, n27238, n27239, n27240, n27241, n27242,
         n27243, n27244, n27245, n27246, n27247, n27248, n27249, n27250,
         n27251, n27252, n27253, n27254, n27255, n27256, n27257, n27258,
         n27259, n27260, n27261, n27262, n27263, n27264, n27265, n27266,
         n27267, n27268, n27269, n27270, n27271, n27272, n27273, n27274,
         n27275, n27276, n27277, n27278, n27279, n27280, n27281, n27282,
         n27283, n27284, n27285, n27286, n27287, n27288, n27289, n27290,
         n27291, n27292, n27293, n27294, n27295, n27296, n27297, n27298,
         n27299, n27300, n27301, n27302, n27303, n27304, n27305, n27306,
         n27307, n27308, n27309, n27310, n27311, n27312, n27313, n27314,
         n27315, n27316, n27317, n27318, n27319, n27320, n27321, n27322,
         n27323, n27324, n27325, n27326, n27327, n27328, n27329, n27330,
         n27331, n27332, n27333, n27334, n27335, n27336, n27337, n27338,
         n27339, n27340, n27341, n27342, n27343, n27344, n27345, n27346,
         n27347, n27348, n27349, n27350, n27351, n27352, n27353, n27354,
         n27355, n27356, n27357, n27358, n27359, n27360, n27361, n27362,
         n27363, n27364, n27365, n27366, n27367, n27368, n27369, n27370,
         n27371, n27372, n27373, n27374, n27375, n27376, n27377, n27378,
         n27379, n27380, n27381, n27382, n27383, n27384, n27385, n27386,
         n27387, n27388, n27389, n27390, n27391, n27392, n27393, n27394,
         n27395, n27396, n27397, n27398, n27399, n27400, n27401, n27402,
         n27403, n27404, n27405, n27406, n27407, n27408, n27409, n27410,
         n27411, n27412, n27413, n27414, n27415, n27416, n27417, n27418,
         n27419, n27420, n27421, n27422, n27423, n27424, n27425, n27426,
         n27427, n27428, n27429, n27430, n27431, n27432, n27433, n27434,
         n27435, n27436, n27437, n27438, n27439, n27440, n27441, n27442,
         n27443, n27444, n27445, n27446, n27447, n27448, n27449, n27450,
         n27451, n27452, n27453, n27454, n27455, n27456, n27457, n27458,
         n27459, n27460, n27461, n27462, n27463, n27464, n27465, n27466,
         n27467, n27468, n27469, n27470, n27471, n27472, n27473, n27474,
         n27475, n27476, n27477, n27478, n27479, n27480, n27481, n27482,
         n27483, n27484, n27485, n27486, n27487, n27488, n27489, n27490,
         n27491, n27492, n27493, n27494, n27495, n27496, n27497, n27498,
         n27499, n27500, n27501, n27502, n27503, n27504, n27505, n27506,
         n27507, n27508, n27509, n27510, n27511, n27512, n27513, n27514,
         n27515, n27516, n27517, n27518, n27519, n27520, n27521, n27522,
         n27523, n27524, n27525, n27526, n27527, n27528, n27529, n27530,
         n27531, n27532, n27533, n27534, n27535, n27536, n27537, n27538,
         n27539, n27540, n27541, n27542, n27543, n27544, n27545, n27546,
         n27547, n27548, n27549, n27550, n27551, n27552, n27553, n27554,
         n27555, n27556, n27557, n27558, n27559, n27560, n27561, n27562,
         n27563, n27564, n27565, n27566, n27567, n27568, n27569, n27570,
         n27571, n27572, n27573, n27574, n27575, n27576, n27577, n27578,
         n27579, n27580, n27581, n27582, n27583, n27584, n27585, n27586,
         n27587, n27588, n27589, n27590, n27591, n27592, n27593, n27594,
         n27595, n27596, n27597, n27598, n27599, n27600, n27601, n27602,
         n27603, n27604, n27605, n27606, n27607, n27608, n27609, n27610,
         n27611, n27612, n27613, n27614, n27615, n27616, n27617, n27618,
         n27619, n27620, n27621, n27622, n27623, n27624, n27625, n27626,
         n27627, n27628, n27629, n27630, n27631, n27632, n27633, n27634,
         n27635, n27636, n27637, n27638, n27639, n27640, n27641, n27642,
         n27643, n27644, n27645, n27646, n27647, n27648, n27649, n27650,
         n27651, n27652, n27653, n27654, n27655, n27656, n27657, n27658,
         n27659, n27660, n27661, n27662, n27663, n27664, n27665, n27666,
         n27667, n27668, n27669, n27670, n27671, n27672, n27673, n27674,
         n27675, n27676, n27677, n27678, n27679, n27680, n27681, n27682,
         n27683, n27684, n27685, n27686, n27687, n27688, n27689, n27690,
         n27691, n27692, n27693, n27694, n27695, n27696, n27697, n27698,
         n27699, n27700, n27701, n27702, n27703, n27704, n27705, n27706,
         n27707, n27708, n27709, n27710, n27711, n27712, n27713, n27714,
         n27715, n27716, n27717, n27718, n27719, n27720, n27721, n27722,
         n27723, n27724, n27725, n27726, n27727, n27728, n27729, n27730,
         n27731, n27732, n27733, n27734, n27735, n27736, n27737, n27738,
         n27739, n27740, n27741, n27742, n27743, n27744, n27745, n27746,
         n27747, n27748, n27749, n27750, n27751, n27752, n27753, n27754,
         n27755, n27756, n27757, n27758, n27759, n27760, n27761, n27762,
         n27763, n27764, n27765, n27766, n27767, n27768, n27769, n27770,
         n27771, n27772, n27773, n27774, n27775, n27776, n27777, n27778,
         n27779, n27780, n27781, n27782, n27783, n27784, n27785, n27786,
         n27787, n27788, n27789, n27790, n27791, n27792, n27793, n27794,
         n27795, n27796, n27797, n27798, n27799, n27800, n27801, n27802,
         n27803, n27804, n27805, n27806, n27807, n27808, n27809, n27810,
         n27811, n27812, n27813, n27814, n27815, n27816, n27817, n27818,
         n27819, n27820, n27821, n27822, n27823, n27824, n27825, n27826,
         n27827, n27828, n27829, n27830, n27831, n27832, n27833, n27834,
         n27835, n27836, n27837, n27838, n27839, n27840, n27841, n27842,
         n27843, n27844, n27845, n27846, n27847, n27848, n27849, n27850,
         n27851, n27852, n27853, n27854, n27855, n27856, n27857, n27858,
         n27859, n27860, n27861, n27862, n27863, n27864, n27865, n27866,
         n27867, n27868, n27869, n27870, n27871, n27872, n27873, n27874,
         n27875, n27876, n27877, n27878, n27879, n27880, n27881, n27882,
         n27883, n27884, n27885, n27886, n27887, n27888, n27889, n27890,
         n27891, n27892, n27893, n27894, n27895, n27896, n27897, n27898,
         n27899, n27900, n27901, n27902, n27903, n27904, n27905, n27906,
         n27907, n27908, n27909, n27910, n27911, n27912, n27913, n27914,
         n27915, n27916, n27917, n27918, n27919, n27920, n27921, n27922,
         n27923, n27924, n27925, n27926, n27927, n27928, n27929, n27930,
         n27931, n27932, n27933, n27934, n27935, n27936, n27937, n27938,
         n27939, n27940, n27941, n27942, n27943, n27944, n27945, n27946,
         n27947, n27948, n27949, n27950, n27951, n27952, n27953, n27954,
         n27955, n27956, n27957, n27958, n27959, n27960, n27961, n27962,
         n27963, n27964, n27965, n27966, n27967, n27968, n27969, n27970,
         n27971, n27972, n27973, n27974, n27975, n27976, n27977, n27978,
         n27979, n27980, n27981, n27982, n27983, n27984, n27985, n27986,
         n27987, n27988, n27989, n27990, n27991, n27992, n27993, n27994,
         n27995, n27996, n27997, n27998, n27999, n28000, n28001, n28002,
         n28003, n28004, n28005, n28006, n28007, n28008, n28009, n28010,
         n28011, n28012, n28013, n28014, n28015, n28016, n28017, n28018,
         n28019, n28020, n28021, n28022, n28023, n28024, n28025, n28026,
         n28027, n28028, n28029, n28030, n28031, n28032, n28033, n28034,
         n28035, n28036, n28037, n28038, n28039, n28040, n28041, n28042,
         n28043, n28044, n28045, n28046, n28047, n28048, n28049, n28050,
         n28051, n28052, n28053, n28054, n28055, n28056, n28057, n28058,
         n28059, n28060, n28061, n28062, n28063, n28064, n28065, n28066,
         n28067, n28068, n28069, n28070, n28071, n28072, n28073, n28074,
         n28075, n28076, n28077, n28078, n28079, n28080, n28081, n28082,
         n28083, n28084, n28085, n28086, n28087, n28088, n28089, n28090,
         n28091, n28092, n28093, n28094, n28095, n28096, n28097, n28098,
         n28099, n28100, n28101, n28102, n28103, n28104, n28105, n28106,
         n28107, n28108, n28109, n28110, n28111, n28112, n28113, n28114,
         n28115, n28116, n28117, n28118, n28119, n28120, n28121, n28122,
         n28123, n28124, n28125, n28126, n28127, n28128, n28129, n28130,
         n28131, n28132, n28133, n28134, n28135, n28136, n28137, n28138,
         n28139, n28140, n28141, n28142, n28143, n28144, n28145, n28146,
         n28147, n28148, n28149, n28150, n28151, n28152, n28153, n28154,
         n28155, n28156, n28157, n28158, n28159, n28160, n28161, n28162,
         n28163, n28164, n28165, n28166, n28167, n28168, n28169, n28170,
         n28171, n28172, n28173, n28174, n28175, n28176, n28177, n28178,
         n28179, n28180, n28181, n28182, n28183, n28184, n28185, n28186,
         n28187, n28188, n28189, n28190, n28191, n28192, n28193, n28194,
         n28195, n28196, n28197, n28198, n28199, n28200, n28201, n28202,
         n28203, n28204, n28205, n28206, n28207, n28208, n28209, n28210,
         n28211, n28212, n28213, n28214, n28215, n28216, n28217, n28218,
         n28219, n28220, n28221, n28222, n28223, n28224, n28225, n28226,
         n28227, n28228, n28229, n28230, n28231, n28232, n28233, n28234,
         n28235, n28236, n28237, n28238, n28239, n28240, n28241, n28242,
         n28243, n28244, n28245, n28246, n28247, n28248, n28249, n28250,
         n28251, n28252, n28253, n28254, n28255, n28256, n28257, n28258,
         n28259, n28260, n28261, n28262, n28263, n28264, n28265, n28266,
         n28267, n28268, n28269, n28270, n28271, n28272, n28273, n28274,
         n28275, n28276, n28277, n28278, n28279, n28280, n28281, n28282,
         n28283, n28284, n28285, n28286, n28287, n28288, n28289, n28290,
         n28291, n28292, n28293, n28294, n28295, n28296, n28297, n28298,
         n28299, n28300, n28301, n28302, n28303, n28304, n28305, n28306,
         n28307, n28308, n28309, n28310, n28311, n28312, n28313, n28314,
         n28315, n28316, n28317, n28318, n28319, n28320, n28321, n28322,
         n28323, n28324, n28325, n28326, n28327, n28328, n28329, n28330,
         n28331, n28332, n28333, n28334, n28335, n28336, n28337, n28338,
         n28339, n28340, n28341, n28342, n28343, n28344, n28345, n28346,
         n28347, n28348, n28349, n28350, n28351, n28352, n28353, n28354,
         n28355, n28356, n28357, n28358, n28359, n28360, n28361, n28362,
         n28363, n28364, n28365, n28366, n28367, n28368, n28369, n28370,
         n28371, n28372, n28373, n28374, n28375, n28376, n28377, n28378,
         n28379, n28380, n28381, n28382, n28383, n28384, n28385, n28386,
         n28387, n28388, n28389, n28390, n28391, n28392, n28393, n28394,
         n28395, n28396, n28397, n28398, n28399, n28400, n28401, n28402,
         n28403, n28404, n28405, n28406, n28407, n28408, n28409, n28410,
         n28411, n28412, n28413, n28414, n28415, n28416, n28417, n28418,
         n28419, n28420, n28421, n28422, n28423, n28424, n28425, n28426,
         n28427, n28428, n28429, n28430, n28431, n28432, n28433, n28434,
         n28435, n28436, n28437, n28438, n28439, n28440, n28441, n28442,
         n28443, n28444, n28445, n28446, n28447, n28448, n28449, n28450,
         n28451, n28452, n28453, n28454, n28455, n28456, n28457, n28458,
         n28459, n28460, n28461, n28462, n28463, n28464, n28465, n28466,
         n28467, n28468, n28469, n28470, n28471, n28472, n28473, n28474,
         n28475, n28476, n28477, n28478, n28479, n28480, n28481, n28482,
         n28483, n28484, n28485, n28486, n28487, n28488, n28489, n28490,
         n28491, n28492, n28493, n28494, n28495, n28496, n28497, n28498,
         n28499, n28500, n28501, n28502, n28503, n28504, n28505, n28506,
         n28507, n28508, n28509, n28510, n28511, n28512, n28513, n28514,
         n28515, n28516, n28517, n28518, n28519, n28520, n28521, n28522,
         n28523, n28524, n28525, n28526, n28527, n28528, n28529, n28530,
         n28531, n28532, n28533, n28534, n28535, n28536, n28537, n28538,
         n28539, n28540, n28541, n28542, n28543, n28544, n28545, n28546,
         n28547, n28548, n28549, n28550, n28551, n28552, n28553, n28554,
         n28555, n28556, n28557, n28558, n28559, n28560, n28561, n28562,
         n28563, n28564, n28565, n28566, n28567, n28568, n28569, n28570,
         n28571, n28572, n28573, n28574, n28575, n28576, n28577, n28578,
         n28579, n28580, n28581, n28582, n28583, n28584, n28585, n28586,
         n28587, n28588, n28589, n28590, n28591, n28592, n28593, n28594,
         n28595, n28596, n28597, n28598, n28599, n28600, n28601, n28602,
         n28603, n28604, n28605, n28606, n28607, n28608, n28609, n28610,
         n28611, n28612, n28613, n28614, n28615, n28616, n28617, n28618,
         n28619, n28620, n28621, n28622, n28623, n28624, n28625, n28626,
         n28627, n28628, n28629, n28630, n28631, n28632, n28633, n28634,
         n28635, n28636, n28637, n28638, n28639, n28640, n28641, n28642,
         n28643, n28644, n28645, n28646, n28647, n28648, n28649, n28650,
         n28651, n28652, n28653, n28654, n28655, n28656, n28657, n28658,
         n28659, n28660, n28661, n28662, n28663, n28664, n28665, n28666,
         n28667, n28668, n28669, n28670, n28671, n28672, n28673, n28674,
         n28675, n28676, n28677, n28678, n28679, n28680, n28681, n28682,
         n28683, n28684, n28685, n28686, n28687, n28688, n28689, n28690,
         n28691, n28692, n28693, n28694, n28695, n28696, n28697, n28698,
         n28699, n28700, n28701, n28702, n28703, n28704, n28705, n28706,
         n28707, n28708, n28709, n28710, n28711, n28712, n28713, n28714,
         n28715, n28716, n28717, n28718, n28719, n28720, n28721, n28722,
         n28723, n28724, n28725, n28726, n28727, n28728, n28729, n28730,
         n28731, n28732, n28733, n28734, n28735, n28736, n28737, n28738,
         n28739, n28740, n28741, n28742, n28743, n28744, n28745, n28746,
         n28747, n28748, n28749, n28750, n28751, n28752, n28753, n28754,
         n28755, n28756, n28757, n28758, n28759, n28760, n28761, n28762,
         n28763, n28764, n28765, n28766, n28767, n28768, n28769, n28770,
         n28771, n28772, n28773, n28774, n28775, n28776, n28777, n28778,
         n28779, n28780, n28781, n28782, n28783, n28784, n28785, n28786,
         n28787, n28788, n28789, n28790, n28791, n28792, n28793, n28794,
         n28795, n28796, n28797, n28798, n28799, n28800, n28801, n28802,
         n28803, n28804, n28805, n28806, n28807, n28808, n28809, n28810,
         n28811, n28812, n28813, n28814, n28815, n28816, n28817, n28818,
         n28819, n28820, n28821, n28822, n28823, n28824, n28825, n28826,
         n28827, n28828, n28829, n28830, n28831, n28832, n28833, n28834,
         n28835, n28836, n28837, n28838, n28839, n28840, n28841, n28842,
         n28843, n28844, n28845, n28846, n28847, n28848, n28849, n28850,
         n28851, n28852, n28853, n28854, n28855, n28856, n28857, n28858,
         n28859, n28860, n28861, n28862, n28863, n28864, n28865, n28866,
         n28867, n28868, n28869, n28870, n28871, n28872, n28873, n28874,
         n28875, n28876, n28877, n28878, n28879, n28880, n28881, n28882,
         n28883, n28884, n28885, n28886, n28887, n28888, n28889, n28890,
         n28891, n28892, n28893, n28894, n28895, n28896, n28897, n28898,
         n28899, n28900, n28901, n28902, n28903, n28904, n28905, n28906,
         n28907, n28908, n28909, n28910, n28911, n28912, n28913, n28914,
         n28915, n28916, n28917, n28918, n28919, n28920, n28921, n28922,
         n28923, n28924, n28925, n28926, n28927, n28928, n28929, n28930,
         n28931, n28932, n28933, n28934, n28935, n28936, n28937, n28938,
         n28939, n28940, n28941, n28942, n28943, n28944, n28945, n28946,
         n28947, n28948, n28949, n28950, n28951, n28952, n28953, n28954,
         n28955, n28956, n28957, n28958, n28959, n28960, n28961, n28962,
         n28963, n28964, n28965, n28966, n28967, n28968, n28969, n28970,
         n28971, n28972, n28973, n28974, n28975, n28976, n28977, n28978,
         n28979, n28980, n28981, n28982, n28983, n28984, n28985, n28986,
         n28987, n28988, n28989, n28990, n28991, n28992, n28993, n28994,
         n28995, n28996, n28997, n28998, n28999, n29000, n29001, n29002,
         n29003, n29004, n29005, n29006, n29007, n29008, n29009, n29010,
         n29011, n29012, n29013, n29014, n29015, n29016, n29017, n29018,
         n29019, n29020, n29021, n29022, n29023, n29024, n29025, n29026,
         n29027, n29028, n29029, n29030, n29031, n29032, n29033, n29034,
         n29035, n29036, n29037, n29038, n29039, n29040, n29041, n29042,
         n29043, n29044, n29045, n29046, n29047, n29048, n29049, n29050,
         n29051, n29052, n29053, n29054, n29055, n29056, n29057, n29058,
         n29059, n29060, n29061, n29062, n29063, n29064, n29065, n29066,
         n29067, n29068, n29069, n29070, n29071, n29072, n29073, n29074,
         n29075, n29076, n29077, n29078, n29079, n29080, n29081, n29082,
         n29083, n29084, n29085, n29086, n29087, n29088, n29089, n29090,
         n29091, n29092, n29093, n29094, n29095, n29096, n29097, n29098,
         n29099, n29100, n29101, n29102, n29103, n29104, n29105, n29106,
         n29107, n29108, n29109, n29110, n29111, n29112, n29113, n29114,
         n29115, n29116, n29117, n29118, n29119, n29120, n29121, n29122,
         n29123, n29124, n29125, n29126, n29127, n29128, n29129, n29130,
         n29131, n29132, n29133, n29134, n29135, n29136, n29137, n29138,
         n29139, n29140, n29141, n29142, n29143, n29144, n29145, n29146,
         n29147, n29148, n29149, n29150, n29151, n29152, n29153, n29154,
         n29155, n29156, n29157, n29158, n29159, n29160, n29161, n29162,
         n29163, n29164, n29165, n29166, n29167, n29168, n29169, n29170,
         n29171, n29172, n29173, n29174, n29175, n29176, n29177, n29178,
         n29179, n29180, n29181, n29182, n29183, n29184, n29185, n29186,
         n29187, n29188, n29189, n29190, n29191, n29192, n29193, n29194,
         n29195, n29196, n29197, n29198, n29199, n29200, n29201, n29202,
         n29203, n29204, n29205, n29206, n29207, n29208, n29209, n29210,
         n29211, n29212, n29213, n29214, n29215, n29216, n29217, n29218,
         n29219, n29220, n29221, n29222, n29223, n29224, n29225, n29226,
         n29227, n29228, n29229, n29230, n29231, n29232, n29233, n29234,
         n29235, n29236, n29237, n29238, n29239, n29240, n29241, n29242,
         n29243, n29244, n29245, n29246, n29247, n29248, n29249, n29250,
         n29251, n29252, n29253, n29254, n29255, n29256, n29257, n29258,
         n29259, n29260, n29261, n29262, n29263, n29264, n29265, n29266,
         n29267, n29268, n29269, n29270, n29271, n29272, n29273, n29274,
         n29275, n29276, n29277, n29278, n29279, n29280, n29281, n29282,
         n29283, n29284, n29285, n29286, n29287, n29288, n29289, n29290,
         n29291, n29292, n29293, n29294, n29295, n29296, n29297, n29298,
         n29299, n29300, n29301, n29302, n29303, n29304, n29305, n29306,
         n29307, n29308, n29309, n29310, n29311, n29312, n29313, n29314,
         n29315, n29316, n29317, n29318, n29319, n29320, n29321, n29322,
         n29323, n29324, n29325, n29326, n29327, n29328, n29329, n29330,
         n29331, n29332, n29333, n29334, n29335, n29336, n29337, n29338,
         n29339, n29340, n29341, n29342, n29343, n29344, n29345, n29346,
         n29347, n29348, n29349, n29350, n29351, n29352, n29353, n29354,
         n29355, n29356, n29357, n29358, n29359, n29360, n29361, n29362,
         n29363, n29364, n29365, n29366, n29367, n29368, n29369, n29370,
         n29371, n29372, n29373, n29374, n29375, n29376, n29377, n29378,
         n29379, n29380, n29381, n29382, n29383, n29384, n29385, n29386,
         n29387, n29388, n29389, n29390, n29391, n29392, n29393, n29394,
         n29395, n29396, n29397, n29398, n29399, n29400, n29401, n29402,
         n29403, n29404, n29405, n29406, n29407, n29408, n29409, n29410,
         n29411, n29412, n29413, n29414, n29415, n29416, n29417, n29418,
         n29419, n29420, n29421, n29422, n29423, n29424, n29425, n29426,
         n29427, n29428, n29429, n29430, n29431, n29432, n29433, n29434,
         n29435, n29436, n29437, n29438, n29439, n29440, n29441, n29442,
         n29443, n29444, n29445, n29446, n29447, n29448, n29449, n29450,
         n29451, n29452, n29453, n29454, n29455, n29456, n29457, n29458,
         n29459, n29460, n29461, n29462, n29463, n29464, n29465, n29466,
         n29467, n29468, n29469, n29470, n29471, n29472, n29473, n29474,
         n29475, n29476, n29477, n29478, n29479, n29480, n29481, n29482,
         n29483, n29484, n29485, n29486, n29487, n29488, n29489, n29490,
         n29491, n29492, n29493, n29494, n29495, n29496, n29497, n29498,
         n29499, n29500, n29501, n29502, n29503, n29504, n29505, n29506,
         n29507, n29508, n29509, n29510, n29511, n29512, n29513, n29514,
         n29515, n29516, n29517, n29518, n29519, n29520, n29521, n29522,
         n29523, n29524, n29525, n29526, n29527, n29528, n29529, n29530,
         n29531, n29532, n29533, n29534, n29535, n29536, n29537, n29538,
         n29539, n29540, n29541, n29542, n29543, n29544, n29545, n29546,
         n29547, n29548, n29549, n29550, n29551, n29552, n29553, n29554,
         n29555, n29556, n29557, n29558, n29559, n29560, n29561, n29562,
         n29563, n29564, n29565, n29566, n29567, n29568, n29569, n29570,
         n29571, n29572, n29573, n29574, n29575, n29576, n29577, n29578,
         n29579, n29580, n29581, n29582, n29583, n29584, n29585, n29586,
         n29587, n29588, n29589, n29590, n29591, n29592, n29593, n29594,
         n29595, n29596, n29597, n29598, n29599, n29600, n29601, n29602,
         n29603, n29604, n29605, n29606, n29607, n29608, n29609, n29610,
         n29611, n29612, n29613, n29614, n29615, n29616, n29617, n29618,
         n29619, n29620, n29621, n29622, n29623, n29624, n29625, n29626,
         n29627, n29628, n29629, n29630, n29631, n29632, n29633, n29634,
         n29635, n29636, n29637, n29638, n29639, n29640, n29641, n29642,
         n29643, n29644, n29645, n29646, n29647, n29648, n29649, n29650,
         n29651, n29652, n29653, n29654, n29655, n29656, n29657, n29658,
         n29659, n29660, n29661, n29662, n29663, n29664, n29665, n29666,
         n29667, n29668, n29669, n29670, n29671, n29672, n29673, n29674,
         n29675, n29676, n29677, n29678, n29679, n29680, n29681, n29682,
         n29683, n29684, n29685, n29686, n29687, n29688, n29689, n29690,
         n29691, n29692, n29693, n29694, n29695, n29696, n29697, n29698,
         n29699, n29700, n29701, n29702, n29703, n29704, n29705, n29706,
         n29707, n29708, n29709, n29710, n29711, n29712, n29713, n29714,
         n29715, n29716, n29717, n29718, n29719, n29720, n29721, n29722,
         n29723, n29724, n29725, n29726, n29727, n29728, n29729, n29730,
         n29731, n29732, n29733, n29734, n29735, n29736, n29737, n29738,
         n29739, n29740, n29741, n29742, n29743, n29744, n29745, n29746,
         n29747, n29748, n29749, n29750, n29751, n29752, n29753, n29754,
         n29755, n29756, n29757, n29758, n29759, n29760, n29761, n29762,
         n29763, n29764, n29765, n29766, n29767, n29768, n29769, n29770,
         n29771, n29772, n29773, n29774, n29775, n29776, n29777, n29778,
         n29779, n29780, n29781, n29782, n29783, n29784, n29785, n29786,
         n29787, n29788, n29789, n29790, n29791, n29792, n29793, n29794,
         n29795, n29796, n29797, n29798, n29799, n29800, n29801, n29802,
         n29803, n29804, n29805, n29806, n29807, n29808, n29809, n29810,
         n29811, n29812, n29813, n29814, n29815, n29816, n29817, n29818,
         n29819, n29820, n29821, n29822, n29823, n29824, n29825, n29826,
         n29827, n29828, n29829, n29830, n29831, n29832, n29833, n29834,
         n29835, n29836, n29837, n29838, n29839, n29840, n29841, n29842,
         n29843, n29844, n29845, n29846, n29847, n29848, n29849, n29850,
         n29851, n29852, n29853, n29854, n29855, n29856, n29857, n29858,
         n29859, n29860, n29861, n29862, n29863, n29864, n29865, n29866,
         n29867, n29868, n29869, n29870, n29871, n29872, n29873, n29874,
         n29875, n29876, n29877, n29878, n29879, n29880, n29881, n29882,
         n29883, n29884, n29885, n29886, n29887, n29888, n29889, n29890,
         n29891, n29892, n29893, n29894, n29895, n29896, n29897, n29898,
         n29899, n29900, n29901, n29902, n29903, n29904, n29905, n29906,
         n29907, n29908, n29909, n29910, n29911, n29912, n29913, n29914,
         n29915, n29916, n29917, n29918, n29919, n29920, n29921, n29922,
         n29923, n29924, n29925, n29926, n29927, n29928, n29929, n29930,
         n29931, n29932, n29933, n29934, n29935, n29936, n29937, n29938,
         n29939, n29940, n29941, n29942, n29943, n29944, n29945, n29946,
         n29947, n29948, n29949, n29950, n29951, n29952, n29953, n29954,
         n29955, n29956, n29957, n29958, n29959, n29960, n29961, n29962,
         n29963, n29964, n29965, n29966, n29967, n29968, n29969, n29970,
         n29971, n29972, n29973, n29974, n29975, n29976, n29977, n29978,
         n29979, n29980, n29981, n29982, n29983, n29984, n29985, n29986,
         n29987, n29988, n29989, n29990, n29991, n29992, n29993, n29994,
         n29995, n29996, n29997, n29998, n29999, n30000, n30001, n30002,
         n30003, n30004, n30005, n30006, n30007, n30008, n30009, n30010,
         n30011, n30012, n30013, n30014, n30015, n30016, n30017, n30018,
         n30019, n30020, n30021, n30022, n30023, n30024, n30025, n30026,
         n30027, n30028, n30029, n30030, n30031, n30032, n30033, n30034,
         n30035, n30036, n30037, n30038, n30039, n30040, n30041, n30042,
         n30043, n30044, n30045, n30046, n30047, n30048, n30049, n30050,
         n30051, n30052, n30053, n30054, n30055, n30056, n30057, n30058,
         n30059, n30060, n30061, n30062, n30063, n30064, n30065, n30066,
         n30067, n30068, n30069, n30070, n30071, n30072, n30073, n30074,
         n30075, n30076, n30077, n30078, n30079, n30080, n30081, n30082,
         n30083, n30084, n30085, n30086, n30087, n30088, n30089, n30090,
         n30091, n30092, n30093, n30094, n30095, n30096, n30097, n30098,
         n30099, n30100, n30101, n30102, n30103, n30104, n30105, n30106,
         n30107, n30108, n30109, n30110, n30111, n30112, n30113, n30114,
         n30115, n30116, n30117, n30118, n30119, n30120, n30121, n30122,
         n30123, n30124, n30125, n30126, n30127, n30128, n30129, n30130,
         n30131, n30132, n30133, n30134, n30135, n30136, n30137, n30138,
         n30139, n30140, n30141, n30142, n30143, n30144, n30145, n30146,
         n30147, n30148, n30149, n30150, n30151, n30152, n30153, n30154,
         n30155, n30156, n30157, n30158, n30159, n30160, n30161, n30162,
         n30163, n30164, n30165, n30166, n30167, n30168, n30169, n30170,
         n30171, n30172, n30173, n30174, n30175, n30176, n30177, n30178,
         n30179, n30180, n30181, n30182, n30183, n30184, n30185, n30186,
         n30187, n30188, n30189, n30190, n30191, n30192, n30193, n30194,
         n30195, n30196, n30197, n30198, n30199, n30200, n30201, n30202,
         n30203, n30204, n30205, n30206, n30207, n30208, n30209, n30210,
         n30211, n30212, n30213, n30214, n30215, n30216, n30217, n30218,
         n30219, n30220, n30221, n30222, n30223, n30224, n30225, n30226,
         n30227, n30228, n30229, n30230, n30231, n30232, n30233, n30234,
         n30235, n30236, n30237, n30238, n30239, n30240, n30241, n30242,
         n30243, n30244, n30245, n30246, n30247, n30248, n30249, n30250,
         n30251, n30252, n30253, n30254, n30255, n30256, n30257, n30258,
         n30259, n30260, n30261, n30262, n30263, n30264, n30265, n30266,
         n30267, n30268, n30269, n30270, n30271, n30272, n30273, n30274,
         n30275, n30276, n30277, n30278, n30279, n30280, n30281, n30282,
         n30283, n30284, n30285, n30286, n30287, n30288, n30289, n30290,
         n30291, n30292, n30293, n30294, n30295, n30296, n30297, n30298,
         n30299, n30300, n30301, n30302, n30303, n30304, n30305, n30306,
         n30307, n30308, n30309, n30310, n30311, n30312, n30313, n30314,
         n30315, n30316, n30317, n30318, n30319, n30320, n30321, n30322,
         n30323, n30324, n30325, n30326, n30327, n30328, n30329, n30330,
         n30331, n30332, n30333, n30334, n30335, n30336, n30337, n30338,
         n30339, n30340, n30341, n30342, n30343, n30344, n30345, n30346,
         n30347, n30348, n30349, n30350, n30351, n30352, n30353, n30354,
         n30355, n30356, n30357, n30358, n30359, n30360, n30361, n30362,
         n30363, n30364, n30365, n30366, n30367, n30368, n30369, n30370,
         n30371, n30372, n30373, n30374, n30375, n30376, n30377, n30378,
         n30379, n30380, n30381, n30382, n30383, n30384, n30385, n30386,
         n30387, n30388, n30389, n30390, n30391, n30392, n30393, n30394,
         n30395, n30396, n30397, n30398, n30399, n30400, n30401, n30402,
         n30403, n30404, n30405, n30406, n30407, n30408, n30409, n30410,
         n30411, n30412, n30413, n30414, n30415, n30416, n30417, n30418,
         n30419, n30420, n30421, n30422, n30423, n30424, n30425, n30426,
         n30427, n30428, n30429, n30430, n30431, n30432, n30433, n30434,
         n30435, n30436, n30437, n30438, n30439, n30440, n30441, n30442,
         n30443, n30444, n30445, n30446, n30447, n30448, n30449, n30450,
         n30451, n30452, n30453, n30454, n30455, n30456, n30457, n30458,
         n30459, n30460, n30461, n30462, n30463, n30464, n30465, n30466,
         n30467, n30468, n30469, n30470, n30471, n30472, n30473, n30474,
         n30475, n30476, n30477, n30478, n30479, n30480, n30481, n30482,
         n30483, n30484, n30485, n30486, n30487, n30488, n30489, n30490,
         n30491, n30492, n30493, n30494, n30495, n30496, n30497, n30498,
         n30499, n30500, n30501, n30502, n30503, n30504, n30505, n30506,
         n30507, n30508, n30509, n30510, n30511, n30512, n30513, n30514,
         n30515, n30516, n30517, n30518, n30519, n30520, n30521, n30522,
         n30523, n30524, n30525, n30526, n30527, n30528, n30529, n30530,
         n30531, n30532, n30533, n30534, n30535, n30536, n30537, n30538,
         n30539, n30540, n30541, n30542, n30543, n30544, n30545, n30546,
         n30547, n30548, n30549, n30550, n30551, n30552, n30553, n30554,
         n30555, n30556, n30557, n30558, n30559, n30560, n30561, n30562,
         n30563, n30564, n30565, n30566, n30567, n30568, n30569, n30570,
         n30571, n30572, n30573, n30574, n30575, n30576, n30577, n30578,
         n30579, n30580, n30581, n30582, n30583, n30584, n30585, n30586,
         n30587, n30588, n30589, n30590, n30591, n30592, n30593, n30594,
         n30595, n30596, n30597, n30598, n30599, n30600, n30601, n30602,
         n30603, n30604, n30605, n30606, n30607, n30608, n30609, n30610,
         n30611, n30612, n30613, n30614, n30615, n30616, n30617, n30618,
         n30619, n30620, n30621, n30622, n30623, n30624, n30625, n30626,
         n30627, n30628, n30629, n30630, n30631, n30632, n30633, n30634,
         n30635, n30636, n30637, n30638, n30639, n30640, n30641, n30642,
         n30643, n30644, n30645, n30646, n30647, n30648, n30649, n30650,
         n30651, n30652, n30653, n30654, n30655, n30656, n30657, n30658,
         n30659, n30660, n30661, n30662, n30663, n30664, n30665, n30666,
         n30667, n30668, n30669, n30670, n30671, n30672, n30673, n30674,
         n30675, n30676, n30677, n30678, n30679, n30680, n30681, n30682,
         n30683, n30684, n30685, n30686, n30687, n30688, n30689, n30690,
         n30691, n30692, n30693, n30694, n30695, n30696, n30697, n30698,
         n30699, n30700, n30701, n30702, n30703, n30704, n30705, n30706,
         n30707, n30708, n30709, n30710, n30711, n30712, n30713, n30714,
         n30715, n30716, n30717, n30718, n30719, n30720, n30721, n30722,
         n30723, n30724, n30725, n30726, n30727, n30728, n30729, n30730,
         n30731, n30732, n30733, n30734, n30735, n30736, n30737, n30738,
         n30739, n30740, n30741, n30742, n30743, n30744, n30745, n30746,
         n30747, n30748, n30749, n30750, n30751, n30752, n30753, n30754,
         n30755, n30756, n30757, n30758, n30759, n30760, n30761, n30762,
         n30763, n30764, n30765, n30766, n30767, n30768, n30769, n30770,
         n30771, n30772, n30773, n30774, n30775, n30776, n30777, n30778,
         n30779, n30780, n30781, n30782, n30783, n30784, n30785, n30786,
         n30787, n30788, n30789, n30790, n30791, n30792, n30793, n30794,
         n30795, n30796, n30797, n30798, n30799, n30800, n30801, n30802,
         n30803, n30804, n30805, n30806, n30807, n30808, n30809, n30810,
         n30811, n30812, n30813, n30814, n30815, n30816, n30817, n30818,
         n30819, n30820, n30821, n30822, n30823, n30824, n30825, n30826,
         n30827, n30828, n30829, n30830, n30831, n30832, n30833, n30834,
         n30835, n30836, n30837, n30838, n30839, n30840, n30841, n30842,
         n30843, n30844, n30845, n30846, n30847, n30848, n30849, n30850,
         n30851, n30852, n30853, n30854, n30855, n30856, n30857, n30858,
         n30859, n30860, n30861, n30862, n30863, n30864, n30865, n30866,
         n30867, n30868, n30869, n30870, n30871, n30872, n30873, n30874,
         n30875, n30876, n30877, n30878, n30879, n30880, n30881, n30882,
         n30883, n30884, n30885, n30886, n30887, n30888, n30889, n30890,
         n30891, n30892, n30893, n30894, n30895, n30896, n30897, n30898,
         n30899, n30900, n30901, n30902, n30903, n30904, n30905, n30906,
         n30907, n30908, n30909, n30910, n30911, n30912, n30913, n30914,
         n30915, n30916, n30917, n30918, n30919, n30920, n30921, n30922,
         n30923, n30924, n30925, n30926, n30927, n30928, n30929, n30930,
         n30931, n30932, n30933, n30934, n30935, n30936, n30937, n30938,
         n30939, n30940, n30941, n30942, n30943, n30944, n30945, n30946,
         n30947, n30948, n30949, n30950, n30951, n30952, n30953, n30954,
         n30955, n30956, n30957, n30958, n30959, n30960, n30961, n30962,
         n30963, n30964, n30965, n30966, n30967, n30968, n30969, n30970,
         n30971, n30972, n30973, n30974, n30975, n30976, n30977, n30978,
         n30979, n30980, n30981, n30982, n30983, n30984, n30985, n30986,
         n30987, n30988, n30989, n30990, n30991, n30992, n30993, n30994,
         n30995, n30996, n30997, n30998, n30999, n31000, n31001, n31002,
         n31003, n31004, n31005, n31006, n31007, n31008, n31009, n31010,
         n31011, n31012, n31013, n31014, n31015, n31016, n31017, n31018,
         n31019, n31020, n31021, n31022, n31023, n31024, n31025, n31026,
         n31027, n31028, n31029, n31030, n31031, n31032, n31033, n31034,
         n31035, n31036, n31037, n31038, n31039, n31040, n31041, n31042,
         n31043, n31044, n31045, n31046, n31047, n31048, n31049, n31050,
         n31051, n31052, n31053, n31054, n31055, n31056, n31057, n31058,
         n31059, n31060, n31061, n31062, n31063, n31064, n31065, n31066,
         n31067, n31068, n31069, n31070, n31071, n31072, n31073, n31074,
         n31075, n31076, n31077, n31078, n31079, n31080, n31081, n31082,
         n31083, n31084, n31085, n31086, n31087, n31088, n31089, n31090,
         n31091, n31092, n31093, n31094, n31095, n31096, n31097, n31098,
         n31099, n31100, n31101, n31102, n31103, n31104, n31105, n31106,
         n31107, n31108, n31109, n31110, n31111, n31112, n31113, n31114,
         n31115, n31116, n31117, n31118, n31119, n31120, n31121, n31122,
         n31123, n31124, n31125, n31126, n31127, n31128, n31129, n31130,
         n31131, n31132, n31133, n31134, n31135, n31136, n31137, n31138,
         n31139, n31140, n31141, n31142, n31143, n31144, n31145, n31146,
         n31147, n31148, n31149, n31150, n31151, n31152, n31153, n31154,
         n31155, n31156, n31157, n31158, n31159, n31160, n31161, n31162,
         n31163, n31164, n31165, n31166, n31167, n31168, n31169, n31170,
         n31171, n31172, n31173, n31174, n31175, n31176, n31177, n31178,
         n31179, n31180, n31181, n31182, n31183, n31184, n31185, n31186,
         n31187, n31188, n31189, n31190, n31191, n31192, n31193, n31194,
         n31195, n31196, n31197, n31198, n31199, n31200, n31201, n31202,
         n31203, n31204, n31205, n31206, n31207, n31208, n31209, n31210,
         n31211, n31212, n31213, n31214, n31215, n31216, n31217, n31218,
         n31219, n31220, n31221, n31222, n31223, n31224, n31225, n31226,
         n31227, n31228, n31229, n31230, n31231, n31232, n31233, n31234,
         n31235, n31236, n31237, n31238, n31239, n31240, n31241, n31242,
         n31243, n31244, n31245, n31246, n31247, n31248, n31249, n31250,
         n31251, n31252, n31253, n31254, n31255, n31256, n31257, n31258,
         n31259, n31260, n31261, n31262, n31263, n31264, n31265, n31266,
         n31267, n31268, n31269, n31270, n31271, n31272, n31273, n31274,
         n31275, n31276, n31277, n31278, n31279, n31280, n31281, n31282,
         n31283, n31284, n31285, n31286, n31287, n31288, n31289, n31290,
         n31291, n31292, n31293, n31294, n31295, n31296, n31297, n31298,
         n31299, n31300, n31301, n31302, n31303, n31304, n31305, n31306,
         n31307, n31308, n31309, n31310, n31311, n31312, n31313, n31314,
         n31315, n31316, n31317, n31318, n31319, n31320, n31321, n31322,
         n31323, n31324, n31325, n31326, n31327, n31328, n31329, n31330,
         n31331, n31332, n31333, n31334, n31335, n31336, n31337, n31338,
         n31339, n31340, n31341, n31342, n31343, n31344, n31345, n31346,
         n31347, n31348, n31349, n31350, n31351, n31352, n31353, n31354,
         n31355, n31356, n31357, n31358, n31359, n31360, n31361, n31362,
         n31363, n31364, n31365, n31366, n31367, n31368, n31369, n31370,
         n31371, n31372, n31373, n31374, n31375, n31376, n31377, n31378,
         n31379, n31380, n31381, n31382, n31383, n31384, n31385, n31386,
         n31387, n31388, n31389, n31390, n31391, n31392, n31393, n31394,
         n31395, n31396, n31397, n31398, n31399, n31400, n31401, n31402,
         n31403, n31404, n31405, n31406, n31407, n31408, n31409, n31410,
         n31411, n31412, n31413, n31414, n31415, n31416, n31417, n31418,
         n31419, n31420, n31421, n31422, n31423, n31424, n31425, n31426,
         n31427, n31428, n31429, n31430, n31431, n31432, n31433, n31434,
         n31435, n31436, n31437, n31438, n31439, n31440, n31441, n31442,
         n31443, n31444, n31445, n31446, n31447, n31448, n31449, n31450,
         n31451, n31452, n31453, n31454, n31455, n31456, n31457, n31458,
         n31459, n31460, n31461, n31462, n31463, n31464, n31465, n31466,
         n31467, n31468, n31469, n31470, n31471, n31472, n31473, n31474,
         n31475, n31476, n31477, n31478, n31479, n31480, n31481, n31482,
         n31483, n31484, n31485, n31486, n31487, n31488, n31489, n31490,
         n31491, n31492, n31493, n31494, n31495, n31496, n31497, n31498,
         n31499, n31500, n31501, n31502, n31503, n31504, n31505, n31506,
         n31507, n31508, n31509, n31510, n31511, n31512, n31513, n31514,
         n31515, n31516, n31517, n31518, n31519, n31520, n31521, n31522,
         n31523, n31524, n31525, n31526, n31527, n31528, n31529, n31530,
         n31531, n31532, n31533, n31534, n31535, n31536, n31537, n31538,
         n31539, n31540, n31541, n31542, n31543, n31544, n31545, n31546,
         n31547, n31548, n31549, n31550, n31551, n31552, n31553, n31554,
         n31555, n31556, n31557, n31558, n31559, n31560, n31561, n31562,
         n31563, n31564, n31565, n31566, n31567, n31568, n31569, n31570,
         n31571, n31572, n31573, n31574, n31575, n31576, n31577, n31578,
         n31579, n31580, n31581, n31582, n31583, n31584, n31585, n31586,
         n31587, n31588, n31589, n31590, n31591, n31592, n31593, n31594,
         n31595, n31596, n31597, n31598, n31599, n31600, n31601, n31602,
         n31603, n31604, n31605, n31606, n31607, n31608, n31609, n31610,
         n31611, n31612, n31613, n31614, n31615, n31616, n31617, n31618,
         n31619, n31620, n31621, n31622, n31623, n31624, n31625, n31626,
         n31627, n31628, n31629, n31630, n31631, n31632, n31633, n31634,
         n31635, n31636, n31637, n31638, n31639, n31640, n31641, n31642,
         n31643, n31644, n31645, n31646, n31647, n31648, n31649, n31650,
         n31651, n31652, n31653, n31654, n31655, n31656, n31657, n31658,
         n31659, n31660, n31661, n31662, n31663, n31664, n31665, n31666,
         n31667, n31668, n31669, n31670, n31671, n31672, n31673, n31674,
         n31675, n31676, n31677, n31678, n31679, n31680, n31681, n31682,
         n31683, n31684, n31685, n31686, n31687, n31688, n31689, n31690,
         n31691, n31692, n31693, n31694, n31695, n31696, n31697, n31698,
         n31699, n31700, n31701, n31702, n31703, n31704, n31705, n31706,
         n31707, n31708, n31709, n31710, n31711, n31712, n31713, n31714,
         n31715, n31716, n31717, n31718, n31719, n31720, n31721, n31722,
         n31723, n31724, n31725, n31726, n31727, n31728, n31729, n31730,
         n31731, n31732, n31733, n31734, n31735, n31736, n31737, n31738,
         n31739, n31740, n31741, n31742, n31743, n31744, n31745, n31746,
         n31747, n31748, n31749, n31750, n31751, n31752, n31753, n31754,
         n31755, n31756, n31757, n31758, n31759, n31760, n31761, n31762,
         n31763, n31764, n31765, n31766, n31767, n31768, n31769, n31770,
         n31771, n31772, n31773, n31774, n31775, n31776, n31777, n31778,
         n31779, n31780, n31781, n31782, n31783, n31784, n31785, n31786,
         n31787, n31788, n31789, n31790, n31791, n31792, n31793, n31794,
         n31795, n31796, n31797, n31798, n31799, n31800, n31801, n31802,
         n31803, n31804, n31805, n31806, n31807, n31808, n31809, n31810,
         n31811, n31812, n31813, n31814, n31815, n31816, n31817, n31818,
         n31819, n31820, n31821, n31822, n31823, n31824, n31825, n31826,
         n31827, n31828, n31829, n31830, n31831, n31832, n31833, n31834,
         n31835, n31836, n31837, n31838, n31839, n31840, n31841, n31842,
         n31843, n31844, n31845, n31846, n31847, n31848, n31849, n31850,
         n31851, n31852, n31853, n31854, n31855, n31856, n31857, n31858,
         n31859, n31860, n31861, n31862, n31863, n31864, n31865, n31866,
         n31867, n31868, n31869, n31870, n31871, n31872, n31873, n31874,
         n31875, n31876, n31877, n31878, n31879, n31880, n31881, n31882,
         n31883, n31884, n31885, n31886, n31887, n31888, n31889, n31890,
         n31891, n31892, n31893, n31894, n31895, n31896, n31897, n31898,
         n31899, n31900, n31901, n31902, n31903, n31904, n31905, n31906,
         n31907, n31908, n31909, n31910, n31911, n31912, n31913, n31914,
         n31915, n31916, n31917, n31918, n31919, n31920, n31921, n31922,
         n31923, n31924, n31925, n31926, n31927, n31928, n31929, n31930,
         n31931, n31932, n31933, n31934, n31935, n31936, n31937, n31938,
         n31939, n31940, n31941, n31942, n31943, n31944, n31945, n31946,
         n31947, n31948, n31949, n31950, n31951, n31952, n31953, n31954,
         n31955, n31956, n31957, n31958, n31959, n31960, n31961, n31962,
         n31963, n31964, n31965, n31966, n31967, n31968, n31969, n31970,
         n31971, n31972, n31973, n31974, n31975, n31976, n31977, n31978,
         n31979, n31980, n31981, n31982, n31983, n31984, n31985, n31986,
         n31987, n31988, n31989, n31990, n31991, n31992, n31993, n31994,
         n31995, n31996, n31997, n31998, n31999, n32000, n32001, n32002,
         n32003, n32004, n32005, n32006, n32007, n32008, n32009, n32010,
         n32011, n32012, n32013, n32014, n32015, n32016, n32017, n32018,
         n32019, n32020, n32021, n32022, n32023, n32024, n32025, n32026,
         n32027, n32028, n32029, n32030, n32031, n32032, n32033, n32034,
         n32035, n32036, n32037, n32038, n32039, n32040, n32041, n32042,
         n32043, n32044, n32045, n32046, n32047, n32048, n32049, n32050,
         n32051, n32052, n32053, n32054, n32055, n32056, n32057, n32058,
         n32059, n32060, n32061, n32062, n32063, n32064, n32065, n32066,
         n32067, n32068, n32069, n32070, n32071, n32072, n32073, n32074,
         n32075, n32076, n32077, n32078, n32079, n32080, n32081, n32082,
         n32083, n32084, n32085, n32086, n32087, n32088, n32089, n32090,
         n32091, n32092, n32093, n32094, n32095, n32096, n32097, n32098,
         n32099, n32100, n32101, n32102, n32103, n32104, n32105, n32106,
         n32107, n32108, n32109, n32110, n32111, n32112, n32113, n32114,
         n32115, n32116, n32117, n32118, n32119, n32120, n32121, n32122,
         n32123, n32124, n32125, n32126, n32127, n32128, n32129, n32130,
         n32131, n32132, n32133, n32134, n32135, n32136, n32137, n32138,
         n32139, n32140, n32141, n32142, n32143, n32144, n32145, n32146,
         n32147, n32148, n32149, n32150, n32151, n32152, n32153, n32154,
         n32155, n32156, n32157, n32158, n32159, n32160, n32161, n32162,
         n32163, n32164, n32165, n32166, n32167, n32168, n32169, n32170,
         n32171, n32172, n32173, n32174, n32175, n32176, n32177, n32178,
         n32179, n32180, n32181, n32182, n32183, n32184, n32185, n32186,
         n32187, n32188, n32189, n32190, n32191, n32192, n32193, n32194,
         n32195, n32196, n32197, n32198, n32199, n32200, n32201, n32202,
         n32203, n32204, n32205, n32206, n32207, n32208, n32209, n32210,
         n32211, n32212, n32213, n32214, n32215, n32216, n32217, n32218,
         n32219, n32220, n32221, n32222, n32223, n32224, n32225, n32226,
         n32227, n32228, n32229, n32230, n32231, n32232, n32233, n32234,
         n32235, n32236, n32237, n32238, n32239, n32240, n32241, n32242,
         n32243, n32244, n32245, n32246, n32247, n32248, n32249, n32250,
         n32251, n32252, n32253, n32254, n32255, n32256, n32257, n32258,
         n32259, n32260, n32261, n32262, n32263, n32264, n32265, n32266,
         n32267, n32268, n32269, n32270, n32271, n32272, n32273, n32274,
         n32275, n32276, n32277, n32278, n32279, n32280, n32281, n32282,
         n32283, n32284, n32285, n32286, n32287, n32288, n32289, n32290,
         n32291, n32292, n32293, n32294, n32295, n32296, n32297, n32298,
         n32299, n32300, n32301, n32302, n32303, n32304, n32305, n32306,
         n32307, n32308, n32309, n32310, n32311, n32312, n32313, n32314,
         n32315, n32316, n32317, n32318, n32319, n32320, n32321, n32322,
         n32323, n32324, n32325, n32326, n32327, n32328, n32329, n32330,
         n32331, n32332, n32333, n32334, n32335, n32336, n32337, n32338,
         n32339, n32340, n32341, n32342, n32343, n32344, n32345, n32346,
         n32347, n32348, n32349, n32350, n32351, n32352, n32353, n32354,
         n32355, n32356, n32357, n32358, n32359, n32360, n32361, n32362,
         n32363, n32364, n32365, n32366, n32367, n32368, n32369, n32370,
         n32371, n32372, n32373, n32374, n32375, n32376, n32377, n32378,
         n32379, n32380, n32381, n32382, n32383, n32384, n32385, n32386,
         n32387, n32388, n32389, n32390, n32391, n32392, n32393, n32394,
         n32395, n32396, n32397, n32398, n32399, n32400, n32401, n32402,
         n32403, n32404, n32405, n32406, n32407, n32408, n32409, n32410,
         n32411, n32412, n32413, n32414, n32415, n32416, n32417, n32418,
         n32419, n32420, n32421, n32422, n32423, n32424, n32425, n32426,
         n32427, n32428, n32429, n32430, n32431, n32432, n32433, n32434,
         n32435, n32436, n32437, n32438, n32439, n32440, n32441, n32442,
         n32443, n32444, n32445, n32446, n32447, n32448, n32449, n32450,
         n32451, n32452, n32453, n32454, n32455, n32456, n32457, n32458,
         n32459, n32460, n32461, n32462, n32463, n32464, n32465, n32466,
         n32467, n32468, n32469, n32470, n32471, n32472, n32473, n32474,
         n32475, n32476, n32477, n32478, n32479, n32480, n32481, n32482,
         n32483, n32484, n32485, n32486, n32487, n32488, n32489, n32490,
         n32491, n32492, n32493, n32494, n32495, n32496, n32497, n32498,
         n32499, n32500, n32501, n32502, n32503, n32504, n32505, n32506,
         n32507, n32508, n32509, n32510, n32511, n32512, n32513, n32514,
         n32515, n32516, n32517, n32518, n32519, n32520, n32521, n32522,
         n32523, n32524, n32525, n32526, n32527, n32528, n32529, n32530,
         n32531, n32532, n32533, n32534, n32535, n32536, n32537, n32538,
         n32539, n32540, n32541, n32542, n32543, n32544, n32545, n32546,
         n32547, n32548, n32549, n32550, n32551, n32552, n32553, n32554,
         n32555, n32556, n32557, n32558, n32559, n32560, n32561, n32562,
         n32563, n32564, n32565, n32566, n32567, n32568, n32569, n32570,
         n32571, n32572, n32573, n32574, n32575, n32576, n32577, n32578,
         n32579, n32580, n32581, n32582, n32583, n32584, n32585, n32586,
         n32587, n32588, n32589, n32590, n32591, n32592, n32593, n32594,
         n32595, n32596, n32597, n32598, n32599, n32600, n32601, n32602,
         n32603, n32604, n32605, n32606, n32607, n32608, n32609, n32610,
         n32611, n32612, n32613, n32614, n32615, n32616, n32617, n32618,
         n32619, n32620, n32621, n32622, n32623, n32624, n32625, n32626,
         n32627, n32628, n32629, n32630, n32631, n32632, n32633, n32634,
         n32635, n32636, n32637, n32638, n32639, n32640, n32641, n32642,
         n32643, n32644, n32645, n32646, n32647, n32648, n32649, n32650,
         n32651, n32652, n32653, n32654, n32655, n32656, n32657, n32658,
         n32659, n32660, n32661, n32662, n32663, n32664, n32665, n32666,
         n32667, n32668, n32669, n32670, n32671, n32672, n32673, n32674,
         n32675, n32676, n32677, n32678, n32679, n32680, n32681, n32682,
         n32683, n32684, n32685, n32686, n32687, n32688, n32689, n32690,
         n32691, n32692, n32693, n32694, n32695, n32696, n32697, n32698,
         n32699, n32700, n32701, n32702, n32703, n32704, n32705, n32706,
         n32707, n32708, n32709, n32710, n32711, n32712, n32713, n32714,
         n32715, n32716, n32717, n32718, n32719, n32720, n32721, n32722,
         n32723, n32724, n32725, n32726, n32727, n32728, n32729, n32730,
         n32731, n32732, n32733, n32734, n32735, n32736, n32737, n32738,
         n32739, n32740, n32741, n32742, n32743, n32744, n32745, n32746,
         n32747, n32748, n32749, n32750, n32751, n32752, n32753, n32754,
         n32755, n32756, n32757, n32758, n32759, n32760, n32761, n32762,
         n32763, n32764, n32765, n32766, n32767, n32768, n32769, n32770,
         n32771, n32772, n32773, n32774, n32775, n32776, n32777, n32778,
         n32779, n32780, n32781, n32782, n32783, n32784, n32785, n32786,
         n32787, n32788, n32789, n32790, n32791, n32792, n32793, n32794,
         n32795, n32796, n32797, n32798, n32799, n32800, n32801, n32802,
         n32803, n32804, n32805, n32806, n32807, n32808, n32809, n32810,
         n32811, n32812, n32813, n32814, n32815, n32816, n32817, n32818,
         n32819, n32820, n32821, n32822, n32823, n32824, n32825, n32826,
         n32827, n32828, n32829, n32830, n32831, n32832, n32833, n32834,
         n32835, n32836, n32837, n32838, n32839, n32840, n32841, n32842,
         n32843, n32844, n32845, n32846, n32847, n32848, n32849, n32850,
         n32851, n32852, n32853, n32854, n32855, n32856, n32857, n32858,
         n32859, n32860, n32861, n32862, n32863, n32864, n32865, n32866,
         n32867, n32868, n32869, n32870, n32871, n32872, n32873, n32874,
         n32875, n32876, n32877, n32878, n32879, n32880, n32881, n32882,
         n32883, n32884, n32885, n32886, n32887, n32888, n32889, n32890,
         n32891, n32892, n32893, n32894, n32895, n32896, n32897, n32898,
         n32899, n32900, n32901, n32902, n32903, n32904, n32905, n32906,
         n32907, n32908, n32909, n32910, n32911, n32912, n32913, n32914,
         n32915, n32916, n32917, n32918, n32919, n32920, n32921, n32922,
         n32923, n32924, n32925, n32926, n32927, n32928, n32929, n32930,
         n32931, n32932, n32933, n32934, n32935, n32936, n32937, n32938,
         n32939, n32940, n32941, n32942, n32943, n32944, n32945, n32946,
         n32947, n32948, n32949, n32950, n32951, n32952, n32953, n32954,
         n32955, n32956, n32957, n32958, n32959, n32960, n32961, n32962,
         n32963, n32964, n32965, n32966, n32967, n32968, n32969, n32970,
         n32971, n32972, n32973, n32974, n32975, n32976, n32977, n32978,
         n32979, n32980, n32981, n32982, n32983, n32984, n32985, n32986,
         n32987, n32988, n32989, n32990, n32991, n32992, n32993, n32994,
         n32995, n32996, n32997, n32998, n32999, n33000, n33001, n33002,
         n33003, n33004, n33005, n33006, n33007, n33008, n33009, n33010,
         n33011, n33012, n33013, n33014, n33015, n33016, n33017, n33018,
         n33019, n33020, n33021, n33022, n33023, n33024, n33025, n33026,
         n33027, n33028, n33029, n33030, n33031, n33032, n33033, n33034,
         n33035, n33036, n33037, n33038, n33039, n33040, n33041, n33042,
         n33043, n33044, n33045, n33046, n33047, n33048, n33049, n33050,
         n33051, n33052, n33053, n33054, n33055, n33056, n33057, n33058,
         n33059, n33060, n33061, n33062, n33063, n33064, n33065, n33066,
         n33067, n33068, n33069, n33070, n33071, n33072, n33073, n33074,
         n33075, n33076, n33077, n33078, n33079, n33080, n33081, n33082,
         n33083, n33084, n33085, n33086, n33087, n33088, n33089, n33090,
         n33091, n33092, n33093, n33094, n33095, n33096, n33097, n33098,
         n33099, n33100, n33101, n33102, n33103, n33104, n33105, n33106,
         n33107, n33108, n33109, n33110, n33111, n33112, n33113, n33114,
         n33115, n33116, n33117, n33118, n33119, n33120, n33121, n33122,
         n33123, n33124, n33125, n33126, n33127, n33128, n33129, n33130,
         n33131, n33132, n33133, n33134, n33135, n33136, n33137, n33138,
         n33139, n33140, n33141, n33142, n33143, n33144, n33145, n33146,
         n33147, n33148, n33149, n33150, n33151, n33152, n33153, n33154,
         n33155, n33156, n33157, n33158, n33159, n33160, n33161, n33162,
         n33163, n33164, n33165, n33166, n33167, n33168, n33169, n33170,
         n33171, n33172, n33173, n33174, n33175, n33176, n33177, n33178,
         n33179, n33180, n33181, n33182, n33183, n33184, n33185, n33186,
         n33187, n33188, n33189, n33190, n33191, n33192, n33193, n33194,
         n33195, n33196, n33197, n33198, n33199, n33200, n33201, n33202,
         n33203, n33204, n33205, n33206, n33207, n33208, n33209, n33210,
         n33211, n33212, n33213, n33214, n33215, n33216, n33217, n33218,
         n33219, n33220, n33221, n33222, n33223, n33224, n33225, n33226,
         n33227, n33228, n33229, n33230, n33231, n33232, n33233, n33234,
         n33235, n33236, n33237, n33238, n33239, n33240, n33241, n33242,
         n33243, n33244, n33245, n33246, n33247, n33248, n33249, n33250,
         n33251, n33252, n33253, n33254, n33255, n33256, n33257, n33258,
         n33259, n33260, n33261, n33262, n33263, n33264, n33265, n33266,
         n33267, n33268, n33269, n33270, n33271, n33272, n33273, n33274,
         n33275, n33276, n33277, n33278, n33279, n33280, n33281, n33282,
         n33283, n33284, n33285, n33286, n33287, n33288, n33289, n33290,
         n33291, n33292, n33293, n33294, n33295, n33296, n33297, n33298,
         n33299, n33300, n33301, n33302, n33303, n33304, n33305, n33306,
         n33307, n33308, n33309, n33310, n33311, n33312, n33313, n33314,
         n33315, n33316, n33317, n33318, n33319, n33320, n33321, n33322,
         n33323, n33324, n33325, n33326, n33327, n33328, n33329, n33330,
         n33331, n33332, n33333, n33334, n33335, n33336, n33337, n33338,
         n33339, n33340, n33341, n33342, n33343, n33344, n33345, n33346,
         n33347, n33348, n33349, n33350, n33351, n33352, n33353, n33354,
         n33355, n33356, n33357, n33358, n33359, n33360, n33361, n33362,
         n33363, n33364, n33365, n33366, n33367, n33368, n33369, n33370,
         n33371, n33372, n33373, n33374, n33375, n33376, n33377, n33378,
         n33379, n33380, n33381, n33382, n33383, n33384, n33385, n33386,
         n33387, n33388, n33389, n33390, n33391, n33392, n33393, n33394,
         n33395, n33396, n33397, n33398, n33399, n33400, n33401, n33402,
         n33403, n33404, n33405, n33406, n33407, n33408, n33409, n33410,
         n33411, n33412, n33413, n33414, n33415, n33416, n33417, n33418,
         n33419, n33420, n33421, n33422, n33423, n33424, n33425, n33426,
         n33427, n33428, n33429, n33430, n33431, n33432, n33433, n33434,
         n33435, n33436, n33437, n33438, n33439, n33440, n33441, n33442,
         n33443, n33444, n33445, n33446, n33447, n33448, n33449, n33450,
         n33451, n33452, n33453, n33454, n33455, n33456, n33457, n33458,
         n33459, n33460, n33461, n33462, n33463, n33464, n33465, n33466,
         n33467, n33468, n33469, n33470, n33471, n33472, n33473, n33474,
         n33475, n33476, n33477, n33478, n33479, n33480, n33481, n33482,
         n33483, n33484, n33485, n33486, n33487, n33488, n33489, n33490,
         n33491, n33492, n33493, n33494, n33495, n33496, n33497, n33498,
         n33499, n33500, n33501, n33502, n33503, n33504, n33505, n33506,
         n33507, n33508, n33509, n33510, n33511, n33512, n33513, n33514,
         n33515, n33516, n33517, n33518, n33519, n33520, n33521, n33522,
         n33523, n33524, n33525, n33526, n33527, n33528, n33529, n33530,
         n33531, n33532, n33533, n33534, n33535, n33536, n33537, n33538,
         n33539, n33540, n33541, n33542, n33543, n33544, n33545, n33546,
         n33547, n33548, n33549, n33550, n33551, n33552, n33553, n33554,
         n33555, n33556, n33557, n33558, n33559, n33560, n33561, n33562,
         n33563, n33564, n33565, n33566, n33567, n33568, n33569, n33570,
         n33571, n33572, n33573, n33574, n33575, n33576, n33577, n33578,
         n33579, n33580, n33581, n33582, n33583, n33584, n33585, n33586,
         n33587, n33588, n33589, n33590, n33591, n33592, n33593, n33594,
         n33595, n33596, n33597, n33598, n33599, n33600, n33601, n33602,
         n33603, n33604, n33605, n33606, n33607, n33608, n33609, n33610,
         n33611, n33612, n33613, n33614, n33615, n33616, n33617, n33618,
         n33619, n33620, n33621, n33622, n33623, n33624, n33625, n33626,
         n33627, n33628, n33629, n33630, n33631, n33632, n33633, n33634,
         n33635, n33636, n33637, n33638, n33639, n33640, n33641, n33642,
         n33643, n33644, n33645, n33646, n33647, n33648, n33649, n33650,
         n33651, n33652, n33653, n33654, n33655, n33656, n33657, n33658,
         n33659, n33660, n33661, n33662, n33663, n33664, n33665, n33666,
         n33667, n33668, n33669, n33670, n33671, n33672, n33673, n33674,
         n33675, n33676, n33677, n33678, n33679, n33680, n33681, n33682,
         n33683, n33684, n33685, n33686, n33687, n33688, n33689, n33690,
         n33691, n33692, n33693, n33694, n33695, n33696, n33697, n33698,
         n33699, n33700, n33701, n33702, n33703, n33704, n33705, n33706,
         n33707, n33708, n33709, n33710, n33711, n33712, n33713, n33714,
         n33715, n33716, n33717, n33718, n33719, n33720, n33721, n33722,
         n33723, n33724, n33725, n33726, n33727, n33728, n33729, n33730,
         n33731, n33732, n33733, n33734, n33735, n33736, n33737, n33738,
         n33739, n33740, n33741, n33742, n33743, n33744, n33745, n33746,
         n33747, n33748, n33749, n33750, n33751, n33752, n33753, n33754,
         n33755, n33756, n33757, n33758, n33759, n33760, n33761, n33762,
         n33763, n33764, n33765, n33766, n33767, n33768, n33769, n33770,
         n33771, n33772, n33773, n33774, n33775, n33776, n33777, n33778,
         n33779, n33780, n33781, n33782, n33783, n33784, n33785, n33786,
         n33787, n33788, n33789, n33790, n33791, n33792, n33793, n33794,
         n33795, n33796, n33797, n33798, n33799, n33800, n33801, n33802,
         n33803, n33804, n33805, n33806, n33807, n33808, n33809, n33810,
         n33811, n33812, n33813, n33814, n33815, n33816, n33817, n33818,
         n33819, n33820, n33821, n33822, n33823, n33824, n33825, n33826,
         n33827, n33828, n33829, n33830, n33831, n33832, n33833, n33834,
         n33835, n33836, n33837, n33838, n33839, n33840, n33841, n33842,
         n33843, n33844, n33845, n33846, n33847, n33848, n33849, n33850,
         n33851, n33852, n33853, n33854, n33855, n33856, n33857, n33858,
         n33859, n33860, n33861, n33862, n33863, n33864, n33865, n33866,
         n33867, n33868, n33869, n33870, n33871, n33872, n33873, n33874,
         n33875, n33876, n33877, n33878, n33879, n33880, n33881, n33882,
         n33883, n33884, n33885, n33886, n33887, n33888, n33889, n33890,
         n33891, n33892, n33893, n33894, n33895, n33896, n33897, n33898,
         n33899, n33900, n33901, n33902, n33903, n33904, n33905, n33906,
         n33907, n33908, n33909, n33910, n33911, n33912, n33913, n33914,
         n33915, n33916, n33917, n33918, n33919, n33920, n33921, n33922,
         n33923, n33924, n33925, n33926, n33927, n33928, n33929, n33930,
         n33931, n33932, n33933, n33934, n33935, n33936, n33937, n33938,
         n33939, n33940, n33941, n33942, n33943, n33944, n33945, n33946,
         n33947, n33948, n33949, n33950, n33951, n33952, n33953, n33954,
         n33955, n33956, n33957, n33958, n33959, n33960, n33961, n33962,
         n33963, n33964, n33965, n33966, n33967, n33968, n33969, n33970,
         n33971, n33972, n33973, n33974, n33975, n33976, n33977, n33978,
         n33979, n33980, n33981, n33982, n33983, n33984, n33985, n33986,
         n33987, n33988, n33989, n33990, n33991, n33992, n33993, n33994,
         n33995, n33996, n33997, n33998, n33999, n34000, n34001, n34002,
         n34003, n34004, n34005, n34006, n34007, n34008, n34009, n34010,
         n34011, n34012, n34013, n34014, n34015, n34016, n34017, n34018,
         n34019, n34020, n34021, n34022, n34023, n34024, n34025, n34026,
         n34027, n34028, n34029, n34030, n34031, n34032, n34033, n34034,
         n34035, n34036, n34037, n34038, n34039, n34040, n34041, n34042,
         n34043, n34044, n34045, n34046, n34047, n34048, n34049, n34050,
         n34051, n34052, n34053, n34054, n34055, n34056, n34057, n34058,
         n34059, n34060, n34061, n34062, n34063, n34064, n34065, n34066,
         n34067, n34068, n34069, n34070, n34071, n34072, n34073, n34074,
         n34075, n34076, n34077, n34078, n34079, n34080, n34081, n34082,
         n34083, n34084, n34085, n34086, n34087, n34088, n34089, n34090,
         n34091, n34092, n34093, n34094, n34095, n34096, n34097, n34098,
         n34099, n34100, n34101, n34102, n34103, n34104, n34105, n34106,
         n34107, n34108, n34109, n34110, n34111, n34112, n34113, n34114,
         n34115, n34116, n34117, n34118, n34119, n34120, n34121, n34122,
         n34123, n34124, n34125, n34126, n34127, n34128, n34129, n34130,
         n34131, n34132, n34133, n34134, n34135, n34136, n34137, n34138,
         n34139, n34140, n34141, n34142, n34143, n34144, n34145, n34146,
         n34147, n34148, n34149, n34150, n34151, n34152, n34153, n34154,
         n34155, n34156, n34157, n34158, n34159, n34160, n34161, n34162,
         n34163, n34164, n34165, n34166, n34167, n34168, n34169, n34170,
         n34171, n34172, n34173, n34174, n34175, n34176, n34177, n34178,
         n34179, n34180, n34181, n34182, n34183, n34184, n34185, n34186,
         n34187, n34188, n34189, n34190, n34191, n34192, n34193, n34194,
         n34195, n34196, n34197, n34198, n34199, n34200, n34201, n34202,
         n34203, n34204, n34205, n34206, n34207, n34208, n34209, n34210,
         n34211, n34212, n34213, n34214, n34215, n34216, n34217, n34218,
         n34219, n34220, n34221, n34222, n34223, n34224, n34225, n34226,
         n34227, n34228, n34229, n34230, n34231, n34232, n34233, n34234,
         n34235, n34236, n34237, n34238, n34239, n34240, n34241, n34242,
         n34243, n34244, n34245, n34246, n34247, n34248, n34249, n34250,
         n34251, n34252, n34253, n34254, n34255, n34256, n34257, n34258,
         n34259, n34260, n34261, n34262, n34263, n34264, n34265, n34266,
         n34267, n34268, n34269, n34270, n34271, n34272, n34273, n34274,
         n34275, n34276, n34277, n34278, n34279, n34280, n34281, n34282,
         n34283, n34284, n34285, n34286, n34287, n34288, n34289, n34290,
         n34291, n34292, n34293, n34294, n34295, n34296, n34297, n34298,
         n34299, n34300, n34301, n34302, n34303, n34304, n34305, n34306,
         n34307, n34308, n34309, n34310, n34311, n34312, n34313, n34314,
         n34315, n34316, n34317, n34318, n34319, n34320, n34321, n34322,
         n34323, n34324, n34325, n34326, n34327, n34328, n34329, n34330,
         n34331, n34332, n34333, n34334, n34335, n34336, n34337, n34338,
         n34339, n34340, n34341, n34342, n34343, n34344, n34345, n34346,
         n34347, n34348, n34349, n34350, n34351, n34352, n34353, n34354,
         n34355, n34356, n34357, n34358, n34359, n34360, n34361, n34362,
         n34363, n34364, n34365, n34366, n34367, n34368, n34369, n34370,
         n34371, n34372, n34373, n34374, n34375, n34376, n34377, n34378,
         n34379, n34380, n34381, n34382, n34383, n34384, n34385, n34386,
         n34387, n34388, n34389, n34390, n34391, n34392, n34393, n34394,
         n34395, n34396, n34397, n34398, n34399, n34400, n34401, n34402,
         n34403, n34404, n34405, n34406, n34407, n34408, n34409, n34410,
         n34411, n34412, n34413, n34414, n34415, n34416, n34417, n34418,
         n34419, n34420, n34421, n34422, n34423, n34424, n34425, n34426,
         n34427, n34428, n34429, n34430, n34431, n34432, n34433, n34434,
         n34435, n34436, n34437, n34438, n34439, n34440, n34441, n34442,
         n34443, n34444, n34445, n34446, n34447, n34448, n34449, n34450,
         n34451, n34452, n34453, n34454, n34455, n34456, n34457, n34458,
         n34459, n34460, n34461, n34462, n34463, n34464, n34465, n34466,
         n34467, n34468, n34469, n34470, n34471, n34472, n34473, n34474,
         n34475, n34476, n34477, n34478, n34479, n34480, n34481, n34482,
         n34483, n34484, n34485, n34486, n34487, n34488, n34489, n34490,
         n34491, n34492, n34493, n34494, n34495, n34496, n34497, n34498,
         n34499, n34500, n34501, n34502, n34503, n34504, n34505, n34506,
         n34507, n34508, n34509, n34510, n34511, n34512, n34513, n34514,
         n34515, n34516, n34517, n34518, n34519, n34520, n34521, n34522,
         n34523, n34524, n34525, n34526, n34527, n34528, n34529, n34530,
         n34531, n34532, n34533, n34534, n34535, n34536, n34537, n34538,
         n34539, n34540, n34541, n34542, n34543, n34544, n34545, n34546,
         n34547, n34548, n34549, n34550, n34551, n34552, n34553, n34554,
         n34555, n34556, n34557, n34558, n34559, n34560, n34561, n34562,
         n34563, n34564, n34565, n34566, n34567, n34568, n34569, n34570,
         n34571, n34572, n34573, n34574, n34575, n34576, n34577, n34578,
         n34579, n34580, n34581, n34582, n34583, n34584, n34585, n34586,
         n34587, n34588, n34589, n34590, n34591, n34592, n34593, n34594,
         n34595, n34596, n34597, n34598, n34599, n34600, n34601, n34602,
         n34603, n34604, n34605, n34606, n34607, n34608, n34609, n34610,
         n34611, n34612, n34613, n34614, n34615, n34616, n34617, n34618,
         n34619, n34620, n34621, n34622, n34623, n34624, n34625, n34626,
         n34627, n34628, n34629, n34630, n34631, n34632, n34633, n34634,
         n34635, n34636, n34637, n34638, n34639, n34640, n34641, n34642,
         n34643, n34644, n34645, n34646, n34647, n34648, n34649, n34650,
         n34651, n34652, n34653, n34654, n34655, n34656, n34657, n34658,
         n34659, n34660, n34661, n34662, n34663, n34664, n34665, n34666,
         n34667, n34668, n34669, n34670, n34671, n34672, n34673, n34674,
         n34675, n34676, n34677, n34678, n34679, n34680, n34681, n34682,
         n34683, n34684, n34685, n34686, n34687, n34688, n34689, n34690,
         n34691, n34692, n34693, n34694, n34695, n34696, n34697, n34698,
         n34699, n34700, n34701, n34702, n34703, n34704, n34705, n34706,
         n34707, n34708, n34709, n34710, n34711, n34712, n34713, n34714,
         n34715, n34716, n34717, n34718, n34719, n34720, n34721, n34722,
         n34723, n34724, n34725, n34726, n34727, n34728, n34729, n34730,
         n34731, n34732, n34733, n34734, n34735, n34736, n34737, n34738,
         n34739, n34740, n34741, n34742, n34743, n34744, n34745, n34746,
         n34747, n34748, n34749, n34750, n34751, n34752, n34753, n34754,
         n34755, n34756, n34757, n34758, n34759, n34760, n34761, n34762,
         n34763, n34764, n34765, n34766, n34767, n34768, n34769, n34770,
         n34771, n34772, n34773, n34774, n34775, n34776, n34777, n34778,
         n34779, n34780, n34781, n34782, n34783, n34784, n34785, n34786,
         n34787, n34788, n34789, n34790, n34791, n34792, n34793, n34794,
         n34795, n34796, n34797, n34798, n34799, n34800, n34801, n34802,
         n34803, n34804, n34805, n34806, n34807, n34808, n34809, n34810,
         n34811, n34812, n34813, n34814, n34815, n34816, n34817, n34818,
         n34819, n34820, n34821, n34822, n34823, n34824, n34825, n34826,
         n34827, n34828, n34829, n34830, n34831, n34832, n34833, n34834,
         n34835, n34836, n34837, n34838, n34839, n34840, n34841, n34842,
         n34843, n34844, n34845, n34846, n34847, n34848, n34849, n34850,
         n34851, n34852, n34853, n34854, n34855, n34856, n34857, n34858,
         n34859, n34860, n34861, n34862, n34863, n34864, n34865, n34866,
         n34867, n34868, n34869, n34870, n34871, n34872, n34873, n34874,
         n34875, n34876, n34877, n34878, n34879, n34880, n34881, n34882,
         n34883, n34884, n34885, n34886, n34887, n34888, n34889, n34890,
         n34891, n34892, n34893, n34894, n34895, n34896, n34897, n34898,
         n34899, n34900, n34901, n34902, n34903, n34904, n34905, n34906,
         n34907, n34908, n34909, n34910, n34911, n34912, n34913, n34914,
         n34915, n34916, n34917, n34918, n34919, n34920, n34921, n34922,
         n34923, n34924, n34925, n34926, n34927, n34928, n34929, n34930,
         n34931, n34932, n34933, n34934, n34935, n34936, n34937, n34938,
         n34939, n34940, n34941, n34942, n34943, n34944, n34945, n34946,
         n34947, n34948, n34949, n34950, n34951, n34952, n34953, n34954,
         n34955, n34956, n34957, n34958, n34959, n34960, n34961, n34962,
         n34963, n34964, n34965, n34966, n34967, n34968, n34969, n34970,
         n34971, n34972, n34973, n34974, n34975, n34976, n34977, n34978,
         n34979, n34980, n34981, n34982, n34983, n34984, n34985, n34986,
         n34987, n34988, n34989, n34990, n34991, n34992, n34993, n34994,
         n34995, n34996, n34997, n34998, n34999, n35000, n35001, n35002,
         n35003, n35004, n35005, n35006, n35007, n35008, n35009, n35010,
         n35011, n35012, n35013, n35014, n35015, n35016, n35017, n35018,
         n35019, n35020, n35021, n35022, n35023, n35024, n35025, n35026,
         n35027, n35028, n35029, n35030, n35031, n35032, n35033, n35034,
         n35035, n35036, n35037, n35038, n35039, n35040, n35041, n35042,
         n35043, n35044, n35045, n35046, n35047, n35048, n35049, n35050,
         n35051, n35052, n35053, n35054, n35055, n35056, n35057, n35058,
         n35059, n35060, n35061, n35062, n35063, n35064, n35065, n35066,
         n35067, n35068, n35069, n35070, n35071, n35072, n35073, n35074,
         n35075, n35076, n35077, n35078, n35079, n35080, n35081, n35082,
         n35083, n35084, n35085, n35086, n35087, n35088, n35089, n35090,
         n35091, n35092, n35093, n35094, n35095, n35096, n35097, n35098,
         n35099, n35100, n35101, n35102, n35103, n35104, n35105, n35106,
         n35107, n35108, n35109, n35110, n35111, n35112, n35113, n35114,
         n35115, n35116, n35117, n35118, n35119, n35120, n35121, n35122,
         n35123, n35124, n35125, n35126, n35127, n35128, n35129, n35130,
         n35131, n35132, n35133, n35134, n35135, n35136, n35137, n35138,
         n35139, n35140, n35141, n35142, n35143, n35144, n35145, n35146,
         n35147, n35148, n35149, n35150, n35151, n35152, n35153, n35154,
         n35155, n35156, n35157, n35158, n35159, n35160, n35161, n35162,
         n35163, n35164, n35165, n35166, n35167, n35168, n35169, n35170,
         n35171, n35172, n35173, n35174, n35175, n35176, n35177, n35178,
         n35179, n35180, n35181, n35182, n35183, n35184, n35185, n35186,
         n35187, n35188, n35189, n35190, n35191, n35192, n35193, n35194,
         n35195, n35196, n35197, n35198, n35199, n35200, n35201, n35202,
         n35203, n35204, n35205, n35206, n35207, n35208, n35209, n35210,
         n35211, n35212, n35213, n35214, n35215, n35216, n35217, n35218,
         n35219, n35220, n35221, n35222, n35223, n35224, n35225, n35226,
         n35227, n35228, n35229, n35230, n35231, n35232, n35233, n35234,
         n35235, n35236, n35237, n35238, n35239, n35240, n35241, n35242,
         n35243, n35244, n35245, n35246, n35247, n35248, n35249, n35250,
         n35251, n35252, n35253, n35254, n35255, n35256, n35257, n35258,
         n35259, n35260, n35261, n35262, n35263, n35264, n35265, n35266,
         n35267, n35268, n35269, n35270, n35271, n35272, n35273, n35274,
         n35275, n35276, n35277, n35278, n35279, n35280, n35281, n35282,
         n35283, n35284, n35285, n35286, n35287, n35288, n35289, n35290,
         n35291, n35292, n35293, n35294, n35295, n35296, n35297, n35298,
         n35299, n35300, n35301, n35302, n35303, n35304, n35305, n35306,
         n35307, n35308, n35309, n35310, n35311, n35312, n35313, n35314,
         n35315, n35316, n35317, n35318, n35319, n35320, n35321, n35322,
         n35323, n35324, n35325, n35326, n35327, n35328, n35329, n35330,
         n35331, n35332, n35333, n35334, n35335, n35336, n35337, n35338,
         n35339, n35340, n35341, n35342, n35343, n35344, n35345, n35346,
         n35347, n35348, n35349, n35350, n35351, n35352, n35353, n35354,
         n35355, n35356, n35357, n35358, n35359, n35360, n35361, n35362,
         n35363, n35364, n35365, n35366, n35367, n35368, n35369, n35370,
         n35371, n35372, n35373, n35374, n35375, n35376, n35377, n35378,
         n35379, n35380, n35381, n35382, n35383, n35384, n35385, n35386,
         n35387, n35388, n35389, n35390, n35391, n35392, n35393, n35394,
         n35395, n35396, n35397, n35398, n35399, n35400, n35401, n35402,
         n35403, n35404, n35405, n35406, n35407, n35408, n35409, n35410,
         n35411, n35412, n35413, n35414, n35415, n35416, n35417, n35418,
         n35419, n35420, n35421, n35422, n35423, n35424, n35425, n35426,
         n35427, n35428, n35429, n35430, n35431, n35432, n35433, n35434,
         n35435, n35436, n35437, n35438, n35439, n35440, n35441, n35442,
         n35443, n35444, n35445, n35446, n35447, n35448, n35449, n35450,
         n35451, n35452, n35453, n35454, n35455, n35456, n35457, n35458,
         n35459, n35460, n35461, n35462, n35463, n35464, n35465, n35466,
         n35467, n35468, n35469, n35470, n35471, n35472, n35473, n35474,
         n35475, n35476, n35477, n35478, n35479, n35480, n35481, n35482,
         n35483, n35484, n35485, n35486, n35487, n35488, n35489, n35490,
         n35491, n35492, n35493, n35494, n35495, n35496, n35497, n35498,
         n35499, n35500, n35501, n35502, n35503, n35504, n35505, n35506,
         n35507, n35508, n35509, n35510, n35511, n35512, n35513, n35514,
         n35515, n35516, n35517, n35518, n35519, n35520, n35521, n35522,
         n35523, n35524, n35525, n35526, n35527, n35528, n35529, n35530,
         n35531, n35532, n35533, n35534, n35535, n35536, n35537, n35538,
         n35539, n35540, n35541, n35542, n35543, n35544, n35545, n35546,
         n35547, n35548, n35549, n35550, n35551, n35552, n35553, n35554,
         n35555, n35556, n35557, n35558, n35559, n35560, n35561, n35562,
         n35563, n35564, n35565, n35566, n35567, n35568, n35569, n35570,
         n35571, n35572, n35573, n35574, n35575, n35576, n35577, n35578,
         n35579, n35580, n35581, n35582, n35583, n35584, n35585, n35586,
         n35587, n35588, n35589, n35590, n35591, n35592, n35593, n35594,
         n35595, n35596, n35597, n35598, n35599, n35600, n35601, n35602,
         n35603, n35604, n35605, n35606, n35607, n35608, n35609, n35610,
         n35611, n35612, n35613, n35614, n35615, n35616, n35617, n35618,
         n35619, n35620, n35621, n35622, n35623, n35624, n35625, n35626,
         n35627, n35628, n35629, n35630, n35631, n35632, n35633, n35634,
         n35635, n35636, n35637, n35638, n35639, n35640, n35641, n35642,
         n35643, n35644, n35645, n35646, n35647, n35648, n35649, n35650,
         n35651, n35652, n35653, n35654, n35655, n35656, n35657, n35658,
         n35659, n35660, n35661, n35662, n35663, n35664, n35665, n35666,
         n35667, n35668, n35669, n35670, n35671, n35672, n35673, n35674,
         n35675, n35676, n35677, n35678, n35679, n35680, n35681, n35682,
         n35683, n35684, n35685, n35686, n35687, n35688, n35689, n35690,
         n35691, n35692, n35693, n35694, n35695, n35696, n35697, n35698,
         n35699, n35700, n35701, n35702, n35703, n35704, n35705, n35706,
         n35707, n35708, n35709, n35710, n35711, n35712, n35713, n35714,
         n35715, n35716, n35717, n35718, n35719, n35720, n35721, n35722,
         n35723, n35724, n35725, n35726, n35727, n35728, n35729, n35730,
         n35731, n35732, n35733, n35734, n35735, n35736, n35737, n35738,
         n35739, n35740, n35741, n35742, n35743, n35744, n35745, n35746,
         n35747, n35748, n35749, n35750, n35751, n35752, n35753, n35754,
         n35755, n35756, n35757, n35758, n35759, n35760, n35761, n35762,
         n35763, n35764, n35765, n35766, n35767, n35768, n35769, n35770,
         n35771, n35772, n35773, n35774, n35775, n35776, n35777, n35778,
         n35779, n35780, n35781, n35782, n35783, n35784, n35785, n35786,
         n35787, n35788, n35789, n35790, n35791, n35792, n35793, n35794,
         n35795, n35796, n35797, n35798, n35799, n35800, n35801, n35802,
         n35803, n35804, n35805, n35806, n35807, n35808, n35809, n35810,
         n35811, n35812, n35813, n35814, n35815, n35816, n35817, n35818,
         n35819, n35820, n35821, n35822, n35823, n35824, n35825, n35826,
         n35827, n35828, n35829, n35830, n35831, n35832, n35833, n35834,
         n35835, n35836, n35837, n35838, n35839, n35840, n35841, n35842,
         n35843, n35844, n35845, n35846, n35847, n35848, n35849, n35850,
         n35851, n35852, n35853, n35854, n35855, n35856, n35857, n35858,
         n35859, n35860, n35861, n35862, n35863, n35864, n35865, n35866,
         n35867, n35868, n35869, n35870, n35871, n35872, n35873, n35874,
         n35875, n35876, n35877, n35878, n35879, n35880, n35881, n35882,
         n35883, n35884, n35885, n35886, n35887, n35888, n35889, n35890,
         n35891, n35892, n35893, n35894, n35895, n35896, n35897, n35898,
         n35899, n35900, n35901, n35902, n35903, n35904, n35905, n35906,
         n35907, n35908, n35909, n35910, n35911, n35912, n35913, n35914,
         n35915, n35916, n35917, n35918, n35919, n35920, n35921, n35922,
         n35923, n35924, n35925, n35926, n35927, n35928, n35929, n35930,
         n35931, n35932, n35933, n35934, n35935, n35936, n35937, n35938,
         n35939, n35940, n35941, n35942, n35943, n35944, n35945, n35946,
         n35947, n35948, n35949, n35950, n35951, n35952, n35953, n35954,
         n35955, n35956, n35957, n35958, n35959, n35960, n35961, n35962,
         n35963, n35964, n35965, n35966, n35967, n35968, n35969, n35970,
         n35971, n35972, n35973, n35974, n35975, n35976, n35977, n35978,
         n35979, n35980, n35981, n35982, n35983, n35984, n35985, n35986,
         n35987, n35988, n35989, n35990, n35991, n35992, n35993, n35994,
         n35995, n35996, n35997, n35998, n35999, n36000, n36001, n36002,
         n36003, n36004, n36005, n36006, n36007, n36008, n36009, n36010,
         n36011, n36012, n36013, n36014, n36015, n36016, n36017, n36018,
         n36019, n36020, n36021, n36022, n36023, n36024, n36025, n36026,
         n36027, n36028, n36029, n36030, n36031, n36032, n36033, n36034,
         n36035, n36036, n36037, n36038, n36039, n36040, n36041, n36042,
         n36043, n36044, n36045, n36046, n36047, n36048, n36049, n36050,
         n36051, n36052, n36053, n36054, n36055, n36056, n36057, n36058,
         n36059, n36060, n36061, n36062, n36063, n36064, n36065, n36066,
         n36067, n36068, n36069, n36070, n36071, n36072, n36073, n36074,
         n36075, n36076, n36077, n36078, n36079, n36080, n36081, n36082,
         n36083, n36084, n36085, n36086, n36087, n36088, n36089, n36090,
         n36091, n36092, n36093, n36094, n36095, n36096, n36097, n36098,
         n36099, n36100, n36101, n36102, n36103, n36104, n36105, n36106,
         n36107, n36108, n36109, n36110, n36111, n36112, n36113, n36114,
         n36115, n36116, n36117, n36118, n36119, n36120, n36121, n36122,
         n36123, n36124, n36125, n36126, n36127, n36128, n36129, n36130,
         n36131, n36132, n36133, n36134, n36135, n36136, n36137, n36138,
         n36139, n36140, n36141, n36142, n36143, n36144, n36145, n36146,
         n36147, n36148, n36149, n36150, n36151, n36152, n36153, n36154,
         n36155, n36156, n36157, n36158, n36159, n36160, n36161, n36162,
         n36163, n36164, n36165, n36166, n36167, n36168, n36169, n36170,
         n36171, n36172, n36173, n36174, n36175, n36176, n36177, n36178,
         n36179, n36180, n36181, n36182, n36183, n36184, n36185, n36186,
         n36187, n36188, n36189, n36190, n36191, n36192, n36193, n36194,
         n36195, n36196, n36197, n36198, n36199, n36200, n36201, n36202,
         n36203, n36204, n36205, n36206, n36207, n36208, n36209, n36210,
         n36211, n36212, n36213, n36214, n36215, n36216, n36217, n36218,
         n36219, n36220, n36221, n36222, n36223, n36224, n36225, n36226,
         n36227, n36228, n36229, n36230, n36231, n36232, n36233, n36234,
         n36235, n36236, n36237, n36238, n36239, n36240, n36241, n36242,
         n36243, n36244, n36245, n36246, n36247, n36248, n36249, n36250,
         n36251, n36252, n36253, n36254, n36255, n36256, n36257, n36258,
         n36259, n36260, n36261, n36262, n36263, n36264, n36265, n36266,
         n36267, n36268, n36269, n36270, n36271, n36272, n36273, n36274,
         n36275, n36276, n36277, n36278, n36279, n36280, n36281, n36282,
         n36283, n36284, n36285, n36286, n36287, n36288, n36289, n36290,
         n36291, n36292, n36293, n36294, n36295, n36296, n36297, n36298,
         n36299, n36300, n36301, n36302, n36303, n36304, n36305, n36306,
         n36307, n36308, n36309, n36310, n36311, n36312, n36313, n36314,
         n36315, n36316, n36317, n36318, n36319, n36320, n36321, n36322,
         n36323, n36324, n36325, n36326, n36327, n36328, n36329, n36330,
         n36331, n36332, n36333, n36334, n36335, n36336, n36337, n36338,
         n36339, n36340, n36341, n36342, n36343, n36344, n36345, n36346,
         n36347, n36348, n36349, n36350, n36351, n36352, n36353, n36354,
         n36355, n36356, n36357, n36358, n36359, n36360, n36361, n36362,
         n36363, n36364, n36365, n36366, n36367, n36368, n36369, n36370,
         n36371, n36372, n36373, n36374, n36375, n36376, n36377, n36378,
         n36379, n36380, n36381, n36382, n36383, n36384, n36385, n36386,
         n36387, n36388, n36389, n36390, n36391, n36392, n36393, n36394,
         n36395, n36396, n36397, n36398, n36399, n36400, n36401, n36402,
         n36403, n36404, n36405, n36406, n36407, n36408, n36409, n36410,
         n36411, n36412, n36413, n36414, n36415, n36416, n36417, n36418,
         n36419, n36420, n36421, n36422, n36423, n36424, n36425, n36426,
         n36427, n36428, n36429, n36430, n36431, n36432, n36433, n36434,
         n36435, n36436, n36437, n36438, n36439, n36440, n36441, n36442,
         n36443, n36444, n36445, n36446, n36447, n36448, n36449, n36450,
         n36451, n36452, n36453, n36454, n36455, n36456, n36457, n36458,
         n36459, n36460, n36461, n36462, n36463, n36464, n36465, n36466,
         n36467, n36468, n36469, n36470, n36471, n36472, n36473, n36474,
         n36475, n36476, n36477, n36478, n36479, n36480, n36481, n36482,
         n36483, n36484, n36485, n36486, n36487, n36488, n36489, n36490,
         n36491, n36492, n36493, n36494, n36495, n36496, n36497, n36498,
         n36499, n36500, n36501, n36502, n36503, n36504, n36505, n36506,
         n36507, n36508, n36509, n36510, n36511, n36512, n36513, n36514,
         n36515, n36516, n36517, n36518, n36519, n36520, n36521, n36522,
         n36523, n36524, n36525, n36526, n36527, n36528, n36529, n36530,
         n36531, n36532, n36533, n36534, n36535, n36536, n36537, n36538,
         n36539, n36540, n36541, n36542, n36543, n36544, n36545, n36546,
         n36547, n36548, n36549, n36550, n36551, n36552, n36553, n36554,
         n36555, n36556, n36557, n36558, n36559, n36560, n36561, n36562,
         n36563, n36564, n36565, n36566, n36567, n36568, n36569, n36570,
         n36571, n36572, n36573, n36574, n36575, n36576, n36577, n36578,
         n36579, n36580, n36581, n36582, n36583, n36584, n36585, n36586,
         n36587, n36588, n36589, n36590, n36591, n36592, n36593, n36594,
         n36595, n36596, n36597, n36598, n36599, n36600, n36601, n36602,
         n36603, n36604, n36605, n36606, n36607, n36608, n36609, n36610,
         n36611, n36612, n36613, n36614, n36615, n36616, n36617, n36618,
         n36619, n36620, n36621, n36622, n36623, n36624, n36625, n36626,
         n36627, n36628, n36629, n36630, n36631, n36632, n36633, n36634,
         n36635, n36636, n36637, n36638, n36639, n36640, n36641, n36642,
         n36643, n36644, n36645, n36646, n36647, n36648, n36649, n36650,
         n36651, n36652, n36653, n36654, n36655, n36656, n36657, n36658,
         n36659, n36660, n36661, n36662, n36663, n36664, n36665, n36666,
         n36667, n36668, n36669, n36670, n36671, n36672, n36673, n36674,
         n36675, n36676, n36677, n36678, n36679, n36680, n36681, n36682,
         n36683, n36684, n36685, n36686, n36687, n36688, n36689, n36690,
         n36691, n36692, n36693, n36694, n36695, n36696, n36697, n36698,
         n36699, n36700, n36701, n36702, n36703, n36704, n36705, n36706,
         n36707, n36708, n36709, n36710, n36711, n36712, n36713, n36714,
         n36715, n36716, n36717, n36718, n36719, n36720, n36721, n36722,
         n36723, n36724, n36725, n36726, n36727, n36728, n36729, n36730,
         n36731, n36732, n36733, n36734, n36735, n36736, n36737, n36738,
         n36739, n36740, n36741, n36742, n36743, n36744, n36745, n36746,
         n36747, n36748, n36749, n36750, n36751, n36752, n36753, n36754,
         n36755, n36756, n36757, n36758, n36759, n36760, n36761, n36762,
         n36763, n36764, n36765, n36766, n36767, n36768, n36769, n36770,
         n36771, n36772, n36773, n36774, n36775, n36776, n36777, n36778,
         n36779, n36780, n36781, n36782, n36783, n36784, n36785, n36786,
         n36787, n36788, n36789, n36790, n36791, n36792, n36793, n36794,
         n36795, n36796, n36797, n36798, n36799, n36800, n36801, n36802,
         n36803, n36804, n36805, n36806, n36807, n36808, n36809, n36810,
         n36811, n36812, n36813, n36814, n36815, n36816, n36817, n36818,
         n36819, n36820, n36821, n36822, n36823, n36824, n36825, n36826,
         n36827, n36828, n36829, n36830, n36831, n36832, n36833, n36834,
         n36835, n36836, n36837, n36838, n36839, n36840, n36841, n36842,
         n36843, n36844, n36845, n36846, n36847, n36848, n36849, n36850,
         n36851, n36852, n36853, n36854, n36855, n36856, n36857, n36858,
         n36859, n36860, n36861, n36862, n36863, n36864, n36865, n36866,
         n36867, n36868, n36869, n36870, n36871, n36872, n36873, n36874,
         n36875, n36876, n36877, n36878, n36879, n36880, n36881, n36882,
         n36883, n36884, n36885, n36886, n36887, n36888, n36889, n36890,
         n36891, n36892, n36893, n36894, n36895, n36896, n36897, n36898,
         n36899, n36900, n36901, n36902, n36903, n36904, n36905, n36906,
         n36907, n36908, n36909, n36910, n36911, n36912, n36913, n36914,
         n36915, n36916, n36917, n36918, n36919, n36920, n36921, n36922,
         n36923, n36924, n36925, n36926, n36927, n36928, n36929, n36930,
         n36931, n36932, n36933, n36934, n36935, n36936, n36937, n36938,
         n36939, n36940, n36941, n36942, n36943, n36944, n36945, n36946,
         n36947, n36948, n36949, n36950, n36951, n36952, n36953, n36954,
         n36955, n36956, n36957, n36958, n36959, n36960, n36961, n36962,
         n36963, n36964, n36965, n36966, n36967, n36968, n36969, n36970,
         n36971, n36972, n36973, n36974, n36975, n36976, n36977, n36978,
         n36979, n36980, n36981, n36982, n36983, n36984, n36985, n36986,
         n36987, n36988, n36989, n36990, n36991, n36992, n36993, n36994,
         n36995, n36996, n36997, n36998, n36999, n37000, n37001, n37002,
         n37003, n37004, n37005, n37006, n37007, n37008, n37009, n37010,
         n37011, n37012, n37013, n37014, n37015, n37016, n37017, n37018,
         n37019, n37020, n37021, n37022, n37023, n37024, n37025, n37026,
         n37027, n37028, n37029, n37030, n37031, n37032, n37033, n37034,
         n37035, n37036, n37037, n37038, n37039, n37040, n37041, n37042,
         n37043, n37044, n37045, n37046, n37047, n37048, n37049, n37050,
         n37051, n37052, n37053, n37054, n37055, n37056, n37057, n37058,
         n37059, n37060, n37061, n37062, n37063, n37064, n37065, n37066,
         n37067, n37068, n37069, n37070, n37071, n37072, n37073, n37074,
         n37075, n37076, n37077, n37078, n37079, n37080, n37081, n37082,
         n37083, n37084, n37085, n37086, n37087, n37088, n37089, n37090,
         n37091, n37092, n37093, n37094, n37095, n37096, n37097, n37098,
         n37099, n37100, n37101, n37102, n37103, n37104, n37105, n37106,
         n37107, n37108, n37109, n37110, n37111, n37112, n37113, n37114,
         n37115, n37116, n37117, n37118, n37119, n37120, n37121, n37122,
         n37123, n37124, n37125, n37126, n37127, n37128, n37129, n37130,
         n37131, n37132, n37133, n37134, n37135, n37136, n37137, n37138,
         n37139, n37140, n37141, n37142, n37143, n37144, n37145, n37146,
         n37147, n37148, n37149, n37150, n37151, n37152, n37153, n37154,
         n37155, n37156, n37157, n37158, n37159, n37160, n37161, n37162,
         n37163, n37164, n37165, n37166, n37167, n37168, n37169, n37170,
         n37171, n37172, n37173, n37174, n37175, n37176, n37177, n37178,
         n37179, n37180, n37181, n37182, n37183, n37184, n37185, n37186,
         n37187, n37188, n37189, n37190, n37191, n37192, n37193, n37194,
         n37195, n37196, n37197, n37198, n37199, n37200, n37201, n37202,
         n37203, n37204, n37205, n37206, n37207, n37208, n37209, n37210,
         n37211, n37212, n37213, n37214, n37215, n37216, n37217, n37218,
         n37219, n37220, n37221, n37222, n37223, n37224, n37225, n37226,
         n37227, n37228, n37229, n37230, n37231, n37232, n37233, n37234,
         n37235, n37236, n37237, n37238, n37239, n37240, n37241, n37242,
         n37243, n37244, n37245, n37246, n37247, n37248, n37249, n37250,
         n37251, n37252, n37253, n37254, n37255, n37256, n37257, n37258,
         n37259, n37260, n37261, n37262, n37263, n37264, n37265, n37266,
         n37267, n37268, n37269, n37270, n37271, n37272, n37273, n37274,
         n37275, n37276, n37277, n37278, n37279, n37280, n37281, n37282,
         n37283, n37284, n37285, n37286, n37287, n37288, n37289, n37290,
         n37291, n37292, n37293, n37294, n37295, n37296, n37297, n37298,
         n37299, n37300, n37301, n37302, n37303, n37304, n37305, n37306,
         n37307, n37308, n37309, n37310, n37311, n37312, n37313, n37314,
         n37315, n37316, n37317, n37318, n37319, n37320, n37321, n37322,
         n37323, n37324, n37325, n37326, n37327, n37328, n37329, n37330,
         n37331, n37332, n37333, n37334, n37335, n37336, n37337, n37338,
         n37339, n37340, n37341, n37342, n37343, n37344, n37345, n37346,
         n37347, n37348, n37349, n37350, n37351, n37352, n37353, n37354,
         n37355, n37356, n37357, n37358, n37359, n37360, n37361, n37362,
         n37363, n37364, n37365, n37366, n37367, n37368, n37369, n37370,
         n37371, n37372, n37373, n37374, n37375, n37376, n37377, n37378,
         n37379, n37380, n37381, n37382, n37383, n37384, n37385, n37386,
         n37387, n37388, n37389, n37390, n37391, n37392, n37393, n37394,
         n37395, n37396, n37397, n37398, n37399, n37400, n37401, n37402,
         n37403, n37404, n37405, n37406, n37407, n37408, n37409, n37410,
         n37411, n37412, n37413, n37414, n37415, n37416, n37417, n37418,
         n37419, n37420, n37421, n37422, n37423, n37424, n37425, n37426,
         n37427, n37428, n37429, n37430, n37431, n37432, n37433, n37434,
         n37435, n37436, n37437, n37438, n37439, n37440, n37441, n37442,
         n37443, n37444, n37445, n37446, n37447, n37448, n37449, n37450,
         n37451, n37452, n37453, n37454, n37455, n37456, n37457, n37458,
         n37459, n37460, n37461, n37462, n37463, n37464, n37465, n37466,
         n37467, n37468, n37469, n37470, n37471, n37472, n37473, n37474,
         n37475, n37476, n37477, n37478, n37479, n37480, n37481, n37482,
         n37483, n37484, n37485, n37486, n37487, n37488, n37489, n37490,
         n37491, n37492, n37493, n37494, n37495, n37496, n37497, n37498,
         n37499, n37500, n37501, n37502, n37503, n37504, n37505, n37506,
         n37507, n37508, n37509, n37510, n37511, n37512, n37513, n37514,
         n37515, n37516, n37517, n37518, n37519, n37520, n37521, n37522,
         n37523, n37524, n37525, n37526, n37527, n37528, n37529, n37530,
         n37531, n37532, n37533, n37534, n37535, n37536, n37537, n37538,
         n37539, n37540, n37541, n37542, n37543, n37544, n37545, n37546,
         n37547, n37548, n37549, n37550, n37551, n37552, n37553, n37554,
         n37555, n37556, n37557, n37558, n37559, n37560, n37561, n37562,
         n37563, n37564, n37565, n37566, n37567, n37568, n37569, n37570,
         n37571, n37572, n37573, n37574, n37575, n37576, n37577, n37578,
         n37579, n37580, n37581, n37582, n37583, n37584, n37585, n37586,
         n37587, n37588, n37589, n37590, n37591, n37592, n37593, n37594,
         n37595, n37596, n37597, n37598, n37599, n37600, n37601, n37602,
         n37603, n37604, n37605, n37606, n37607, n37608, n37609, n37610,
         n37611, n37612, n37613, n37614, n37615, n37616, n37617, n37618,
         n37619, n37620, n37621, n37622, n37623, n37624, n37625, n37626,
         n37627, n37628, n37629, n37630, n37631, n37632, n37633, n37634,
         n37635, n37636, n37637, n37638, n37639, n37640, n37641, n37642,
         n37643, n37644, n37645, n37646, n37647, n37648, n37649, n37650,
         n37651, n37652, n37653, n37654, n37655, n37656, n37657, n37658,
         n37659, n37660, n37661, n37662, n37663, n37664, n37665, n37666,
         n37667, n37668, n37669, n37670, n37671, n37672, n37673, n37674,
         n37675, n37676, n37677, n37678, n37679, n37680, n37681, n37682,
         n37683, n37684, n37685, n37686, n37687, n37688, n37689, n37690,
         n37691, n37692, n37693, n37694, n37695, n37696, n37697, n37698,
         n37699, n37700, n37701, n37702, n37703, n37704, n37705, n37706,
         n37707, n37708, n37709, n37710, n37711, n37712, n37713, n37714,
         n37715, n37716, n37717, n37718, n37719, n37720, n37721, n37722,
         n37723, n37724, n37725, n37726, n37727, n37728, n37729, n37730,
         n37731, n37732, n37733, n37734, n37735, n37736, n37737, n37738,
         n37739, n37740, n37741, n37742, n37743, n37744, n37745, n37746,
         n37747, n37748, n37749, n37750, n37751, n37752, n37753, n37754,
         n37755, n37756, n37757, n37758, n37759, n37760, n37761, n37762,
         n37763, n37764, n37765, n37766, n37767, n37768, n37769, n37770,
         n37771, n37772, n37773, n37774, n37775, n37776, n37777, n37778,
         n37779, n37780, n37781, n37782, n37783, n37784, n37785, n37786,
         n37787, n37788, n37789, n37790, n37791, n37792, n37793, n37794,
         n37795, n37796, n37797, n37798, n37799, n37800, n37801, n37802,
         n37803, n37804, n37805, n37806, n37807, n37808, n37809, n37810,
         n37811, n37812, n37813, n37814, n37815, n37816, n37817, n37818,
         n37819, n37820, n37821, n37822, n37823, n37824, n37825, n37826,
         n37827, n37828, n37829, n37830, n37831, n37832, n37833, n37834,
         n37835, n37836, n37837, n37838, n37839, n37840, n37841, n37842,
         n37843, n37844, n37845, n37846, n37847, n37848, n37849, n37850,
         n37851, n37852, n37853, n37854, n37855, n37856, n37857, n37858,
         n37859, n37860, n37861, n37862, n37863, n37864, n37865, n37866,
         n37867, n37868, n37869, n37870, n37871, n37872, n37873, n37874,
         n37875, n37876, n37877, n37878, n37879, n37880, n37881, n37882,
         n37883, n37884, n37885, n37886, n37887, n37888, n37889, n37890,
         n37891, n37892, n37893, n37894, n37895, n37896, n37897, n37898,
         n37899, n37900, n37901, n37902, n37903, n37904, n37905, n37906,
         n37907, n37908, n37909, n37910, n37911, n37912, n37913, n37914,
         n37915, n37916, n37917, n37918, n37919, n37920, n37921, n37922,
         n37923, n37924, n37925, n37926, n37927, n37928, n37929, n37930,
         n37931, n37932, n37933, n37934, n37935, n37936, n37937, n37938,
         n37939, n37940, n37941, n37942, n37943, n37944, n37945, n37946,
         n37947, n37948, n37949, n37950, n37951, n37952, n37953, n37954,
         n37955, n37956, n37957, n37958, n37959, n37960, n37961, n37962,
         n37963, n37964, n37965, n37966, n37967, n37968, n37969, n37970,
         n37971, n37972, n37973, n37974, n37975, n37976, n37977, n37978,
         n37979, n37980, n37981, n37982, n37983, n37984, n37985, n37986,
         n37987, n37988, n37989, n37990, n37991, n37992, n37993, n37994,
         n37995, n37996, n37997, n37998, n37999, n38000, n38001, n38002,
         n38003, n38004, n38005, n38006, n38007, n38008, n38009, n38010,
         n38011, n38012, n38013, n38014, n38015, n38016, n38017, n38018,
         n38019, n38020, n38021, n38022, n38023, n38024, n38025, n38026,
         n38027, n38028, n38029, n38030, n38031, n38032, n38033, n38034,
         n38035, n38036, n38037, n38038, n38039, n38040, n38041, n38042,
         n38043, n38044, n38045, n38046, n38047, n38048, n38049, n38050,
         n38051, n38052, n38053, n38054, n38055, n38056, n38057, n38058,
         n38059, n38060, n38061, n38062, n38063, n38064, n38065, n38066,
         n38067, n38068, n38069, n38070, n38071, n38072, n38073, n38074,
         n38075, n38076, n38077, n38078, n38079, n38080, n38081, n38082,
         n38083, n38084, n38085, n38086, n38087, n38088, n38089, n38090,
         n38091, n38092, n38093, n38094, n38095, n38096, n38097, n38098,
         n38099, n38100, n38101, n38102, n38103, n38104, n38105, n38106,
         n38107, n38108, n38109, n38110, n38111, n38112, n38113, n38114,
         n38115, n38116, n38117, n38118, n38119, n38120, n38121, n38122,
         n38123, n38124, n38125, n38126, n38127, n38128, n38129, n38130,
         n38131, n38132, n38133, n38134, n38135, n38136, n38137, n38138,
         n38139, n38140, n38141, n38142, n38143, n38144, n38145, n38146,
         n38147, n38148, n38149, n38150, n38151, n38152, n38153, n38154,
         n38155, n38156, n38157, n38158, n38159, n38160, n38161, n38162,
         n38163, n38164, n38165, n38166, n38167, n38168, n38169, n38170,
         n38171, n38172, n38173, n38174, n38175, n38176, n38177, n38178,
         n38179, n38180, n38181, n38182, n38183, n38184, n38185, n38186,
         n38187, n38188, n38189, n38190, n38191, n38192, n38193, n38194,
         n38195, n38196, n38197, n38198, n38199, n38200, n38201, n38202,
         n38203, n38204, n38205, n38206, n38207, n38208, n38209, n38210,
         n38211, n38212, n38213, n38214, n38215, n38216, n38217, n38218,
         n38219, n38220, n38221, n38222, n38223, n38224, n38225, n38226,
         n38227, n38228, n38229, n38230, n38231, n38232, n38233, n38234,
         n38235, n38236, n38237, n38238, n38239, n38240, n38241, n38242,
         n38243, n38244, n38245, n38246, n38247, n38248, n38249, n38250,
         n38251, n38252, n38253, n38254, n38255, n38256, n38257, n38258,
         n38259, n38260, n38261, n38262, n38263, n38264, n38265, n38266,
         n38267, n38268, n38269, n38270, n38271, n38272, n38273, n38274,
         n38275, n38276, n38277, n38278, n38279, n38280, n38281, n38282,
         n38283, n38284, n38285, n38286, n38287, n38288, n38289, n38290,
         n38291, n38292, n38293, n38294, n38295, n38296, n38297, n38298,
         n38299, n38300, n38301, n38302, n38303, n38304, n38305, n38306,
         n38307, n38308, n38309, n38310, n38311, n38312, n38313, n38314,
         n38315, n38316, n38317, n38318, n38319, n38320, n38321, n38322,
         n38323, n38324, n38325, n38326, n38327, n38328, n38329, n38330,
         n38331, n38332, n38333, n38334, n38335, n38336, n38337, n38338,
         n38339, n38340, n38341, n38342, n38343, n38344, n38345, n38346,
         n38347, n38348, n38349, n38350, n38351, n38352, n38353, n38354,
         n38355, n38356, n38357, n38358, n38359, n38360, n38361, n38362,
         n38363, n38364, n38365, n38366, n38367, n38368, n38369, n38370,
         n38371, n38372, n38373, n38374, n38375, n38376, n38377, n38378,
         n38379, n38380, n38381, n38382, n38383, n38384, n38385, n38386,
         n38387, n38388, n38389, n38390, n38391, n38392, n38393, n38394,
         n38395, n38396, n38397, n38398, n38399, n38400, n38401, n38402,
         n38403, n38404, n38405, n38406, n38407, n38408, n38409, n38410,
         n38411, n38412, n38413, n38414, n38415, n38416, n38417, n38418,
         n38419, n38420, n38421, n38422, n38423, n38424, n38425, n38426,
         n38427, n38428, n38429, n38430, n38431, n38432, n38433, n38434,
         n38435, n38436, n38437, n38438, n38439, n38440, n38441, n38442,
         n38443, n38444, n38445, n38446, n38447, n38448, n38449, n38450,
         n38451, n38452, n38453, n38454, n38455, n38456, n38457, n38458,
         n38459, n38460, n38461, n38462, n38463, n38464, n38465, n38466,
         n38467, n38468, n38469, n38470, n38471, n38472, n38473, n38474,
         n38475, n38476, n38477, n38478, n38479, n38480, n38481, n38482,
         n38483, n38484, n38485, n38486, n38487, n38488, n38489, n38490,
         n38491, n38492, n38493, n38494, n38495, n38496, n38497, n38498,
         n38499, n38500, n38501, n38502, n38503, n38504, n38505, n38506,
         n38507, n38508, n38509, n38510, n38511, n38512, n38513, n38514,
         n38515, n38516, n38517, n38518, n38519, n38520, n38521, n38522,
         n38523, n38524, n38525, n38526, n38527, n38528, n38529, n38530,
         n38531, n38532, n38533, n38534, n38535, n38536, n38537, n38538,
         n38539, n38540, n38541, n38542, n38543, n38544, n38545, n38546,
         n38547, n38548, n38549, n38550, n38551, n38552, n38553, n38554,
         n38555, n38556, n38557, n38558, n38559, n38560, n38561, n38562,
         n38563, n38564, n38565, n38566, n38567, n38568, n38569, n38570,
         n38571, n38572, n38573, n38574, n38575, n38576, n38577, n38578,
         n38579, n38580, n38581, n38582, n38583, n38584, n38585, n38586,
         n38587, n38588, n38589, n38590, n38591, n38592, n38593, n38594,
         n38595, n38596, n38597, n38598, n38599, n38600, n38601, n38602,
         n38603, n38604, n38605, n38606, n38607, n38608, n38609, n38610,
         n38611, n38612, n38613, n38614, n38615, n38616, n38617, n38618,
         n38619, n38620, n38621, n38622, n38623, n38624, n38625, n38626,
         n38627, n38628, n38629, n38630, n38631, n38632, n38633, n38634,
         n38635, n38636, n38637, n38638, n38639, n38640, n38641, n38642,
         n38643, n38644, n38645, n38646, n38647, n38648, n38649, n38650,
         n38651, n38652, n38653, n38654, n38655, n38656, n38657, n38658,
         n38659, n38660, n38661, n38662, n38663, n38664, n38665, n38666,
         n38667, n38668, n38669, n38670, n38671, n38672, n38673, n38674,
         n38675, n38676, n38677, n38678, n38679, n38680, n38681, n38682,
         n38683, n38684, n38685, n38686, n38687, n38688, n38689, n38690,
         n38691, n38692, n38693, n38694, n38695, n38696, n38697, n38698,
         n38699, n38700, n38701, n38702, n38703, n38704, n38705, n38706,
         n38707, n38708, n38709, n38710, n38711, n38712, n38713, n38714,
         n38715, n38716, n38717, n38718, n38719, n38720, n38721, n38722,
         n38723, n38724, n38725, n38726, n38727, n38728, n38729, n38730,
         n38731, n38732, n38733, n38734, n38735, n38736, n38737, n38738,
         n38739, n38740, n38741, n38742, n38743, n38744, n38745, n38746,
         n38747, n38748, n38749, n38750, n38751, n38752, n38753, n38754,
         n38755, n38756, n38757, n38758, n38759, n38760, n38761, n38762,
         n38763, n38764, n38765, n38766, n38767, n38768, n38769, n38770,
         n38771, n38772, n38773, n38774, n38775, n38776, n38777, n38778,
         n38779, n38780, n38781, n38782, n38783, n38784, n38785, n38786,
         n38787, n38788, n38789, n38790, n38791, n38792, n38793, n38794,
         n38795, n38796, n38797, n38798, n38799, n38800, n38801, n38802,
         n38803, n38804, n38805, n38806, n38807, n38808, n38809, n38810,
         n38811, n38812, n38813, n38814, n38815, n38816, n38817, n38818,
         n38819, n38820, n38821, n38822, n38823, n38824, n38825, n38826,
         n38827, n38828, n38829, n38830, n38831, n38832, n38833, n38834,
         n38835, n38836, n38837, n38838, n38839, n38840, n38841, n38842,
         n38843, n38844, n38845, n38846, n38847, n38848, n38849, n38850,
         n38851, n38852, n38853, n38854, n38855, n38856, n38857, n38858,
         n38859, n38860, n38861, n38862, n38863, n38864, n38865, n38866,
         n38867, n38868, n38869, n38870, n38871, n38872, n38873, n38874,
         n38875, n38876, n38877, n38878, n38879, n38880, n38881, n38882,
         n38883, n38884, n38885, n38886, n38887, n38888, n38889, n38890,
         n38891, n38892, n38893, n38894, n38895, n38896, n38897, n38898,
         n38899, n38900, n38901, n38902, n38903, n38904, n38905, n38906,
         n38907, n38908, n38909, n38910, n38911, n38912, n38913, n38914,
         n38915, n38916, n38917, n38918, n38919, n38920, n38921, n38922,
         n38923, n38924, n38925, n38926, n38927, n38928, n38929, n38930,
         n38931, n38932, n38933, n38934, n38935, n38936, n38937, n38938,
         n38939, n38940, n38941, n38942, n38943, n38944, n38945, n38946,
         n38947, n38948, n38949, n38950, n38951, n38952, n38953, n38954,
         n38955, n38956, n38957, n38958, n38959, n38960, n38961, n38962,
         n38963, n38964, n38965, n38966, n38967, n38968, n38969, n38970,
         n38971, n38972, n38973, n38974, n38975, n38976, n38977, n38978,
         n38979, n38980, n38981, n38982, n38983, n38984, n38985, n38986,
         n38987, n38988, n38989, n38990, n38991, n38992, n38993, n38994,
         n38995, n38996, n38997, n38998, n38999, n39000, n39001, n39002,
         n39003, n39004, n39005, n39006, n39007, n39008, n39009, n39010,
         n39011, n39012, n39013, n39014, n39015, n39016, n39017, n39018,
         n39019, n39020, n39021, n39022, n39023, n39024, n39025, n39026,
         n39027, n39028, n39029, n39030, n39031, n39032, n39033, n39034,
         n39035, n39036, n39037, n39038, n39039, n39040, n39041, n39042,
         n39043, n39044, n39045, n39046, n39047, n39048, n39049, n39050,
         n39051, n39052, n39053, n39054, n39055, n39056, n39057, n39058,
         n39059, n39060, n39061, n39062, n39063, n39064, n39065, n39066,
         n39067, n39068, n39069, n39070, n39071, n39072, n39073, n39074,
         n39075, n39076, n39077, n39078, n39079, n39080, n39081, n39082,
         n39083, n39084, n39085, n39086, n39087, n39088, n39089, n39090,
         n39091, n39092, n39093, n39094, n39095, n39096, n39097, n39098,
         n39099, n39100, n39101, n39102, n39103, n39104, n39105, n39106,
         n39107, n39108, n39109, n39110, n39111, n39112, n39113, n39114,
         n39115, n39116, n39117, n39118, n39119, n39120, n39121, n39122,
         n39123, n39124, n39125, n39126, n39127, n39128, n39129, n39130,
         n39131, n39132, n39133, n39134, n39135, n39136, n39137, n39138,
         n39139, n39140, n39141, n39142, n39143, n39144, n39145, n39146,
         n39147, n39148, n39149, n39150, n39151, n39152, n39153, n39154,
         n39155, n39156, n39157, n39158, n39159, n39160, n39161, n39162,
         n39163, n39164, n39165, n39166, n39167, n39168, n39169, n39170,
         n39171, n39172, n39173, n39174, n39175, n39176, n39177, n39178,
         n39179, n39180, n39181, n39182, n39183, n39184, n39185, n39186,
         n39187, n39188, n39189, n39190, n39191, n39192, n39193, n39194,
         n39195, n39196, n39197, n39198, n39199, n39200, n39201, n39202,
         n39203, n39204, n39205, n39206, n39207, n39208, n39209, n39210,
         n39211, n39212, n39213, n39214, n39215, n39216, n39217, n39218,
         n39219, n39220, n39221, n39222, n39223, n39224, n39225, n39226,
         n39227, n39228, n39229, n39230, n39231, n39232, n39233, n39234,
         n39235, n39236, n39237, n39238, n39239, n39240, n39241, n39242,
         n39243, n39244, n39245, n39246, n39247, n39248, n39249, n39250,
         n39251, n39252, n39253, n39254, n39255, n39256, n39257, n39258,
         n39259, n39260, n39261, n39262, n39263, n39264, n39265, n39266,
         n39267, n39268, n39269, n39270, n39271, n39272, n39273, n39274,
         n39275, n39276, n39277, n39278, n39279, n39280, n39281, n39282,
         n39283, n39284, n39285, n39286, n39287, n39288, n39289, n39290,
         n39291, n39292, n39293, n39294, n39295, n39296, n39297, n39298,
         n39299, n39300, n39301, n39302, n39303, n39304, n39305, n39306,
         n39307, n39308, n39309, n39310, n39311, n39312, n39313, n39314,
         n39315, n39316, n39317, n39318, n39319, n39320, n39321, n39322,
         n39323, n39324, n39325, n39326, n39327, n39328, n39329, n39330,
         n39331, n39332, n39333, n39334, n39335, n39336, n39337, n39338,
         n39339, n39340, n39341, n39342, n39343, n39344, n39345, n39346,
         n39347, n39348, n39349, n39350, n39351, n39352, n39353, n39354,
         n39355, n39356, n39357, n39358, n39359, n39360, n39361, n39362,
         n39363, n39364, n39365, n39366, n39367, n39368, n39369, n39370,
         n39371, n39372, n39373, n39374, n39375, n39376, n39377, n39378,
         n39379, n39380, n39381, n39382, n39383, n39384, n39385, n39386,
         n39387, n39388, n39389, n39390, n39391, n39392, n39393, n39394,
         n39395, n39396, n39397, n39398, n39399, n39400, n39401, n39402,
         n39403, n39404, n39405, n39406, n39407, n39408, n39409, n39410,
         n39411, n39412, n39413, n39414, n39415, n39416, n39417, n39418,
         n39419, n39420, n39421, n39422, n39423, n39424, n39425, n39426,
         n39427, n39428, n39429, n39430, n39431, n39432, n39433, n39434,
         n39435, n39436, n39437, n39438, n39439, n39440, n39441, n39442,
         n39443, n39444, n39445, n39446, n39447, n39448, n39449, n39450,
         n39451, n39452, n39453, n39454, n39455, n39456, n39457, n39458,
         n39459, n39460, n39461, n39462, n39463, n39464, n39465, n39466,
         n39467, n39468, n39469, n39470, n39471, n39472, n39473, n39474,
         n39475, n39476, n39477, n39478, n39479, n39480, n39481, n39482,
         n39483, n39484, n39485, n39486, n39487, n39488, n39489, n39490,
         n39491, n39492, n39493, n39494, n39495, n39496, n39497, n39498,
         n39499, n39500, n39501, n39502, n39503, n39504, n39505, n39506,
         n39507, n39508, n39509, n39510, n39511, n39512, n39513, n39514,
         n39515, n39516, n39517, n39518, n39519, n39520, n39521, n39522,
         n39523, n39524, n39525, n39526, n39527, n39528, n39529, n39530,
         n39531, n39532, n39533, n39534, n39535, n39536, n39537, n39538,
         n39539, n39540, n39541, n39542, n39543, n39544, n39545, n39546,
         n39547, n39548, n39549, n39550, n39551, n39552, n39553, n39554,
         n39555, n39556, n39557, n39558, n39559, n39560, n39561, n39562,
         n39563, n39564, n39565, n39566, n39567, n39568, n39569, n39570,
         n39571, n39572, n39573, n39574, n39575, n39576, n39577, n39578,
         n39579, n39580, n39581, n39582, n39583, n39584, n39585, n39586,
         n39587, n39588, n39589, n39590, n39591, n39592, n39593, n39594,
         n39595, n39596, n39597, n39598, n39599, n39600, n39601, n39602,
         n39603, n39604, n39605, n39606, n39607, n39608, n39609, n39610,
         n39611, n39612, n39613, n39614, n39615, n39616, n39617, n39618,
         n39619, n39620, n39621, n39622, n39623, n39624, n39625, n39626,
         n39627, n39628, n39629, n39630, n39631, n39632, n39633, n39634,
         n39635, n39636, n39637, n39638, n39639, n39640, n39641, n39642,
         n39643, n39644, n39645, n39646, n39647, n39648, n39649, n39650,
         n39651, n39652, n39653, n39654, n39655, n39656, n39657, n39658,
         n39659, n39660, n39661, n39662, n39663, n39664, n39665, n39666,
         n39667, n39668, n39669, n39670, n39671, n39672, n39673, n39674,
         n39675, n39676, n39677, n39678, n39679, n39680, n39681, n39682,
         n39683, n39684, n39685, n39686, n39687, n39688, n39689, n39690,
         n39691, n39692, n39693, n39694, n39695, n39696, n39697, n39698,
         n39699, n39700, n39701, n39702, n39703, n39704, n39705, n39706,
         n39707, n39708, n39709, n39710, n39711, n39712, n39713, n39714,
         n39715, n39716, n39717, n39718, n39719, n39720, n39721, n39722,
         n39723, n39724, n39725, n39726, n39727, n39728, n39729, n39730,
         n39731, n39732, n39733, n39734, n39735, n39736, n39737, n39738,
         n39739, n39740, n39741, n39742, n39743, n39744, n39745, n39746,
         n39747, n39748, n39749, n39750, n39751, n39752, n39753, n39754,
         n39755, n39756, n39757, n39758, n39759, n39760, n39761, n39762,
         n39763, n39764, n39765, n39766, n39767, n39768, n39769, n39770,
         n39771, n39772, n39773, n39774, n39775, n39776, n39777, n39778,
         n39779, n39780, n39781, n39782, n39783, n39784, n39785, n39786,
         n39787, n39788, n39789, n39790, n39791, n39792, n39793, n39794,
         n39795, n39796, n39797, n39798, n39799, n39800, n39801, n39802,
         n39803, n39804, n39805, n39806, n39807, n39808, n39809, n39810,
         n39811, n39812, n39813, n39814, n39815, n39816, n39817, n39818,
         n39819, n39820, n39821, n39822, n39823, n39824, n39825, n39826,
         n39827, n39828, n39829, n39830, n39831, n39832, n39833, n39834,
         n39835, n39836, n39837, n39838, n39839, n39840, n39841, n39842,
         n39843, n39844, n39845, n39846, n39847, n39848, n39849, n39850,
         n39851, n39852, n39853, n39854, n39855, n39856, n39857, n39858,
         n39859, n39860, n39861, n39862, n39863, n39864, n39865, n39866,
         n39867, n39868, n39869, n39870, n39871, n39872, n39873, n39874,
         n39875, n39876, n39877, n39878, n39879, n39880, n39881, n39882,
         n39883, n39884, n39885, n39886, n39887, n39888, n39889, n39890,
         n39891, n39892, n39893, n39894, n39895, n39896, n39897, n39898,
         n39899, n39900, n39901, n39902, n39903, n39904, n39905, n39906,
         n39907, n39908, n39909, n39910, n39911, n39912, n39913, n39914,
         n39915, n39916, n39917, n39918, n39919, n39920, n39921, n39922,
         n39923, n39924, n39925, n39926, n39927, n39928, n39929, n39930,
         n39931, n39932, n39933, n39934, n39935, n39936, n39937, n39938,
         n39939, n39940, n39941, n39942, n39943, n39944, n39945, n39946,
         n39947, n39948, n39949, n39950, n39951, n39952, n39953, n39954,
         n39955, n39956, n39957, n39958, n39959, n39960, n39961, n39962,
         n39963, n39964, n39965, n39966, n39967, n39968, n39969, n39970,
         n39971, n39972, n39973, n39974, n39975, n39976, n39977, n39978,
         n39979, n39980, n39981, n39982, n39983, n39984, n39985, n39986,
         n39987, n39988, n39989, n39990, n39991, n39992, n39993, n39994,
         n39995, n39996, n39997, n39998, n39999, n40000, n40001, n40002,
         n40003, n40004, n40005, n40006, n40007, n40008, n40009, n40010,
         n40011, n40012, n40013, n40014, n40015, n40016, n40017, n40018,
         n40019, n40020, n40021, n40022, n40023, n40024, n40025, n40026,
         n40027, n40028, n40029, n40030, n40031, n40032, n40033, n40034,
         n40035, n40036, n40037, n40038, n40039, n40040, n40041, n40042,
         n40043, n40044, n40045, n40046, n40047, n40048, n40049, n40050,
         n40051, n40052, n40053, n40054, n40055, n40056, n40057, n40058,
         n40059, n40060, n40061, n40062, n40063, n40064, n40065, n40066,
         n40067, n40068, n40069, n40070, n40071, n40072, n40073, n40074,
         n40075, n40076, n40077, n40078, n40079, n40080, n40081, n40082,
         n40083, n40084, n40085, n40086, n40087, n40088, n40089, n40090,
         n40091, n40092, n40093, n40094, n40095, n40096, n40097, n40098,
         n40099, n40100, n40101, n40102, n40103, n40104, n40105, n40106,
         n40107, n40108, n40109, n40110, n40111, n40112, n40113, n40114,
         n40115, n40116, n40117, n40118, n40119, n40120, n40121, n40122,
         n40123, n40124, n40125, n40126, n40127, n40128, n40129, n40130,
         n40131, n40132, n40133, n40134, n40135, n40136, n40137, n40138,
         n40139, n40140, n40141, n40142, n40143, n40144, n40145, n40146,
         n40147, n40148, n40149, n40150, n40151, n40152, n40153, n40154,
         n40155, n40156, n40157, n40158, n40159, n40160, n40161, n40162,
         n40163, n40164, n40165, n40166, n40167, n40168, n40169, n40170,
         n40171, n40172, n40173, n40174, n40175, n40176, n40177, n40178,
         n40179, n40180, n40181, n40182, n40183, n40184, n40185, n40186,
         n40187, n40188, n40189, n40190, n40191, n40192, n40193, n40194,
         n40195, n40196, n40197, n40198, n40199, n40200, n40201, n40202,
         n40203, n40204, n40205, n40206, n40207, n40208, n40209, n40210,
         n40211, n40212, n40213, n40214, n40215, n40216, n40217, n40218,
         n40219, n40220, n40221, n40222, n40223, n40224, n40225, n40226,
         n40227, n40228, n40229, n40230, n40231, n40232, n40233, n40234,
         n40235, n40236, n40237, n40238, n40239, n40240, n40241, n40242,
         n40243, n40244, n40245, n40246, n40247, n40248, n40249, n40250,
         n40251, n40252, n40253, n40254, n40255, n40256, n40257, n40258,
         n40259, n40260, n40261, n40262, n40263, n40264, n40265, n40266,
         n40267, n40268, n40269, n40270, n40271, n40272, n40273, n40274,
         n40275, n40276, n40277, n40278, n40279, n40280, n40281, n40282,
         n40283, n40284, n40285, n40286, n40287, n40288, n40289, n40290,
         n40291, n40292, n40293, n40294, n40295, n40296, n40297, n40298,
         n40299, n40300, n40301, n40302, n40303, n40304, n40305, n40306,
         n40307, n40308, n40309, n40310, n40311, n40312, n40313, n40314,
         n40315, n40316, n40317, n40318, n40319, n40320, n40321, n40322,
         n40323, n40324, n40325, n40326, n40327, n40328, n40329, n40330,
         n40331, n40332, n40333, n40334, n40335, n40336, n40337, n40338,
         n40339, n40340, n40341, n40342, n40343, n40344, n40345, n40346,
         n40347, n40348, n40349, n40350, n40351, n40352, n40353, n40354,
         n40355, n40356, n40357, n40358, n40359, n40360, n40361, n40362,
         n40363, n40364, n40365, n40366, n40367, n40368, n40369, n40370,
         n40371, n40372, n40373, n40374, n40375, n40376, n40377, n40378,
         n40379, n40380, n40381, n40382, n40383, n40384, n40385, n40386,
         n40387, n40388, n40389, n40390, n40391, n40392, n40393, n40394,
         n40395, n40396, n40397, n40398, n40399, n40400, n40401, n40402,
         n40403, n40404, n40405, n40406, n40407, n40408, n40409, n40410,
         n40411, n40412, n40413, n40414, n40415, n40416, n40417, n40418,
         n40419, n40420, n40421, n40422, n40423, n40424, n40425, n40426,
         n40427, n40428, n40429, n40430, n40431, n40432, n40433, n40434,
         n40435, n40436, n40437, n40438, n40439, n40440, n40441, n40442,
         n40443, n40444, n40445, n40446, n40447, n40448, n40449, n40450,
         n40451, n40452, n40453, n40454, n40455, n40456, n40457, n40458,
         n40459, n40460, n40461, n40462, n40463, n40464, n40465, n40466,
         n40467, n40468, n40469, n40470, n40471, n40472, n40473, n40474,
         n40475, n40476, n40477, n40478, n40479, n40480, n40481, n40482,
         n40483, n40484, n40485, n40486, n40487, n40488, n40489, n40490,
         n40491, n40492, n40493, n40494, n40495, n40496, n40497, n40498,
         n40499, n40500, n40501, n40502, n40503, n40504, n40505, n40506,
         n40507, n40508, n40509, n40510, n40511, n40512, n40513, n40514,
         n40515, n40516, n40517, n40518, n40519, n40520, n40521, n40522,
         n40523, n40524, n40525, n40526, n40527, n40528, n40529, n40530,
         n40531, n40532, n40533, n40534, n40535, n40536, n40537, n40538,
         n40539, n40540, n40541, n40542, n40543, n40544, n40545, n40546,
         n40547, n40548, n40549, n40550, n40551, n40552, n40553, n40554,
         n40555, n40556, n40557, n40558, n40559, n40560, n40561, n40562,
         n40563, n40564, n40565, n40566, n40567, n40568, n40569, n40570,
         n40571, n40572, n40573, n40574, n40575, n40576, n40577, n40578,
         n40579, n40580, n40581, n40582, n40583, n40584, n40585, n40586,
         n40587, n40588, n40589, n40590, n40591, n40592, n40593, n40594,
         n40595, n40596, n40597, n40598, n40599, n40600, n40601, n40602,
         n40603, n40604, n40605, n40606, n40607, n40608, n40609, n40610,
         n40611, n40612, n40613, n40614, n40615, n40616, n40617, n40618,
         n40619, n40620, n40621, n40622, n40623, n40624, n40625, n40626,
         n40627, n40628, n40629, n40630, n40631, n40632, n40633, n40634,
         n40635, n40636, n40637, n40638, n40639, n40640, n40641, n40642,
         n40643, n40644, n40645, n40646, n40647, n40648, n40649, n40650,
         n40651, n40652, n40653, n40654, n40655, n40656, n40657, n40658,
         n40659, n40660, n40661, n40662, n40663, n40664, n40665, n40666,
         n40667, n40668, n40669, n40670, n40671, n40672, n40673, n40674,
         n40675, n40676, n40677, n40678, n40679, n40680, n40681, n40682,
         n40683, n40684, n40685, n40686, n40687, n40688, n40689, n40690,
         n40691, n40692, n40693, n40694, n40695, n40696, n40697, n40698,
         n40699, n40700, n40701, n40702, n40703, n40704, n40705, n40706,
         n40707, n40708, n40709, n40710, n40711, n40712, n40713, n40714,
         n40715, n40716, n40717, n40718, n40719, n40720, n40721, n40722,
         n40723, n40724, n40725, n40726, n40727, n40728, n40729, n40730,
         n40731, n40732, n40733, n40734, n40735, n40736, n40737, n40738,
         n40739, n40740, n40741, n40742, n40743, n40744, n40745, n40746,
         n40747, n40748, n40749, n40750, n40751, n40752, n40753, n40754,
         n40755, n40756, n40757, n40758, n40759, n40760, n40761, n40762,
         n40763, n40764, n40765, n40766, n40767, n40768, n40769, n40770,
         n40771, n40772, n40773, n40774, n40775, n40776, n40777, n40778,
         n40779, n40780, n40781, n40782, n40783, n40784, n40785, n40786,
         n40787, n40788, n40789, n40790, n40791, n40792, n40793, n40794,
         n40795, n40796, n40797, n40798, n40799, n40800, n40801, n40802,
         n40803, n40804, n40805, n40806, n40807, n40808, n40809, n40810,
         n40811, n40812, n40813, n40814, n40815, n40816, n40817, n40818,
         n40819, n40820, n40821, n40822, n40823, n40824, n40825, n40826,
         n40827, n40828, n40829, n40830, n40831, n40832, n40833, n40834,
         n40835, n40836, n40837, n40838, n40839, n40840, n40841, n40842,
         n40843, n40844, n40845, n40846, n40847, n40848, n40849, n40850,
         n40851, n40852, n40853, n40854, n40855, n40856, n40857, n40858,
         n40859, n40860, n40861, n40862, n40863, n40864, n40865, n40866,
         n40867, n40868, n40869, n40870, n40871, n40872, n40873, n40874,
         n40875, n40876, n40877, n40878, n40879, n40880, n40881, n40882,
         n40883, n40884, n40885, n40886, n40887, n40888, n40889, n40890,
         n40891, n40892, n40893, n40894, n40895, n40896, n40897, n40898,
         n40899, n40900, n40901, n40902, n40903, n40904, n40905, n40906,
         n40907, n40908, n40909, n40910, n40911, n40912, n40913, n40914,
         n40915, n40916, n40917, n40918, n40919, n40920, n40921, n40922,
         n40923, n40924, n40925, n40926, n40927, n40928, n40929, n40930,
         n40931, n40932, n40933, n40934, n40935, n40936, n40937, n40938,
         n40939, n40940, n40941, n40942, n40943, n40944, n40945, n40946,
         n40947, n40948, n40949, n40950, n40951, n40952, n40953, n40954,
         n40955, n40956, n40957, n40958, n40959, n40960, n40961, n40962,
         n40963, n40964, n40965, n40966, n40967, n40968, n40969, n40970,
         n40971, n40972, n40973, n40974, n40975, n40976, n40977, n40978,
         n40979, n40980, n40981, n40982, n40983, n40984, n40985, n40986,
         n40987, n40988, n40989, n40990, n40991, n40992, n40993, n40994,
         n40995, n40996, n40997, n40998, n40999, n41000, n41001, n41002,
         n41003, n41004, n41005, n41006, n41007, n41008, n41009, n41010,
         n41011, n41012, n41013, n41014, n41015, n41016, n41017, n41018,
         n41019, n41020, n41021, n41022, n41023, n41024, n41025, n41026,
         n41027, n41028, n41029, n41030, n41031, n41032, n41033, n41034,
         n41035, n41036, n41037, n41038, n41039, n41040, n41041, n41042,
         n41043, n41044, n41045, n41046, n41047, n41048, n41049, n41050,
         n41051, n41052, n41053, n41054, n41055, n41056, n41057, n41058,
         n41059, n41060, n41061, n41062, n41063, n41064, n41065, n41066,
         n41067, n41068, n41069, n41070, n41071, n41072, n41073, n41074,
         n41075, n41076, n41077, n41078, n41079, n41080, n41081, n41082,
         n41083, n41084, n41085, n41086, n41087, n41088, n41089, n41090,
         n41091, n41092, n41093, n41094, n41095, n41096, n41097, n41098,
         n41099, n41100, n41101, n41102, n41103, n41104, n41105, n41106,
         n41107, n41108, n41109, n41110, n41111, n41112, n41113, n41114,
         n41115, n41116, n41117, n41118, n41119, n41120, n41121, n41122,
         n41123, n41124, n41125, n41126, n41127, n41128, n41129, n41130,
         n41131, n41132, n41133, n41134, n41135, n41136, n41137, n41138,
         n41139, n41140, n41141, n41142, n41143, n41144, n41145, n41146,
         n41147, n41148, n41149, n41150, n41151, n41152, n41153, n41154,
         n41155, n41156, n41157, n41158, n41159, n41160, n41161, n41162,
         n41163, n41164, n41165, n41166, n41167, n41168, n41169, n41170,
         n41171, n41172, n41173, n41174, n41175, n41176, n41177, n41178,
         n41179, n41180, n41181, n41182, n41183, n41184, n41185, n41186,
         n41187, n41188, n41189, n41190, n41191, n41192, n41193, n41194,
         n41195, n41196, n41197, n41198, n41199, n41200, n41201, n41202,
         n41203, n41204, n41205, n41206, n41207, n41208, n41209, n41210,
         n41211, n41212, n41213, n41214, n41215, n41216, n41217, n41218,
         n41219, n41220, n41221, n41222, n41223, n41224, n41225, n41226,
         n41227, n41228, n41229, n41230, n41231, n41232, n41233, n41234,
         n41235, n41236, n41237, n41238, n41239, n41240, n41241, n41242,
         n41243, n41244, n41245, n41246, n41247, n41248, n41249, n41250,
         n41251, n41252, n41253, n41254, n41255, n41256, n41257, n41258,
         n41259, n41260, n41261, n41262, n41263, n41264, n41265, n41266,
         n41267, n41268, n41269, n41270, n41271, n41272, n41273, n41274,
         n41275, n41276, n41277, n41278, n41279, n41280, n41281, n41282,
         n41283, n41284, n41285, n41286, n41287, n41288, n41289, n41290,
         n41291, n41292, n41293, n41294, n41295, n41296, n41297, n41298,
         n41299, n41300, n41301, n41302, n41303, n41304, n41305, n41306,
         n41307, n41308, n41309, n41310, n41311, n41312, n41313, n41314,
         n41315, n41316, n41317, n41318, n41319, n41320, n41321, n41322,
         n41323, n41324, n41325, n41326, n41327, n41328, n41329, n41330,
         n41331, n41332, n41333, n41334, n41335, n41336, n41337, n41338,
         n41339, n41340, n41341, n41342, n41343, n41344, n41345, n41346,
         n41347, n41348, n41349, n41350, n41351, n41352, n41353, n41354,
         n41355, n41356, n41357, n41358, n41359, n41360, n41361, n41362,
         n41363, n41364, n41365, n41366, n41367, n41368, n41369, n41370,
         n41371, n41372, n41373, n41374, n41375, n41376, n41377, n41378,
         n41379, n41380, n41381, n41382, n41383, n41384, n41385, n41386,
         n41387, n41388, n41389, n41390, n41391, n41392, n41393, n41394,
         n41395, n41396, n41397, n41398, n41399, n41400, n41401, n41402,
         n41403, n41404, n41405, n41406, n41407, n41408, n41409, n41410,
         n41411, n41412, n41413, n41414, n41415, n41416, n41417, n41418,
         n41419, n41420, n41421, n41422, n41423, n41424, n41425, n41426,
         n41427, n41428, n41429, n41430, n41431, n41432, n41433, n41434,
         n41435, n41436, n41437, n41438, n41439, n41440, n41441, n41442,
         n41443, n41444, n41445, n41446, n41447, n41448, n41449, n41450,
         n41451, n41452, n41453, n41454, n41455, n41456, n41457, n41458,
         n41459, n41460, n41461, n41462, n41463, n41464, n41465, n41466,
         n41467, n41468, n41469, n41470, n41471, n41472, n41473, n41474,
         n41475, n41476, n41477, n41478, n41479, n41480, n41481, n41482,
         n41483, n41484, n41485, n41486, n41487, n41488, n41489, n41490,
         n41491, n41492, n41493, n41494, n41495, n41496, n41497, n41498,
         n41499, n41500, n41501, n41502, n41503, n41504, n41505, n41506,
         n41507, n41508, n41509, n41510, n41511, n41512, n41513, n41514,
         n41515, n41516, n41517, n41518, n41519, n41520, n41521, n41522,
         n41523, n41524, n41525, n41526, n41527, n41528, n41529, n41530,
         n41531, n41532, n41533, n41534, n41535, n41536, n41537, n41538,
         n41539, n41540, n41541, n41542, n41543, n41544, n41545, n41546,
         n41547, n41548, n41549, n41550, n41551, n41552, n41553, n41554,
         n41555, n41556, n41557, n41558, n41559, n41560, n41561, n41562,
         n41563, n41564, n41565, n41566, n41567, n41568, n41569, n41570,
         n41571, n41572, n41573, n41574, n41575, n41576, n41577, n41578,
         n41579, n41580, n41581, n41582, n41583, n41584, n41585, n41586,
         n41587, n41588, n41589, n41590, n41591, n41592, n41593, n41594,
         n41595, n41596, n41597, n41598, n41599, n41600, n41601, n41602,
         n41603, n41604, n41605, n41606, n41607, n41608, n41609, n41610,
         n41611, n41612, n41613, n41614, n41615, n41616, n41617, n41618,
         n41619, n41620, n41621, n41622, n41623, n41624, n41625, n41626,
         n41627, n41628, n41629, n41630, n41631, n41632, n41633, n41634,
         n41635, n41636, n41637, n41638, n41639, n41640, n41641, n41642,
         n41643, n41644, n41645, n41646, n41647, n41648, n41649, n41650,
         n41651, n41652, n41653, n41654, n41655, n41656, n41657, n41658,
         n41659, n41660, n41661, n41662, n41663, n41664, n41665, n41666,
         n41667, n41668, n41669, n41670, n41671, n41672, n41673, n41674,
         n41675, n41676, n41677, n41678, n41679, n41680, n41681, n41682,
         n41683, n41684, n41685, n41686, n41687, n41688, n41689, n41690,
         n41691, n41692, n41693, n41694, n41695, n41696, n41697, n41698,
         n41699, n41700, n41701, n41702, n41703, n41704, n41705, n41706,
         n41707, n41708, n41709, n41710, n41711, n41712, n41713, n41714,
         n41715, n41716, n41717, n41718, n41719, n41720, n41721, n41722,
         n41723, n41724, n41725, n41726, n41727, n41728, n41729, n41730,
         n41731, n41732, n41733, n41734, n41735, n41736, n41737, n41738,
         n41739, n41740, n41741, n41742, n41743, n41744, n41745, n41746,
         n41747, n41748, n41749, n41750, n41751, n41752, n41753, n41754,
         n41755, n41756, n41757, n41758, n41759, n41760, n41761, n41762,
         n41763, n41764, n41765, n41766, n41767, n41768, n41769, n41770,
         n41771, n41772, n41773, n41774, n41775, n41776, n41777, n41778,
         n41779, n41780, n41781, n41782, n41783, n41784, n41785, n41786,
         n41787, n41788, n41789, n41790, n41791, n41792, n41793, n41794,
         n41795, n41796, n41797, n41798, n41799, n41800, n41801, n41802,
         n41803, n41804, n41805, n41806, n41807, n41808, n41809, n41810,
         n41811, n41812, n41813, n41814, n41815, n41816, n41817, n41818,
         n41819, n41820, n41821, n41822, n41823, n41824, n41825, n41826,
         n41827, n41828, n41829, n41830, n41831, n41832, n41833, n41834,
         n41835, n41836, n41837, n41838, n41839, n41840, n41841, n41842,
         n41843, n41844, n41845, n41846, n41847, n41848, n41849, n41850,
         n41851, n41852, n41853, n41854, n41855, n41856, n41857, n41858,
         n41859, n41860, n41861, n41862, n41863, n41864, n41865, n41866,
         n41867, n41868, n41869, n41870, n41871, n41872, n41873, n41874,
         n41875, n41876, n41877, n41878, n41879, n41880, n41881, n41882,
         n41883, n41884, n41885, n41886, n41887, n41888, n41889, n41890,
         n41891, n41892, n41893, n41894, n41895, n41896, n41897, n41898,
         n41899, n41900, n41901, n41902, n41903, n41904, n41905, n41906,
         n41907, n41908, n41909, n41910, n41911, n41912, n41913, n41914,
         n41915, n41916, n41917, n41918, n41919, n41920, n41921, n41922,
         n41923, n41924, n41925, n41926, n41927, n41928, n41929, n41930,
         n41931, n41932, n41933, n41934, n41935, n41936, n41937, n41938,
         n41939, n41940, n41941, n41942, n41943, n41944, n41945, n41946,
         n41947, n41948, n41949, n41950, n41951, n41952, n41953, n41954,
         n41955, n41956, n41957, n41958, n41959, n41960, n41961, n41962,
         n41963, n41964, n41965, n41966, n41967, n41968, n41969, n41970,
         n41971, n41972, n41973, n41974, n41975, n41976, n41977, n41978,
         n41979, n41980, n41981, n41982, n41983, n41984, n41985, n41986,
         n41987, n41988, n41989, n41990, n41991, n41992, n41993, n41994,
         n41995, n41996, n41997, n41998, n41999, n42000, n42001, n42002,
         n42003, n42004, n42005, n42006, n42007, n42008, n42009, n42010,
         n42011, n42012, n42013, n42014, n42015, n42016, n42017, n42018,
         n42019, n42020, n42021, n42022, n42023, n42024, n42025, n42026,
         n42027, n42028, n42029, n42030, n42031, n42032, n42033, n42034,
         n42035, n42036, n42037, n42038, n42039, n42040, n42041, n42042,
         n42043, n42044, n42045, n42046, n42047, n42048, n42049, n42050,
         n42051, n42052, n42053, n42054, n42055, n42056, n42057, n42058,
         n42059, n42060, n42061, n42062, n42063, n42064, n42065, n42066,
         n42067, n42068, n42069, n42070, n42071, n42072, n42073, n42074,
         n42075, n42076, n42077, n42078, n42079, n42080, n42081, n42082,
         n42083, n42084, n42085, n42086, n42087, n42088, n42089, n42090,
         n42091, n42092, n42093, n42094, n42095, n42096, n42097, n42098,
         n42099, n42100, n42101, n42102, n42103, n42104, n42105, n42106,
         n42107, n42108, n42109, n42110, n42111, n42112, n42113, n42114,
         n42115, n42116, n42117, n42118, n42119, n42120, n42121, n42122,
         n42123, n42124, n42125, n42126, n42127, n42128, n42129, n42130,
         n42131, n42132, n42133, n42134, n42135, n42136, n42137, n42138,
         n42139, n42140, n42141, n42142, n42143, n42144, n42145, n42146,
         n42147, n42148, n42149, n42150, n42151, n42152, n42153, n42154,
         n42155, n42156, n42157, n42158, n42159, n42160, n42161, n42162,
         n42163, n42164, n42165, n42166, n42167, n42168, n42169, n42170,
         n42171, n42172, n42173, n42174, n42175, n42176, n42177, n42178,
         n42179, n42180, n42181, n42182, n42183, n42184, n42185, n42186,
         n42187, n42188, n42189, n42190, n42191, n42192, n42193, n42194,
         n42195, n42196, n42197, n42198, n42199, n42200, n42201, n42202,
         n42203, n42204, n42205, n42206, n42207, n42208, n42209, n42210,
         n42211, n42212, n42213, n42214, n42215, n42216, n42217, n42218,
         n42219, n42220, n42221, n42222, n42223, n42224, n42225, n42226,
         n42227, n42228, n42229, n42230, n42231, n42232, n42233, n42234,
         n42235, n42236, n42237, n42238, n42239, n42240, n42241, n42242,
         n42243, n42244, n42245, n42246, n42247, n42248, n42249, n42250,
         n42251, n42252, n42253, n42254, n42255, n42256, n42257, n42258,
         n42259, n42260, n42261, n42262, n42263, n42264, n42265, n42266,
         n42267, n42268, n42269, n42270, n42271, n42272, n42273, n42274,
         n42275, n42276, n42277, n42278, n42279, n42280, n42281, n42282,
         n42283, n42284, n42285, n42286, n42287, n42288, n42289, n42290,
         n42291, n42292, n42293, n42294, n42295, n42296, n42297, n42298,
         n42299, n42300, n42301, n42302, n42303, n42304, n42305, n42306,
         n42307, n42308, n42309, n42310, n42311, n42312, n42313, n42314,
         n42315, n42316, n42317, n42318, n42319, n42320, n42321, n42322,
         n42323, n42324, n42325, n42326, n42327, n42328, n42329, n42330,
         n42331, n42332, n42333, n42334, n42335, n42336, n42337, n42338,
         n42339, n42340, n42341, n42342, n42343, n42344, n42345, n42346,
         n42347, n42348, n42349, n42350, n42351, n42352, n42353, n42354,
         n42355, n42356, n42357, n42358, n42359, n42360, n42361, n42362,
         n42363, n42364, n42365, n42366, n42367, n42368, n42369, n42370,
         n42371, n42372, n42373, n42374, n42375, n42376, n42377, n42378,
         n42379, n42380, n42381, n42382, n42383, n42384, n42385, n42386,
         n42387, n42388, n42389, n42390, n42391, n42392, n42393, n42394,
         n42395, n42396, n42397, n42398, n42399, n42400, n42401, n42402,
         n42403, n42404, n42405, n42406, n42407, n42408, n42409, n42410,
         n42411, n42412, n42413, n42414, n42415, n42416, n42417, n42418,
         n42419, n42420, n42421, n42422, n42423, n42424, n42425, n42426,
         n42427, n42428, n42429, n42430, n42431, n42432, n42433, n42434,
         n42435, n42436, n42437, n42438, n42439, n42440, n42441, n42442,
         n42443, n42444, n42445, n42446, n42447, n42448, n42449, n42450,
         n42451, n42452, n42453, n42454, n42455, n42456, n42457, n42458,
         n42459, n42460, n42461, n42462, n42463, n42464, n42465, n42466,
         n42467, n42468, n42469, n42470, n42471, n42472, n42473, n42474,
         n42475, n42476, n42477, n42478, n42479, n42480, n42481, n42482,
         n42483, n42484, n42485, n42486, n42487, n42488, n42489, n42490,
         n42491, n42492, n42493, n42494, n42495, n42496, n42497, n42498,
         n42499, n42500, n42501, n42502, n42503, n42504, n42505, n42506,
         n42507, n42508, n42509, n42510, n42511, n42512, n42513, n42514,
         n42515, n42516, n42517, n42518, n42519, n42520, n42521, n42522,
         n42523, n42524, n42525, n42526, n42527, n42528, n42529, n42530,
         n42531, n42532, n42533, n42534, n42535, n42536, n42537, n42538,
         n42539, n42540, n42541, n42542, n42543, n42544, n42545, n42546,
         n42547, n42548, n42549, n42550, n42551, n42552, n42553, n42554,
         n42555, n42556, n42557, n42558, n42559, n42560, n42561, n42562,
         n42563, n42564, n42565, n42566, n42567, n42568, n42569, n42570,
         n42571, n42572, n42573, n42574, n42575, n42576, n42577, n42578,
         n42579, n42580, n42581, n42582, n42583, n42584, n42585, n42586,
         n42587, n42588, n42589, n42590, n42591, n42592, n42593, n42594,
         n42595, n42596, n42597, n42598, n42599, n42600, n42601, n42602,
         n42603, n42604, n42605, n42606, n42607, n42608, n42609, n42610,
         n42611, n42612, n42613, n42614, n42615, n42616, n42617, n42618,
         n42619, n42620, n42621, n42622, n42623, n42624, n42625, n42626,
         n42627, n42628, n42629, n42630, n42631, n42632, n42633, n42634,
         n42635, n42636, n42637, n42638, n42639, n42640, n42641, n42642,
         n42643, n42644, n42645, n42646, n42647, n42648, n42649, n42650,
         n42651, n42652, n42653, n42654, n42655, n42656, n42657, n42658,
         n42659, n42660, n42661, n42662, n42663, n42664, n42665, n42666,
         n42667, n42668, n42669, n42670, n42671, n42672, n42673, n42674,
         n42675, n42676, n42677, n42678, n42679, n42680, n42681, n42682,
         n42683, n42684, n42685, n42686, n42687, n42688, n42689, n42690,
         n42691, n42692, n42693, n42694, n42695, n42696, n42697, n42698,
         n42699, n42700, n42701, n42702, n42703, n42704, n42705, n42706,
         n42707, n42708, n42709, n42710, n42711, n42712, n42713, n42714,
         n42715, n42716, n42717, n42718, n42719, n42720, n42721, n42722,
         n42723, n42724, n42725, n42726, n42727, n42728, n42729, n42730,
         n42731, n42732, n42733, n42734, n42735, n42736, n42737, n42738,
         n42739, n42740, n42741, n42742, n42743, n42744, n42745, n42746,
         n42747, n42748, n42749, n42750, n42751, n42752, n42753, n42754,
         n42755, n42756, n42757, n42758, n42759, n42760, n42761, n42762,
         n42763, n42764, n42765, n42766, n42767, n42768, n42769, n42770,
         n42771, n42772, n42773, n42774, n42775, n42776, n42777, n42778,
         n42779, n42780, n42781, n42782, n42783, n42784, n42785, n42786,
         n42787, n42788, n42789, n42790, n42791, n42792, n42793, n42794,
         n42795, n42796, n42797, n42798, n42799, n42800, n42801, n42802,
         n42803, n42804, n42805, n42806, n42807, n42808, n42809, n42810,
         n42811, n42812, n42813, n42814, n42815, n42816, n42817, n42818,
         n42819, n42820, n42821, n42822, n42823, n42824, n42825, n42826,
         n42827, n42828, n42829, n42830, n42831, n42832, n42833, n42834,
         n42835, n42836, n42837, n42838, n42839, n42840, n42841, n42842,
         n42843, n42844, n42845, n42846, n42847, n42848, n42849, n42850,
         n42851, n42852, n42853, n42854, n42855, n42856, n42857, n42858,
         n42859, n42860, n42861, n42862, n42863, n42864, n42865, n42866,
         n42867, n42868, n42869, n42870, n42871, n42872, n42873, n42874,
         n42875, n42876, n42877, n42878, n42879, n42880, n42881, n42882,
         n42883, n42884, n42885, n42886, n42887, n42888, n42889, n42890,
         n42891, n42892, n42893, n42894, n42895, n42896, n42897, n42898,
         n42899, n42900, n42901, n42902, n42903, n42904, n42905, n42906,
         n42907, n42908, n42909, n42910, n42911, n42912, n42913, n42914,
         n42915, n42916, n42917, n42918, n42919, n42920, n42921, n42922,
         n42923, n42924, n42925, n42926, n42927, n42928, n42929, n42930,
         n42931, n42932, n42933, n42934, n42935, n42936, n42937, n42938,
         n42939, n42940, n42941, n42942, n42943, n42944, n42945, n42946,
         n42947, n42948, n42949, n42950, n42951, n42952, n42953, n42954,
         n42955, n42956, n42957, n42958, n42959, n42960, n42961, n42962,
         n42963, n42964, n42965, n42966, n42967, n42968, n42969, n42970,
         n42971, n42972, n42973, n42974, n42975, n42976, n42977, n42978,
         n42979, n42980, n42981, n42982, n42983, n42984, n42985, n42986,
         n42987, n42988, n42989, n42990, n42991, n42992, n42993, n42994,
         n42995, n42996, n42997, n42998, n42999, n43000, n43001, n43002,
         n43003, n43004, n43005, n43006, n43007, n43008, n43009, n43010,
         n43011, n43012, n43013, n43014, n43015, n43016, n43017, n43018,
         n43019, n43020, n43021, n43022, n43023, n43024, n43025, n43026,
         n43027, n43028, n43029, n43030, n43031, n43032, n43033, n43034,
         n43035, n43036, n43037, n43038, n43039, n43040, n43041, n43042,
         n43043, n43044, n43045, n43046, n43047, n43048, n43049, n43050,
         n43051, n43052, n43053, n43054, n43055, n43056, n43057, n43058,
         n43059, n43060, n43061, n43062, n43063, n43064, n43065, n43066,
         n43067, n43068, n43069, n43070, n43071, n43072, n43073, n43074,
         n43075, n43076, n43077, n43078, n43079, n43080, n43081, n43082,
         n43083, n43084, n43085, n43086, n43087, n43088, n43089, n43090,
         n43091, n43092, n43093, n43094, n43095, n43096, n43097, n43098,
         n43099, n43100, n43101, n43102, n43103, n43104, n43105, n43106,
         n43107, n43108, n43109, n43110, n43111, n43112, n43113, n43114,
         n43115, n43116, n43117, n43118, n43119, n43120, n43121, n43122,
         n43123, n43124, n43125, n43126, n43127, n43128, n43129, n43130,
         n43131, n43132, n43133, n43134, n43135, n43136, n43137, n43138,
         n43139, n43140, n43141, n43142, n43143, n43144, n43145, n43146,
         n43147, n43148, n43149, n43150, n43151, n43152, n43153, n43154,
         n43155, n43156, n43157, n43158, n43159, n43160, n43161, n43162,
         n43163, n43164, n43165, n43166, n43167, n43168, n43169, n43170,
         n43171, n43172, n43173, n43174, n43175, n43176, n43177, n43178,
         n43179, n43180, n43181, n43182, n43183, n43184, n43185, n43186,
         n43187, n43188, n43189, n43190, n43191, n43192, n43193, n43194,
         n43195, n43196, n43197, n43198, n43199, n43200, n43201, n43202,
         n43203, n43204, n43205, n43206, n43207, n43208, n43209, n43210,
         n43211, n43212, n43213, n43214, n43215, n43216, n43217, n43218,
         n43219, n43220, n43221, n43222, n43223, n43224, n43225, n43226,
         n43227, n43228, n43229, n43230, n43231, n43232, n43233, n43234,
         n43235, n43236, n43237, n43238, n43239, n43240, n43241, n43242,
         n43243, n43244, n43245, n43246, n43247, n43248, n43249, n43250,
         n43251, n43252, n43253, n43254, n43255, n43256, n43257, n43258,
         n43259, n43260, n43261, n43262, n43263, n43264, n43265, n43266,
         n43267, n43268, n43269, n43270, n43271, n43272, n43273, n43274,
         n43275, n43276, n43277, n43278, n43279, n43280, n43281, n43282,
         n43283, n43284, n43285, n43286, n43287, n43288, n43289, n43290,
         n43291, n43292, n43293, n43294, n43295, n43296, n43297, n43298,
         n43299, n43300, n43301, n43302, n43303, n43304, n43305, n43306,
         n43307, n43308, n43309, n43310, n43311, n43312, n43313, n43314,
         n43315, n43316, n43317, n43318, n43319, n43320, n43321, n43322,
         n43323, n43324, n43325, n43326, n43327, n43328, n43329, n43330,
         n43331, n43332, n43333, n43334, n43335, n43336, n43337, n43338,
         n43339, n43340, n43341, n43342, n43343, n43344, n43345, n43346,
         n43347, n43348, n43349, n43350, n43351, n43352, n43353, n43354,
         n43355, n43356, n43357, n43358, n43359, n43360, n43361, n43362,
         n43363, n43364, n43365, n43366, n43367, n43368, n43369, n43370,
         n43371, n43372, n43373, n43374, n43375, n43376, n43377, n43378,
         n43379, n43380, n43381, n43382, n43383, n43384, n43385, n43386,
         n43387, n43388, n43389, n43390, n43391, n43392, n43393, n43394,
         n43395, n43396, n43397, n43398, n43399, n43400, n43401, n43402,
         n43403, n43404, n43405, n43406, n43407, n43408, n43409, n43410,
         n43411, n43412, n43413, n43414, n43415, n43416, n43417, n43418,
         n43419, n43420, n43421, n43422, n43423, n43424, n43425, n43426,
         n43427, n43428, n43429, n43430, n43431, n43432, n43433, n43434,
         n43435, n43436, n43437, n43438, n43439, n43440, n43441, n43442,
         n43443, n43444, n43445, n43446, n43447, n43448, n43449, n43450,
         n43451, n43452, n43453, n43454, n43455, n43456, n43457, n43458,
         n43459, n43460, n43461, n43462, n43463, n43464, n43465, n43466,
         n43467, n43468, n43469, n43470, n43471, n43472, n43473, n43474,
         n43475, n43476, n43477, n43478, n43479, n43480, n43481, n43482,
         n43483, n43484, n43485, n43486, n43487, n43488, n43489, n43490,
         n43491, n43492, n43493, n43494, n43495, n43496, n43497, n43498,
         n43499, n43500, n43501, n43502, n43503, n43504, n43505, n43506,
         n43507, n43508, n43509, n43510, n43511, n43512, n43513, n43514,
         n43515, n43516, n43517, n43518, n43519, n43520, n43521, n43522,
         n43523, n43524, n43525, n43526, n43527, n43528, n43529, n43530,
         n43531, n43532, n43533, n43534, n43535, n43536, n43537, n43538,
         n43539, n43540, n43541, n43542, n43543, n43544, n43545, n43546,
         n43547, n43548, n43549, n43550, n43551, n43552, n43553, n43554,
         n43555, n43556, n43557, n43558, n43559, n43560, n43561, n43562,
         n43563, n43564, n43565, n43566, n43567, n43568, n43569, n43570,
         n43571, n43572, n43573, n43574, n43575, n43576, n43577, n43578,
         n43579, n43580, n43581, n43582, n43583, n43584, n43585, n43586,
         n43587, n43588, n43589, n43590, n43591, n43592, n43593, n43594,
         n43595, n43596, n43597, n43598, n43599, n43600, n43601, n43602,
         n43603, n43604, n43605, n43606, n43607, n43608, n43609, n43610,
         n43611, n43612, n43613, n43614, n43615, n43616, n43617, n43618,
         n43619, n43620, n43621, n43622, n43623, n43624, n43625, n43626,
         n43627, n43628, n43629, n43630, n43631, n43632, n43633, n43634,
         n43635, n43636, n43637, n43638, n43639, n43640, n43641, n43642,
         n43643, n43644, n43645, n43646, n43647, n43648, n43649, n43650,
         n43651, n43652, n43653, n43654, n43655, n43656, n43657, n43658,
         n43659, n43660, n43661, n43662, n43663, n43664, n43665, n43666,
         n43667, n43668, n43669, n43670, n43671, n43672, n43673, n43674,
         n43675, n43676, n43677, n43678, n43679, n43680, n43681, n43682,
         n43683, n43684, n43685, n43686, n43687, n43688, n43689, n43690,
         n43691, n43692, n43693, n43694, n43695, n43696, n43697, n43698,
         n43699, n43700, n43701, n43702, n43703, n43704, n43705, n43706,
         n43707, n43708, n43709, n43710, n43711, n43712, n43713, n43714,
         n43715, n43716, n43717, n43718, n43719, n43720, n43721, n43722,
         n43723, n43724, n43725, n43726, n43727, n43728, n43729, n43730,
         n43731, n43732, n43733, n43734, n43735, n43736, n43737, n43738,
         n43739, n43740, n43741, n43742, n43743, n43744, n43745, n43746,
         n43747, n43748, n43749, n43750, n43751, n43752, n43753, n43754,
         n43755, n43756, n43757, n43758, n43759, n43760, n43761, n43762,
         n43763, n43764, n43765, n43766, n43767, n43768, n43769, n43770,
         n43771, n43772, n43773, n43774, n43775, n43776, n43777, n43778,
         n43779, n43780, n43781, n43782, n43783, n43784, n43785, n43786,
         n43787, n43788, n43789, n43790, n43791, n43792, n43793, n43794,
         n43795, n43796, n43797, n43798, n43799, n43800, n43801, n43802,
         n43803, n43804, n43805, n43806, n43807, n43808, n43809, n43810,
         n43811, n43812, n43813, n43814, n43815, n43816, n43817, n43818,
         n43819, n43820, n43821, n43822, n43823, n43824, n43825, n43826,
         n43827, n43828, n43829, n43830, n43831, n43832, n43833, n43834,
         n43835, n43836, n43837, n43838, n43839, n43840, n43841, n43842,
         n43843, n43844, n43845, n43846, n43847, n43848, n43849, n43850,
         n43851, n43852, n43853, n43854, n43855, n43856, n43857, n43858,
         n43859, n43860, n43861, n43862, n43863, n43864, n43865, n43866,
         n43867, n43868, n43869, n43870, n43871, n43872, n43873, n43874,
         n43875, n43876, n43877, n43878, n43879, n43880, n43881, n43882,
         n43883, n43884, n43885, n43886, n43887, n43888, n43889, n43890,
         n43891, n43892, n43893, n43894, n43895, n43896, n43897, n43898,
         n43899, n43900, n43901, n43902, n43903, n43904, n43905, n43906,
         n43907, n43908, n43909, n43910, n43911, n43912, n43913, n43914,
         n43915, n43916, n43917, n43918, n43919, n43920, n43921, n43922,
         n43923, n43924, n43925, n43926, n43927, n43928, n43929, n43930,
         n43931, n43932, n43933, n43934, n43935, n43936, n43937, n43938,
         n43939, n43940, n43941, n43942, n43943, n43944, n43945, n43946,
         n43947, n43948, n43949, n43950, n43951, n43952, n43953, n43954,
         n43955, n43956, n43957, n43958, n43959, n43960, n43961, n43962,
         n43963, n43964, n43965, n43966, n43967, n43968, n43969, n43970,
         n43971, n43972, n43973, n43974, n43975, n43976, n43977, n43978,
         n43979, n43980, n43981, n43982, n43983, n43984, n43985, n43986,
         n43987, n43988, n43989, n43990, n43991, n43992, n43993, n43994,
         n43995, n43996, n43997, n43998, n43999, n44000, n44001, n44002,
         n44003, n44004, n44005, n44006, n44007, n44008, n44009, n44010,
         n44011, n44012, n44013, n44014, n44015, n44016, n44017, n44018,
         n44019, n44020, n44021, n44022, n44023, n44024, n44025, n44026,
         n44027, n44028, n44029, n44030, n44031, n44032, n44033, n44034,
         n44035, n44036, n44037, n44038, n44039, n44040, n44041, n44042,
         n44043, n44044, n44045, n44046, n44047, n44048, n44049, n44050,
         n44051, n44052, n44053, n44054, n44055, n44056, n44057, n44058,
         n44059, n44060, n44061, n44062, n44063, n44064, n44065, n44066,
         n44067, n44068, n44069, n44070, n44071, n44072, n44073, n44074,
         n44075, n44076, n44077, n44078, n44079, n44080, n44081, n44082,
         n44083, n44084, n44085, n44086, n44087, n44088, n44089, n44090,
         n44091, n44092, n44093, n44094, n44095, n44096, n44097, n44098,
         n44099, n44100, n44101, n44102, n44103, n44104, n44105, n44106,
         n44107, n44108, n44109, n44110, n44111, n44112, n44113, n44114,
         n44115, n44116, n44117, n44118, n44119, n44120, n44121, n44122,
         n44123, n44124, n44125, n44126, n44127, n44128, n44129, n44130,
         n44131, n44132, n44133, n44134, n44135, n44136, n44137, n44138,
         n44139, n44140, n44141, n44142, n44143, n44144, n44145, n44146,
         n44147, n44148, n44149, n44150, n44151, n44152, n44153, n44154,
         n44155, n44156, n44157, n44158, n44159, n44160, n44161, n44162,
         n44163, n44164, n44165, n44166, n44167, n44168, n44169, n44170,
         n44171, n44172, n44173, n44174, n44175, n44176, n44177, n44178,
         n44179, n44180, n44181, n44182, n44183, n44184, n44185, n44186,
         n44187, n44188, n44189, n44190, n44191, n44192, n44193, n44194,
         n44195, n44196, n44197, n44198, n44199, n44200, n44201, n44202,
         n44203, n44204, n44205, n44206, n44207, n44208, n44209, n44210,
         n44211, n44212, n44213, n44214, n44215, n44216, n44217, n44218,
         n44219, n44220, n44221, n44222, n44223, n44224, n44225, n44226,
         n44227, n44228, n44229, n44230, n44231, n44232, n44233, n44234,
         n44235, n44236, n44237, n44238, n44239, n44240, n44241, n44242,
         n44243, n44244, n44245, n44246, n44247, n44248, n44249, n44250,
         n44251, n44252, n44253, n44254, n44255, n44256, n44257, n44258,
         n44259, n44260, n44261, n44262, n44263, n44264, n44265, n44266,
         n44267, n44268, n44269, n44270, n44271, n44272, n44273, n44274,
         n44275, n44276, n44277, n44278, n44279, n44280, n44281, n44282,
         n44283, n44284, n44285, n44286, n44287, n44288, n44289, n44290,
         n44291, n44292, n44293, n44294, n44295, n44296, n44297, n44298,
         n44299, n44300, n44301, n44302, n44303, n44304, n44305, n44306,
         n44307, n44308, n44309, n44310, n44311, n44312, n44313, n44314,
         n44315, n44316, n44317, n44318, n44319, n44320, n44321, n44322,
         n44323, n44324, n44325, n44326, n44327, n44328, n44329, n44330,
         n44331, n44332, n44333, n44334, n44335, n44336, n44337, n44338,
         n44339, n44340, n44341, n44342, n44343, n44344, n44345, n44346,
         n44347, n44348, n44349, n44350, n44351, n44352, n44353, n44354,
         n44355, n44356, n44357, n44358, n44359, n44360, n44361, n44362,
         n44363, n44364, n44365, n44366, n44367, n44368, n44369, n44370,
         n44371, n44372, n44373, n44374, n44375, n44376, n44377, n44378,
         n44379, n44380, n44381, n44382, n44383, n44384, n44385, n44386,
         n44387, n44388, n44389, n44390, n44391, n44392, n44393, n44394,
         n44395, n44396, n44397, n44398, n44399, n44400, n44401, n44402,
         n44403, n44404, n44405, n44406, n44407, n44408, n44409, n44410,
         n44411, n44412, n44413, n44414, n44415, n44416, n44417, n44418,
         n44419, n44420, n44421, n44422, n44423, n44424, n44425, n44426,
         n44427, n44428, n44429, n44430, n44431, n44432, n44433, n44434,
         n44435, n44436, n44437, n44438, n44439, n44440, n44441, n44442,
         n44443, n44444, n44445, n44446, n44447, n44448, n44449, n44450,
         n44451, n44452, n44453, n44454, n44455, n44456, n44457, n44458,
         n44459, n44460, n44461, n44462, n44463, n44464, n44465, n44466,
         n44467, n44468, n44469, n44470, n44471, n44472, n44473, n44474,
         n44475, n44476, n44477, n44478, n44479, n44480, n44481, n44482,
         n44483, n44484, n44485, n44486, n44487, n44488, n44489, n44490,
         n44491, n44492, n44493, n44494, n44495, n44496, n44497, n44498,
         n44499, n44500, n44501, n44502, n44503, n44504, n44505, n44506,
         n44507, n44508, n44509, n44510, n44511, n44512, n44513, n44514,
         n44515, n44516, n44517, n44518, n44519, n44520, n44521, n44522,
         n44523, n44524, n44525, n44526, n44527, n44528, n44529, n44530,
         n44531, n44532, n44533, n44534, n44535, n44536, n44537, n44538,
         n44539, n44540, n44541, n44542, n44543, n44544, n44545, n44546,
         n44547, n44548, n44549, n44550, n44551, n44552, n44553, n44554,
         n44555, n44556, n44557, n44558, n44559, n44560, n44561, n44562,
         n44563, n44564, n44565, n44566, n44567, n44568, n44569, n44570,
         n44571, n44572, n44573, n44574, n44575, n44576, n44577, n44578,
         n44579, n44580, n44581, n44582, n44583, n44584, n44585, n44586,
         n44587, n44588, n44589, n44590, n44591, n44592, n44593, n44594,
         n44595, n44596, n44597, n44598, n44599, n44600, n44601, n44602,
         n44603, n44604, n44605, n44606, n44607, n44608, n44609, n44610,
         n44611, n44612, n44613, n44614, n44615, n44616, n44617, n44618,
         n44619, n44620, n44621, n44622, n44623, n44624, n44625, n44626,
         n44627, n44628, n44629, n44630, n44631, n44632, n44633, n44634,
         n44635, n44636, n44637, n44638, n44639, n44640, n44641, n44642,
         n44643, n44644, n44645, n44646, n44647, n44648, n44649, n44650,
         n44651, n44652, n44653, n44654, n44655, n44656, n44657, n44658,
         n44659, n44660, n44661, n44662, n44663, n44664, n44665, n44666,
         n44667, n44668, n44669, n44670, n44671, n44672, n44673, n44674,
         n44675, n44676, n44677, n44678, n44679, n44680, n44681, n44682,
         n44683, n44684, n44685, n44686, n44687, n44688, n44689, n44690,
         n44691, n44692, n44693, n44694, n44695, n44696, n44697, n44698,
         n44699, n44700, n44701, n44702, n44703, n44704, n44705, n44706,
         n44707, n44708, n44709, n44710, n44711, n44712, n44713, n44714,
         n44715, n44716, n44717, n44718, n44719, n44720, n44721, n44722,
         n44723, n44724, n44725, n44726, n44727, n44728, n44729, n44730,
         n44731, n44732, n44733, n44734, n44735, n44736, n44737, n44738,
         n44739, n44740, n44741, n44742, n44743, n44744, n44745, n44746,
         n44747, n44748, n44749, n44750, n44751, n44752, n44753, n44754,
         n44755, n44756, n44757, n44758, n44759, n44760, n44761, n44762,
         n44763, n44764, n44765, n44766, n44767, n44768, n44769, n44770,
         n44771, n44772, n44773, n44774, n44775, n44776, n44777, n44778,
         n44779, n44780, n44781, n44782, n44783, n44784, n44785, n44786,
         n44787, n44788, n44789, n44790, n44791, n44792, n44793, n44794,
         n44795, n44796, n44797, n44798, n44799, n44800, n44801, n44802,
         n44803, n44804, n44805, n44806, n44807, n44808, n44809, n44810,
         n44811, n44812, n44813, n44814, n44815, n44816, n44817, n44818,
         n44819, n44820, n44821, n44822, n44823, n44824, n44825, n44826,
         n44827, n44828, n44829, n44830, n44831, n44832, n44833, n44834,
         n44835, n44836, n44837, n44838, n44839, n44840, n44841, n44842,
         n44843, n44844, n44845, n44846, n44847, n44848, n44849, n44850,
         n44851, n44852, n44853, n44854, n44855, n44856, n44857, n44858,
         n44859, n44860, n44861, n44862, n44863, n44864, n44865, n44866,
         n44867, n44868, n44869, n44870, n44871, n44872, n44873, n44874,
         n44875, n44876, n44877, n44878, n44879, n44880, n44881, n44882,
         n44883, n44884, n44885, n44886, n44887, n44888, n44889, n44890,
         n44891, n44892, n44893, n44894, n44895, n44896, n44897, n44898,
         n44899, n44900, n44901, n44902, n44903, n44904, n44905, n44906,
         n44907, n44908, n44909, n44910, n44911, n44912, n44913, n44914,
         n44915, n44916, n44917, n44918, n44919, n44920, n44921, n44922,
         n44923, n44924, n44925, n44926, n44927, n44928, n44929, n44930,
         n44931, n44932, n44933, n44934, n44935, n44936, n44937, n44938,
         n44939, n44940, n44941, n44942, n44943, n44944, n44945, n44946,
         n44947, n44948, n44949, n44950, n44951, n44952, n44953, n44954,
         n44955, n44956, n44957, n44958, n44959, n44960, n44961, n44962,
         n44963, n44964, n44965, n44966, n44967, n44968, n44969, n44970,
         n44971, n44972, n44973, n44974, n44975, n44976, n44977, n44978,
         n44979, n44980, n44981, n44982, n44983, n44984, n44985, n44986,
         n44987, n44988, n44989, n44990, n44991, n44992, n44993, n44994,
         n44995, n44996, n44997, n44998, n44999, n45000, n45001, n45002,
         n45003, n45004, n45005, n45006, n45007, n45008, n45009, n45010,
         n45011, n45012, n45013, n45014, n45015, n45016, n45017, n45018,
         n45019, n45020, n45021, n45022, n45023, n45024, n45025, n45026,
         n45027, n45028, n45029, n45030, n45031, n45032, n45033, n45034,
         n45035, n45036, n45037, n45038, n45039, n45040, n45041, n45042,
         n45043, n45044, n45045, n45046, n45047, n45048, n45049, n45050,
         n45051, n45052, n45053, n45054, n45055, n45056, n45057, n45058,
         n45059, n45060, n45061, n45062, n45063, n45064, n45065, n45066,
         n45067, n45068, n45069, n45070, n45071, n45072, n45073, n45074,
         n45075, n45076, n45077, n45078, n45079, n45080, n45081, n45082,
         n45083, n45084, n45085, n45086, n45087, n45088, n45089, n45090,
         n45091, n45092, n45093, n45094, n45095, n45096, n45097, n45098,
         n45099, n45100, n45101, n45102, n45103, n45104, n45105, n45106,
         n45107, n45108, n45109, n45110, n45111, n45112, n45113, n45114,
         n45115, n45116, n45117, n45118, n45119, n45120, n45121, n45122,
         n45123, n45124, n45125, n45126, n45127, n45128, n45129, n45130,
         n45131, n45132, n45133, n45134, n45135, n45136, n45137, n45138,
         n45139, n45140, n45141, n45142, n45143, n45144, n45145, n45146,
         n45147, n45148, n45149, n45150, n45151, n45152, n45153, n45154,
         n45155, n45156, n45157, n45158, n45159, n45160, n45161, n45162,
         n45163, n45164, n45165, n45166, n45167, n45168, n45169, n45170,
         n45171, n45172, n45173, n45174, n45175, n45176, n45177, n45178,
         n45179, n45180, n45181, n45182, n45183, n45184, n45185, n45186,
         n45187, n45188, n45189, n45190, n45191, n45192, n45193, n45194,
         n45195, n45196, n45197, n45198, n45199, n45200, n45201, n45202,
         n45203, n45204, n45205, n45206, n45207, n45208, n45209, n45210,
         n45211, n45212, n45213, n45214, n45215, n45216, n45217, n45218,
         n45219, n45220, n45221, n45222, n45223, n45224, n45225, n45226,
         n45227, n45228, n45229, n45230, n45231, n45232, n45233, n45234,
         n45235, n45236, n45237, n45238, n45239, n45240, n45241, n45242,
         n45243, n45244, n45245, n45246, n45247, n45248, n45249, n45250,
         n45251, n45252, n45253, n45254, n45255, n45256, n45257, n45258,
         n45259, n45260, n45261, n45262, n45263, n45264, n45265, n45266,
         n45267, n45268, n45269, n45270, n45271, n45272, n45273, n45274,
         n45275, n45276, n45277, n45278, n45279, n45280, n45281, n45282,
         n45283, n45284, n45285, n45286, n45287, n45288, n45289, n45290,
         n45291, n45292, n45293, n45294, n45295, n45296, n45297, n45298,
         n45299, n45300, n45301, n45302, n45303, n45304, n45305, n45306,
         n45307, n45308, n45309, n45310, n45311, n45312, n45313, n45314,
         n45315, n45316, n45317, n45318, n45319, n45320, n45321, n45322,
         n45323, n45324, n45325, n45326, n45327, n45328, n45329, n45330,
         n45331, n45332, n45333, n45334, n45335, n45336, n45337, n45338,
         n45339, n45340, n45341, n45342, n45343, n45344, n45345, n45346,
         n45347, n45348, n45349, n45350, n45351, n45352, n45353, n45354,
         n45355, n45356, n45357, n45358, n45359, n45360, n45361, n45362,
         n45363, n45364, n45365, n45366, n45367, n45368, n45369, n45370,
         n45371, n45372, n45373, n45374, n45375, n45376, n45377, n45378,
         n45379, n45380, n45381, n45382, n45383, n45384, n45385, n45386,
         n45387, n45388, n45389, n45390, n45391, n45392, n45393, n45394,
         n45395, n45396, n45397, n45398, n45399, n45400, n45401, n45402,
         n45403, n45404, n45405, n45406, n45407, n45408, n45409, n45410,
         n45411, n45412, n45413, n45414, n45415, n45416, n45417, n45418,
         n45419, n45420, n45421, n45422, n45423, n45424, n45425, n45426,
         n45427, n45428, n45429, n45430, n45431, n45432, n45433, n45434,
         n45435, n45436, n45437, n45438, n45439, n45440, n45441, n45442,
         n45443, n45444, n45445, n45446, n45447, n45448, n45449, n45450,
         n45451, n45452, n45453, n45454, n45455, n45456, n45457, n45458,
         n45459, n45460, n45461, n45462, n45463, n45464, n45465, n45466,
         n45467, n45468, n45469, n45470, n45471, n45472, n45473, n45474,
         n45475, n45476, n45477, n45478, n45479, n45480, n45481, n45482,
         n45483, n45484, n45485, n45486, n45487, n45488, n45489, n45490,
         n45491, n45492, n45493, n45494, n45495, n45496, n45497, n45498,
         n45499, n45500, n45501, n45502, n45503, n45504, n45505, n45506,
         n45507, n45508, n45509, n45510, n45511, n45512, n45513, n45514,
         n45515, n45516, n45517, n45518, n45519, n45520, n45521, n45522,
         n45523, n45524, n45525, n45526, n45527, n45528, n45529, n45530,
         n45531, n45532, n45533, n45534, n45535, n45536, n45537, n45538,
         n45539, n45540, n45541, n45542, n45543, n45544, n45545, n45546,
         n45547, n45548, n45549, n45550, n45551, n45552, n45553, n45554,
         n45555, n45556, n45557, n45558, n45559, n45560, n45561, n45562,
         n45563, n45564, n45565, n45566, n45567, n45568, n45569, n45570,
         n45571, n45572, n45573, n45574, n45575, n45576, n45577, n45578,
         n45579, n45580, n45581, n45582, n45583, n45584, n45585, n45586,
         n45587, n45588, n45589, n45590, n45591, n45592, n45593, n45594,
         n45595, n45596, n45597, n45598, n45599, n45600, n45601, n45602,
         n45603, n45604, n45605, n45606, n45607, n45608, n45609, n45610,
         n45611, n45612, n45613, n45614, n45615, n45616, n45617, n45618,
         n45619, n45620, n45621, n45622, n45623, n45624, n45625, n45626,
         n45627, n45628, n45629, n45630, n45631, n45632, n45633, n45634,
         n45635, n45636, n45637, n45638, n45639, n45640, n45641, n45642,
         n45643, n45644, n45645, n45646, n45647, n45648, n45649, n45650,
         n45651, n45652, n45653, n45654, n45655, n45656, n45657, n45658,
         n45659, n45660, n45661, n45662, n45663, n45664, n45665, n45666,
         n45667, n45668, n45669, n45670, n45671, n45672, n45673, n45674,
         n45675, n45676, n45677, n45678, n45679, n45680, n45681, n45682,
         n45683, n45684, n45685, n45686, n45687, n45688, n45689, n45690,
         n45691, n45692, n45693, n45694, n45695, n45696, n45697, n45698,
         n45699, n45700, n45701, n45702, n45703, n45704, n45705, n45706,
         n45707, n45708, n45709, n45710, n45711, n45712, n45713, n45714,
         n45715, n45716, n45717, n45718, n45719, n45720, n45721, n45722,
         n45723, n45724, n45725, n45726, n45727, n45728, n45729, n45730,
         n45731, n45732, n45733, n45734, n45735, n45736, n45737, n45738,
         n45739, n45740, n45741, n45742, n45743, n45744, n45745, n45746,
         n45747, n45748, n45749, n45750, n45751, n45752, n45753, n45754,
         n45755, n45756, n45757, n45758, n45759, n45760, n45761, n45762,
         n45763, n45764, n45765, n45766, n45767, n45768, n45769, n45770,
         n45771, n45772, n45773, n45774, n45775, n45776, n45777, n45778,
         n45779, n45780, n45781, n45782, n45783, n45784, n45785, n45786,
         n45787, n45788, n45789, n45790, n45791, n45792, n45793, n45794,
         n45795, n45796, n45797, n45798, n45799, n45800, n45801, n45802,
         n45803, n45804, n45805, n45806, n45807, n45808, n45809, n45810,
         n45811, n45812, n45813, n45814, n45815, n45816, n45817, n45818,
         n45819, n45820, n45821, n45822, n45823, n45824, n45825, n45826,
         n45827, n45828, n45829, n45830, n45831, n45832, n45833, n45834,
         n45835, n45836, n45837, n45838, n45839, n45840, n45841, n45842,
         n45843, n45844, n45845, n45846, n45847, n45848, n45849, n45850,
         n45851, n45852, n45853, n45854, n45855, n45856, n45857, n45858,
         n45859, n45860, n45861, n45862, n45863, n45864, n45865, n45866,
         n45867, n45868, n45869, n45870, n45871, n45872, n45873, n45874,
         n45875, n45876, n45877, n45878, n45879, n45880, n45881, n45882,
         n45883, n45884, n45885, n45886, n45887, n45888, n45889, n45890,
         n45891, n45892, n45893, n45894, n45895, n45896, n45897, n45898,
         n45899, n45900, n45901, n45902, n45903, n45904, n45905, n45906,
         n45907, n45908, n45909, n45910, n45911, n45912, n45913, n45914,
         n45915, n45916, n45917, n45918, n45919, n45920, n45921, n45922,
         n45923, n45924, n45925, n45926, n45927, n45928, n45929, n45930,
         n45931, n45932, n45933, n45934, n45935, n45936, n45937, n45938,
         n45939, n45940, n45941, n45942, n45943, n45944, n45945, n45946,
         n45947, n45948, n45949, n45950, n45951, n45952, n45953, n45954,
         n45955, n45956, n45957, n45958, n45959, n45960, n45961, n45962,
         n45963, n45964, n45965, n45966, n45967, n45968, n45969, n45970,
         n45971, n45972, n45973, n45974, n45975, n45976, n45977, n45978,
         n45979, n45980, n45981, n45982, n45983, n45984, n45985, n45986,
         n45987, n45988, n45989, n45990, n45991, n45992, n45993, n45994,
         n45995, n45996, n45997, n45998, n45999, n46000, n46001, n46002,
         n46003, n46004, n46005, n46006, n46007, n46008, n46009, n46010,
         n46011, n46012, n46013, n46014, n46015, n46016, n46017, n46018,
         n46019, n46020, n46021, n46022, n46023, n46024, n46025, n46026,
         n46027, n46028, n46029, n46030, n46031, n46032, n46033, n46034,
         n46035, n46036, n46037, n46038, n46039, n46040, n46041, n46042,
         n46043, n46044, n46045, n46046, n46047, n46048, n46049, n46050,
         n46051, n46052, n46053, n46054, n46055, n46056, n46057, n46058,
         n46059, n46060, n46061, n46062, n46063, n46064, n46065, n46066,
         n46067, n46068, n46069, n46070, n46071, n46072, n46073, n46074,
         n46075, n46076, n46077, n46078, n46079, n46080, n46081, n46082,
         n46083, n46084, n46085, n46086, n46087, n46088, n46089, n46090,
         n46091, n46092, n46093, n46094, n46095, n46096, n46097, n46098,
         n46099, n46100, n46101, n46102, n46103, n46104, n46105, n46106,
         n46107, n46108, n46109, n46110, n46111, n46112, n46113, n46114,
         n46115, n46116, n46117, n46118, n46119, n46120, n46121, n46122,
         n46123, n46124, n46125, n46126, n46127, n46128, n46129, n46130,
         n46131, n46132, n46133, n46134, n46135, n46136, n46137, n46138,
         n46139, n46140, n46141, n46142, n46143, n46144, n46145, n46146,
         n46147, n46148, n46149, n46150, n46151, n46152, n46153, n46154,
         n46155, n46156, n46157, n46158, n46159, n46160, n46161, n46162,
         n46163, n46164, n46165, n46166, n46167, n46168, n46169, n46170,
         n46171, n46172, n46173, n46174, n46175, n46176, n46177, n46178,
         n46179, n46180, n46181, n46182, n46183, n46184, n46185, n46186,
         n46187, n46188, n46189, n46190, n46191, n46192, n46193, n46194,
         n46195, n46196, n46197, n46198, n46199, n46200, n46201, n46202,
         n46203, n46204, n46205, n46206, n46207, n46208, n46209, n46210,
         n46211, n46212, n46213, n46214, n46215, n46216, n46217, n46218,
         n46219, n46220, n46221, n46222, n46223, n46224, n46225, n46226,
         n46227, n46228, n46229, n46230, n46231, n46232, n46233, n46234,
         n46235, n46236, n46237, n46238, n46239, n46240, n46241, n46242,
         n46243, n46244, n46245, n46246, n46247, n46248, n46249, n46250,
         n46251, n46252, n46253, n46254, n46255, n46256, n46257, n46258,
         n46259, n46260, n46261, n46262, n46263, n46264, n46265, n46266,
         n46267, n46268, n46269, n46270, n46271, n46272, n46273, n46274,
         n46275, n46276, n46277, n46278, n46279, n46280, n46281, n46282,
         n46283, n46284, n46285, n46286, n46287, n46288, n46289, n46290,
         n46291, n46292, n46293, n46294, n46295, n46296, n46297, n46298,
         n46299, n46300, n46301, n46302, n46303, n46304, n46305, n46306,
         n46307, n46308, n46309, n46310, n46311, n46312, n46313, n46314,
         n46315, n46316, n46317, n46318, n46319, n46320, n46321, n46322,
         n46323, n46324, n46325, n46326, n46327, n46328, n46329, n46330,
         n46331, n46332, n46333, n46334, n46335, n46336, n46337, n46338,
         n46339, n46340, n46341, n46342, n46343, n46344, n46345, n46346,
         n46347, n46348, n46349, n46350, n46351, n46352, n46353, n46354,
         n46355, n46356, n46357, n46358, n46359, n46360, n46361, n46362,
         n46363, n46364, n46365, n46366, n46367, n46368, n46369, n46370,
         n46371, n46372, n46373, n46374, n46375, n46376, n46377, n46378,
         n46379, n46380, n46381, n46382, n46383, n46384, n46385, n46386,
         n46387, n46388, n46389, n46390, n46391, n46392, n46393, n46394,
         n46395, n46396, n46397, n46398, n46399, n46400, n46401, n46402,
         n46403, n46404, n46405, n46406, n46407, n46408, n46409, n46410,
         n46411, n46412, n46413, n46414, n46415, n46416, n46417, n46418,
         n46419, n46420, n46421, n46422, n46423, n46424, n46425, n46426,
         n46427, n46428, n46429, n46430, n46431, n46432, n46433, n46434,
         n46435, n46436, n46437, n46438, n46439, n46440, n46441, n46442,
         n46443, n46444, n46445, n46446, n46447, n46448, n46449, n46450,
         n46451, n46452, n46453, n46454, n46455, n46456, n46457, n46458,
         n46459, n46460, n46461, n46462, n46463, n46464, n46465, n46466,
         n46467, n46468, n46469, n46470, n46471, n46472, n46473, n46474,
         n46475, n46476, n46477, n46478, n46479, n46480, n46481, n46482,
         n46483, n46484, n46485, n46486, n46487, n46488, n46489, n46490,
         n46491, n46492, n46493, n46494, n46495, n46496, n46497, n46498,
         n46499, n46500, n46501, n46502, n46503, n46504, n46505, n46506,
         n46507, n46508, n46509, n46510, n46511, n46512, n46513, n46514,
         n46515, n46516, n46517, n46518, n46519, n46520, n46521, n46522,
         n46523, n46524, n46525, n46526, n46527, n46528, n46529, n46530,
         n46531, n46532, n46533, n46534, n46535, n46536, n46537, n46538,
         n46539, n46540, n46541, n46542, n46543, n46544, n46545, n46546,
         n46547, n46548, n46549, n46550, n46551, n46552, n46553, n46554,
         n46555, n46556, n46557, n46558, n46559, n46560, n46561, n46562,
         n46563, n46564, n46565, n46566, n46567, n46568, n46569, n46570,
         n46571, n46572, n46573, n46574, n46575, n46576, n46577, n46578,
         n46579, n46580, n46581, n46582, n46583, n46584, n46585, n46586,
         n46587, n46588, n46589, n46590, n46591, n46592, n46593, n46594,
         n46595, n46596, n46597, n46598, n46599, n46600, n46601, n46602,
         n46603, n46604, n46605, n46606, n46607, n46608, n46609, n46610,
         n46611, n46612, n46613, n46614, n46615, n46616, n46617, n46618,
         n46619, n46620, n46621, n46622, n46623, n46624, n46625, n46626,
         n46627, n46628, n46629, n46630, n46631, n46632, n46633, n46634,
         n46635, n46636, n46637, n46638, n46639, n46640, n46641, n46642,
         n46643, n46644, n46645, n46646, n46647, n46648, n46649, n46650,
         n46651, n46652, n46653, n46654, n46655, n46656, n46657, n46658,
         n46659, n46660, n46661, n46662, n46663, n46664, n46665, n46666,
         n46667, n46668, n46669, n46670, n46671, n46672, n46673, n46674,
         n46675, n46676, n46677, n46678, n46679, n46680, n46681, n46682,
         n46683, n46684, n46685, n46686, n46687, n46688, n46689, n46690,
         n46691, n46692, n46693, n46694, n46695, n46696, n46697, n46698,
         n46699, n46700, n46701, n46702, n46703, n46704, n46705, n46706,
         n46707, n46708, n46709, n46710, n46711, n46712, n46713, n46714,
         n46715, n46716, n46717, n46718, n46719, n46720, n46721, n46722,
         n46723, n46724, n46725, n46726, n46727, n46728, n46729, n46730,
         n46731, n46732, n46733, n46734, n46735, n46736, n46737, n46738,
         n46739, n46740, n46741, n46742, n46743, n46744, n46745, n46746,
         n46747, n46748, n46749, n46750, n46751, n46752, n46753, n46754,
         n46755, n46756, n46757, n46758, n46759, n46760, n46761, n46762,
         n46763, n46764, n46765, n46766, n46767, n46768, n46769, n46770,
         n46771, n46772, n46773, n46774, n46775, n46776, n46777, n46778,
         n46779, n46780, n46781, n46782, n46783, n46784, n46785, n46786,
         n46787, n46788, n46789, n46790, n46791, n46792, n46793, n46794,
         n46795, n46796, n46797, n46798, n46799, n46800, n46801, n46802,
         n46803, n46804, n46805, n46806, n46807, n46808, n46809, n46810,
         n46811, n46812, n46813, n46814, n46815, n46816, n46817, n46818,
         n46819, n46820, n46821, n46822, n46823, n46824, n46825, n46826,
         n46827, n46828, n46829, n46830, n46831, n46832, n46833, n46834,
         n46835, n46836, n46837, n46838, n46839, n46840, n46841, n46842,
         n46843, n46844, n46845, n46846, n46847, n46848, n46849, n46850,
         n46851, n46852, n46853, n46854, n46855, n46856, n46857, n46858,
         n46859, n46860, n46861, n46862, n46863, n46864, n46865, n46866,
         n46867, n46868, n46869, n46870, n46871, n46872, n46873, n46874,
         n46875, n46876, n46877, n46878, n46879, n46880, n46881, n46882,
         n46883, n46884, n46885, n46886, n46887, n46888, n46889, n46890,
         n46891, n46892, n46893, n46894, n46895, n46896, n46897, n46898,
         n46899, n46900, n46901, n46902, n46903, n46904, n46905, n46906,
         n46907, n46908, n46909, n46910, n46911, n46912, n46913, n46914,
         n46915, n46916, n46917, n46918, n46919, n46920, n46921, n46922,
         n46923, n46924, n46925, n46926, n46927, n46928, n46929, n46930,
         n46931, n46932, n46933, n46934, n46935, n46936, n46937, n46938,
         n46939, n46940, n46941, n46942, n46943, n46944, n46945, n46946,
         n46947, n46948, n46949, n46950, n46951, n46952, n46953, n46954,
         n46955, n46956, n46957, n46958, n46959, n46960, n46961, n46962,
         n46963, n46964, n46965, n46966, n46967, n46968, n46969, n46970,
         n46971, n46972, n46973, n46974, n46975, n46976, n46977, n46978,
         n46979, n46980, n46981, n46982, n46983, n46984, n46985, n46986,
         n46987, n46988, n46989, n46990, n46991, n46992, n46993, n46994,
         n46995, n46996, n46997, n46998, n46999, n47000, n47001, n47002,
         n47003, n47004, n47005, n47006, n47007, n47008, n47009, n47010,
         n47011, n47012, n47013, n47014, n47015, n47016, n47017, n47018,
         n47019, n47020, n47021, n47022, n47023, n47024, n47025, n47026,
         n47027, n47028, n47029, n47030, n47031, n47032, n47033, n47034,
         n47035, n47036, n47037, n47038, n47039, n47040, n47041, n47042,
         n47043, n47044, n47045, n47046, n47047, n47048, n47049, n47050,
         n47051, n47052, n47053, n47054, n47055, n47056, n47057, n47058,
         n47059, n47060, n47061, n47062, n47063, n47064, n47065, n47066,
         n47067, n47068, n47069, n47070, n47071, n47072, n47073, n47074,
         n47075, n47076, n47077, n47078, n47079, n47080, n47081, n47082,
         n47083, n47084, n47085, n47086, n47087, n47088, n47089, n47090,
         n47091, n47092, n47093, n47094, n47095, n47096, n47097, n47098,
         n47099, n47100, n47101, n47102, n47103, n47104, n47105, n47106,
         n47107, n47108, n47109, n47110, n47111, n47112, n47113, n47114,
         n47115, n47116, n47117, n47118, n47119, n47120, n47121, n47122,
         n47123, n47124, n47125, n47126, n47127, n47128, n47129, n47130,
         n47131, n47132, n47133, n47134, n47135, n47136, n47137, n47138,
         n47139, n47140, n47141, n47142, n47143, n47144, n47145, n47146,
         n47147, n47148, n47149, n47150, n47151, n47152, n47153, n47154,
         n47155, n47156, n47157, n47158, n47159, n47160, n47161, n47162,
         n47163, n47164, n47165, n47166, n47167, n47168, n47169, n47170,
         n47171, n47172, n47173, n47174, n47175, n47176, n47177, n47178,
         n47179, n47180, n47181, n47182, n47183, n47184, n47185, n47186,
         n47187, n47188, n47189, n47190, n47191, n47192, n47193, n47194,
         n47195, n47196, n47197, n47198, n47199, n47200, n47201, n47202,
         n47203, n47204, n47205, n47206, n47207, n47208, n47209, n47210,
         n47211, n47212, n47213, n47214, n47215, n47216, n47217, n47218,
         n47219, n47220, n47221, n47222, n47223, n47224, n47225, n47226,
         n47227, n47228, n47229, n47230, n47231, n47232, n47233, n47234,
         n47235, n47236, n47237, n47238, n47239, n47240, n47241, n47242,
         n47243, n47244, n47245, n47246, n47247, n47248, n47249, n47250,
         n47251, n47252, n47253, n47254, n47255, n47256, n47257, n47258,
         n47259, n47260, n47261, n47262, n47263, n47264, n47265, n47266,
         n47267, n47268, n47269, n47270, n47271, n47272, n47273, n47274,
         n47275, n47276, n47277, n47278, n47279, n47280, n47281, n47282,
         n47283, n47284, n47285, n47286, n47287, n47288, n47289, n47290,
         n47291, n47292, n47293, n47294, n47295, n47296, n47297, n47298,
         n47299, n47300, n47301, n47302, n47303, n47304, n47305, n47306,
         n47307, n47308, n47309, n47310, n47311, n47312, n47313, n47314,
         n47315, n47316, n47317, n47318, n47319, n47320, n47321, n47322,
         n47323, n47324, n47325, n47326, n47327, n47328, n47329, n47330,
         n47331, n47332, n47333, n47334, n47335, n47336, n47337, n47338,
         n47339, n47340, n47341, n47342, n47343, n47344, n47345, n47346,
         n47347, n47348, n47349, n47350, n47351, n47352, n47353, n47354,
         n47355, n47356, n47357, n47358, n47359, n47360, n47361, n47362,
         n47363, n47364, n47365, n47366, n47367, n47368, n47369, n47370,
         n47371, n47372, n47373, n47374, n47375, n47376, n47377, n47378,
         n47379, n47380, n47381, n47382, n47383, n47384, n47385, n47386,
         n47387, n47388, n47389, n47390, n47391, n47392, n47393, n47394,
         n47395, n47396, n47397, n47398, n47399, n47400, n47401, n47402,
         n47403, n47404, n47405, n47406, n47407, n47408, n47409, n47410,
         n47411, n47412, n47413, n47414, n47415, n47416, n47417, n47418,
         n47419, n47420, n47421, n47422, n47423, n47424, n47425, n47426,
         n47427, n47428, n47429, n47430, n47431, n47432, n47433, n47434,
         n47435, n47436, n47437, n47438, n47439, n47440, n47441, n47442,
         n47443, n47444, n47445, n47446, n47447, n47448, n47449, n47450,
         n47451, n47452, n47453, n47454, n47455, n47456, n47457, n47458,
         n47459, n47460, n47461, n47462, n47463, n47464, n47465, n47466,
         n47467, n47468, n47469, n47470, n47471, n47472, n47473, n47474,
         n47475, n47476, n47477, n47478, n47479, n47480, n47481, n47482,
         n47483, n47484, n47485, n47486, n47487, n47488, n47489, n47490,
         n47491, n47492, n47493, n47494, n47495, n47496, n47497, n47498,
         n47499, n47500, n47501, n47502, n47503, n47504, n47505, n47506,
         n47507, n47508, n47509, n47510, n47511, n47512, n47513, n47514,
         n47515, n47516, n47517, n47518, n47519, n47520, n47521, n47522,
         n47523, n47524, n47525, n47526, n47527, n47528, n47529, n47530,
         n47531, n47532, n47533, n47534, n47535, n47536, n47537, n47538,
         n47539, n47540, n47541, n47542, n47543, n47544, n47545, n47546,
         n47547, n47548, n47549, n47550, n47551, n47552, n47553, n47554,
         n47555, n47556, n47557, n47558, n47559, n47560, n47561, n47562,
         n47563, n47564, n47565, n47566, n47567, n47568, n47569, n47570,
         n47571, n47572, n47573, n47574, n47575, n47576, n47577, n47578,
         n47579, n47580, n47581, n47582, n47583, n47584, n47585, n47586,
         n47587, n47588, n47589, n47590, n47591, n47592, n47593, n47594,
         n47595, n47596, n47597, n47598, n47599, n47600, n47601, n47602,
         n47603, n47604, n47605, n47606, n47607, n47608, n47609, n47610,
         n47611, n47612, n47613, n47614, n47615, n47616, n47617, n47618,
         n47619, n47620, n47621, n47622, n47623, n47624, n47625, n47626,
         n47627, n47628, n47629, n47630, n47631, n47632, n47633, n47634,
         n47635, n47636, n47637, n47638, n47639, n47640, n47641, n47642,
         n47643, n47644, n47645, n47646, n47647, n47648, n47649, n47650,
         n47651, n47652, n47653, n47654, n47655, n47656, n47657, n47658,
         n47659, n47660, n47661, n47662, n47663, n47664, n47665, n47666,
         n47667, n47668, n47669, n47670, n47671, n47672, n47673, n47674,
         n47675, n47676, n47677, n47678, n47679, n47680, n47681, n47682,
         n47683, n47684, n47685, n47686, n47687, n47688, n47689, n47690,
         n47691, n47692, n47693, n47694, n47695, n47696, n47697, n47698,
         n47699, n47700, n47701, n47702, n47703, n47704, n47705, n47706,
         n47707, n47708, n47709, n47710, n47711, n47712, n47713, n47714,
         n47715, n47716, n47717, n47718, n47719, n47720, n47721, n47722,
         n47723, n47724, n47725, n47726, n47727, n47728, n47729, n47730,
         n47731, n47732, n47733, n47734, n47735, n47736, n47737, n47738,
         n47739, n47740, n47741, n47742, n47743, n47744, n47745, n47746,
         n47747, n47748, n47749, n47750, n47751, n47752, n47753, n47754,
         n47755, n47756, n47757, n47758, n47759, n47760, n47761, n47762,
         n47763, n47764, n47765, n47766, n47767, n47768, n47769, n47770,
         n47771, n47772, n47773, n47774, n47775, n47776, n47777, n47778,
         n47779, n47780, n47781, n47782, n47783, n47784, n47785, n47786,
         n47787, n47788, n47789, n47790, n47791, n47792, n47793, n47794,
         n47795, n47796, n47797, n47798, n47799, n47800, n47801, n47802,
         n47803, n47804, n47805, n47806, n47807, n47808, n47809, n47810,
         n47811, n47812, n47813, n47814, n47815, n47816, n47817, n47818,
         n47819, n47820, n47821, n47822, n47823, n47824, n47825, n47826,
         n47827, n47828, n47829, n47830, n47831, n47832, n47833, n47834,
         n47835, n47836, n47837, n47838, n47839, n47840, n47841, n47842,
         n47843, n47844, n47845, n47846, n47847, n47848, n47849, n47850,
         n47851, n47852, n47853, n47854, n47855, n47856, n47857, n47858,
         n47859, n47860, n47861, n47862, n47863, n47864, n47865, n47866,
         n47867, n47868, n47869, n47870, n47871, n47872, n47873, n47874,
         n47875, n47876, n47877, n47878, n47879, n47880, n47881, n47882,
         n47883, n47884, n47885, n47886, n47887, n47888, n47889, n47890,
         n47891, n47892, n47893, n47894, n47895, n47896, n47897, n47898,
         n47899, n47900, n47901, n47902, n47903, n47904, n47905, n47906,
         n47907, n47908, n47909, n47910, n47911, n47912, n47913, n47914,
         n47915, n47916, n47917, n47918, n47919, n47920, n47921, n47922,
         n47923, n47924, n47925, n47926, n47927, n47928, n47929, n47930,
         n47931, n47932, n47933, n47934, n47935, n47936, n47937, n47938,
         n47939, n47940, n47941, n47942, n47943, n47944, n47945, n47946,
         n47947, n47948, n47949, n47950, n47951, n47952, n47953, n47954,
         n47955, n47956, n47957, n47958, n47959, n47960, n47961, n47962,
         n47963, n47964, n47965, n47966, n47967, n47968, n47969, n47970,
         n47971, n47972, n47973, n47974, n47975, n47976, n47977, n47978,
         n47979, n47980, n47981, n47982, n47983, n47984, n47985, n47986,
         n47987, n47988, n47989, n47990, n47991, n47992, n47993, n47994,
         n47995, n47996, n47997, n47998, n47999, n48000, n48001, n48002,
         n48003, n48004, n48005, n48006, n48007, n48008, n48009, n48010,
         n48011, n48012, n48013, n48014, n48015, n48016, n48017, n48018,
         n48019, n48020, n48021, n48022, n48023, n48024, n48025, n48026,
         n48027, n48028, n48029, n48030, n48031, n48032, n48033, n48034,
         n48035, n48036, n48037, n48038, n48039, n48040, n48041, n48042,
         n48043, n48044, n48045, n48046, n48047, n48048, n48049, n48050,
         n48051, n48052, n48053, n48054, n48055, n48056, n48057, n48058,
         n48059, n48060, n48061, n48062, n48063, n48064, n48065, n48066,
         n48067, n48068, n48069, n48070, n48071, n48072, n48073, n48074,
         n48075, n48076, n48077, n48078, n48079, n48080, n48081, n48082,
         n48083, n48084, n48085, n48086, n48087, n48088, n48089, n48090,
         n48091, n48092, n48093, n48094, n48095, n48096, n48097, n48098,
         n48099, n48100, n48101, n48102, n48103, n48104, n48105, n48106,
         n48107, n48108, n48109, n48110, n48111, n48112, n48113, n48114,
         n48115, n48116, n48117, n48118, n48119, n48120, n48121, n48122,
         n48123, n48124, n48125, n48126, n48127, n48128, n48129, n48130,
         n48131, n48132, n48133, n48134, n48135, n48136, n48137, n48138,
         n48139, n48140, n48141, n48142, n48143, n48144, n48145, n48146,
         n48147, n48148, n48149, n48150, n48151, n48152, n48153, n48154,
         n48155, n48156, n48157, n48158, n48159, n48160, n48161, n48162,
         n48163, n48164, n48165, n48166, n48167, n48168, n48169, n48170,
         n48171, n48172, n48173, n48174, n48175, n48176, n48177, n48178,
         n48179, n48180, n48181, n48182, n48183, n48184, n48185, n48186,
         n48187, n48188, n48189, n48190, n48191, n48192, n48193, n48194,
         n48195, n48196, n48197, n48198, n48199, n48200, n48201, n48202,
         n48203, n48204, n48205, n48206, n48207, n48208, n48209, n48210,
         n48211, n48212, n48213, n48214, n48215, n48216, n48217, n48218,
         n48219, n48220, n48221, n48222, n48223, n48224, n48225, n48226,
         n48227, n48228, n48229, n48230, n48231, n48232, n48233, n48234,
         n48235, n48236, n48237, n48238, n48239, n48240, n48241, n48242,
         n48243, n48244, n48245, n48246, n48247, n48248, n48249, n48250,
         n48251, n48252, n48253, n48254, n48255, n48256, n48257, n48258,
         n48259, n48260, n48261, n48262, n48263, n48264, n48265, n48266,
         n48267, n48268, n48269, n48270, n48271, n48272, n48273, n48274,
         n48275, n48276, n48277, n48278, n48279, n48280, n48281, n48282,
         n48283, n48284, n48285, n48286, n48287, n48288, n48289, n48290,
         n48291, n48292, n48293, n48294, n48295, n48296, n48297, n48298,
         n48299, n48300, n48301, n48302, n48303, n48304, n48305, n48306,
         n48307, n48308, n48309, n48310, n48311, n48312, n48313, n48314,
         n48315, n48316, n48317, n48318, n48319, n48320, n48321, n48322,
         n48323, n48324, n48325, n48326, n48327, n48328, n48329, n48330,
         n48331, n48332, n48333, n48334, n48335, n48336, n48337, n48338,
         n48339, n48340, n48341, n48342, n48343, n48344, n48345, n48346,
         n48347, n48348, n48349, n48350, n48351, n48352, n48353, n48354,
         n48355, n48356, n48357, n48358, n48359, n48360, n48361, n48362,
         n48363, n48364, n48365, n48366, n48367, n48368, n48369, n48370,
         n48371, n48372, n48373, n48374, n48375, n48376, n48377, n48378,
         n48379, n48380, n48381, n48382, n48383, n48384, n48385, n48386,
         n48387, n48388, n48389, n48390, n48391, n48392, n48393, n48394,
         n48395, n48396, n48397, n48398, n48399, n48400, n48401, n48402,
         n48403, n48404, n48405, n48406, n48407, n48408, n48409, n48410,
         n48411, n48412, n48413, n48414, n48415, n48416, n48417, n48418,
         n48419, n48420, n48421, n48422, n48423, n48424, n48425, n48426,
         n48427, n48428, n48429, n48430, n48431, n48432, n48433, n48434,
         n48435, n48436, n48437, n48438, n48439, n48440, n48441, n48442,
         n48443, n48444, n48445, n48446, n48447, n48448, n48449, n48450,
         n48451, n48452, n48453, n48454, n48455, n48456, n48457, n48458,
         n48459, n48460, n48461, n48462, n48463, n48464, n48465, n48466,
         n48467, n48468, n48469, n48470, n48471, n48472, n48473, n48474,
         n48475, n48476, n48477, n48478, n48479, n48480, n48481, n48482,
         n48483, n48484, n48485, n48486, n48487, n48488, n48489, n48490,
         n48491, n48492, n48493, n48494, n48495, n48496, n48497, n48498,
         n48499, n48500, n48501, n48502, n48503, n48504, n48505, n48506,
         n48507, n48508, n48509, n48510, n48511, n48512, n48513, n48514,
         n48515, n48516, n48517, n48518, n48519, n48520, n48521, n48522,
         n48523, n48524, n48525, n48526, n48527, n48528, n48529, n48530,
         n48531, n48532, n48533, n48534, n48535, n48536, n48537, n48538,
         n48539, n48540, n48541, n48542, n48543, n48544, n48545, n48546,
         n48547, n48548, n48549, n48550, n48551, n48552, n48553, n48554,
         n48555, n48556, n48557, n48558, n48559, n48560, n48561, n48562,
         n48563, n48564, n48565, n48566, n48567, n48568, n48569, n48570,
         n48571, n48572, n48573, n48574, n48575, n48576, n48577, n48578,
         n48579, n48580, n48581, n48582, n48583, n48584, n48585, n48586,
         n48587, n48588, n48589, n48590, n48591, n48592, n48593, n48594,
         n48595, n48596, n48597, n48598, n48599, n48600, n48601, n48602,
         n48603, n48604, n48605, n48606, n48607, n48608, n48609, n48610,
         n48611, n48612, n48613, n48614, n48615, n48616, n48617, n48618,
         n48619, n48620, n48621, n48622, n48623, n48624, n48625, n48626,
         n48627, n48628, n48629, n48630, n48631, n48632, n48633, n48634,
         n48635, n48636, n48637, n48638, n48639, n48640, n48641, n48642,
         n48643, n48644, n48645, n48646, n48647, n48648, n48649, n48650,
         n48651, n48652, n48653, n48654, n48655, n48656, n48657, n48658,
         n48659, n48660, n48661, n48662, n48663, n48664, n48665, n48666,
         n48667, n48668, n48669, n48670, n48671, n48672, n48673, n48674,
         n48675, n48676, n48677, n48678, n48679, n48680, n48681, n48682,
         n48683, n48684, n48685, n48686, n48687, n48688, n48689, n48690,
         n48691, n48692, n48693, n48694, n48695, n48696, n48697, n48698,
         n48699, n48700, n48701, n48702, n48703, n48704, n48705, n48706,
         n48707, n48708, n48709, n48710, n48711, n48712, n48713, n48714,
         n48715, n48716, n48717, n48718, n48719, n48720, n48721, n48722,
         n48723, n48724, n48725, n48726, n48727, n48728, n48729, n48730,
         n48731, n48732, n48733, n48734, n48735, n48736, n48737, n48738,
         n48739, n48740, n48741, n48742, n48743, n48744, n48745, n48746,
         n48747, n48748, n48749, n48750, n48751, n48752, n48753, n48754,
         n48755, n48756, n48757, n48758, n48759, n48760, n48761, n48762,
         n48763, n48764, n48765, n48766, n48767, n48768, n48769, n48770,
         n48771, n48772, n48773, n48774, n48775, n48776, n48777, n48778,
         n48779, n48780, n48781, n48782, n48783, n48784, n48785, n48786,
         n48787, n48788, n48789, n48790, n48791, n48792, n48793, n48794,
         n48795, n48796, n48797, n48798, n48799, n48800, n48801, n48802,
         n48803, n48804, n48805, n48806, n48807, n48808, n48809, n48810,
         n48811, n48812, n48813, n48814, n48815, n48816, n48817, n48818,
         n48819, n48820, n48821, n48822, n48823, n48824, n48825, n48826,
         n48827, n48828, n48829, n48830, n48831, n48832, n48833, n48834,
         n48835, n48836, n48837, n48838, n48839, n48840, n48841, n48842,
         n48843, n48844, n48845, n48846, n48847, n48848, n48849, n48850,
         n48851, n48852, n48853, n48854, n48855, n48856, n48857, n48858,
         n48859, n48860, n48861, n48862, n48863, n48864, n48865, n48866,
         n48867, n48868, n48869, n48870, n48871, n48872, n48873, n48874,
         n48875, n48876, n48877, n48878, n48879, n48880, n48881, n48882,
         n48883, n48884, n48885, n48886, n48887, n48888, n48889, n48890,
         n48891, n48892, n48893, n48894, n48895, n48896, n48897, n48898,
         n48899, n48900, n48901, n48902, n48903, n48904, n48905, n48906,
         n48907, n48908, n48909, n48910, n48911, n48912, n48913, n48914,
         n48915, n48916, n48917, n48918, n48919, n48920, n48921, n48922,
         n48923, n48924, n48925, n48926, n48927, n48928, n48929, n48930,
         n48931, n48932, n48933, n48934, n48935, n48936, n48937, n48938,
         n48939, n48940, n48941, n48942, n48943, n48944, n48945, n48946,
         n48947, n48948, n48949, n48950, n48951, n48952, n48953, n48954,
         n48955, n48956, n48957, n48958, n48959, n48960, n48961, n48962,
         n48963, n48964, n48965, n48966, n48967, n48968, n48969, n48970,
         n48971, n48972, n48973, n48974, n48975, n48976, n48977, n48978,
         n48979, n48980, n48981, n48982, n48983, n48984, n48985, n48986,
         n48987, n48988, n48989, n48990, n48991, n48992, n48993, n48994,
         n48995, n48996, n48997, n48998, n48999, n49000, n49001, n49002,
         n49003, n49004, n49005, n49006, n49007, n49008, n49009, n49010,
         n49011, n49012, n49013, n49014, n49015, n49016, n49017, n49018,
         n49019, n49020, n49021, n49022, n49023, n49024, n49025, n49026,
         n49027, n49028, n49029, n49030, n49031, n49032, n49033, n49034,
         n49035, n49036, n49037, n49038, n49039, n49040, n49041, n49042,
         n49043, n49044, n49045, n49046, n49047, n49048, n49049, n49050,
         n49051, n49052, n49053, n49054, n49055, n49056, n49057, n49058,
         n49059, n49060, n49061, n49062, n49063, n49064, n49065, n49066,
         n49067, n49068, n49069, n49070, n49071, n49072, n49073, n49074,
         n49075, n49076, n49077, n49078, n49079, n49080, n49081, n49082,
         n49083, n49084, n49085, n49086, n49087, n49088, n49089, n49090,
         n49091, n49092, n49093, n49094, n49095, n49096, n49097, n49098,
         n49099, n49100, n49101, n49102, n49103, n49104, n49105, n49106,
         n49107, n49108, n49109, n49110, n49111, n49112, n49113, n49114,
         n49115, n49116, n49117, n49118, n49119, n49120, n49121, n49122,
         n49123, n49124, n49125, n49126, n49127, n49128, n49129, n49130,
         n49131, n49132, n49133, n49134, n49135, n49136, n49137, n49138,
         n49139, n49140, n49141, n49142, n49143, n49144, n49145, n49146,
         n49147, n49148, n49149, n49150, n49151, n49152, n49153, n49154,
         n49155, n49156, n49157, n49158, n49159, n49160, n49161, n49162,
         n49163, n49164, n49165, n49166, n49167, n49168, n49169, n49170,
         n49171, n49172, n49173, n49174, n49175, n49176, n49177, n49178,
         n49179, n49180, n49181, n49182, n49183, n49184, n49185, n49186,
         n49187, n49188, n49189, n49190, n49191, n49192, n49193, n49194,
         n49195, n49196, n49197, n49198, n49199, n49200, n49201, n49202,
         n49203, n49204, n49205, n49206, n49207, n49208, n49209, n49210,
         n49211, n49212, n49213, n49214, n49215, n49216, n49217, n49218,
         n49219, n49220, n49221, n49222, n49223, n49224, n49225, n49226,
         n49227, n49228, n49229, n49230, n49231, n49232, n49233, n49234,
         n49235, n49236, n49237, n49238, n49239, n49240, n49241, n49242,
         n49243, n49244, n49245, n49246, n49247, n49248, n49249, n49250,
         n49251, n49252, n49253, n49254, n49255, n49256, n49257, n49258,
         n49259, n49260, n49261, n49262, n49263, n49264, n49265, n49266,
         n49267, n49268, n49269, n49270, n49271, n49272, n49273, n49274,
         n49275, n49276, n49277, n49278, n49279, n49280, n49281, n49282,
         n49283, n49284, n49285, n49286, n49287, n49288, n49289, n49290,
         n49291, n49292, n49293, n49294, n49295, n49296, n49297, n49298,
         n49299, n49300, n49301, n49302, n49303, n49304, n49305, n49306,
         n49307, n49308, n49309, n49310, n49311, n49312, n49313, n49314,
         n49315, n49316, n49317, n49318, n49319, n49320, n49321, n49322,
         n49323, n49324, n49325, n49326, n49327, n49328, n49329, n49330,
         n49331, n49332, n49333, n49334, n49335, n49336, n49337, n49338,
         n49339, n49340, n49341, n49342, n49343, n49344, n49345, n49346,
         n49347, n49348, n49349, n49350, n49351, n49352, n49353, n49354,
         n49355, n49356, n49357, n49358, n49359, n49360, n49361, n49362,
         n49363, n49364, n49365, n49366, n49367, n49368, n49369, n49370,
         n49371, n49372, n49373, n49374, n49375, n49376, n49377, n49378,
         n49379, n49380, n49381, n49382, n49383, n49384, n49385, n49386,
         n49387, n49388, n49389, n49390, n49391, n49392, n49393, n49394,
         n49395, n49396, n49397, n49398, n49399, n49400, n49401, n49402,
         n49403, n49404, n49405, n49406, n49407, n49408, n49409, n49410,
         n49411, n49412, n49413, n49414, n49415, n49416, n49417, n49418,
         n49419, n49420, n49421, n49422, n49423, n49424, n49425, n49426,
         n49427, n49428, n49429, n49430, n49431, n49432, n49433, n49434,
         n49435, n49436, n49437, n49438, n49439, n49440, n49441, n49442,
         n49443, n49444, n49445, n49446, n49447, n49448, n49449, n49450,
         n49451, n49452, n49453, n49454, n49455, n49456, n49457, n49458,
         n49459, n49460, n49461, n49462, n49463, n49464, n49465, n49466,
         n49467, n49468, n49469, n49470, n49471, n49472, n49473, n49474,
         n49475, n49476, n49477, n49478, n49479, n49480, n49481, n49482,
         n49483, n49484, n49485, n49486, n49487, n49488, n49489, n49490,
         n49491, n49492, n49493, n49494, n49495, n49496, n49497, n49498,
         n49499, n49500, n49501, n49502, n49503, n49504, n49505, n49506,
         n49507, n49508, n49509, n49510, n49511, n49512, n49513, n49514,
         n49515, n49516, n49517, n49518, n49519, n49520, n49521, n49522,
         n49523, n49524, n49525, n49526, n49527, n49528, n49529, n49530,
         n49531, n49532, n49533, n49534, n49535, n49536, n49537, n49538,
         n49539, n49540, n49541, n49542, n49543, n49544, n49545, n49546,
         n49547, n49548, n49549, n49550, n49551, n49552, n49553, n49554,
         n49555, n49556, n49557, n49558, n49559, n49560, n49561, n49562,
         n49563, n49564, n49565, n49566, n49567, n49568, n49569, n49570,
         n49571, n49572, n49573, n49574, n49575, n49576, n49577, n49578,
         n49579, n49580, n49581, n49582, n49583, n49584, n49585, n49586,
         n49587, n49588, n49589, n49590, n49591, n49592, n49593, n49594,
         n49595, n49596, n49597, n49598, n49599, n49600, n49601, n49602,
         n49603, n49604, n49605, n49606, n49607, n49608, n49609, n49610,
         n49611, n49612, n49613, n49614, n49615, n49616, n49617, n49618,
         n49619, n49620, n49621, n49622, n49623, n49624, n49625, n49626,
         n49627, n49628, n49629, n49630, n49631, n49632, n49633, n49634,
         n49635, n49636, n49637, n49638, n49639, n49640, n49641, n49642,
         n49643, n49644, n49645, n49646, n49647, n49648, n49649, n49650,
         n49651, n49652, n49653, n49654, n49655, n49656, n49657, n49658,
         n49659, n49660, n49661, n49662, n49663, n49664, n49665, n49666,
         n49667, n49668, n49669, n49670, n49671, n49672, n49673, n49674,
         n49675, n49676, n49677, n49678, n49679, n49680, n49681, n49682,
         n49683, n49684, n49685, n49686, n49687, n49688, n49689, n49690,
         n49691, n49692, n49693, n49694, n49695, n49696, n49697, n49698,
         n49699, n49700, n49701, n49702, n49703, n49704, n49705, n49706,
         n49707, n49708, n49709, n49710, n49711, n49712, n49713, n49714,
         n49715, n49716, n49717, n49718, n49719, n49720, n49721, n49722,
         n49723, n49724, n49725, n49726, n49727, n49728, n49729, n49730,
         n49731, n49732, n49733, n49734, n49735, n49736, n49737, n49738,
         n49739, n49740, n49741, n49742, n49743, n49744, n49745, n49746,
         n49747, n49748, n49749, n49750, n49751, n49752, n49753, n49754,
         n49755, n49756, n49757, n49758, n49759, n49760, n49761, n49762,
         n49763, n49764, n49765, n49766, n49767, n49768, n49769, n49770,
         n49771, n49772, n49773, n49774, n49775, n49776, n49777, n49778,
         n49779, n49780, n49781, n49782, n49783, n49784, n49785, n49786,
         n49787, n49788, n49789, n49790, n49791, n49792, n49793, n49794,
         n49795, n49796, n49797, n49798, n49799, n49800, n49801, n49802,
         n49803, n49804, n49805, n49806, n49807, n49808, n49809, n49810,
         n49811, n49812, n49813, n49814, n49815, n49816, n49817, n49818,
         n49819, n49820, n49821, n49822, n49823, n49824, n49825, n49826,
         n49827, n49828, n49829, n49830, n49831, n49832, n49833, n49834,
         n49835, n49836, n49837, n49838, n49839, n49840, n49841, n49842,
         n49843, n49844, n49845, n49846, n49847, n49848, n49849, n49850,
         n49851, n49852, n49853, n49854, n49855, n49856, n49857, n49858,
         n49859, n49860, n49861, n49862, n49863, n49864, n49865, n49866,
         n49867, n49868, n49869, n49870, n49871, n49872, n49873, n49874,
         n49875, n49876, n49877, n49878, n49879, n49880, n49881, n49882,
         n49883, n49884, n49885, n49886, n49887, n49888, n49889, n49890,
         n49891, n49892, n49893, n49894, n49895, n49896, n49897, n49898,
         n49899, n49900, n49901, n49902, n49903, n49904, n49905, n49906,
         n49907, n49908, n49909, n49910, n49911, n49912, n49913, n49914,
         n49915, n49916, n49917, n49918, n49919, n49920, n49921, n49922,
         n49923, n49924, n49925, n49926, n49927, n49928, n49929, n49930,
         n49931, n49932, n49933, n49934, n49935, n49936, n49937, n49938,
         n49939, n49940, n49941, n49942, n49943, n49944, n49945, n49946,
         n49947, n49948, n49949, n49950, n49951, n49952, n49953, n49954,
         n49955, n49956, n49957, n49958, n49959, n49960, n49961, n49962,
         n49963, n49964, n49965, n49966, n49967, n49968, n49969, n49970,
         n49971, n49972, n49973, n49974, n49975, n49976, n49977, n49978,
         n49979, n49980, n49981, n49982, n49983, n49984, n49985, n49986,
         n49987, n49988, n49989, n49990, n49991, n49992, n49993, n49994,
         n49995, n49996, n49997, n49998, n49999, n50000, n50001, n50002,
         n50003, n50004, n50005, n50006, n50007, n50008, n50009, n50010,
         n50011, n50012, n50013, n50014, n50015, n50016, n50017, n50018,
         n50019, n50020, n50021, n50022, n50023, n50024, n50025, n50026,
         n50027, n50028, n50029, n50030, n50031, n50032, n50033, n50034,
         n50035, n50036, n50037, n50038, n50039, n50040, n50041, n50042,
         n50043, n50044, n50045, n50046, n50047, n50048, n50049, n50050,
         n50051, n50052, n50053, n50054, n50055, n50056, n50057, n50058,
         n50059, n50060, n50061, n50062, n50063, n50064, n50065, n50066,
         n50067, n50068, n50069, n50070, n50071, n50072, n50073, n50074,
         n50075, n50076, n50077, n50078, n50079, n50080, n50081, n50082,
         n50083, n50084, n50085, n50086, n50087, n50088, n50089, n50090,
         n50091, n50092, n50093, n50094, n50095, n50096, n50097, n50098,
         n50099, n50100, n50101, n50102, n50103, n50104, n50105, n50106,
         n50107, n50108, n50109, n50110, n50111, n50112, n50113, n50114,
         n50115, n50116, n50117, n50118, n50119, n50120, n50121, n50122,
         n50123, n50124, n50125, n50126, n50127, n50128, n50129, n50130,
         n50131, n50132, n50133, n50134, n50135, n50136, n50137, n50138,
         n50139, n50140, n50141, n50142, n50143, n50144, n50145, n50146,
         n50147, n50148, n50149, n50150, n50151, n50152, n50153, n50154,
         n50155, n50156, n50157, n50158, n50159, n50160, n50161, n50162,
         n50163, n50164, n50165, n50166, n50167, n50168, n50169, n50170,
         n50171, n50172, n50173, n50174, n50175, n50176, n50177, n50178,
         n50179, n50180, n50181, n50182, n50183, n50184, n50185, n50186,
         n50187, n50188, n50189, n50190, n50191, n50192, n50193, n50194,
         n50195, n50196, n50197, n50198, n50199, n50200, n50201, n50202,
         n50203, n50204, n50205, n50206, n50207, n50208, n50209, n50210,
         n50211, n50212, n50213, n50214, n50215, n50216, n50217, n50218,
         n50219, n50220, n50221, n50222, n50223, n50224, n50225, n50226,
         n50227, n50228, n50229, n50230, n50231, n50232, n50233, n50234,
         n50235, n50236, n50237, n50238, n50239, n50240, n50241, n50242,
         n50243, n50244, n50245, n50246, n50247, n50248, n50249, n50250,
         n50251, n50252, n50253, n50254, n50255, n50256, n50257, n50258,
         n50259, n50260, n50261, n50262, n50263, n50264, n50265, n50266,
         n50267, n50268, n50269, n50270, n50271, n50272, n50273, n50274,
         n50275, n50276, n50277, n50278, n50279, n50280, n50281, n50282,
         n50283, n50284, n50285, n50286, n50287, n50288, n50289, n50290,
         n50291, n50292, n50293, n50294, n50295, n50296, n50297, n50298,
         n50299, n50300, n50301, n50302, n50303, n50304, n50305, n50306,
         n50307, n50308, n50309, n50310, n50311, n50312, n50313, n50314,
         n50315, n50316, n50317, n50318, n50319, n50320, n50321, n50322,
         n50323, n50324, n50325, n50326, n50327, n50328, n50329, n50330,
         n50331, n50332, n50333, n50334, n50335, n50336, n50337, n50338,
         n50339, n50340, n50341, n50342, n50343, n50344, n50345, n50346,
         n50347, n50348, n50349, n50350, n50351, n50352, n50353, n50354,
         n50355, n50356, n50357, n50358, n50359, n50360, n50361, n50362,
         n50363, n50364, n50365, n50366, n50367, n50368, n50369, n50370,
         n50371, n50372, n50373, n50374, n50375, n50376, n50377, n50378,
         n50379, n50380, n50381, n50382, n50383, n50384, n50385, n50386,
         n50387, n50388, n50389, n50390, n50391, n50392, n50393, n50394,
         n50395, n50396, n50397, n50398, n50399, n50400, n50401, n50402,
         n50403, n50404, n50405, n50406, n50407, n50408, n50409, n50410,
         n50411, n50412, n50413, n50414, n50415, n50416, n50417, n50418,
         n50419, n50420, n50421, n50422, n50423, n50424, n50425, n50426,
         n50427, n50428, n50429, n50430, n50431, n50432, n50433, n50434,
         n50435, n50436, n50437, n50438, n50439, n50440, n50441, n50442,
         n50443, n50444, n50445, n50446, n50447, n50448, n50449, n50450,
         n50451, n50452, n50453, n50454, n50455, n50456, n50457, n50458,
         n50459, n50460, n50461, n50462, n50463, n50464, n50465, n50466,
         n50467, n50468, n50469, n50470, n50471, n50472, n50473, n50474,
         n50475, n50476, n50477, n50478, n50479, n50480, n50481, n50482,
         n50483, n50484, n50485, n50486, n50487, n50488, n50489, n50490,
         n50491, n50492, n50493, n50494, n50495, n50496, n50497, n50498,
         n50499, n50500, n50501, n50502, n50503, n50504, n50505, n50506,
         n50507, n50508, n50509, n50510, n50511, n50512, n50513, n50514,
         n50515, n50516, n50517, n50518, n50519, n50520, n50521, n50522,
         n50523, n50524, n50525, n50526, n50527, n50528, n50529, n50530,
         n50531, n50532, n50533, n50534, n50535, n50536, n50537, n50538,
         n50539, n50540, n50541, n50542, n50543, n50544, n50545, n50546,
         n50547, n50548, n50549, n50550, n50551, n50552, n50553, n50554,
         n50555, n50556, n50557, n50558, n50559, n50560, n50561, n50562,
         n50563, n50564, n50565, n50566, n50567, n50568, n50569, n50570,
         n50571, n50572, n50573, n50574, n50575, n50576, n50577, n50578,
         n50579, n50580, n50581, n50582, n50583, n50584, n50585, n50586,
         n50587, n50588, n50589, n50590, n50591, n50592, n50593, n50594,
         n50595, n50596, n50597, n50598, n50599, n50600, n50601, n50602,
         n50603, n50604, n50605, n50606, n50607, n50608, n50609, n50610,
         n50611, n50612, n50613, n50614, n50615, n50616, n50617, n50618,
         n50619, n50620, n50621, n50622, n50623, n50624, n50625, n50626,
         n50627, n50628, n50629, n50630, n50631, n50632, n50633, n50634,
         n50635, n50636, n50637, n50638, n50639, n50640, n50641, n50642,
         n50643, n50644, n50645, n50646, n50647, n50648, n50649, n50650,
         n50651, n50652, n50653, n50654, n50655, n50656, n50657, n50658,
         n50659, n50660, n50661, n50662, n50663, n50664, n50665, n50666,
         n50667, n50668, n50669, n50670, n50671, n50672, n50673, n50674,
         n50675, n50676, n50677, n50678, n50679, n50680, n50681, n50682,
         n50683, n50684, n50685, n50686, n50687, n50688, n50689, n50690,
         n50691, n50692, n50693, n50694, n50695, n50696, n50697, n50698,
         n50699, n50700, n50701, n50702, n50703, n50704, n50705, n50706,
         n50707, n50708, n50709, n50710, n50711, n50712, n50713, n50714,
         n50715, n50716, n50717, n50718, n50719, n50720, n50721, n50722,
         n50723, n50724, n50725, n50726, n50727, n50728, n50729, n50730,
         n50731, n50732, n50733, n50734, n50735, n50736, n50737, n50738,
         n50739, n50740, n50741, n50742, n50743, n50744, n50745, n50746,
         n50747, n50748, n50749, n50750, n50751, n50752, n50753, n50754,
         n50755, n50756, n50757, n50758, n50759, n50760, n50761, n50762,
         n50763, n50764, n50765, n50766, n50767, n50768, n50769, n50770,
         n50771, n50772, n50773, n50774, n50775, n50776, n50777, n50778,
         n50779, n50780, n50781, n50782, n50783, n50784, n50785, n50786,
         n50787, n50788, n50789, n50790, n50791, n50792, n50793, n50794,
         n50795, n50796, n50797, n50798, n50799, n50800, n50801, n50802,
         n50803, n50804, n50805, n50806, n50807, n50808, n50809, n50810,
         n50811, n50812, n50813, n50814, n50815, n50816, n50817, n50818,
         n50819, n50820, n50821, n50822, n50823, n50824, n50825, n50826,
         n50827, n50828, n50829, n50830, n50831, n50832, n50833, n50834,
         n50835, n50836, n50837, n50838, n50839, n50840, n50841, n50842,
         n50843, n50844, n50845, n50846, n50847, n50848, n50849, n50850,
         n50851, n50852, n50853, n50854, n50855, n50856, n50857, n50858,
         n50859, n50860, n50861, n50862, n50863, n50864, n50865, n50866,
         n50867, n50868, n50869, n50870, n50871, n50872, n50873, n50874,
         n50875, n50876, n50877, n50878, n50879, n50880, n50881, n50882,
         n50883, n50884, n50885, n50886, n50887, n50888, n50889, n50890,
         n50891, n50892, n50893, n50894, n50895, n50896, n50897, n50898,
         n50899, n50900, n50901, n50902, n50903, n50904, n50905, n50906,
         n50907, n50908, n50909, n50910, n50911, n50912, n50913, n50914,
         n50915, n50916, n50917, n50918, n50919, n50920, n50921, n50922,
         n50923, n50924, n50925, n50926, n50927, n50928, n50929, n50930,
         n50931, n50932, n50933, n50934, n50935, n50936, n50937, n50938,
         n50939, n50940, n50941, n50942, n50943, n50944, n50945, n50946,
         n50947, n50948, n50949, n50950, n50951, n50952, n50953, n50954,
         n50955, n50956, n50957, n50958, n50959, n50960, n50961, n50962,
         n50963, n50964, n50965, n50966, n50967, n50968, n50969, n50970,
         n50971, n50972, n50973, n50974, n50975, n50976, n50977, n50978,
         n50979, n50980, n50981, n50982, n50983, n50984, n50985, n50986,
         n50987, n50988, n50989, n50990, n50991, n50992, n50993, n50994,
         n50995, n50996, n50997, n50998, n50999, n51000, n51001, n51002,
         n51003, n51004, n51005, n51006, n51007, n51008, n51009, n51010,
         n51011, n51012, n51013, n51014, n51015, n51016, n51017, n51018,
         n51019, n51020, n51021, n51022, n51023, n51024, n51025, n51026,
         n51027, n51028, n51029, n51030, n51031, n51032, n51033, n51034,
         n51035, n51036, n51037, n51038, n51039, n51040, n51041, n51042,
         n51043, n51044, n51045, n51046, n51047, n51048, n51049, n51050,
         n51051, n51052, n51053, n51054, n51055, n51056, n51057, n51058,
         n51059, n51060, n51061, n51062, n51063, n51064, n51065, n51066,
         n51067, n51068, n51069, n51070, n51071, n51072, n51073, n51074,
         n51075, n51076, n51077, n51078, n51079, n51080, n51081, n51082,
         n51083, n51084, n51085, n51086, n51087, n51088, n51089, n51090,
         n51091, n51092, n51093, n51094, n51095, n51096, n51097, n51098,
         n51099, n51100, n51101, n51102, n51103, n51104, n51105, n51106,
         n51107, n51108, n51109, n51110, n51111, n51112, n51113, n51114,
         n51115, n51116, n51117, n51118, n51119, n51120, n51121, n51122,
         n51123, n51124, n51125, n51126, n51127, n51128, n51129, n51130,
         n51131, n51132, n51133, n51134, n51135, n51136, n51137, n51138,
         n51139, n51140, n51141, n51142, n51143, n51144, n51145, n51146,
         n51147, n51148, n51149, n51150, n51151, n51152, n51153, n51154,
         n51155, n51156, n51157, n51158, n51159, n51160, n51161, n51162,
         n51163, n51164, n51165, n51166, n51167, n51168, n51169, n51170,
         n51171, n51172, n51173, n51174, n51175, n51176, n51177, n51178,
         n51179, n51180, n51181, n51182, n51183, n51184, n51185, n51186,
         n51187, n51188, n51189, n51190, n51191, n51192, n51193, n51194,
         n51195, n51196, n51197, n51198, n51199, n51200, n51201, n51202,
         n51203, n51204, n51205, n51206, n51207, n51208, n51209, n51210,
         n51211, n51212, n51213, n51214, n51215, n51216, n51217, n51218,
         n51219, n51220, n51221, n51222, n51223, n51224, n51225, n51226,
         n51227, n51228, n51229, n51230, n51231, n51232, n51233, n51234,
         n51235, n51236, n51237, n51238, n51239, n51240, n51241, n51242,
         n51243, n51244, n51245, n51246, n51247, n51248, n51249, n51250,
         n51251, n51252, n51253, n51254, n51255, n51256, n51257, n51258,
         n51259, n51260, n51261, n51262, n51263, n51264, n51265, n51266,
         n51267, n51268, n51269, n51270, n51271, n51272, n51273, n51274,
         n51275, n51276, n51277, n51278, n51279, n51280, n51281, n51282,
         n51283, n51284, n51285, n51286, n51287, n51288, n51289, n51290,
         n51291, n51292, n51293, n51294, n51295, n51296, n51297, n51298,
         n51299, n51300, n51301, n51302, n51303, n51304, n51305, n51306,
         n51307, n51308, n51309, n51310, n51311, n51312, n51313, n51314,
         n51315, n51316, n51317, n51318, n51319, n51320, n51321, n51322,
         n51323, n51324, n51325, n51326, n51327, n51328, n51329, n51330,
         n51331, n51332, n51333, n51334, n51335, n51336, n51337, n51338,
         n51339, n51340, n51341, n51342, n51343, n51344, n51345, n51346,
         n51347, n51348, n51349, n51350, n51351, n51352, n51353, n51354,
         n51355, n51356, n51357, n51358, n51359, n51360, n51361, n51362,
         n51363, n51364, n51365, n51366, n51367, n51368, n51369, n51370,
         n51371, n51372, n51373, n51374, n51375, n51376, n51377, n51378,
         n51379, n51380, n51381, n51382, n51383, n51384, n51385, n51386,
         n51387, n51388, n51389, n51390, n51391, n51392, n51393, n51394,
         n51395, n51396, n51397, n51398, n51399, n51400, n51401, n51402,
         n51403, n51404, n51405, n51406, n51407, n51408, n51409, n51410,
         n51411, n51412, n51413, n51414, n51415, n51416, n51417, n51418,
         n51419, n51420, n51421, n51422, n51423, n51424, n51425, n51426,
         n51427, n51428, n51429, n51430, n51431, n51432, n51433, n51434,
         n51435, n51436, n51437, n51438, n51439, n51440, n51441, n51442,
         n51443, n51444, n51445, n51446, n51447, n51448, n51449, n51450,
         n51451, n51452, n51453, n51454, n51455, n51456, n51457, n51458,
         n51459, n51460, n51461, n51462, n51463, n51464, n51465, n51466,
         n51467, n51468, n51469, n51470, n51471, n51472, n51473, n51474,
         n51475, n51476, n51477, n51478, n51479, n51480, n51481, n51482,
         n51483, n51484, n51485, n51486, n51487, n51488, n51489, n51490,
         n51491, n51492, n51493, n51494, n51495, n51496, n51497, n51498,
         n51499, n51500, n51501, n51502, n51503, n51504, n51505, n51506,
         n51507, n51508, n51509, n51510, n51511, n51512, n51513, n51514,
         n51515, n51516, n51517, n51518, n51519, n51520, n51521, n51522,
         n51523, n51524, n51525, n51526, n51527, n51528, n51529, n51530,
         n51531, n51532, n51533, n51534, n51535, n51536, n51537, n51538,
         n51539, n51540, n51541, n51542, n51543, n51544, n51545, n51546,
         n51547, n51548, n51549, n51550, n51551, n51552, n51553, n51554,
         n51555, n51556, n51557, n51558, n51559, n51560, n51561, n51562,
         n51563, n51564, n51565, n51566, n51567, n51568, n51569, n51570,
         n51571, n51572, n51573, n51574, n51575, n51576, n51577, n51578,
         n51579, n51580, n51581, n51582, n51583, n51584, n51585, n51586,
         n51587, n51588, n51589, n51590, n51591, n51592, n51593, n51594,
         n51595, n51596, n51597, n51598, n51599, n51600, n51601, n51602,
         n51603, n51604, n51605, n51606, n51607, n51608, n51609, n51610,
         n51611, n51612, n51613, n51614, n51615, n51616, n51617, n51618,
         n51619, n51620, n51621, n51622, n51623, n51624, n51625, n51626,
         n51627, n51628, n51629, n51630, n51631, n51632, n51633, n51634,
         n51635, n51636, n51637, n51638, n51639, n51640, n51641, n51642,
         n51643, n51644, n51645, n51646, n51647, n51648, n51649, n51650,
         n51651, n51652, n51653, n51654, n51655, n51656, n51657, n51658,
         n51659, n51660, n51661, n51662, n51663, n51664, n51665, n51666,
         n51667, n51668, n51669, n51670, n51671, n51672, n51673, n51674,
         n51675, n51676, n51677, n51678, n51679, n51680, n51681, n51682,
         n51683, n51684, n51685, n51686, n51687, n51688, n51689, n51690,
         n51691, n51692, n51693, n51694, n51695, n51696, n51697, n51698,
         n51699, n51700, n51701, n51702, n51703, n51704, n51705, n51706,
         n51707, n51708, n51709, n51710, n51711, n51712, n51713, n51714,
         n51715, n51716, n51717, n51718, n51719, n51720, n51721, n51722,
         n51723, n51724, n51725, n51726, n51727, n51728, n51729, n51730,
         n51731, n51732, n51733, n51734, n51735, n51736, n51737, n51738,
         n51739, n51740, n51741, n51742, n51743, n51744, n51745, n51746,
         n51747, n51748, n51749, n51750, n51751, n51752, n51753, n51754,
         n51755, n51756, n51757, n51758, n51759, n51760, n51761, n51762,
         n51763, n51764, n51765, n51766, n51767, n51768, n51769, n51770,
         n51771, n51772, n51773, n51774, n51775, n51776, n51777, n51778,
         n51779, n51780, n51781, n51782, n51783, n51784, n51785, n51786,
         n51787, n51788, n51789, n51790, n51791, n51792, n51793, n51794,
         n51795, n51796, n51797, n51798, n51799, n51800, n51801, n51802,
         n51803, n51804, n51805, n51806, n51807, n51808, n51809, n51810,
         n51811, n51812, n51813, n51814, n51815, n51816, n51817, n51818,
         n51819, n51820, n51821, n51822, n51823, n51824, n51825, n51826,
         n51827, n51828, n51829, n51830, n51831, n51832, n51833, n51834,
         n51835, n51836, n51837, n51838, n51839, n51840, n51841, n51842,
         n51843, n51844, n51845, n51846, n51847, n51848, n51849, n51850,
         n51851, n51852, n51853, n51854, n51855, n51856, n51857, n51858,
         n51859, n51860, n51861, n51862, n51863, n51864, n51865, n51866,
         n51867, n51868, n51869, n51870, n51871, n51872, n51873, n51874,
         n51875, n51876, n51877, n51878, n51879, n51880, n51881, n51882,
         n51883, n51884, n51885, n51886, n51887, n51888, n51889, n51890,
         n51891, n51892, n51893, n51894, n51895, n51896, n51897, n51898,
         n51899, n51900, n51901, n51902, n51903, n51904, n51905, n51906,
         n51907, n51908, n51909, n51910, n51911, n51912, n51913, n51914,
         n51915, n51916, n51917, n51918, n51919, n51920, n51921, n51922,
         n51923, n51924, n51925, n51926, n51927, n51928, n51929, n51930,
         n51931, n51932, n51933, n51934, n51935, n51936, n51937, n51938,
         n51939, n51940, n51941, n51942, n51943, n51944, n51945, n51946,
         n51947, n51948, n51949, n51950, n51951, n51952, n51953, n51954,
         n51955, n51956, n51957, n51958, n51959, n51960, n51961, n51962,
         n51963, n51964, n51965, n51966, n51967, n51968, n51969, n51970,
         n51971, n51972, n51973, n51974, n51975, n51976, n51977, n51978,
         n51979, n51980, n51981, n51982, n51983, n51984, n51985, n51986,
         n51987, n51988, n51989, n51990, n51991, n51992, n51993, n51994,
         n51995, n51996, n51997, n51998, n51999, n52000, n52001, n52002,
         n52003, n52004, n52005, n52006, n52007, n52008, n52009, n52010,
         n52011, n52012, n52013, n52014, n52015, n52016, n52017, n52018,
         n52019, n52020, n52021, n52022, n52023, n52024, n52025, n52026,
         n52027, n52028, n52029, n52030, n52031, n52032, n52033, n52034,
         n52035, n52036, n52037, n52038, n52039, n52040, n52041, n52042,
         n52043, n52044, n52045, n52046, n52047, n52048, n52049, n52050,
         n52051, n52052, n52053, n52054, n52055, n52056, n52057, n52058,
         n52059, n52060, n52061, n52062, n52063, n52064, n52065, n52066,
         n52067, n52068, n52069, n52070, n52071, n52072, n52073, n52074,
         n52075, n52076, n52077, n52078, n52079, n52080, n52081, n52082,
         n52083, n52084, n52085, n52086, n52087, n52088, n52089, n52090,
         n52091, n52092, n52093, n52094, n52095, n52096, n52097, n52098,
         n52099, n52100, n52101, n52102, n52103, n52104, n52105, n52106,
         n52107, n52108, n52109, n52110, n52111, n52112, n52113, n52114,
         n52115, n52116, n52117, n52118, n52119, n52120, n52121, n52122,
         n52123, n52124, n52125, n52126, n52127, n52128, n52129, n52130,
         n52131, n52132, n52133, n52134, n52135, n52136, n52137, n52138,
         n52139, n52140, n52141, n52142, n52143, n52144, n52145, n52146,
         n52147, n52148, n52149, n52150, n52151, n52152, n52153, n52154,
         n52155, n52156, n52157, n52158, n52159, n52160, n52161, n52162,
         n52163, n52164, n52165, n52166, n52167, n52168, n52169, n52170,
         n52171, n52172, n52173, n52174, n52175, n52176, n52177, n52178,
         n52179, n52180, n52181, n52182, n52183, n52184, n52185, n52186,
         n52187, n52188, n52189, n52190, n52191, n52192, n52193, n52194,
         n52195, n52196, n52197, n52198, n52199, n52200, n52201, n52202,
         n52203, n52204, n52205, n52206, n52207, n52208, n52209, n52210,
         n52211, n52212, n52213, n52214, n52215, n52216, n52217, n52218,
         n52219, n52220, n52221, n52222, n52223, n52224, n52225, n52226,
         n52227, n52228, n52229, n52230, n52231, n52232, n52233, n52234,
         n52235, n52236, n52237, n52238, n52239, n52240, n52241, n52242,
         n52243, n52244, n52245, n52246, n52247, n52248, n52249, n52250,
         n52251, n52252, n52253, n52254, n52255, n52256, n52257, n52258,
         n52259, n52260, n52261, n52262, n52263, n52264, n52265, n52266,
         n52267, n52268, n52269, n52270, n52271, n52272, n52273, n52274,
         n52275, n52276, n52277, n52278, n52279, n52280, n52281, n52282,
         n52283, n52284, n52285, n52286, n52287, n52288, n52289, n52290,
         n52291, n52292, n52293, n52294, n52295, n52296, n52297, n52298,
         n52299, n52300, n52301, n52302, n52303, n52304, n52305, n52306,
         n52307, n52308, n52309, n52310, n52311, n52312, n52313, n52314,
         n52315, n52316, n52317, n52318, n52319, n52320, n52321, n52322,
         n52323, n52324, n52325, n52326, n52327, n52328, n52329, n52330,
         n52331, n52332, n52333, n52334, n52335, n52336, n52337, n52338,
         n52339, n52340, n52341, n52342, n52343, n52344, n52345, n52346,
         n52347, n52348, n52349, n52350, n52351, n52352, n52353, n52354,
         n52355, n52356, n52357, n52358, n52359, n52360, n52361, n52362,
         n52363, n52364, n52365, n52366, n52367, n52368, n52369, n52370,
         n52371, n52372, n52373, n52374, n52375, n52376, n52377, n52378,
         n52379, n52380, n52381, n52382, n52383, n52384, n52385, n52386,
         n52387, n52388, n52389, n52390, n52391, n52392, n52393, n52394,
         n52395, n52396, n52397, n52398, n52399, n52400, n52401, n52402,
         n52403, n52404, n52405, n52406, n52407, n52408, n52409, n52410,
         n52411, n52412, n52413, n52414, n52415, n52416, n52417, n52418,
         n52419, n52420, n52421, n52422, n52423, n52424, n52425, n52426,
         n52427, n52428, n52429, n52430, n52431, n52432, n52433, n52434,
         n52435, n52436, n52437, n52438, n52439, n52440, n52441, n52442,
         n52443, n52444, n52445, n52446, n52447, n52448, n52449, n52450,
         n52451, n52452, n52453, n52454, n52455, n52456, n52457, n52458,
         n52459, n52460, n52461, n52462, n52463, n52464, n52465, n52466,
         n52467, n52468, n52469, n52470, n52471, n52472, n52473, n52474,
         n52475, n52476, n52477, n52478, n52479, n52480, n52481, n52482,
         n52483, n52484, n52485, n52486, n52487, n52488, n52489, n52490,
         n52491, n52492, n52493, n52494, n52495, n52496, n52497, n52498,
         n52499, n52500, n52501, n52502, n52503, n52504, n52505, n52506,
         n52507, n52508, n52509, n52510, n52511, n52512, n52513, n52514,
         n52515, n52516, n52517, n52518, n52519, n52520, n52521, n52522,
         n52523, n52524, n52525, n52526, n52527, n52528, n52529, n52530,
         n52531, n52532, n52533, n52534, n52535, n52536, n52537, n52538,
         n52539, n52540, n52541, n52542, n52543, n52544, n52545, n52546,
         n52547, n52548, n52549, n52550, n52551, n52552, n52553, n52554,
         n52555, n52556, n52557, n52558, n52559, n52560, n52561, n52562,
         n52563, n52564, n52565, n52566, n52567, n52568, n52569, n52570,
         n52571, n52572, n52573, n52574, n52575, n52576, n52577, n52578,
         n52579, n52580, n52581, n52582, n52583, n52584, n52585, n52586,
         n52587, n52588, n52589, n52590, n52591, n52592, n52593, n52594,
         n52595, n52596, n52597, n52598, n52599, n52600, n52601, n52602,
         n52603, n52604, n52605, n52606, n52607, n52608, n52609, n52610,
         n52611, n52612, n52613, n52614, n52615, n52616, n52617, n52618,
         n52619, n52620, n52621, n52622, n52623, n52624, n52625, n52626,
         n52627, n52628, n52629, n52630, n52631, n52632, n52633, n52634,
         n52635, n52636, n52637, n52638, n52639, n52640, n52641, n52642,
         n52643, n52644, n52645, n52646, n52647, n52648, n52649, n52650,
         n52651, n52652, n52653, n52654, n52655, n52656, n52657, n52658,
         n52659, n52660, n52661, n52662, n52663, n52664, n52665, n52666,
         n52667, n52668, n52669, n52670, n52671, n52672, n52673, n52674,
         n52675, n52676, n52677, n52678, n52679, n52680, n52681, n52682,
         n52683, n52684, n52685, n52686, n52687, n52688, n52689, n52690,
         n52691, n52692, n52693, n52694, n52695, n52696, n52697, n52698,
         n52699, n52700, n52701, n52702, n52703, n52704, n52705, n52706,
         n52707, n52708, n52709, n52710, n52711, n52712, n52713, n52714,
         n52715, n52716, n52717, n52718, n52719, n52720, n52721, n52722,
         n52723, n52724, n52725, n52726, n52727, n52728, n52729, n52730,
         n52731, n52732, n52733, n52734, n52735, n52736, n52737, n52738,
         n52739, n52740, n52741, n52742, n52743, n52744, n52745, n52746,
         n52747, n52748, n52749, n52750, n52751, n52752, n52753, n52754,
         n52755, n52756, n52757, n52758, n52759, n52760, n52761, n52762,
         n52763, n52764, n52765, n52766, n52767, n52768, n52769, n52770,
         n52771, n52772, n52773, n52774, n52775, n52776, n52777, n52778,
         n52779, n52780, n52781, n52782, n52783, n52784, n52785, n52786,
         n52787, n52788, n52789, n52790, n52791, n52792, n52793, n52794,
         n52795, n52796, n52797, n52798, n52799, n52800, n52801, n52802,
         n52803, n52804, n52805, n52806, n52807, n52808, n52809, n52810,
         n52811, n52812, n52813, n52814, n52815, n52816, n52817, n52818,
         n52819, n52820, n52821, n52822, n52823, n52824, n52825, n52826,
         n52827, n52828, n52829, n52830, n52831, n52832, n52833, n52834,
         n52835, n52836, n52837, n52838, n52839, n52840, n52841, n52842,
         n52843, n52844, n52845, n52846, n52847, n52848, n52849, n52850,
         n52851, n52852, n52853, n52854, n52855, n52856, n52857, n52858,
         n52859, n52860, n52861, n52862, n52863, n52864, n52865, n52866,
         n52867, n52868, n52869, n52870, n52871, n52872, n52873, n52874,
         n52875, n52876, n52877, n52878, n52879, n52880, n52881, n52882,
         n52883, n52884, n52885, n52886, n52887, n52888, n52889, n52890,
         n52891, n52892, n52893, n52894, n52895, n52896, n52897, n52898,
         n52899, n52900, n52901, n52902, n52903, n52904, n52905, n52906,
         n52907, n52908, n52909, n52910, n52911, n52912, n52913, n52914,
         n52915, n52916, n52917, n52918, n52919, n52920, n52921, n52922,
         n52923, n52924, n52925, n52926, n52927, n52928, n52929, n52930,
         n52931, n52932, n52933, n52934, n52935, n52936, n52937, n52938,
         n52939, n52940, n52941, n52942, n52943, n52944, n52945, n52946,
         n52947, n52948, n52949, n52950, n52951, n52952, n52953, n52954,
         n52955, n52956, n52957, n52958, n52959, n52960, n52961, n52962,
         n52963, n52964, n52965, n52966, n52967, n52968, n52969, n52970,
         n52971, n52972, n52973, n52974, n52975, n52976, n52977, n52978,
         n52979, n52980, n52981, n52982, n52983, n52984, n52985, n52986,
         n52987, n52988, n52989, n52990, n52991, n52992, n52993, n52994,
         n52995, n52996, n52997, n52998, n52999, n53000, n53001, n53002,
         n53003, n53004, n53005, n53006, n53007, n53008, n53009, n53010,
         n53011, n53012, n53013, n53014, n53015, n53016, n53017, n53018,
         n53019, n53020, n53021, n53022, n53023, n53024, n53025, n53026,
         n53027, n53028, n53029, n53030, n53031, n53032, n53033, n53034,
         n53035, n53036, n53037, n53038, n53039, n53040, n53041, n53042,
         n53043, n53044, n53045, n53046, n53047, n53048, n53049, n53050,
         n53051, n53052, n53053, n53054, n53055, n53056, n53057, n53058,
         n53059, n53060, n53061, n53062, n53063, n53064, n53065, n53066,
         n53067, n53068, n53069, n53070, n53071, n53072, n53073, n53074,
         n53075, n53076, n53077, n53078, n53079, n53080, n53081, n53082,
         n53083, n53084, n53085, n53086, n53087, n53088, n53089, n53090,
         n53091, n53092, n53093, n53094, n53095, n53096, n53097, n53098,
         n53099, n53100, n53101, n53102, n53103, n53104, n53105, n53106,
         n53107, n53108, n53109, n53110, n53111, n53112, n53113, n53114,
         n53115, n53116, n53117, n53118, n53119, n53120, n53121, n53122,
         n53123, n53124, n53125, n53126, n53127, n53128, n53129, n53130,
         n53131, n53132, n53133, n53134, n53135, n53136, n53137, n53138,
         n53139, n53140, n53141, n53142, n53143, n53144, n53145, n53146,
         n53147, n53148, n53149, n53150, n53151, n53152, n53153, n53154,
         n53155, n53156, n53157, n53158, n53159, n53160, n53161, n53162,
         n53163, n53164, n53165, n53166, n53167, n53168, n53169, n53170,
         n53171, n53172, n53173, n53174, n53175, n53176, n53177, n53178,
         n53179, n53180, n53181, n53182, n53183, n53184, n53185, n53186,
         n53187, n53188, n53189, n53190, n53191, n53192, n53193, n53194,
         n53195, n53196, n53197, n53198, n53199, n53200, n53201, n53202,
         n53203, n53204, n53205, n53206, n53207, n53208, n53209, n53210,
         n53211, n53212, n53213, n53214, n53215, n53216, n53217, n53218,
         n53219, n53220, n53221, n53222, n53223, n53224, n53225, n53226,
         n53227, n53228, n53229, n53230, n53231, n53232, n53233, n53234,
         n53235, n53236, n53237, n53238, n53239, n53240, n53241, n53242,
         n53243, n53244, n53245, n53246, n53247, n53248, n53249, n53250,
         n53251, n53252, n53253, n53254, n53255, n53256, n53257, n53258,
         n53259, n53260, n53261, n53262, n53263, n53264, n53265, n53266,
         n53267, n53268, n53269, n53270, n53271, n53272, n53273, n53274,
         n53275, n53276, n53277, n53278, n53279, n53280, n53281, n53282,
         n53283, n53284, n53285, n53286, n53287, n53288, n53289, n53290,
         n53291, n53292, n53293, n53294, n53295, n53296, n53297, n53298,
         n53299, n53300, n53301, n53302, n53303, n53304, n53305, n53306,
         n53307, n53308, n53309, n53310, n53311, n53312, n53313, n53314,
         n53315, n53316, n53317, n53318, n53319, n53320, n53321, n53322,
         n53323, n53324, n53325, n53326, n53327, n53328, n53329, n53330,
         n53331, n53332, n53333, n53334, n53335, n53336, n53337, n53338,
         n53339, n53340, n53341, n53342, n53343, n53344, n53345, n53346,
         n53347, n53348, n53349, n53350, n53351, n53352, n53353, n53354,
         n53355, n53356, n53357, n53358, n53359, n53360, n53361, n53362,
         n53363, n53364, n53365, n53366, n53367, n53368, n53369, n53370,
         n53371, n53372, n53373, n53374, n53375, n53376, n53377, n53378,
         n53379, n53380, n53381, n53382, n53383, n53384, n53385, n53386,
         n53387, n53388, n53389, n53390, n53391, n53392, n53393, n53394,
         n53395, n53396, n53397, n53398, n53399, n53400, n53401, n53402,
         n53403, n53404, n53405, n53406, n53407, n53408, n53409, n53410,
         n53411, n53412, n53413, n53414, n53415, n53416, n53417, n53418,
         n53419, n53420, n53421, n53422, n53423, n53424, n53425, n53426,
         n53427, n53428, n53429, n53430, n53431, n53432, n53433, n53434,
         n53435, n53436, n53437, n53438, n53439, n53440, n53441, n53442,
         n53443, n53444, n53445, n53446, n53447, n53448, n53449, n53450,
         n53451, n53452, n53453, n53454, n53455, n53456, n53457, n53458,
         n53459, n53460, n53461, n53462, n53463, n53464, n53465, n53466,
         n53467, n53468, n53469, n53470, n53471, n53472, n53473, n53474,
         n53475, n53476, n53477, n53478, n53479, n53480, n53481, n53482,
         n53483, n53484, n53485, n53486, n53487, n53488, n53489, n53490,
         n53491, n53492, n53493, n53494, n53495, n53496, n53497, n53498,
         n53499, n53500, n53501, n53502, n53503, n53504, n53505, n53506,
         n53507, n53508, n53509, n53510, n53511, n53512, n53513, n53514,
         n53515, n53516, n53517, n53518, n53519, n53520, n53521, n53522,
         n53523, n53524, n53525, n53526, n53527, n53528, n53529, n53530,
         n53531, n53532, n53533, n53534, n53535, n53536, n53537, n53538,
         n53539, n53540, n53541, n53542, n53543, n53544, n53545, n53546,
         n53547, n53548, n53549, n53550, n53551, n53552, n53553, n53554,
         n53555, n53556, n53557, n53558, n53559, n53560, n53561, n53562,
         n53563, n53564, n53565, n53566, n53567, n53568, n53569, n53570,
         n53571, n53572, n53573, n53574, n53575, n53576, n53577, n53578,
         n53579, n53580, n53581, n53582, n53583, n53584, n53585, n53586,
         n53587, n53588, n53589, n53590, n53591, n53592, n53593, n53594,
         n53595, n53596, n53597, n53598, n53599, n53600, n53601, n53602,
         n53603, n53604, n53605, n53606, n53607, n53608, n53609, n53610,
         n53611, n53612, n53613, n53614, n53615, n53616, n53617, n53618,
         n53619, n53620, n53621, n53622, n53623, n53624, n53625, n53626,
         n53627, n53628, n53629, n53630, n53631, n53632, n53633, n53634,
         n53635, n53636, n53637, n53638, n53639, n53640, n53641, n53642,
         n53643, n53644, n53645, n53646, n53647, n53648, n53649, n53650,
         n53651, n53652, n53653, n53654, n53655, n53656, n53657, n53658,
         n53659, n53660, n53661, n53662, n53663, n53664, n53665, n53666,
         n53667, n53668, n53669, n53670, n53671, n53672, n53673, n53674,
         n53675, n53676, n53677, n53678, n53679, n53680, n53681, n53682,
         n53683, n53684, n53685, n53686, n53687, n53688, n53689, n53690,
         n53691, n53692, n53693, n53694, n53695, n53696, n53697, n53698,
         n53699, n53700, n53701, n53702, n53703, n53704, n53705, n53706,
         n53707, n53708, n53709, n53710, n53711, n53712, n53713, n53714,
         n53715, n53716, n53717, n53718, n53719, n53720, n53721, n53722,
         n53723, n53724, n53725, n53726, n53727, n53728, n53729, n53730,
         n53731, n53732, n53733, n53734, n53735, n53736, n53737, n53738,
         n53739, n53740, n53741, n53742, n53743, n53744, n53745, n53746,
         n53747, n53748, n53749, n53750, n53751, n53752, n53753, n53754,
         n53755, n53756, n53757, n53758, n53759, n53760, n53761, n53762,
         n53763, n53764, n53765, n53766, n53767, n53768, n53769, n53770,
         n53771, n53772, n53773, n53774, n53775, n53776, n53777, n53778,
         n53779, n53780, n53781, n53782, n53783, n53784, n53785, n53786,
         n53787, n53788, n53789, n53790, n53791, n53792, n53793, n53794,
         n53795, n53796, n53797, n53798, n53799, n53800, n53801, n53802,
         n53803, n53804, n53805, n53806, n53807, n53808, n53809, n53810,
         n53811, n53812, n53813, n53814, n53815, n53816, n53817, n53818,
         n53819, n53820, n53821, n53822, n53823, n53824, n53825, n53826,
         n53827, n53828, n53829, n53830, n53831, n53832, n53833, n53834,
         n53835, n53836, n53837, n53838, n53839, n53840, n53841, n53842,
         n53843, n53844, n53845, n53846, n53847, n53848, n53849, n53850,
         n53851, n53852, n53853, n53854, n53855, n53856, n53857, n53858,
         n53859, n53860, n53861, n53862, n53863, n53864, n53865, n53866,
         n53867, n53868, n53869, n53870, n53871, n53872, n53873, n53874,
         n53875, n53876, n53877, n53878, n53879, n53880, n53881, n53882,
         n53883, n53884, n53885, n53886, n53887, n53888, n53889, n53890,
         n53891, n53892, n53893, n53894, n53895, n53896, n53897, n53898,
         n53899, n53900, n53901, n53902, n53903, n53904, n53905, n53906,
         n53907, n53908, n53909, n53910, n53911, n53912, n53913, n53914,
         n53915, n53916, n53917, n53918, n53919, n53920, n53921, n53922,
         n53923, n53924, n53925, n53926, n53927, n53928, n53929, n53930,
         n53931, n53932, n53933, n53934, n53935, n53936, n53937, n53938,
         n53939, n53940, n53941, n53942, n53943, n53944, n53945, n53946,
         n53947, n53948, n53949, n53950, n53951, n53952, n53953, n53954,
         n53955, n53956, n53957, n53958, n53959, n53960, n53961, n53962,
         n53963, n53964, n53965, n53966, n53967, n53968, n53969, n53970,
         n53971, n53972, n53973, n53974, n53975, n53976, n53977, n53978,
         n53979, n53980, n53981, n53982, n53983, n53984, n53985, n53986,
         n53987, n53988, n53989, n53990, n53991, n53992, n53993, n53994,
         n53995, n53996, n53997, n53998, n53999, n54000, n54001, n54002,
         n54003, n54004, n54005, n54006, n54007, n54008, n54009, n54010,
         n54011, n54012, n54013, n54014, n54015, n54016, n54017, n54018,
         n54019, n54020, n54021, n54022, n54023, n54024, n54025, n54026,
         n54027, n54028, n54029, n54030, n54031, n54032, n54033, n54034,
         n54035, n54036, n54037, n54038, n54039, n54040, n54041, n54042,
         n54043, n54044, n54045, n54046, n54047, n54048, n54049, n54050,
         n54051, n54052, n54053, n54054, n54055, n54056, n54057, n54058,
         n54059, n54060, n54061, n54062, n54063, n54064, n54065, n54066,
         n54067, n54068, n54069, n54070, n54071, n54072, n54073, n54074,
         n54075, n54076, n54077, n54078, n54079, n54080, n54081, n54082,
         n54083, n54084, n54085, n54086, n54087, n54088, n54089, n54090,
         n54091, n54092, n54093, n54094, n54095, n54096, n54097, n54098,
         n54099, n54100, n54101, n54102, n54103, n54104, n54105, n54106,
         n54107, n54108, n54109, n54110, n54111, n54112, n54113, n54114,
         n54115, n54116, n54117, n54118, n54119, n54120, n54121, n54122,
         n54123, n54124, n54125, n54126, n54127, n54128, n54129, n54130,
         n54131, n54132, n54133, n54134, n54135, n54136, n54137, n54138,
         n54139, n54140, n54141, n54142, n54143, n54144, n54145, n54146,
         n54147, n54148, n54149, n54150, n54151, n54152, n54153, n54154,
         n54155, n54156, n54157, n54158, n54159, n54160, n54161, n54162,
         n54163, n54164, n54165, n54166, n54167, n54168, n54169, n54170,
         n54171, n54172, n54173, n54174, n54175, n54176, n54177, n54178,
         n54179, n54180, n54181, n54182, n54183, n54184, n54185, n54186,
         n54187, n54188, n54189, n54190, n54191, n54192, n54193, n54194,
         n54195, n54196, n54197, n54198, n54199, n54200, n54201, n54202,
         n54203, n54204, n54205, n54206, n54207, n54208, n54209, n54210,
         n54211, n54212, n54213, n54214, n54215, n54216, n54217, n54218,
         n54219, n54220, n54221, n54222, n54223, n54224, n54225, n54226,
         n54227, n54228, n54229, n54230, n54231, n54232, n54233, n54234,
         n54235, n54236, n54237, n54238, n54239, n54240, n54241, n54242,
         n54243, n54244, n54245, n54246, n54247, n54248, n54249, n54250,
         n54251, n54252, n54253, n54254, n54255, n54256, n54257, n54258,
         n54259, n54260, n54261, n54262, n54263, n54264, n54265, n54266,
         n54267, n54268, n54269, n54270, n54271, n54272, n54273, n54274,
         n54275, n54276, n54277, n54278, n54279, n54280, n54281, n54282,
         n54283, n54284, n54285, n54286, n54287, n54288, n54289, n54290,
         n54291, n54292, n54293, n54294, n54295, n54296, n54297, n54298,
         n54299, n54300, n54301, n54302, n54303, n54304, n54305, n54306,
         n54307, n54308, n54309, n54310, n54311, n54312, n54313, n54314,
         n54315, n54316, n54317, n54318, n54319, n54320, n54321, n54322,
         n54323, n54324, n54325, n54326, n54327, n54328, n54329, n54330,
         n54331, n54332, n54333, n54334, n54335, n54336, n54337, n54338,
         n54339, n54340, n54341, n54342, n54343, n54344, n54345, n54346,
         n54347, n54348, n54349, n54350, n54351, n54352, n54353, n54354,
         n54355, n54356, n54357, n54358, n54359, n54360, n54361, n54362,
         n54363, n54364, n54365, n54366, n54367, n54368, n54369, n54370,
         n54371, n54372, n54373, n54374, n54375, n54376, n54377, n54378,
         n54379, n54380, n54381, n54382, n54383, n54384, n54385, n54386,
         n54387, n54388, n54389, n54390, n54391, n54392, n54393, n54394,
         n54395, n54396, n54397, n54398, n54399, n54400, n54401, n54402,
         n54403, n54404, n54405, n54406, n54407, n54408, n54409, n54410,
         n54411, n54412, n54413, n54414, n54415, n54416, n54417, n54418,
         n54419, n54420, n54421, n54422, n54423, n54424, n54425, n54426,
         n54427, n54428, n54429, n54430, n54431, n54432, n54433, n54434,
         n54435, n54436, n54437, n54438, n54439, n54440, n54441, n54442,
         n54443, n54444, n54445, n54446, n54447, n54448, n54449, n54450,
         n54451, n54452, n54453, n54454, n54455, n54456, n54457, n54458,
         n54459, n54460, n54461, n54462, n54463, n54464, n54465, n54466,
         n54467, n54468, n54469, n54470, n54471, n54472, n54473, n54474,
         n54475, n54476, n54477, n54478, n54479, n54480, n54481, n54482,
         n54483, n54484, n54485, n54486, n54487, n54488, n54489, n54490,
         n54491, n54492, n54493, n54494, n54495, n54496, n54497, n54498,
         n54499, n54500, n54501, n54502, n54503, n54504, n54505, n54506,
         n54507, n54508, n54509, n54510, n54511, n54512, n54513, n54514,
         n54515, n54516, n54517, n54518, n54519, n54520, n54521, n54522,
         n54523, n54524, n54525, n54526, n54527, n54528, n54529, n54530,
         n54531, n54532, n54533, n54534, n54535, n54536, n54537, n54538,
         n54539, n54540, n54541, n54542, n54543, n54544, n54545, n54546,
         n54547, n54548, n54549, n54550, n54551, n54552, n54553, n54554,
         n54555, n54556, n54557, n54558, n54559, n54560, n54561, n54562,
         n54563, n54564, n54565, n54566, n54567, n54568, n54569, n54570,
         n54571, n54572, n54573, n54574, n54575, n54576, n54577, n54578,
         n54579, n54580, n54581, n54582, n54583, n54584, n54585, n54586,
         n54587, n54588, n54589, n54590, n54591, n54592, n54593, n54594,
         n54595, n54596, n54597, n54598, n54599, n54600, n54601, n54602,
         n54603, n54604, n54605, n54606, n54607, n54608, n54609, n54610,
         n54611, n54612, n54613, n54614, n54615, n54616, n54617, n54618,
         n54619, n54620, n54621, n54622, n54623, n54624, n54625, n54626,
         n54627, n54628, n54629, n54630, n54631, n54632, n54633, n54634,
         n54635, n54636, n54637, n54638, n54639, n54640, n54641, n54642,
         n54643, n54644, n54645, n54646, n54647, n54648, n54649, n54650,
         n54651, n54652, n54653, n54654, n54655, n54656, n54657, n54658,
         n54659, n54660, n54661, n54662, n54663, n54664, n54665, n54666,
         n54667, n54668, n54669, n54670, n54671, n54672, n54673, n54674,
         n54675, n54676, n54677, n54678, n54679, n54680, n54681, n54682,
         n54683, n54684, n54685, n54686, n54687, n54688, n54689, n54690,
         n54691, n54692, n54693, n54694, n54695, n54696, n54697, n54698,
         n54699, n54700, n54701, n54702, n54703, n54704, n54705, n54706,
         n54707, n54708, n54709, n54710, n54711, n54712, n54713, n54714,
         n54715, n54716, n54717, n54718, n54719, n54720, n54721, n54722,
         n54723, n54724, n54725, n54726, n54727, n54728, n54729, n54730,
         n54731, n54732, n54733, n54734, n54735, n54736, n54737, n54738,
         n54739, n54740, n54741, n54742, n54743, n54744, n54745, n54746,
         n54747, n54748, n54749, n54750, n54751, n54752, n54753, n54754,
         n54755, n54756, n54757, n54758, n54759, n54760, n54761, n54762,
         n54763, n54764, n54765, n54766, n54767, n54768, n54769, n54770,
         n54771, n54772, n54773, n54774, n54775, n54776, n54777, n54778,
         n54779, n54780, n54781, n54782, n54783, n54784, n54785, n54786,
         n54787, n54788, n54789, n54790, n54791, n54792, n54793, n54794,
         n54795, n54796, n54797, n54798, n54799, n54800, n54801, n54802,
         n54803, n54804, n54805, n54806, n54807, n54808, n54809, n54810,
         n54811, n54812, n54813, n54814, n54815, n54816, n54817, n54818,
         n54819, n54820, n54821, n54822, n54823, n54824, n54825, n54826,
         n54827, n54828, n54829, n54830, n54831, n54832, n54833, n54834,
         n54835, n54836, n54837, n54838, n54839, n54840, n54841, n54842,
         n54843, n54844, n54845, n54846, n54847, n54848, n54849, n54850,
         n54851, n54852, n54853, n54854, n54855, n54856, n54857, n54858,
         n54859, n54860, n54861, n54862, n54863, n54864, n54865, n54866,
         n54867, n54868, n54869, n54870, n54871, n54872, n54873, n54874,
         n54875, n54876, n54877, n54878, n54879, n54880, n54881, n54882,
         n54883, n54884, n54885, n54886, n54887, n54888, n54889, n54890,
         n54891, n54892, n54893, n54894, n54895, n54896, n54897, n54898,
         n54899, n54900, n54901, n54902, n54903, n54904, n54905, n54906,
         n54907, n54908, n54909, n54910, n54911, n54912, n54913, n54914,
         n54915, n54916, n54917, n54918, n54919, n54920, n54921, n54922,
         n54923, n54924, n54925, n54926, n54927, n54928, n54929, n54930,
         n54931, n54932, n54933, n54934, n54935, n54936, n54937, n54938,
         n54939, n54940, n54941, n54942, n54943, n54944, n54945, n54946,
         n54947, n54948, n54949, n54950, n54951, n54952, n54953, n54954,
         n54955, n54956, n54957, n54958, n54959, n54960, n54961, n54962,
         n54963, n54964, n54965, n54966, n54967, n54968, n54969, n54970,
         n54971, n54972, n54973, n54974, n54975, n54976, n54977, n54978,
         n54979, n54980, n54981, n54982, n54983, n54984, n54985, n54986,
         n54987, n54988, n54989, n54990, n54991, n54992, n54993, n54994,
         n54995, n54996, n54997, n54998, n54999, n55000, n55001, n55002,
         n55003, n55004, n55005, n55006, n55007, n55008, n55009, n55010,
         n55011, n55012, n55013, n55014, n55015, n55016, n55017, n55018,
         n55019, n55020, n55021, n55022, n55023, n55024, n55025, n55026,
         n55027, n55028, n55029, n55030, n55031, n55032, n55033, n55034,
         n55035, n55036, n55037, n55038, n55039, n55040, n55041, n55042,
         n55043, n55044, n55045, n55046, n55047, n55048, n55049, n55050,
         n55051, n55052, n55053, n55054, n55055, n55056, n55057, n55058,
         n55059, n55060, n55061, n55062, n55063, n55064, n55065, n55066,
         n55067, n55068, n55069, n55070, n55071, n55072, n55073, n55074,
         n55075, n55076, n55077, n55078, n55079, n55080, n55081, n55082,
         n55083, n55084, n55085, n55086, n55087, n55088, n55089, n55090,
         n55091, n55092, n55093, n55094, n55095, n55096, n55097, n55098,
         n55099, n55100, n55101, n55102, n55103, n55104, n55105, n55106,
         n55107, n55108, n55109, n55110, n55111, n55112, n55113, n55114,
         n55115, n55116, n55117, n55118, n55119, n55120, n55121, n55122,
         n55123, n55124, n55125, n55126, n55127, n55128, n55129, n55130,
         n55131, n55132, n55133, n55134, n55135, n55136, n55137, n55138,
         n55139, n55140, n55141, n55142, n55143, n55144, n55145, n55146,
         n55147, n55148, n55149, n55150, n55151, n55152, n55153, n55154,
         n55155, n55156, n55157, n55158, n55159, n55160, n55161, n55162,
         n55163, n55164, n55165, n55166, n55167, n55168, n55169, n55170,
         n55171, n55172, n55173, n55174, n55175, n55176, n55177, n55178,
         n55179, n55180, n55181, n55182, n55183, n55184, n55185, n55186,
         n55187, n55188, n55189, n55190, n55191, n55192, n55193, n55194,
         n55195, n55196, n55197, n55198, n55199, n55200, n55201, n55202,
         n55203, n55204, n55205, n55206, n55207, n55208, n55209, n55210,
         n55211, n55212, n55213, n55214, n55215, n55216, n55217, n55218,
         n55219, n55220, n55221, n55222, n55223, n55224, n55225, n55226,
         n55227, n55228, n55229, n55230, n55231, n55232, n55233, n55234,
         n55235, n55236, n55237, n55238, n55239, n55240, n55241, n55242,
         n55243, n55244, n55245, n55246, n55247, n55248, n55249, n55250,
         n55251, n55252, n55253, n55254, n55255, n55256, n55257, n55258,
         n55259, n55260, n55261, n55262, n55263, n55264, n55265, n55266,
         n55267, n55268, n55269, n55270, n55271, n55272, n55273, n55274,
         n55275, n55276, n55277, n55278, n55279, n55280, n55281, n55282,
         n55283, n55284, n55285, n55286, n55287, n55288, n55289, n55290,
         n55291, n55292, n55293, n55294, n55295, n55296, n55297, n55298,
         n55299, n55300, n55301, n55302, n55303, n55304, n55305, n55306,
         n55307, n55308, n55309, n55310, n55311, n55312, n55313, n55314,
         n55315, n55316, n55317, n55318, n55319, n55320, n55321, n55322,
         n55323, n55324, n55325, n55326, n55327, n55328, n55329, n55330,
         n55331, n55332, n55333, n55334, n55335, n55336, n55337, n55338,
         n55339, n55340, n55341, n55342, n55343, n55344, n55345, n55346,
         n55347, n55348, n55349, n55350, n55351, n55352, n55353, n55354,
         n55355, n55356, n55357, n55358, n55359, n55360, n55361, n55362,
         n55363, n55364, n55365, n55366, n55367, n55368, n55369, n55370,
         n55371, n55372, n55373, n55374, n55375, n55376, n55377, n55378,
         n55379, n55380, n55381, n55382, n55383, n55384, n55385, n55386,
         n55387, n55388, n55389, n55390, n55391, n55392, n55393, n55394,
         n55395, n55396, n55397, n55398, n55399, n55400, n55401, n55402,
         n55403, n55404, n55405, n55406, n55407, n55408, n55409, n55410,
         n55411, n55412, n55413, n55414, n55415, n55416, n55417, n55418,
         n55419, n55420, n55421, n55422, n55423, n55424, n55425, n55426,
         n55427, n55428, n55429, n55430, n55431, n55432, n55433, n55434,
         n55435, n55436, n55437, n55438, n55439, n55440, n55441, n55442,
         n55443, n55444, n55445, n55446, n55447, n55448, n55449, n55450,
         n55451, n55452, n55453, n55454, n55455, n55456, n55457, n55458,
         n55459, n55460, n55461, n55462, n55463, n55464, n55465, n55466,
         n55467, n55468, n55469, n55470, n55471, n55472, n55473, n55474,
         n55475, n55476, n55477, n55478, n55479, n55480, n55481, n55482,
         n55483, n55484, n55485, n55486, n55487, n55488, n55489, n55490,
         n55491, n55492, n55493, n55494, n55495, n55496, n55497, n55498,
         n55499, n55500, n55501, n55502, n55503, n55504, n55505, n55506,
         n55507, n55508, n55509, n55510, n55511, n55512, n55513, n55514,
         n55515, n55516, n55517, n55518, n55519, n55520, n55521, n55522,
         n55523, n55524, n55525, n55526, n55527, n55528, n55529, n55530,
         n55531, n55532, n55533, n55534, n55535, n55536, n55537, n55538,
         n55539, n55540, n55541, n55542, n55543, n55544, n55545, n55546,
         n55547, n55548, n55549, n55550, n55551, n55552, n55553, n55554,
         n55555, n55556, n55557, n55558, n55559, n55560, n55561, n55562,
         n55563, n55564, n55565, n55566, n55567, n55568, n55569, n55570,
         n55571, n55572, n55573, n55574, n55575, n55576, n55577, n55578,
         n55579, n55580, n55581, n55582, n55583, n55584, n55585, n55586,
         n55587, n55588, n55589, n55590, n55591, n55592, n55593, n55594,
         n55595, n55596, n55597, n55598, n55599, n55600, n55601, n55602,
         n55603, n55604, n55605, n55606, n55607, n55608, n55609, n55610,
         n55611, n55612, n55613, n55614, n55615, n55616, n55617, n55618,
         n55619, n55620, n55621, n55622, n55623, n55624, n55625, n55626,
         n55627, n55628, n55629, n55630, n55631, n55632, n55633, n55634,
         n55635, n55636, n55637, n55638, n55639, n55640, n55641, n55642,
         n55643, n55644, n55645, n55646, n55647, n55648, n55649, n55650,
         n55651, n55652, n55653, n55654, n55655, n55656, n55657, n55658,
         n55659, n55660, n55661, n55662, n55663, n55664, n55665, n55666,
         n55667, n55668, n55669, n55670, n55671, n55672, n55673, n55674,
         n55675, n55676, n55677, n55678, n55679, n55680, n55681, n55682,
         n55683, n55684, n55685, n55686, n55687, n55688, n55689, n55690,
         n55691, n55692, n55693, n55694, n55695, n55696, n55697, n55698,
         n55699, n55700, n55701, n55702, n55703, n55704, n55705, n55706,
         n55707, n55708, n55709, n55710, n55711, n55712, n55713, n55714,
         n55715, n55716, n55717, n55718, n55719, n55720, n55721, n55722,
         n55723, n55724, n55725, n55726, n55727, n55728, n55729, n55730,
         n55731, n55732, n55733, n55734, n55735, n55736, n55737, n55738,
         n55739, n55740, n55741, n55742, n55743, n55744, n55745, n55746,
         n55747, n55748, n55749, n55750, n55751, n55752, n55753, n55754,
         n55755, n55756, n55757, n55758, n55759, n55760, n55761, n55762,
         n55763, n55764, n55765, n55766, n55767, n55768, n55769, n55770,
         n55771, n55772, n55773, n55774, n55775, n55776, n55777, n55778,
         n55779, n55780, n55781, n55782, n55783, n55784, n55785, n55786,
         n55787, n55788, n55789, n55790, n55791, n55792, n55793, n55794,
         n55795, n55796, n55797, n55798, n55799, n55800, n55801, n55802,
         n55803, n55804, n55805, n55806, n55807, n55808, n55809, n55810,
         n55811, n55812, n55813, n55814, n55815, n55816, n55817, n55818,
         n55819, n55820, n55821, n55822, n55823, n55824, n55825, n55826,
         n55827, n55828, n55829, n55830, n55831, n55832, n55833, n55834,
         n55835, n55836, n55837, n55838, n55839, n55840, n55841, n55842,
         n55843, n55844, n55845, n55846, n55847, n55848, n55849, n55850,
         n55851, n55852, n55853, n55854, n55855, n55856, n55857, n55858,
         n55859, n55860, n55861, n55862, n55863, n55864, n55865, n55866,
         n55867, n55868, n55869, n55870, n55871, n55872, n55873, n55874,
         n55875, n55876, n55877, n55878, n55879, n55880, n55881, n55882,
         n55883, n55884, n55885, n55886, n55887, n55888, n55889, n55890,
         n55891, n55892, n55893, n55894, n55895, n55896, n55897, n55898,
         n55899, n55900, n55901, n55902, n55903, n55904, n55905, n55906,
         n55907, n55908, n55909, n55910, n55911, n55912, n55913, n55914,
         n55915, n55916, n55917, n55918, n55919, n55920, n55921, n55922,
         n55923, n55924, n55925, n55926, n55927, n55928, n55929, n55930,
         n55931, n55932, n55933, n55934, n55935, n55936, n55937, n55938,
         n55939, n55940, n55941, n55942, n55943, n55944, n55945, n55946,
         n55947, n55948, n55949, n55950, n55951, n55952, n55953, n55954,
         n55955, n55956, n55957, n55958, n55959, n55960, n55961, n55962,
         n55963, n55964, n55965, n55966, n55967, n55968, n55969, n55970,
         n55971, n55972, n55973, n55974, n55975, n55976, n55977, n55978,
         n55979, n55980, n55981, n55982, n55983, n55984, n55985, n55986,
         n55987, n55988, n55989, n55990, n55991, n55992, n55993, n55994,
         n55995, n55996, n55997, n55998, n55999, n56000, n56001, n56002,
         n56003, n56004, n56005, n56006, n56007, n56008, n56009, n56010,
         n56011, n56012, n56013, n56014, n56015, n56016, n56017, n56018,
         n56019, n56020, n56021, n56022, n56023, n56024, n56025, n56026,
         n56027, n56028, n56029, n56030, n56031, n56032, n56033, n56034,
         n56035, n56036, n56037, n56038, n56039, n56040, n56041, n56042,
         n56043, n56044, n56045, n56046, n56047, n56048, n56049, n56050,
         n56051, n56052, n56053, n56054, n56055, n56056, n56057, n56058,
         n56059, n56060, n56061, n56062, n56063, n56064, n56065, n56066,
         n56067, n56068, n56069, n56070, n56071, n56072, n56073, n56074,
         n56075, n56076, n56077, n56078, n56079, n56080, n56081, n56082,
         n56083, n56084, n56085, n56086, n56087, n56088, n56089, n56090,
         n56091, n56092, n56093, n56094, n56095, n56096, n56097, n56098,
         n56099, n56100, n56101, n56102, n56103, n56104, n56105, n56106,
         n56107, n56108, n56109, n56110, n56111, n56112, n56113, n56114,
         n56115, n56116, n56117, n56118, n56119, n56120, n56121, n56122,
         n56123, n56124, n56125, n56126, n56127, n56128, n56129, n56130,
         n56131, n56132, n56133, n56134, n56135, n56136, n56137, n56138,
         n56139, n56140, n56141, n56142, n56143, n56144, n56145, n56146,
         n56147, n56148, n56149, n56150, n56151, n56152, n56153, n56154,
         n56155, n56156, n56157, n56158, n56159, n56160, n56161, n56162,
         n56163, n56164, n56165, n56166, n56167, n56168, n56169, n56170,
         n56171, n56172, n56173, n56174, n56175, n56176, n56177, n56178,
         n56179, n56180, n56181, n56182, n56183, n56184, n56185, n56186,
         n56187, n56188, n56189, n56190, n56191, n56192, n56193, n56194,
         n56195, n56196, n56197, n56198, n56199, n56200, n56201, n56202,
         n56203, n56204, n56205, n56206, n56207, n56208, n56209, n56210,
         n56211, n56212, n56213, n56214, n56215, n56216, n56217, n56218,
         n56219, n56220, n56221, n56222, n56223, n56224, n56225, n56226,
         n56227, n56228, n56229, n56230, n56231, n56232, n56233, n56234,
         n56235, n56236, n56237, n56238, n56239, n56240, n56241, n56242,
         n56243, n56244, n56245, n56246, n56247, n56248, n56249, n56250,
         n56251, n56252, n56253, n56254, n56255, n56256, n56257, n56258,
         n56259, n56260, n56261, n56262, n56263, n56264, n56265, n56266,
         n56267, n56268, n56269, n56270, n56271, n56272, n56273, n56274,
         n56275, n56276, n56277, n56278, n56279, n56280, n56281, n56282,
         n56283, n56284, n56285, n56286, n56287, n56288, n56289, n56290,
         n56291, n56292, n56293, n56294, n56295, n56296, n56297, n56298,
         n56299, n56300, n56301, n56302, n56303, n56304, n56305, n56306,
         n56307, n56308, n56309, n56310, n56311, n56312, n56313, n56314,
         n56315, n56316, n56317, n56318, n56319, n56320, n56321, n56322,
         n56323, n56324, n56325, n56326, n56327, n56328, n56329, n56330,
         n56331, n56332, n56333, n56334, n56335, n56336, n56337, n56338,
         n56339, n56340, n56341, n56342, n56343, n56344, n56345, n56346,
         n56347, n56348, n56349, n56350, n56351, n56352, n56353, n56354,
         n56355, n56356, n56357, n56358, n56359, n56360, n56361, n56362,
         n56363, n56364, n56365, n56366, n56367, n56368, n56369, n56370,
         n56371, n56372, n56373, n56374, n56375, n56376, n56377, n56378,
         n56379, n56380, n56381, n56382, n56383, n56384, n56385, n56386,
         n56387, n56388, n56389, n56390, n56391, n56392, n56393, n56394,
         n56395, n56396, n56397, n56398, n56399, n56400, n56401, n56402,
         n56403, n56404, n56405, n56406, n56407, n56408, n56409, n56410,
         n56411, n56412, n56413, n56414, n56415, n56416, n56417, n56418,
         n56419, n56420, n56421, n56422, n56423, n56424, n56425, n56426,
         n56427, n56428, n56429, n56430, n56431, n56432, n56433, n56434,
         n56435, n56436, n56437, n56438, n56439, n56440, n56441, n56442,
         n56443, n56444, n56445, n56446, n56447, n56448, n56449, n56450,
         n56451, n56452, n56453, n56454, n56455, n56456, n56457, n56458,
         n56459, n56460, n56461, n56462, n56463, n56464, n56465, n56466,
         n56467, n56468, n56469, n56470, n56471, n56472, n56473, n56474,
         n56475, n56476, n56477, n56478, n56479, n56480, n56481, n56482,
         n56483, n56484, n56485, n56486, n56487, n56488, n56489, n56490,
         n56491, n56492, n56493, n56494, n56495, n56496, n56497, n56498,
         n56499, n56500, n56501, n56502, n56503, n56504, n56505, n56506,
         n56507, n56508, n56509, n56510, n56511, n56512, n56513, n56514,
         n56515, n56516, n56517, n56518, n56519, n56520, n56521, n56522,
         n56523, n56524, n56525, n56526, n56527, n56528, n56529, n56530,
         n56531, n56532, n56533, n56534, n56535, n56536, n56537, n56538,
         n56539, n56540, n56541, n56542, n56543, n56544, n56545, n56546,
         n56547, n56548, n56549, n56550, n56551, n56552, n56553, n56554,
         n56555, n56556, n56557, n56558, n56559, n56560, n56561, n56562,
         n56563, n56564, n56565, n56566, n56567, n56568, n56569, n56570,
         n56571, n56572, n56573, n56574, n56575, n56576, n56577, n56578,
         n56579, n56580, n56581, n56582, n56583, n56584, n56585, n56586,
         n56587, n56588, n56589, n56590, n56591, n56592, n56593, n56594,
         n56595, n56596, n56597, n56598, n56599, n56600, n56601, n56602,
         n56603, n56604, n56605, n56606, n56607, n56608, n56609, n56610,
         n56611, n56612, n56613, n56614, n56615, n56616, n56617, n56618,
         n56619, n56620, n56621, n56622, n56623, n56624, n56625, n56626,
         n56627, n56628, n56629, n56630, n56631, n56632, n56633, n56634,
         n56635, n56636, n56637, n56638, n56639, n56640, n56641, n56642,
         n56643, n56644, n56645, n56646, n56647, n56648, n56649, n56650,
         n56651, n56652, n56653, n56654, n56655, n56656, n56657, n56658,
         n56659, n56660, n56661, n56662, n56663, n56664, n56665, n56666,
         n56667, n56668, n56669, n56670, n56671, n56672, n56673, n56674,
         n56675, n56676, n56677, n56678, n56679, n56680, n56681, n56682,
         n56683, n56684, n56685, n56686, n56687, n56688, n56689, n56690,
         n56691, n56692, n56693, n56694, n56695, n56696, n56697, n56698,
         n56699, n56700, n56701, n56702, n56703, n56704, n56705, n56706,
         n56707, n56708, n56709, n56710, n56711, n56712, n56713, n56714,
         n56715, n56716, n56717, n56718, n56719, n56720, n56721, n56722,
         n56723, n56724, n56725, n56726, n56727, n56728, n56729, n56730,
         n56731, n56732, n56733, n56734, n56735, n56736, n56737, n56738,
         n56739, n56740, n56741, n56742, n56743, n56744, n56745, n56746,
         n56747, n56748, n56749, n56750, n56751, n56752, n56753, n56754,
         n56755, n56756, n56757, n56758, n56759, n56760, n56761, n56762,
         n56763, n56764, n56765, n56766, n56767, n56768, n56769, n56770,
         n56771, n56772, n56773, n56774, n56775, n56776, n56777, n56778,
         n56779, n56780, n56781, n56782, n56783, n56784, n56785, n56786,
         n56787, n56788, n56789, n56790, n56791, n56792, n56793, n56794,
         n56795, n56796, n56797, n56798, n56799, n56800, n56801, n56802,
         n56803, n56804, n56805, n56806, n56807, n56808, n56809, n56810,
         n56811, n56812, n56813, n56814, n56815, n56816, n56817, n56818,
         n56819, n56820, n56821, n56822, n56823, n56824, n56825, n56826,
         n56827, n56828, n56829, n56830, n56831, n56832, n56833, n56834,
         n56835, n56836, n56837, n56838, n56839, n56840, n56841, n56842,
         n56843, n56844, n56845, n56846, n56847, n56848, n56849, n56850,
         n56851, n56852, n56853, n56854, n56855, n56856, n56857, n56858,
         n56859, n56860, n56861, n56862, n56863, n56864, n56865, n56866,
         n56867, n56868, n56869, n56870, n56871, n56872, n56873, n56874,
         n56875, n56876, n56877, n56878, n56879, n56880, n56881, n56882,
         n56883, n56884, n56885, n56886, n56887, n56888, n56889, n56890,
         n56891, n56892, n56893, n56894, n56895, n56896, n56897, n56898,
         n56899, n56900, n56901, n56902, n56903, n56904, n56905, n56906,
         n56907, n56908, n56909, n56910, n56911, n56912, n56913, n56914,
         n56915, n56916, n56917, n56918, n56919, n56920, n56921, n56922,
         n56923, n56924, n56925, n56926, n56927, n56928, n56929, n56930,
         n56931, n56932, n56933, n56934, n56935, n56936, n56937, n56938,
         n56939, n56940, n56941, n56942, n56943, n56944, n56945, n56946,
         n56947, n56948, n56949, n56950, n56951, n56952, n56953, n56954,
         n56955, n56956, n56957, n56958, n56959, n56960, n56961, n56962,
         n56963, n56964, n56965, n56966, n56967, n56968, n56969, n56970,
         n56971, n56972, n56973, n56974, n56975, n56976, n56977, n56978,
         n56979, n56980, n56981, n56982, n56983, n56984, n56985, n56986,
         n56987, n56988, n56989, n56990, n56991, n56992, n56993, n56994,
         n56995, n56996, n56997, n56998, n56999, n57000, n57001, n57002,
         n57003, n57004, n57005, n57006, n57007, n57008, n57009, n57010,
         n57011, n57012, n57013, n57014, n57015, n57016, n57017, n57018,
         n57019, n57020, n57021, n57022, n57023, n57024, n57025, n57026,
         n57027, n57028, n57029, n57030, n57031, n57032, n57033, n57034,
         n57035, n57036, n57037, n57038, n57039, n57040, n57041, n57042,
         n57043, n57044, n57045, n57046, n57047, n57048, n57049, n57050,
         n57051, n57052, n57053, n57054, n57055, n57056, n57057, n57058,
         n57059, n57060, n57061, n57062, n57063, n57064, n57065, n57066,
         n57067, n57068, n57069, n57070, n57071, n57072, n57073, n57074,
         n57075, n57076, n57077, n57078, n57079, n57080, n57081, n57082,
         n57083, n57084, n57085, n57086, n57087, n57088, n57089, n57090,
         n57091, n57092, n57093, n57094, n57095, n57096, n57097, n57098,
         n57099, n57100, n57101, n57102, n57103, n57104, n57105, n57106,
         n57107, n57108, n57109, n57110, n57111, n57112, n57113, n57114,
         n57115, n57116, n57117, n57118, n57119, n57120, n57121, n57122,
         n57123, n57124, n57125, n57126, n57127, n57128, n57129, n57130,
         n57131, n57132, n57133, n57134, n57135, n57136, n57137, n57138,
         n57139, n57140, n57141, n57142, n57143, n57144, n57145, n57146,
         n57147, n57148, n57149, n57150, n57151, n57152, n57153, n57154,
         n57155, n57156, n57157, n57158, n57159, n57160, n57161, n57162,
         n57163, n57164, n57165, n57166, n57167, n57168, n57169, n57170,
         n57171, n57172, n57173, n57174, n57175, n57176, n57177, n57178,
         n57179, n57180, n57181, n57182, n57183, n57184, n57185, n57186,
         n57187, n57188, n57189, n57190, n57191, n57192, n57193, n57194,
         n57195, n57196, n57197, n57198, n57199, n57200, n57201, n57202,
         n57203, n57204, n57205, n57206, n57207, n57208, n57209, n57210,
         n57211, n57212, n57213, n57214, n57215, n57216, n57217, n57218,
         n57219, n57220, n57221, n57222, n57223, n57224, n57225, n57226,
         n57227, n57228, n57229, n57230, n57231, n57232, n57233, n57234,
         n57235, n57236, n57237, n57238, n57239, n57240, n57241, n57242,
         n57243, n57244, n57245, n57246, n57247, n57248, n57249, n57250,
         n57251, n57252, n57253, n57254, n57255, n57256, n57257, n57258,
         n57259, n57260, n57261, n57262, n57263, n57264, n57265, n57266,
         n57267, n57268, n57269, n57270, n57271, n57272, n57273, n57274,
         n57275, n57276, n57277, n57278, n57279, n57280, n57281, n57282,
         n57283, n57284, n57285, n57286, n57287, n57288, n57289, n57290,
         n57291, n57292, n57293, n57294, n57295, n57296, n57297, n57298,
         n57299, n57300, n57301, n57302, n57303, n57304, n57305, n57306,
         n57307, n57308, n57309, n57310, n57311, n57312, n57313, n57314,
         n57315, n57316, n57317, n57318, n57319, n57320, n57321, n57322,
         n57323, n57324, n57325, n57326, n57327, n57328, n57329, n57330,
         n57331, n57332, n57333, n57334, n57335, n57336, n57337, n57338,
         n57339, n57340, n57341, n57342, n57343, n57344, n57345, n57346,
         n57347, n57348, n57349, n57350, n57351, n57352, n57353, n57354,
         n57355, n57356, n57357, n57358, n57359, n57360, n57361, n57362,
         n57363, n57364, n57365, n57366, n57367, n57368, n57369, n57370,
         n57371, n57372, n57373, n57374, n57375, n57376, n57377, n57378,
         n57379, n57380, n57381, n57382, n57383, n57384, n57385, n57386,
         n57387, n57388, n57389, n57390, n57391, n57392, n57393, n57394,
         n57395, n57396, n57397, n57398, n57399, n57400, n57401, n57402,
         n57403, n57404, n57405, n57406, n57407, n57408, n57409, n57410,
         n57411, n57412, n57413, n57414, n57415, n57416, n57417, n57418,
         n57419, n57420, n57421, n57422, n57423, n57424, n57425, n57426,
         n57427, n57428, n57429, n57430, n57431, n57432, n57433, n57434,
         n57435, n57436, n57437, n57438, n57439, n57440, n57441, n57442,
         n57443, n57444, n57445, n57446, n57447, n57448, n57449, n57450,
         n57451, n57452, n57453, n57454, n57455, n57456, n57457, n57458,
         n57459, n57460, n57461, n57462, n57463, n57464, n57465, n57466,
         n57467, n57468, n57469, n57470, n57471, n57472, n57473, n57474,
         n57475, n57476, n57477, n57478, n57479, n57480, n57481, n57482,
         n57483, n57484, n57485, n57486, n57487, n57488, n57489, n57490,
         n57491, n57492, n57493, n57494, n57495, n57496, n57497, n57498,
         n57499, n57500, n57501, n57502, n57503, n57504, n57505, n57506,
         n57507, n57508, n57509, n57510, n57511, n57512, n57513, n57514,
         n57515, n57516, n57517, n57518, n57519, n57520, n57521, n57522,
         n57523, n57524, n57525, n57526, n57527, n57528, n57529, n57530,
         n57531, n57532, n57533, n57534, n57535, n57536, n57537, n57538,
         n57539, n57540, n57541, n57542, n57543, n57544, n57545, n57546,
         n57547, n57548, n57549, n57550, n57551, n57552, n57553, n57554,
         n57555, n57556, n57557, n57558, n57559, n57560, n57561, n57562,
         n57563, n57564, n57565, n57566, n57567, n57568, n57569, n57570,
         n57571, n57572, n57573, n57574, n57575, n57576, n57577, n57578,
         n57579, n57580, n57581, n57582, n57583, n57584, n57585, n57586,
         n57587, n57588, n57589, n57590, n57591, n57592, n57593, n57594,
         n57595, n57596, n57597, n57598, n57599, n57600, n57601, n57602,
         n57603, n57604, n57605, n57606, n57607, n57608, n57609, n57610,
         n57611, n57612, n57613, n57614, n57615, n57616, n57617, n57618,
         n57619, n57620, n57621, n57622, n57623, n57624, n57625, n57626,
         n57627, n57628, n57629, n57630, n57631, n57632, n57633, n57634,
         n57635, n57636, n57637, n57638, n57639, n57640, n57641, n57642,
         n57643, n57644, n57645, n57646, n57647, n57648, n57649, n57650,
         n57651, n57652, n57653, n57654, n57655, n57656, n57657, n57658,
         n57659, n57660, n57661, n57662, n57663, n57664, n57665, n57666,
         n57667, n57668, n57669, n57670, n57671, n57672, n57673, n57674,
         n57675, n57676, n57677, n57678, n57679, n57680, n57681, n57682,
         n57683, n57684, n57685, n57686, n57687, n57688, n57689, n57690,
         n57691, n57692, n57693, n57694, n57695, n57696, n57697, n57698,
         n57699, n57700, n57701, n57702, n57703, n57704, n57705, n57706,
         n57707, n57708, n57709, n57710, n57711, n57712, n57713, n57714,
         n57715, n57716, n57717, n57718, n57719, n57720, n57721, n57722,
         n57723, n57724, n57725, n57726, n57727, n57728, n57729, n57730,
         n57731, n57732, n57733, n57734, n57735, n57736, n57737, n57738,
         n57739, n57740, n57741, n57742, n57743, n57744, n57745, n57746,
         n57747, n57748, n57749, n57750, n57751, n57752, n57753, n57754,
         n57755, n57756, n57757, n57758, n57759, n57760, n57761, n57762,
         n57763, n57764, n57765, n57766, n57767, n57768, n57769, n57770,
         n57771, n57772, n57773, n57774, n57775, n57776, n57777, n57778,
         n57779, n57780, n57781, n57782, n57783, n57784, n57785, n57786,
         n57787, n57788, n57789, n57790, n57791, n57792, n57793, n57794,
         n57795, n57796, n57797, n57798, n57799, n57800, n57801, n57802,
         n57803, n57804, n57805, n57806, n57807, n57808, n57809, n57810,
         n57811, n57812, n57813, n57814, n57815, n57816, n57817, n57818,
         n57819, n57820, n57821, n57822, n57823, n57824, n57825, n57826,
         n57827, n57828, n57829, n57830, n57831, n57832, n57833, n57834,
         n57835, n57836, n57837, n57838, n57839, n57840, n57841, n57842,
         n57843, n57844, n57845, n57846, n57847, n57848, n57849, n57850,
         n57851, n57852, n57853, n57854, n57855, n57856, n57857, n57858,
         n57859, n57860, n57861, n57862, n57863, n57864, n57865, n57866,
         n57867, n57868, n57869, n57870, n57871, n57872, n57873, n57874,
         n57875, n57876, n57877, n57878, n57879, n57880, n57881, n57882,
         n57883, n57884, n57885, n57886, n57887, n57888, n57889, n57890,
         n57891, n57892, n57893, n57894, n57895, n57896, n57897, n57898,
         n57899, n57900, n57901, n57902, n57903, n57904, n57905, n57906,
         n57907, n57908, n57909, n57910, n57911, n57912, n57913, n57914,
         n57915, n57916, n57917, n57918, n57919, n57920, n57921, n57922,
         n57923, n57924, n57925, n57926, n57927, n57928, n57929, n57930,
         n57931, n57932, n57933, n57934, n57935, n57936, n57937, n57938,
         n57939, n57940, n57941, n57942, n57943, n57944, n57945, n57946,
         n57947, n57948, n57949, n57950, n57951, n57952, n57953, n57954,
         n57955, n57956, n57957, n57958, n57959, n57960, n57961, n57962,
         n57963, n57964, n57965, n57966, n57967, n57968, n57969, n57970,
         n57971, n57972, n57973, n57974, n57975, n57976, n57977, n57978,
         n57979, n57980, n57981, n57982, n57983, n57984, n57985, n57986,
         n57987, n57988, n57989, n57990, n57991, n57992, n57993, n57994,
         n57995, n57996, n57997, n57998, n57999, n58000, n58001, n58002,
         n58003, n58004, n58005, n58006, n58007, n58008, n58009, n58010,
         n58011, n58012, n58013, n58014, n58015, n58016, n58017, n58018,
         n58019, n58020, n58021, n58022, n58023, n58024, n58025, n58026,
         n58027, n58028, n58029, n58030, n58031, n58032, n58033, n58034,
         n58035, n58036, n58037, n58038, n58039, n58040, n58041, n58042,
         n58043, n58044, n58045, n58046, n58047, n58048, n58049, n58050,
         n58051, n58052, n58053, n58054, n58055, n58056, n58057, n58058,
         n58059, n58060, n58061, n58062, n58063, n58064, n58065, n58066,
         n58067, n58068, n58069, n58070, n58071, n58072, n58073, n58074,
         n58075, n58076, n58077, n58078, n58079, n58080, n58081, n58082,
         n58083, n58084, n58085, n58086, n58087, n58088, n58089, n58090,
         n58091, n58092, n58093, n58094, n58095, n58096, n58097, n58098,
         n58099, n58100, n58101, n58102, n58103, n58104, n58105, n58106,
         n58107, n58108, n58109, n58110, n58111, n58112, n58113, n58114,
         n58115, n58116, n58117, n58118, n58119, n58120, n58121, n58122,
         n58123, n58124, n58125, n58126, n58127, n58128, n58129, n58130,
         n58131, n58132, n58133, n58134, n58135, n58136, n58137, n58138,
         n58139, n58140, n58141, n58142, n58143, n58144, n58145, n58146,
         n58147, n58148, n58149, n58150, n58151, n58152, n58153, n58154,
         n58155, n58156, n58157, n58158, n58159, n58160, n58161, n58162,
         n58163, n58164, n58165, n58166, n58167, n58168, n58169, n58170,
         n58171, n58172, n58173, n58174, n58175, n58176, n58177, n58178,
         n58179, n58180, n58181, n58182, n58183, n58184, n58185, n58186,
         n58187, n58188, n58189, n58190, n58191, n58192, n58193, n58194,
         n58195, n58196, n58197, n58198, n58199, n58200, n58201, n58202,
         n58203, n58204, n58205, n58206, n58207, n58208, n58209, n58210,
         n58211, n58212, n58213, n58214, n58215, n58216, n58217, n58218,
         n58219, n58220, n58221, n58222, n58223, n58224, n58225, n58226,
         n58227, n58228, n58229, n58230, n58231, n58232, n58233, n58234,
         n58235, n58236, n58237, n58238, n58239, n58240, n58241, n58242,
         n58243, n58244, n58245, n58246, n58247, n58248, n58249, n58250,
         n58251, n58252, n58253, n58254, n58255, n58256, n58257, n58258,
         n58259, n58260, n58261, n58262, n58263, n58264, n58265, n58266,
         n58267, n58268, n58269, n58270, n58271, n58272, n58273, n58274,
         n58275, n58276, n58277, n58278, n58279, n58280, n58281, n58282,
         n58283, n58284, n58285, n58286, n58287, n58288, n58289, n58290,
         n58291, n58292, n58293, n58294, n58295, n58296, n58297, n58298,
         n58299, n58300, n58301, n58302, n58303, n58304, n58305, n58306,
         n58307, n58308, n58309, n58310, n58311, n58312, n58313, n58314,
         n58315, n58316, n58317, n58318, n58319, n58320, n58321, n58322,
         n58323, n58324, n58325, n58326, n58327, n58328, n58329, n58330,
         n58331, n58332, n58333, n58334, n58335, n58336, n58337, n58338,
         n58339, n58340, n58341, n58342, n58343, n58344, n58345, n58346,
         n58347, n58348, n58349, n58350, n58351, n58352, n58353, n58354,
         n58355, n58356, n58357, n58358, n58359, n58360, n58361, n58362,
         n58363, n58364, n58365, n58366, n58367, n58368, n58369, n58370,
         n58371, n58372, n58373, n58374, n58375, n58376, n58377, n58378,
         n58379, n58380, n58381, n58382, n58383, n58384, n58385, n58386,
         n58387, n58388, n58389, n58390, n58391, n58392, n58393, n58394,
         n58395, n58396, n58397, n58398, n58399, n58400, n58401, n58402,
         n58403, n58404, n58405, n58406, n58407, n58408, n58409, n58410,
         n58411, n58412, n58413, n58414, n58415, n58416, n58417, n58418,
         n58419, n58420, n58421, n58422, n58423, n58424, n58425, n58426,
         n58427, n58428, n58429, n58430, n58431, n58432, n58433, n58434,
         n58435, n58436, n58437, n58438, n58439, n58440, n58441, n58442,
         n58443, n58444, n58445, n58446, n58447, n58448, n58449, n58450,
         n58451, n58452, n58453, n58454, n58455, n58456, n58457, n58458,
         n58459, n58460, n58461, n58462, n58463, n58464, n58465, n58466,
         n58467, n58468, n58469, n58470, n58471, n58472, n58473, n58474,
         n58475, n58476, n58477, n58478, n58479, n58480, n58481, n58482,
         n58483, n58484, n58485, n58486, n58487, n58488, n58489, n58490,
         n58491, n58492, n58493, n58494, n58495, n58496, n58497, n58498,
         n58499, n58500, n58501, n58502, n58503, n58504, n58505, n58506,
         n58507, n58508, n58509, n58510, n58511, n58512, n58513, n58514,
         n58515, n58516, n58517, n58518, n58519, n58520, n58521, n58522,
         n58523, n58524, n58525, n58526, n58527, n58528, n58529, n58530,
         n58531, n58532, n58533, n58534, n58535, n58536, n58537, n58538,
         n58539, n58540, n58541, n58542, n58543, n58544, n58545, n58546,
         n58547, n58548, n58549, n58550, n58551, n58552, n58553, n58554,
         n58555, n58556, n58557, n58558, n58559, n58560, n58561, n58562,
         n58563, n58564, n58565, n58566, n58567, n58568, n58569, n58570,
         n58571, n58572, n58573, n58574, n58575, n58576, n58577, n58578,
         n58579, n58580, n58581, n58582, n58583, n58584, n58585, n58586,
         n58587, n58588, n58589, n58590, n58591, n58592, n58593, n58594,
         n58595, n58596, n58597, n58598, n58599, n58600, n58601, n58602,
         n58603, n58604, n58605, n58606, n58607, n58608, n58609, n58610,
         n58611, n58612, n58613, n58614, n58615, n58616, n58617, n58618,
         n58619, n58620, n58621, n58622, n58623, n58624, n58625, n58626,
         n58627, n58628, n58629, n58630, n58631, n58632, n58633, n58634,
         n58635, n58636, n58637, n58638, n58639, n58640, n58641, n58642,
         n58643, n58644, n58645, n58646, n58647, n58648, n58649, n58650,
         n58651, n58652, n58653, n58654, n58655, n58656, n58657, n58658,
         n58659, n58660, n58661, n58662, n58663, n58664, n58665, n58666,
         n58667, n58668, n58669, n58670, n58671, n58672, n58673, n58674,
         n58675, n58676, n58677, n58678, n58679, n58680, n58681, n58682,
         n58683, n58684, n58685, n58686, n58687, n58688, n58689, n58690,
         n58691, n58692, n58693, n58694, n58695, n58696, n58697, n58698,
         n58699, n58700, n58701, n58702, n58703, n58704, n58705, n58706,
         n58707, n58708, n58709, n58710, n58711, n58712, n58713, n58714,
         n58715, n58716, n58717, n58718, n58719, n58720, n58721, n58722,
         n58723, n58724, n58725, n58726, n58727, n58728, n58729, n58730,
         n58731, n58732, n58733, n58734, n58735, n58736, n58737, n58738,
         n58739, n58740, n58741, n58742, n58743, n58744, n58745, n58746,
         n58747, n58748, n58749, n58750, n58751, n58752, n58753, n58754,
         n58755, n58756, n58757, n58758, n58759, n58760, n58761, n58762,
         n58763, n58764, n58765, n58766, n58767, n58768, n58769, n58770,
         n58771, n58772, n58773, n58774, n58775, n58776, n58777, n58778,
         n58779, n58780, n58781, n58782, n58783, n58784, n58785, n58786,
         n58787, n58788, n58789, n58790, n58791, n58792, n58793, n58794,
         n58795, n58796, n58797, n58798, n58799, n58800, n58801, n58802,
         n58803, n58804, n58805, n58806, n58807, n58808, n58809, n58810,
         n58811, n58812, n58813, n58814, n58815, n58816, n58817, n58818,
         n58819, n58820, n58821, n58822, n58823, n58824, n58825, n58826,
         n58827, n58828, n58829, n58830, n58831, n58832, n58833, n58834,
         n58835, n58836, n58837, n58838, n58839, n58840, n58841, n58842,
         n58843, n58844, n58845, n58846, n58847, n58848, n58849, n58850,
         n58851, n58852, n58853, n58854, n58855, n58856, n58857, n58858,
         n58859, n58860, n58861, n58862, n58863, n58864, n58865, n58866,
         n58867, n58868, n58869, n58870, n58871, n58872, n58873, n58874,
         n58875, n58876, n58877, n58878, n58879, n58880, n58881, n58882,
         n58883, n58884, n58885, n58886, n58887, n58888, n58889, n58890,
         n58891, n58892, n58893, n58894, n58895, n58896, n58897, n58898,
         n58899, n58900, n58901, n58902, n58903, n58904, n58905, n58906,
         n58907, n58908, n58909, n58910, n58911, n58912, n58913, n58914,
         n58915, n58916, n58917, n58918, n58919, n58920, n58921, n58922,
         n58923, n58924, n58925, n58926, n58927, n58928, n58929, n58930,
         n58931, n58932, n58933, n58934, n58935, n58936, n58937, n58938,
         n58939, n58940, n58941, n58942, n58943, n58944, n58945, n58946,
         n58947, n58948, n58949, n58950, n58951, n58952, n58953, n58954,
         n58955, n58956, n58957, n58958, n58959, n58960, n58961, n58962,
         n58963, n58964, n58965, n58966, n58967, n58968, n58969, n58970,
         n58971, n58972, n58973, n58974, n58975, n58976, n58977, n58978,
         n58979, n58980, n58981, n58982, n58983, n58984, n58985, n58986,
         n58987, n58988, n58989, n58990, n58991, n58992, n58993, n58994,
         n58995, n58996, n58997, n58998, n58999, n59000, n59001, n59002,
         n59003, n59004, n59005, n59006, n59007, n59008, n59009, n59010,
         n59011, n59012, n59013, n59014, n59015, n59016, n59017, n59018,
         n59019, n59020, n59021, n59022, n59023, n59024, n59025, n59026,
         n59027, n59028, n59029, n59030, n59031, n59032, n59033, n59034,
         n59035, n59036, n59037, n59038, n59039, n59040, n59041, n59042,
         n59043, n59044, n59045, n59046, n59047, n59048, n59049, n59050,
         n59051, n59052, n59053, n59054, n59055, n59056, n59057, n59058,
         n59059, n59060, n59061, n59062, n59063, n59064, n59065, n59066,
         n59067, n59068, n59069, n59070, n59071, n59072, n59073, n59074,
         n59075, n59076, n59077, n59078, n59079, n59080, n59081, n59082,
         n59083, n59084, n59085, n59086, n59087, n59088, n59089, n59090,
         n59091, n59092, n59093, n59094, n59095, n59096, n59097, n59098,
         n59099, n59100, n59101, n59102, n59103, n59104, n59105, n59106,
         n59107, n59108, n59109, n59110, n59111, n59112, n59113, n59114,
         n59115, n59116, n59117, n59118, n59119, n59120, n59121, n59122,
         n59123, n59124, n59125, n59126, n59127, n59128, n59129, n59130,
         n59131, n59132, n59133, n59134, n59135, n59136, n59137, n59138,
         n59139, n59140, n59141, n59142, n59143, n59144, n59145, n59146,
         n59147, n59148, n59149, n59150, n59151, n59152, n59153, n59154,
         n59155, n59156, n59157, n59158, n59159, n59160, n59161, n59162,
         n59163, n59164, n59165, n59166, n59167, n59168, n59169, n59170,
         n59171, n59172, n59173, n59174, n59175, n59176, n59177, n59178,
         n59179, n59180, n59181, n59182, n59183, n59184, n59185, n59186,
         n59187, n59188, n59189, n59190, n59191, n59192, n59193, n59194,
         n59195, n59196, n59197, n59198, n59199, n59200, n59201, n59202,
         n59203, n59204, n59205, n59206, n59207, n59208, n59209, n59210,
         n59211, n59212, n59213, n59214, n59215, n59216, n59217, n59218,
         n59219, n59220, n59221, n59222, n59223, n59224, n59225, n59226,
         n59227, n59228, n59229, n59230, n59231, n59232, n59233, n59234,
         n59235, n59236, n59237, n59238, n59239, n59240, n59241, n59242,
         n59243, n59244, n59245, n59246, n59247, n59248, n59249, n59250,
         n59251, n59252, n59253, n59254, n59255, n59256, n59257, n59258,
         n59259, n59260, n59261, n59262, n59263, n59264, n59265, n59266,
         n59267, n59268, n59269, n59270, n59271, n59272, n59273, n59274,
         n59275, n59276, n59277, n59278, n59279, n59280, n59281, n59282,
         n59283, n59284, n59285, n59286, n59287, n59288, n59289, n59290,
         n59291, n59292, n59293, n59294, n59295, n59296, n59297, n59298,
         n59299, n59300, n59301, n59302, n59303, n59304, n59305, n59306,
         n59307, n59308, n59309, n59310, n59311, n59312, n59313, n59314,
         n59315, n59316, n59317, n59318, n59319, n59320, n59321, n59322,
         n59323, n59324, n59325, n59326, n59327, n59328, n59329, n59330,
         n59331, n59332, n59333, n59334, n59335, n59336, n59337, n59338,
         n59339, n59340, n59341, n59342, n59343, n59344, n59345, n59346,
         n59347, n59348, n59349, n59350, n59351, n59352, n59353, n59354,
         n59355, n59356, n59357, n59358, n59359, n59360, n59361, n59362,
         n59363, n59364, n59365, n59366, n59367, n59368, n59369, n59370,
         n59371, n59372, n59373, n59374, n59375, n59376, n59377, n59378,
         n59379, n59380, n59381, n59382, n59383, n59384, n59385, n59386,
         n59387, n59388, n59389, n59390, n59391, n59392, n59393, n59394,
         n59395, n59396, n59397, n59398, n59399, n59400, n59401, n59402,
         n59403, n59404, n59405, n59406, n59407, n59408, n59409, n59410,
         n59411, n59412, n59413, n59414, n59415, n59416, n59417, n59418,
         n59419, n59420, n59421, n59422, n59423, n59424, n59425, n59426,
         n59427, n59428, n59429, n59430, n59431, n59432, n59433, n59434,
         n59435, n59436, n59437, n59438, n59439, n59440, n59441, n59442,
         n59443, n59444, n59445, n59446, n59447, n59448, n59449, n59450,
         n59451, n59452, n59453, n59454, n59455, n59456, n59457, n59458,
         n59459, n59460, n59461, n59462, n59463, n59464, n59465, n59466,
         n59467, n59468, n59469, n59470, n59471, n59472, n59473, n59474,
         n59475, n59476, n59477, n59478, n59479, n59480, n59481, n59482,
         n59483, n59484, n59485, n59486, n59487, n59488, n59489, n59490,
         n59491, n59492, n59493, n59494, n59495, n59496, n59497, n59498,
         n59499, n59500, n59501, n59502, n59503, n59504, n59505, n59506,
         n59507, n59508, n59509, n59510, n59511, n59512, n59513, n59514,
         n59515, n59516, n59517, n59518, n59519, n59520, n59521, n59522,
         n59523, n59524, n59525, n59526, n59527, n59528, n59529, n59530,
         n59531, n59532, n59533, n59534, n59535, n59536, n59537, n59538,
         n59539, n59540, n59541, n59542, n59543, n59544, n59545, n59546,
         n59547, n59548, n59549, n59550, n59551, n59552, n59553, n59554,
         n59555, n59556, n59557, n59558, n59559, n59560, n59561, n59562,
         n59563, n59564, n59565, n59566, n59567, n59568, n59569, n59570,
         n59571, n59572, n59573, n59574, n59575, n59576, n59577, n59578,
         n59579, n59580, n59581, n59582, n59583, n59584, n59585, n59586,
         n59587, n59588, n59589, n59590, n59591, n59592, n59593, n59594,
         n59595, n59596, n59597, n59598, n59599, n59600, n59601, n59602,
         n59603, n59604, n59605, n59606, n59607, n59608, n59609, n59610,
         n59611, n59612, n59613, n59614, n59615, n59616, n59617, n59618,
         n59619, n59620, n59621, n59622, n59623, n59624, n59625, n59626,
         n59627, n59628, n59629, n59630, n59631, n59632, n59633, n59634,
         n59635, n59636, n59637, n59638, n59639, n59640, n59641, n59642,
         n59643, n59644, n59645, n59646, n59647, n59648, n59649, n59650,
         n59651, n59652, n59653, n59654, n59655, n59656, n59657, n59658,
         n59659, n59660, n59661, n59662, n59663, n59664, n59665, n59666,
         n59667, n59668, n59669, n59670, n59671, n59672, n59673, n59674,
         n59675, n59676, n59677, n59678, n59679, n59680, n59681, n59682,
         n59683, n59684, n59685, n59686, n59687, n59688, n59689, n59690,
         n59691, n59692, n59693, n59694, n59695, n59696, n59697, n59698,
         n59699, n59700, n59701, n59702, n59703, n59704, n59705, n59706,
         n59707, n59708, n59709, n59710, n59711, n59712, n59713, n59714,
         n59715, n59716, n59717, n59718, n59719, n59720, n59721, n59722,
         n59723, n59724, n59725, n59726, n59727, n59728, n59729, n59730,
         n59731, n59732, n59733, n59734, n59735, n59736, n59737, n59738,
         n59739, n59740, n59741, n59742, n59743, n59744, n59745, n59746,
         n59747, n59748, n59749, n59750, n59751, n59752, n59753, n59754,
         n59755, n59756, n59757, n59758, n59759, n59760, n59761, n59762,
         n59763, n59764, n59765, n59766, n59767, n59768, n59769, n59770,
         n59771, n59772, n59773, n59774, n59775, n59776, n59777, n59778,
         n59779, n59780, n59781, n59782, n59783, n59784, n59785, n59786,
         n59787, n59788, n59789, n59790, n59791, n59792, n59793, n59794,
         n59795, n59796, n59797, n59798, n59799, n59800, n59801, n59802,
         n59803, n59804, n59805, n59806, n59807, n59808, n59809, n59810,
         n59811, n59812, n59813, n59814, n59815, n59816, n59817, n59818,
         n59819, n59820, n59821, n59822, n59823, n59824, n59825, n59826,
         n59827, n59828, n59829, n59830, n59831, n59832, n59833, n59834,
         n59835, n59836, n59837, n59838, n59839, n59840, n59841, n59842,
         n59843, n59844, n59845, n59846, n59847, n59848, n59849, n59850,
         n59851, n59852, n59853, n59854, n59855, n59856, n59857, n59858,
         n59859, n59860, n59861, n59862, n59863, n59864, n59865, n59866,
         n59867, n59868, n59869, n59870, n59871, n59872, n59873, n59874,
         n59875, n59876, n59877, n59878, n59879, n59880, n59881, n59882,
         n59883, n59884, n59885, n59886, n59887, n59888, n59889, n59890,
         n59891, n59892, n59893, n59894, n59895, n59896, n59897, n59898,
         n59899, n59900, n59901, n59902, n59903, n59904, n59905, n59906,
         n59907, n59908, n59909, n59910, n59911, n59912, n59913, n59914,
         n59915, n59916, n59917, n59918, n59919, n59920, n59921, n59922,
         n59923, n59924, n59925, n59926, n59927, n59928, n59929, n59930,
         n59931, n59932, n59933, n59934, n59935, n59936, n59937, n59938,
         n59939, n59940, n59941, n59942, n59943, n59944, n59945, n59946,
         n59947, n59948, n59949, n59950, n59951, n59952, n59953, n59954,
         n59955, n59956, n59957, n59958, n59959, n59960, n59961, n59962,
         n59963, n59964, n59965, n59966, n59967, n59968, n59969, n59970,
         n59971, n59972, n59973, n59974, n59975, n59976, n59977, n59978,
         n59979, n59980, n59981, n59982, n59983, n59984, n59985, n59986,
         n59987, n59988, n59989, n59990, n59991, n59992, n59993, n59994,
         n59995, n59996, n59997, n59998, n59999, n60000, n60001, n60002,
         n60003, n60004, n60005, n60006, n60007, n60008, n60009, n60010,
         n60011, n60012, n60013, n60014, n60015, n60016, n60017, n60018,
         n60019, n60020, n60021, n60022, n60023, n60024, n60025, n60026,
         n60027, n60028, n60029, n60030, n60031, n60032, n60033, n60034,
         n60035, n60036, n60037, n60038, n60039, n60040, n60041, n60042,
         n60043, n60044, n60045, n60046, n60047, n60048, n60049, n60050,
         n60051, n60052, n60053, n60054, n60055, n60056, n60057, n60058,
         n60059, n60060, n60061, n60062, n60063, n60064, n60065, n60066,
         n60067, n60068, n60069, n60070, n60071, n60072, n60073, n60074,
         n60075, n60076, n60077, n60078, n60079, n60080, n60081, n60082,
         n60083, n60084, n60085, n60086, n60087, n60088, n60089, n60090,
         n60091, n60092, n60093, n60094, n60095, n60096, n60097, n60098,
         n60099, n60100, n60101, n60102, n60103, n60104, n60105, n60106,
         n60107, n60108, n60109, n60110, n60111, n60112, n60113, n60114,
         n60115, n60116, n60117, n60118, n60119, n60120, n60121, n60122,
         n60123, n60124, n60125, n60126, n60127, n60128, n60129, n60130,
         n60131, n60132, n60133, n60134, n60135, n60136, n60137, n60138,
         n60139, n60140, n60141, n60142, n60143, n60144, n60145, n60146,
         n60147, n60148, n60149, n60150, n60151, n60152, n60153, n60154,
         n60155, n60156, n60157, n60158, n60159, n60160, n60161, n60162,
         n60163, n60164, n60165, n60166, n60167, n60168, n60169, n60170,
         n60171, n60172, n60173, n60174, n60175, n60176, n60177, n60178,
         n60179, n60180, n60181, n60182, n60183, n60184, n60185, n60186,
         n60187, n60188, n60189, n60190, n60191, n60192, n60193, n60194,
         n60195, n60196, n60197, n60198, n60199, n60200, n60201, n60202,
         n60203, n60204, n60205, n60206, n60207, n60208, n60209, n60210,
         n60211, n60212, n60213, n60214, n60215, n60216, n60217, n60218,
         n60219, n60220, n60221, n60222, n60223, n60224, n60225, n60226,
         n60227, n60228, n60229, n60230, n60231, n60232, n60233, n60234,
         n60235, n60236, n60237, n60238, n60239, n60240, n60241, n60242,
         n60243, n60244, n60245, n60246, n60247, n60248, n60249, n60250,
         n60251, n60252, n60253, n60254, n60255, n60256, n60257, n60258,
         n60259, n60260, n60261, n60262, n60263, n60264, n60265, n60266,
         n60267, n60268, n60269, n60270, n60271, n60272, n60273, n60274,
         n60275, n60276, n60277, n60278, n60279, n60280, n60281, n60282,
         n60283, n60284, n60285, n60286, n60287, n60288, n60289, n60290,
         n60291, n60292, n60293, n60294, n60295, n60296, n60297, n60298,
         n60299, n60300, n60301, n60302, n60303, n60304, n60305, n60306,
         n60307, n60308, n60309, n60310, n60311, n60312, n60313, n60314,
         n60315, n60316, n60317, n60318, n60319, n60320, n60321, n60322,
         n60323, n60324, n60325, n60326, n60327, n60328, n60329, n60330,
         n60331, n60332, n60333, n60334, n60335, n60336, n60337, n60338,
         n60339, n60340, n60341, n60342, n60343, n60344, n60345, n60346,
         n60347, n60348, n60349, n60350, n60351, n60352, n60353, n60354,
         n60355, n60356, n60357, n60358, n60359, n60360, n60361, n60362,
         n60363, n60364, n60365, n60366, n60367, n60368, n60369, n60370,
         n60371, n60372, n60373, n60374, n60375, n60376, n60377, n60378,
         n60379, n60380, n60381, n60382, n60383, n60384, n60385, n60386,
         n60387, n60388, n60389, n60390, n60391, n60392, n60393, n60394,
         n60395, n60396, n60397, n60398, n60399, n60400, n60401, n60402,
         n60403, n60404, n60405, n60406, n60407, n60408, n60409, n60410,
         n60411, n60412, n60413, n60414, n60415, n60416, n60417, n60418,
         n60419, n60420, n60421, n60422, n60423, n60424, n60425, n60426,
         n60427, n60428, n60429, n60430, n60431, n60432, n60433, n60434,
         n60435, n60436, n60437, n60438, n60439, n60440, n60441, n60442,
         n60443, n60444, n60445, n60446, n60447, n60448, n60449, n60450,
         n60451, n60452, n60453, n60454, n60455, n60456, n60457, n60458,
         n60459, n60460, n60461, n60462, n60463, n60464, n60465, n60466,
         n60467, n60468, n60469, n60470, n60471, n60472, n60473, n60474,
         n60475, n60476, n60477, n60478, n60479, n60480, n60481, n60482,
         n60483, n60484, n60485, n60486, n60487, n60488, n60489, n60490,
         n60491, n60492, n60493, n60494, n60495, n60496, n60497, n60498,
         n60499, n60500, n60501, n60502, n60503, n60504, n60505, n60506,
         n60507, n60508, n60509, n60510, n60511, n60512, n60513, n60514,
         n60515, n60516, n60517, n60518, n60519, n60520, n60521, n60522,
         n60523, n60524, n60525, n60526, n60527, n60528, n60529, n60530,
         n60531, n60532, n60533, n60534, n60535, n60536, n60537, n60538,
         n60539, n60540, n60541, n60542, n60543, n60544, n60545, n60546,
         n60547, n60548, n60549, n60550, n60551, n60552, n60553, n60554,
         n60555, n60556, n60557, n60558, n60559, n60560, n60561, n60562,
         n60563, n60564, n60565, n60566, n60567, n60568, n60569, n60570,
         n60571, n60572, n60573, n60574, n60575, n60576, n60577, n60578,
         n60579, n60580, n60581, n60582, n60583, n60584, n60585, n60586,
         n60587, n60588, n60589, n60590, n60591, n60592, n60593, n60594,
         n60595, n60596, n60597, n60598, n60599, n60600, n60601, n60602,
         n60603, n60604, n60605, n60606, n60607, n60608, n60609, n60610,
         n60611, n60612, n60613, n60614, n60615, n60616, n60617, n60618,
         n60619, n60620, n60621, n60622, n60623, n60624, n60625, n60626,
         n60627, n60628, n60629, n60630, n60631, n60632, n60633, n60634,
         n60635, n60636, n60637, n60638, n60639, n60640, n60641, n60642,
         n60643, n60644, n60645, n60646, n60647, n60648, n60649, n60650,
         n60651, n60652, n60653, n60654, n60655, n60656, n60657, n60658,
         n60659, n60660, n60661, n60662, n60663, n60664, n60665, n60666,
         n60667, n60668, n60669, n60670, n60671, n60672, n60673, n60674,
         n60675, n60676, n60677, n60678, n60679, n60680, n60681, n60682,
         n60683, n60684, n60685, n60686, n60687, n60688, n60689, n60690,
         n60691, n60692, n60693, n60694, n60695, n60696, n60697, n60698,
         n60699, n60700, n60701, n60702, n60703, n60704, n60705, n60706,
         n60707, n60708, n60709, n60710, n60711, n60712, n60713, n60714,
         n60715, n60716, n60717, n60718, n60719, n60720, n60721, n60722,
         n60723, n60724, n60725, n60726, n60727, n60728, n60729, n60730,
         n60731, n60732, n60733, n60734, n60735, n60736, n60737, n60738,
         n60739, n60740, n60741, n60742, n60743, n60744, n60745, n60746,
         n60747, n60748, n60749, n60750, n60751, n60752, n60753, n60754,
         n60755, n60756, n60757, n60758, n60759, n60760, n60761, n60762,
         n60763, n60764, n60765, n60766, n60767, n60768, n60769, n60770,
         n60771, n60772, n60773, n60774, n60775, n60776, n60777, n60778,
         n60779, n60780, n60781, n60782, n60783, n60784, n60785, n60786,
         n60787, n60788, n60789, n60790, n60791, n60792, n60793, n60794,
         n60795, n60796, n60797, n60798, n60799, n60800, n60801, n60802,
         n60803, n60804, n60805, n60806, n60807, n60808, n60809, n60810,
         n60811, n60812, n60813, n60814, n60815, n60816, n60817, n60818,
         n60819, n60820, n60821, n60822, n60823, n60824, n60825, n60826,
         n60827, n60828, n60829, n60830, n60831, n60832, n60833, n60834,
         n60835, n60836, n60837, n60838, n60839, n60840, n60841, n60842,
         n60843, n60844, n60845, n60846, n60847, n60848, n60849, n60850,
         n60851, n60852, n60853, n60854, n60855, n60856, n60857, n60858,
         n60859, n60860, n60861, n60862, n60863, n60864, n60865, n60866,
         n60867, n60868, n60869, n60870, n60871, n60872, n60873, n60874,
         n60875, n60876, n60877, n60878, n60879, n60880, n60881, n60882,
         n60883, n60884, n60885, n60886, n60887, n60888, n60889, n60890,
         n60891, n60892, n60893, n60894, n60895, n60896, n60897, n60898,
         n60899, n60900, n60901, n60902, n60903, n60904, n60905, n60906,
         n60907, n60908, n60909, n60910, n60911, n60912, n60913, n60914,
         n60915, n60916, n60917, n60918, n60919, n60920, n60921, n60922,
         n60923, n60924, n60925, n60926, n60927, n60928, n60929, n60930,
         n60931, n60932, n60933, n60934, n60935, n60936, n60937, n60938,
         n60939, n60940, n60941, n60942, n60943, n60944, n60945, n60946,
         n60947, n60948, n60949, n60950, n60951, n60952, n60953, n60954,
         n60955, n60956, n60957, n60958, n60959, n60960, n60961, n60962,
         n60963, n60964, n60965, n60966, n60967, n60968, n60969, n60970,
         n60971, n60972, n60973, n60974, n60975, n60976, n60977, n60978,
         n60979, n60980, n60981, n60982, n60983, n60984, n60985, n60986,
         n60987, n60988, n60989, n60990, n60991, n60992, n60993, n60994,
         n60995, n60996, n60997, n60998, n60999, n61000, n61001, n61002,
         n61003, n61004, n61005, n61006, n61007, n61008, n61009, n61010,
         n61011, n61012, n61013, n61014, n61015, n61016, n61017, n61018,
         n61019, n61020, n61021, n61022, n61023, n61024, n61025, n61026,
         n61027, n61028, n61029, n61030, n61031, n61032, n61033, n61034,
         n61035, n61036, n61037, n61038, n61039, n61040, n61041, n61042,
         n61043, n61044, n61045, n61046, n61047, n61048, n61049, n61050,
         n61051, n61052, n61053, n61054, n61055, n61056, n61057, n61058,
         n61059, n61060, n61061, n61062, n61063, n61064, n61065, n61066,
         n61067, n61068, n61069, n61070, n61071, n61072, n61073, n61074,
         n61075, n61076, n61077, n61078, n61079, n61080, n61081, n61082,
         n61083, n61084, n61085, n61086, n61087, n61088, n61089, n61090,
         n61091, n61092, n61093, n61094, n61095, n61096, n61097, n61098,
         n61099, n61100, n61101, n61102, n61103, n61104, n61105, n61106,
         n61107, n61108, n61109, n61110, n61111, n61112, n61113, n61114,
         n61115, n61116, n61117, n61118, n61119, n61120, n61121, n61122,
         n61123, n61124, n61125, n61126, n61127, n61128, n61129, n61130,
         n61131, n61132, n61133, n61134, n61135, n61136, n61137, n61138,
         n61139, n61140, n61141, n61142, n61143, n61144, n61145, n61146,
         n61147, n61148, n61149, n61150, n61151, n61152, n61153, n61154,
         n61155, n61156, n61157, n61158, n61159, n61160, n61161, n61162,
         n61163, n61164, n61165, n61166, n61167, n61168, n61169, n61170,
         n61171, n61172, n61173, n61174, n61175, n61176, n61177, n61178,
         n61179, n61180, n61181, n61182, n61183, n61184, n61185, n61186,
         n61187, n61188, n61189, n61190, n61191, n61192, n61193, n61194,
         n61195, n61196, n61197, n61198, n61199, n61200, n61201, n61202,
         n61203, n61204, n61205, n61206, n61207, n61208, n61209, n61210,
         n61211, n61212, n61213, n61214, n61215, n61216, n61217, n61218,
         n61219, n61220, n61221, n61222, n61223, n61224, n61225, n61226,
         n61227, n61228, n61229, n61230, n61231, n61232, n61233, n61234,
         n61235, n61236, n61237, n61238, n61239, n61240, n61241, n61242,
         n61243, n61244, n61245, n61246, n61247, n61248, n61249, n61250,
         n61251, n61252, n61253, n61254, n61255, n61256, n61257, n61258,
         n61259, n61260, n61261, n61262, n61263, n61264, n61265, n61266,
         n61267, n61268, n61269, n61270, n61271, n61272, n61273, n61274,
         n61275, n61276, n61277, n61278, n61279, n61280, n61281, n61282,
         n61283;

  DFF ebreg_reg ( .D(n5), .CLK(clk), .RST(rst), .Q(ebreg) );
  DFF greg_reg ( .D(n4), .CLK(clk), .RST(rst), .Q(g) );
  ANDN U10 ( .B(n28359), .A(n28358), .Z(n52447) );
  ANDN U11 ( .B(n28346), .A(n28345), .Z(n52464) );
  NANDN U12 ( .A(n28327), .B(n28328), .Z(n52482) );
  ANDN U13 ( .B(n28311), .A(n28310), .Z(n52500) );
  ANDN U14 ( .B(n28296), .A(n28295), .Z(n52515) );
  ANDN U15 ( .B(n28032), .A(n28031), .Z(n53204) );
  ANDN U16 ( .B(n28012), .A(n28011), .Z(n53234) );
  ANDN U17 ( .B(n27999), .A(n27998), .Z(n53260) );
  ANDN U18 ( .B(n27984), .A(n27983), .Z(n53288) );
  NANDN U19 ( .A(n27966), .B(n27967), .Z(n53316) );
  NANDN U20 ( .A(n27960), .B(n27961), .Z(n53327) );
  ANDN U21 ( .B(n27882), .A(n27881), .Z(n53454) );
  NANDN U22 ( .A(x[1422]), .B(y[1422]), .Z(n8) );
  ANDN U23 ( .B(n8), .A(n33075), .Z(n53495) );
  NOR U24 ( .A(n33097), .B(n33098), .Z(n53507) );
  ANDN U25 ( .B(n27773), .A(n27772), .Z(n53586) );
  NOR U26 ( .A(n33419), .B(n33420), .Z(n53627) );
  ANDN U27 ( .B(n27703), .A(n27702), .Z(n53701) );
  NOR U28 ( .A(n27634), .B(n27635), .Z(n53816) );
  XNOR U29 ( .A(y[1808]), .B(x[1808]), .Z(n9) );
  NAND U30 ( .A(n27541), .B(n9), .Z(n53937) );
  NANDN U31 ( .A(n27524), .B(n27525), .Z(n53951) );
  NANDN U32 ( .A(n27501), .B(n27502), .Z(n53996) );
  NANDN U33 ( .A(n27466), .B(n27467), .Z(n54025) );
  ANDN U34 ( .B(n27454), .A(n27453), .Z(n54041) );
  ANDN U35 ( .B(n34337), .A(n34336), .Z(n54070) );
  NANDN U36 ( .A(n27348), .B(n27349), .Z(n54154) );
  NANDN U37 ( .A(n27300), .B(n27299), .Z(n10) );
  NAND U38 ( .A(n27301), .B(n10), .Z(n11) );
  NANDN U39 ( .A(n27302), .B(n11), .Z(n54238) );
  NANDN U40 ( .A(x[2148]), .B(y[2148]), .Z(n12) );
  ANDN U41 ( .B(n12), .A(n27264), .Z(n54309) );
  ANDN U42 ( .B(n27218), .A(n27217), .Z(n54415) );
  NANDN U43 ( .A(x[2270]), .B(y[2270]), .Z(n13) );
  NANDN U44 ( .A(n27202), .B(n13), .Z(n54437) );
  ANDN U45 ( .B(n35398), .A(n35397), .Z(n54501) );
  ANDN U46 ( .B(n27091), .A(n27090), .Z(n54558) );
  NOR U47 ( .A(n35577), .B(n35578), .Z(n54572) );
  ANDN U48 ( .B(n27054), .A(n27053), .Z(n54631) );
  ANDN U49 ( .B(n35880), .A(n35879), .Z(n54688) );
  ANDN U50 ( .B(n26953), .A(n26952), .Z(n54753) );
  ANDN U51 ( .B(n25082), .A(n25081), .Z(n56729) );
  ANDN U52 ( .B(n28357), .A(n28356), .Z(n52449) );
  ANDN U53 ( .B(n28342), .A(n28341), .Z(n52467) );
  ANDN U54 ( .B(n28335), .A(n28334), .Z(n52475) );
  ANDN U55 ( .B(n28318), .A(n28317), .Z(n52492) );
  ANDN U56 ( .B(n28294), .A(n28293), .Z(n52521) );
  NOR U57 ( .A(n28271), .B(n28272), .Z(n52597) );
  NOR U58 ( .A(n28179), .B(n28180), .Z(n52882) );
  NOR U59 ( .A(n31479), .B(n31480), .Z(n52889) );
  ANDN U60 ( .B(n28153), .A(n28152), .Z(n52923) );
  ANDN U61 ( .B(n28114), .A(n28113), .Z(n53026) );
  ANDN U62 ( .B(n28089), .A(n28088), .Z(n53090) );
  NANDN U63 ( .A(n28065), .B(n28066), .Z(n53150) );
  NANDN U64 ( .A(n28029), .B(n28030), .Z(n53205) );
  NOR U65 ( .A(n32413), .B(n32414), .Z(n53235) );
  NANDN U66 ( .A(n27996), .B(n27997), .Z(n53261) );
  ANDN U67 ( .B(n27982), .A(n27981), .Z(n53290) );
  NANDN U68 ( .A(n27962), .B(n27963), .Z(n53318) );
  NANDN U69 ( .A(n53437), .B(n53436), .Z(n14) );
  NAND U70 ( .A(n53439), .B(n14), .Z(n15) );
  AND U71 ( .A(n53440), .B(n15), .Z(n16) );
  OR U72 ( .A(n52288), .B(n16), .Z(n17) );
  NAND U73 ( .A(n52287), .B(n17), .Z(n18) );
  NANDN U74 ( .A(n53441), .B(n18), .Z(n19) );
  NAND U75 ( .A(n53442), .B(n19), .Z(n20) );
  NAND U76 ( .A(n53443), .B(n20), .Z(n21) );
  ANDN U77 ( .B(n21), .A(n52286), .Z(n22) );
  OR U78 ( .A(n53444), .B(n22), .Z(n23) );
  AND U79 ( .A(n53445), .B(n23), .Z(n24) );
  NANDN U80 ( .A(n24), .B(n53446), .Z(n25) );
  NANDN U81 ( .A(n53447), .B(n25), .Z(n26) );
  NAND U82 ( .A(n53448), .B(n26), .Z(n53451) );
  ANDN U83 ( .B(n27867), .A(n27866), .Z(n53469) );
  NOR U84 ( .A(n27842), .B(n27843), .Z(n53497) );
  ANDN U85 ( .B(n27833), .A(n27832), .Z(n53514) );
  ANDN U86 ( .B(n27814), .A(n27813), .Z(n53532) );
  ANDN U87 ( .B(n27788), .A(n27787), .Z(n53568) );
  ANDN U88 ( .B(n27771), .A(n27770), .Z(n53587) );
  NANDN U89 ( .A(n27764), .B(n27765), .Z(n53596) );
  ANDN U90 ( .B(n27739), .A(n27738), .Z(n53628) );
  NAND U91 ( .A(n53689), .B(n53690), .Z(n27) );
  NANDN U92 ( .A(n53692), .B(n27), .Z(n28) );
  AND U93 ( .A(n53693), .B(n28), .Z(n29) );
  OR U94 ( .A(n53694), .B(n29), .Z(n30) );
  NANDN U95 ( .A(n53695), .B(n30), .Z(n31) );
  NAND U96 ( .A(n53696), .B(n31), .Z(n32) );
  NANDN U97 ( .A(n53697), .B(n32), .Z(n33) );
  NANDN U98 ( .A(n53698), .B(n33), .Z(n34) );
  AND U99 ( .A(n53699), .B(n34), .Z(n35) );
  OR U100 ( .A(n52246), .B(n35), .Z(n36) );
  NAND U101 ( .A(n53700), .B(n36), .Z(n37) );
  NAND U102 ( .A(n53701), .B(n37), .Z(n38) );
  NAND U103 ( .A(n53702), .B(n38), .Z(n39) );
  NANDN U104 ( .A(n53703), .B(n39), .Z(n40) );
  AND U105 ( .A(n53704), .B(n40), .Z(n41) );
  NANDN U106 ( .A(n41), .B(n53705), .Z(n42) );
  NANDN U107 ( .A(n53706), .B(n42), .Z(n43) );
  NAND U108 ( .A(n53707), .B(n43), .Z(n44) );
  NAND U109 ( .A(n53708), .B(n44), .Z(n53709) );
  ANDN U110 ( .B(n27691), .A(n27690), .Z(n53740) );
  NOR U111 ( .A(n27683), .B(n27684), .Z(n53746) );
  NANDN U112 ( .A(n27630), .B(n27631), .Z(n53818) );
  ANDN U113 ( .B(n27609), .A(n27608), .Z(n53838) );
  NANDN U114 ( .A(n27600), .B(n27601), .Z(n45) );
  NAND U115 ( .A(n27602), .B(n45), .Z(n46) );
  ANDN U116 ( .B(n46), .A(n27603), .Z(n53845) );
  ANDN U117 ( .B(n27589), .A(n27588), .Z(n53861) );
  NANDN U118 ( .A(n27578), .B(n27579), .Z(n53881) );
  NOR U119 ( .A(n33954), .B(n33955), .Z(n53894) );
  ANDN U120 ( .B(n27565), .A(n27564), .Z(n53902) );
  ANDN U121 ( .B(n27540), .A(n27539), .Z(n53938) );
  ANDN U122 ( .B(n27523), .A(n27522), .Z(n53952) );
  ANDN U123 ( .B(n27516), .A(n27515), .Z(n53967) );
  ANDN U124 ( .B(n27508), .A(n27507), .Z(n53987) );
  NANDN U125 ( .A(n27505), .B(n27506), .Z(n53994) );
  NANDN U126 ( .A(n27462), .B(n27463), .Z(n54027) );
  ANDN U127 ( .B(n27452), .A(n27451), .Z(n54042) );
  ANDN U128 ( .B(n27431), .A(n27430), .Z(n54071) );
  ANDN U129 ( .B(n27406), .A(n27405), .Z(n52170) );
  ANDN U130 ( .B(n27362), .A(n27361), .Z(n54141) );
  ANDN U131 ( .B(n27347), .A(n27346), .Z(n54155) );
  NANDN U132 ( .A(n34734), .B(n34735), .Z(n54252) );
  ANDN U133 ( .B(n34914), .A(n34913), .Z(n54310) );
  NANDN U134 ( .A(n27240), .B(n27241), .Z(n47) );
  NAND U135 ( .A(n27242), .B(n47), .Z(n48) );
  AND U136 ( .A(n27243), .B(n48), .Z(n52129) );
  NAND U137 ( .A(n54423), .B(n54422), .Z(n49) );
  NAND U138 ( .A(n54424), .B(n49), .Z(n50) );
  ANDN U139 ( .B(n50), .A(n52116), .Z(n51) );
  OR U140 ( .A(n51), .B(n54425), .Z(n52) );
  NAND U141 ( .A(n54426), .B(n52), .Z(n53) );
  NANDN U142 ( .A(n54427), .B(n53), .Z(n54) );
  NAND U143 ( .A(n54428), .B(n54), .Z(n55) );
  NANDN U144 ( .A(n52115), .B(n55), .Z(n56) );
  ANDN U145 ( .B(n56), .A(n54429), .Z(n57) );
  NANDN U146 ( .A(n57), .B(n54430), .Z(n58) );
  NANDN U147 ( .A(n54431), .B(n58), .Z(n59) );
  NAND U148 ( .A(n54432), .B(n59), .Z(n60) );
  NAND U149 ( .A(n54433), .B(n60), .Z(n61) );
  NANDN U150 ( .A(n54434), .B(n61), .Z(n62) );
  AND U151 ( .A(n54435), .B(n62), .Z(n54436) );
  NAND U152 ( .A(n54466), .B(n54467), .Z(n63) );
  NAND U153 ( .A(n54470), .B(n63), .Z(n64) );
  NANDN U154 ( .A(n54471), .B(n64), .Z(n65) );
  NAND U155 ( .A(n54472), .B(n65), .Z(n66) );
  NANDN U156 ( .A(n52109), .B(n66), .Z(n67) );
  AND U157 ( .A(n52108), .B(n67), .Z(n68) );
  ANDN U158 ( .B(n52106), .A(n52105), .Z(n69) );
  OR U159 ( .A(n52107), .B(n68), .Z(n70) );
  AND U160 ( .A(n69), .B(n70), .Z(n71) );
  OR U161 ( .A(n71), .B(n54473), .Z(n72) );
  AND U162 ( .A(n54474), .B(n72), .Z(n73) );
  OR U163 ( .A(n73), .B(n54475), .Z(n74) );
  NAND U164 ( .A(n54476), .B(n74), .Z(n75) );
  NANDN U165 ( .A(n54477), .B(n75), .Z(n54478) );
  NANDN U166 ( .A(n27140), .B(n27141), .Z(n54502) );
  NANDN U167 ( .A(n54534), .B(n54533), .Z(n76) );
  NANDN U168 ( .A(n54535), .B(n76), .Z(n77) );
  AND U169 ( .A(n54536), .B(n77), .Z(n78) );
  OR U170 ( .A(n78), .B(n54537), .Z(n79) );
  NAND U171 ( .A(n54538), .B(n79), .Z(n80) );
  ANDN U172 ( .B(n80), .A(n54539), .Z(n81) );
  OR U173 ( .A(n81), .B(n54540), .Z(n82) );
  NAND U174 ( .A(n54541), .B(n82), .Z(n83) );
  NANDN U175 ( .A(n54542), .B(n83), .Z(n84) );
  NAND U176 ( .A(n54543), .B(n84), .Z(n85) );
  NANDN U177 ( .A(n54544), .B(n85), .Z(n86) );
  ANDN U178 ( .B(n86), .A(n54545), .Z(n87) );
  NANDN U179 ( .A(n87), .B(n54546), .Z(n88) );
  NANDN U180 ( .A(n52092), .B(n88), .Z(n89) );
  NAND U181 ( .A(n52091), .B(n89), .Z(n90) );
  ANDN U182 ( .B(n90), .A(n54547), .Z(n54550) );
  ANDN U183 ( .B(n27084), .A(n27083), .Z(n54575) );
  NAND U184 ( .A(n35604), .B(n35603), .Z(n91) );
  ANDN U185 ( .B(n91), .A(n35605), .Z(n54584) );
  ANDN U186 ( .B(n27058), .A(n27057), .Z(n54629) );
  NAND U187 ( .A(n54670), .B(n54671), .Z(n92) );
  NANDN U188 ( .A(n54672), .B(n92), .Z(n93) );
  NAND U189 ( .A(n54673), .B(n93), .Z(n94) );
  NANDN U190 ( .A(n54674), .B(n94), .Z(n95) );
  NAND U191 ( .A(n54675), .B(n95), .Z(n96) );
  AND U192 ( .A(n54676), .B(n96), .Z(n97) );
  OR U193 ( .A(n54677), .B(n97), .Z(n98) );
  NAND U194 ( .A(n54678), .B(n98), .Z(n99) );
  NANDN U195 ( .A(n54679), .B(n99), .Z(n100) );
  NAND U196 ( .A(n54680), .B(n100), .Z(n101) );
  NANDN U197 ( .A(n54681), .B(n101), .Z(n102) );
  AND U198 ( .A(n54682), .B(n102), .Z(n103) );
  OR U199 ( .A(n54683), .B(n103), .Z(n104) );
  NAND U200 ( .A(n54684), .B(n104), .Z(n105) );
  NAND U201 ( .A(n54685), .B(n105), .Z(n106) );
  NAND U202 ( .A(n54686), .B(n106), .Z(n54687) );
  ANDN U203 ( .B(n26984), .A(n26983), .Z(n52062) );
  ANDN U204 ( .B(n36006), .A(n36005), .Z(n54729) );
  ANDN U205 ( .B(n26969), .A(n26968), .Z(n54738) );
  ANDN U206 ( .B(n26949), .A(n26948), .Z(n54755) );
  NAND U207 ( .A(n55150), .B(n55151), .Z(n107) );
  NANDN U208 ( .A(n55152), .B(n107), .Z(n108) );
  NANDN U209 ( .A(n55153), .B(n108), .Z(n109) );
  NAND U210 ( .A(n55154), .B(n109), .Z(n110) );
  NAND U211 ( .A(n55155), .B(n110), .Z(n111) );
  ANDN U212 ( .B(n111), .A(n51989), .Z(n112) );
  NANDN U213 ( .A(n112), .B(n51988), .Z(n113) );
  NANDN U214 ( .A(n55156), .B(n113), .Z(n114) );
  NAND U215 ( .A(n55157), .B(n114), .Z(n115) );
  NAND U216 ( .A(n55158), .B(n115), .Z(n116) );
  NANDN U217 ( .A(n55159), .B(n116), .Z(n117) );
  AND U218 ( .A(n55160), .B(n117), .Z(n118) );
  NANDN U219 ( .A(n118), .B(n55161), .Z(n119) );
  AND U220 ( .A(n55162), .B(n119), .Z(n120) );
  OR U221 ( .A(n120), .B(n55163), .Z(n121) );
  NAND U222 ( .A(n55164), .B(n121), .Z(n122) );
  NANDN U223 ( .A(n55165), .B(n122), .Z(n55168) );
  NANDN U224 ( .A(x[3496]), .B(y[3496]), .Z(n123) );
  ANDN U225 ( .B(n123), .A(n26039), .Z(n51877) );
  ANDN U226 ( .B(n25727), .A(n25726), .Z(n56051) );
  NANDN U227 ( .A(x[3952]), .B(y[3952]), .Z(n124) );
  ANDN U228 ( .B(n124), .A(n25571), .Z(n51753) );
  AND U229 ( .A(n56246), .B(n56245), .Z(n56247) );
  AND U230 ( .A(n56723), .B(n56722), .Z(n56724) );
  AND U231 ( .A(n56839), .B(n56838), .Z(n56840) );
  ANDN U232 ( .B(n24965), .A(n24964), .Z(n56919) );
  NAND U233 ( .A(n56955), .B(n56954), .Z(n125) );
  ANDN U234 ( .B(n125), .A(n56957), .Z(n126) );
  ANDN U235 ( .B(n51577), .A(n126), .Z(n127) );
  NAND U236 ( .A(n51578), .B(n127), .Z(n128) );
  NANDN U237 ( .A(n56958), .B(n128), .Z(n129) );
  NAND U238 ( .A(n56959), .B(n129), .Z(n130) );
  NANDN U239 ( .A(n56960), .B(n130), .Z(n131) );
  AND U240 ( .A(n56961), .B(n131), .Z(n132) );
  AND U241 ( .A(n51575), .B(n51576), .Z(n133) );
  NANDN U242 ( .A(n132), .B(n56962), .Z(n134) );
  AND U243 ( .A(n133), .B(n134), .Z(n135) );
  ANDN U244 ( .B(n56965), .A(n56964), .Z(n136) );
  NANDN U245 ( .A(n135), .B(n56963), .Z(n137) );
  AND U246 ( .A(n136), .B(n137), .Z(n138) );
  OR U247 ( .A(n56966), .B(n138), .Z(n139) );
  AND U248 ( .A(n56967), .B(n139), .Z(n140) );
  NANDN U249 ( .A(n56968), .B(n140), .Z(n141) );
  NAND U250 ( .A(n56969), .B(n141), .Z(n142) );
  NANDN U251 ( .A(n56970), .B(n142), .Z(n56971) );
  ANDN U252 ( .B(n24825), .A(n24824), .Z(n57095) );
  NAND U253 ( .A(n57125), .B(n57126), .Z(n143) );
  ANDN U254 ( .B(n143), .A(n51545), .Z(n144) );
  ANDN U255 ( .B(n51544), .A(n144), .Z(n145) );
  NAND U256 ( .A(n57127), .B(n145), .Z(n146) );
  NANDN U257 ( .A(n57128), .B(n146), .Z(n147) );
  AND U258 ( .A(n57129), .B(n57130), .Z(n148) );
  NAND U259 ( .A(n147), .B(n148), .Z(n149) );
  NANDN U260 ( .A(n57131), .B(n149), .Z(n150) );
  AND U261 ( .A(n57133), .B(n57132), .Z(n151) );
  NAND U262 ( .A(n150), .B(n151), .Z(n152) );
  NAND U263 ( .A(n57134), .B(n152), .Z(n153) );
  AND U264 ( .A(n57135), .B(n57136), .Z(n154) );
  NAND U265 ( .A(n153), .B(n154), .Z(n155) );
  NANDN U266 ( .A(n57137), .B(n155), .Z(n156) );
  NAND U267 ( .A(n57138), .B(n156), .Z(n57141) );
  NAND U268 ( .A(n57282), .B(n57283), .Z(n157) );
  NAND U269 ( .A(n57284), .B(n157), .Z(n158) );
  NAND U270 ( .A(n57285), .B(n158), .Z(n159) );
  NAND U271 ( .A(n57286), .B(n159), .Z(n160) );
  AND U272 ( .A(n57288), .B(n160), .Z(n161) );
  NAND U273 ( .A(n161), .B(n57287), .Z(n162) );
  NAND U274 ( .A(n57289), .B(n162), .Z(n163) );
  NANDN U275 ( .A(n57290), .B(n163), .Z(n164) );
  AND U276 ( .A(n57291), .B(n164), .Z(n165) );
  OR U277 ( .A(n165), .B(n57292), .Z(n166) );
  NAND U278 ( .A(n57293), .B(n166), .Z(n167) );
  ANDN U279 ( .B(n167), .A(n51514), .Z(n168) );
  NANDN U280 ( .A(n168), .B(n51513), .Z(n169) );
  NANDN U281 ( .A(n57294), .B(n169), .Z(n170) );
  NAND U282 ( .A(n57295), .B(n170), .Z(n57296) );
  ANDN U283 ( .B(n57360), .A(n57361), .Z(n57362) );
  ANDN U284 ( .B(n57539), .A(n57540), .Z(n57541) );
  ANDN U285 ( .B(n57586), .A(n57585), .Z(n171) );
  NAND U286 ( .A(n57584), .B(n57583), .Z(n172) );
  AND U287 ( .A(n171), .B(n172), .Z(n173) );
  NANDN U288 ( .A(n173), .B(n51446), .Z(n174) );
  ANDN U289 ( .B(n174), .A(n57587), .Z(n175) );
  ANDN U290 ( .B(n51444), .A(n51445), .Z(n176) );
  NANDN U291 ( .A(n175), .B(n57588), .Z(n177) );
  AND U292 ( .A(n176), .B(n177), .Z(n178) );
  ANDN U293 ( .B(n57590), .A(n57591), .Z(n179) );
  NANDN U294 ( .A(n178), .B(n57589), .Z(n180) );
  AND U295 ( .A(n179), .B(n180), .Z(n181) );
  NANDN U296 ( .A(n181), .B(n51443), .Z(n182) );
  NANDN U297 ( .A(n57592), .B(n182), .Z(n183) );
  NAND U298 ( .A(n57593), .B(n183), .Z(n57594) );
  NAND U299 ( .A(n57656), .B(n57655), .Z(n184) );
  NANDN U300 ( .A(n57659), .B(n184), .Z(n185) );
  NANDN U301 ( .A(n57660), .B(n185), .Z(n186) );
  NAND U302 ( .A(n57661), .B(n186), .Z(n187) );
  NANDN U303 ( .A(n51432), .B(n187), .Z(n188) );
  AND U304 ( .A(n51431), .B(n188), .Z(n189) );
  ANDN U305 ( .B(n57664), .A(n57663), .Z(n190) );
  OR U306 ( .A(n57662), .B(n189), .Z(n191) );
  AND U307 ( .A(n190), .B(n191), .Z(n192) );
  OR U308 ( .A(n57665), .B(n192), .Z(n193) );
  NAND U309 ( .A(n57666), .B(n193), .Z(n194) );
  NANDN U310 ( .A(n51430), .B(n194), .Z(n57667) );
  AND U311 ( .A(n57757), .B(n57758), .Z(n195) );
  NAND U312 ( .A(n57759), .B(n195), .Z(n196) );
  NAND U313 ( .A(n57760), .B(n196), .Z(n197) );
  ANDN U314 ( .B(n51399), .A(n51398), .Z(n198) );
  NAND U315 ( .A(n197), .B(n198), .Z(n199) );
  NANDN U316 ( .A(n57761), .B(n199), .Z(n200) );
  AND U317 ( .A(n57762), .B(n57763), .Z(n201) );
  NAND U318 ( .A(n200), .B(n201), .Z(n202) );
  NAND U319 ( .A(n51397), .B(n202), .Z(n203) );
  NANDN U320 ( .A(n57764), .B(n203), .Z(n204) );
  NAND U321 ( .A(n57765), .B(n204), .Z(n205) );
  AND U322 ( .A(n51395), .B(n205), .Z(n206) );
  NANDN U323 ( .A(n51396), .B(n206), .Z(n57768) );
  ANDN U324 ( .B(n57850), .A(n57851), .Z(n207) );
  OR U325 ( .A(n57848), .B(n57849), .Z(n208) );
  AND U326 ( .A(n207), .B(n208), .Z(n209) );
  ANDN U327 ( .B(n51380), .A(n51379), .Z(n210) );
  OR U328 ( .A(n209), .B(n57852), .Z(n211) );
  AND U329 ( .A(n210), .B(n211), .Z(n212) );
  ANDN U330 ( .B(n57855), .A(n57854), .Z(n213) );
  NANDN U331 ( .A(n212), .B(n57853), .Z(n214) );
  AND U332 ( .A(n213), .B(n214), .Z(n215) );
  ANDN U333 ( .B(n57858), .A(n57857), .Z(n216) );
  OR U334 ( .A(n57856), .B(n215), .Z(n217) );
  AND U335 ( .A(n216), .B(n217), .Z(n218) );
  ANDN U336 ( .B(n57860), .A(n57861), .Z(n219) );
  OR U337 ( .A(n57859), .B(n218), .Z(n220) );
  AND U338 ( .A(n219), .B(n220), .Z(n221) );
  ANDN U339 ( .B(n51378), .A(n51377), .Z(n222) );
  OR U340 ( .A(n221), .B(n57862), .Z(n223) );
  NAND U341 ( .A(n222), .B(n223), .Z(n57863) );
  AND U342 ( .A(n57919), .B(n57918), .Z(n57920) );
  AND U343 ( .A(n58030), .B(n51340), .Z(n224) );
  NAND U344 ( .A(n51341), .B(n224), .Z(n225) );
  NANDN U345 ( .A(n58031), .B(n225), .Z(n226) );
  NAND U346 ( .A(n58032), .B(n226), .Z(n227) );
  NANDN U347 ( .A(n58033), .B(n227), .Z(n228) );
  AND U348 ( .A(n58034), .B(n228), .Z(n229) );
  OR U349 ( .A(n58035), .B(n229), .Z(n230) );
  NAND U350 ( .A(n58036), .B(n230), .Z(n231) );
  NANDN U351 ( .A(n58037), .B(n231), .Z(n232) );
  AND U352 ( .A(n58038), .B(n58039), .Z(n233) );
  NAND U353 ( .A(n232), .B(n233), .Z(n234) );
  NANDN U354 ( .A(n58040), .B(n234), .Z(n235) );
  NAND U355 ( .A(n58041), .B(n235), .Z(n236) );
  AND U356 ( .A(n51339), .B(n51338), .Z(n237) );
  NANDN U357 ( .A(n58042), .B(n236), .Z(n238) );
  NAND U358 ( .A(n237), .B(n238), .Z(n58043) );
  NAND U359 ( .A(n58120), .B(n58121), .Z(n239) );
  ANDN U360 ( .B(n239), .A(n58122), .Z(n240) );
  ANDN U361 ( .B(n58124), .A(n240), .Z(n241) );
  NAND U362 ( .A(n58123), .B(n241), .Z(n242) );
  NAND U363 ( .A(n58125), .B(n242), .Z(n243) );
  AND U364 ( .A(n51315), .B(n51316), .Z(n244) );
  NAND U365 ( .A(n243), .B(n244), .Z(n245) );
  NAND U366 ( .A(n58126), .B(n245), .Z(n246) );
  NANDN U367 ( .A(n51314), .B(n246), .Z(n247) );
  NAND U368 ( .A(n51313), .B(n247), .Z(n248) );
  AND U369 ( .A(n58127), .B(n248), .Z(n249) );
  NAND U370 ( .A(n249), .B(n51312), .Z(n250) );
  NAND U371 ( .A(n58128), .B(n250), .Z(n251) );
  AND U372 ( .A(n58129), .B(n251), .Z(n252) );
  NAND U373 ( .A(n58130), .B(n252), .Z(n58133) );
  NAND U374 ( .A(n58335), .B(n58334), .Z(n253) );
  NAND U375 ( .A(n58336), .B(n253), .Z(n254) );
  NAND U376 ( .A(n58337), .B(n254), .Z(n255) );
  NAND U377 ( .A(n58338), .B(n255), .Z(n256) );
  AND U378 ( .A(n58340), .B(n256), .Z(n257) );
  NAND U379 ( .A(n257), .B(n58339), .Z(n258) );
  NAND U380 ( .A(n51259), .B(n258), .Z(n259) );
  AND U381 ( .A(n58341), .B(n259), .Z(n260) );
  NAND U382 ( .A(n260), .B(n58342), .Z(n261) );
  AND U383 ( .A(n58344), .B(n58345), .Z(n262) );
  NANDN U384 ( .A(n58343), .B(n261), .Z(n263) );
  NAND U385 ( .A(n262), .B(n263), .Z(n264) );
  AND U386 ( .A(n51257), .B(n51258), .Z(n265) );
  NANDN U387 ( .A(n58346), .B(n264), .Z(n266) );
  NAND U388 ( .A(n265), .B(n266), .Z(n267) );
  NAND U389 ( .A(n58347), .B(n267), .Z(n268) );
  AND U390 ( .A(n58349), .B(n268), .Z(n269) );
  NAND U391 ( .A(n269), .B(n58348), .Z(n58350) );
  NAND U392 ( .A(n58492), .B(n58491), .Z(n270) );
  ANDN U393 ( .B(n270), .A(n58493), .Z(n271) );
  ANDN U394 ( .B(n51223), .A(n271), .Z(n272) );
  NAND U395 ( .A(n51222), .B(n272), .Z(n273) );
  ANDN U396 ( .B(n273), .A(n58494), .Z(n274) );
  NANDN U397 ( .A(n274), .B(n58495), .Z(n275) );
  NAND U398 ( .A(n51221), .B(n275), .Z(n276) );
  NAND U399 ( .A(n58496), .B(n276), .Z(n277) );
  NANDN U400 ( .A(n277), .B(n58497), .Z(n278) );
  ANDN U401 ( .B(n278), .A(n58498), .Z(n279) );
  ANDN U402 ( .B(n51220), .A(n279), .Z(n280) );
  NAND U403 ( .A(n51219), .B(n280), .Z(n281) );
  ANDN U404 ( .B(n281), .A(n58499), .Z(n282) );
  NANDN U405 ( .A(n282), .B(n58500), .Z(n283) );
  NANDN U406 ( .A(n58501), .B(n283), .Z(n284) );
  NAND U407 ( .A(n58502), .B(n284), .Z(n285) );
  AND U408 ( .A(n51218), .B(n51217), .Z(n286) );
  NANDN U409 ( .A(n58503), .B(n285), .Z(n287) );
  NAND U410 ( .A(n286), .B(n287), .Z(n58506) );
  AND U411 ( .A(n58550), .B(n58549), .Z(n58551) );
  AND U412 ( .A(n58753), .B(n58754), .Z(n288) );
  NANDN U413 ( .A(n58752), .B(n58751), .Z(n289) );
  AND U414 ( .A(n288), .B(n289), .Z(n290) );
  OR U415 ( .A(n51158), .B(n290), .Z(n291) );
  NAND U416 ( .A(n51157), .B(n291), .Z(n292) );
  NAND U417 ( .A(n58755), .B(n292), .Z(n293) );
  AND U418 ( .A(n58756), .B(n58757), .Z(n294) );
  NAND U419 ( .A(n293), .B(n294), .Z(n295) );
  NAND U420 ( .A(n51156), .B(n295), .Z(n296) );
  AND U421 ( .A(n58758), .B(n58759), .Z(n297) );
  NAND U422 ( .A(n296), .B(n297), .Z(n298) );
  NANDN U423 ( .A(n58760), .B(n298), .Z(n299) );
  AND U424 ( .A(n58761), .B(n58762), .Z(n300) );
  NAND U425 ( .A(n299), .B(n300), .Z(n301) );
  NANDN U426 ( .A(n58763), .B(n301), .Z(n58764) );
  AND U427 ( .A(n51140), .B(n51141), .Z(n302) );
  OR U428 ( .A(n58803), .B(n58804), .Z(n303) );
  NAND U429 ( .A(n302), .B(n303), .Z(n304) );
  NAND U430 ( .A(n58805), .B(n304), .Z(n305) );
  AND U431 ( .A(n58806), .B(n305), .Z(n306) );
  NANDN U432 ( .A(n51139), .B(n306), .Z(n307) );
  NAND U433 ( .A(n51138), .B(n307), .Z(n308) );
  AND U434 ( .A(n58808), .B(n308), .Z(n309) );
  NAND U435 ( .A(n309), .B(n58807), .Z(n310) );
  ANDN U436 ( .B(n58811), .A(n58810), .Z(n311) );
  NANDN U437 ( .A(n58809), .B(n310), .Z(n312) );
  NAND U438 ( .A(n311), .B(n312), .Z(n313) );
  NAND U439 ( .A(n58812), .B(n313), .Z(n314) );
  AND U440 ( .A(n51137), .B(n314), .Z(n315) );
  NANDN U441 ( .A(n51136), .B(n315), .Z(n58813) );
  AND U442 ( .A(n51120), .B(n51121), .Z(n316) );
  AND U443 ( .A(n58855), .B(n51122), .Z(n317) );
  NAND U444 ( .A(n51123), .B(n317), .Z(n318) );
  NANDN U445 ( .A(n58856), .B(n318), .Z(n319) );
  AND U446 ( .A(n58858), .B(n58857), .Z(n320) );
  NAND U447 ( .A(n319), .B(n320), .Z(n321) );
  NANDN U448 ( .A(n58859), .B(n321), .Z(n322) );
  AND U449 ( .A(n58861), .B(n58860), .Z(n323) );
  NAND U450 ( .A(n322), .B(n323), .Z(n324) );
  NAND U451 ( .A(n58862), .B(n324), .Z(n325) );
  NOR U452 ( .A(n58864), .B(n58863), .Z(n326) );
  NAND U453 ( .A(n325), .B(n326), .Z(n327) );
  NAND U454 ( .A(n58865), .B(n327), .Z(n328) );
  NAND U455 ( .A(n316), .B(n328), .Z(n58868) );
  AND U456 ( .A(n58915), .B(n58914), .Z(n329) );
  OR U457 ( .A(n58912), .B(n58913), .Z(n330) );
  NAND U458 ( .A(n329), .B(n330), .Z(n331) );
  NAND U459 ( .A(n58916), .B(n331), .Z(n332) );
  AND U460 ( .A(n51110), .B(n332), .Z(n333) );
  NANDN U461 ( .A(n51109), .B(n333), .Z(n334) );
  NAND U462 ( .A(n58917), .B(n334), .Z(n335) );
  AND U463 ( .A(n58918), .B(n335), .Z(n336) );
  NAND U464 ( .A(n336), .B(n58919), .Z(n337) );
  AND U465 ( .A(n58921), .B(n58922), .Z(n338) );
  NANDN U466 ( .A(n58920), .B(n337), .Z(n339) );
  NAND U467 ( .A(n338), .B(n339), .Z(n340) );
  AND U468 ( .A(n58925), .B(n58924), .Z(n341) );
  NANDN U469 ( .A(n58923), .B(n340), .Z(n342) );
  NAND U470 ( .A(n341), .B(n342), .Z(n343) );
  NAND U471 ( .A(n58926), .B(n343), .Z(n58927) );
  NAND U472 ( .A(n59031), .B(n59032), .Z(n344) );
  ANDN U473 ( .B(n51081), .A(n51080), .Z(n345) );
  NANDN U474 ( .A(n59033), .B(n344), .Z(n346) );
  NAND U475 ( .A(n345), .B(n346), .Z(n347) );
  ANDN U476 ( .B(n51078), .A(n51079), .Z(n348) );
  NANDN U477 ( .A(n59034), .B(n347), .Z(n349) );
  NAND U478 ( .A(n348), .B(n349), .Z(n350) );
  ANDN U479 ( .B(n59036), .A(n59035), .Z(n351) );
  NANDN U480 ( .A(n51077), .B(n350), .Z(n352) );
  NAND U481 ( .A(n351), .B(n352), .Z(n353) );
  NAND U482 ( .A(n59037), .B(n353), .Z(n354) );
  AND U483 ( .A(n59039), .B(n354), .Z(n355) );
  NAND U484 ( .A(n355), .B(n59038), .Z(n356) );
  AND U485 ( .A(n51076), .B(n51075), .Z(n357) );
  NANDN U486 ( .A(n59040), .B(n356), .Z(n358) );
  NAND U487 ( .A(n357), .B(n358), .Z(n59043) );
  ANDN U488 ( .B(n59395), .A(n50995), .Z(n359) );
  NAND U489 ( .A(n50996), .B(n359), .Z(n360) );
  AND U490 ( .A(n59396), .B(n360), .Z(n361) );
  NANDN U491 ( .A(n361), .B(n59397), .Z(n362) );
  NANDN U492 ( .A(n59398), .B(n362), .Z(n363) );
  NAND U493 ( .A(n59399), .B(n363), .Z(n364) );
  NAND U494 ( .A(n59400), .B(n364), .Z(n365) );
  AND U495 ( .A(n59401), .B(n365), .Z(n366) );
  NAND U496 ( .A(n366), .B(n59402), .Z(n367) );
  NAND U497 ( .A(n59403), .B(n367), .Z(n368) );
  AND U498 ( .A(n59404), .B(n368), .Z(n369) );
  NAND U499 ( .A(n369), .B(n59405), .Z(n370) );
  NAND U500 ( .A(n59406), .B(n370), .Z(n371) );
  AND U501 ( .A(n50993), .B(n371), .Z(n372) );
  NAND U502 ( .A(n372), .B(n50994), .Z(n373) );
  NAND U503 ( .A(n59407), .B(n373), .Z(n374) );
  AND U504 ( .A(n59409), .B(n374), .Z(n375) );
  NAND U505 ( .A(n375), .B(n59408), .Z(n376) );
  NANDN U506 ( .A(n59410), .B(n376), .Z(n59411) );
  AND U507 ( .A(n59597), .B(n59599), .Z(n377) );
  NAND U508 ( .A(n59598), .B(n377), .Z(n378) );
  AND U509 ( .A(n59600), .B(n378), .Z(n379) );
  NOR U510 ( .A(n59601), .B(n379), .Z(n380) );
  NAND U511 ( .A(n59602), .B(n380), .Z(n381) );
  ANDN U512 ( .B(n381), .A(n59603), .Z(n382) );
  NOR U513 ( .A(n50949), .B(n50950), .Z(n383) );
  NANDN U514 ( .A(n382), .B(n383), .Z(n384) );
  AND U515 ( .A(n59604), .B(n384), .Z(n385) );
  NOR U516 ( .A(n59605), .B(n385), .Z(n386) );
  NAND U517 ( .A(n59606), .B(n386), .Z(n387) );
  AND U518 ( .A(n59607), .B(n387), .Z(n388) );
  ANDN U519 ( .B(n50948), .A(n388), .Z(n389) );
  NAND U520 ( .A(n50947), .B(n389), .Z(n390) );
  AND U521 ( .A(n59608), .B(n390), .Z(n391) );
  NANDN U522 ( .A(n391), .B(n59609), .Z(n392) );
  ANDN U523 ( .B(n392), .A(n59610), .Z(n59611) );
  NAND U524 ( .A(n59819), .B(n59820), .Z(n393) );
  ANDN U525 ( .B(n393), .A(n59823), .Z(n394) );
  NANDN U526 ( .A(n59822), .B(n394), .Z(n395) );
  ANDN U527 ( .B(n59826), .A(n59825), .Z(n396) );
  NANDN U528 ( .A(n59824), .B(n395), .Z(n397) );
  NAND U529 ( .A(n396), .B(n397), .Z(n398) );
  NAND U530 ( .A(n59827), .B(n398), .Z(n399) );
  AND U531 ( .A(n59829), .B(n399), .Z(n400) );
  NAND U532 ( .A(n400), .B(n59828), .Z(n401) );
  NAND U533 ( .A(n59830), .B(n401), .Z(n402) );
  AND U534 ( .A(n59832), .B(n402), .Z(n403) );
  NANDN U535 ( .A(n59831), .B(n403), .Z(n404) );
  NAND U536 ( .A(n59833), .B(n404), .Z(n405) );
  AND U537 ( .A(n50886), .B(n405), .Z(n406) );
  NANDN U538 ( .A(n50885), .B(n406), .Z(n407) );
  NAND U539 ( .A(n59834), .B(n407), .Z(n408) );
  AND U540 ( .A(n59836), .B(n408), .Z(n409) );
  NANDN U541 ( .A(n59835), .B(n409), .Z(n410) );
  NANDN U542 ( .A(n59837), .B(n410), .Z(n59838) );
  NAND U543 ( .A(n60520), .B(n60519), .Z(n411) );
  AND U544 ( .A(n60521), .B(n411), .Z(n412) );
  NOR U545 ( .A(n60522), .B(n412), .Z(n413) );
  NAND U546 ( .A(n60523), .B(n413), .Z(n414) );
  NANDN U547 ( .A(n60524), .B(n414), .Z(n415) );
  AND U548 ( .A(n60526), .B(n60525), .Z(n416) );
  NAND U549 ( .A(n415), .B(n416), .Z(n417) );
  NAND U550 ( .A(n60527), .B(n417), .Z(n418) );
  ANDN U551 ( .B(n60529), .A(n60528), .Z(n419) );
  NAND U552 ( .A(n418), .B(n419), .Z(n420) );
  NANDN U553 ( .A(n60530), .B(n420), .Z(n421) );
  ANDN U554 ( .B(n50676), .A(n50677), .Z(n422) );
  NAND U555 ( .A(n421), .B(n422), .Z(n423) );
  NAND U556 ( .A(n60531), .B(n423), .Z(n424) );
  ANDN U557 ( .B(n60533), .A(n60532), .Z(n425) );
  NAND U558 ( .A(n424), .B(n425), .Z(n426) );
  NAND U559 ( .A(n60534), .B(n426), .Z(n60535) );
  AND U560 ( .A(n60992), .B(n60991), .Z(n60993) );
  AND U561 ( .A(n61036), .B(n61037), .Z(n427) );
  NAND U562 ( .A(n61039), .B(n427), .Z(n428) );
  NAND U563 ( .A(n61040), .B(n428), .Z(n429) );
  ANDN U564 ( .B(n50517), .A(n50516), .Z(n430) );
  NAND U565 ( .A(n429), .B(n430), .Z(n431) );
  NANDN U566 ( .A(n61041), .B(n431), .Z(n432) );
  AND U567 ( .A(n61043), .B(n61042), .Z(n433) );
  NAND U568 ( .A(n432), .B(n433), .Z(n434) );
  NAND U569 ( .A(n61044), .B(n434), .Z(n435) );
  AND U570 ( .A(n61046), .B(n61045), .Z(n436) );
  NAND U571 ( .A(n435), .B(n436), .Z(n437) );
  NANDN U572 ( .A(n61047), .B(n437), .Z(n438) );
  AND U573 ( .A(n61049), .B(n61048), .Z(n439) );
  NAND U574 ( .A(n438), .B(n439), .Z(n440) );
  NAND U575 ( .A(n61050), .B(n440), .Z(n441) );
  AND U576 ( .A(n61052), .B(n61051), .Z(n442) );
  NAND U577 ( .A(n441), .B(n442), .Z(n443) );
  NANDN U578 ( .A(n61053), .B(n443), .Z(n61054) );
  NOR U579 ( .A(n50456), .B(n50457), .Z(n444) );
  NANDN U580 ( .A(n61250), .B(n61249), .Z(n445) );
  AND U581 ( .A(n444), .B(n445), .Z(n446) );
  ANDN U582 ( .B(n50453), .A(n50454), .Z(n447) );
  OR U583 ( .A(n61251), .B(n446), .Z(n448) );
  AND U584 ( .A(n447), .B(n448), .Z(n449) );
  ANDN U585 ( .B(n50452), .A(n50451), .Z(n450) );
  NANDN U586 ( .A(n449), .B(n61252), .Z(n451) );
  AND U587 ( .A(n450), .B(n451), .Z(n452) );
  ANDN U588 ( .B(n61255), .A(n61254), .Z(n453) );
  NANDN U589 ( .A(n452), .B(n61253), .Z(n454) );
  AND U590 ( .A(n453), .B(n454), .Z(n455) );
  AND U591 ( .A(n50450), .B(n50449), .Z(n456) );
  NANDN U592 ( .A(n455), .B(n61256), .Z(n457) );
  AND U593 ( .A(n456), .B(n457), .Z(n458) );
  AND U594 ( .A(n61258), .B(n61259), .Z(n459) );
  OR U595 ( .A(n458), .B(n61257), .Z(n460) );
  NAND U596 ( .A(n459), .B(n460), .Z(n61260) );
  NANDN U597 ( .A(n52438), .B(n52439), .Z(n461) );
  NAND U598 ( .A(n52440), .B(n461), .Z(n462) );
  ANDN U599 ( .B(n462), .A(n52441), .Z(n52443) );
  NAND U600 ( .A(n52475), .B(n52474), .Z(n463) );
  NANDN U601 ( .A(n52432), .B(n463), .Z(n464) );
  AND U602 ( .A(n52476), .B(n464), .Z(n465) );
  OR U603 ( .A(n52477), .B(n465), .Z(n466) );
  NAND U604 ( .A(n52478), .B(n466), .Z(n467) );
  NAND U605 ( .A(n52479), .B(n467), .Z(n468) );
  NAND U606 ( .A(n52480), .B(n468), .Z(n469) );
  NAND U607 ( .A(n52481), .B(n469), .Z(n470) );
  ANDN U608 ( .B(n470), .A(n52482), .Z(n471) );
  NANDN U609 ( .A(n471), .B(n52483), .Z(n472) );
  NANDN U610 ( .A(n52484), .B(n472), .Z(n473) );
  NAND U611 ( .A(n52485), .B(n473), .Z(n474) );
  NANDN U612 ( .A(n52486), .B(n474), .Z(n475) );
  NAND U613 ( .A(n52487), .B(n475), .Z(n476) );
  AND U614 ( .A(n52488), .B(n476), .Z(n477) );
  OR U615 ( .A(n52489), .B(n477), .Z(n478) );
  NAND U616 ( .A(n52490), .B(n478), .Z(n479) );
  NANDN U617 ( .A(n52431), .B(n479), .Z(n52491) );
  ANDN U618 ( .B(n28290), .A(n28289), .Z(n52523) );
  NAND U619 ( .A(n52584), .B(n52583), .Z(n480) );
  NANDN U620 ( .A(n52585), .B(n480), .Z(n481) );
  AND U621 ( .A(n52586), .B(n481), .Z(n482) );
  NANDN U622 ( .A(n482), .B(n52587), .Z(n483) );
  NANDN U623 ( .A(n52588), .B(n483), .Z(n484) );
  NAND U624 ( .A(n52589), .B(n484), .Z(n485) );
  NANDN U625 ( .A(n52590), .B(n485), .Z(n486) );
  NAND U626 ( .A(n52426), .B(n486), .Z(n487) );
  ANDN U627 ( .B(n487), .A(n52425), .Z(n488) );
  NANDN U628 ( .A(n488), .B(n52424), .Z(n489) );
  AND U629 ( .A(n52591), .B(n489), .Z(n490) );
  NANDN U630 ( .A(n490), .B(n52592), .Z(n491) );
  NANDN U631 ( .A(n52423), .B(n491), .Z(n492) );
  NAND U632 ( .A(n52422), .B(n492), .Z(n52593) );
  ANDN U633 ( .B(n28268), .A(n28267), .Z(n52605) );
  NAND U634 ( .A(n52727), .B(n52728), .Z(n493) );
  NANDN U635 ( .A(n52729), .B(n493), .Z(n494) );
  NAND U636 ( .A(n52730), .B(n494), .Z(n495) );
  NANDN U637 ( .A(n52731), .B(n495), .Z(n496) );
  NAND U638 ( .A(n52732), .B(n496), .Z(n497) );
  ANDN U639 ( .B(n497), .A(n52733), .Z(n498) );
  OR U640 ( .A(n52734), .B(n498), .Z(n499) );
  NAND U641 ( .A(n52735), .B(n499), .Z(n500) );
  NANDN U642 ( .A(n52736), .B(n500), .Z(n501) );
  NAND U643 ( .A(n52737), .B(n501), .Z(n502) );
  NANDN U644 ( .A(n52738), .B(n502), .Z(n503) );
  ANDN U645 ( .B(n503), .A(n52409), .Z(n504) );
  NANDN U646 ( .A(n504), .B(n52739), .Z(n505) );
  ANDN U647 ( .B(n505), .A(n52408), .Z(n506) );
  NANDN U648 ( .A(n506), .B(n52740), .Z(n507) );
  NANDN U649 ( .A(n52741), .B(n507), .Z(n508) );
  NAND U650 ( .A(n52742), .B(n508), .Z(n52743) );
  NAND U651 ( .A(n52863), .B(n52862), .Z(n509) );
  NANDN U652 ( .A(n52864), .B(n509), .Z(n510) );
  NAND U653 ( .A(n52865), .B(n510), .Z(n511) );
  NANDN U654 ( .A(n52395), .B(n511), .Z(n512) );
  NAND U655 ( .A(n52394), .B(n512), .Z(n513) );
  ANDN U656 ( .B(n513), .A(n52393), .Z(n514) );
  NANDN U657 ( .A(n514), .B(n52392), .Z(n515) );
  ANDN U658 ( .B(n515), .A(n52866), .Z(n516) );
  NANDN U659 ( .A(n516), .B(n52867), .Z(n517) );
  NANDN U660 ( .A(n52391), .B(n517), .Z(n518) );
  NAND U661 ( .A(n52390), .B(n518), .Z(n52868) );
  NAND U662 ( .A(n52377), .B(n52885), .Z(n519) );
  NANDN U663 ( .A(n52886), .B(n519), .Z(n520) );
  AND U664 ( .A(n52887), .B(n520), .Z(n521) );
  OR U665 ( .A(n52376), .B(n521), .Z(n522) );
  NAND U666 ( .A(n52888), .B(n522), .Z(n523) );
  NANDN U667 ( .A(n52375), .B(n523), .Z(n524) );
  NAND U668 ( .A(n52374), .B(n524), .Z(n525) );
  NAND U669 ( .A(n52889), .B(n525), .Z(n526) );
  AND U670 ( .A(n52890), .B(n526), .Z(n527) );
  NANDN U671 ( .A(n527), .B(n52891), .Z(n528) );
  NAND U672 ( .A(n52373), .B(n528), .Z(n529) );
  NANDN U673 ( .A(n52372), .B(n529), .Z(n52892) );
  NAND U674 ( .A(n52915), .B(n52916), .Z(n530) );
  NANDN U675 ( .A(n52917), .B(n530), .Z(n531) );
  NAND U676 ( .A(n52918), .B(n531), .Z(n532) );
  NANDN U677 ( .A(n52362), .B(n532), .Z(n533) );
  NAND U678 ( .A(n52919), .B(n533), .Z(n534) );
  ANDN U679 ( .B(n534), .A(n52361), .Z(n535) );
  NANDN U680 ( .A(n535), .B(n52920), .Z(n536) );
  NANDN U681 ( .A(n52921), .B(n536), .Z(n537) );
  NAND U682 ( .A(n52922), .B(n537), .Z(n538) );
  NAND U683 ( .A(n52923), .B(n538), .Z(n539) );
  NANDN U684 ( .A(n52924), .B(n539), .Z(n540) );
  AND U685 ( .A(n52925), .B(n540), .Z(n541) );
  NANDN U686 ( .A(n541), .B(n52926), .Z(n542) );
  NAND U687 ( .A(n52927), .B(n542), .Z(n543) );
  NANDN U688 ( .A(n52928), .B(n543), .Z(n52929) );
  NAND U689 ( .A(n52961), .B(n52962), .Z(n544) );
  NANDN U690 ( .A(n52963), .B(n544), .Z(n545) );
  AND U691 ( .A(n52964), .B(n545), .Z(n546) );
  OR U692 ( .A(n546), .B(n52965), .Z(n547) );
  NAND U693 ( .A(n52966), .B(n547), .Z(n548) );
  NANDN U694 ( .A(n52967), .B(n548), .Z(n549) );
  NAND U695 ( .A(n52355), .B(n549), .Z(n550) );
  NAND U696 ( .A(n52968), .B(n550), .Z(n551) );
  AND U697 ( .A(n52969), .B(n551), .Z(n552) );
  OR U698 ( .A(n52970), .B(n552), .Z(n553) );
  NAND U699 ( .A(n52971), .B(n553), .Z(n554) );
  NANDN U700 ( .A(n52972), .B(n554), .Z(n555) );
  NAND U701 ( .A(n52973), .B(n555), .Z(n556) );
  NANDN U702 ( .A(n52974), .B(n556), .Z(n557) );
  AND U703 ( .A(n52975), .B(n557), .Z(n558) );
  OR U704 ( .A(n558), .B(n52976), .Z(n559) );
  NAND U705 ( .A(n52977), .B(n559), .Z(n560) );
  NAND U706 ( .A(n52978), .B(n560), .Z(n52979) );
  NAND U707 ( .A(n53016), .B(n53015), .Z(n561) );
  NANDN U708 ( .A(n53017), .B(n561), .Z(n562) );
  AND U709 ( .A(n53018), .B(n562), .Z(n563) );
  OR U710 ( .A(n53019), .B(n563), .Z(n564) );
  NAND U711 ( .A(n53020), .B(n564), .Z(n565) );
  NANDN U712 ( .A(n53021), .B(n565), .Z(n566) );
  NAND U713 ( .A(n53022), .B(n566), .Z(n567) );
  NAND U714 ( .A(n53023), .B(n567), .Z(n568) );
  AND U715 ( .A(n53024), .B(n568), .Z(n569) );
  OR U716 ( .A(n53025), .B(n569), .Z(n570) );
  NAND U717 ( .A(n53026), .B(n570), .Z(n571) );
  NANDN U718 ( .A(n53027), .B(n571), .Z(n572) );
  NAND U719 ( .A(n53028), .B(n572), .Z(n573) );
  NAND U720 ( .A(n53029), .B(n573), .Z(n574) );
  ANDN U721 ( .B(n574), .A(n52352), .Z(n575) );
  NANDN U722 ( .A(n575), .B(n53030), .Z(n576) );
  NAND U723 ( .A(n53031), .B(n576), .Z(n577) );
  NANDN U724 ( .A(n53032), .B(n577), .Z(n578) );
  NAND U725 ( .A(n53033), .B(n578), .Z(n53034) );
  NAND U726 ( .A(n53071), .B(n53070), .Z(n579) );
  NAND U727 ( .A(n53073), .B(n579), .Z(n580) );
  AND U728 ( .A(n53074), .B(n580), .Z(n581) );
  OR U729 ( .A(n52349), .B(n581), .Z(n582) );
  NAND U730 ( .A(n53075), .B(n582), .Z(n583) );
  NANDN U731 ( .A(n52348), .B(n583), .Z(n584) );
  NAND U732 ( .A(n53076), .B(n584), .Z(n585) );
  NANDN U733 ( .A(n53077), .B(n585), .Z(n586) );
  AND U734 ( .A(n53078), .B(n586), .Z(n587) );
  OR U735 ( .A(n52347), .B(n587), .Z(n588) );
  NAND U736 ( .A(n53079), .B(n588), .Z(n589) );
  NANDN U737 ( .A(n53080), .B(n589), .Z(n590) );
  NAND U738 ( .A(n53081), .B(n590), .Z(n591) );
  NANDN U739 ( .A(n53082), .B(n591), .Z(n592) );
  AND U740 ( .A(n53083), .B(n592), .Z(n53085) );
  ANDN U741 ( .B(n28064), .A(n28063), .Z(n53152) );
  NOR U742 ( .A(n28060), .B(n28061), .Z(n53165) );
  NAND U743 ( .A(n53180), .B(n53179), .Z(n593) );
  NAND U744 ( .A(n53181), .B(n593), .Z(n594) );
  ANDN U745 ( .B(n594), .A(n52333), .Z(n595) );
  NANDN U746 ( .A(n595), .B(n52332), .Z(n596) );
  NANDN U747 ( .A(n52331), .B(n596), .Z(n597) );
  NAND U748 ( .A(n52330), .B(n597), .Z(n598) );
  NANDN U749 ( .A(n53182), .B(n598), .Z(n599) );
  NAND U750 ( .A(n53183), .B(n599), .Z(n600) );
  ANDN U751 ( .B(n600), .A(n53184), .Z(n601) );
  NANDN U752 ( .A(n601), .B(n53185), .Z(n602) );
  NANDN U753 ( .A(n53186), .B(n602), .Z(n603) );
  NAND U754 ( .A(n53187), .B(n603), .Z(n604) );
  NANDN U755 ( .A(n53188), .B(n604), .Z(n53189) );
  NAND U756 ( .A(n53227), .B(n53226), .Z(n605) );
  NANDN U757 ( .A(n52326), .B(n605), .Z(n606) );
  NAND U758 ( .A(n53228), .B(n606), .Z(n607) );
  NAND U759 ( .A(n53229), .B(n607), .Z(n608) );
  NANDN U760 ( .A(n53230), .B(n608), .Z(n609) );
  ANDN U761 ( .B(n609), .A(n53231), .Z(n610) );
  NANDN U762 ( .A(n610), .B(n53232), .Z(n611) );
  NANDN U763 ( .A(n53233), .B(n611), .Z(n612) );
  NAND U764 ( .A(n53234), .B(n612), .Z(n613) );
  NAND U765 ( .A(n53235), .B(n613), .Z(n614) );
  NAND U766 ( .A(n52325), .B(n614), .Z(n615) );
  AND U767 ( .A(n53236), .B(n615), .Z(n616) );
  NANDN U768 ( .A(n616), .B(n52324), .Z(n617) );
  NANDN U769 ( .A(n53237), .B(n617), .Z(n618) );
  NAND U770 ( .A(n53238), .B(n618), .Z(n53239) );
  NANDN U771 ( .A(n53270), .B(n53271), .Z(n619) );
  NANDN U772 ( .A(n53273), .B(n619), .Z(n620) );
  ANDN U773 ( .B(n620), .A(n52317), .Z(n621) );
  NANDN U774 ( .A(n621), .B(n52316), .Z(n622) );
  NANDN U775 ( .A(n53274), .B(n622), .Z(n623) );
  NANDN U776 ( .A(n53275), .B(n623), .Z(n624) );
  NAND U777 ( .A(n53276), .B(n624), .Z(n625) );
  NANDN U778 ( .A(n53277), .B(n625), .Z(n626) );
  AND U779 ( .A(n53278), .B(n626), .Z(n627) );
  OR U780 ( .A(n53279), .B(n627), .Z(n628) );
  AND U781 ( .A(n53280), .B(n628), .Z(n629) );
  OR U782 ( .A(n52315), .B(n629), .Z(n630) );
  NAND U783 ( .A(n53281), .B(n630), .Z(n631) );
  NANDN U784 ( .A(n52314), .B(n631), .Z(n53282) );
  OR U785 ( .A(n53318), .B(n53319), .Z(n632) );
  NAND U786 ( .A(n53320), .B(n632), .Z(n633) );
  NANDN U787 ( .A(n53321), .B(n633), .Z(n634) );
  NAND U788 ( .A(n52311), .B(n634), .Z(n635) );
  NANDN U789 ( .A(n53322), .B(n635), .Z(n636) );
  AND U790 ( .A(n53323), .B(n636), .Z(n637) );
  NANDN U791 ( .A(n637), .B(n53324), .Z(n638) );
  NANDN U792 ( .A(n53325), .B(n638), .Z(n639) );
  NAND U793 ( .A(n53326), .B(n639), .Z(n640) );
  NANDN U794 ( .A(n53327), .B(n640), .Z(n641) );
  NAND U795 ( .A(n53328), .B(n641), .Z(n642) );
  ANDN U796 ( .B(n642), .A(n53329), .Z(n643) );
  NANDN U797 ( .A(n643), .B(n53330), .Z(n644) );
  ANDN U798 ( .B(n644), .A(n53331), .Z(n645) );
  NANDN U799 ( .A(n645), .B(n53332), .Z(n646) );
  NANDN U800 ( .A(n53333), .B(n646), .Z(n647) );
  NAND U801 ( .A(n53334), .B(n647), .Z(n53335) );
  ANDN U802 ( .B(n27943), .A(n27942), .Z(n53357) );
  NAND U803 ( .A(n53431), .B(n53432), .Z(n648) );
  NAND U804 ( .A(n53433), .B(n648), .Z(n649) );
  NANDN U805 ( .A(n52296), .B(n649), .Z(n650) );
  NAND U806 ( .A(n52295), .B(n650), .Z(n651) );
  NANDN U807 ( .A(n52294), .B(n651), .Z(n652) );
  AND U808 ( .A(n52293), .B(n652), .Z(n653) );
  OR U809 ( .A(n53434), .B(n653), .Z(n654) );
  AND U810 ( .A(n53435), .B(n654), .Z(n655) );
  OR U811 ( .A(n52292), .B(n655), .Z(n656) );
  NAND U812 ( .A(n52291), .B(n656), .Z(n657) );
  NANDN U813 ( .A(n52290), .B(n657), .Z(n53436) );
  NAND U814 ( .A(n53464), .B(n53463), .Z(n658) );
  NAND U815 ( .A(n53465), .B(n658), .Z(n659) );
  NANDN U816 ( .A(n53466), .B(n659), .Z(n660) );
  NAND U817 ( .A(n53467), .B(n660), .Z(n661) );
  NANDN U818 ( .A(n53468), .B(n661), .Z(n662) );
  AND U819 ( .A(n53469), .B(n662), .Z(n663) );
  OR U820 ( .A(n53470), .B(n663), .Z(n664) );
  NANDN U821 ( .A(n53471), .B(n664), .Z(n665) );
  NAND U822 ( .A(n53472), .B(n665), .Z(n666) );
  NANDN U823 ( .A(n53473), .B(n666), .Z(n667) );
  NAND U824 ( .A(n53474), .B(n667), .Z(n668) );
  ANDN U825 ( .B(n668), .A(n52282), .Z(n669) );
  NANDN U826 ( .A(n669), .B(n53475), .Z(n670) );
  AND U827 ( .A(n53476), .B(n670), .Z(n671) );
  NANDN U828 ( .A(n671), .B(n53477), .Z(n672) );
  NAND U829 ( .A(n53478), .B(n672), .Z(n673) );
  NANDN U830 ( .A(n53479), .B(n673), .Z(n53482) );
  NAND U831 ( .A(n53509), .B(n52276), .Z(n674) );
  NANDN U832 ( .A(n53510), .B(n674), .Z(n675) );
  NAND U833 ( .A(n53511), .B(n675), .Z(n676) );
  NANDN U834 ( .A(n53512), .B(n676), .Z(n677) );
  NANDN U835 ( .A(n53513), .B(n677), .Z(n678) );
  AND U836 ( .A(n53514), .B(n678), .Z(n679) );
  OR U837 ( .A(n52275), .B(n679), .Z(n680) );
  NAND U838 ( .A(n53515), .B(n680), .Z(n681) );
  NANDN U839 ( .A(n53516), .B(n681), .Z(n682) );
  NANDN U840 ( .A(n52274), .B(n682), .Z(n683) );
  NANDN U841 ( .A(n53517), .B(n683), .Z(n684) );
  ANDN U842 ( .B(n684), .A(n53518), .Z(n685) );
  NANDN U843 ( .A(n685), .B(n53519), .Z(n686) );
  NANDN U844 ( .A(n52273), .B(n686), .Z(n687) );
  NAND U845 ( .A(n53520), .B(n687), .Z(n53521) );
  NAND U846 ( .A(n53548), .B(n53549), .Z(n688) );
  NAND U847 ( .A(n53550), .B(n688), .Z(n689) );
  ANDN U848 ( .B(n689), .A(n53551), .Z(n690) );
  NANDN U849 ( .A(n690), .B(n53552), .Z(n691) );
  NAND U850 ( .A(n53553), .B(n691), .Z(n692) );
  NAND U851 ( .A(n52266), .B(n692), .Z(n693) );
  NANDN U852 ( .A(n52265), .B(n693), .Z(n694) );
  NAND U853 ( .A(n53554), .B(n694), .Z(n695) );
  ANDN U854 ( .B(n695), .A(n53555), .Z(n696) );
  NANDN U855 ( .A(n696), .B(n53556), .Z(n697) );
  NANDN U856 ( .A(n52264), .B(n697), .Z(n698) );
  NAND U857 ( .A(n53557), .B(n698), .Z(n699) );
  NAND U858 ( .A(n53558), .B(n699), .Z(n700) );
  NANDN U859 ( .A(n53559), .B(n700), .Z(n701) );
  AND U860 ( .A(n53560), .B(n701), .Z(n53561) );
  NANDN U861 ( .A(n53592), .B(n53591), .Z(n702) );
  NAND U862 ( .A(n53593), .B(n702), .Z(n703) );
  NANDN U863 ( .A(n53594), .B(n703), .Z(n704) );
  NAND U864 ( .A(n53595), .B(n704), .Z(n705) );
  NANDN U865 ( .A(n52258), .B(n705), .Z(n706) );
  AND U866 ( .A(n52257), .B(n706), .Z(n707) );
  OR U867 ( .A(n53596), .B(n707), .Z(n708) );
  NAND U868 ( .A(n53597), .B(n708), .Z(n709) );
  NANDN U869 ( .A(n53598), .B(n709), .Z(n710) );
  NANDN U870 ( .A(n53599), .B(n710), .Z(n711) );
  NANDN U871 ( .A(n53600), .B(n711), .Z(n712) );
  AND U872 ( .A(n53601), .B(n712), .Z(n713) );
  OR U873 ( .A(n53602), .B(n713), .Z(n714) );
  NAND U874 ( .A(n53603), .B(n714), .Z(n715) );
  NANDN U875 ( .A(n53604), .B(n715), .Z(n716) );
  NAND U876 ( .A(n53605), .B(n716), .Z(n53606) );
  ANDN U877 ( .B(n27737), .A(n27736), .Z(n53629) );
  NANDN U878 ( .A(n53710), .B(n53709), .Z(n717) );
  NAND U879 ( .A(n53711), .B(n717), .Z(n718) );
  ANDN U880 ( .B(n718), .A(n53712), .Z(n719) );
  NANDN U881 ( .A(n719), .B(n53713), .Z(n720) );
  NANDN U882 ( .A(n53714), .B(n720), .Z(n721) );
  NANDN U883 ( .A(n53715), .B(n721), .Z(n722) );
  NAND U884 ( .A(n53716), .B(n722), .Z(n723) );
  NANDN U885 ( .A(n53717), .B(n723), .Z(n724) );
  AND U886 ( .A(n53718), .B(n724), .Z(n725) );
  OR U887 ( .A(n53719), .B(n725), .Z(n726) );
  NAND U888 ( .A(n53720), .B(n726), .Z(n727) );
  NANDN U889 ( .A(n53721), .B(n727), .Z(n728) );
  NAND U890 ( .A(n53722), .B(n728), .Z(n729) );
  NANDN U891 ( .A(n53723), .B(n729), .Z(n730) );
  AND U892 ( .A(n53724), .B(n730), .Z(n731) );
  OR U893 ( .A(n53725), .B(n731), .Z(n732) );
  NAND U894 ( .A(n53726), .B(n732), .Z(n733) );
  NANDN U895 ( .A(n53727), .B(n733), .Z(n734) );
  NAND U896 ( .A(n53728), .B(n734), .Z(n53729) );
  NOR U897 ( .A(n33647), .B(n33648), .Z(n53743) );
  NAND U898 ( .A(n53789), .B(n53790), .Z(n735) );
  NANDN U899 ( .A(n53791), .B(n735), .Z(n736) );
  AND U900 ( .A(n53792), .B(n736), .Z(n737) );
  OR U901 ( .A(n53793), .B(n737), .Z(n738) );
  NAND U902 ( .A(n53794), .B(n738), .Z(n739) );
  NANDN U903 ( .A(n53795), .B(n739), .Z(n740) );
  NAND U904 ( .A(n53796), .B(n740), .Z(n741) );
  NAND U905 ( .A(n53797), .B(n741), .Z(n742) );
  ANDN U906 ( .B(n742), .A(n53798), .Z(n743) );
  NANDN U907 ( .A(n743), .B(n53799), .Z(n744) );
  NANDN U908 ( .A(n52235), .B(n744), .Z(n745) );
  NAND U909 ( .A(n53800), .B(n745), .Z(n746) );
  NANDN U910 ( .A(n53801), .B(n746), .Z(n747) );
  NANDN U911 ( .A(n53802), .B(n747), .Z(n748) );
  AND U912 ( .A(n53803), .B(n748), .Z(n749) );
  OR U913 ( .A(n53804), .B(n749), .Z(n750) );
  NAND U914 ( .A(n53805), .B(n750), .Z(n751) );
  NANDN U915 ( .A(n53806), .B(n751), .Z(n53807) );
  OR U916 ( .A(n53830), .B(n53831), .Z(n752) );
  NANDN U917 ( .A(n52224), .B(n752), .Z(n753) );
  NAND U918 ( .A(n53832), .B(n753), .Z(n754) );
  NANDN U919 ( .A(n52223), .B(n754), .Z(n755) );
  NAND U920 ( .A(n53833), .B(n755), .Z(n756) );
  ANDN U921 ( .B(n756), .A(n53834), .Z(n757) );
  OR U922 ( .A(n52222), .B(n757), .Z(n758) );
  NAND U923 ( .A(n53835), .B(n758), .Z(n759) );
  NAND U924 ( .A(n53836), .B(n759), .Z(n760) );
  NANDN U925 ( .A(n53837), .B(n760), .Z(n761) );
  NAND U926 ( .A(n53838), .B(n761), .Z(n762) );
  AND U927 ( .A(n52221), .B(n762), .Z(n763) );
  NANDN U928 ( .A(n763), .B(n52220), .Z(n764) );
  NAND U929 ( .A(n53839), .B(n764), .Z(n765) );
  NANDN U930 ( .A(n53840), .B(n765), .Z(n53841) );
  NANDN U931 ( .A(n53867), .B(n53866), .Z(n766) );
  NAND U932 ( .A(n53868), .B(n766), .Z(n767) );
  ANDN U933 ( .B(n767), .A(n53869), .Z(n768) );
  NOR U934 ( .A(n53871), .B(n768), .Z(n769) );
  NAND U935 ( .A(n53870), .B(n769), .Z(n770) );
  AND U936 ( .A(n53872), .B(n770), .Z(n771) );
  NANDN U937 ( .A(n771), .B(n53873), .Z(n772) );
  NAND U938 ( .A(n53874), .B(n772), .Z(n773) );
  NAND U939 ( .A(n52213), .B(n773), .Z(n774) );
  NAND U940 ( .A(n53875), .B(n774), .Z(n775) );
  NAND U941 ( .A(n53876), .B(n775), .Z(n776) );
  ANDN U942 ( .B(n776), .A(n53877), .Z(n777) );
  NANDN U943 ( .A(n777), .B(n53878), .Z(n778) );
  NANDN U944 ( .A(n53879), .B(n778), .Z(n779) );
  NAND U945 ( .A(n53880), .B(n779), .Z(n780) );
  NANDN U946 ( .A(n53881), .B(n780), .Z(n53882) );
  OR U947 ( .A(n53914), .B(n53915), .Z(n781) );
  NAND U948 ( .A(n53917), .B(n781), .Z(n782) );
  AND U949 ( .A(n53918), .B(n782), .Z(n783) );
  OR U950 ( .A(n52207), .B(n783), .Z(n784) );
  NAND U951 ( .A(n52206), .B(n784), .Z(n785) );
  NAND U952 ( .A(n53919), .B(n785), .Z(n786) );
  NANDN U953 ( .A(n52205), .B(n786), .Z(n787) );
  NAND U954 ( .A(n52204), .B(n787), .Z(n788) );
  ANDN U955 ( .B(n788), .A(n53920), .Z(n789) );
  NANDN U956 ( .A(n789), .B(n53921), .Z(n790) );
  AND U957 ( .A(n53922), .B(n790), .Z(n791) );
  NANDN U958 ( .A(n791), .B(n53923), .Z(n792) );
  NAND U959 ( .A(n53924), .B(n792), .Z(n793) );
  NAND U960 ( .A(n53925), .B(n793), .Z(n53926) );
  NANDN U961 ( .A(n53957), .B(n53956), .Z(n794) );
  NAND U962 ( .A(n53958), .B(n794), .Z(n795) );
  ANDN U963 ( .B(n795), .A(n53959), .Z(n796) );
  NANDN U964 ( .A(n796), .B(n53960), .Z(n797) );
  NANDN U965 ( .A(n53961), .B(n797), .Z(n798) );
  NAND U966 ( .A(n53962), .B(n798), .Z(n799) );
  NANDN U967 ( .A(n53963), .B(n799), .Z(n800) );
  NAND U968 ( .A(n53964), .B(n800), .Z(n801) );
  AND U969 ( .A(n53965), .B(n801), .Z(n802) );
  NANDN U970 ( .A(n802), .B(n53966), .Z(n803) );
  NAND U971 ( .A(n53967), .B(n803), .Z(n804) );
  NANDN U972 ( .A(n53968), .B(n804), .Z(n805) );
  NAND U973 ( .A(n53969), .B(n805), .Z(n806) );
  NAND U974 ( .A(n53970), .B(n806), .Z(n807) );
  ANDN U975 ( .B(n807), .A(n53971), .Z(n808) );
  NANDN U976 ( .A(n808), .B(n53972), .Z(n809) );
  NAND U977 ( .A(n53973), .B(n809), .Z(n810) );
  NANDN U978 ( .A(n53974), .B(n810), .Z(n53975) );
  NANDN U979 ( .A(n54009), .B(n54008), .Z(n811) );
  NAND U980 ( .A(n54010), .B(n811), .Z(n812) );
  NANDN U981 ( .A(n54011), .B(n812), .Z(n813) );
  NANDN U982 ( .A(n52195), .B(n813), .Z(n814) );
  NAND U983 ( .A(n52194), .B(n814), .Z(n815) );
  ANDN U984 ( .B(n815), .A(n52193), .Z(n816) );
  NANDN U985 ( .A(n816), .B(n54012), .Z(n817) );
  NANDN U986 ( .A(n54013), .B(n817), .Z(n818) );
  NANDN U987 ( .A(n52192), .B(n818), .Z(n819) );
  NAND U988 ( .A(n54014), .B(n819), .Z(n820) );
  NAND U989 ( .A(n54015), .B(n820), .Z(n821) );
  AND U990 ( .A(n54016), .B(n821), .Z(n822) );
  NANDN U991 ( .A(n822), .B(n54017), .Z(n823) );
  NANDN U992 ( .A(n54018), .B(n823), .Z(n824) );
  NAND U993 ( .A(n54019), .B(n824), .Z(n825) );
  NANDN U994 ( .A(n54020), .B(n825), .Z(n54021) );
  NANDN U995 ( .A(n54043), .B(n54044), .Z(n826) );
  NANDN U996 ( .A(n54045), .B(n826), .Z(n827) );
  NAND U997 ( .A(n54046), .B(n827), .Z(n828) );
  NANDN U998 ( .A(n54047), .B(n828), .Z(n829) );
  NANDN U999 ( .A(n52184), .B(n829), .Z(n830) );
  AND U1000 ( .A(n54048), .B(n830), .Z(n831) );
  OR U1001 ( .A(n54049), .B(n831), .Z(n832) );
  AND U1002 ( .A(n54050), .B(n832), .Z(n833) );
  OR U1003 ( .A(n54051), .B(n833), .Z(n834) );
  NANDN U1004 ( .A(n54052), .B(n834), .Z(n835) );
  NAND U1005 ( .A(n54053), .B(n835), .Z(n836) );
  ANDN U1006 ( .B(n54054), .A(n54055), .Z(n837) );
  NAND U1007 ( .A(n836), .B(n837), .Z(n838) );
  NAND U1008 ( .A(n54056), .B(n838), .Z(n839) );
  ANDN U1009 ( .B(n52183), .A(n52182), .Z(n840) );
  NAND U1010 ( .A(n839), .B(n840), .Z(n841) );
  NAND U1011 ( .A(n54057), .B(n841), .Z(n54058) );
  NAND U1012 ( .A(n54085), .B(n54084), .Z(n842) );
  NANDN U1013 ( .A(n54086), .B(n842), .Z(n843) );
  NAND U1014 ( .A(n52175), .B(n843), .Z(n844) );
  NANDN U1015 ( .A(n54087), .B(n844), .Z(n845) );
  NAND U1016 ( .A(n54088), .B(n845), .Z(n846) );
  ANDN U1017 ( .B(n846), .A(n52174), .Z(n847) );
  OR U1018 ( .A(n847), .B(n54089), .Z(n848) );
  NAND U1019 ( .A(n54090), .B(n848), .Z(n849) );
  ANDN U1020 ( .B(n849), .A(n54091), .Z(n850) );
  NANDN U1021 ( .A(n850), .B(n54092), .Z(n851) );
  NANDN U1022 ( .A(n52173), .B(n851), .Z(n852) );
  NANDN U1023 ( .A(n54093), .B(n852), .Z(n853) );
  NAND U1024 ( .A(n52172), .B(n853), .Z(n54096) );
  OR U1025 ( .A(n54115), .B(n54116), .Z(n854) );
  NANDN U1026 ( .A(n54117), .B(n854), .Z(n855) );
  NAND U1027 ( .A(n54118), .B(n855), .Z(n856) );
  NAND U1028 ( .A(n54119), .B(n856), .Z(n857) );
  NAND U1029 ( .A(n54120), .B(n857), .Z(n858) );
  AND U1030 ( .A(n54121), .B(n858), .Z(n859) );
  OR U1031 ( .A(n52161), .B(n859), .Z(n860) );
  NAND U1032 ( .A(n54122), .B(n860), .Z(n861) );
  NANDN U1033 ( .A(n54123), .B(n861), .Z(n862) );
  NAND U1034 ( .A(n54124), .B(n862), .Z(n863) );
  NANDN U1035 ( .A(n54125), .B(n863), .Z(n864) );
  ANDN U1036 ( .B(n864), .A(n52160), .Z(n865) );
  NANDN U1037 ( .A(n865), .B(n52159), .Z(n866) );
  NANDN U1038 ( .A(n54126), .B(n866), .Z(n867) );
  NAND U1039 ( .A(n54127), .B(n867), .Z(n868) );
  NANDN U1040 ( .A(n54128), .B(n868), .Z(n54129) );
  NANDN U1041 ( .A(n54163), .B(n54162), .Z(n869) );
  AND U1042 ( .A(n54164), .B(n869), .Z(n870) );
  OR U1043 ( .A(n54165), .B(n54166), .Z(n871) );
  NAND U1044 ( .A(n870), .B(n871), .Z(n872) );
  ANDN U1045 ( .B(n872), .A(n54167), .Z(n873) );
  NANDN U1046 ( .A(n873), .B(n54168), .Z(n874) );
  NANDN U1047 ( .A(n54169), .B(n874), .Z(n875) );
  NAND U1048 ( .A(n52154), .B(n875), .Z(n876) );
  NANDN U1049 ( .A(n54170), .B(n876), .Z(n877) );
  NANDN U1050 ( .A(n54171), .B(n877), .Z(n878) );
  AND U1051 ( .A(n54172), .B(n878), .Z(n879) );
  OR U1052 ( .A(n879), .B(n54173), .Z(n880) );
  AND U1053 ( .A(n52153), .B(n880), .Z(n881) );
  OR U1054 ( .A(n54174), .B(n881), .Z(n882) );
  NAND U1055 ( .A(n54175), .B(n882), .Z(n883) );
  NANDN U1056 ( .A(n54176), .B(n883), .Z(n54177) );
  OR U1057 ( .A(n54249), .B(n54250), .Z(n884) );
  NAND U1058 ( .A(n54251), .B(n884), .Z(n885) );
  ANDN U1059 ( .B(n885), .A(n54252), .Z(n886) );
  NANDN U1060 ( .A(n886), .B(n54253), .Z(n887) );
  NANDN U1061 ( .A(n54254), .B(n887), .Z(n888) );
  NANDN U1062 ( .A(n54255), .B(n888), .Z(n889) );
  NAND U1063 ( .A(n54256), .B(n889), .Z(n890) );
  NANDN U1064 ( .A(n52148), .B(n890), .Z(n891) );
  AND U1065 ( .A(n54257), .B(n891), .Z(n892) );
  OR U1066 ( .A(n892), .B(n54258), .Z(n893) );
  NAND U1067 ( .A(n54259), .B(n893), .Z(n894) );
  ANDN U1068 ( .B(n894), .A(n54260), .Z(n895) );
  NANDN U1069 ( .A(n895), .B(n54261), .Z(n896) );
  ANDN U1070 ( .B(n896), .A(n54262), .Z(n897) );
  NANDN U1071 ( .A(n897), .B(n54263), .Z(n898) );
  NANDN U1072 ( .A(n54264), .B(n898), .Z(n899) );
  NAND U1073 ( .A(n54265), .B(n899), .Z(n54266) );
  NAND U1074 ( .A(n54303), .B(n54304), .Z(n900) );
  NAND U1075 ( .A(n54305), .B(n900), .Z(n901) );
  NANDN U1076 ( .A(n52145), .B(n901), .Z(n902) );
  NAND U1077 ( .A(n52144), .B(n902), .Z(n903) );
  NANDN U1078 ( .A(n54306), .B(n903), .Z(n904) );
  AND U1079 ( .A(n54307), .B(n904), .Z(n905) );
  NANDN U1080 ( .A(n905), .B(n54308), .Z(n906) );
  NAND U1081 ( .A(n54309), .B(n906), .Z(n907) );
  NAND U1082 ( .A(n54310), .B(n907), .Z(n908) );
  NAND U1083 ( .A(n54311), .B(n908), .Z(n909) );
  NAND U1084 ( .A(n54312), .B(n909), .Z(n910) );
  ANDN U1085 ( .B(n910), .A(n54313), .Z(n911) );
  OR U1086 ( .A(n911), .B(n54314), .Z(n912) );
  NAND U1087 ( .A(n54315), .B(n912), .Z(n913) );
  NANDN U1088 ( .A(n54316), .B(n913), .Z(n54317) );
  OR U1089 ( .A(n54350), .B(n54351), .Z(n914) );
  NANDN U1090 ( .A(n52140), .B(n914), .Z(n915) );
  AND U1091 ( .A(n52139), .B(n915), .Z(n916) );
  OR U1092 ( .A(n916), .B(n54352), .Z(n917) );
  NANDN U1093 ( .A(n54353), .B(n917), .Z(n918) );
  NAND U1094 ( .A(n54354), .B(n918), .Z(n919) );
  NANDN U1095 ( .A(n52138), .B(n919), .Z(n920) );
  NAND U1096 ( .A(n52137), .B(n920), .Z(n921) );
  ANDN U1097 ( .B(n921), .A(n52136), .Z(n922) );
  NANDN U1098 ( .A(n922), .B(n52135), .Z(n923) );
  NAND U1099 ( .A(n54355), .B(n923), .Z(n924) );
  NANDN U1100 ( .A(n54356), .B(n924), .Z(n925) );
  AND U1101 ( .A(n54357), .B(n925), .Z(n54359) );
  NANDN U1102 ( .A(n52128), .B(n54385), .Z(n926) );
  NAND U1103 ( .A(n54386), .B(n926), .Z(n927) );
  ANDN U1104 ( .B(n927), .A(n54387), .Z(n928) );
  OR U1105 ( .A(n54388), .B(n928), .Z(n929) );
  NAND U1106 ( .A(n54389), .B(n929), .Z(n930) );
  NANDN U1107 ( .A(n52127), .B(n930), .Z(n931) );
  NAND U1108 ( .A(n54390), .B(n931), .Z(n932) );
  NAND U1109 ( .A(n54391), .B(n932), .Z(n933) );
  ANDN U1110 ( .B(n933), .A(n54392), .Z(n934) );
  NANDN U1111 ( .A(n934), .B(n54393), .Z(n935) );
  NAND U1112 ( .A(n54394), .B(n935), .Z(n936) );
  NANDN U1113 ( .A(n52126), .B(n936), .Z(n937) );
  NAND U1114 ( .A(n52125), .B(n937), .Z(n54395) );
  ANDN U1115 ( .B(n27216), .A(n27215), .Z(n54417) );
  ANDN U1116 ( .B(n27201), .A(n27200), .Z(n54438) );
  NANDN U1117 ( .A(n54493), .B(n54492), .Z(n938) );
  NANDN U1118 ( .A(n54494), .B(n938), .Z(n939) );
  ANDN U1119 ( .B(n939), .A(n54495), .Z(n940) );
  NANDN U1120 ( .A(n940), .B(n54496), .Z(n941) );
  NANDN U1121 ( .A(n52101), .B(n941), .Z(n942) );
  NAND U1122 ( .A(n54497), .B(n942), .Z(n943) );
  NANDN U1123 ( .A(n52100), .B(n943), .Z(n944) );
  NANDN U1124 ( .A(n54498), .B(n944), .Z(n945) );
  ANDN U1125 ( .B(n945), .A(n54499), .Z(n946) );
  NANDN U1126 ( .A(n946), .B(n54500), .Z(n947) );
  NAND U1127 ( .A(n54501), .B(n947), .Z(n948) );
  NAND U1128 ( .A(n52099), .B(n948), .Z(n949) );
  NANDN U1129 ( .A(n54502), .B(n949), .Z(n54503) );
  ANDN U1130 ( .B(n35533), .A(n35532), .Z(n54551) );
  NANDN U1131 ( .A(n54580), .B(n54579), .Z(n950) );
  NAND U1132 ( .A(n54581), .B(n950), .Z(n951) );
  NANDN U1133 ( .A(n54582), .B(n951), .Z(n952) );
  NAND U1134 ( .A(n54583), .B(n952), .Z(n953) );
  NAND U1135 ( .A(n54584), .B(n953), .Z(n954) );
  AND U1136 ( .A(n54585), .B(n954), .Z(n955) );
  OR U1137 ( .A(n54586), .B(n955), .Z(n956) );
  NAND U1138 ( .A(n54587), .B(n956), .Z(n957) );
  NAND U1139 ( .A(n54588), .B(n957), .Z(n958) );
  NANDN U1140 ( .A(n54589), .B(n958), .Z(n959) );
  NAND U1141 ( .A(n54590), .B(n959), .Z(n960) );
  ANDN U1142 ( .B(n960), .A(n54591), .Z(n961) );
  OR U1143 ( .A(n54592), .B(n961), .Z(n962) );
  NAND U1144 ( .A(n54593), .B(n962), .Z(n963) );
  NANDN U1145 ( .A(n52087), .B(n963), .Z(n964) );
  NAND U1146 ( .A(n54594), .B(n964), .Z(n965) );
  AND U1147 ( .A(n54595), .B(n965), .Z(n966) );
  NAND U1148 ( .A(n966), .B(n54596), .Z(n54599) );
  NAND U1149 ( .A(n54629), .B(n54628), .Z(n967) );
  NANDN U1150 ( .A(n54630), .B(n967), .Z(n968) );
  AND U1151 ( .A(n54631), .B(n968), .Z(n969) );
  NANDN U1152 ( .A(n969), .B(n54632), .Z(n970) );
  NAND U1153 ( .A(n54633), .B(n970), .Z(n971) );
  NANDN U1154 ( .A(n54634), .B(n971), .Z(n972) );
  NAND U1155 ( .A(n54635), .B(n972), .Z(n973) );
  NANDN U1156 ( .A(n54636), .B(n973), .Z(n974) );
  AND U1157 ( .A(n52080), .B(n974), .Z(n975) );
  OR U1158 ( .A(n54637), .B(n975), .Z(n976) );
  ANDN U1159 ( .B(n976), .A(n54638), .Z(n977) );
  NANDN U1160 ( .A(n977), .B(n54639), .Z(n978) );
  NANDN U1161 ( .A(n54640), .B(n978), .Z(n979) );
  NAND U1162 ( .A(n52079), .B(n979), .Z(n54643) );
  NAND U1163 ( .A(n54687), .B(n54688), .Z(n980) );
  NAND U1164 ( .A(n54689), .B(n980), .Z(n981) );
  AND U1165 ( .A(n54690), .B(n981), .Z(n982) );
  NANDN U1166 ( .A(n982), .B(n54691), .Z(n983) );
  NANDN U1167 ( .A(n54692), .B(n983), .Z(n984) );
  NANDN U1168 ( .A(n54693), .B(n984), .Z(n985) );
  NAND U1169 ( .A(n54694), .B(n985), .Z(n986) );
  NANDN U1170 ( .A(n54695), .B(n986), .Z(n987) );
  AND U1171 ( .A(n52069), .B(n987), .Z(n988) );
  OR U1172 ( .A(n54696), .B(n988), .Z(n989) );
  AND U1173 ( .A(n54697), .B(n989), .Z(n990) );
  OR U1174 ( .A(n54698), .B(n990), .Z(n991) );
  NAND U1175 ( .A(n54699), .B(n991), .Z(n992) );
  NANDN U1176 ( .A(n52068), .B(n992), .Z(n54700) );
  AND U1177 ( .A(n52058), .B(n52059), .Z(n993) );
  NANDN U1178 ( .A(n54720), .B(n54719), .Z(n994) );
  NAND U1179 ( .A(n993), .B(n994), .Z(n995) );
  NANDN U1180 ( .A(n54721), .B(n995), .Z(n996) );
  NAND U1181 ( .A(n54722), .B(n996), .Z(n997) );
  ANDN U1182 ( .B(n997), .A(n54723), .Z(n998) );
  NANDN U1183 ( .A(n998), .B(n54724), .Z(n999) );
  NANDN U1184 ( .A(n54725), .B(n999), .Z(n1000) );
  NAND U1185 ( .A(n54726), .B(n1000), .Z(n1001) );
  NANDN U1186 ( .A(n54727), .B(n1001), .Z(n1002) );
  NAND U1187 ( .A(n54728), .B(n1002), .Z(n1003) );
  AND U1188 ( .A(n54729), .B(n1003), .Z(n1004) );
  NANDN U1189 ( .A(n1004), .B(n54730), .Z(n1005) );
  NANDN U1190 ( .A(n54731), .B(n1005), .Z(n1006) );
  NANDN U1191 ( .A(n54732), .B(n1006), .Z(n54733) );
  NANDN U1192 ( .A(n54765), .B(n54764), .Z(n1007) );
  NAND U1193 ( .A(n54766), .B(n1007), .Z(n1008) );
  AND U1194 ( .A(n54767), .B(n1008), .Z(n1009) );
  OR U1195 ( .A(n52052), .B(n1009), .Z(n1010) );
  NAND U1196 ( .A(n54768), .B(n1010), .Z(n1011) );
  NANDN U1197 ( .A(n54769), .B(n1011), .Z(n1012) );
  NAND U1198 ( .A(n54770), .B(n1012), .Z(n1013) );
  NANDN U1199 ( .A(n54771), .B(n1013), .Z(n1014) );
  AND U1200 ( .A(n54772), .B(n1014), .Z(n1015) );
  OR U1201 ( .A(n1015), .B(n54773), .Z(n1016) );
  NANDN U1202 ( .A(n54774), .B(n1016), .Z(n1017) );
  AND U1203 ( .A(n54775), .B(n1017), .Z(n1018) );
  OR U1204 ( .A(n1018), .B(n54776), .Z(n1019) );
  NAND U1205 ( .A(n54777), .B(n1019), .Z(n1020) );
  ANDN U1206 ( .B(n1020), .A(n54778), .Z(n1021) );
  OR U1207 ( .A(n1021), .B(n54779), .Z(n1022) );
  NAND U1208 ( .A(n54780), .B(n1022), .Z(n1023) );
  NANDN U1209 ( .A(n54781), .B(n1023), .Z(n1024) );
  NAND U1210 ( .A(n54782), .B(n1024), .Z(n54783) );
  NAND U1211 ( .A(n54810), .B(n52045), .Z(n1025) );
  NANDN U1212 ( .A(n54811), .B(n1025), .Z(n1026) );
  AND U1213 ( .A(n54812), .B(n1026), .Z(n1027) );
  OR U1214 ( .A(n1027), .B(n52044), .Z(n1028) );
  NANDN U1215 ( .A(n54813), .B(n1028), .Z(n1029) );
  AND U1216 ( .A(n52043), .B(n1029), .Z(n1030) );
  OR U1217 ( .A(n54814), .B(n1030), .Z(n1031) );
  AND U1218 ( .A(n54815), .B(n1031), .Z(n1032) );
  OR U1219 ( .A(n1032), .B(n52042), .Z(n1033) );
  NANDN U1220 ( .A(n54816), .B(n1033), .Z(n1034) );
  NAND U1221 ( .A(n52041), .B(n1034), .Z(n54819) );
  AND U1222 ( .A(n54838), .B(n54837), .Z(n1035) );
  NANDN U1223 ( .A(n54835), .B(n54834), .Z(n1036) );
  NAND U1224 ( .A(n1035), .B(n1036), .Z(n1037) );
  NAND U1225 ( .A(n54839), .B(n1037), .Z(n1038) );
  NANDN U1226 ( .A(n54840), .B(n1038), .Z(n1039) );
  AND U1227 ( .A(n54841), .B(n1039), .Z(n1040) );
  OR U1228 ( .A(n1040), .B(n54842), .Z(n1041) );
  NANDN U1229 ( .A(n54843), .B(n1041), .Z(n1042) );
  AND U1230 ( .A(n54844), .B(n1042), .Z(n1043) );
  OR U1231 ( .A(n1043), .B(n54845), .Z(n1044) );
  NAND U1232 ( .A(n54846), .B(n1044), .Z(n1045) );
  ANDN U1233 ( .B(n1045), .A(n54847), .Z(n1046) );
  OR U1234 ( .A(n54848), .B(n1046), .Z(n1047) );
  NAND U1235 ( .A(n54849), .B(n1047), .Z(n1048) );
  NANDN U1236 ( .A(n52027), .B(n1048), .Z(n1049) );
  NAND U1237 ( .A(n52026), .B(n1049), .Z(n54850) );
  NANDN U1238 ( .A(n55015), .B(n55014), .Z(n1050) );
  NAND U1239 ( .A(n55016), .B(n1050), .Z(n1051) );
  ANDN U1240 ( .B(n1051), .A(n55017), .Z(n1052) );
  NANDN U1241 ( .A(n1052), .B(n52014), .Z(n1053) );
  NANDN U1242 ( .A(n55018), .B(n1053), .Z(n1054) );
  NANDN U1243 ( .A(n55019), .B(n1054), .Z(n1055) );
  NAND U1244 ( .A(n55020), .B(n1055), .Z(n1056) );
  NANDN U1245 ( .A(n55021), .B(n1056), .Z(n1057) );
  AND U1246 ( .A(n55022), .B(n1057), .Z(n1058) );
  OR U1247 ( .A(n1058), .B(n55023), .Z(n1059) );
  NANDN U1248 ( .A(n55024), .B(n1059), .Z(n1060) );
  AND U1249 ( .A(n55025), .B(n1060), .Z(n1061) );
  OR U1250 ( .A(n1061), .B(n55026), .Z(n1062) );
  AND U1251 ( .A(n55027), .B(n1062), .Z(n1063) );
  AND U1252 ( .A(n55029), .B(n55030), .Z(n1064) );
  OR U1253 ( .A(n1063), .B(n55028), .Z(n1065) );
  NAND U1254 ( .A(n1064), .B(n1065), .Z(n55031) );
  NANDN U1255 ( .A(n55059), .B(n55058), .Z(n1066) );
  NANDN U1256 ( .A(n55060), .B(n1066), .Z(n1067) );
  AND U1257 ( .A(n55061), .B(n1067), .Z(n1068) );
  OR U1258 ( .A(n52008), .B(n1068), .Z(n1069) );
  NAND U1259 ( .A(n52007), .B(n1069), .Z(n1070) );
  NANDN U1260 ( .A(n55062), .B(n1070), .Z(n1071) );
  NANDN U1261 ( .A(n55063), .B(n1071), .Z(n1072) );
  NAND U1262 ( .A(n55064), .B(n1072), .Z(n1073) );
  AND U1263 ( .A(n55065), .B(n1073), .Z(n1074) );
  OR U1264 ( .A(n1074), .B(n55066), .Z(n1075) );
  NAND U1265 ( .A(n52006), .B(n1075), .Z(n1076) );
  NANDN U1266 ( .A(n55067), .B(n1076), .Z(n1077) );
  NAND U1267 ( .A(n55068), .B(n1077), .Z(n55069) );
  NAND U1268 ( .A(n55089), .B(n55090), .Z(n1078) );
  NANDN U1269 ( .A(n55091), .B(n1078), .Z(n1079) );
  NAND U1270 ( .A(n51996), .B(n1079), .Z(n1080) );
  NANDN U1271 ( .A(n55092), .B(n1080), .Z(n1081) );
  NAND U1272 ( .A(n55093), .B(n1081), .Z(n1082) );
  ANDN U1273 ( .B(n1082), .A(n51995), .Z(n1083) );
  NANDN U1274 ( .A(n1083), .B(n51994), .Z(n1084) );
  NAND U1275 ( .A(n55094), .B(n1084), .Z(n1085) );
  NAND U1276 ( .A(n51993), .B(n1085), .Z(n1086) );
  NANDN U1277 ( .A(n55095), .B(n1086), .Z(n1087) );
  NAND U1278 ( .A(n55096), .B(n1087), .Z(n1088) );
  ANDN U1279 ( .B(n1088), .A(n55097), .Z(n55100) );
  NANDN U1280 ( .A(n55131), .B(n55130), .Z(n1089) );
  NAND U1281 ( .A(n55132), .B(n1089), .Z(n1090) );
  ANDN U1282 ( .B(n1090), .A(n55133), .Z(n1091) );
  NANDN U1283 ( .A(n1091), .B(n55134), .Z(n1092) );
  NANDN U1284 ( .A(n55135), .B(n1092), .Z(n1093) );
  NANDN U1285 ( .A(n55136), .B(n1093), .Z(n1094) );
  NAND U1286 ( .A(n55137), .B(n1094), .Z(n1095) );
  NANDN U1287 ( .A(n55138), .B(n1095), .Z(n1096) );
  AND U1288 ( .A(n55139), .B(n1096), .Z(n1097) );
  OR U1289 ( .A(n1097), .B(n55140), .Z(n1098) );
  NANDN U1290 ( .A(n55141), .B(n1098), .Z(n1099) );
  AND U1291 ( .A(n55142), .B(n1099), .Z(n1100) );
  OR U1292 ( .A(n1100), .B(n55143), .Z(n1101) );
  NAND U1293 ( .A(n55144), .B(n1101), .Z(n1102) );
  AND U1294 ( .A(n55145), .B(n1102), .Z(n1103) );
  NAND U1295 ( .A(n55146), .B(n1103), .Z(n1104) );
  NANDN U1296 ( .A(n55147), .B(n1104), .Z(n1105) );
  NAND U1297 ( .A(n55148), .B(n1105), .Z(n1106) );
  NANDN U1298 ( .A(n55149), .B(n1106), .Z(n55150) );
  NAND U1299 ( .A(n55178), .B(n55177), .Z(n1107) );
  NAND U1300 ( .A(n55179), .B(n1107), .Z(n1108) );
  ANDN U1301 ( .B(n1108), .A(n55180), .Z(n1109) );
  NANDN U1302 ( .A(n1109), .B(n55181), .Z(n1110) );
  NANDN U1303 ( .A(n55182), .B(n1110), .Z(n1111) );
  NANDN U1304 ( .A(n55183), .B(n1111), .Z(n1112) );
  NAND U1305 ( .A(n55184), .B(n1112), .Z(n1113) );
  NANDN U1306 ( .A(n55185), .B(n1113), .Z(n1114) );
  AND U1307 ( .A(n55186), .B(n1114), .Z(n1115) );
  OR U1308 ( .A(n1115), .B(n55187), .Z(n1116) );
  NANDN U1309 ( .A(n55188), .B(n1116), .Z(n1117) );
  AND U1310 ( .A(n55189), .B(n1117), .Z(n1118) );
  OR U1311 ( .A(n1118), .B(n55190), .Z(n1119) );
  NAND U1312 ( .A(n51981), .B(n1119), .Z(n1120) );
  ANDN U1313 ( .B(n1120), .A(n55191), .Z(n1121) );
  OR U1314 ( .A(n55192), .B(n1121), .Z(n1122) );
  AND U1315 ( .A(n55193), .B(n1122), .Z(n55194) );
  NAND U1316 ( .A(n55289), .B(n55288), .Z(n1123) );
  NANDN U1317 ( .A(n55290), .B(n1123), .Z(n1124) );
  NAND U1318 ( .A(n51975), .B(n1124), .Z(n1125) );
  NANDN U1319 ( .A(n55291), .B(n1125), .Z(n1126) );
  NAND U1320 ( .A(n55292), .B(n1126), .Z(n1127) );
  ANDN U1321 ( .B(n1127), .A(n51974), .Z(n1128) );
  OR U1322 ( .A(n1128), .B(n55293), .Z(n1129) );
  NAND U1323 ( .A(n51973), .B(n1129), .Z(n1130) );
  ANDN U1324 ( .B(n1130), .A(n55294), .Z(n1131) );
  NANDN U1325 ( .A(n1131), .B(n55295), .Z(n1132) );
  NANDN U1326 ( .A(n51972), .B(n1132), .Z(n1133) );
  NANDN U1327 ( .A(n55296), .B(n1133), .Z(n55297) );
  NAND U1328 ( .A(n55361), .B(n55362), .Z(n1134) );
  NANDN U1329 ( .A(n55363), .B(n1134), .Z(n1135) );
  AND U1330 ( .A(n55364), .B(n1135), .Z(n1136) );
  OR U1331 ( .A(n55365), .B(n1136), .Z(n1137) );
  NANDN U1332 ( .A(n55366), .B(n1137), .Z(n1138) );
  NAND U1333 ( .A(n55367), .B(n1138), .Z(n1139) );
  NANDN U1334 ( .A(n55368), .B(n1139), .Z(n1140) );
  NAND U1335 ( .A(n55369), .B(n1140), .Z(n1141) );
  AND U1336 ( .A(n55370), .B(n1141), .Z(n1142) );
  OR U1337 ( .A(n55371), .B(n1142), .Z(n1143) );
  NAND U1338 ( .A(n55372), .B(n1143), .Z(n1144) );
  NANDN U1339 ( .A(n55373), .B(n1144), .Z(n1145) );
  NAND U1340 ( .A(n55374), .B(n1145), .Z(n1146) );
  NANDN U1341 ( .A(n55375), .B(n1146), .Z(n1147) );
  AND U1342 ( .A(n55376), .B(n1147), .Z(n1148) );
  OR U1343 ( .A(n55377), .B(n1148), .Z(n1149) );
  NANDN U1344 ( .A(n55378), .B(n1149), .Z(n1150) );
  NAND U1345 ( .A(n55379), .B(n1150), .Z(n1151) );
  NANDN U1346 ( .A(n55380), .B(n1151), .Z(n55381) );
  AND U1347 ( .A(n55417), .B(n55416), .Z(n1152) );
  NAND U1348 ( .A(n51961), .B(n1152), .Z(n1153) );
  AND U1349 ( .A(n55418), .B(n1153), .Z(n1154) );
  NOR U1350 ( .A(n1154), .B(n55420), .Z(n1155) );
  NAND U1351 ( .A(n55419), .B(n1155), .Z(n1156) );
  AND U1352 ( .A(n55421), .B(n1156), .Z(n1157) );
  OR U1353 ( .A(n1157), .B(n55422), .Z(n1158) );
  NAND U1354 ( .A(n55423), .B(n1158), .Z(n1159) );
  ANDN U1355 ( .B(n1159), .A(n55424), .Z(n1160) );
  OR U1356 ( .A(n1160), .B(n55425), .Z(n1161) );
  NAND U1357 ( .A(n55426), .B(n1161), .Z(n1162) );
  NANDN U1358 ( .A(n55427), .B(n1162), .Z(n1163) );
  NAND U1359 ( .A(n55428), .B(n1163), .Z(n1164) );
  NANDN U1360 ( .A(n55429), .B(n1164), .Z(n1165) );
  ANDN U1361 ( .B(n1165), .A(n55430), .Z(n1166) );
  NANDN U1362 ( .A(n1166), .B(n55431), .Z(n1167) );
  NANDN U1363 ( .A(n55432), .B(n1167), .Z(n1168) );
  NAND U1364 ( .A(n55433), .B(n1168), .Z(n1169) );
  NANDN U1365 ( .A(n55434), .B(n1169), .Z(n55435) );
  NANDN U1366 ( .A(n55454), .B(n55453), .Z(n1170) );
  NAND U1367 ( .A(n55455), .B(n1170), .Z(n1171) );
  ANDN U1368 ( .B(n1171), .A(n55456), .Z(n1172) );
  NANDN U1369 ( .A(n1172), .B(n55457), .Z(n1173) );
  NANDN U1370 ( .A(n55458), .B(n1173), .Z(n1174) );
  NAND U1371 ( .A(n51947), .B(n1174), .Z(n1175) );
  NANDN U1372 ( .A(n55459), .B(n1175), .Z(n1176) );
  NAND U1373 ( .A(n55460), .B(n1176), .Z(n1177) );
  ANDN U1374 ( .B(n1177), .A(n51946), .Z(n1178) );
  NANDN U1375 ( .A(n1178), .B(n51945), .Z(n1179) );
  NANDN U1376 ( .A(n55461), .B(n1179), .Z(n1180) );
  NANDN U1377 ( .A(n55462), .B(n1180), .Z(n1181) );
  NAND U1378 ( .A(n55463), .B(n1181), .Z(n55464) );
  NAND U1379 ( .A(n55490), .B(n55489), .Z(n1182) );
  NAND U1380 ( .A(n55491), .B(n1182), .Z(n1183) );
  ANDN U1381 ( .B(n1183), .A(n51936), .Z(n1184) );
  OR U1382 ( .A(n1184), .B(n55492), .Z(n1185) );
  NAND U1383 ( .A(n51935), .B(n1185), .Z(n1186) );
  NANDN U1384 ( .A(n55493), .B(n1186), .Z(n1187) );
  NAND U1385 ( .A(n55494), .B(n1187), .Z(n1188) );
  NANDN U1386 ( .A(n51934), .B(n1188), .Z(n1189) );
  ANDN U1387 ( .B(n1189), .A(n55495), .Z(n1190) );
  NANDN U1388 ( .A(n1190), .B(n51933), .Z(n1191) );
  NANDN U1389 ( .A(n55496), .B(n1191), .Z(n1192) );
  NAND U1390 ( .A(n55497), .B(n1192), .Z(n55498) );
  NAND U1391 ( .A(n55521), .B(n51925), .Z(n1193) );
  NANDN U1392 ( .A(n55522), .B(n1193), .Z(n1194) );
  ANDN U1393 ( .B(n1194), .A(n55523), .Z(n1195) );
  NANDN U1394 ( .A(n1195), .B(n55524), .Z(n1196) );
  NANDN U1395 ( .A(n55525), .B(n1196), .Z(n1197) );
  NAND U1396 ( .A(n51924), .B(n1197), .Z(n1198) );
  NANDN U1397 ( .A(n55526), .B(n1198), .Z(n1199) );
  NANDN U1398 ( .A(n55527), .B(n1199), .Z(n1200) );
  AND U1399 ( .A(n55528), .B(n1200), .Z(n1201) );
  OR U1400 ( .A(n1201), .B(n55529), .Z(n1202) );
  AND U1401 ( .A(n51923), .B(n1202), .Z(n1203) );
  OR U1402 ( .A(n55530), .B(n1203), .Z(n1204) );
  NANDN U1403 ( .A(n55531), .B(n1204), .Z(n1205) );
  NAND U1404 ( .A(n55532), .B(n1205), .Z(n55533) );
  NAND U1405 ( .A(n55553), .B(n51914), .Z(n1206) );
  NANDN U1406 ( .A(n55554), .B(n1206), .Z(n1207) );
  AND U1407 ( .A(n55555), .B(n1207), .Z(n1208) );
  OR U1408 ( .A(n51913), .B(n1208), .Z(n1209) );
  NANDN U1409 ( .A(n55556), .B(n1209), .Z(n1210) );
  NAND U1410 ( .A(n55557), .B(n1210), .Z(n1211) );
  NANDN U1411 ( .A(n55558), .B(n1211), .Z(n1212) );
  NAND U1412 ( .A(n55559), .B(n1212), .Z(n1213) );
  ANDN U1413 ( .B(n1213), .A(n51912), .Z(n1214) );
  OR U1414 ( .A(n1214), .B(n55560), .Z(n1215) );
  NAND U1415 ( .A(n55561), .B(n1215), .Z(n1216) );
  NANDN U1416 ( .A(n55562), .B(n1216), .Z(n1217) );
  NAND U1417 ( .A(n55563), .B(n1217), .Z(n55564) );
  OR U1418 ( .A(n55581), .B(n55582), .Z(n1218) );
  NANDN U1419 ( .A(n51899), .B(n1218), .Z(n1219) );
  NAND U1420 ( .A(n51898), .B(n1219), .Z(n1220) );
  NANDN U1421 ( .A(n55583), .B(n1220), .Z(n1221) );
  NANDN U1422 ( .A(n55584), .B(n1221), .Z(n1222) );
  AND U1423 ( .A(n55585), .B(n1222), .Z(n1223) );
  OR U1424 ( .A(n1223), .B(n55586), .Z(n1224) );
  NAND U1425 ( .A(n55587), .B(n1224), .Z(n1225) );
  ANDN U1426 ( .B(n1225), .A(n55588), .Z(n1226) );
  OR U1427 ( .A(n55589), .B(n1226), .Z(n1227) );
  NAND U1428 ( .A(n55590), .B(n1227), .Z(n1228) );
  NANDN U1429 ( .A(n51897), .B(n1228), .Z(n1229) );
  NAND U1430 ( .A(n51896), .B(n1229), .Z(n55591) );
  NAND U1431 ( .A(n55614), .B(n55613), .Z(n1230) );
  NANDN U1432 ( .A(n55616), .B(n1230), .Z(n1231) );
  NANDN U1433 ( .A(n51887), .B(n1231), .Z(n1232) );
  NAND U1434 ( .A(n51886), .B(n1232), .Z(n1233) );
  AND U1435 ( .A(n55618), .B(n1233), .Z(n1234) );
  NAND U1436 ( .A(n1234), .B(n55617), .Z(n1235) );
  AND U1437 ( .A(n55620), .B(n55621), .Z(n1236) );
  NANDN U1438 ( .A(n55619), .B(n1235), .Z(n1237) );
  NAND U1439 ( .A(n1236), .B(n1237), .Z(n1238) );
  NANDN U1440 ( .A(n55622), .B(n1238), .Z(n1239) );
  NAND U1441 ( .A(n55623), .B(n1239), .Z(n1240) );
  ANDN U1442 ( .B(n1240), .A(n55624), .Z(n1241) );
  NANDN U1443 ( .A(n1241), .B(n55625), .Z(n1242) );
  NANDN U1444 ( .A(n55626), .B(n1242), .Z(n1243) );
  NAND U1445 ( .A(n51885), .B(n1243), .Z(n1244) );
  ANDN U1446 ( .B(n1244), .A(n55627), .Z(n55630) );
  NAND U1447 ( .A(n55778), .B(n55779), .Z(n1245) );
  NANDN U1448 ( .A(n55780), .B(n1245), .Z(n1246) );
  ANDN U1449 ( .B(n1246), .A(n55781), .Z(n1247) );
  NANDN U1450 ( .A(n1247), .B(n55782), .Z(n1248) );
  NANDN U1451 ( .A(n51876), .B(n1248), .Z(n1249) );
  NAND U1452 ( .A(n51875), .B(n1249), .Z(n1250) );
  NANDN U1453 ( .A(n51874), .B(n1250), .Z(n1251) );
  NANDN U1454 ( .A(n55783), .B(n1251), .Z(n1252) );
  AND U1455 ( .A(n55784), .B(n1252), .Z(n1253) );
  OR U1456 ( .A(n1253), .B(n55785), .Z(n1254) );
  NAND U1457 ( .A(n55786), .B(n1254), .Z(n1255) );
  ANDN U1458 ( .B(n1255), .A(n55787), .Z(n1256) );
  OR U1459 ( .A(n1256), .B(n55788), .Z(n1257) );
  NAND U1460 ( .A(n55789), .B(n1257), .Z(n1258) );
  NANDN U1461 ( .A(n55790), .B(n1258), .Z(n55791) );
  ANDN U1462 ( .B(n55813), .A(n55816), .Z(n1259) );
  NAND U1463 ( .A(n55814), .B(n1259), .Z(n1260) );
  AND U1464 ( .A(n55817), .B(n1260), .Z(n1261) );
  OR U1465 ( .A(n55818), .B(n1261), .Z(n1262) );
  NAND U1466 ( .A(n55819), .B(n1262), .Z(n1263) );
  NANDN U1467 ( .A(n51863), .B(n1263), .Z(n1264) );
  NAND U1468 ( .A(n51862), .B(n1264), .Z(n1265) );
  NANDN U1469 ( .A(n55820), .B(n1265), .Z(n1266) );
  AND U1470 ( .A(n55821), .B(n1266), .Z(n1267) );
  OR U1471 ( .A(n1267), .B(n55822), .Z(n1268) );
  NAND U1472 ( .A(n55823), .B(n1268), .Z(n1269) );
  AND U1473 ( .A(n51861), .B(n1269), .Z(n1270) );
  OR U1474 ( .A(n1270), .B(n55824), .Z(n1271) );
  NAND U1475 ( .A(n55825), .B(n1271), .Z(n1272) );
  NANDN U1476 ( .A(n55826), .B(n1272), .Z(n1273) );
  NAND U1477 ( .A(n55827), .B(n1273), .Z(n55828) );
  NAND U1478 ( .A(n55861), .B(n55862), .Z(n1274) );
  NAND U1479 ( .A(n55863), .B(n1274), .Z(n1275) );
  NANDN U1480 ( .A(n51856), .B(n1275), .Z(n1276) );
  NAND U1481 ( .A(n51855), .B(n1276), .Z(n1277) );
  NANDN U1482 ( .A(n55864), .B(n1277), .Z(n1278) );
  AND U1483 ( .A(n55865), .B(n1278), .Z(n1279) );
  OR U1484 ( .A(n1279), .B(n55866), .Z(n1280) );
  NAND U1485 ( .A(n55867), .B(n1280), .Z(n1281) );
  AND U1486 ( .A(n51854), .B(n1281), .Z(n1282) );
  OR U1487 ( .A(n1282), .B(n55868), .Z(n1283) );
  NAND U1488 ( .A(n55869), .B(n1283), .Z(n1284) );
  ANDN U1489 ( .B(n1284), .A(n55870), .Z(n1285) );
  NANDN U1490 ( .A(n1285), .B(n55871), .Z(n1286) );
  NANDN U1491 ( .A(n55872), .B(n1286), .Z(n1287) );
  NAND U1492 ( .A(n55873), .B(n1287), .Z(n1288) );
  NANDN U1493 ( .A(n55874), .B(n1288), .Z(n55875) );
  NANDN U1494 ( .A(n55891), .B(n55890), .Z(n1289) );
  NAND U1495 ( .A(n55893), .B(n1289), .Z(n1290) );
  NAND U1496 ( .A(n55894), .B(n1290), .Z(n1291) );
  NANDN U1497 ( .A(n55895), .B(n1291), .Z(n1292) );
  NAND U1498 ( .A(n55896), .B(n1292), .Z(n1293) );
  ANDN U1499 ( .B(n1293), .A(n51841), .Z(n1294) );
  NANDN U1500 ( .A(n1294), .B(n51840), .Z(n1295) );
  ANDN U1501 ( .B(n1295), .A(n55897), .Z(n1296) );
  NANDN U1502 ( .A(n1296), .B(n55898), .Z(n1297) );
  NANDN U1503 ( .A(n51839), .B(n1297), .Z(n1298) );
  NAND U1504 ( .A(n51838), .B(n1298), .Z(n55901) );
  NANDN U1505 ( .A(n55923), .B(n55922), .Z(n1299) );
  NANDN U1506 ( .A(n51832), .B(n1299), .Z(n1300) );
  NAND U1507 ( .A(n51831), .B(n1300), .Z(n1301) );
  NANDN U1508 ( .A(n55924), .B(n1301), .Z(n1302) );
  NAND U1509 ( .A(n55925), .B(n1302), .Z(n1303) );
  ANDN U1510 ( .B(n1303), .A(n55926), .Z(n1304) );
  NANDN U1511 ( .A(n1304), .B(n55927), .Z(n1305) );
  ANDN U1512 ( .B(n1305), .A(n51830), .Z(n1306) );
  NANDN U1513 ( .A(n1306), .B(n51829), .Z(n1307) );
  NAND U1514 ( .A(n55928), .B(n1307), .Z(n1308) );
  NANDN U1515 ( .A(n51828), .B(n1308), .Z(n55929) );
  NAND U1516 ( .A(n51820), .B(n55950), .Z(n1309) );
  NANDN U1517 ( .A(n55951), .B(n1309), .Z(n1310) );
  AND U1518 ( .A(n55952), .B(n1310), .Z(n1311) );
  OR U1519 ( .A(n55953), .B(n1311), .Z(n1312) );
  NAND U1520 ( .A(n55954), .B(n1312), .Z(n1313) );
  NANDN U1521 ( .A(n51819), .B(n1313), .Z(n1314) );
  NAND U1522 ( .A(n51818), .B(n1314), .Z(n1315) );
  NAND U1523 ( .A(n55955), .B(n1315), .Z(n1316) );
  AND U1524 ( .A(n55956), .B(n1316), .Z(n1317) );
  NAND U1525 ( .A(n1317), .B(n55957), .Z(n1318) );
  NANDN U1526 ( .A(n55958), .B(n1318), .Z(n1319) );
  AND U1527 ( .A(n55959), .B(n1319), .Z(n1320) );
  OR U1528 ( .A(n55960), .B(n1320), .Z(n1321) );
  AND U1529 ( .A(n55961), .B(n1321), .Z(n55962) );
  NANDN U1530 ( .A(n55989), .B(n55988), .Z(n1322) );
  NANDN U1531 ( .A(n55990), .B(n1322), .Z(n1323) );
  NAND U1532 ( .A(n55991), .B(n1323), .Z(n1324) );
  NANDN U1533 ( .A(n51810), .B(n1324), .Z(n1325) );
  NAND U1534 ( .A(n51809), .B(n1325), .Z(n1326) );
  ANDN U1535 ( .B(n1326), .A(n55992), .Z(n1327) );
  NANDN U1536 ( .A(n1327), .B(n55993), .Z(n1328) );
  AND U1537 ( .A(n51808), .B(n1328), .Z(n1329) );
  OR U1538 ( .A(n55994), .B(n1329), .Z(n1330) );
  NAND U1539 ( .A(n55995), .B(n1330), .Z(n1331) );
  NANDN U1540 ( .A(n51807), .B(n1331), .Z(n55996) );
  NAND U1541 ( .A(n56018), .B(n51799), .Z(n1332) );
  ANDN U1542 ( .B(n1332), .A(n56019), .Z(n1333) );
  ANDN U1543 ( .B(n56021), .A(n1333), .Z(n1334) );
  NAND U1544 ( .A(n56020), .B(n1334), .Z(n1335) );
  NANDN U1545 ( .A(n56022), .B(n1335), .Z(n1336) );
  ANDN U1546 ( .B(n56023), .A(n56024), .Z(n1337) );
  NAND U1547 ( .A(n1336), .B(n1337), .Z(n1338) );
  NANDN U1548 ( .A(n56025), .B(n1338), .Z(n1339) );
  ANDN U1549 ( .B(n56027), .A(n56026), .Z(n1340) );
  NAND U1550 ( .A(n1339), .B(n1340), .Z(n1341) );
  NANDN U1551 ( .A(n56028), .B(n1341), .Z(n1342) );
  NAND U1552 ( .A(n56029), .B(n1342), .Z(n1343) );
  NANDN U1553 ( .A(n56030), .B(n1343), .Z(n1344) );
  AND U1554 ( .A(n56031), .B(n1344), .Z(n1345) );
  OR U1555 ( .A(n56032), .B(n1345), .Z(n1346) );
  AND U1556 ( .A(n56033), .B(n1346), .Z(n56035) );
  OR U1557 ( .A(n56062), .B(n56063), .Z(n1347) );
  NAND U1558 ( .A(n56064), .B(n1347), .Z(n1348) );
  ANDN U1559 ( .B(n1348), .A(n56065), .Z(n1349) );
  NANDN U1560 ( .A(n1349), .B(n56066), .Z(n1350) );
  NANDN U1561 ( .A(n56067), .B(n1350), .Z(n1351) );
  NAND U1562 ( .A(n51793), .B(n1351), .Z(n1352) );
  NANDN U1563 ( .A(n56068), .B(n1352), .Z(n1353) );
  NAND U1564 ( .A(n56069), .B(n1353), .Z(n1354) );
  ANDN U1565 ( .B(n1354), .A(n51792), .Z(n1355) );
  NANDN U1566 ( .A(n1355), .B(n51791), .Z(n1356) );
  NANDN U1567 ( .A(n56070), .B(n1356), .Z(n1357) );
  NAND U1568 ( .A(n56071), .B(n1357), .Z(n56074) );
  NAND U1569 ( .A(n56095), .B(n56096), .Z(n1358) );
  NAND U1570 ( .A(n56097), .B(n1358), .Z(n1359) );
  NANDN U1571 ( .A(n56098), .B(n1359), .Z(n1360) );
  NAND U1572 ( .A(n56099), .B(n1360), .Z(n1361) );
  NANDN U1573 ( .A(n51781), .B(n1361), .Z(n1362) );
  AND U1574 ( .A(n56100), .B(n1362), .Z(n1363) );
  NOR U1575 ( .A(n56102), .B(n1363), .Z(n1364) );
  NAND U1576 ( .A(n56101), .B(n1364), .Z(n1365) );
  AND U1577 ( .A(n56103), .B(n1365), .Z(n1366) );
  OR U1578 ( .A(n56104), .B(n1366), .Z(n1367) );
  NAND U1579 ( .A(n56105), .B(n1367), .Z(n1368) );
  NANDN U1580 ( .A(n51780), .B(n1368), .Z(n56106) );
  NAND U1581 ( .A(n56133), .B(n56134), .Z(n1369) );
  NANDN U1582 ( .A(n56135), .B(n1369), .Z(n1370) );
  AND U1583 ( .A(n56136), .B(n1370), .Z(n1371) );
  NAND U1584 ( .A(n1371), .B(n56137), .Z(n1372) );
  NANDN U1585 ( .A(n56138), .B(n1372), .Z(n1373) );
  AND U1586 ( .A(n56139), .B(n1373), .Z(n1374) );
  OR U1587 ( .A(n1374), .B(n56140), .Z(n1375) );
  NAND U1588 ( .A(n56141), .B(n1375), .Z(n1376) );
  AND U1589 ( .A(n51772), .B(n1376), .Z(n1377) );
  OR U1590 ( .A(n56142), .B(n1377), .Z(n1378) );
  AND U1591 ( .A(n56143), .B(n1378), .Z(n1379) );
  OR U1592 ( .A(n56144), .B(n1379), .Z(n1380) );
  NAND U1593 ( .A(n56145), .B(n1380), .Z(n1381) );
  NANDN U1594 ( .A(n51771), .B(n1381), .Z(n56146) );
  NANDN U1595 ( .A(n56170), .B(n56169), .Z(n1382) );
  NAND U1596 ( .A(n56172), .B(n1382), .Z(n1383) );
  AND U1597 ( .A(n56173), .B(n1383), .Z(n1384) );
  NANDN U1598 ( .A(n1384), .B(n56174), .Z(n1385) );
  NAND U1599 ( .A(n56175), .B(n1385), .Z(n1386) );
  NANDN U1600 ( .A(n56176), .B(n1386), .Z(n1387) );
  AND U1601 ( .A(n51762), .B(n51761), .Z(n1388) );
  NAND U1602 ( .A(n1387), .B(n1388), .Z(n1389) );
  NANDN U1603 ( .A(n56177), .B(n1389), .Z(n1390) );
  AND U1604 ( .A(n56179), .B(n56178), .Z(n1391) );
  NAND U1605 ( .A(n1390), .B(n1391), .Z(n1392) );
  NANDN U1606 ( .A(n56180), .B(n1392), .Z(n1393) );
  NAND U1607 ( .A(n56181), .B(n1393), .Z(n56182) );
  NAND U1608 ( .A(n56209), .B(n56208), .Z(n1394) );
  NANDN U1609 ( .A(n56210), .B(n1394), .Z(n1395) );
  AND U1610 ( .A(n56211), .B(n1395), .Z(n1396) );
  OR U1611 ( .A(n1396), .B(n56212), .Z(n1397) );
  NAND U1612 ( .A(n56213), .B(n1397), .Z(n1398) );
  NANDN U1613 ( .A(n56214), .B(n1398), .Z(n1399) );
  NAND U1614 ( .A(n56215), .B(n1399), .Z(n1400) );
  NAND U1615 ( .A(n56216), .B(n1400), .Z(n1401) );
  ANDN U1616 ( .B(n1401), .A(n56217), .Z(n1402) );
  NANDN U1617 ( .A(n1402), .B(n56218), .Z(n1403) );
  ANDN U1618 ( .B(n1403), .A(n51751), .Z(n1404) );
  NANDN U1619 ( .A(n1404), .B(n51750), .Z(n1405) );
  NANDN U1620 ( .A(n56219), .B(n1405), .Z(n1406) );
  NAND U1621 ( .A(n56220), .B(n1406), .Z(n56221) );
  NANDN U1622 ( .A(n56248), .B(n56247), .Z(n1407) );
  NAND U1623 ( .A(n56250), .B(n1407), .Z(n1408) );
  NAND U1624 ( .A(n56251), .B(n1408), .Z(n1409) );
  NANDN U1625 ( .A(n51740), .B(n1409), .Z(n1410) );
  NAND U1626 ( .A(n51739), .B(n1410), .Z(n1411) );
  ANDN U1627 ( .B(n1411), .A(n56252), .Z(n1412) );
  NANDN U1628 ( .A(n1412), .B(n56253), .Z(n1413) );
  NANDN U1629 ( .A(n56254), .B(n1413), .Z(n1414) );
  NAND U1630 ( .A(n56255), .B(n1414), .Z(n1415) );
  NANDN U1631 ( .A(n56256), .B(n1415), .Z(n1416) );
  NAND U1632 ( .A(n56257), .B(n1416), .Z(n1417) );
  ANDN U1633 ( .B(n1417), .A(n56258), .Z(n56261) );
  NANDN U1634 ( .A(n51730), .B(n56282), .Z(n1418) );
  NAND U1635 ( .A(n51729), .B(n1418), .Z(n1419) );
  ANDN U1636 ( .B(n1419), .A(n51728), .Z(n1420) );
  NANDN U1637 ( .A(n1420), .B(n56283), .Z(n1421) );
  NANDN U1638 ( .A(n51727), .B(n1421), .Z(n1422) );
  NAND U1639 ( .A(n56284), .B(n1422), .Z(n1423) );
  NANDN U1640 ( .A(n51726), .B(n1423), .Z(n1424) );
  NAND U1641 ( .A(n51725), .B(n1424), .Z(n1425) );
  AND U1642 ( .A(n56285), .B(n1425), .Z(n1426) );
  OR U1643 ( .A(n56286), .B(n1426), .Z(n1427) );
  NAND U1644 ( .A(n56287), .B(n1427), .Z(n1428) );
  NANDN U1645 ( .A(n56288), .B(n1428), .Z(n1429) );
  NAND U1646 ( .A(n56289), .B(n1429), .Z(n56290) );
  NAND U1647 ( .A(n56317), .B(n56316), .Z(n1430) );
  NAND U1648 ( .A(n51718), .B(n1430), .Z(n1431) );
  AND U1649 ( .A(n56318), .B(n1431), .Z(n1432) );
  NOR U1650 ( .A(n56319), .B(n1432), .Z(n1433) );
  NAND U1651 ( .A(n56320), .B(n1433), .Z(n1434) );
  AND U1652 ( .A(n51717), .B(n1434), .Z(n1435) );
  NOR U1653 ( .A(n56321), .B(n51716), .Z(n1436) );
  NANDN U1654 ( .A(n1435), .B(n1436), .Z(n1437) );
  AND U1655 ( .A(n51715), .B(n1437), .Z(n1438) );
  OR U1656 ( .A(n56322), .B(n1438), .Z(n1439) );
  NAND U1657 ( .A(n56323), .B(n1439), .Z(n1440) );
  NANDN U1658 ( .A(n51714), .B(n1440), .Z(n56324) );
  NANDN U1659 ( .A(n56347), .B(n56346), .Z(n1441) );
  NAND U1660 ( .A(n56348), .B(n1441), .Z(n1442) );
  ANDN U1661 ( .B(n1442), .A(n56349), .Z(n1443) );
  NANDN U1662 ( .A(n1443), .B(n56350), .Z(n1444) );
  NAND U1663 ( .A(n56351), .B(n1444), .Z(n1445) );
  NANDN U1664 ( .A(n51705), .B(n1445), .Z(n1446) );
  NAND U1665 ( .A(n51704), .B(n1446), .Z(n1447) );
  NANDN U1666 ( .A(n56352), .B(n1447), .Z(n1448) );
  AND U1667 ( .A(n56353), .B(n1448), .Z(n1449) );
  OR U1668 ( .A(n1449), .B(n56354), .Z(n1450) );
  NAND U1669 ( .A(n56355), .B(n1450), .Z(n1451) );
  NANDN U1670 ( .A(n56356), .B(n1451), .Z(n1452) );
  NAND U1671 ( .A(n56357), .B(n1452), .Z(n1453) );
  NAND U1672 ( .A(n51703), .B(n1453), .Z(n1454) );
  AND U1673 ( .A(n56358), .B(n1454), .Z(n56360) );
  NAND U1674 ( .A(n56377), .B(n56376), .Z(n1455) );
  NANDN U1675 ( .A(n56378), .B(n1455), .Z(n1456) );
  AND U1676 ( .A(n56379), .B(n1456), .Z(n1457) );
  AND U1677 ( .A(n56381), .B(n56380), .Z(n1458) );
  NANDN U1678 ( .A(n1457), .B(n51694), .Z(n1459) );
  AND U1679 ( .A(n1458), .B(n1459), .Z(n1460) );
  AND U1680 ( .A(n51692), .B(n51693), .Z(n1461) );
  OR U1681 ( .A(n56382), .B(n1460), .Z(n1462) );
  AND U1682 ( .A(n1461), .B(n1462), .Z(n1463) );
  NANDN U1683 ( .A(n1463), .B(n56383), .Z(n1464) );
  ANDN U1684 ( .B(n1464), .A(n51691), .Z(n1465) );
  NANDN U1685 ( .A(n1465), .B(n51690), .Z(n1466) );
  NANDN U1686 ( .A(n56384), .B(n1466), .Z(n1467) );
  NAND U1687 ( .A(n56385), .B(n1467), .Z(n56386) );
  NANDN U1688 ( .A(n56412), .B(n56411), .Z(n1468) );
  NAND U1689 ( .A(n56413), .B(n1468), .Z(n1469) );
  ANDN U1690 ( .B(n1469), .A(n56414), .Z(n1470) );
  NANDN U1691 ( .A(n1470), .B(n51682), .Z(n1471) );
  NANDN U1692 ( .A(n56415), .B(n1471), .Z(n1472) );
  NAND U1693 ( .A(n56416), .B(n1472), .Z(n1473) );
  NAND U1694 ( .A(n56417), .B(n1473), .Z(n1474) );
  NANDN U1695 ( .A(n56418), .B(n1474), .Z(n1475) );
  AND U1696 ( .A(n56419), .B(n1475), .Z(n1476) );
  OR U1697 ( .A(n56420), .B(n1476), .Z(n1477) );
  NAND U1698 ( .A(n56421), .B(n1477), .Z(n1478) );
  NANDN U1699 ( .A(n56422), .B(n1478), .Z(n1479) );
  NAND U1700 ( .A(n56423), .B(n1479), .Z(n1480) );
  AND U1701 ( .A(n51681), .B(n1480), .Z(n1481) );
  NANDN U1702 ( .A(n51680), .B(n1481), .Z(n56426) );
  NANDN U1703 ( .A(n56498), .B(n56497), .Z(n1482) );
  NANDN U1704 ( .A(n56499), .B(n1482), .Z(n1483) );
  AND U1705 ( .A(n56500), .B(n1483), .Z(n1484) );
  AND U1706 ( .A(n56503), .B(n56502), .Z(n1485) );
  OR U1707 ( .A(n1484), .B(n56501), .Z(n1486) );
  AND U1708 ( .A(n1485), .B(n1486), .Z(n1487) );
  OR U1709 ( .A(n56504), .B(n1487), .Z(n1488) );
  NAND U1710 ( .A(n56505), .B(n1488), .Z(n1489) );
  NAND U1711 ( .A(n56506), .B(n1489), .Z(n1490) );
  NANDN U1712 ( .A(n51671), .B(n1490), .Z(n1491) );
  NAND U1713 ( .A(n51670), .B(n1491), .Z(n1492) );
  ANDN U1714 ( .B(n1492), .A(n56507), .Z(n1493) );
  NANDN U1715 ( .A(n1493), .B(n56508), .Z(n1494) );
  NAND U1716 ( .A(n56509), .B(n1494), .Z(n1495) );
  NANDN U1717 ( .A(n56510), .B(n1495), .Z(n56511) );
  NAND U1718 ( .A(n56538), .B(n56539), .Z(n1496) );
  NAND U1719 ( .A(n56540), .B(n1496), .Z(n1497) );
  NANDN U1720 ( .A(n51663), .B(n1497), .Z(n1498) );
  NAND U1721 ( .A(n56541), .B(n1498), .Z(n1499) );
  NANDN U1722 ( .A(n56542), .B(n1499), .Z(n1500) );
  AND U1723 ( .A(n56543), .B(n1500), .Z(n1501) );
  AND U1724 ( .A(n56546), .B(n56545), .Z(n1502) );
  NANDN U1725 ( .A(n1501), .B(n56544), .Z(n1503) );
  AND U1726 ( .A(n1502), .B(n1503), .Z(n1504) );
  AND U1727 ( .A(n51662), .B(n51661), .Z(n1505) );
  OR U1728 ( .A(n56547), .B(n1504), .Z(n1506) );
  AND U1729 ( .A(n1505), .B(n1506), .Z(n1507) );
  OR U1730 ( .A(n56548), .B(n1507), .Z(n1508) );
  AND U1731 ( .A(n56549), .B(n1508), .Z(n1509) );
  OR U1732 ( .A(n56550), .B(n1509), .Z(n1510) );
  NAND U1733 ( .A(n56551), .B(n1510), .Z(n1511) );
  NANDN U1734 ( .A(n51660), .B(n1511), .Z(n56552) );
  NANDN U1735 ( .A(n56583), .B(n56582), .Z(n1512) );
  NAND U1736 ( .A(n56585), .B(n1512), .Z(n1513) );
  NAND U1737 ( .A(n56586), .B(n1513), .Z(n1514) );
  NANDN U1738 ( .A(n56587), .B(n1514), .Z(n1515) );
  NAND U1739 ( .A(n56588), .B(n1515), .Z(n1516) );
  ANDN U1740 ( .B(n1516), .A(n51654), .Z(n1517) );
  NANDN U1741 ( .A(n1517), .B(n51653), .Z(n1518) );
  ANDN U1742 ( .B(n1518), .A(n56589), .Z(n1519) );
  NANDN U1743 ( .A(n1519), .B(n56590), .Z(n1520) );
  NANDN U1744 ( .A(n51652), .B(n1520), .Z(n1521) );
  NAND U1745 ( .A(n51651), .B(n1521), .Z(n56593) );
  NAND U1746 ( .A(n56617), .B(n56616), .Z(n1522) );
  NANDN U1747 ( .A(n56619), .B(n1522), .Z(n1523) );
  ANDN U1748 ( .B(n1523), .A(n51642), .Z(n1524) );
  NANDN U1749 ( .A(n1524), .B(n51641), .Z(n1525) );
  NANDN U1750 ( .A(n56620), .B(n1525), .Z(n1526) );
  NAND U1751 ( .A(n56621), .B(n1526), .Z(n1527) );
  NANDN U1752 ( .A(n56622), .B(n1527), .Z(n1528) );
  NAND U1753 ( .A(n56623), .B(n1528), .Z(n1529) );
  ANDN U1754 ( .B(n1529), .A(n51640), .Z(n1530) );
  NANDN U1755 ( .A(n1530), .B(n51639), .Z(n1531) );
  ANDN U1756 ( .B(n1531), .A(n56624), .Z(n56626) );
  ANDN U1757 ( .B(n56652), .A(n56653), .Z(n1532) );
  NANDN U1758 ( .A(n56651), .B(n56650), .Z(n1533) );
  NAND U1759 ( .A(n1532), .B(n1533), .Z(n1534) );
  NAND U1760 ( .A(n56654), .B(n1534), .Z(n1535) );
  AND U1761 ( .A(n56656), .B(n1535), .Z(n1536) );
  NAND U1762 ( .A(n1536), .B(n56655), .Z(n1537) );
  NAND U1763 ( .A(n56657), .B(n1537), .Z(n1538) );
  NANDN U1764 ( .A(n51631), .B(n1538), .Z(n1539) );
  AND U1765 ( .A(n51630), .B(n1539), .Z(n1540) );
  OR U1766 ( .A(n56658), .B(n1540), .Z(n1541) );
  NAND U1767 ( .A(n56659), .B(n1541), .Z(n1542) );
  NANDN U1768 ( .A(n56660), .B(n1542), .Z(n1543) );
  NAND U1769 ( .A(n56661), .B(n1543), .Z(n56662) );
  NAND U1770 ( .A(n51624), .B(n56687), .Z(n1544) );
  NANDN U1771 ( .A(n51623), .B(n1544), .Z(n1545) );
  AND U1772 ( .A(n56688), .B(n1545), .Z(n1546) );
  NAND U1773 ( .A(n1546), .B(n56689), .Z(n1547) );
  NANDN U1774 ( .A(n51622), .B(n1547), .Z(n1548) );
  AND U1775 ( .A(n56690), .B(n1548), .Z(n1549) );
  OR U1776 ( .A(n51621), .B(n1549), .Z(n1550) );
  NAND U1777 ( .A(n51620), .B(n1550), .Z(n1551) );
  NANDN U1778 ( .A(n56691), .B(n1551), .Z(n1552) );
  NAND U1779 ( .A(n56692), .B(n1552), .Z(n1553) );
  NAND U1780 ( .A(n56693), .B(n1553), .Z(n1554) );
  AND U1781 ( .A(n56694), .B(n1554), .Z(n56697) );
  NANDN U1782 ( .A(n56725), .B(n56724), .Z(n1555) );
  NAND U1783 ( .A(n51611), .B(n1555), .Z(n1556) );
  AND U1784 ( .A(n56726), .B(n1556), .Z(n1557) );
  NANDN U1785 ( .A(n1557), .B(n56727), .Z(n1558) );
  NAND U1786 ( .A(n56728), .B(n1558), .Z(n1559) );
  NAND U1787 ( .A(n56729), .B(n1559), .Z(n1560) );
  NANDN U1788 ( .A(n56730), .B(n1560), .Z(n1561) );
  NAND U1789 ( .A(n56731), .B(n1561), .Z(n1562) );
  AND U1790 ( .A(n56732), .B(n1562), .Z(n1563) );
  NANDN U1791 ( .A(n1563), .B(n56733), .Z(n1564) );
  ANDN U1792 ( .B(n1564), .A(n56734), .Z(n1565) );
  NANDN U1793 ( .A(n1565), .B(n56735), .Z(n1566) );
  NANDN U1794 ( .A(n51610), .B(n1566), .Z(n1567) );
  NAND U1795 ( .A(n56736), .B(n1567), .Z(n56737) );
  NAND U1796 ( .A(n56821), .B(n56822), .Z(n1568) );
  NANDN U1797 ( .A(n56823), .B(n1568), .Z(n1569) );
  NAND U1798 ( .A(n56824), .B(n1569), .Z(n1570) );
  ANDN U1799 ( .B(n51602), .A(n51601), .Z(n1571) );
  NANDN U1800 ( .A(n56825), .B(n1570), .Z(n1572) );
  NAND U1801 ( .A(n1571), .B(n1572), .Z(n1573) );
  NAND U1802 ( .A(n56826), .B(n1573), .Z(n1574) );
  AND U1803 ( .A(n56828), .B(n1574), .Z(n1575) );
  NAND U1804 ( .A(n1575), .B(n56827), .Z(n1576) );
  ANDN U1805 ( .B(n56830), .A(n56831), .Z(n1577) );
  NANDN U1806 ( .A(n56829), .B(n1576), .Z(n1578) );
  NAND U1807 ( .A(n1577), .B(n1578), .Z(n1579) );
  ANDN U1808 ( .B(n56834), .A(n56833), .Z(n1580) );
  NANDN U1809 ( .A(n56832), .B(n1579), .Z(n1581) );
  NAND U1810 ( .A(n1580), .B(n1581), .Z(n1582) );
  NANDN U1811 ( .A(n56835), .B(n1582), .Z(n1583) );
  NAND U1812 ( .A(n56836), .B(n1583), .Z(n1584) );
  AND U1813 ( .A(n56837), .B(n1584), .Z(n56841) );
  NAND U1814 ( .A(n56872), .B(n56871), .Z(n1585) );
  NANDN U1815 ( .A(n56874), .B(n1585), .Z(n1586) );
  NANDN U1816 ( .A(n51597), .B(n1586), .Z(n1587) );
  NAND U1817 ( .A(n51596), .B(n1587), .Z(n1588) );
  NAND U1818 ( .A(n56875), .B(n1588), .Z(n1589) );
  AND U1819 ( .A(n56876), .B(n1589), .Z(n1590) );
  NAND U1820 ( .A(n1590), .B(n56877), .Z(n1591) );
  NANDN U1821 ( .A(n56878), .B(n1591), .Z(n1592) );
  AND U1822 ( .A(n56879), .B(n1592), .Z(n1593) );
  ANDN U1823 ( .B(n51594), .A(n51595), .Z(n1594) );
  OR U1824 ( .A(n56880), .B(n1593), .Z(n1595) );
  AND U1825 ( .A(n1594), .B(n1595), .Z(n1596) );
  OR U1826 ( .A(n56881), .B(n1596), .Z(n1597) );
  NAND U1827 ( .A(n56882), .B(n1597), .Z(n1598) );
  NAND U1828 ( .A(n56883), .B(n1598), .Z(n56884) );
  NANDN U1829 ( .A(n56910), .B(n56909), .Z(n1599) );
  NANDN U1830 ( .A(n56911), .B(n1599), .Z(n1600) );
  AND U1831 ( .A(n56912), .B(n1600), .Z(n1601) );
  NANDN U1832 ( .A(n1601), .B(n56913), .Z(n1602) );
  NAND U1833 ( .A(n51586), .B(n1602), .Z(n1603) );
  NANDN U1834 ( .A(n56914), .B(n1603), .Z(n1604) );
  NANDN U1835 ( .A(n1604), .B(n56915), .Z(n1605) );
  AND U1836 ( .A(n56916), .B(n1605), .Z(n1606) );
  ANDN U1837 ( .B(n51585), .A(n1606), .Z(n1607) );
  NAND U1838 ( .A(n51584), .B(n1607), .Z(n1608) );
  ANDN U1839 ( .B(n1608), .A(n56917), .Z(n1609) );
  NANDN U1840 ( .A(n1609), .B(n56918), .Z(n1610) );
  NAND U1841 ( .A(n56919), .B(n1610), .Z(n1611) );
  NAND U1842 ( .A(n51583), .B(n1611), .Z(n56921) );
  OR U1843 ( .A(n56991), .B(n56992), .Z(n1612) );
  NAND U1844 ( .A(n56993), .B(n1612), .Z(n1613) );
  NANDN U1845 ( .A(n56994), .B(n1613), .Z(n1614) );
  NAND U1846 ( .A(n56995), .B(n1614), .Z(n1615) );
  NANDN U1847 ( .A(n56996), .B(n1615), .Z(n1616) );
  AND U1848 ( .A(n56997), .B(n1616), .Z(n1617) );
  OR U1849 ( .A(n1617), .B(n56998), .Z(n1618) );
  NAND U1850 ( .A(n56999), .B(n1618), .Z(n1619) );
  ANDN U1851 ( .B(n1619), .A(n57000), .Z(n1620) );
  NANDN U1852 ( .A(n1620), .B(n57001), .Z(n1621) );
  NANDN U1853 ( .A(n57002), .B(n1621), .Z(n1622) );
  NAND U1854 ( .A(n57003), .B(n1622), .Z(n1623) );
  AND U1855 ( .A(n57005), .B(n57006), .Z(n1624) );
  NANDN U1856 ( .A(n57004), .B(n1623), .Z(n1625) );
  NAND U1857 ( .A(n1624), .B(n1625), .Z(n1626) );
  NAND U1858 ( .A(n51573), .B(n1626), .Z(n1627) );
  AND U1859 ( .A(n57007), .B(n1627), .Z(n1628) );
  NAND U1860 ( .A(n1628), .B(n57008), .Z(n1629) );
  NANDN U1861 ( .A(n57009), .B(n1629), .Z(n57010) );
  NAND U1862 ( .A(n57042), .B(n57041), .Z(n1630) );
  NANDN U1863 ( .A(n57043), .B(n1630), .Z(n1631) );
  AND U1864 ( .A(n57044), .B(n1631), .Z(n1632) );
  OR U1865 ( .A(n1632), .B(n57045), .Z(n1633) );
  NAND U1866 ( .A(n51566), .B(n1633), .Z(n1634) );
  ANDN U1867 ( .B(n1634), .A(n57046), .Z(n1635) );
  NANDN U1868 ( .A(n1635), .B(n57047), .Z(n1636) );
  NANDN U1869 ( .A(n51565), .B(n1636), .Z(n1637) );
  NAND U1870 ( .A(n51564), .B(n1637), .Z(n1638) );
  AND U1871 ( .A(n51563), .B(n57048), .Z(n1639) );
  NAND U1872 ( .A(n1638), .B(n1639), .Z(n1640) );
  NANDN U1873 ( .A(n51562), .B(n1640), .Z(n57049) );
  NAND U1874 ( .A(n57083), .B(n57082), .Z(n1641) );
  AND U1875 ( .A(n57084), .B(n1641), .Z(n1642) );
  NANDN U1876 ( .A(n51556), .B(n51557), .Z(n1643) );
  NAND U1877 ( .A(n1642), .B(n1643), .Z(n1644) );
  NANDN U1878 ( .A(n57085), .B(n1644), .Z(n1645) );
  NAND U1879 ( .A(n57086), .B(n1645), .Z(n1646) );
  NANDN U1880 ( .A(n57087), .B(n1646), .Z(n1647) );
  AND U1881 ( .A(n57088), .B(n1647), .Z(n1648) );
  OR U1882 ( .A(n57089), .B(n1648), .Z(n1649) );
  NAND U1883 ( .A(n57090), .B(n1649), .Z(n1650) );
  NANDN U1884 ( .A(n57091), .B(n1650), .Z(n1651) );
  NAND U1885 ( .A(n57092), .B(n1651), .Z(n1652) );
  NAND U1886 ( .A(n57093), .B(n1652), .Z(n1653) );
  ANDN U1887 ( .B(n1653), .A(n57094), .Z(n1654) );
  NANDN U1888 ( .A(n1654), .B(n57095), .Z(n1655) );
  NAND U1889 ( .A(n51555), .B(n1655), .Z(n1656) );
  NAND U1890 ( .A(n57096), .B(n1656), .Z(n1657) );
  NAND U1891 ( .A(n57097), .B(n1657), .Z(n57098) );
  NAND U1892 ( .A(n57141), .B(n57140), .Z(n1658) );
  AND U1893 ( .A(n57144), .B(n1658), .Z(n1659) );
  OR U1894 ( .A(n57145), .B(n1659), .Z(n1660) );
  NAND U1895 ( .A(n57146), .B(n1660), .Z(n1661) );
  NANDN U1896 ( .A(n57147), .B(n1661), .Z(n1662) );
  AND U1897 ( .A(n51542), .B(n51543), .Z(n1663) );
  NAND U1898 ( .A(n1662), .B(n1663), .Z(n1664) );
  NANDN U1899 ( .A(n57148), .B(n1664), .Z(n1665) );
  AND U1900 ( .A(n57150), .B(n57149), .Z(n1666) );
  NAND U1901 ( .A(n1665), .B(n1666), .Z(n1667) );
  NANDN U1902 ( .A(n57151), .B(n1667), .Z(n1668) );
  AND U1903 ( .A(n57153), .B(n57152), .Z(n1669) );
  NAND U1904 ( .A(n1668), .B(n1669), .Z(n1670) );
  NAND U1905 ( .A(n57154), .B(n1670), .Z(n1671) );
  AND U1906 ( .A(n57155), .B(n1671), .Z(n57157) );
  NAND U1907 ( .A(n57184), .B(n57183), .Z(n1672) );
  NANDN U1908 ( .A(n57186), .B(n1672), .Z(n1673) );
  AND U1909 ( .A(n57187), .B(n1673), .Z(n1674) );
  AND U1910 ( .A(n57190), .B(n57189), .Z(n1675) );
  OR U1911 ( .A(n1674), .B(n57188), .Z(n1676) );
  AND U1912 ( .A(n1675), .B(n1676), .Z(n1677) );
  OR U1913 ( .A(n1677), .B(n57191), .Z(n1678) );
  NAND U1914 ( .A(n57192), .B(n1678), .Z(n1679) );
  ANDN U1915 ( .B(n1679), .A(n57193), .Z(n1680) );
  NANDN U1916 ( .A(n1680), .B(n57194), .Z(n1681) );
  NANDN U1917 ( .A(n57195), .B(n1681), .Z(n1682) );
  NAND U1918 ( .A(n57196), .B(n1682), .Z(n1683) );
  NAND U1919 ( .A(n57197), .B(n1683), .Z(n1684) );
  NANDN U1920 ( .A(n57198), .B(n1684), .Z(n1685) );
  AND U1921 ( .A(n57199), .B(n1685), .Z(n1686) );
  NANDN U1922 ( .A(n1686), .B(n57200), .Z(n1687) );
  NAND U1923 ( .A(n57201), .B(n1687), .Z(n1688) );
  NANDN U1924 ( .A(n57202), .B(n1688), .Z(n57203) );
  OR U1925 ( .A(n57226), .B(n57227), .Z(n1689) );
  ANDN U1926 ( .B(n1689), .A(n51527), .Z(n1690) );
  ANDN U1927 ( .B(n57229), .A(n1690), .Z(n1691) );
  NAND U1928 ( .A(n57228), .B(n1691), .Z(n1692) );
  NAND U1929 ( .A(n57230), .B(n1692), .Z(n1693) );
  AND U1930 ( .A(n51526), .B(n51525), .Z(n1694) );
  NAND U1931 ( .A(n1693), .B(n1694), .Z(n1695) );
  NANDN U1932 ( .A(n57231), .B(n1695), .Z(n1696) );
  ANDN U1933 ( .B(n57232), .A(n57233), .Z(n1697) );
  NAND U1934 ( .A(n1696), .B(n1697), .Z(n1698) );
  NANDN U1935 ( .A(n57234), .B(n1698), .Z(n1699) );
  ANDN U1936 ( .B(n57235), .A(n57236), .Z(n1700) );
  NAND U1937 ( .A(n1699), .B(n1700), .Z(n1701) );
  NANDN U1938 ( .A(n51524), .B(n1701), .Z(n57237) );
  ANDN U1939 ( .B(n57269), .A(n57270), .Z(n1702) );
  NANDN U1940 ( .A(n57268), .B(n57267), .Z(n1703) );
  AND U1941 ( .A(n1702), .B(n1703), .Z(n1704) );
  ANDN U1942 ( .B(n57273), .A(n57272), .Z(n1705) );
  OR U1943 ( .A(n57271), .B(n1704), .Z(n1706) );
  AND U1944 ( .A(n1705), .B(n1706), .Z(n1707) );
  AND U1945 ( .A(n51518), .B(n51517), .Z(n1708) );
  OR U1946 ( .A(n57274), .B(n1707), .Z(n1709) );
  AND U1947 ( .A(n1708), .B(n1709), .Z(n1710) );
  AND U1948 ( .A(n51516), .B(n51515), .Z(n1711) );
  NANDN U1949 ( .A(n1710), .B(n57275), .Z(n1712) );
  AND U1950 ( .A(n1711), .B(n1712), .Z(n1713) );
  AND U1951 ( .A(n57277), .B(n57278), .Z(n1714) );
  NANDN U1952 ( .A(n1713), .B(n57276), .Z(n1715) );
  AND U1953 ( .A(n1714), .B(n1715), .Z(n1716) );
  OR U1954 ( .A(n57279), .B(n1716), .Z(n1717) );
  ANDN U1955 ( .B(n1717), .A(n57280), .Z(n57283) );
  ANDN U1956 ( .B(n51511), .A(n51512), .Z(n57297) );
  NANDN U1957 ( .A(n57332), .B(n57331), .Z(n1718) );
  NANDN U1958 ( .A(n51508), .B(n1718), .Z(n1719) );
  AND U1959 ( .A(n57333), .B(n1719), .Z(n1720) );
  ANDN U1960 ( .B(n57336), .A(n57335), .Z(n1721) );
  NANDN U1961 ( .A(n1720), .B(n57334), .Z(n1722) );
  AND U1962 ( .A(n1721), .B(n1722), .Z(n1723) );
  NANDN U1963 ( .A(n1723), .B(n51507), .Z(n1724) );
  ANDN U1964 ( .B(n1724), .A(n57337), .Z(n1725) );
  NAND U1965 ( .A(n1725), .B(n57338), .Z(n1726) );
  NAND U1966 ( .A(n57339), .B(n1726), .Z(n1727) );
  NAND U1967 ( .A(n57340), .B(n1727), .Z(n1728) );
  NANDN U1968 ( .A(n1728), .B(n57341), .Z(n1729) );
  NANDN U1969 ( .A(n57342), .B(n1729), .Z(n1730) );
  NAND U1970 ( .A(n57343), .B(n1730), .Z(n1731) );
  NAND U1971 ( .A(n57344), .B(n1731), .Z(n1732) );
  AND U1972 ( .A(n57346), .B(n1732), .Z(n1733) );
  NANDN U1973 ( .A(n57345), .B(n1733), .Z(n57347) );
  AND U1974 ( .A(n57379), .B(n51499), .Z(n1734) );
  AND U1975 ( .A(n57381), .B(n57382), .Z(n1735) );
  OR U1976 ( .A(n57380), .B(n1734), .Z(n1736) );
  AND U1977 ( .A(n1735), .B(n1736), .Z(n1737) );
  OR U1978 ( .A(n57383), .B(n1737), .Z(n1738) );
  NAND U1979 ( .A(n57384), .B(n1738), .Z(n1739) );
  NANDN U1980 ( .A(n57385), .B(n1739), .Z(n1740) );
  AND U1981 ( .A(n51498), .B(n51497), .Z(n1741) );
  NAND U1982 ( .A(n1740), .B(n1741), .Z(n1742) );
  NANDN U1983 ( .A(n57386), .B(n1742), .Z(n1743) );
  ANDN U1984 ( .B(n57387), .A(n57388), .Z(n1744) );
  NAND U1985 ( .A(n1743), .B(n1744), .Z(n1745) );
  NANDN U1986 ( .A(n57389), .B(n1745), .Z(n57391) );
  ANDN U1987 ( .B(n57423), .A(n57424), .Z(n1746) );
  NANDN U1988 ( .A(n57422), .B(n57421), .Z(n1747) );
  AND U1989 ( .A(n1746), .B(n1747), .Z(n1748) );
  ANDN U1990 ( .B(n51491), .A(n51492), .Z(n1749) );
  NANDN U1991 ( .A(n1748), .B(n57425), .Z(n1750) );
  AND U1992 ( .A(n1749), .B(n1750), .Z(n1751) );
  ANDN U1993 ( .B(n57427), .A(n57428), .Z(n1752) );
  NANDN U1994 ( .A(n1751), .B(n57426), .Z(n1753) );
  AND U1995 ( .A(n1752), .B(n1753), .Z(n1754) );
  ANDN U1996 ( .B(n57430), .A(n57429), .Z(n1755) );
  NANDN U1997 ( .A(n1754), .B(n51490), .Z(n1756) );
  AND U1998 ( .A(n1755), .B(n1756), .Z(n1757) );
  AND U1999 ( .A(n57433), .B(n57432), .Z(n1758) );
  OR U2000 ( .A(n57431), .B(n1757), .Z(n1759) );
  AND U2001 ( .A(n1758), .B(n1759), .Z(n57436) );
  NAND U2002 ( .A(n57465), .B(n57466), .Z(n1760) );
  AND U2003 ( .A(n57469), .B(n1760), .Z(n1761) );
  NANDN U2004 ( .A(n57468), .B(n1761), .Z(n1762) );
  NAND U2005 ( .A(n57470), .B(n1762), .Z(n1763) );
  NANDN U2006 ( .A(n57471), .B(n1763), .Z(n1764) );
  AND U2007 ( .A(n57472), .B(n1764), .Z(n1765) );
  OR U2008 ( .A(n57473), .B(n1765), .Z(n1766) );
  AND U2009 ( .A(n57474), .B(n1766), .Z(n1767) );
  OR U2010 ( .A(n57475), .B(n1767), .Z(n1768) );
  NAND U2011 ( .A(n57476), .B(n1768), .Z(n1769) );
  NANDN U2012 ( .A(n57477), .B(n1769), .Z(n1770) );
  NAND U2013 ( .A(n57478), .B(n1770), .Z(n1771) );
  AND U2014 ( .A(n51480), .B(n1771), .Z(n1772) );
  NANDN U2015 ( .A(n51481), .B(n1772), .Z(n1773) );
  NAND U2016 ( .A(n57479), .B(n1773), .Z(n1774) );
  AND U2017 ( .A(n57480), .B(n1774), .Z(n1775) );
  NANDN U2018 ( .A(n57481), .B(n1775), .Z(n57482) );
  NANDN U2019 ( .A(n57508), .B(n57507), .Z(n1776) );
  ANDN U2020 ( .B(n1776), .A(n57509), .Z(n1777) );
  ANDN U2021 ( .B(n57510), .A(n1777), .Z(n1778) );
  NAND U2022 ( .A(n57511), .B(n1778), .Z(n1779) );
  NANDN U2023 ( .A(n57512), .B(n1779), .Z(n1780) );
  AND U2024 ( .A(n57513), .B(n57514), .Z(n1781) );
  NAND U2025 ( .A(n1780), .B(n1781), .Z(n1782) );
  NANDN U2026 ( .A(n57515), .B(n1782), .Z(n1783) );
  NAND U2027 ( .A(n57516), .B(n1783), .Z(n1784) );
  NANDN U2028 ( .A(n57517), .B(n1784), .Z(n1785) );
  AND U2029 ( .A(n57518), .B(n1785), .Z(n1786) );
  AND U2030 ( .A(n57521), .B(n57520), .Z(n1787) );
  OR U2031 ( .A(n57519), .B(n1786), .Z(n1788) );
  AND U2032 ( .A(n1787), .B(n1788), .Z(n1789) );
  AND U2033 ( .A(n51468), .B(n51469), .Z(n1790) );
  NANDN U2034 ( .A(n1789), .B(n57522), .Z(n1791) );
  AND U2035 ( .A(n1790), .B(n1791), .Z(n57523) );
  NAND U2036 ( .A(n57552), .B(n57551), .Z(n1792) );
  AND U2037 ( .A(n57554), .B(n1792), .Z(n1793) );
  ANDN U2038 ( .B(n51460), .A(n1793), .Z(n1794) );
  NAND U2039 ( .A(n51461), .B(n1794), .Z(n1795) );
  NANDN U2040 ( .A(n57555), .B(n1795), .Z(n1796) );
  AND U2041 ( .A(n57556), .B(n57557), .Z(n1797) );
  NAND U2042 ( .A(n1796), .B(n1797), .Z(n1798) );
  NAND U2043 ( .A(n51459), .B(n1798), .Z(n1799) );
  ANDN U2044 ( .B(n57558), .A(n57559), .Z(n1800) );
  NAND U2045 ( .A(n1799), .B(n1800), .Z(n1801) );
  NANDN U2046 ( .A(n57560), .B(n1801), .Z(n1802) );
  ANDN U2047 ( .B(n57562), .A(n57561), .Z(n1803) );
  NAND U2048 ( .A(n1802), .B(n1803), .Z(n1804) );
  NAND U2049 ( .A(n57563), .B(n1804), .Z(n57564) );
  NAND U2050 ( .A(n57595), .B(n57594), .Z(n1805) );
  AND U2051 ( .A(n57596), .B(n1805), .Z(n1806) );
  NOR U2052 ( .A(n57597), .B(n1806), .Z(n1807) );
  NAND U2053 ( .A(n57598), .B(n1807), .Z(n1808) );
  NAND U2054 ( .A(n57599), .B(n1808), .Z(n1809) );
  NAND U2055 ( .A(n57600), .B(n1809), .Z(n1810) );
  NAND U2056 ( .A(n57601), .B(n1810), .Z(n1811) );
  ANDN U2057 ( .B(n1811), .A(n57602), .Z(n1812) );
  ANDN U2058 ( .B(n57605), .A(n57606), .Z(n1813) );
  NAND U2059 ( .A(n1812), .B(n57603), .Z(n1814) );
  NAND U2060 ( .A(n57604), .B(n1814), .Z(n1815) );
  AND U2061 ( .A(n1813), .B(n1815), .Z(n1816) );
  ANDN U2062 ( .B(n57608), .A(n57609), .Z(n1817) );
  OR U2063 ( .A(n57607), .B(n1816), .Z(n1818) );
  AND U2064 ( .A(n1817), .B(n1818), .Z(n1819) );
  ANDN U2065 ( .B(n57612), .A(n57611), .Z(n1820) );
  OR U2066 ( .A(n57610), .B(n1819), .Z(n1821) );
  AND U2067 ( .A(n1820), .B(n1821), .Z(n57614) );
  NANDN U2068 ( .A(n57645), .B(n57644), .Z(n1822) );
  NAND U2069 ( .A(n57647), .B(n1822), .Z(n1823) );
  NAND U2070 ( .A(n57648), .B(n1823), .Z(n1824) );
  NANDN U2071 ( .A(n51436), .B(n1824), .Z(n1825) );
  NAND U2072 ( .A(n51435), .B(n1825), .Z(n1826) );
  ANDN U2073 ( .B(n1826), .A(n57649), .Z(n1827) );
  ANDN U2074 ( .B(n57651), .A(n1827), .Z(n1828) );
  NAND U2075 ( .A(n57650), .B(n1828), .Z(n1829) );
  ANDN U2076 ( .B(n1829), .A(n57652), .Z(n1830) );
  NANDN U2077 ( .A(n1830), .B(n57653), .Z(n1831) );
  NANDN U2078 ( .A(n51434), .B(n1831), .Z(n1832) );
  NAND U2079 ( .A(n51433), .B(n1832), .Z(n57656) );
  ANDN U2080 ( .B(n57685), .A(n57686), .Z(n1833) );
  NAND U2081 ( .A(n57684), .B(n1833), .Z(n1834) );
  ANDN U2082 ( .B(n1834), .A(n57687), .Z(n1835) );
  NOR U2083 ( .A(n51424), .B(n1835), .Z(n1836) );
  NAND U2084 ( .A(n51425), .B(n1836), .Z(n1837) );
  ANDN U2085 ( .B(n1837), .A(n51423), .Z(n1838) );
  ANDN U2086 ( .B(n57688), .A(n1838), .Z(n1839) );
  NAND U2087 ( .A(n57689), .B(n1839), .Z(n1840) );
  ANDN U2088 ( .B(n1840), .A(n57690), .Z(n1841) );
  NANDN U2089 ( .A(n1841), .B(n57691), .Z(n1842) );
  ANDN U2090 ( .B(n1842), .A(n57692), .Z(n1843) );
  ANDN U2091 ( .B(n51422), .A(n1843), .Z(n1844) );
  NAND U2092 ( .A(n51421), .B(n1844), .Z(n1845) );
  NANDN U2093 ( .A(n57693), .B(n1845), .Z(n1846) );
  NAND U2094 ( .A(n57694), .B(n1846), .Z(n1847) );
  NAND U2095 ( .A(n51420), .B(n1847), .Z(n1848) );
  AND U2096 ( .A(n57695), .B(n1848), .Z(n57697) );
  NOR U2097 ( .A(n57726), .B(n57727), .Z(n1849) );
  NAND U2098 ( .A(n57724), .B(n57723), .Z(n1850) );
  AND U2099 ( .A(n1849), .B(n1850), .Z(n1851) );
  OR U2100 ( .A(n57728), .B(n1851), .Z(n1852) );
  NAND U2101 ( .A(n57729), .B(n1852), .Z(n1853) );
  NANDN U2102 ( .A(n51411), .B(n1853), .Z(n1854) );
  NAND U2103 ( .A(n51410), .B(n1854), .Z(n1855) );
  NANDN U2104 ( .A(n57730), .B(n1855), .Z(n1856) );
  AND U2105 ( .A(n57731), .B(n1856), .Z(n1857) );
  NANDN U2106 ( .A(n1857), .B(n57732), .Z(n1858) );
  NAND U2107 ( .A(n57733), .B(n1858), .Z(n1859) );
  NANDN U2108 ( .A(n51409), .B(n1859), .Z(n1860) );
  AND U2109 ( .A(n57734), .B(n1860), .Z(n57735) );
  AND U2110 ( .A(n57770), .B(n57769), .Z(n57771) );
  ANDN U2111 ( .B(n57803), .A(n57802), .Z(n1861) );
  NAND U2112 ( .A(n57804), .B(n1861), .Z(n1862) );
  NAND U2113 ( .A(n57805), .B(n1862), .Z(n1863) );
  ANDN U2114 ( .B(n57806), .A(n57807), .Z(n1864) );
  NAND U2115 ( .A(n1863), .B(n1864), .Z(n1865) );
  NAND U2116 ( .A(n57808), .B(n1865), .Z(n1866) );
  ANDN U2117 ( .B(n51390), .A(n51389), .Z(n1867) );
  NAND U2118 ( .A(n1866), .B(n1867), .Z(n1868) );
  NANDN U2119 ( .A(n57809), .B(n1868), .Z(n1869) );
  ANDN U2120 ( .B(n57810), .A(n57811), .Z(n1870) );
  NAND U2121 ( .A(n1869), .B(n1870), .Z(n1871) );
  NANDN U2122 ( .A(n57812), .B(n1871), .Z(n1872) );
  ANDN U2123 ( .B(n1872), .A(n57813), .Z(n1873) );
  NAND U2124 ( .A(n57814), .B(n1873), .Z(n57815) );
  NAND U2125 ( .A(n57864), .B(n57863), .Z(n1874) );
  NAND U2126 ( .A(n57867), .B(n1874), .Z(n1875) );
  NANDN U2127 ( .A(n57868), .B(n1875), .Z(n1876) );
  AND U2128 ( .A(n57869), .B(n57870), .Z(n1877) );
  NAND U2129 ( .A(n1876), .B(n1877), .Z(n1878) );
  NANDN U2130 ( .A(n57871), .B(n1878), .Z(n1879) );
  ANDN U2131 ( .B(n57872), .A(n57873), .Z(n1880) );
  NAND U2132 ( .A(n1879), .B(n1880), .Z(n1881) );
  NANDN U2133 ( .A(n57874), .B(n1881), .Z(n1882) );
  ANDN U2134 ( .B(n51376), .A(n51375), .Z(n1883) );
  NAND U2135 ( .A(n1882), .B(n1883), .Z(n1884) );
  NAND U2136 ( .A(n57875), .B(n1884), .Z(n1885) );
  ANDN U2137 ( .B(n57877), .A(n57876), .Z(n1886) );
  NAND U2138 ( .A(n1885), .B(n1886), .Z(n1887) );
  NANDN U2139 ( .A(n57878), .B(n1887), .Z(n1888) );
  AND U2140 ( .A(n57879), .B(n1888), .Z(n1889) );
  AND U2141 ( .A(n51373), .B(n51374), .Z(n1890) );
  OR U2142 ( .A(n1889), .B(n57880), .Z(n1891) );
  AND U2143 ( .A(n1890), .B(n1891), .Z(n57881) );
  NAND U2144 ( .A(n57905), .B(n57906), .Z(n1892) );
  ANDN U2145 ( .B(n1892), .A(n57907), .Z(n1893) );
  ANDN U2146 ( .B(n57908), .A(n1893), .Z(n1894) );
  NAND U2147 ( .A(n57909), .B(n1894), .Z(n1895) );
  AND U2148 ( .A(n51365), .B(n1895), .Z(n1896) );
  NOR U2149 ( .A(n57911), .B(n1896), .Z(n1897) );
  NAND U2150 ( .A(n57910), .B(n1897), .Z(n1898) );
  AND U2151 ( .A(n57912), .B(n1898), .Z(n1899) );
  NOR U2152 ( .A(n57913), .B(n57914), .Z(n1900) );
  NANDN U2153 ( .A(n1899), .B(n1900), .Z(n1901) );
  ANDN U2154 ( .B(n1901), .A(n57915), .Z(n1902) );
  NANDN U2155 ( .A(n1902), .B(n57916), .Z(n1903) );
  ANDN U2156 ( .B(n1903), .A(n57917), .Z(n57921) );
  NAND U2157 ( .A(n57940), .B(n57941), .Z(n1904) );
  ANDN U2158 ( .B(n1904), .A(n57943), .Z(n1905) );
  OR U2159 ( .A(n57946), .B(n57945), .Z(n1906) );
  NAND U2160 ( .A(n1905), .B(n1906), .Z(n1907) );
  NANDN U2161 ( .A(n57947), .B(n1907), .Z(n1908) );
  AND U2162 ( .A(n57949), .B(n57948), .Z(n1909) );
  NAND U2163 ( .A(n1908), .B(n1909), .Z(n1910) );
  NAND U2164 ( .A(n57950), .B(n1910), .Z(n1911) );
  AND U2165 ( .A(n51354), .B(n51355), .Z(n1912) );
  NAND U2166 ( .A(n1911), .B(n1912), .Z(n1913) );
  NANDN U2167 ( .A(n57951), .B(n1913), .Z(n1914) );
  ANDN U2168 ( .B(n57952), .A(n57953), .Z(n1915) );
  NAND U2169 ( .A(n1914), .B(n1915), .Z(n1916) );
  NAND U2170 ( .A(n51353), .B(n1916), .Z(n1917) );
  ANDN U2171 ( .B(n1917), .A(n57954), .Z(n57956) );
  NAND U2172 ( .A(n57981), .B(n57982), .Z(n1918) );
  NAND U2173 ( .A(n57983), .B(n1918), .Z(n1919) );
  AND U2174 ( .A(n51347), .B(n1919), .Z(n1920) );
  NAND U2175 ( .A(n1920), .B(n51346), .Z(n1921) );
  NAND U2176 ( .A(n57984), .B(n1921), .Z(n1922) );
  AND U2177 ( .A(n57985), .B(n1922), .Z(n1923) );
  NANDN U2178 ( .A(n57986), .B(n1923), .Z(n1924) );
  ANDN U2179 ( .B(n57988), .A(n57989), .Z(n1925) );
  NANDN U2180 ( .A(n57987), .B(n1924), .Z(n1926) );
  NAND U2181 ( .A(n1925), .B(n1926), .Z(n1927) );
  ANDN U2182 ( .B(n57992), .A(n57991), .Z(n1928) );
  NANDN U2183 ( .A(n57990), .B(n1927), .Z(n1929) );
  NAND U2184 ( .A(n1928), .B(n1929), .Z(n1930) );
  NAND U2185 ( .A(n57993), .B(n1930), .Z(n1931) );
  AND U2186 ( .A(n51345), .B(n1931), .Z(n1932) );
  NAND U2187 ( .A(n1932), .B(n51344), .Z(n57994) );
  AND U2188 ( .A(n58046), .B(n58045), .Z(n58047) );
  AND U2189 ( .A(n58072), .B(n58073), .Z(n1933) );
  NAND U2190 ( .A(n58075), .B(n1933), .Z(n1934) );
  NANDN U2191 ( .A(n58076), .B(n1934), .Z(n1935) );
  AND U2192 ( .A(n58078), .B(n58077), .Z(n1936) );
  NAND U2193 ( .A(n1935), .B(n1936), .Z(n1937) );
  NAND U2194 ( .A(n58079), .B(n1937), .Z(n1938) );
  AND U2195 ( .A(n51327), .B(n51326), .Z(n1939) );
  NAND U2196 ( .A(n1938), .B(n1939), .Z(n1940) );
  NAND U2197 ( .A(n58080), .B(n1940), .Z(n1941) );
  AND U2198 ( .A(n58081), .B(n58082), .Z(n1942) );
  NAND U2199 ( .A(n1941), .B(n1942), .Z(n1943) );
  NANDN U2200 ( .A(n58083), .B(n1943), .Z(n1944) );
  AND U2201 ( .A(n58085), .B(n58084), .Z(n1945) );
  NAND U2202 ( .A(n1944), .B(n1945), .Z(n1946) );
  NANDN U2203 ( .A(n58086), .B(n1946), .Z(n1947) );
  AND U2204 ( .A(n58088), .B(n58087), .Z(n1948) );
  NAND U2205 ( .A(n1947), .B(n1948), .Z(n1949) );
  NAND U2206 ( .A(n58089), .B(n1949), .Z(n58090) );
  AND U2207 ( .A(n58135), .B(n58134), .Z(n58136) );
  NAND U2208 ( .A(n58161), .B(n58160), .Z(n1950) );
  NANDN U2209 ( .A(n58162), .B(n1950), .Z(n1951) );
  NAND U2210 ( .A(n58163), .B(n1951), .Z(n1952) );
  NANDN U2211 ( .A(n1952), .B(n58164), .Z(n1953) );
  ANDN U2212 ( .B(n1953), .A(n58165), .Z(n1954) );
  NANDN U2213 ( .A(n1954), .B(n58166), .Z(n1955) );
  NANDN U2214 ( .A(n58167), .B(n1955), .Z(n1956) );
  NAND U2215 ( .A(n58168), .B(n1956), .Z(n1957) );
  AND U2216 ( .A(n58170), .B(n58171), .Z(n1958) );
  NANDN U2217 ( .A(n58169), .B(n1957), .Z(n1959) );
  NAND U2218 ( .A(n1958), .B(n1959), .Z(n1960) );
  AND U2219 ( .A(n51302), .B(n51303), .Z(n1961) );
  NANDN U2220 ( .A(n58172), .B(n1960), .Z(n1962) );
  NAND U2221 ( .A(n1961), .B(n1962), .Z(n1963) );
  ANDN U2222 ( .B(n58175), .A(n58174), .Z(n1964) );
  NANDN U2223 ( .A(n58173), .B(n1963), .Z(n1965) );
  NAND U2224 ( .A(n1964), .B(n1965), .Z(n58176) );
  AND U2225 ( .A(n58199), .B(n58198), .Z(n1966) );
  NAND U2226 ( .A(n58200), .B(n1966), .Z(n1967) );
  NAND U2227 ( .A(n58201), .B(n1967), .Z(n1968) );
  ANDN U2228 ( .B(n58203), .A(n58202), .Z(n1969) );
  NAND U2229 ( .A(n1968), .B(n1969), .Z(n1970) );
  NANDN U2230 ( .A(n58204), .B(n1970), .Z(n1971) );
  AND U2231 ( .A(n51291), .B(n51290), .Z(n1972) );
  NAND U2232 ( .A(n1971), .B(n1972), .Z(n1973) );
  NANDN U2233 ( .A(n58205), .B(n1973), .Z(n1974) );
  AND U2234 ( .A(n58207), .B(n58206), .Z(n1975) );
  NAND U2235 ( .A(n1974), .B(n1975), .Z(n1976) );
  NANDN U2236 ( .A(n58208), .B(n1976), .Z(n1977) );
  AND U2237 ( .A(n51289), .B(n58209), .Z(n1978) );
  NAND U2238 ( .A(n1977), .B(n1978), .Z(n1979) );
  NAND U2239 ( .A(n58210), .B(n1979), .Z(n1980) );
  AND U2240 ( .A(n58211), .B(n1980), .Z(n58213) );
  NAND U2241 ( .A(n58236), .B(n58235), .Z(n1981) );
  NANDN U2242 ( .A(n58238), .B(n1981), .Z(n1982) );
  ANDN U2243 ( .B(n1982), .A(n51279), .Z(n1983) );
  NANDN U2244 ( .A(n1983), .B(n58239), .Z(n1984) );
  NANDN U2245 ( .A(n58240), .B(n1984), .Z(n1985) );
  NAND U2246 ( .A(n58241), .B(n1985), .Z(n1986) );
  NANDN U2247 ( .A(n51278), .B(n1986), .Z(n1987) );
  NAND U2248 ( .A(n51277), .B(n1987), .Z(n1988) );
  AND U2249 ( .A(n58242), .B(n1988), .Z(n1989) );
  NAND U2250 ( .A(n1989), .B(n58243), .Z(n1990) );
  NANDN U2251 ( .A(n58244), .B(n1990), .Z(n1991) );
  AND U2252 ( .A(n58245), .B(n1991), .Z(n1992) );
  OR U2253 ( .A(n1992), .B(n58246), .Z(n1993) );
  NAND U2254 ( .A(n58247), .B(n1993), .Z(n1994) );
  NANDN U2255 ( .A(n58248), .B(n1994), .Z(n58249) );
  ANDN U2256 ( .B(n51265), .A(n51264), .Z(n1995) );
  NANDN U2257 ( .A(n58320), .B(n58319), .Z(n1996) );
  AND U2258 ( .A(n1995), .B(n1996), .Z(n1997) );
  AND U2259 ( .A(n58323), .B(n58322), .Z(n1998) );
  NANDN U2260 ( .A(n1997), .B(n58321), .Z(n1999) );
  AND U2261 ( .A(n1998), .B(n1999), .Z(n2000) );
  OR U2262 ( .A(n58324), .B(n2000), .Z(n2001) );
  NAND U2263 ( .A(n58325), .B(n2001), .Z(n2002) );
  NAND U2264 ( .A(n58326), .B(n2002), .Z(n2003) );
  ANDN U2265 ( .B(n51262), .A(n51261), .Z(n2004) );
  NAND U2266 ( .A(n2003), .B(n2004), .Z(n2005) );
  NAND U2267 ( .A(n58327), .B(n2005), .Z(n2006) );
  AND U2268 ( .A(n58328), .B(n58329), .Z(n2007) );
  NAND U2269 ( .A(n2006), .B(n2007), .Z(n2008) );
  NAND U2270 ( .A(n51260), .B(n2008), .Z(n2009) );
  AND U2271 ( .A(n58330), .B(n58331), .Z(n2010) );
  NAND U2272 ( .A(n2009), .B(n2010), .Z(n2011) );
  NANDN U2273 ( .A(n58332), .B(n2011), .Z(n2012) );
  AND U2274 ( .A(n58333), .B(n2012), .Z(n58335) );
  OR U2275 ( .A(n58365), .B(n58366), .Z(n2013) );
  NAND U2276 ( .A(n58367), .B(n2013), .Z(n2014) );
  ANDN U2277 ( .B(n2014), .A(n58368), .Z(n2015) );
  NANDN U2278 ( .A(n2015), .B(n58369), .Z(n2016) );
  NANDN U2279 ( .A(n58370), .B(n2016), .Z(n2017) );
  NAND U2280 ( .A(n58371), .B(n2017), .Z(n2018) );
  NANDN U2281 ( .A(n2018), .B(n58372), .Z(n2019) );
  NANDN U2282 ( .A(n51252), .B(n2019), .Z(n2020) );
  NAND U2283 ( .A(n58373), .B(n2020), .Z(n2021) );
  NANDN U2284 ( .A(n2021), .B(n58374), .Z(n2022) );
  NANDN U2285 ( .A(n58375), .B(n2022), .Z(n2023) );
  NAND U2286 ( .A(n58376), .B(n2023), .Z(n2024) );
  NAND U2287 ( .A(n51251), .B(n2024), .Z(n2025) );
  AND U2288 ( .A(n58378), .B(n2025), .Z(n2026) );
  NAND U2289 ( .A(n2026), .B(n58377), .Z(n2027) );
  NANDN U2290 ( .A(n58379), .B(n2027), .Z(n58380) );
  AND U2291 ( .A(n51239), .B(n51240), .Z(n2028) );
  AND U2292 ( .A(n58404), .B(n58405), .Z(n2029) );
  NAND U2293 ( .A(n58403), .B(n2029), .Z(n2030) );
  NANDN U2294 ( .A(n58406), .B(n2030), .Z(n2031) );
  AND U2295 ( .A(n51241), .B(n51242), .Z(n2032) );
  NAND U2296 ( .A(n2031), .B(n2032), .Z(n2033) );
  NANDN U2297 ( .A(n58407), .B(n2033), .Z(n2034) );
  AND U2298 ( .A(n58408), .B(n58409), .Z(n2035) );
  NAND U2299 ( .A(n2034), .B(n2035), .Z(n2036) );
  NANDN U2300 ( .A(n58410), .B(n2036), .Z(n2037) );
  AND U2301 ( .A(n58412), .B(n58411), .Z(n2038) );
  NAND U2302 ( .A(n2037), .B(n2038), .Z(n2039) );
  NAND U2303 ( .A(n58413), .B(n2039), .Z(n2040) );
  AND U2304 ( .A(n58414), .B(n58415), .Z(n2041) );
  NAND U2305 ( .A(n2040), .B(n2041), .Z(n2042) );
  NANDN U2306 ( .A(n58416), .B(n2042), .Z(n2043) );
  NAND U2307 ( .A(n2028), .B(n2043), .Z(n58419) );
  AND U2308 ( .A(n58449), .B(n58448), .Z(n2044) );
  NAND U2309 ( .A(n58450), .B(n2044), .Z(n2045) );
  NANDN U2310 ( .A(n58451), .B(n2045), .Z(n2046) );
  AND U2311 ( .A(n58453), .B(n58452), .Z(n2047) );
  NAND U2312 ( .A(n2046), .B(n2047), .Z(n2048) );
  NAND U2313 ( .A(n58454), .B(n2048), .Z(n2049) );
  AND U2314 ( .A(n58456), .B(n58455), .Z(n2050) );
  NAND U2315 ( .A(n2049), .B(n2050), .Z(n2051) );
  NAND U2316 ( .A(n58457), .B(n2051), .Z(n2052) );
  AND U2317 ( .A(n51231), .B(n51232), .Z(n2053) );
  NAND U2318 ( .A(n2052), .B(n2053), .Z(n2054) );
  NANDN U2319 ( .A(n58458), .B(n2054), .Z(n2055) );
  AND U2320 ( .A(n58460), .B(n58459), .Z(n2056) );
  NAND U2321 ( .A(n2055), .B(n2056), .Z(n2057) );
  NANDN U2322 ( .A(n58461), .B(n2057), .Z(n2058) );
  AND U2323 ( .A(n58462), .B(n2058), .Z(n58463) );
  AND U2324 ( .A(n58526), .B(n58527), .Z(n2059) );
  OR U2325 ( .A(n58523), .B(n58524), .Z(n2060) );
  NAND U2326 ( .A(n2059), .B(n2060), .Z(n2061) );
  ANDN U2327 ( .B(n51213), .A(n51212), .Z(n2062) );
  NANDN U2328 ( .A(n58528), .B(n2061), .Z(n2063) );
  NAND U2329 ( .A(n2062), .B(n2063), .Z(n2064) );
  AND U2330 ( .A(n58530), .B(n58531), .Z(n2065) );
  NANDN U2331 ( .A(n58529), .B(n2064), .Z(n2066) );
  NAND U2332 ( .A(n2065), .B(n2066), .Z(n2067) );
  NAND U2333 ( .A(n51211), .B(n2067), .Z(n2068) );
  AND U2334 ( .A(n58533), .B(n2068), .Z(n2069) );
  NAND U2335 ( .A(n2069), .B(n58532), .Z(n2070) );
  NAND U2336 ( .A(n58534), .B(n2070), .Z(n2071) );
  AND U2337 ( .A(n58536), .B(n2071), .Z(n2072) );
  NAND U2338 ( .A(n2072), .B(n58535), .Z(n2073) );
  NANDN U2339 ( .A(n58537), .B(n2073), .Z(n58538) );
  NAND U2340 ( .A(n58564), .B(n58563), .Z(n2074) );
  AND U2341 ( .A(n58565), .B(n2074), .Z(n2075) );
  ANDN U2342 ( .B(n58567), .A(n2075), .Z(n2076) );
  NAND U2343 ( .A(n58566), .B(n2076), .Z(n2077) );
  NANDN U2344 ( .A(n58568), .B(n2077), .Z(n2078) );
  AND U2345 ( .A(n51200), .B(n51201), .Z(n2079) );
  NAND U2346 ( .A(n2078), .B(n2079), .Z(n2080) );
  NANDN U2347 ( .A(n58569), .B(n2080), .Z(n2081) );
  AND U2348 ( .A(n58570), .B(n58571), .Z(n2082) );
  NAND U2349 ( .A(n2081), .B(n2082), .Z(n2083) );
  NANDN U2350 ( .A(n58572), .B(n2083), .Z(n2084) );
  NAND U2351 ( .A(n58573), .B(n2084), .Z(n2085) );
  AND U2352 ( .A(n51199), .B(n51198), .Z(n2086) );
  NANDN U2353 ( .A(n58574), .B(n2085), .Z(n2087) );
  NAND U2354 ( .A(n2086), .B(n2087), .Z(n58577) );
  NAND U2355 ( .A(n58612), .B(n58611), .Z(n2088) );
  NANDN U2356 ( .A(n58613), .B(n2088), .Z(n2089) );
  AND U2357 ( .A(n58614), .B(n2089), .Z(n2090) );
  NANDN U2358 ( .A(n2090), .B(n58615), .Z(n2091) );
  NANDN U2359 ( .A(n58616), .B(n2091), .Z(n2092) );
  NAND U2360 ( .A(n58617), .B(n2092), .Z(n2093) );
  NANDN U2361 ( .A(n2093), .B(n58618), .Z(n2094) );
  ANDN U2362 ( .B(n2094), .A(n58619), .Z(n2095) );
  ANDN U2363 ( .B(n51192), .A(n2095), .Z(n2096) );
  NAND U2364 ( .A(n51191), .B(n2096), .Z(n2097) );
  ANDN U2365 ( .B(n2097), .A(n58620), .Z(n2098) );
  NANDN U2366 ( .A(n2098), .B(n58621), .Z(n2099) );
  NANDN U2367 ( .A(n58622), .B(n2099), .Z(n2100) );
  NAND U2368 ( .A(n58623), .B(n2100), .Z(n2101) );
  AND U2369 ( .A(n51189), .B(n51190), .Z(n2102) );
  NANDN U2370 ( .A(n58624), .B(n2101), .Z(n2103) );
  NAND U2371 ( .A(n2102), .B(n2103), .Z(n2104) );
  NANDN U2372 ( .A(n58625), .B(n2104), .Z(n58626) );
  AND U2373 ( .A(n58662), .B(n58663), .Z(n2105) );
  OR U2374 ( .A(n58660), .B(n58661), .Z(n2106) );
  AND U2375 ( .A(n2105), .B(n2106), .Z(n2107) );
  AND U2376 ( .A(n51181), .B(n51182), .Z(n2108) );
  OR U2377 ( .A(n58664), .B(n2107), .Z(n2109) );
  AND U2378 ( .A(n2108), .B(n2109), .Z(n2110) );
  AND U2379 ( .A(n51179), .B(n51180), .Z(n2111) );
  NANDN U2380 ( .A(n2110), .B(n58665), .Z(n2112) );
  AND U2381 ( .A(n2111), .B(n2112), .Z(n2113) );
  AND U2382 ( .A(n58667), .B(n58666), .Z(n2114) );
  OR U2383 ( .A(n51178), .B(n2113), .Z(n2115) );
  AND U2384 ( .A(n2114), .B(n2115), .Z(n2116) );
  AND U2385 ( .A(n58670), .B(n58669), .Z(n2117) );
  OR U2386 ( .A(n58668), .B(n2116), .Z(n2118) );
  AND U2387 ( .A(n2117), .B(n2118), .Z(n2119) );
  AND U2388 ( .A(n51177), .B(n51176), .Z(n2120) );
  OR U2389 ( .A(n2119), .B(n58671), .Z(n2121) );
  NAND U2390 ( .A(n2120), .B(n2121), .Z(n2122) );
  AND U2391 ( .A(n58672), .B(n2122), .Z(n58676) );
  AND U2392 ( .A(n58710), .B(n58709), .Z(n2123) );
  OR U2393 ( .A(n58707), .B(n58708), .Z(n2124) );
  NAND U2394 ( .A(n2123), .B(n2124), .Z(n2125) );
  AND U2395 ( .A(n51169), .B(n51168), .Z(n2126) );
  NANDN U2396 ( .A(n58711), .B(n2125), .Z(n2127) );
  NAND U2397 ( .A(n2126), .B(n2127), .Z(n2128) );
  NAND U2398 ( .A(n58712), .B(n2128), .Z(n2129) );
  AND U2399 ( .A(n58713), .B(n2129), .Z(n2130) );
  NAND U2400 ( .A(n2130), .B(n58714), .Z(n2131) );
  NAND U2401 ( .A(n51167), .B(n2131), .Z(n2132) );
  AND U2402 ( .A(n58716), .B(n2132), .Z(n2133) );
  NAND U2403 ( .A(n2133), .B(n58715), .Z(n2134) );
  AND U2404 ( .A(n58719), .B(n58718), .Z(n2135) );
  NANDN U2405 ( .A(n58717), .B(n2134), .Z(n2136) );
  NAND U2406 ( .A(n2135), .B(n2136), .Z(n2137) );
  NAND U2407 ( .A(n58720), .B(n2137), .Z(n2138) );
  NAND U2408 ( .A(n58721), .B(n2138), .Z(n2139) );
  AND U2409 ( .A(n58722), .B(n2139), .Z(n58726) );
  NAND U2410 ( .A(n58764), .B(n58765), .Z(n2140) );
  NAND U2411 ( .A(n58767), .B(n2140), .Z(n2141) );
  AND U2412 ( .A(n58770), .B(n2141), .Z(n2142) );
  NANDN U2413 ( .A(n58769), .B(n2142), .Z(n2143) );
  NAND U2414 ( .A(n51153), .B(n2143), .Z(n2144) );
  AND U2415 ( .A(n58771), .B(n2144), .Z(n2145) );
  NANDN U2416 ( .A(n58772), .B(n2145), .Z(n2146) );
  ANDN U2417 ( .B(n58775), .A(n58774), .Z(n2147) );
  NANDN U2418 ( .A(n58773), .B(n2146), .Z(n2148) );
  NAND U2419 ( .A(n2147), .B(n2148), .Z(n2149) );
  ANDN U2420 ( .B(n51152), .A(n51151), .Z(n2150) );
  NANDN U2421 ( .A(n58776), .B(n2149), .Z(n2151) );
  NAND U2422 ( .A(n2150), .B(n2151), .Z(n2152) );
  NAND U2423 ( .A(n58777), .B(n2152), .Z(n2153) );
  AND U2424 ( .A(n58778), .B(n2153), .Z(n2154) );
  NANDN U2425 ( .A(n58779), .B(n2154), .Z(n58780) );
  NAND U2426 ( .A(n58813), .B(n58814), .Z(n2155) );
  AND U2427 ( .A(n58817), .B(n2155), .Z(n2156) );
  ANDN U2428 ( .B(n58818), .A(n58819), .Z(n2157) );
  NANDN U2429 ( .A(n2156), .B(n51135), .Z(n2158) );
  AND U2430 ( .A(n2157), .B(n2158), .Z(n2159) );
  ANDN U2431 ( .B(n58822), .A(n58821), .Z(n2160) );
  OR U2432 ( .A(n58820), .B(n2159), .Z(n2161) );
  AND U2433 ( .A(n2160), .B(n2161), .Z(n2162) );
  AND U2434 ( .A(n51134), .B(n51133), .Z(n2163) );
  OR U2435 ( .A(n58823), .B(n2162), .Z(n2164) );
  AND U2436 ( .A(n2163), .B(n2164), .Z(n2165) );
  OR U2437 ( .A(n58824), .B(n2165), .Z(n2166) );
  NAND U2438 ( .A(n58825), .B(n2166), .Z(n2167) );
  NANDN U2439 ( .A(n58826), .B(n2167), .Z(n2168) );
  AND U2440 ( .A(n58828), .B(n58827), .Z(n2169) );
  NAND U2441 ( .A(n2168), .B(n2169), .Z(n2170) );
  NANDN U2442 ( .A(n58829), .B(n2170), .Z(n58830) );
  NAND U2443 ( .A(n58868), .B(n58867), .Z(n2171) );
  AND U2444 ( .A(n58871), .B(n2171), .Z(n2172) );
  AND U2445 ( .A(n51119), .B(n58873), .Z(n2173) );
  OR U2446 ( .A(n58872), .B(n2172), .Z(n2174) );
  AND U2447 ( .A(n2173), .B(n2174), .Z(n2175) );
  OR U2448 ( .A(n51118), .B(n2175), .Z(n2176) );
  NAND U2449 ( .A(n51117), .B(n2176), .Z(n2177) );
  NANDN U2450 ( .A(n58874), .B(n2177), .Z(n2178) );
  ANDN U2451 ( .B(n58875), .A(n58876), .Z(n2179) );
  NAND U2452 ( .A(n2178), .B(n2179), .Z(n2180) );
  NANDN U2453 ( .A(n58877), .B(n2180), .Z(n2181) );
  ANDN U2454 ( .B(n58879), .A(n58878), .Z(n2182) );
  NAND U2455 ( .A(n2181), .B(n2182), .Z(n2183) );
  NANDN U2456 ( .A(n58880), .B(n2183), .Z(n2184) );
  AND U2457 ( .A(n58881), .B(n2184), .Z(n58883) );
  ANDN U2458 ( .B(n58941), .A(n58940), .Z(n2185) );
  NAND U2459 ( .A(n58942), .B(n2185), .Z(n2186) );
  ANDN U2460 ( .B(n2186), .A(n58943), .Z(n2187) );
  ANDN U2461 ( .B(n58945), .A(n2187), .Z(n2188) );
  NAND U2462 ( .A(n58944), .B(n2188), .Z(n2189) );
  AND U2463 ( .A(n58946), .B(n2189), .Z(n2190) );
  NOR U2464 ( .A(n51100), .B(n2190), .Z(n2191) );
  NAND U2465 ( .A(n51101), .B(n2191), .Z(n2192) );
  AND U2466 ( .A(n58947), .B(n2192), .Z(n2193) );
  NOR U2467 ( .A(n58948), .B(n2193), .Z(n2194) );
  NAND U2468 ( .A(n58949), .B(n2194), .Z(n2195) );
  ANDN U2469 ( .B(n2195), .A(n58950), .Z(n2196) );
  NOR U2470 ( .A(n58951), .B(n2196), .Z(n2197) );
  NAND U2471 ( .A(n58952), .B(n2197), .Z(n2198) );
  ANDN U2472 ( .B(n2198), .A(n58953), .Z(n2199) );
  NANDN U2473 ( .A(n2199), .B(n58954), .Z(n2200) );
  NANDN U2474 ( .A(n58955), .B(n2200), .Z(n2201) );
  NAND U2475 ( .A(n58956), .B(n2201), .Z(n58957) );
  NAND U2476 ( .A(n58991), .B(n58990), .Z(n2202) );
  AND U2477 ( .A(n58992), .B(n2202), .Z(n2203) );
  NOR U2478 ( .A(n2203), .B(n51093), .Z(n2204) );
  NAND U2479 ( .A(n51094), .B(n2204), .Z(n2205) );
  NANDN U2480 ( .A(n58993), .B(n2205), .Z(n2206) );
  NAND U2481 ( .A(n58994), .B(n2206), .Z(n2207) );
  NANDN U2482 ( .A(n58995), .B(n2207), .Z(n2208) );
  AND U2483 ( .A(n58996), .B(n2208), .Z(n2209) );
  AND U2484 ( .A(n58997), .B(n2209), .Z(n2210) );
  ANDN U2485 ( .B(n51092), .A(n51091), .Z(n2211) );
  OR U2486 ( .A(n58998), .B(n2210), .Z(n2212) );
  AND U2487 ( .A(n2211), .B(n2212), .Z(n2213) );
  OR U2488 ( .A(n58999), .B(n2213), .Z(n2214) );
  NAND U2489 ( .A(n59000), .B(n2214), .Z(n2215) );
  NAND U2490 ( .A(n59001), .B(n2215), .Z(n2216) );
  AND U2491 ( .A(n59003), .B(n59002), .Z(n2217) );
  NAND U2492 ( .A(n2216), .B(n2217), .Z(n2218) );
  NANDN U2493 ( .A(n59004), .B(n2218), .Z(n59005) );
  NAND U2494 ( .A(n59042), .B(n59043), .Z(n2219) );
  NAND U2495 ( .A(n59046), .B(n2219), .Z(n2220) );
  NANDN U2496 ( .A(n59047), .B(n2220), .Z(n2221) );
  ANDN U2497 ( .B(n51074), .A(n59048), .Z(n2222) );
  NAND U2498 ( .A(n2221), .B(n2222), .Z(n2223) );
  NAND U2499 ( .A(n59049), .B(n2223), .Z(n2224) );
  ANDN U2500 ( .B(n59050), .A(n59051), .Z(n2225) );
  NAND U2501 ( .A(n2224), .B(n2225), .Z(n2226) );
  NANDN U2502 ( .A(n59052), .B(n2226), .Z(n2227) );
  ANDN U2503 ( .B(n51073), .A(n51072), .Z(n2228) );
  NAND U2504 ( .A(n2227), .B(n2228), .Z(n2229) );
  NANDN U2505 ( .A(n59053), .B(n2229), .Z(n2230) );
  AND U2506 ( .A(n59055), .B(n59054), .Z(n2231) );
  NAND U2507 ( .A(n2230), .B(n2231), .Z(n2232) );
  NANDN U2508 ( .A(n59056), .B(n2232), .Z(n2233) );
  AND U2509 ( .A(n59057), .B(n2233), .Z(n59059) );
  NAND U2510 ( .A(n59084), .B(n59083), .Z(n2234) );
  NAND U2511 ( .A(n59085), .B(n2234), .Z(n2235) );
  ANDN U2512 ( .B(n2235), .A(n51062), .Z(n2236) );
  AND U2513 ( .A(n59088), .B(n59087), .Z(n2237) );
  NANDN U2514 ( .A(n2236), .B(n59086), .Z(n2238) );
  AND U2515 ( .A(n2237), .B(n2238), .Z(n2239) );
  AND U2516 ( .A(n59091), .B(n59090), .Z(n2240) );
  NANDN U2517 ( .A(n2239), .B(n59089), .Z(n2241) );
  AND U2518 ( .A(n2240), .B(n2241), .Z(n2242) );
  OR U2519 ( .A(n59092), .B(n2242), .Z(n2243) );
  AND U2520 ( .A(n59093), .B(n2243), .Z(n2244) );
  OR U2521 ( .A(n59094), .B(n2244), .Z(n2245) );
  NAND U2522 ( .A(n59095), .B(n2245), .Z(n2246) );
  NANDN U2523 ( .A(n59096), .B(n2246), .Z(n2247) );
  AND U2524 ( .A(n59098), .B(n59097), .Z(n2248) );
  NAND U2525 ( .A(n2247), .B(n2248), .Z(n2249) );
  NAND U2526 ( .A(n59099), .B(n2249), .Z(n59100) );
  ANDN U2527 ( .B(n59175), .A(n59174), .Z(n2250) );
  NAND U2528 ( .A(n59171), .B(n59172), .Z(n2251) );
  AND U2529 ( .A(n2250), .B(n2251), .Z(n2252) );
  AND U2530 ( .A(n59177), .B(n59178), .Z(n2253) );
  OR U2531 ( .A(n59176), .B(n2252), .Z(n2254) );
  AND U2532 ( .A(n2253), .B(n2254), .Z(n2255) );
  AND U2533 ( .A(n59180), .B(n59181), .Z(n2256) );
  NANDN U2534 ( .A(n2255), .B(n59179), .Z(n2257) );
  AND U2535 ( .A(n2256), .B(n2257), .Z(n2258) );
  AND U2536 ( .A(n51051), .B(n51050), .Z(n2259) );
  NANDN U2537 ( .A(n2258), .B(n59182), .Z(n2260) );
  AND U2538 ( .A(n2259), .B(n2260), .Z(n2261) );
  AND U2539 ( .A(n59184), .B(n59185), .Z(n2262) );
  NANDN U2540 ( .A(n2261), .B(n59183), .Z(n2263) );
  AND U2541 ( .A(n2262), .B(n2263), .Z(n2264) );
  NANDN U2542 ( .A(n2264), .B(n59186), .Z(n2265) );
  AND U2543 ( .A(n59187), .B(n2265), .Z(n59189) );
  AND U2544 ( .A(n59220), .B(n59222), .Z(n2266) );
  NAND U2545 ( .A(n59221), .B(n2266), .Z(n2267) );
  AND U2546 ( .A(n59223), .B(n2267), .Z(n2268) );
  ANDN U2547 ( .B(n59225), .A(n2268), .Z(n2269) );
  NAND U2548 ( .A(n59224), .B(n2269), .Z(n2270) );
  AND U2549 ( .A(n59226), .B(n2270), .Z(n2271) );
  ANDN U2550 ( .B(n51042), .A(n2271), .Z(n2272) );
  NAND U2551 ( .A(n51041), .B(n2272), .Z(n2273) );
  AND U2552 ( .A(n59227), .B(n2273), .Z(n2274) );
  NANDN U2553 ( .A(n2274), .B(n59228), .Z(n2275) );
  NANDN U2554 ( .A(n59229), .B(n2275), .Z(n2276) );
  NAND U2555 ( .A(n59230), .B(n2276), .Z(n2277) );
  AND U2556 ( .A(n51039), .B(n51040), .Z(n2278) );
  NANDN U2557 ( .A(n59231), .B(n2277), .Z(n2279) );
  NAND U2558 ( .A(n2278), .B(n2279), .Z(n2280) );
  NAND U2559 ( .A(n59232), .B(n2280), .Z(n2281) );
  AND U2560 ( .A(n59234), .B(n2281), .Z(n2282) );
  NAND U2561 ( .A(n2282), .B(n59233), .Z(n59235) );
  AND U2562 ( .A(n59263), .B(n59264), .Z(n2283) );
  NAND U2563 ( .A(n59265), .B(n2283), .Z(n2284) );
  NANDN U2564 ( .A(n59266), .B(n2284), .Z(n2285) );
  NAND U2565 ( .A(n59267), .B(n2285), .Z(n2286) );
  NAND U2566 ( .A(n59268), .B(n2286), .Z(n2287) );
  AND U2567 ( .A(n59269), .B(n2287), .Z(n2288) );
  AND U2568 ( .A(n59271), .B(n59270), .Z(n2289) );
  NANDN U2569 ( .A(n2288), .B(n51031), .Z(n2290) );
  AND U2570 ( .A(n2289), .B(n2290), .Z(n2291) );
  ANDN U2571 ( .B(n51030), .A(n51029), .Z(n2292) );
  OR U2572 ( .A(n59272), .B(n2291), .Z(n2293) );
  AND U2573 ( .A(n2292), .B(n2293), .Z(n2294) );
  AND U2574 ( .A(n59275), .B(n59274), .Z(n2295) );
  NANDN U2575 ( .A(n2294), .B(n59273), .Z(n2296) );
  AND U2576 ( .A(n2295), .B(n2296), .Z(n2297) );
  OR U2577 ( .A(n59276), .B(n2297), .Z(n2298) );
  AND U2578 ( .A(n59277), .B(n2298), .Z(n59279) );
  NAND U2579 ( .A(n59308), .B(n59309), .Z(n2299) );
  AND U2580 ( .A(n59311), .B(n2299), .Z(n2300) );
  NAND U2581 ( .A(n2300), .B(n59310), .Z(n2301) );
  AND U2582 ( .A(n59313), .B(n59314), .Z(n2302) );
  NANDN U2583 ( .A(n59312), .B(n2301), .Z(n2303) );
  NAND U2584 ( .A(n2302), .B(n2303), .Z(n2304) );
  AND U2585 ( .A(n51021), .B(n51020), .Z(n2305) );
  NANDN U2586 ( .A(n59315), .B(n2304), .Z(n2306) );
  NAND U2587 ( .A(n2305), .B(n2306), .Z(n2307) );
  NAND U2588 ( .A(n59316), .B(n2307), .Z(n2308) );
  AND U2589 ( .A(n59317), .B(n2308), .Z(n2309) );
  NAND U2590 ( .A(n2309), .B(n59318), .Z(n2310) );
  AND U2591 ( .A(n59320), .B(n59321), .Z(n2311) );
  NANDN U2592 ( .A(n59319), .B(n2310), .Z(n2312) );
  NAND U2593 ( .A(n2311), .B(n2312), .Z(n2313) );
  NAND U2594 ( .A(n59322), .B(n2313), .Z(n2314) );
  AND U2595 ( .A(n59323), .B(n2314), .Z(n2315) );
  NAND U2596 ( .A(n2315), .B(n59324), .Z(n2316) );
  NAND U2597 ( .A(n59325), .B(n2316), .Z(n59327) );
  OR U2598 ( .A(n59355), .B(n59354), .Z(n2317) );
  AND U2599 ( .A(n59356), .B(n2317), .Z(n2318) );
  AND U2600 ( .A(n59359), .B(n59358), .Z(n2319) );
  NANDN U2601 ( .A(n2318), .B(n59357), .Z(n2320) );
  NAND U2602 ( .A(n2319), .B(n2320), .Z(n2321) );
  NAND U2603 ( .A(n59360), .B(n2321), .Z(n2322) );
  AND U2604 ( .A(n59362), .B(n2322), .Z(n2323) );
  NANDN U2605 ( .A(n59361), .B(n2323), .Z(n2324) );
  NAND U2606 ( .A(n59363), .B(n2324), .Z(n2325) );
  AND U2607 ( .A(n51010), .B(n2325), .Z(n2326) );
  NANDN U2608 ( .A(n51011), .B(n2326), .Z(n2327) );
  NAND U2609 ( .A(n59364), .B(n2327), .Z(n2328) );
  AND U2610 ( .A(n59366), .B(n2328), .Z(n2329) );
  NANDN U2611 ( .A(n59365), .B(n2329), .Z(n2330) );
  NAND U2612 ( .A(n59367), .B(n2330), .Z(n2331) );
  AND U2613 ( .A(n51009), .B(n2331), .Z(n2332) );
  NANDN U2614 ( .A(n51008), .B(n2332), .Z(n59368) );
  NAND U2615 ( .A(n59411), .B(n59412), .Z(n2333) );
  ANDN U2616 ( .B(n2333), .A(n59413), .Z(n2334) );
  NOR U2617 ( .A(n59414), .B(n2334), .Z(n2335) );
  NAND U2618 ( .A(n59415), .B(n2335), .Z(n2336) );
  NANDN U2619 ( .A(n59416), .B(n2336), .Z(n2337) );
  AND U2620 ( .A(n50990), .B(n50989), .Z(n2338) );
  NAND U2621 ( .A(n2337), .B(n2338), .Z(n2339) );
  NAND U2622 ( .A(n59417), .B(n2339), .Z(n2340) );
  AND U2623 ( .A(n50988), .B(n50987), .Z(n2341) );
  NAND U2624 ( .A(n2340), .B(n2341), .Z(n2342) );
  NAND U2625 ( .A(n59418), .B(n2342), .Z(n2343) );
  ANDN U2626 ( .B(n59419), .A(n59420), .Z(n2344) );
  NAND U2627 ( .A(n2343), .B(n2344), .Z(n2345) );
  NAND U2628 ( .A(n59421), .B(n2345), .Z(n2346) );
  ANDN U2629 ( .B(n50986), .A(n50985), .Z(n2347) );
  NAND U2630 ( .A(n2346), .B(n2347), .Z(n2348) );
  NAND U2631 ( .A(n59422), .B(n2348), .Z(n2349) );
  AND U2632 ( .A(n59423), .B(n2349), .Z(n59425) );
  NAND U2633 ( .A(n59452), .B(n59453), .Z(n2350) );
  AND U2634 ( .A(n59454), .B(n2350), .Z(n2351) );
  NANDN U2635 ( .A(n59455), .B(n2351), .Z(n2352) );
  NAND U2636 ( .A(n59456), .B(n2352), .Z(n2353) );
  AND U2637 ( .A(n50977), .B(n2353), .Z(n2354) );
  NANDN U2638 ( .A(n50976), .B(n2354), .Z(n2355) );
  AND U2639 ( .A(n59459), .B(n59458), .Z(n2356) );
  NANDN U2640 ( .A(n59457), .B(n2355), .Z(n2357) );
  NAND U2641 ( .A(n2356), .B(n2357), .Z(n2358) );
  NAND U2642 ( .A(n59460), .B(n2358), .Z(n2359) );
  AND U2643 ( .A(n59461), .B(n2359), .Z(n2360) );
  NAND U2644 ( .A(n2360), .B(n59462), .Z(n2361) );
  AND U2645 ( .A(n59464), .B(n59465), .Z(n2362) );
  NANDN U2646 ( .A(n59463), .B(n2361), .Z(n2363) );
  NAND U2647 ( .A(n2362), .B(n2363), .Z(n2364) );
  NAND U2648 ( .A(n59466), .B(n2364), .Z(n2365) );
  AND U2649 ( .A(n59468), .B(n2365), .Z(n2366) );
  NANDN U2650 ( .A(n59467), .B(n2366), .Z(n2367) );
  NAND U2651 ( .A(n59469), .B(n2367), .Z(n59470) );
  ANDN U2652 ( .B(n50969), .A(n50968), .Z(n2368) );
  OR U2653 ( .A(n59501), .B(n59502), .Z(n2369) );
  NAND U2654 ( .A(n2368), .B(n2369), .Z(n2370) );
  ANDN U2655 ( .B(n59505), .A(n59504), .Z(n2371) );
  NANDN U2656 ( .A(n59503), .B(n2370), .Z(n2372) );
  NAND U2657 ( .A(n2371), .B(n2372), .Z(n2373) );
  NAND U2658 ( .A(n59506), .B(n2373), .Z(n2374) );
  AND U2659 ( .A(n59507), .B(n2374), .Z(n2375) );
  NANDN U2660 ( .A(n50967), .B(n2375), .Z(n2376) );
  ANDN U2661 ( .B(n59510), .A(n59509), .Z(n2377) );
  NANDN U2662 ( .A(n59508), .B(n2376), .Z(n2378) );
  NAND U2663 ( .A(n2377), .B(n2378), .Z(n2379) );
  NAND U2664 ( .A(n59511), .B(n2379), .Z(n2380) );
  AND U2665 ( .A(n59512), .B(n2380), .Z(n2381) );
  NAND U2666 ( .A(n2381), .B(n59513), .Z(n2382) );
  NAND U2667 ( .A(n59514), .B(n2382), .Z(n2383) );
  AND U2668 ( .A(n50966), .B(n2383), .Z(n2384) );
  NANDN U2669 ( .A(n50965), .B(n2384), .Z(n59515) );
  NAND U2670 ( .A(n59550), .B(n59551), .Z(n2385) );
  ANDN U2671 ( .B(n2385), .A(n59552), .Z(n2386) );
  ANDN U2672 ( .B(n50956), .A(n2386), .Z(n2387) );
  NAND U2673 ( .A(n50957), .B(n2387), .Z(n2388) );
  NAND U2674 ( .A(n59553), .B(n2388), .Z(n2389) );
  ANDN U2675 ( .B(n59554), .A(n59555), .Z(n2390) );
  NAND U2676 ( .A(n2389), .B(n2390), .Z(n2391) );
  NAND U2677 ( .A(n59556), .B(n2391), .Z(n2392) );
  ANDN U2678 ( .B(n50955), .A(n50954), .Z(n2393) );
  NAND U2679 ( .A(n2392), .B(n2393), .Z(n2394) );
  NAND U2680 ( .A(n59557), .B(n2394), .Z(n2395) );
  AND U2681 ( .A(n59559), .B(n59558), .Z(n2396) );
  NAND U2682 ( .A(n2395), .B(n2396), .Z(n2397) );
  NAND U2683 ( .A(n59560), .B(n2397), .Z(n2398) );
  ANDN U2684 ( .B(n2398), .A(n59561), .Z(n59563) );
  NAND U2685 ( .A(n59625), .B(n59624), .Z(n2399) );
  NAND U2686 ( .A(n59626), .B(n2399), .Z(n2400) );
  AND U2687 ( .A(n59627), .B(n2400), .Z(n2401) );
  AND U2688 ( .A(n50937), .B(n50938), .Z(n2402) );
  OR U2689 ( .A(n2401), .B(n59628), .Z(n2403) );
  NAND U2690 ( .A(n2402), .B(n2403), .Z(n2404) );
  NAND U2691 ( .A(n59629), .B(n2404), .Z(n2405) );
  AND U2692 ( .A(n59631), .B(n2405), .Z(n2406) );
  NAND U2693 ( .A(n2406), .B(n59630), .Z(n2407) );
  ANDN U2694 ( .B(n50936), .A(n50935), .Z(n2408) );
  NANDN U2695 ( .A(n59632), .B(n2407), .Z(n2409) );
  NAND U2696 ( .A(n2408), .B(n2409), .Z(n2410) );
  NAND U2697 ( .A(n59633), .B(n2410), .Z(n2411) );
  AND U2698 ( .A(n59635), .B(n2411), .Z(n2412) );
  NANDN U2699 ( .A(n59634), .B(n2412), .Z(n2413) );
  NAND U2700 ( .A(n59636), .B(n2413), .Z(n2414) );
  AND U2701 ( .A(n59638), .B(n2414), .Z(n2415) );
  NAND U2702 ( .A(n2415), .B(n59637), .Z(n2416) );
  NANDN U2703 ( .A(n59639), .B(n2416), .Z(n59640) );
  ANDN U2704 ( .B(n59672), .A(n59671), .Z(n2417) );
  NANDN U2705 ( .A(n59670), .B(n59669), .Z(n2418) );
  AND U2706 ( .A(n2417), .B(n2418), .Z(n2419) );
  ANDN U2707 ( .B(n59674), .A(n50925), .Z(n2420) );
  NANDN U2708 ( .A(n2419), .B(n59673), .Z(n2421) );
  AND U2709 ( .A(n2420), .B(n2421), .Z(n2422) );
  ANDN U2710 ( .B(n59677), .A(n59676), .Z(n2423) );
  OR U2711 ( .A(n2422), .B(n59675), .Z(n2424) );
  AND U2712 ( .A(n2423), .B(n2424), .Z(n2425) );
  ANDN U2713 ( .B(n59679), .A(n59680), .Z(n2426) );
  NANDN U2714 ( .A(n2425), .B(n59678), .Z(n2427) );
  AND U2715 ( .A(n2426), .B(n2427), .Z(n2428) );
  ANDN U2716 ( .B(n50924), .A(n50923), .Z(n2429) );
  NANDN U2717 ( .A(n2428), .B(n59681), .Z(n2430) );
  AND U2718 ( .A(n2429), .B(n2430), .Z(n2431) );
  NANDN U2719 ( .A(n2431), .B(n59682), .Z(n2432) );
  AND U2720 ( .A(n59683), .B(n2432), .Z(n59686) );
  NOR U2721 ( .A(n50916), .B(n50917), .Z(n2433) );
  NAND U2722 ( .A(n59717), .B(n2433), .Z(n2434) );
  NAND U2723 ( .A(n59718), .B(n2434), .Z(n2435) );
  ANDN U2724 ( .B(n59720), .A(n59719), .Z(n2436) );
  NAND U2725 ( .A(n2435), .B(n2436), .Z(n2437) );
  NAND U2726 ( .A(n59721), .B(n2437), .Z(n2438) );
  AND U2727 ( .A(n50914), .B(n50913), .Z(n2439) );
  NAND U2728 ( .A(n2438), .B(n2439), .Z(n2440) );
  NANDN U2729 ( .A(n59722), .B(n2440), .Z(n2441) );
  AND U2730 ( .A(n59724), .B(n59723), .Z(n2442) );
  NAND U2731 ( .A(n2441), .B(n2442), .Z(n2443) );
  NAND U2732 ( .A(n59725), .B(n2443), .Z(n2444) );
  ANDN U2733 ( .B(n59726), .A(n50912), .Z(n2445) );
  NAND U2734 ( .A(n2444), .B(n2445), .Z(n2446) );
  NAND U2735 ( .A(n50911), .B(n2446), .Z(n2447) );
  ANDN U2736 ( .B(n59728), .A(n59727), .Z(n2448) );
  NAND U2737 ( .A(n2447), .B(n2448), .Z(n2449) );
  NAND U2738 ( .A(n59729), .B(n2449), .Z(n59730) );
  ANDN U2739 ( .B(n50902), .A(n50903), .Z(n2450) );
  NANDN U2740 ( .A(n50904), .B(n59763), .Z(n2451) );
  NAND U2741 ( .A(n2450), .B(n2451), .Z(n2452) );
  NAND U2742 ( .A(n59764), .B(n2452), .Z(n2453) );
  AND U2743 ( .A(n59765), .B(n2453), .Z(n2454) );
  NANDN U2744 ( .A(n59766), .B(n2454), .Z(n2455) );
  ANDN U2745 ( .B(n50901), .A(n50900), .Z(n2456) );
  NANDN U2746 ( .A(n59767), .B(n2455), .Z(n2457) );
  NAND U2747 ( .A(n2456), .B(n2457), .Z(n2458) );
  AND U2748 ( .A(n59769), .B(n59770), .Z(n2459) );
  NANDN U2749 ( .A(n59768), .B(n2458), .Z(n2460) );
  NAND U2750 ( .A(n2459), .B(n2460), .Z(n2461) );
  NAND U2751 ( .A(n59771), .B(n2461), .Z(n2462) );
  AND U2752 ( .A(n59773), .B(n2462), .Z(n2463) );
  NANDN U2753 ( .A(n59772), .B(n2463), .Z(n2464) );
  AND U2754 ( .A(n59776), .B(n59775), .Z(n2465) );
  NANDN U2755 ( .A(n59774), .B(n2464), .Z(n2466) );
  NAND U2756 ( .A(n2465), .B(n2466), .Z(n59777) );
  AND U2757 ( .A(n59805), .B(n59806), .Z(n2467) );
  NAND U2758 ( .A(n50890), .B(n2467), .Z(n2468) );
  NAND U2759 ( .A(n59807), .B(n2468), .Z(n2469) );
  NAND U2760 ( .A(n50889), .B(n2469), .Z(n2470) );
  AND U2761 ( .A(n59809), .B(n59810), .Z(n2471) );
  NANDN U2762 ( .A(n59808), .B(n2470), .Z(n2472) );
  NAND U2763 ( .A(n2471), .B(n2472), .Z(n2473) );
  NAND U2764 ( .A(n59811), .B(n2473), .Z(n2474) );
  AND U2765 ( .A(n59812), .B(n2474), .Z(n2475) );
  NAND U2766 ( .A(n2475), .B(n59813), .Z(n2476) );
  AND U2767 ( .A(n59815), .B(n59816), .Z(n2477) );
  NANDN U2768 ( .A(n59814), .B(n2476), .Z(n2478) );
  NAND U2769 ( .A(n2477), .B(n2478), .Z(n2479) );
  NAND U2770 ( .A(n59817), .B(n2479), .Z(n2480) );
  AND U2771 ( .A(n50887), .B(n2480), .Z(n2481) );
  NAND U2772 ( .A(n2481), .B(n50888), .Z(n59820) );
  ANDN U2773 ( .B(n59851), .A(n59852), .Z(n2482) );
  NAND U2774 ( .A(n59850), .B(n59849), .Z(n2483) );
  AND U2775 ( .A(n2482), .B(n2483), .Z(n2484) );
  ANDN U2776 ( .B(n50876), .A(n50875), .Z(n2485) );
  OR U2777 ( .A(n59853), .B(n2484), .Z(n2486) );
  AND U2778 ( .A(n2485), .B(n2486), .Z(n2487) );
  AND U2779 ( .A(n59855), .B(n59854), .Z(n2488) );
  NANDN U2780 ( .A(n2487), .B(n50874), .Z(n2489) );
  AND U2781 ( .A(n2488), .B(n2489), .Z(n2490) );
  ANDN U2782 ( .B(n59858), .A(n59857), .Z(n2491) );
  NANDN U2783 ( .A(n2490), .B(n59856), .Z(n2492) );
  AND U2784 ( .A(n2491), .B(n2492), .Z(n2493) );
  AND U2785 ( .A(n59860), .B(n59861), .Z(n2494) );
  NANDN U2786 ( .A(n2493), .B(n59859), .Z(n2495) );
  AND U2787 ( .A(n2494), .B(n2495), .Z(n2496) );
  NANDN U2788 ( .A(n2496), .B(n59862), .Z(n2497) );
  ANDN U2789 ( .B(n2497), .A(n59863), .Z(n59865) );
  NAND U2790 ( .A(n59891), .B(n59892), .Z(n2498) );
  AND U2791 ( .A(n59894), .B(n2498), .Z(n2499) );
  NANDN U2792 ( .A(n59893), .B(n2499), .Z(n2500) );
  NAND U2793 ( .A(n59895), .B(n2500), .Z(n2501) );
  AND U2794 ( .A(n59896), .B(n2501), .Z(n2502) );
  NAND U2795 ( .A(n2502), .B(n59897), .Z(n2503) );
  NAND U2796 ( .A(n59898), .B(n2503), .Z(n2504) );
  AND U2797 ( .A(n59900), .B(n2504), .Z(n2505) );
  NANDN U2798 ( .A(n59899), .B(n2505), .Z(n2506) );
  NAND U2799 ( .A(n59901), .B(n2506), .Z(n2507) );
  AND U2800 ( .A(n50865), .B(n2507), .Z(n2508) );
  NANDN U2801 ( .A(n50866), .B(n2508), .Z(n2509) );
  NAND U2802 ( .A(n59902), .B(n2509), .Z(n2510) );
  AND U2803 ( .A(n59904), .B(n2510), .Z(n2511) );
  NANDN U2804 ( .A(n59903), .B(n2511), .Z(n2512) );
  NAND U2805 ( .A(n59905), .B(n2512), .Z(n2513) );
  AND U2806 ( .A(n50864), .B(n2513), .Z(n2514) );
  NANDN U2807 ( .A(n50863), .B(n2514), .Z(n59906) );
  AND U2808 ( .A(n50854), .B(n50855), .Z(n2515) );
  OR U2809 ( .A(n59934), .B(n59935), .Z(n2516) );
  NAND U2810 ( .A(n2515), .B(n2516), .Z(n2517) );
  NAND U2811 ( .A(n50852), .B(n2517), .Z(n2518) );
  AND U2812 ( .A(n59937), .B(n2518), .Z(n2519) );
  NANDN U2813 ( .A(n59936), .B(n2519), .Z(n2520) );
  NAND U2814 ( .A(n59938), .B(n2520), .Z(n2521) );
  AND U2815 ( .A(n59939), .B(n2521), .Z(n2522) );
  NANDN U2816 ( .A(n50851), .B(n2522), .Z(n2523) );
  ANDN U2817 ( .B(n59942), .A(n59941), .Z(n2524) );
  NANDN U2818 ( .A(n59940), .B(n2523), .Z(n2525) );
  NAND U2819 ( .A(n2524), .B(n2525), .Z(n2526) );
  NAND U2820 ( .A(n59943), .B(n2526), .Z(n2527) );
  AND U2821 ( .A(n59944), .B(n2527), .Z(n2528) );
  NAND U2822 ( .A(n2528), .B(n59945), .Z(n2529) );
  NAND U2823 ( .A(n59946), .B(n2529), .Z(n2530) );
  AND U2824 ( .A(n50850), .B(n2530), .Z(n2531) );
  NANDN U2825 ( .A(n50849), .B(n2531), .Z(n59947) );
  NAND U2826 ( .A(n59980), .B(n59979), .Z(n2532) );
  AND U2827 ( .A(n59981), .B(n2532), .Z(n2533) );
  NOR U2828 ( .A(n59983), .B(n2533), .Z(n2534) );
  NAND U2829 ( .A(n59982), .B(n2534), .Z(n2535) );
  NANDN U2830 ( .A(n50841), .B(n2535), .Z(n2536) );
  ANDN U2831 ( .B(n59985), .A(n59984), .Z(n2537) );
  NAND U2832 ( .A(n2536), .B(n2537), .Z(n2538) );
  NAND U2833 ( .A(n59986), .B(n2538), .Z(n2539) );
  ANDN U2834 ( .B(n59987), .A(n59988), .Z(n2540) );
  NAND U2835 ( .A(n2539), .B(n2540), .Z(n2541) );
  NAND U2836 ( .A(n59989), .B(n2541), .Z(n2542) );
  ANDN U2837 ( .B(n50840), .A(n50839), .Z(n2543) );
  NAND U2838 ( .A(n2542), .B(n2543), .Z(n2544) );
  NANDN U2839 ( .A(n59990), .B(n2544), .Z(n2545) );
  NAND U2840 ( .A(n59991), .B(n2545), .Z(n2546) );
  NAND U2841 ( .A(n59992), .B(n2546), .Z(n2547) );
  AND U2842 ( .A(n50838), .B(n2547), .Z(n2548) );
  NAND U2843 ( .A(n2548), .B(n50837), .Z(n59993) );
  NAND U2844 ( .A(n60016), .B(n60017), .Z(n2549) );
  AND U2845 ( .A(n60019), .B(n2549), .Z(n2550) );
  NANDN U2846 ( .A(n60018), .B(n2550), .Z(n2551) );
  NAND U2847 ( .A(n60020), .B(n2551), .Z(n2552) );
  ANDN U2848 ( .B(n2552), .A(n50824), .Z(n2553) );
  NANDN U2849 ( .A(n50825), .B(n2553), .Z(n2554) );
  NAND U2850 ( .A(n60021), .B(n2554), .Z(n2555) );
  AND U2851 ( .A(n60023), .B(n2555), .Z(n2556) );
  NANDN U2852 ( .A(n60022), .B(n2556), .Z(n2557) );
  AND U2853 ( .A(n50822), .B(n50823), .Z(n2558) );
  NANDN U2854 ( .A(n60024), .B(n2557), .Z(n2559) );
  NAND U2855 ( .A(n2558), .B(n2559), .Z(n2560) );
  NAND U2856 ( .A(n50821), .B(n2560), .Z(n2561) );
  AND U2857 ( .A(n60025), .B(n2561), .Z(n2562) );
  NAND U2858 ( .A(n2562), .B(n60026), .Z(n2563) );
  NAND U2859 ( .A(n60027), .B(n2563), .Z(n2564) );
  AND U2860 ( .A(n60028), .B(n2564), .Z(n2565) );
  NAND U2861 ( .A(n2565), .B(n60029), .Z(n60030) );
  NAND U2862 ( .A(n60059), .B(n60058), .Z(n2566) );
  NAND U2863 ( .A(n60060), .B(n2566), .Z(n2567) );
  AND U2864 ( .A(n60061), .B(n2567), .Z(n2568) );
  AND U2865 ( .A(n60064), .B(n60063), .Z(n2569) );
  NANDN U2866 ( .A(n2568), .B(n60062), .Z(n2570) );
  AND U2867 ( .A(n2569), .B(n2570), .Z(n2571) );
  AND U2868 ( .A(n60066), .B(n60067), .Z(n2572) );
  NANDN U2869 ( .A(n2571), .B(n60065), .Z(n2573) );
  AND U2870 ( .A(n2572), .B(n2573), .Z(n2574) );
  ANDN U2871 ( .B(n60070), .A(n60069), .Z(n2575) );
  NANDN U2872 ( .A(n2574), .B(n60068), .Z(n2576) );
  AND U2873 ( .A(n2575), .B(n2576), .Z(n2577) );
  AND U2874 ( .A(n60071), .B(n60072), .Z(n2578) );
  NANDN U2875 ( .A(n2577), .B(n50811), .Z(n2579) );
  AND U2876 ( .A(n2578), .B(n2579), .Z(n2580) );
  NANDN U2877 ( .A(n2580), .B(n60073), .Z(n2581) );
  ANDN U2878 ( .B(n2581), .A(n60074), .Z(n60076) );
  NAND U2879 ( .A(n60100), .B(n60099), .Z(n2582) );
  NAND U2880 ( .A(n60101), .B(n2582), .Z(n2583) );
  ANDN U2881 ( .B(n2583), .A(n60102), .Z(n2584) );
  NAND U2882 ( .A(n60103), .B(n2584), .Z(n2585) );
  NANDN U2883 ( .A(n60104), .B(n2585), .Z(n2586) );
  AND U2884 ( .A(n60105), .B(n2586), .Z(n2587) );
  NAND U2885 ( .A(n60106), .B(n2587), .Z(n2588) );
  NAND U2886 ( .A(n60107), .B(n2588), .Z(n2589) );
  NANDN U2887 ( .A(n60108), .B(n2589), .Z(n2590) );
  NAND U2888 ( .A(n60109), .B(n2590), .Z(n2591) );
  AND U2889 ( .A(n50799), .B(n2591), .Z(n2592) );
  NANDN U2890 ( .A(n50798), .B(n2592), .Z(n2593) );
  NAND U2891 ( .A(n60110), .B(n2593), .Z(n2594) );
  AND U2892 ( .A(n60112), .B(n2594), .Z(n2595) );
  NANDN U2893 ( .A(n60111), .B(n2595), .Z(n2596) );
  NAND U2894 ( .A(n50797), .B(n2596), .Z(n60113) );
  NANDN U2895 ( .A(n50788), .B(n60145), .Z(n2597) );
  ANDN U2896 ( .B(n2597), .A(n60146), .Z(n2598) );
  NOR U2897 ( .A(n60147), .B(n2598), .Z(n2599) );
  NAND U2898 ( .A(n60148), .B(n2599), .Z(n2600) );
  NAND U2899 ( .A(n60149), .B(n2600), .Z(n2601) );
  AND U2900 ( .A(n60151), .B(n60150), .Z(n2602) );
  NAND U2901 ( .A(n2601), .B(n2602), .Z(n2603) );
  NAND U2902 ( .A(n60152), .B(n2603), .Z(n2604) );
  ANDN U2903 ( .B(n50787), .A(n50786), .Z(n2605) );
  NAND U2904 ( .A(n2604), .B(n2605), .Z(n2606) );
  NAND U2905 ( .A(n60153), .B(n2606), .Z(n2607) );
  AND U2906 ( .A(n60155), .B(n60154), .Z(n2608) );
  NAND U2907 ( .A(n2607), .B(n2608), .Z(n2609) );
  NAND U2908 ( .A(n60156), .B(n2609), .Z(n2610) );
  NAND U2909 ( .A(n60157), .B(n2610), .Z(n2611) );
  NANDN U2910 ( .A(n60158), .B(n2611), .Z(n2612) );
  AND U2911 ( .A(n60159), .B(n2612), .Z(n2613) );
  NANDN U2912 ( .A(n2613), .B(n60160), .Z(n2614) );
  AND U2913 ( .A(n60161), .B(n2614), .Z(n60163) );
  NAND U2914 ( .A(n60189), .B(n60188), .Z(n2615) );
  AND U2915 ( .A(n60190), .B(n2615), .Z(n2616) );
  ANDN U2916 ( .B(n50775), .A(n2616), .Z(n2617) );
  NAND U2917 ( .A(n50774), .B(n2617), .Z(n2618) );
  NAND U2918 ( .A(n60191), .B(n2618), .Z(n2619) );
  AND U2919 ( .A(n60192), .B(n60193), .Z(n2620) );
  NAND U2920 ( .A(n2619), .B(n2620), .Z(n2621) );
  NAND U2921 ( .A(n60194), .B(n2621), .Z(n2622) );
  ANDN U2922 ( .B(n50773), .A(n50772), .Z(n2623) );
  NAND U2923 ( .A(n2622), .B(n2623), .Z(n2624) );
  NANDN U2924 ( .A(n60195), .B(n2624), .Z(n2625) );
  ANDN U2925 ( .B(n60197), .A(n60196), .Z(n2626) );
  NAND U2926 ( .A(n2625), .B(n2626), .Z(n2627) );
  NAND U2927 ( .A(n60198), .B(n2627), .Z(n2628) );
  ANDN U2928 ( .B(n60199), .A(n50771), .Z(n2629) );
  NAND U2929 ( .A(n2628), .B(n2629), .Z(n2630) );
  NAND U2930 ( .A(n60200), .B(n2630), .Z(n60202) );
  NAND U2931 ( .A(n50762), .B(n60229), .Z(n2631) );
  AND U2932 ( .A(n60230), .B(n2631), .Z(n2632) );
  NAND U2933 ( .A(n2632), .B(n60231), .Z(n2633) );
  NAND U2934 ( .A(n60232), .B(n2633), .Z(n2634) );
  AND U2935 ( .A(n60233), .B(n2634), .Z(n2635) );
  NANDN U2936 ( .A(n60234), .B(n2635), .Z(n2636) );
  NAND U2937 ( .A(n60235), .B(n2636), .Z(n2637) );
  AND U2938 ( .A(n50760), .B(n2637), .Z(n2638) );
  NANDN U2939 ( .A(n50761), .B(n2638), .Z(n2639) );
  NAND U2940 ( .A(n60236), .B(n2639), .Z(n2640) );
  AND U2941 ( .A(n60238), .B(n2640), .Z(n2641) );
  NAND U2942 ( .A(n2641), .B(n60237), .Z(n2642) );
  AND U2943 ( .A(n60241), .B(n60240), .Z(n2643) );
  NANDN U2944 ( .A(n60239), .B(n2642), .Z(n2644) );
  NAND U2945 ( .A(n2643), .B(n2644), .Z(n60242) );
  NAND U2946 ( .A(n60267), .B(n60268), .Z(n2645) );
  NAND U2947 ( .A(n60269), .B(n2645), .Z(n2646) );
  NAND U2948 ( .A(n60270), .B(n2646), .Z(n2647) );
  ANDN U2949 ( .B(n50749), .A(n50748), .Z(n2648) );
  NAND U2950 ( .A(n2647), .B(n2648), .Z(n2649) );
  NAND U2951 ( .A(n60271), .B(n2649), .Z(n2650) );
  ANDN U2952 ( .B(n60273), .A(n60272), .Z(n2651) );
  NAND U2953 ( .A(n2650), .B(n2651), .Z(n2652) );
  NAND U2954 ( .A(n60274), .B(n2652), .Z(n2653) );
  AND U2955 ( .A(n50746), .B(n50747), .Z(n2654) );
  NAND U2956 ( .A(n2653), .B(n2654), .Z(n2655) );
  NAND U2957 ( .A(n50745), .B(n2655), .Z(n2656) );
  ANDN U2958 ( .B(n60276), .A(n60275), .Z(n2657) );
  NAND U2959 ( .A(n2656), .B(n2657), .Z(n2658) );
  NAND U2960 ( .A(n60277), .B(n2658), .Z(n2659) );
  NAND U2961 ( .A(n60278), .B(n2659), .Z(n60279) );
  NAND U2962 ( .A(n60309), .B(n60310), .Z(n2660) );
  AND U2963 ( .A(n60311), .B(n2660), .Z(n2661) );
  NAND U2964 ( .A(n2661), .B(n60312), .Z(n2662) );
  AND U2965 ( .A(n60313), .B(n60314), .Z(n2663) );
  NANDN U2966 ( .A(n50739), .B(n2662), .Z(n2664) );
  NAND U2967 ( .A(n2663), .B(n2664), .Z(n2665) );
  ANDN U2968 ( .B(n50738), .A(n50737), .Z(n2666) );
  NANDN U2969 ( .A(n60315), .B(n2665), .Z(n2667) );
  NAND U2970 ( .A(n2666), .B(n2667), .Z(n2668) );
  NAND U2971 ( .A(n50736), .B(n2668), .Z(n2669) );
  AND U2972 ( .A(n60316), .B(n2669), .Z(n2670) );
  NANDN U2973 ( .A(n60317), .B(n2670), .Z(n2671) );
  AND U2974 ( .A(n60320), .B(n60319), .Z(n2672) );
  NANDN U2975 ( .A(n60318), .B(n2671), .Z(n2673) );
  NAND U2976 ( .A(n2672), .B(n2673), .Z(n2674) );
  AND U2977 ( .A(n60321), .B(n2674), .Z(n60322) );
  NANDN U2978 ( .A(n60351), .B(n60350), .Z(n2675) );
  AND U2979 ( .A(n60352), .B(n2675), .Z(n2676) );
  NOR U2980 ( .A(n60354), .B(n2676), .Z(n2677) );
  NAND U2981 ( .A(n60353), .B(n2677), .Z(n2678) );
  NAND U2982 ( .A(n60355), .B(n2678), .Z(n2679) );
  ANDN U2983 ( .B(n60357), .A(n60356), .Z(n2680) );
  NAND U2984 ( .A(n2679), .B(n2680), .Z(n2681) );
  NAND U2985 ( .A(n60358), .B(n2681), .Z(n2682) );
  ANDN U2986 ( .B(n60360), .A(n60359), .Z(n2683) );
  NAND U2987 ( .A(n2682), .B(n2683), .Z(n2684) );
  NANDN U2988 ( .A(n60361), .B(n2684), .Z(n2685) );
  ANDN U2989 ( .B(n60363), .A(n60362), .Z(n2686) );
  NAND U2990 ( .A(n2685), .B(n2686), .Z(n2687) );
  NAND U2991 ( .A(n60364), .B(n2687), .Z(n2688) );
  ANDN U2992 ( .B(n60365), .A(n60366), .Z(n2689) );
  NAND U2993 ( .A(n2688), .B(n2689), .Z(n2690) );
  NANDN U2994 ( .A(n60367), .B(n2690), .Z(n60368) );
  NAND U2995 ( .A(n60391), .B(n60392), .Z(n2691) );
  NAND U2996 ( .A(n60393), .B(n2691), .Z(n2692) );
  NAND U2997 ( .A(n60394), .B(n2692), .Z(n2693) );
  NAND U2998 ( .A(n60395), .B(n2693), .Z(n2694) );
  NANDN U2999 ( .A(n60396), .B(n2694), .Z(n2695) );
  AND U3000 ( .A(n60397), .B(n2695), .Z(n2696) );
  NANDN U3001 ( .A(n2696), .B(n60398), .Z(n2697) );
  AND U3002 ( .A(n60399), .B(n2697), .Z(n2698) );
  NANDN U3003 ( .A(n2698), .B(n60400), .Z(n2699) );
  NAND U3004 ( .A(n60401), .B(n2699), .Z(n2700) );
  NANDN U3005 ( .A(n60402), .B(n2700), .Z(n2701) );
  AND U3006 ( .A(n50710), .B(n50711), .Z(n2702) );
  NAND U3007 ( .A(n2701), .B(n2702), .Z(n2703) );
  NAND U3008 ( .A(n60403), .B(n2703), .Z(n2704) );
  ANDN U3009 ( .B(n60404), .A(n60405), .Z(n2705) );
  NAND U3010 ( .A(n2704), .B(n2705), .Z(n2706) );
  NANDN U3011 ( .A(n60406), .B(n2706), .Z(n60407) );
  NAND U3012 ( .A(n60436), .B(n60437), .Z(n2707) );
  AND U3013 ( .A(n60439), .B(n2707), .Z(n2708) );
  NANDN U3014 ( .A(n60438), .B(n2708), .Z(n2709) );
  ANDN U3015 ( .B(n50700), .A(n50701), .Z(n2710) );
  NANDN U3016 ( .A(n60440), .B(n2709), .Z(n2711) );
  NAND U3017 ( .A(n2710), .B(n2711), .Z(n2712) );
  NAND U3018 ( .A(n60441), .B(n2712), .Z(n2713) );
  AND U3019 ( .A(n60443), .B(n2713), .Z(n2714) );
  NANDN U3020 ( .A(n60442), .B(n2714), .Z(n2715) );
  NAND U3021 ( .A(n60444), .B(n2715), .Z(n2716) );
  AND U3022 ( .A(n50699), .B(n2716), .Z(n2717) );
  NANDN U3023 ( .A(n50698), .B(n2717), .Z(n2718) );
  ANDN U3024 ( .B(n60447), .A(n60446), .Z(n2719) );
  NANDN U3025 ( .A(n60445), .B(n2718), .Z(n2720) );
  NAND U3026 ( .A(n2719), .B(n2720), .Z(n2721) );
  NAND U3027 ( .A(n60448), .B(n2721), .Z(n60449) );
  NAND U3028 ( .A(n60479), .B(n60478), .Z(n2722) );
  ANDN U3029 ( .B(n2722), .A(n60481), .Z(n2723) );
  NOR U3030 ( .A(n50688), .B(n2723), .Z(n2724) );
  NAND U3031 ( .A(n50689), .B(n2724), .Z(n2725) );
  NANDN U3032 ( .A(n60482), .B(n2725), .Z(n2726) );
  ANDN U3033 ( .B(n60484), .A(n60483), .Z(n2727) );
  NAND U3034 ( .A(n2726), .B(n2727), .Z(n2728) );
  NAND U3035 ( .A(n60485), .B(n2728), .Z(n2729) );
  AND U3036 ( .A(n60487), .B(n60486), .Z(n2730) );
  NAND U3037 ( .A(n2729), .B(n2730), .Z(n2731) );
  NAND U3038 ( .A(n50687), .B(n2731), .Z(n2732) );
  ANDN U3039 ( .B(n60489), .A(n60488), .Z(n2733) );
  NAND U3040 ( .A(n2732), .B(n2733), .Z(n2734) );
  NAND U3041 ( .A(n60490), .B(n2734), .Z(n2735) );
  ANDN U3042 ( .B(n60492), .A(n60491), .Z(n2736) );
  NAND U3043 ( .A(n2735), .B(n2736), .Z(n2737) );
  NANDN U3044 ( .A(n60493), .B(n2737), .Z(n60495) );
  AND U3045 ( .A(n50669), .B(n50670), .Z(n2738) );
  NANDN U3046 ( .A(n60553), .B(n60552), .Z(n2739) );
  AND U3047 ( .A(n2738), .B(n2739), .Z(n2740) );
  NANDN U3048 ( .A(n2740), .B(n50667), .Z(n2741) );
  AND U3049 ( .A(n60554), .B(n2741), .Z(n2742) );
  AND U3050 ( .A(n50666), .B(n50665), .Z(n2743) );
  NANDN U3051 ( .A(n2742), .B(n60555), .Z(n2744) );
  NAND U3052 ( .A(n2743), .B(n2744), .Z(n2745) );
  AND U3053 ( .A(n50662), .B(n50663), .Z(n2746) );
  NANDN U3054 ( .A(n50664), .B(n2745), .Z(n2747) );
  NAND U3055 ( .A(n2746), .B(n2747), .Z(n2748) );
  NAND U3056 ( .A(n60556), .B(n2748), .Z(n2749) );
  AND U3057 ( .A(n60558), .B(n2749), .Z(n2750) );
  NANDN U3058 ( .A(n60557), .B(n2750), .Z(n2751) );
  NAND U3059 ( .A(n60559), .B(n2751), .Z(n2752) );
  AND U3060 ( .A(n50661), .B(n2752), .Z(n2753) );
  NAND U3061 ( .A(n2753), .B(n50660), .Z(n60560) );
  NAND U3062 ( .A(n60587), .B(n60586), .Z(n2754) );
  AND U3063 ( .A(n60589), .B(n2754), .Z(n2755) );
  NOR U3064 ( .A(n60591), .B(n60592), .Z(n2756) );
  NANDN U3065 ( .A(n2755), .B(n2756), .Z(n2757) );
  NANDN U3066 ( .A(n60593), .B(n2757), .Z(n2758) );
  ANDN U3067 ( .B(n60595), .A(n60594), .Z(n2759) );
  NAND U3068 ( .A(n2758), .B(n2759), .Z(n2760) );
  NAND U3069 ( .A(n60596), .B(n2760), .Z(n2761) );
  ANDN U3070 ( .B(n60597), .A(n60598), .Z(n2762) );
  NAND U3071 ( .A(n2761), .B(n2762), .Z(n2763) );
  NANDN U3072 ( .A(n50651), .B(n2763), .Z(n2764) );
  ANDN U3073 ( .B(n60600), .A(n60599), .Z(n2765) );
  NAND U3074 ( .A(n2764), .B(n2765), .Z(n2766) );
  NAND U3075 ( .A(n60601), .B(n2766), .Z(n2767) );
  AND U3076 ( .A(n50650), .B(n50649), .Z(n2768) );
  NAND U3077 ( .A(n2767), .B(n2768), .Z(n2769) );
  NAND U3078 ( .A(n60602), .B(n2769), .Z(n2770) );
  AND U3079 ( .A(n60603), .B(n2770), .Z(n60604) );
  AND U3080 ( .A(n50635), .B(n50634), .Z(n2771) );
  NAND U3081 ( .A(n60627), .B(n2771), .Z(n2772) );
  NAND U3082 ( .A(n60628), .B(n2772), .Z(n2773) );
  ANDN U3083 ( .B(n60630), .A(n60629), .Z(n2774) );
  NAND U3084 ( .A(n2773), .B(n2774), .Z(n2775) );
  NANDN U3085 ( .A(n60631), .B(n2775), .Z(n2776) );
  NOR U3086 ( .A(n60633), .B(n60632), .Z(n2777) );
  NAND U3087 ( .A(n2776), .B(n2777), .Z(n2778) );
  NAND U3088 ( .A(n50632), .B(n2778), .Z(n2779) );
  ANDN U3089 ( .B(n60635), .A(n60634), .Z(n2780) );
  NAND U3090 ( .A(n2779), .B(n2780), .Z(n2781) );
  NAND U3091 ( .A(n60636), .B(n2781), .Z(n2782) );
  ANDN U3092 ( .B(n50631), .A(n50630), .Z(n2783) );
  NAND U3093 ( .A(n2782), .B(n2783), .Z(n2784) );
  NAND U3094 ( .A(n60637), .B(n2784), .Z(n2785) );
  NAND U3095 ( .A(n60638), .B(n2785), .Z(n2786) );
  NAND U3096 ( .A(n60639), .B(n2786), .Z(n60641) );
  ANDN U3097 ( .B(n60709), .A(n60708), .Z(n2787) );
  NAND U3098 ( .A(n60710), .B(n2787), .Z(n2788) );
  NAND U3099 ( .A(n60711), .B(n2788), .Z(n2789) );
  ANDN U3100 ( .B(n50615), .A(n50616), .Z(n2790) );
  NAND U3101 ( .A(n2789), .B(n2790), .Z(n2791) );
  NAND U3102 ( .A(n60712), .B(n2791), .Z(n2792) );
  ANDN U3103 ( .B(n60714), .A(n60713), .Z(n2793) );
  NAND U3104 ( .A(n2792), .B(n2793), .Z(n2794) );
  NAND U3105 ( .A(n60715), .B(n2794), .Z(n2795) );
  ANDN U3106 ( .B(n50614), .A(n50613), .Z(n2796) );
  NAND U3107 ( .A(n2795), .B(n2796), .Z(n2797) );
  NAND U3108 ( .A(n50612), .B(n2797), .Z(n2798) );
  ANDN U3109 ( .B(n60717), .A(n60716), .Z(n2799) );
  NAND U3110 ( .A(n2798), .B(n2799), .Z(n2800) );
  NAND U3111 ( .A(n60718), .B(n2800), .Z(n2801) );
  AND U3112 ( .A(n60719), .B(n2801), .Z(n60720) );
  NAND U3113 ( .A(n60747), .B(n50602), .Z(n2802) );
  AND U3114 ( .A(n60748), .B(n2802), .Z(n2803) );
  NAND U3115 ( .A(n2803), .B(n60749), .Z(n2804) );
  NAND U3116 ( .A(n60750), .B(n2804), .Z(n2805) );
  AND U3117 ( .A(n60751), .B(n2805), .Z(n2806) );
  NAND U3118 ( .A(n2806), .B(n60752), .Z(n2807) );
  ANDN U3119 ( .B(n50601), .A(n50600), .Z(n2808) );
  NANDN U3120 ( .A(n60753), .B(n2807), .Z(n2809) );
  NAND U3121 ( .A(n2808), .B(n2809), .Z(n2810) );
  NAND U3122 ( .A(n60754), .B(n2810), .Z(n2811) );
  AND U3123 ( .A(n60755), .B(n2811), .Z(n2812) );
  NANDN U3124 ( .A(n60756), .B(n2812), .Z(n2813) );
  NAND U3125 ( .A(n60757), .B(n2813), .Z(n2814) );
  AND U3126 ( .A(n50599), .B(n2814), .Z(n2815) );
  NANDN U3127 ( .A(n50598), .B(n2815), .Z(n2816) );
  NANDN U3128 ( .A(n60758), .B(n2816), .Z(n60759) );
  AND U3129 ( .A(n50582), .B(n50583), .Z(n2817) );
  OR U3130 ( .A(n60822), .B(n60823), .Z(n2818) );
  NAND U3131 ( .A(n2817), .B(n2818), .Z(n2819) );
  ANDN U3132 ( .B(n60826), .A(n60825), .Z(n2820) );
  NANDN U3133 ( .A(n60824), .B(n2819), .Z(n2821) );
  NAND U3134 ( .A(n2820), .B(n2821), .Z(n2822) );
  NAND U3135 ( .A(n60827), .B(n2822), .Z(n2823) );
  AND U3136 ( .A(n60828), .B(n2823), .Z(n2824) );
  NANDN U3137 ( .A(n50580), .B(n2824), .Z(n2825) );
  ANDN U3138 ( .B(n60831), .A(n60830), .Z(n2826) );
  NANDN U3139 ( .A(n60829), .B(n2825), .Z(n2827) );
  NAND U3140 ( .A(n2826), .B(n2827), .Z(n2828) );
  NAND U3141 ( .A(n60832), .B(n2828), .Z(n2829) );
  AND U3142 ( .A(n60834), .B(n2829), .Z(n2830) );
  NAND U3143 ( .A(n2830), .B(n60833), .Z(n2831) );
  ANDN U3144 ( .B(n50579), .A(n50578), .Z(n2832) );
  NANDN U3145 ( .A(n60835), .B(n2831), .Z(n2833) );
  NAND U3146 ( .A(n2832), .B(n2833), .Z(n60836) );
  AND U3147 ( .A(n60871), .B(n60870), .Z(n2834) );
  OR U3148 ( .A(n60868), .B(n60869), .Z(n2835) );
  AND U3149 ( .A(n2834), .B(n2835), .Z(n2836) );
  ANDN U3150 ( .B(n60873), .A(n60874), .Z(n2837) );
  OR U3151 ( .A(n60872), .B(n2836), .Z(n2838) );
  AND U3152 ( .A(n2837), .B(n2838), .Z(n2839) );
  AND U3153 ( .A(n60876), .B(n60877), .Z(n2840) );
  NANDN U3154 ( .A(n2839), .B(n60875), .Z(n2841) );
  AND U3155 ( .A(n2840), .B(n2841), .Z(n2842) );
  NANDN U3156 ( .A(n2842), .B(n50568), .Z(n2843) );
  NANDN U3157 ( .A(n60878), .B(n2843), .Z(n2844) );
  NAND U3158 ( .A(n60879), .B(n2844), .Z(n2845) );
  AND U3159 ( .A(n50566), .B(n50567), .Z(n2846) );
  NAND U3160 ( .A(n2845), .B(n2846), .Z(n2847) );
  NANDN U3161 ( .A(n60880), .B(n2847), .Z(n2848) );
  AND U3162 ( .A(n60881), .B(n2848), .Z(n60884) );
  AND U3163 ( .A(n60909), .B(n60910), .Z(n2849) );
  NAND U3164 ( .A(n60911), .B(n2849), .Z(n2850) );
  NAND U3165 ( .A(n60912), .B(n2850), .Z(n2851) );
  AND U3166 ( .A(n60914), .B(n60913), .Z(n2852) );
  NAND U3167 ( .A(n2851), .B(n2852), .Z(n2853) );
  NAND U3168 ( .A(n50556), .B(n2853), .Z(n2854) );
  AND U3169 ( .A(n60915), .B(n60916), .Z(n2855) );
  NAND U3170 ( .A(n2854), .B(n2855), .Z(n2856) );
  NAND U3171 ( .A(n60917), .B(n2856), .Z(n2857) );
  ANDN U3172 ( .B(n60919), .A(n60918), .Z(n2858) );
  NAND U3173 ( .A(n2857), .B(n2858), .Z(n2859) );
  NANDN U3174 ( .A(n60920), .B(n2859), .Z(n2860) );
  ANDN U3175 ( .B(n50554), .A(n50555), .Z(n2861) );
  NAND U3176 ( .A(n2860), .B(n2861), .Z(n2862) );
  NAND U3177 ( .A(n60921), .B(n2862), .Z(n2863) );
  ANDN U3178 ( .B(n2863), .A(n60922), .Z(n2864) );
  AND U3179 ( .A(n60923), .B(n2864), .Z(n60926) );
  ANDN U3180 ( .B(n60954), .A(n60953), .Z(n2865) );
  NAND U3181 ( .A(n60955), .B(n2865), .Z(n2866) );
  NANDN U3182 ( .A(n60956), .B(n2866), .Z(n2867) );
  ANDN U3183 ( .B(n50543), .A(n50544), .Z(n2868) );
  NAND U3184 ( .A(n2867), .B(n2868), .Z(n2869) );
  NAND U3185 ( .A(n60957), .B(n2869), .Z(n2870) );
  ANDN U3186 ( .B(n60959), .A(n60958), .Z(n2871) );
  NAND U3187 ( .A(n2870), .B(n2871), .Z(n2872) );
  NAND U3188 ( .A(n60960), .B(n2872), .Z(n2873) );
  ANDN U3189 ( .B(n50542), .A(n50541), .Z(n2874) );
  NAND U3190 ( .A(n2873), .B(n2874), .Z(n2875) );
  NAND U3191 ( .A(n50540), .B(n2875), .Z(n2876) );
  ANDN U3192 ( .B(n60962), .A(n60961), .Z(n2877) );
  NAND U3193 ( .A(n2876), .B(n2877), .Z(n2878) );
  NAND U3194 ( .A(n60963), .B(n2878), .Z(n60964) );
  NANDN U3195 ( .A(n60994), .B(n60993), .Z(n2879) );
  NANDN U3196 ( .A(n60995), .B(n2879), .Z(n2880) );
  NANDN U3197 ( .A(n60996), .B(n2880), .Z(n2881) );
  NANDN U3198 ( .A(n2881), .B(n60997), .Z(n2882) );
  AND U3199 ( .A(n60998), .B(n2882), .Z(n2883) );
  NOR U3200 ( .A(n2883), .B(n50528), .Z(n2884) );
  NAND U3201 ( .A(n50529), .B(n2884), .Z(n2885) );
  NANDN U3202 ( .A(n50527), .B(n2885), .Z(n2886) );
  NAND U3203 ( .A(n60999), .B(n2886), .Z(n2887) );
  NAND U3204 ( .A(n61000), .B(n2887), .Z(n2888) );
  AND U3205 ( .A(n61001), .B(n2888), .Z(n2889) );
  AND U3206 ( .A(n61004), .B(n61003), .Z(n2890) );
  NANDN U3207 ( .A(n2889), .B(n61002), .Z(n2891) );
  AND U3208 ( .A(n2890), .B(n2891), .Z(n2892) );
  NANDN U3209 ( .A(n2892), .B(n50526), .Z(n2893) );
  AND U3210 ( .A(n61005), .B(n2893), .Z(n61007) );
  ANDN U3211 ( .B(n50514), .A(n50515), .Z(n61055) );
  NAND U3212 ( .A(n61083), .B(n50506), .Z(n2894) );
  AND U3213 ( .A(n61085), .B(n2894), .Z(n2895) );
  NAND U3214 ( .A(n2895), .B(n61084), .Z(n2896) );
  NAND U3215 ( .A(n61086), .B(n2896), .Z(n2897) );
  AND U3216 ( .A(n61088), .B(n2897), .Z(n2898) );
  NANDN U3217 ( .A(n61087), .B(n2898), .Z(n2899) );
  ANDN U3218 ( .B(n50504), .A(n50505), .Z(n2900) );
  NANDN U3219 ( .A(n61089), .B(n2899), .Z(n2901) );
  NAND U3220 ( .A(n2900), .B(n2901), .Z(n2902) );
  NAND U3221 ( .A(n61090), .B(n2902), .Z(n2903) );
  AND U3222 ( .A(n61092), .B(n2903), .Z(n2904) );
  NANDN U3223 ( .A(n61091), .B(n2904), .Z(n2905) );
  NAND U3224 ( .A(n61093), .B(n2905), .Z(n2906) );
  AND U3225 ( .A(n50503), .B(n2906), .Z(n2907) );
  NAND U3226 ( .A(n2907), .B(n50502), .Z(n2908) );
  NANDN U3227 ( .A(n61094), .B(n2908), .Z(n61096) );
  NAND U3228 ( .A(n61122), .B(n61121), .Z(n2909) );
  NAND U3229 ( .A(n50491), .B(n2909), .Z(n2910) );
  NAND U3230 ( .A(n61123), .B(n2910), .Z(n2911) );
  ANDN U3231 ( .B(n50490), .A(n50489), .Z(n2912) );
  NANDN U3232 ( .A(n61124), .B(n2911), .Z(n2913) );
  NAND U3233 ( .A(n2912), .B(n2913), .Z(n2914) );
  NAND U3234 ( .A(n61125), .B(n2914), .Z(n2915) );
  AND U3235 ( .A(n50487), .B(n2915), .Z(n2916) );
  NANDN U3236 ( .A(n50488), .B(n2916), .Z(n2917) );
  NAND U3237 ( .A(n61126), .B(n2917), .Z(n2918) );
  AND U3238 ( .A(n61127), .B(n2918), .Z(n2919) );
  NANDN U3239 ( .A(n61128), .B(n2919), .Z(n2920) );
  NAND U3240 ( .A(n61129), .B(n2920), .Z(n2921) );
  AND U3241 ( .A(n50486), .B(n2921), .Z(n2922) );
  NANDN U3242 ( .A(n50485), .B(n2922), .Z(n61130) );
  NAND U3243 ( .A(n61157), .B(n61156), .Z(n2923) );
  ANDN U3244 ( .B(n2923), .A(n61158), .Z(n2924) );
  NOR U3245 ( .A(n50475), .B(n2924), .Z(n2925) );
  NAND U3246 ( .A(n61159), .B(n2925), .Z(n2926) );
  NAND U3247 ( .A(n61160), .B(n2926), .Z(n2927) );
  ANDN U3248 ( .B(n61162), .A(n61161), .Z(n2928) );
  NAND U3249 ( .A(n2927), .B(n2928), .Z(n2929) );
  NAND U3250 ( .A(n61163), .B(n2929), .Z(n2930) );
  AND U3251 ( .A(n50474), .B(n50473), .Z(n2931) );
  NAND U3252 ( .A(n2930), .B(n2931), .Z(n2932) );
  NAND U3253 ( .A(n61164), .B(n2932), .Z(n2933) );
  ANDN U3254 ( .B(n61166), .A(n61165), .Z(n2934) );
  NAND U3255 ( .A(n2933), .B(n2934), .Z(n2935) );
  NAND U3256 ( .A(n61167), .B(n2935), .Z(n2936) );
  AND U3257 ( .A(n61168), .B(n61169), .Z(n2937) );
  NAND U3258 ( .A(n2936), .B(n2937), .Z(n2938) );
  NAND U3259 ( .A(n61170), .B(n2938), .Z(n2939) );
  AND U3260 ( .A(n61171), .B(n2939), .Z(n61173) );
  AND U3261 ( .A(n61261), .B(n61262), .Z(n2940) );
  NANDN U3262 ( .A(n50448), .B(n61260), .Z(n2941) );
  NAND U3263 ( .A(n2940), .B(n2941), .Z(n2942) );
  AND U3264 ( .A(n61264), .B(n61265), .Z(n2943) );
  NANDN U3265 ( .A(n61263), .B(n2942), .Z(n2944) );
  NAND U3266 ( .A(n2943), .B(n2944), .Z(n2945) );
  NAND U3267 ( .A(n61266), .B(n2945), .Z(n2946) );
  AND U3268 ( .A(n61267), .B(n2946), .Z(n2947) );
  NANDN U3269 ( .A(n61268), .B(n2947), .Z(n2948) );
  NAND U3270 ( .A(n61269), .B(n2948), .Z(n2949) );
  AND U3271 ( .A(n50446), .B(n2949), .Z(n2950) );
  NAND U3272 ( .A(n2950), .B(n50447), .Z(n2951) );
  NAND U3273 ( .A(n61270), .B(n2951), .Z(n2952) );
  AND U3274 ( .A(n61271), .B(n2952), .Z(n2953) );
  NANDN U3275 ( .A(n61272), .B(n2953), .Z(n2954) );
  NANDN U3276 ( .A(n61273), .B(n2954), .Z(n61274) );
  AND U3277 ( .A(n53901), .B(n27566), .Z(n2955) );
  AND U3278 ( .A(n33966), .B(n27567), .Z(n2956) );
  NAND U3279 ( .A(n53900), .B(n2956), .Z(n2957) );
  AND U3280 ( .A(n2955), .B(n2957), .Z(n2958) );
  NANDN U3281 ( .A(n2958), .B(n53902), .Z(n2959) );
  ANDN U3282 ( .B(n2959), .A(n33967), .Z(n2960) );
  NOR U3283 ( .A(n53904), .B(n27563), .Z(n2961) );
  NANDN U3284 ( .A(n53903), .B(n2960), .Z(n2962) );
  NAND U3285 ( .A(n2961), .B(n2962), .Z(n2963) );
  AND U3286 ( .A(n33968), .B(n33969), .Z(n2964) );
  NAND U3287 ( .A(n2963), .B(n2964), .Z(n2965) );
  NANDN U3288 ( .A(n33970), .B(n2965), .Z(n2966) );
  AND U3289 ( .A(n27560), .B(n27561), .Z(n2967) );
  OR U3290 ( .A(n2966), .B(n33971), .Z(n2968) );
  AND U3291 ( .A(n2967), .B(n2968), .Z(n2969) );
  NOR U3292 ( .A(n2969), .B(n33972), .Z(n2970) );
  XNOR U3293 ( .A(y[1782]), .B(x[1782]), .Z(n2971) );
  NAND U3294 ( .A(n2970), .B(n2971), .Z(n2972) );
  NANDN U3295 ( .A(n33973), .B(n2972), .Z(n33975) );
  ANDN U3296 ( .B(n28361), .A(n28360), .Z(n52440) );
  NANDN U3297 ( .A(n52461), .B(n52460), .Z(n2973) );
  NANDN U3298 ( .A(n52462), .B(n2973), .Z(n2974) );
  AND U3299 ( .A(n52463), .B(n2974), .Z(n2975) );
  OR U3300 ( .A(n52436), .B(n2975), .Z(n2976) );
  NAND U3301 ( .A(n52464), .B(n2976), .Z(n2977) );
  NANDN U3302 ( .A(n52465), .B(n2977), .Z(n2978) );
  NAND U3303 ( .A(n52466), .B(n2978), .Z(n2979) );
  AND U3304 ( .A(n52435), .B(n2979), .Z(n2980) );
  NANDN U3305 ( .A(n52434), .B(n2980), .Z(n2981) );
  NAND U3306 ( .A(n52467), .B(n2981), .Z(n2982) );
  NANDN U3307 ( .A(n52433), .B(n2982), .Z(n2983) );
  AND U3308 ( .A(n52468), .B(n2983), .Z(n2984) );
  OR U3309 ( .A(n52469), .B(n2984), .Z(n2985) );
  AND U3310 ( .A(n52470), .B(n2985), .Z(n2986) );
  NANDN U3311 ( .A(n2986), .B(n52471), .Z(n2987) );
  NANDN U3312 ( .A(n52472), .B(n2987), .Z(n2988) );
  NANDN U3313 ( .A(n52473), .B(n2988), .Z(n52474) );
  NAND U3314 ( .A(n52509), .B(n52510), .Z(n2989) );
  NAND U3315 ( .A(n52511), .B(n2989), .Z(n2990) );
  ANDN U3316 ( .B(n2990), .A(n52512), .Z(n2991) );
  OR U3317 ( .A(n52513), .B(n2991), .Z(n2992) );
  NAND U3318 ( .A(n52514), .B(n2992), .Z(n2993) );
  NANDN U3319 ( .A(n52429), .B(n2993), .Z(n2994) );
  NAND U3320 ( .A(n52515), .B(n2994), .Z(n2995) );
  NANDN U3321 ( .A(n52516), .B(n2995), .Z(n2996) );
  AND U3322 ( .A(n52517), .B(n2996), .Z(n2997) );
  NANDN U3323 ( .A(n2997), .B(n52518), .Z(n2998) );
  NAND U3324 ( .A(n52519), .B(n2998), .Z(n2999) );
  NANDN U3325 ( .A(n52520), .B(n2999), .Z(n3000) );
  NAND U3326 ( .A(n52521), .B(n3000), .Z(n3001) );
  NANDN U3327 ( .A(n52522), .B(n3001), .Z(n3002) );
  AND U3328 ( .A(n52523), .B(n3002), .Z(n3003) );
  OR U3329 ( .A(n52524), .B(n3003), .Z(n3004) );
  NAND U3330 ( .A(n52525), .B(n3004), .Z(n3005) );
  NAND U3331 ( .A(n52526), .B(n3005), .Z(n52527) );
  NANDN U3332 ( .A(n52421), .B(n52593), .Z(n3006) );
  NAND U3333 ( .A(n52420), .B(n3006), .Z(n3007) );
  NANDN U3334 ( .A(n52594), .B(n3007), .Z(n3008) );
  NAND U3335 ( .A(n52595), .B(n3008), .Z(n3009) );
  NANDN U3336 ( .A(n52419), .B(n3009), .Z(n3010) );
  AND U3337 ( .A(n52418), .B(n3010), .Z(n3011) );
  NANDN U3338 ( .A(n3011), .B(n52596), .Z(n3012) );
  AND U3339 ( .A(n52417), .B(n3012), .Z(n3013) );
  NANDN U3340 ( .A(n3013), .B(n52597), .Z(n3014) );
  NAND U3341 ( .A(n52598), .B(n3014), .Z(n3015) );
  NANDN U3342 ( .A(n52416), .B(n3015), .Z(n52599) );
  OR U3343 ( .A(n52651), .B(n52650), .Z(n3016) );
  NAND U3344 ( .A(n52652), .B(n3016), .Z(n3017) );
  ANDN U3345 ( .B(n3017), .A(n52653), .Z(n3018) );
  NANDN U3346 ( .A(n3018), .B(n52654), .Z(n3019) );
  NANDN U3347 ( .A(n52655), .B(n3019), .Z(n3020) );
  NAND U3348 ( .A(n52656), .B(n3020), .Z(n3021) );
  NANDN U3349 ( .A(n52657), .B(n3021), .Z(n3022) );
  NAND U3350 ( .A(n52658), .B(n3022), .Z(n3023) );
  AND U3351 ( .A(n52659), .B(n3023), .Z(n3024) );
  NANDN U3352 ( .A(n3024), .B(n52660), .Z(n3025) );
  NANDN U3353 ( .A(n52661), .B(n3025), .Z(n3026) );
  NAND U3354 ( .A(n52662), .B(n3026), .Z(n3027) );
  NANDN U3355 ( .A(n52663), .B(n3027), .Z(n3028) );
  NAND U3356 ( .A(n52664), .B(n3028), .Z(n3029) );
  ANDN U3357 ( .B(n3029), .A(n52665), .Z(n3030) );
  NANDN U3358 ( .A(n3030), .B(n52666), .Z(n3031) );
  NANDN U3359 ( .A(n52667), .B(n3031), .Z(n3032) );
  NANDN U3360 ( .A(n52668), .B(n3032), .Z(n3033) );
  NAND U3361 ( .A(n52669), .B(n3033), .Z(n52670) );
  NAND U3362 ( .A(n52744), .B(n52743), .Z(n3034) );
  NAND U3363 ( .A(n52406), .B(n3034), .Z(n3035) );
  ANDN U3364 ( .B(n3035), .A(n52745), .Z(n3036) );
  NANDN U3365 ( .A(n3036), .B(n52405), .Z(n3037) );
  NAND U3366 ( .A(n52746), .B(n3037), .Z(n3038) );
  NAND U3367 ( .A(n52747), .B(n3038), .Z(n3039) );
  NANDN U3368 ( .A(n52404), .B(n3039), .Z(n3040) );
  NAND U3369 ( .A(n52403), .B(n3040), .Z(n3041) );
  ANDN U3370 ( .B(n3041), .A(n52402), .Z(n3042) );
  NANDN U3371 ( .A(n3042), .B(n52401), .Z(n3043) );
  NAND U3372 ( .A(n52748), .B(n3043), .Z(n3044) );
  NAND U3373 ( .A(n52749), .B(n3044), .Z(n3045) );
  NANDN U3374 ( .A(n52750), .B(n3045), .Z(n52751) );
  NAND U3375 ( .A(n52868), .B(n52869), .Z(n3046) );
  NAND U3376 ( .A(n52388), .B(n3046), .Z(n3047) );
  NANDN U3377 ( .A(n52870), .B(n3047), .Z(n3048) );
  NAND U3378 ( .A(n52871), .B(n3048), .Z(n3049) );
  NANDN U3379 ( .A(n52387), .B(n3049), .Z(n3050) );
  AND U3380 ( .A(n52386), .B(n3050), .Z(n3051) );
  OR U3381 ( .A(n52385), .B(n3051), .Z(n3052) );
  AND U3382 ( .A(n52384), .B(n3052), .Z(n3053) );
  NANDN U3383 ( .A(n3053), .B(n52872), .Z(n3054) );
  NAND U3384 ( .A(n52873), .B(n3054), .Z(n3055) );
  NANDN U3385 ( .A(n52383), .B(n3055), .Z(n52874) );
  NANDN U3386 ( .A(n52893), .B(n52892), .Z(n3056) );
  NANDN U3387 ( .A(n52894), .B(n3056), .Z(n3057) );
  AND U3388 ( .A(n52895), .B(n3057), .Z(n3058) );
  OR U3389 ( .A(n52370), .B(n3058), .Z(n3059) );
  NAND U3390 ( .A(n52896), .B(n3059), .Z(n3060) );
  NANDN U3391 ( .A(n52369), .B(n3060), .Z(n3061) );
  NAND U3392 ( .A(n52897), .B(n3061), .Z(n3062) );
  NANDN U3393 ( .A(n52898), .B(n3062), .Z(n3063) );
  AND U3394 ( .A(n52899), .B(n3063), .Z(n3064) );
  OR U3395 ( .A(n52368), .B(n3064), .Z(n3065) );
  NAND U3396 ( .A(n52900), .B(n3065), .Z(n3066) );
  NANDN U3397 ( .A(n52367), .B(n3066), .Z(n3067) );
  NAND U3398 ( .A(n52366), .B(n3067), .Z(n52903) );
  NAND U3399 ( .A(n52930), .B(n52929), .Z(n3068) );
  NANDN U3400 ( .A(n52931), .B(n3068), .Z(n3069) );
  NANDN U3401 ( .A(n52360), .B(n3069), .Z(n3070) );
  NAND U3402 ( .A(n52932), .B(n3070), .Z(n3071) );
  NAND U3403 ( .A(n52933), .B(n3071), .Z(n3072) );
  AND U3404 ( .A(n52934), .B(n3072), .Z(n3073) );
  NANDN U3405 ( .A(n3073), .B(n52935), .Z(n3074) );
  NAND U3406 ( .A(n52359), .B(n3074), .Z(n3075) );
  NANDN U3407 ( .A(n52358), .B(n3075), .Z(n3076) );
  NANDN U3408 ( .A(n52936), .B(n3076), .Z(n3077) );
  NAND U3409 ( .A(n52937), .B(n3077), .Z(n3078) );
  ANDN U3410 ( .B(n3078), .A(n52938), .Z(n3079) );
  NANDN U3411 ( .A(n3079), .B(n52939), .Z(n3080) );
  NANDN U3412 ( .A(n52940), .B(n3080), .Z(n3081) );
  NAND U3413 ( .A(n52941), .B(n3081), .Z(n3082) );
  NANDN U3414 ( .A(n52942), .B(n3082), .Z(n52944) );
  NAND U3415 ( .A(n52979), .B(n52980), .Z(n3083) );
  NAND U3416 ( .A(n52981), .B(n3083), .Z(n3084) );
  AND U3417 ( .A(n52982), .B(n3084), .Z(n3085) );
  OR U3418 ( .A(n52983), .B(n3085), .Z(n3086) );
  NAND U3419 ( .A(n52984), .B(n3086), .Z(n3087) );
  NANDN U3420 ( .A(n52985), .B(n3087), .Z(n3088) );
  NAND U3421 ( .A(n52986), .B(n3088), .Z(n3089) );
  NANDN U3422 ( .A(n52987), .B(n3089), .Z(n3090) );
  AND U3423 ( .A(n52988), .B(n3090), .Z(n3091) );
  OR U3424 ( .A(n52989), .B(n3091), .Z(n3092) );
  NANDN U3425 ( .A(n52990), .B(n3092), .Z(n3093) );
  NAND U3426 ( .A(n52991), .B(n3093), .Z(n3094) );
  NAND U3427 ( .A(n52992), .B(n3094), .Z(n3095) );
  NAND U3428 ( .A(n52993), .B(n3095), .Z(n3096) );
  AND U3429 ( .A(n52994), .B(n3096), .Z(n3097) );
  OR U3430 ( .A(n52995), .B(n3097), .Z(n3098) );
  NAND U3431 ( .A(n52996), .B(n3098), .Z(n3099) );
  NANDN U3432 ( .A(n52997), .B(n3099), .Z(n3100) );
  NAND U3433 ( .A(n52998), .B(n3100), .Z(n52999) );
  NANDN U3434 ( .A(n53035), .B(n53034), .Z(n3101) );
  NANDN U3435 ( .A(n53036), .B(n3101), .Z(n3102) );
  NAND U3436 ( .A(n53037), .B(n3102), .Z(n3103) );
  NANDN U3437 ( .A(n53038), .B(n3103), .Z(n3104) );
  NAND U3438 ( .A(n53039), .B(n3104), .Z(n3105) );
  ANDN U3439 ( .B(n3105), .A(n53040), .Z(n3106) );
  OR U3440 ( .A(n3106), .B(n53041), .Z(n3107) );
  NAND U3441 ( .A(n53042), .B(n3107), .Z(n3108) );
  ANDN U3442 ( .B(n3108), .A(n53043), .Z(n3109) );
  NANDN U3443 ( .A(n3109), .B(n53044), .Z(n3110) );
  NANDN U3444 ( .A(n53045), .B(n3110), .Z(n3111) );
  NAND U3445 ( .A(n53046), .B(n3111), .Z(n3112) );
  NANDN U3446 ( .A(n53047), .B(n3112), .Z(n3113) );
  NANDN U3447 ( .A(n53048), .B(n3113), .Z(n3114) );
  AND U3448 ( .A(n53049), .B(n3114), .Z(n3115) );
  OR U3449 ( .A(n3115), .B(n53050), .Z(n3116) );
  NAND U3450 ( .A(n53051), .B(n3116), .Z(n3117) );
  NAND U3451 ( .A(n53052), .B(n3117), .Z(n3118) );
  NANDN U3452 ( .A(n53053), .B(n3118), .Z(n53054) );
  OR U3453 ( .A(n53084), .B(n53085), .Z(n3119) );
  NANDN U3454 ( .A(n53086), .B(n3119), .Z(n3120) );
  ANDN U3455 ( .B(n3120), .A(n53087), .Z(n3121) );
  NANDN U3456 ( .A(n3121), .B(n53088), .Z(n3122) );
  NANDN U3457 ( .A(n53089), .B(n3122), .Z(n3123) );
  NAND U3458 ( .A(n53090), .B(n3123), .Z(n3124) );
  NANDN U3459 ( .A(n53091), .B(n3124), .Z(n3125) );
  NAND U3460 ( .A(n53092), .B(n3125), .Z(n3126) );
  ANDN U3461 ( .B(n3126), .A(n53093), .Z(n3127) );
  OR U3462 ( .A(n53094), .B(n3127), .Z(n3128) );
  NAND U3463 ( .A(n53095), .B(n3128), .Z(n3129) );
  NANDN U3464 ( .A(n53096), .B(n3129), .Z(n3130) );
  NAND U3465 ( .A(n53097), .B(n3130), .Z(n3131) );
  NANDN U3466 ( .A(n53098), .B(n3131), .Z(n3132) );
  AND U3467 ( .A(n53099), .B(n3132), .Z(n3133) );
  OR U3468 ( .A(n53100), .B(n3133), .Z(n3134) );
  NAND U3469 ( .A(n53101), .B(n3134), .Z(n3135) );
  NANDN U3470 ( .A(n53102), .B(n3135), .Z(n53103) );
  NAND U3471 ( .A(n53162), .B(n53161), .Z(n3136) );
  NAND U3472 ( .A(n52344), .B(n3136), .Z(n3137) );
  ANDN U3473 ( .B(n3137), .A(n52343), .Z(n3138) );
  NANDN U3474 ( .A(n3138), .B(n52342), .Z(n3139) );
  NANDN U3475 ( .A(n53163), .B(n3139), .Z(n3140) );
  NAND U3476 ( .A(n53164), .B(n3140), .Z(n3141) );
  NAND U3477 ( .A(n53165), .B(n3141), .Z(n3142) );
  NAND U3478 ( .A(n53166), .B(n3142), .Z(n3143) );
  AND U3479 ( .A(n53167), .B(n3143), .Z(n3144) );
  NANDN U3480 ( .A(n3144), .B(n53168), .Z(n3145) );
  NANDN U3481 ( .A(n52341), .B(n3145), .Z(n3146) );
  NAND U3482 ( .A(n52340), .B(n3146), .Z(n53171) );
  NANDN U3483 ( .A(n53190), .B(n53189), .Z(n3147) );
  NAND U3484 ( .A(n53191), .B(n3147), .Z(n3148) );
  ANDN U3485 ( .B(n3148), .A(n53192), .Z(n3149) );
  NANDN U3486 ( .A(n3149), .B(n53193), .Z(n3150) );
  NANDN U3487 ( .A(n53194), .B(n3150), .Z(n3151) );
  NAND U3488 ( .A(n53195), .B(n3151), .Z(n3152) );
  NANDN U3489 ( .A(n53196), .B(n3152), .Z(n3153) );
  NAND U3490 ( .A(n53197), .B(n3153), .Z(n3154) );
  ANDN U3491 ( .B(n3154), .A(n53198), .Z(n3155) );
  NANDN U3492 ( .A(n3155), .B(n53199), .Z(n3156) );
  NANDN U3493 ( .A(n53200), .B(n3156), .Z(n3157) );
  NANDN U3494 ( .A(n52329), .B(n3157), .Z(n3158) );
  NAND U3495 ( .A(n53201), .B(n3158), .Z(n3159) );
  NAND U3496 ( .A(n53202), .B(n3159), .Z(n3160) );
  ANDN U3497 ( .B(n3160), .A(n53203), .Z(n3161) );
  NANDN U3498 ( .A(n3161), .B(n53204), .Z(n3162) );
  NANDN U3499 ( .A(n53205), .B(n3162), .Z(n3163) );
  NAND U3500 ( .A(n53206), .B(n3163), .Z(n3164) );
  NANDN U3501 ( .A(n53207), .B(n3164), .Z(n53208) );
  NAND U3502 ( .A(n53239), .B(n53240), .Z(n3165) );
  NANDN U3503 ( .A(n53241), .B(n3165), .Z(n3166) );
  NAND U3504 ( .A(n53242), .B(n3166), .Z(n3167) );
  NANDN U3505 ( .A(n52322), .B(n3167), .Z(n3168) );
  NAND U3506 ( .A(n52321), .B(n3168), .Z(n3169) );
  AND U3507 ( .A(n53243), .B(n3169), .Z(n3170) );
  NANDN U3508 ( .A(n52320), .B(n3170), .Z(n3171) );
  NANDN U3509 ( .A(n53244), .B(n3171), .Z(n3172) );
  ANDN U3510 ( .B(n3172), .A(n53245), .Z(n3173) );
  NANDN U3511 ( .A(n53246), .B(n3173), .Z(n3174) );
  NANDN U3512 ( .A(n53247), .B(n3174), .Z(n3175) );
  AND U3513 ( .A(n53248), .B(n3175), .Z(n3176) );
  NANDN U3514 ( .A(n3176), .B(n53249), .Z(n3177) );
  NANDN U3515 ( .A(n53250), .B(n3177), .Z(n3178) );
  NAND U3516 ( .A(n53251), .B(n3178), .Z(n53252) );
  NAND U3517 ( .A(n53283), .B(n53282), .Z(n3179) );
  NANDN U3518 ( .A(n53284), .B(n3179), .Z(n3180) );
  NAND U3519 ( .A(n53285), .B(n3180), .Z(n3181) );
  NAND U3520 ( .A(n53286), .B(n3181), .Z(n3182) );
  NANDN U3521 ( .A(n53287), .B(n3182), .Z(n3183) );
  AND U3522 ( .A(n53288), .B(n3183), .Z(n3184) );
  OR U3523 ( .A(n3184), .B(n53289), .Z(n3185) );
  NAND U3524 ( .A(n53290), .B(n3185), .Z(n3186) );
  NAND U3525 ( .A(n53291), .B(n3186), .Z(n3187) );
  NAND U3526 ( .A(n53292), .B(n3187), .Z(n3188) );
  NAND U3527 ( .A(n53293), .B(n3188), .Z(n3189) );
  AND U3528 ( .A(n53294), .B(n3189), .Z(n3190) );
  NANDN U3529 ( .A(n3190), .B(n53295), .Z(n3191) );
  NANDN U3530 ( .A(n53296), .B(n3191), .Z(n3192) );
  NANDN U3531 ( .A(n53297), .B(n3192), .Z(n3193) );
  NAND U3532 ( .A(n53298), .B(n3193), .Z(n3194) );
  NANDN U3533 ( .A(n53299), .B(n3194), .Z(n3195) );
  AND U3534 ( .A(n53300), .B(n3195), .Z(n53302) );
  NANDN U3535 ( .A(n53336), .B(n53335), .Z(n3196) );
  NAND U3536 ( .A(n53337), .B(n3196), .Z(n3197) );
  NANDN U3537 ( .A(n53338), .B(n3197), .Z(n3198) );
  NAND U3538 ( .A(n53339), .B(n3198), .Z(n3199) );
  NANDN U3539 ( .A(n53340), .B(n3199), .Z(n3200) );
  AND U3540 ( .A(n53341), .B(n3200), .Z(n3201) );
  OR U3541 ( .A(n53342), .B(n3201), .Z(n3202) );
  NAND U3542 ( .A(n53343), .B(n3202), .Z(n3203) );
  NANDN U3543 ( .A(n53344), .B(n3203), .Z(n3204) );
  NAND U3544 ( .A(n53345), .B(n3204), .Z(n3205) );
  NAND U3545 ( .A(n53346), .B(n3205), .Z(n3206) );
  ANDN U3546 ( .B(n3206), .A(n52310), .Z(n3207) );
  OR U3547 ( .A(n53347), .B(n3207), .Z(n3208) );
  NAND U3548 ( .A(n53348), .B(n3208), .Z(n3209) );
  NANDN U3549 ( .A(n52309), .B(n3209), .Z(n3210) );
  NAND U3550 ( .A(n52308), .B(n3210), .Z(n53349) );
  NAND U3551 ( .A(n53403), .B(n53404), .Z(n3211) );
  NANDN U3552 ( .A(n53405), .B(n3211), .Z(n3212) );
  AND U3553 ( .A(n53406), .B(n3212), .Z(n3213) );
  NANDN U3554 ( .A(n3213), .B(n53407), .Z(n3214) );
  ANDN U3555 ( .B(n3214), .A(n52303), .Z(n3215) );
  OR U3556 ( .A(n53408), .B(n3215), .Z(n3216) );
  NANDN U3557 ( .A(n53409), .B(n3216), .Z(n3217) );
  NANDN U3558 ( .A(n53410), .B(n3217), .Z(n3218) );
  NAND U3559 ( .A(n53412), .B(n53411), .Z(n3219) );
  NANDN U3560 ( .A(n3218), .B(n3219), .Z(n3220) );
  AND U3561 ( .A(n53413), .B(n3220), .Z(n3221) );
  OR U3562 ( .A(n52302), .B(n3221), .Z(n3222) );
  AND U3563 ( .A(n53414), .B(n3222), .Z(n3223) );
  OR U3564 ( .A(n53415), .B(n3223), .Z(n3224) );
  NAND U3565 ( .A(n53416), .B(n3224), .Z(n3225) );
  NANDN U3566 ( .A(n53417), .B(n3225), .Z(n53418) );
  NAND U3567 ( .A(n53450), .B(n53451), .Z(n3226) );
  NAND U3568 ( .A(n53452), .B(n3226), .Z(n3227) );
  NANDN U3569 ( .A(n52285), .B(n3227), .Z(n3228) );
  NAND U3570 ( .A(n52284), .B(n3228), .Z(n3229) );
  NAND U3571 ( .A(n53453), .B(n3229), .Z(n3230) );
  AND U3572 ( .A(n53454), .B(n3230), .Z(n3231) );
  NANDN U3573 ( .A(n3231), .B(n53455), .Z(n3232) );
  NAND U3574 ( .A(n53456), .B(n3232), .Z(n3233) );
  NAND U3575 ( .A(n53457), .B(n3233), .Z(n3234) );
  NANDN U3576 ( .A(n53458), .B(n3234), .Z(n3235) );
  NAND U3577 ( .A(n53459), .B(n3235), .Z(n3236) );
  ANDN U3578 ( .B(n3236), .A(n53460), .Z(n3237) );
  NANDN U3579 ( .A(n3237), .B(n53461), .Z(n3238) );
  NANDN U3580 ( .A(n53462), .B(n3238), .Z(n3239) );
  NANDN U3581 ( .A(n52283), .B(n3239), .Z(n53463) );
  NAND U3582 ( .A(n52279), .B(n53496), .Z(n3240) );
  NAND U3583 ( .A(n53497), .B(n3240), .Z(n3241) );
  NAND U3584 ( .A(n53498), .B(n3241), .Z(n3242) );
  NANDN U3585 ( .A(n52278), .B(n3242), .Z(n3243) );
  NAND U3586 ( .A(n53499), .B(n3243), .Z(n3244) );
  ANDN U3587 ( .B(n3244), .A(n53500), .Z(n3245) );
  NANDN U3588 ( .A(n3245), .B(n53501), .Z(n3246) );
  NAND U3589 ( .A(n53502), .B(n3246), .Z(n3247) );
  NANDN U3590 ( .A(n53503), .B(n3247), .Z(n3248) );
  NAND U3591 ( .A(n53504), .B(n3248), .Z(n3249) );
  NAND U3592 ( .A(n53505), .B(n3249), .Z(n3250) );
  AND U3593 ( .A(n53506), .B(n3250), .Z(n3251) );
  NANDN U3594 ( .A(n3251), .B(n53507), .Z(n3252) );
  NAND U3595 ( .A(n53508), .B(n3252), .Z(n3253) );
  NANDN U3596 ( .A(n52277), .B(n3253), .Z(n53509) );
  NAND U3597 ( .A(n53529), .B(n53530), .Z(n3254) );
  NANDN U3598 ( .A(n53531), .B(n3254), .Z(n3255) );
  AND U3599 ( .A(n53532), .B(n3255), .Z(n3256) );
  NANDN U3600 ( .A(n3256), .B(n53533), .Z(n3257) );
  NAND U3601 ( .A(n53534), .B(n3257), .Z(n3258) );
  NANDN U3602 ( .A(n52267), .B(n3258), .Z(n3259) );
  NANDN U3603 ( .A(n53535), .B(n3259), .Z(n3260) );
  NAND U3604 ( .A(n53536), .B(n3260), .Z(n3261) );
  ANDN U3605 ( .B(n3261), .A(n53537), .Z(n3262) );
  NANDN U3606 ( .A(n3262), .B(n53538), .Z(n3263) );
  NANDN U3607 ( .A(n53539), .B(n3263), .Z(n3264) );
  NAND U3608 ( .A(n53540), .B(n3264), .Z(n3265) );
  NANDN U3609 ( .A(n53541), .B(n3265), .Z(n3266) );
  NAND U3610 ( .A(n53542), .B(n3266), .Z(n3267) );
  ANDN U3611 ( .B(n3267), .A(n53543), .Z(n3268) );
  NANDN U3612 ( .A(n3268), .B(n53544), .Z(n3269) );
  NANDN U3613 ( .A(n53545), .B(n3269), .Z(n3270) );
  NAND U3614 ( .A(n53546), .B(n3270), .Z(n3271) );
  NANDN U3615 ( .A(n53547), .B(n3271), .Z(n53548) );
  NANDN U3616 ( .A(n53579), .B(n53578), .Z(n3272) );
  NANDN U3617 ( .A(n53580), .B(n3272), .Z(n3273) );
  NAND U3618 ( .A(n53581), .B(n3273), .Z(n3274) );
  NANDN U3619 ( .A(n52261), .B(n3274), .Z(n3275) );
  NAND U3620 ( .A(n52260), .B(n3275), .Z(n3276) );
  ANDN U3621 ( .B(n3276), .A(n53582), .Z(n3277) );
  NANDN U3622 ( .A(n3277), .B(n53583), .Z(n3278) );
  NANDN U3623 ( .A(n53584), .B(n3278), .Z(n3279) );
  NANDN U3624 ( .A(n53585), .B(n3279), .Z(n3280) );
  NAND U3625 ( .A(n53586), .B(n3280), .Z(n3281) );
  NANDN U3626 ( .A(n52259), .B(n3281), .Z(n3282) );
  AND U3627 ( .A(n53587), .B(n3282), .Z(n3283) );
  OR U3628 ( .A(n53588), .B(n3283), .Z(n3284) );
  NAND U3629 ( .A(n53589), .B(n3284), .Z(n3285) );
  NANDN U3630 ( .A(n53590), .B(n3285), .Z(n53591) );
  NANDN U3631 ( .A(n53624), .B(n53623), .Z(n3286) );
  NAND U3632 ( .A(n52254), .B(n3286), .Z(n3287) );
  ANDN U3633 ( .B(n3287), .A(n53625), .Z(n3288) );
  NANDN U3634 ( .A(n3288), .B(n53626), .Z(n3289) );
  NANDN U3635 ( .A(n52253), .B(n3289), .Z(n3290) );
  NAND U3636 ( .A(n52252), .B(n3290), .Z(n3291) );
  NAND U3637 ( .A(n53627), .B(n3291), .Z(n3292) );
  NAND U3638 ( .A(n53628), .B(n3292), .Z(n3293) );
  AND U3639 ( .A(n53629), .B(n3293), .Z(n3294) );
  OR U3640 ( .A(n53630), .B(n3294), .Z(n3295) );
  AND U3641 ( .A(n53631), .B(n3295), .Z(n3296) );
  ANDN U3642 ( .B(n52251), .A(n3296), .Z(n3297) );
  NAND U3643 ( .A(n52250), .B(n3297), .Z(n3298) );
  AND U3644 ( .A(n53632), .B(n3298), .Z(n3299) );
  NANDN U3645 ( .A(n53633), .B(n3299), .Z(n53634) );
  ANDN U3646 ( .B(n27701), .A(n27700), .Z(n53702) );
  NANDN U3647 ( .A(n53730), .B(n53729), .Z(n3300) );
  NAND U3648 ( .A(n53731), .B(n3300), .Z(n3301) );
  NANDN U3649 ( .A(n53732), .B(n3301), .Z(n3302) );
  NAND U3650 ( .A(n53733), .B(n3302), .Z(n3303) );
  NANDN U3651 ( .A(n53734), .B(n3303), .Z(n3304) );
  AND U3652 ( .A(n53735), .B(n3304), .Z(n3305) );
  NANDN U3653 ( .A(n3305), .B(n53736), .Z(n3306) );
  NANDN U3654 ( .A(n53737), .B(n3306), .Z(n3307) );
  NAND U3655 ( .A(n53738), .B(n3307), .Z(n3308) );
  OR U3656 ( .A(n53739), .B(n53740), .Z(n3309) );
  NANDN U3657 ( .A(n3308), .B(n3309), .Z(n3310) );
  AND U3658 ( .A(n53741), .B(n3310), .Z(n3311) );
  OR U3659 ( .A(n52245), .B(n3311), .Z(n3312) );
  NAND U3660 ( .A(n53742), .B(n3312), .Z(n3313) );
  NANDN U3661 ( .A(n52244), .B(n3313), .Z(n3314) );
  NAND U3662 ( .A(n52243), .B(n3314), .Z(n53744) );
  NAND U3663 ( .A(n53807), .B(n53808), .Z(n3315) );
  NANDN U3664 ( .A(n53809), .B(n3315), .Z(n3316) );
  NAND U3665 ( .A(n53810), .B(n3316), .Z(n3317) );
  NANDN U3666 ( .A(n53811), .B(n3317), .Z(n3318) );
  NAND U3667 ( .A(n53812), .B(n3318), .Z(n3319) );
  ANDN U3668 ( .B(n3319), .A(n53813), .Z(n3320) );
  NANDN U3669 ( .A(n3320), .B(n53814), .Z(n3321) );
  AND U3670 ( .A(n53815), .B(n3321), .Z(n3322) );
  NAND U3671 ( .A(n52233), .B(n52232), .Z(n3323) );
  AND U3672 ( .A(n52234), .B(n3323), .Z(n3324) );
  NANDN U3673 ( .A(n3322), .B(n3324), .Z(n3325) );
  NAND U3674 ( .A(n53816), .B(n3325), .Z(n3326) );
  NAND U3675 ( .A(n53817), .B(n3326), .Z(n3327) );
  ANDN U3676 ( .B(n3327), .A(n53818), .Z(n3328) );
  NANDN U3677 ( .A(n3328), .B(n53819), .Z(n3329) );
  NAND U3678 ( .A(n53820), .B(n3329), .Z(n3330) );
  NAND U3679 ( .A(n53821), .B(n3330), .Z(n3331) );
  NAND U3680 ( .A(n53822), .B(n3331), .Z(n53823) );
  NAND U3681 ( .A(n53842), .B(n53841), .Z(n3332) );
  NAND U3682 ( .A(n53843), .B(n3332), .Z(n3333) );
  NANDN U3683 ( .A(n53844), .B(n3333), .Z(n3334) );
  NAND U3684 ( .A(n53845), .B(n3334), .Z(n3335) );
  NANDN U3685 ( .A(n53846), .B(n3335), .Z(n3336) );
  AND U3686 ( .A(n53847), .B(n3336), .Z(n3337) );
  OR U3687 ( .A(n53848), .B(n3337), .Z(n3338) );
  ANDN U3688 ( .B(n3338), .A(n53849), .Z(n3339) );
  NOR U3689 ( .A(n53850), .B(n3339), .Z(n3340) );
  NAND U3690 ( .A(n53851), .B(n3340), .Z(n3341) );
  ANDN U3691 ( .B(n3341), .A(n53852), .Z(n3342) );
  NANDN U3692 ( .A(n3342), .B(n53853), .Z(n3343) );
  ANDN U3693 ( .B(n3343), .A(n53854), .Z(n3344) );
  NANDN U3694 ( .A(n3344), .B(n53855), .Z(n3345) );
  NANDN U3695 ( .A(n53856), .B(n3345), .Z(n3346) );
  NANDN U3696 ( .A(n53857), .B(n3346), .Z(n53858) );
  NAND U3697 ( .A(n53882), .B(n53883), .Z(n3347) );
  NANDN U3698 ( .A(n53884), .B(n3347), .Z(n3348) );
  ANDN U3699 ( .B(n3348), .A(n53885), .Z(n3349) );
  NANDN U3700 ( .A(n3349), .B(n53886), .Z(n3350) );
  ANDN U3701 ( .B(n3350), .A(n53887), .Z(n3351) );
  NANDN U3702 ( .A(n3351), .B(n53888), .Z(n3352) );
  NANDN U3703 ( .A(n53889), .B(n3352), .Z(n3353) );
  NAND U3704 ( .A(n53890), .B(n3353), .Z(n3354) );
  AND U3705 ( .A(n52211), .B(n52212), .Z(n3355) );
  NAND U3706 ( .A(n3354), .B(n3355), .Z(n3356) );
  NANDN U3707 ( .A(n53891), .B(n3356), .Z(n3357) );
  NAND U3708 ( .A(n53892), .B(n3357), .Z(n3358) );
  NANDN U3709 ( .A(n53893), .B(n3358), .Z(n3359) );
  AND U3710 ( .A(n52210), .B(n3359), .Z(n3360) );
  NANDN U3711 ( .A(n3360), .B(n53894), .Z(n3361) );
  NAND U3712 ( .A(n53895), .B(n3361), .Z(n3362) );
  NANDN U3713 ( .A(n52209), .B(n3362), .Z(n53896) );
  AND U3714 ( .A(n53926), .B(n52203), .Z(n3363) );
  NAND U3715 ( .A(n53927), .B(n3363), .Z(n3364) );
  NAND U3716 ( .A(n53928), .B(n3364), .Z(n3365) );
  NANDN U3717 ( .A(n53929), .B(n3365), .Z(n3366) );
  NAND U3718 ( .A(n53930), .B(n3366), .Z(n3367) );
  AND U3719 ( .A(n53931), .B(n3367), .Z(n3368) );
  OR U3720 ( .A(n53932), .B(n3368), .Z(n3369) );
  NANDN U3721 ( .A(n53933), .B(n3369), .Z(n3370) );
  NAND U3722 ( .A(n53934), .B(n3370), .Z(n3371) );
  NANDN U3723 ( .A(n53935), .B(n3371), .Z(n3372) );
  NAND U3724 ( .A(n53936), .B(n3372), .Z(n3373) );
  ANDN U3725 ( .B(n3373), .A(n53937), .Z(n3374) );
  NANDN U3726 ( .A(n3374), .B(n53938), .Z(n3375) );
  AND U3727 ( .A(n53939), .B(n3375), .Z(n3376) );
  NANDN U3728 ( .A(n3376), .B(n53940), .Z(n3377) );
  NANDN U3729 ( .A(n53941), .B(n3377), .Z(n3378) );
  NAND U3730 ( .A(n53942), .B(n3378), .Z(n53943) );
  NAND U3731 ( .A(n53976), .B(n53975), .Z(n3379) );
  NANDN U3732 ( .A(n53977), .B(n3379), .Z(n3380) );
  ANDN U3733 ( .B(n3380), .A(n53978), .Z(n3381) );
  OR U3734 ( .A(n3381), .B(n53979), .Z(n3382) );
  NAND U3735 ( .A(n53980), .B(n3382), .Z(n3383) );
  ANDN U3736 ( .B(n3383), .A(n53981), .Z(n3384) );
  NANDN U3737 ( .A(n3384), .B(n53982), .Z(n3385) );
  NANDN U3738 ( .A(n53983), .B(n3385), .Z(n3386) );
  NAND U3739 ( .A(n53984), .B(n3386), .Z(n3387) );
  NANDN U3740 ( .A(n53985), .B(n3387), .Z(n3388) );
  NANDN U3741 ( .A(n53986), .B(n3388), .Z(n3389) );
  AND U3742 ( .A(n53987), .B(n3389), .Z(n3390) );
  OR U3743 ( .A(n52198), .B(n3390), .Z(n3391) );
  NAND U3744 ( .A(n53988), .B(n3391), .Z(n3392) );
  NANDN U3745 ( .A(n53989), .B(n3392), .Z(n3393) );
  NAND U3746 ( .A(n53990), .B(n3393), .Z(n3394) );
  NANDN U3747 ( .A(n53991), .B(n3394), .Z(n3395) );
  AND U3748 ( .A(n53992), .B(n3395), .Z(n53993) );
  NAND U3749 ( .A(n54021), .B(n52191), .Z(n3396) );
  NANDN U3750 ( .A(n54022), .B(n3396), .Z(n3397) );
  NAND U3751 ( .A(n54023), .B(n3397), .Z(n3398) );
  NAND U3752 ( .A(n54024), .B(n3398), .Z(n3399) );
  NANDN U3753 ( .A(n54025), .B(n3399), .Z(n3400) );
  AND U3754 ( .A(n54026), .B(n3400), .Z(n3401) );
  OR U3755 ( .A(n54027), .B(n3401), .Z(n3402) );
  NAND U3756 ( .A(n54028), .B(n3402), .Z(n3403) );
  NAND U3757 ( .A(n54029), .B(n3403), .Z(n3404) );
  NAND U3758 ( .A(n54030), .B(n3404), .Z(n3405) );
  NANDN U3759 ( .A(n54031), .B(n3405), .Z(n3406) );
  AND U3760 ( .A(n54032), .B(n3406), .Z(n3407) );
  OR U3761 ( .A(n54033), .B(n3407), .Z(n3408) );
  NAND U3762 ( .A(n54034), .B(n3408), .Z(n3409) );
  NANDN U3763 ( .A(n54035), .B(n3409), .Z(n3410) );
  NANDN U3764 ( .A(n52190), .B(n3410), .Z(n54036) );
  NANDN U3765 ( .A(n52181), .B(n54058), .Z(n3411) );
  NAND U3766 ( .A(n52180), .B(n3411), .Z(n3412) );
  NANDN U3767 ( .A(n54059), .B(n3412), .Z(n3413) );
  NAND U3768 ( .A(n54060), .B(n3413), .Z(n3414) );
  NAND U3769 ( .A(n54061), .B(n3414), .Z(n3415) );
  AND U3770 ( .A(n54062), .B(n3415), .Z(n3416) );
  OR U3771 ( .A(n54063), .B(n3416), .Z(n3417) );
  NANDN U3772 ( .A(n54064), .B(n3417), .Z(n3418) );
  NAND U3773 ( .A(n54065), .B(n3418), .Z(n3419) );
  NANDN U3774 ( .A(n54066), .B(n3419), .Z(n3420) );
  NAND U3775 ( .A(n54067), .B(n3420), .Z(n3421) );
  AND U3776 ( .A(n54068), .B(n3421), .Z(n3422) );
  NANDN U3777 ( .A(n3422), .B(n54069), .Z(n3423) );
  NAND U3778 ( .A(n54070), .B(n3423), .Z(n3424) );
  NAND U3779 ( .A(n54071), .B(n3424), .Z(n3425) );
  NANDN U3780 ( .A(n54072), .B(n3425), .Z(n54073) );
  NAND U3781 ( .A(n54096), .B(n54095), .Z(n3426) );
  NANDN U3782 ( .A(n54098), .B(n3426), .Z(n3427) );
  ANDN U3783 ( .B(n3427), .A(n54099), .Z(n3428) );
  OR U3784 ( .A(n52170), .B(n52169), .Z(n3429) );
  ANDN U3785 ( .B(n3429), .A(n52171), .Z(n3430) );
  NANDN U3786 ( .A(n3428), .B(n54100), .Z(n3431) );
  NAND U3787 ( .A(n3430), .B(n3431), .Z(n3432) );
  NAND U3788 ( .A(n54101), .B(n3432), .Z(n3433) );
  NANDN U3789 ( .A(n52168), .B(n3433), .Z(n3434) );
  NAND U3790 ( .A(n52167), .B(n3434), .Z(n3435) );
  ANDN U3791 ( .B(n3435), .A(n52166), .Z(n3436) );
  ANDN U3792 ( .B(n52165), .A(n3436), .Z(n3437) );
  NAND U3793 ( .A(n54102), .B(n3437), .Z(n3438) );
  AND U3794 ( .A(n54103), .B(n3438), .Z(n54104) );
  NAND U3795 ( .A(n54130), .B(n54129), .Z(n3439) );
  NAND U3796 ( .A(n54131), .B(n3439), .Z(n3440) );
  ANDN U3797 ( .B(n3440), .A(n54132), .Z(n3441) );
  OR U3798 ( .A(n3441), .B(n54133), .Z(n3442) );
  NANDN U3799 ( .A(n52157), .B(n3442), .Z(n3443) );
  AND U3800 ( .A(n52156), .B(n3443), .Z(n3444) );
  NANDN U3801 ( .A(n54134), .B(n54135), .Z(n3445) );
  NAND U3802 ( .A(n3444), .B(n3445), .Z(n3446) );
  NANDN U3803 ( .A(n54136), .B(n3446), .Z(n3447) );
  NAND U3804 ( .A(n54137), .B(n3447), .Z(n3448) );
  NANDN U3805 ( .A(n54138), .B(n3448), .Z(n3449) );
  AND U3806 ( .A(n54139), .B(n3449), .Z(n3450) );
  OR U3807 ( .A(n54140), .B(n3450), .Z(n3451) );
  NAND U3808 ( .A(n54141), .B(n3451), .Z(n3452) );
  NANDN U3809 ( .A(n54142), .B(n3452), .Z(n3453) );
  AND U3810 ( .A(n54143), .B(n3453), .Z(n54145) );
  NAND U3811 ( .A(n54177), .B(n54178), .Z(n3454) );
  NANDN U3812 ( .A(n54179), .B(n3454), .Z(n3455) );
  NAND U3813 ( .A(n54180), .B(n3455), .Z(n3456) );
  NANDN U3814 ( .A(n54181), .B(n3456), .Z(n3457) );
  NAND U3815 ( .A(n54182), .B(n3457), .Z(n3458) );
  ANDN U3816 ( .B(n3458), .A(n54183), .Z(n3459) );
  NANDN U3817 ( .A(n3459), .B(n54184), .Z(n3460) );
  NANDN U3818 ( .A(n54185), .B(n3460), .Z(n3461) );
  NANDN U3819 ( .A(n54186), .B(n3461), .Z(n3462) );
  NANDN U3820 ( .A(n54187), .B(n3462), .Z(n3463) );
  NAND U3821 ( .A(n54188), .B(n3463), .Z(n3464) );
  ANDN U3822 ( .B(n3464), .A(n54189), .Z(n3465) );
  NANDN U3823 ( .A(n3465), .B(n54190), .Z(n3466) );
  NANDN U3824 ( .A(n54191), .B(n3466), .Z(n3467) );
  NANDN U3825 ( .A(n54192), .B(n3467), .Z(n3468) );
  NAND U3826 ( .A(n54193), .B(n3468), .Z(n3469) );
  NANDN U3827 ( .A(n54194), .B(n3469), .Z(n3470) );
  ANDN U3828 ( .B(n3470), .A(n54195), .Z(n54198) );
  NANDN U3829 ( .A(n27293), .B(n27294), .Z(n54250) );
  NAND U3830 ( .A(n54283), .B(n54282), .Z(n3471) );
  NANDN U3831 ( .A(n54284), .B(n3471), .Z(n3472) );
  NANDN U3832 ( .A(n54285), .B(n3472), .Z(n3473) );
  NAND U3833 ( .A(n54286), .B(n3473), .Z(n3474) );
  NAND U3834 ( .A(n54287), .B(n3474), .Z(n3475) );
  AND U3835 ( .A(n54288), .B(n3475), .Z(n3476) );
  OR U3836 ( .A(n3476), .B(n54289), .Z(n3477) );
  NAND U3837 ( .A(n54290), .B(n3477), .Z(n3478) );
  ANDN U3838 ( .B(n3478), .A(n54291), .Z(n3479) );
  OR U3839 ( .A(n3479), .B(n54292), .Z(n3480) );
  NAND U3840 ( .A(n54293), .B(n3480), .Z(n3481) );
  NANDN U3841 ( .A(n54294), .B(n3481), .Z(n3482) );
  NAND U3842 ( .A(n54295), .B(n3482), .Z(n3483) );
  NANDN U3843 ( .A(n54296), .B(n3483), .Z(n3484) );
  ANDN U3844 ( .B(n3484), .A(n54297), .Z(n3485) );
  NANDN U3845 ( .A(n3485), .B(n54298), .Z(n3486) );
  NANDN U3846 ( .A(n54299), .B(n3486), .Z(n3487) );
  NAND U3847 ( .A(n54300), .B(n3487), .Z(n3488) );
  NANDN U3848 ( .A(n54301), .B(n3488), .Z(n54304) );
  NANDN U3849 ( .A(n54336), .B(n54335), .Z(n3489) );
  ANDN U3850 ( .B(n3489), .A(n54337), .Z(n3490) );
  NANDN U3851 ( .A(n54339), .B(n54338), .Z(n3491) );
  NAND U3852 ( .A(n3490), .B(n3491), .Z(n3492) );
  ANDN U3853 ( .B(n3492), .A(n54340), .Z(n3493) );
  NANDN U3854 ( .A(n3493), .B(n54341), .Z(n3494) );
  NANDN U3855 ( .A(n54342), .B(n3494), .Z(n3495) );
  NAND U3856 ( .A(n54343), .B(n3495), .Z(n3496) );
  AND U3857 ( .A(n52143), .B(n52142), .Z(n3497) );
  NANDN U3858 ( .A(n54344), .B(n3496), .Z(n3498) );
  NAND U3859 ( .A(n3497), .B(n3498), .Z(n3499) );
  ANDN U3860 ( .B(n54346), .A(n54345), .Z(n3500) );
  NAND U3861 ( .A(n3499), .B(n3500), .Z(n3501) );
  NAND U3862 ( .A(n54347), .B(n3501), .Z(n3502) );
  NANDN U3863 ( .A(n3502), .B(n52141), .Z(n3503) );
  ANDN U3864 ( .B(n3503), .A(n54348), .Z(n54351) );
  NAND U3865 ( .A(n54371), .B(n54370), .Z(n3504) );
  NANDN U3866 ( .A(n54373), .B(n3504), .Z(n3505) );
  NANDN U3867 ( .A(n52131), .B(n3505), .Z(n3506) );
  NAND U3868 ( .A(n54374), .B(n3506), .Z(n3507) );
  NANDN U3869 ( .A(n52130), .B(n3507), .Z(n3508) );
  AND U3870 ( .A(n54375), .B(n3508), .Z(n3509) );
  NANDN U3871 ( .A(n3509), .B(n52129), .Z(n3510) );
  NANDN U3872 ( .A(n54376), .B(n3510), .Z(n3511) );
  NAND U3873 ( .A(n54377), .B(n3511), .Z(n3512) );
  NANDN U3874 ( .A(n54378), .B(n3512), .Z(n3513) );
  NAND U3875 ( .A(n54379), .B(n3513), .Z(n3514) );
  ANDN U3876 ( .B(n3514), .A(n54380), .Z(n3515) );
  OR U3877 ( .A(n54381), .B(n3515), .Z(n3516) );
  NAND U3878 ( .A(n54382), .B(n3516), .Z(n3517) );
  NAND U3879 ( .A(n54383), .B(n3517), .Z(n3518) );
  NANDN U3880 ( .A(n54384), .B(n3518), .Z(n54385) );
  NAND U3881 ( .A(n54407), .B(n54408), .Z(n3519) );
  AND U3882 ( .A(n54409), .B(n3519), .Z(n3520) );
  NAND U3883 ( .A(n3520), .B(n52118), .Z(n3521) );
  NANDN U3884 ( .A(n54410), .B(n3521), .Z(n3522) );
  NAND U3885 ( .A(n54411), .B(n3522), .Z(n3523) );
  ANDN U3886 ( .B(n3523), .A(n52117), .Z(n3524) );
  NANDN U3887 ( .A(n3524), .B(n54412), .Z(n3525) );
  NAND U3888 ( .A(n54413), .B(n3525), .Z(n3526) );
  NANDN U3889 ( .A(n54414), .B(n3526), .Z(n3527) );
  NAND U3890 ( .A(n54415), .B(n3527), .Z(n3528) );
  NANDN U3891 ( .A(n54416), .B(n3528), .Z(n3529) );
  AND U3892 ( .A(n54417), .B(n3529), .Z(n3530) );
  OR U3893 ( .A(n3530), .B(n54418), .Z(n3531) );
  NAND U3894 ( .A(n54419), .B(n3531), .Z(n3532) );
  NANDN U3895 ( .A(n54420), .B(n3532), .Z(n54423) );
  NANDN U3896 ( .A(n52112), .B(n54451), .Z(n3533) );
  NAND U3897 ( .A(n52111), .B(n3533), .Z(n3534) );
  NAND U3898 ( .A(n54452), .B(n3534), .Z(n3535) );
  NANDN U3899 ( .A(n54453), .B(n3535), .Z(n3536) );
  NAND U3900 ( .A(n54454), .B(n3536), .Z(n3537) );
  ANDN U3901 ( .B(n3537), .A(n54455), .Z(n3538) );
  NANDN U3902 ( .A(n3538), .B(n54456), .Z(n3539) );
  NANDN U3903 ( .A(n54457), .B(n3539), .Z(n3540) );
  NANDN U3904 ( .A(n54458), .B(n3540), .Z(n3541) );
  NAND U3905 ( .A(n54459), .B(n3541), .Z(n3542) );
  NANDN U3906 ( .A(n54460), .B(n3542), .Z(n3543) );
  AND U3907 ( .A(n54461), .B(n3543), .Z(n3544) );
  OR U3908 ( .A(n54462), .B(n3544), .Z(n3545) );
  ANDN U3909 ( .B(n3545), .A(n54463), .Z(n3546) );
  NANDN U3910 ( .A(n3546), .B(n54464), .Z(n3547) );
  NANDN U3911 ( .A(n54465), .B(n3547), .Z(n3548) );
  NANDN U3912 ( .A(n52110), .B(n3548), .Z(n54466) );
  ANDN U3913 ( .B(n27160), .A(n27159), .Z(n54483) );
  NAND U3914 ( .A(n54504), .B(n54503), .Z(n3549) );
  NANDN U3915 ( .A(n54505), .B(n3549), .Z(n3550) );
  NAND U3916 ( .A(n54506), .B(n3550), .Z(n3551) );
  NANDN U3917 ( .A(n54507), .B(n3551), .Z(n3552) );
  NAND U3918 ( .A(n54508), .B(n3552), .Z(n3553) );
  ANDN U3919 ( .B(n3553), .A(n54509), .Z(n3554) );
  OR U3920 ( .A(n52098), .B(n3554), .Z(n3555) );
  NAND U3921 ( .A(n52097), .B(n3555), .Z(n3556) );
  NANDN U3922 ( .A(n54510), .B(n3556), .Z(n3557) );
  NAND U3923 ( .A(n54511), .B(n3557), .Z(n3558) );
  NANDN U3924 ( .A(n54512), .B(n3558), .Z(n3559) );
  ANDN U3925 ( .B(n3559), .A(n52096), .Z(n3560) );
  NANDN U3926 ( .A(n3560), .B(n52095), .Z(n3561) );
  NANDN U3927 ( .A(n54513), .B(n3561), .Z(n3562) );
  NAND U3928 ( .A(n54514), .B(n3562), .Z(n3563) );
  NANDN U3929 ( .A(n54515), .B(n3563), .Z(n54516) );
  OR U3930 ( .A(n54549), .B(n54550), .Z(n3564) );
  NAND U3931 ( .A(n54551), .B(n3564), .Z(n3565) );
  NANDN U3932 ( .A(n54552), .B(n3565), .Z(n3566) );
  NAND U3933 ( .A(n54553), .B(n3566), .Z(n3567) );
  NANDN U3934 ( .A(n52090), .B(n3567), .Z(n3568) );
  AND U3935 ( .A(n54554), .B(n3568), .Z(n3569) );
  OR U3936 ( .A(n54555), .B(n3569), .Z(n3570) );
  NAND U3937 ( .A(n54556), .B(n3570), .Z(n3571) );
  NANDN U3938 ( .A(n54557), .B(n3571), .Z(n3572) );
  NAND U3939 ( .A(n54558), .B(n3572), .Z(n3573) );
  NANDN U3940 ( .A(n54559), .B(n3573), .Z(n3574) );
  AND U3941 ( .A(n54560), .B(n3574), .Z(n3575) );
  OR U3942 ( .A(n54561), .B(n3575), .Z(n3576) );
  ANDN U3943 ( .B(n3576), .A(n54562), .Z(n3577) );
  NANDN U3944 ( .A(n3577), .B(n54563), .Z(n3578) );
  NANDN U3945 ( .A(n54564), .B(n3578), .Z(n3579) );
  NAND U3946 ( .A(n54565), .B(n3579), .Z(n54568) );
  NAND U3947 ( .A(n54599), .B(n54598), .Z(n3580) );
  NANDN U3948 ( .A(n54601), .B(n3580), .Z(n3581) );
  NANDN U3949 ( .A(n52086), .B(n3581), .Z(n3582) );
  NANDN U3950 ( .A(n54602), .B(n3582), .Z(n3583) );
  NAND U3951 ( .A(n54603), .B(n3583), .Z(n3584) );
  ANDN U3952 ( .B(n3584), .A(n54604), .Z(n3585) );
  OR U3953 ( .A(n54605), .B(n3585), .Z(n3586) );
  NANDN U3954 ( .A(n54606), .B(n3586), .Z(n3587) );
  NAND U3955 ( .A(n54607), .B(n3587), .Z(n3588) );
  NANDN U3956 ( .A(n54608), .B(n3588), .Z(n3589) );
  NAND U3957 ( .A(n54609), .B(n3589), .Z(n3590) );
  ANDN U3958 ( .B(n3590), .A(n54610), .Z(n3591) );
  NANDN U3959 ( .A(n3591), .B(n54611), .Z(n3592) );
  ANDN U3960 ( .B(n3592), .A(n54612), .Z(n3593) );
  NANDN U3961 ( .A(n3593), .B(n54613), .Z(n3594) );
  NANDN U3962 ( .A(n54614), .B(n3594), .Z(n3595) );
  NAND U3963 ( .A(n52085), .B(n3595), .Z(n54616) );
  NAND U3964 ( .A(n54643), .B(n54642), .Z(n3596) );
  NANDN U3965 ( .A(n54644), .B(n3596), .Z(n3597) );
  NAND U3966 ( .A(n54645), .B(n3597), .Z(n3598) );
  NANDN U3967 ( .A(n54646), .B(n3598), .Z(n3599) );
  NAND U3968 ( .A(n54647), .B(n3599), .Z(n3600) );
  ANDN U3969 ( .B(n3600), .A(n54648), .Z(n3601) );
  ANDN U3970 ( .B(n54649), .A(n3601), .Z(n3602) );
  NAND U3971 ( .A(n54650), .B(n3602), .Z(n3603) );
  AND U3972 ( .A(n52078), .B(n3603), .Z(n3604) );
  AND U3973 ( .A(n52077), .B(n52076), .Z(n3605) );
  NANDN U3974 ( .A(n54651), .B(n3604), .Z(n3606) );
  NAND U3975 ( .A(n3605), .B(n3606), .Z(n3607) );
  NANDN U3976 ( .A(n54652), .B(n3607), .Z(n3608) );
  NAND U3977 ( .A(n54653), .B(n3608), .Z(n3609) );
  ANDN U3978 ( .B(n3609), .A(n54654), .Z(n3610) );
  NANDN U3979 ( .A(n3610), .B(n54655), .Z(n3611) );
  NANDN U3980 ( .A(n54656), .B(n3611), .Z(n3612) );
  NANDN U3981 ( .A(n52075), .B(n3612), .Z(n54657) );
  ANDN U3982 ( .B(n27002), .A(n27001), .Z(n54689) );
  AND U3983 ( .A(n54709), .B(n52063), .Z(n3613) );
  OR U3984 ( .A(n52061), .B(n52062), .Z(n3614) );
  AND U3985 ( .A(n3613), .B(n3614), .Z(n3615) );
  NANDN U3986 ( .A(n3615), .B(n54710), .Z(n3616) );
  NANDN U3987 ( .A(n54711), .B(n3616), .Z(n3617) );
  NAND U3988 ( .A(n54712), .B(n3617), .Z(n3618) );
  NANDN U3989 ( .A(n52060), .B(n3618), .Z(n3619) );
  NANDN U3990 ( .A(n54713), .B(n3619), .Z(n3620) );
  AND U3991 ( .A(n54714), .B(n3620), .Z(n3621) );
  OR U3992 ( .A(n54715), .B(n3621), .Z(n3622) );
  NAND U3993 ( .A(n54716), .B(n3622), .Z(n3623) );
  NANDN U3994 ( .A(n54717), .B(n3623), .Z(n3624) );
  ANDN U3995 ( .B(n3624), .A(n54718), .Z(n54720) );
  NANDN U3996 ( .A(n54748), .B(n54749), .Z(n3625) );
  NANDN U3997 ( .A(n54750), .B(n3625), .Z(n3626) );
  NAND U3998 ( .A(n54751), .B(n3626), .Z(n3627) );
  NANDN U3999 ( .A(n54752), .B(n3627), .Z(n3628) );
  NAND U4000 ( .A(n54753), .B(n3628), .Z(n3629) );
  ANDN U4001 ( .B(n3629), .A(n54754), .Z(n3630) );
  NANDN U4002 ( .A(n3630), .B(n54755), .Z(n3631) );
  NANDN U4003 ( .A(n54756), .B(n3631), .Z(n3632) );
  NAND U4004 ( .A(n54757), .B(n3632), .Z(n3633) );
  NANDN U4005 ( .A(n54758), .B(n3633), .Z(n3634) );
  NAND U4006 ( .A(n54759), .B(n3634), .Z(n3635) );
  ANDN U4007 ( .B(n3635), .A(n54760), .Z(n3636) );
  OR U4008 ( .A(n54761), .B(n3636), .Z(n3637) );
  AND U4009 ( .A(n54762), .B(n3637), .Z(n3638) );
  NANDN U4010 ( .A(n3638), .B(n54763), .Z(n3639) );
  NANDN U4011 ( .A(n52054), .B(n3639), .Z(n3640) );
  NAND U4012 ( .A(n52053), .B(n3640), .Z(n54764) );
  NANDN U4013 ( .A(n54798), .B(n54797), .Z(n3641) );
  NANDN U4014 ( .A(n54799), .B(n3641), .Z(n3642) );
  NAND U4015 ( .A(n54800), .B(n3642), .Z(n3643) );
  NANDN U4016 ( .A(n54801), .B(n3643), .Z(n3644) );
  NAND U4017 ( .A(n54802), .B(n3644), .Z(n3645) );
  ANDN U4018 ( .B(n3645), .A(n54803), .Z(n3646) );
  ANDN U4019 ( .B(n52049), .A(n52048), .Z(n3647) );
  NANDN U4020 ( .A(n3646), .B(n54804), .Z(n3648) );
  AND U4021 ( .A(n3647), .B(n3648), .Z(n3649) );
  AND U4022 ( .A(n52047), .B(n54806), .Z(n3650) );
  OR U4023 ( .A(n54805), .B(n3649), .Z(n3651) );
  AND U4024 ( .A(n3650), .B(n3651), .Z(n3652) );
  OR U4025 ( .A(n54807), .B(n3652), .Z(n3653) );
  NAND U4026 ( .A(n54808), .B(n3653), .Z(n3654) );
  NANDN U4027 ( .A(n52046), .B(n3654), .Z(n3655) );
  NANDN U4028 ( .A(n54809), .B(n3655), .Z(n54810) );
  NAND U4029 ( .A(n54829), .B(n54828), .Z(n3656) );
  NAND U4030 ( .A(n52035), .B(n3656), .Z(n3657) );
  ANDN U4031 ( .B(n3657), .A(n54830), .Z(n3658) );
  OR U4032 ( .A(n54831), .B(n3658), .Z(n3659) );
  AND U4033 ( .A(n54832), .B(n3659), .Z(n3660) );
  OR U4034 ( .A(n52034), .B(n3660), .Z(n3661) );
  NAND U4035 ( .A(n52033), .B(n3661), .Z(n3662) );
  NANDN U4036 ( .A(n52032), .B(n3662), .Z(n3663) );
  AND U4037 ( .A(n52031), .B(n52030), .Z(n3664) );
  NAND U4038 ( .A(n3663), .B(n3664), .Z(n3665) );
  NAND U4039 ( .A(n54833), .B(n3665), .Z(n3666) );
  NANDN U4040 ( .A(n52029), .B(n3666), .Z(n54834) );
  ANDN U4041 ( .B(n54866), .A(n54869), .Z(n3667) );
  NAND U4042 ( .A(n54867), .B(n3667), .Z(n3668) );
  AND U4043 ( .A(n54870), .B(n3668), .Z(n3669) );
  OR U4044 ( .A(n3669), .B(n54871), .Z(n3670) );
  NAND U4045 ( .A(n54872), .B(n3670), .Z(n3671) );
  NANDN U4046 ( .A(n54873), .B(n3671), .Z(n3672) );
  NANDN U4047 ( .A(n54874), .B(n3672), .Z(n3673) );
  NAND U4048 ( .A(n54875), .B(n3673), .Z(n3674) );
  ANDN U4049 ( .B(n3674), .A(n54876), .Z(n3675) );
  NOR U4050 ( .A(n3675), .B(n52023), .Z(n3676) );
  NAND U4051 ( .A(n52024), .B(n3676), .Z(n3677) );
  ANDN U4052 ( .B(n3677), .A(n54877), .Z(n3678) );
  NANDN U4053 ( .A(n3678), .B(n54878), .Z(n3679) );
  NAND U4054 ( .A(n54879), .B(n3679), .Z(n3680) );
  NAND U4055 ( .A(n54880), .B(n3680), .Z(n3681) );
  OR U4056 ( .A(n3681), .B(n54881), .Z(n3682) );
  NAND U4057 ( .A(n54882), .B(n3682), .Z(n3683) );
  NANDN U4058 ( .A(n54883), .B(n3683), .Z(n54886) );
  OR U4059 ( .A(n54942), .B(n54941), .Z(n3684) );
  NAND U4060 ( .A(n54943), .B(n3684), .Z(n3685) );
  ANDN U4061 ( .B(n3685), .A(n54944), .Z(n3686) );
  OR U4062 ( .A(n3686), .B(n54945), .Z(n3687) );
  NAND U4063 ( .A(n54946), .B(n3687), .Z(n3688) );
  ANDN U4064 ( .B(n3688), .A(n54947), .Z(n3689) );
  NANDN U4065 ( .A(n3689), .B(n54948), .Z(n3690) );
  NANDN U4066 ( .A(n54949), .B(n3690), .Z(n3691) );
  NANDN U4067 ( .A(n54950), .B(n3691), .Z(n3692) );
  NAND U4068 ( .A(n54951), .B(n3692), .Z(n3693) );
  NANDN U4069 ( .A(n54952), .B(n3693), .Z(n3694) );
  AND U4070 ( .A(n52018), .B(n3694), .Z(n3695) );
  OR U4071 ( .A(n54953), .B(n3695), .Z(n3696) );
  ANDN U4072 ( .B(n3696), .A(n54954), .Z(n3697) );
  NANDN U4073 ( .A(n3697), .B(n54955), .Z(n3698) );
  NANDN U4074 ( .A(n54956), .B(n3698), .Z(n3699) );
  NAND U4075 ( .A(n54957), .B(n3699), .Z(n54958) );
  AND U4076 ( .A(n55033), .B(n55034), .Z(n3700) );
  NANDN U4077 ( .A(n55032), .B(n55031), .Z(n3701) );
  NAND U4078 ( .A(n3700), .B(n3701), .Z(n3702) );
  NAND U4079 ( .A(n52013), .B(n3702), .Z(n3703) );
  NANDN U4080 ( .A(n55035), .B(n3703), .Z(n3704) );
  AND U4081 ( .A(n55036), .B(n3704), .Z(n3705) );
  ANDN U4082 ( .B(n55037), .A(n3705), .Z(n3706) );
  NAND U4083 ( .A(n52012), .B(n3706), .Z(n3707) );
  AND U4084 ( .A(n55038), .B(n3707), .Z(n3708) );
  OR U4085 ( .A(n3708), .B(n55039), .Z(n3709) );
  NAND U4086 ( .A(n55040), .B(n3709), .Z(n3710) );
  ANDN U4087 ( .B(n3710), .A(n55041), .Z(n3711) );
  OR U4088 ( .A(n3711), .B(n55042), .Z(n3712) );
  NAND U4089 ( .A(n55043), .B(n3712), .Z(n3713) );
  NANDN U4090 ( .A(n55044), .B(n3713), .Z(n3714) );
  NAND U4091 ( .A(n55045), .B(n3714), .Z(n55046) );
  NAND U4092 ( .A(n55070), .B(n55069), .Z(n3715) );
  NAND U4093 ( .A(n55071), .B(n3715), .Z(n3716) );
  ANDN U4094 ( .B(n3716), .A(n55072), .Z(n3717) );
  OR U4095 ( .A(n55073), .B(n3717), .Z(n3718) );
  NAND U4096 ( .A(n55074), .B(n3718), .Z(n3719) );
  NANDN U4097 ( .A(n52004), .B(n3719), .Z(n3720) );
  NAND U4098 ( .A(n52003), .B(n3720), .Z(n3721) );
  NANDN U4099 ( .A(n55075), .B(n3721), .Z(n3722) );
  ANDN U4100 ( .B(n3722), .A(n55076), .Z(n3723) );
  NANDN U4101 ( .A(n3723), .B(n55077), .Z(n3724) );
  NANDN U4102 ( .A(n52002), .B(n3724), .Z(n3725) );
  NAND U4103 ( .A(n52001), .B(n3725), .Z(n55078) );
  OR U4104 ( .A(n55099), .B(n55100), .Z(n3726) );
  NANDN U4105 ( .A(n55101), .B(n3726), .Z(n3727) );
  ANDN U4106 ( .B(n3727), .A(n55102), .Z(n3728) );
  NANDN U4107 ( .A(n3728), .B(n55103), .Z(n3729) );
  NANDN U4108 ( .A(n55104), .B(n3729), .Z(n3730) );
  NAND U4109 ( .A(n51992), .B(n3730), .Z(n3731) );
  NANDN U4110 ( .A(n55105), .B(n3731), .Z(n3732) );
  NANDN U4111 ( .A(n55106), .B(n3732), .Z(n3733) );
  AND U4112 ( .A(n55107), .B(n3733), .Z(n3734) );
  OR U4113 ( .A(n3734), .B(n55108), .Z(n3735) );
  NAND U4114 ( .A(n51991), .B(n3735), .Z(n3736) );
  ANDN U4115 ( .B(n3736), .A(n55109), .Z(n3737) );
  OR U4116 ( .A(n3737), .B(n55110), .Z(n3738) );
  NAND U4117 ( .A(n55111), .B(n3738), .Z(n3739) );
  NANDN U4118 ( .A(n55112), .B(n3739), .Z(n55113) );
  NAND U4119 ( .A(n55168), .B(n55167), .Z(n3740) );
  NANDN U4120 ( .A(n55170), .B(n3740), .Z(n3741) );
  NANDN U4121 ( .A(n51987), .B(n3741), .Z(n3742) );
  NAND U4122 ( .A(n51986), .B(n3742), .Z(n3743) );
  NANDN U4123 ( .A(n51985), .B(n3743), .Z(n3744) );
  AND U4124 ( .A(n55171), .B(n3744), .Z(n3745) );
  NAND U4125 ( .A(n3745), .B(n55172), .Z(n3746) );
  NAND U4126 ( .A(n51984), .B(n3746), .Z(n3747) );
  ANDN U4127 ( .B(n3747), .A(n55173), .Z(n3748) );
  NANDN U4128 ( .A(n3748), .B(n55174), .Z(n3749) );
  NANDN U4129 ( .A(n51983), .B(n3749), .Z(n3750) );
  NAND U4130 ( .A(n51982), .B(n3750), .Z(n55178) );
  NANDN U4131 ( .A(n55211), .B(n55210), .Z(n3751) );
  NAND U4132 ( .A(n55213), .B(n3751), .Z(n3752) );
  NAND U4133 ( .A(n55214), .B(n3752), .Z(n3753) );
  NAND U4134 ( .A(n55215), .B(n3753), .Z(n3754) );
  AND U4135 ( .A(n55216), .B(n3754), .Z(n3755) );
  NAND U4136 ( .A(n3755), .B(n55217), .Z(n3756) );
  NAND U4137 ( .A(n55218), .B(n3756), .Z(n3757) );
  NANDN U4138 ( .A(n55219), .B(n3757), .Z(n3758) );
  AND U4139 ( .A(n55220), .B(n3758), .Z(n3759) );
  OR U4140 ( .A(n55221), .B(n3759), .Z(n3760) );
  AND U4141 ( .A(n55222), .B(n3760), .Z(n3761) );
  NOR U4142 ( .A(n51977), .B(n3761), .Z(n3762) );
  NAND U4143 ( .A(n51978), .B(n3762), .Z(n3763) );
  ANDN U4144 ( .B(n3763), .A(n55223), .Z(n3764) );
  NANDN U4145 ( .A(n3764), .B(n55224), .Z(n3765) );
  NANDN U4146 ( .A(n55225), .B(n3765), .Z(n3766) );
  NANDN U4147 ( .A(n55226), .B(n3766), .Z(n3767) );
  AND U4148 ( .A(n55227), .B(n3767), .Z(n55228) );
  NANDN U4149 ( .A(n55273), .B(n55272), .Z(n55275) );
  NAND U4150 ( .A(n55297), .B(n55298), .Z(n3768) );
  NANDN U4151 ( .A(n55299), .B(n3768), .Z(n3769) );
  NAND U4152 ( .A(n51971), .B(n3769), .Z(n3770) );
  NANDN U4153 ( .A(n55300), .B(n3770), .Z(n3771) );
  NANDN U4154 ( .A(n55301), .B(n3771), .Z(n3772) );
  AND U4155 ( .A(n55302), .B(n3772), .Z(n3773) );
  OR U4156 ( .A(n3773), .B(n55303), .Z(n3774) );
  NAND U4157 ( .A(n51970), .B(n3774), .Z(n3775) );
  NANDN U4158 ( .A(n55304), .B(n3775), .Z(n3776) );
  NAND U4159 ( .A(n55305), .B(n3776), .Z(n3777) );
  NANDN U4160 ( .A(n51969), .B(n3777), .Z(n3778) );
  AND U4161 ( .A(n55306), .B(n3778), .Z(n3779) );
  NANDN U4162 ( .A(n55307), .B(n3779), .Z(n55308) );
  NANDN U4163 ( .A(n55382), .B(n55381), .Z(n3780) );
  NAND U4164 ( .A(n55384), .B(n3780), .Z(n3781) );
  ANDN U4165 ( .B(n3781), .A(n55385), .Z(n3782) );
  NANDN U4166 ( .A(n3782), .B(n55386), .Z(n3783) );
  NAND U4167 ( .A(n55387), .B(n3783), .Z(n3784) );
  NANDN U4168 ( .A(n51965), .B(n3784), .Z(n3785) );
  NAND U4169 ( .A(n51964), .B(n3785), .Z(n3786) );
  NANDN U4170 ( .A(n55388), .B(n3786), .Z(n3787) );
  AND U4171 ( .A(n55389), .B(n3787), .Z(n3788) );
  OR U4172 ( .A(n3788), .B(n55390), .Z(n3789) );
  AND U4173 ( .A(n55391), .B(n3789), .Z(n3790) );
  AND U4174 ( .A(n55394), .B(n55393), .Z(n3791) );
  OR U4175 ( .A(n3790), .B(n55392), .Z(n3792) );
  AND U4176 ( .A(n3791), .B(n3792), .Z(n3793) );
  NANDN U4177 ( .A(n3793), .B(n55395), .Z(n3794) );
  NANDN U4178 ( .A(n55396), .B(n3794), .Z(n3795) );
  NAND U4179 ( .A(n55397), .B(n3795), .Z(n55398) );
  NANDN U4180 ( .A(n55436), .B(n55435), .Z(n3796) );
  NAND U4181 ( .A(n55437), .B(n3796), .Z(n3797) );
  NANDN U4182 ( .A(n55438), .B(n3797), .Z(n3798) );
  NAND U4183 ( .A(n55439), .B(n3798), .Z(n3799) );
  NANDN U4184 ( .A(n55440), .B(n3799), .Z(n3800) );
  ANDN U4185 ( .B(n3800), .A(n55441), .Z(n3801) );
  NANDN U4186 ( .A(n3801), .B(n55442), .Z(n3802) );
  AND U4187 ( .A(n55443), .B(n3802), .Z(n3803) );
  OR U4188 ( .A(n51960), .B(n3803), .Z(n3804) );
  NAND U4189 ( .A(n51959), .B(n3804), .Z(n3805) );
  NANDN U4190 ( .A(n51958), .B(n3805), .Z(n3806) );
  AND U4191 ( .A(n51957), .B(n51956), .Z(n3807) );
  NAND U4192 ( .A(n3806), .B(n3807), .Z(n3808) );
  NAND U4193 ( .A(n55444), .B(n3808), .Z(n3809) );
  AND U4194 ( .A(n55445), .B(n3809), .Z(n55446) );
  NANDN U4195 ( .A(n51944), .B(n55464), .Z(n3810) );
  NAND U4196 ( .A(n51943), .B(n3810), .Z(n3811) );
  ANDN U4197 ( .B(n3811), .A(n55465), .Z(n3812) );
  OR U4198 ( .A(n55466), .B(n3812), .Z(n3813) );
  NAND U4199 ( .A(n55467), .B(n3813), .Z(n3814) );
  NANDN U4200 ( .A(n51942), .B(n3814), .Z(n3815) );
  NAND U4201 ( .A(n51941), .B(n3815), .Z(n3816) );
  NANDN U4202 ( .A(n55468), .B(n3816), .Z(n3817) );
  AND U4203 ( .A(n55469), .B(n3817), .Z(n3818) );
  OR U4204 ( .A(n3818), .B(n55470), .Z(n3819) );
  NAND U4205 ( .A(n55471), .B(n3819), .Z(n3820) );
  AND U4206 ( .A(n55472), .B(n3820), .Z(n3821) );
  NAND U4207 ( .A(n3821), .B(n55473), .Z(n55474) );
  NANDN U4208 ( .A(n51932), .B(n55498), .Z(n3822) );
  NANDN U4209 ( .A(n55499), .B(n3822), .Z(n3823) );
  AND U4210 ( .A(n51931), .B(n3823), .Z(n3824) );
  OR U4211 ( .A(n55500), .B(n3824), .Z(n3825) );
  NAND U4212 ( .A(n55501), .B(n3825), .Z(n3826) );
  NANDN U4213 ( .A(n55502), .B(n3826), .Z(n3827) );
  NANDN U4214 ( .A(n55503), .B(n3827), .Z(n3828) );
  NAND U4215 ( .A(n55504), .B(n3828), .Z(n3829) );
  ANDN U4216 ( .B(n3829), .A(n55505), .Z(n3830) );
  NANDN U4217 ( .A(n3830), .B(n55506), .Z(n3831) );
  NANDN U4218 ( .A(n51930), .B(n3831), .Z(n3832) );
  NANDN U4219 ( .A(n55507), .B(n3832), .Z(n55508) );
  NANDN U4220 ( .A(n55534), .B(n55533), .Z(n3833) );
  NAND U4221 ( .A(n51922), .B(n3833), .Z(n3834) );
  ANDN U4222 ( .B(n3834), .A(n55535), .Z(n3835) );
  OR U4223 ( .A(n3835), .B(n55536), .Z(n3836) );
  NAND U4224 ( .A(n55537), .B(n3836), .Z(n3837) );
  NANDN U4225 ( .A(n55538), .B(n3837), .Z(n3838) );
  AND U4226 ( .A(n51921), .B(n3838), .Z(n3839) );
  AND U4227 ( .A(n55541), .B(n55540), .Z(n3840) );
  OR U4228 ( .A(n55539), .B(n3839), .Z(n3841) );
  AND U4229 ( .A(n3840), .B(n3841), .Z(n3842) );
  NANDN U4230 ( .A(n3842), .B(n51920), .Z(n3843) );
  NANDN U4231 ( .A(n55542), .B(n3843), .Z(n3844) );
  NAND U4232 ( .A(n55543), .B(n3844), .Z(n55544) );
  NANDN U4233 ( .A(n55565), .B(n55564), .Z(n3845) );
  NANDN U4234 ( .A(n51911), .B(n3845), .Z(n3846) );
  NAND U4235 ( .A(n51910), .B(n3846), .Z(n3847) );
  NANDN U4236 ( .A(n55566), .B(n3847), .Z(n3848) );
  NAND U4237 ( .A(n55567), .B(n3848), .Z(n3849) );
  ANDN U4238 ( .B(n3849), .A(n51909), .Z(n3850) );
  OR U4239 ( .A(n3850), .B(n55568), .Z(n3851) );
  AND U4240 ( .A(n51908), .B(n3851), .Z(n3852) );
  OR U4241 ( .A(n55569), .B(n3852), .Z(n3853) );
  NAND U4242 ( .A(n55570), .B(n3853), .Z(n3854) );
  NANDN U4243 ( .A(n51907), .B(n3854), .Z(n55571) );
  NANDN U4244 ( .A(n55592), .B(n55591), .Z(n3855) );
  NANDN U4245 ( .A(n55593), .B(n3855), .Z(n3856) );
  NAND U4246 ( .A(n55594), .B(n3856), .Z(n3857) );
  NANDN U4247 ( .A(n51895), .B(n3857), .Z(n3858) );
  NAND U4248 ( .A(n51894), .B(n3858), .Z(n3859) );
  ANDN U4249 ( .B(n3859), .A(n55595), .Z(n3860) );
  OR U4250 ( .A(n55596), .B(n3860), .Z(n3861) );
  NAND U4251 ( .A(n55597), .B(n3861), .Z(n3862) );
  NANDN U4252 ( .A(n51893), .B(n3862), .Z(n3863) );
  NAND U4253 ( .A(n51892), .B(n3863), .Z(n3864) );
  NANDN U4254 ( .A(n55598), .B(n3864), .Z(n3865) );
  ANDN U4255 ( .B(n3865), .A(n55599), .Z(n55602) );
  OR U4256 ( .A(n55629), .B(n55630), .Z(n3866) );
  NANDN U4257 ( .A(n51884), .B(n3866), .Z(n3867) );
  AND U4258 ( .A(n51883), .B(n3867), .Z(n3868) );
  NAND U4259 ( .A(n3868), .B(n55631), .Z(n3869) );
  NANDN U4260 ( .A(n55632), .B(n3869), .Z(n3870) );
  AND U4261 ( .A(n55633), .B(n3870), .Z(n3871) );
  OR U4262 ( .A(n55634), .B(n3871), .Z(n3872) );
  NAND U4263 ( .A(n55635), .B(n3872), .Z(n3873) );
  NANDN U4264 ( .A(n55636), .B(n3873), .Z(n3874) );
  NANDN U4265 ( .A(n55637), .B(n3874), .Z(n3875) );
  NAND U4266 ( .A(n55638), .B(n3875), .Z(n3876) );
  ANDN U4267 ( .B(n3876), .A(n55639), .Z(n3877) );
  ANDN U4268 ( .B(n55641), .A(n55642), .Z(n3878) );
  NANDN U4269 ( .A(n3877), .B(n55640), .Z(n3879) );
  AND U4270 ( .A(n3878), .B(n3879), .Z(n3880) );
  OR U4271 ( .A(n55643), .B(n3880), .Z(n3881) );
  AND U4272 ( .A(n55644), .B(n3881), .Z(n55645) );
  NAND U4273 ( .A(n55744), .B(n55743), .Z(n3882) );
  NANDN U4274 ( .A(n55745), .B(n3882), .Z(n3883) );
  AND U4275 ( .A(n55746), .B(n3883), .Z(n3884) );
  ANDN U4276 ( .B(n51882), .A(n3884), .Z(n3885) );
  NAND U4277 ( .A(n51881), .B(n3885), .Z(n3886) );
  ANDN U4278 ( .B(n3886), .A(n55747), .Z(n3887) );
  NANDN U4279 ( .A(n3887), .B(n55748), .Z(n3888) );
  NANDN U4280 ( .A(n55749), .B(n3888), .Z(n3889) );
  NANDN U4281 ( .A(n55750), .B(n3889), .Z(n3890) );
  NAND U4282 ( .A(n55751), .B(n3890), .Z(n3891) );
  NANDN U4283 ( .A(n55752), .B(n3891), .Z(n3892) );
  AND U4284 ( .A(n55753), .B(n3892), .Z(n3893) );
  OR U4285 ( .A(n3893), .B(n55754), .Z(n3894) );
  NANDN U4286 ( .A(n55755), .B(n3894), .Z(n3895) );
  AND U4287 ( .A(n55756), .B(n3895), .Z(n3896) );
  OR U4288 ( .A(n55757), .B(n3896), .Z(n3897) );
  NAND U4289 ( .A(n55758), .B(n3897), .Z(n3898) );
  NANDN U4290 ( .A(n55759), .B(n3898), .Z(n3899) );
  NANDN U4291 ( .A(n51880), .B(n3899), .Z(n55760) );
  NAND U4292 ( .A(n55791), .B(n55792), .Z(n3900) );
  ANDN U4293 ( .B(n3900), .A(n55793), .Z(n3901) );
  NOR U4294 ( .A(n55794), .B(n3901), .Z(n3902) );
  NAND U4295 ( .A(n55795), .B(n3902), .Z(n3903) );
  ANDN U4296 ( .B(n3903), .A(n55796), .Z(n3904) );
  NANDN U4297 ( .A(n3904), .B(n55797), .Z(n3905) );
  NANDN U4298 ( .A(n51873), .B(n3905), .Z(n3906) );
  NAND U4299 ( .A(n51872), .B(n3906), .Z(n3907) );
  AND U4300 ( .A(n51870), .B(n51869), .Z(n3908) );
  NANDN U4301 ( .A(n51871), .B(n3907), .Z(n3909) );
  NAND U4302 ( .A(n3908), .B(n3909), .Z(n3910) );
  NAND U4303 ( .A(n55798), .B(n3910), .Z(n3911) );
  NANDN U4304 ( .A(n51868), .B(n3911), .Z(n55799) );
  NANDN U4305 ( .A(n55829), .B(n55828), .Z(n3912) );
  NAND U4306 ( .A(n51860), .B(n3912), .Z(n3913) );
  NANDN U4307 ( .A(n55830), .B(n3913), .Z(n3914) );
  AND U4308 ( .A(n55831), .B(n55832), .Z(n3915) );
  NAND U4309 ( .A(n3914), .B(n3915), .Z(n3916) );
  NANDN U4310 ( .A(n55833), .B(n3916), .Z(n3917) );
  NAND U4311 ( .A(n55834), .B(n3917), .Z(n3918) );
  NANDN U4312 ( .A(n55835), .B(n3918), .Z(n3919) );
  AND U4313 ( .A(n55836), .B(n3919), .Z(n3920) );
  NAND U4314 ( .A(n3920), .B(n55837), .Z(n3921) );
  NAND U4315 ( .A(n55838), .B(n3921), .Z(n3922) );
  ANDN U4316 ( .B(n3922), .A(n55839), .Z(n3923) );
  NANDN U4317 ( .A(n3923), .B(n55840), .Z(n3924) );
  NANDN U4318 ( .A(n55841), .B(n3924), .Z(n3925) );
  NAND U4319 ( .A(n51859), .B(n3925), .Z(n3926) );
  ANDN U4320 ( .B(n3926), .A(n55842), .Z(n55844) );
  NAND U4321 ( .A(n55876), .B(n55875), .Z(n3927) );
  ANDN U4322 ( .B(n3927), .A(n55878), .Z(n3928) );
  ANDN U4323 ( .B(n51853), .A(n3928), .Z(n3929) );
  NAND U4324 ( .A(n51852), .B(n3929), .Z(n3930) );
  NAND U4325 ( .A(n55879), .B(n3930), .Z(n3931) );
  NANDN U4326 ( .A(n51851), .B(n3931), .Z(n3932) );
  NAND U4327 ( .A(n51850), .B(n3932), .Z(n3933) );
  ANDN U4328 ( .B(n3933), .A(n55880), .Z(n3934) );
  NANDN U4329 ( .A(n3934), .B(n55881), .Z(n3935) );
  NANDN U4330 ( .A(n55882), .B(n3935), .Z(n3936) );
  NAND U4331 ( .A(n55883), .B(n3936), .Z(n3937) );
  NANDN U4332 ( .A(n51849), .B(n3937), .Z(n55884) );
  AND U4333 ( .A(n55900), .B(n55901), .Z(n3938) );
  AND U4334 ( .A(n51836), .B(n51837), .Z(n3939) );
  NANDN U4335 ( .A(n3938), .B(n55902), .Z(n3940) );
  AND U4336 ( .A(n3939), .B(n3940), .Z(n3941) );
  OR U4337 ( .A(n55903), .B(n3941), .Z(n3942) );
  NAND U4338 ( .A(n55904), .B(n3942), .Z(n3943) );
  NANDN U4339 ( .A(n55905), .B(n3943), .Z(n3944) );
  AND U4340 ( .A(n3944), .B(n55908), .Z(n3945) );
  NANDN U4341 ( .A(n55906), .B(n55907), .Z(n3946) );
  AND U4342 ( .A(n3945), .B(n3946), .Z(n3947) );
  OR U4343 ( .A(n55909), .B(n3947), .Z(n3948) );
  NAND U4344 ( .A(n55910), .B(n3948), .Z(n3949) );
  NANDN U4345 ( .A(n51835), .B(n3949), .Z(n55911) );
  NANDN U4346 ( .A(n55930), .B(n55929), .Z(n3950) );
  NAND U4347 ( .A(n55932), .B(n3950), .Z(n3951) );
  AND U4348 ( .A(n55933), .B(n3951), .Z(n3952) );
  OR U4349 ( .A(n51826), .B(n3952), .Z(n3953) );
  NAND U4350 ( .A(n51825), .B(n3953), .Z(n3954) );
  NANDN U4351 ( .A(n55934), .B(n3954), .Z(n3955) );
  NAND U4352 ( .A(n55935), .B(n3955), .Z(n3956) );
  NAND U4353 ( .A(n55936), .B(n3956), .Z(n3957) );
  AND U4354 ( .A(n55937), .B(n3957), .Z(n3958) );
  NANDN U4355 ( .A(n3958), .B(n55938), .Z(n3959) );
  NANDN U4356 ( .A(n55939), .B(n3959), .Z(n3960) );
  NAND U4357 ( .A(n55940), .B(n3960), .Z(n3961) );
  NANDN U4358 ( .A(n55941), .B(n3961), .Z(n55942) );
  OR U4359 ( .A(n55963), .B(n55962), .Z(n3962) );
  NAND U4360 ( .A(n55964), .B(n3962), .Z(n3963) );
  ANDN U4361 ( .B(n3963), .A(n55965), .Z(n3964) );
  NANDN U4362 ( .A(n3964), .B(n55966), .Z(n3965) );
  NANDN U4363 ( .A(n55967), .B(n3965), .Z(n3966) );
  NAND U4364 ( .A(n51817), .B(n3966), .Z(n3967) );
  NANDN U4365 ( .A(n55968), .B(n3967), .Z(n3968) );
  NAND U4366 ( .A(n55969), .B(n3968), .Z(n3969) );
  ANDN U4367 ( .B(n3969), .A(n51816), .Z(n3970) );
  NANDN U4368 ( .A(n3970), .B(n51815), .Z(n3971) );
  AND U4369 ( .A(n55970), .B(n3971), .Z(n3972) );
  ANDN U4370 ( .B(n55972), .A(n3972), .Z(n3973) );
  NAND U4371 ( .A(n55971), .B(n3973), .Z(n3974) );
  AND U4372 ( .A(n55973), .B(n3974), .Z(n55977) );
  NAND U4373 ( .A(n55996), .B(n51806), .Z(n3975) );
  NANDN U4374 ( .A(n51805), .B(n3975), .Z(n3976) );
  AND U4375 ( .A(n55997), .B(n3976), .Z(n3977) );
  OR U4376 ( .A(n3977), .B(n55998), .Z(n3978) );
  NAND U4377 ( .A(n55999), .B(n3978), .Z(n3979) );
  ANDN U4378 ( .B(n3979), .A(n56000), .Z(n3980) );
  NANDN U4379 ( .A(n3980), .B(n51804), .Z(n3981) );
  NANDN U4380 ( .A(n56001), .B(n3981), .Z(n3982) );
  NAND U4381 ( .A(n56002), .B(n3982), .Z(n3983) );
  NAND U4382 ( .A(n56003), .B(n3983), .Z(n3984) );
  NANDN U4383 ( .A(n56004), .B(n3984), .Z(n3985) );
  AND U4384 ( .A(n56005), .B(n3985), .Z(n3986) );
  OR U4385 ( .A(n56006), .B(n3986), .Z(n3987) );
  NAND U4386 ( .A(n56007), .B(n3987), .Z(n3988) );
  NANDN U4387 ( .A(n56008), .B(n3988), .Z(n56009) );
  NANDN U4388 ( .A(n56035), .B(n56034), .Z(n3989) );
  NANDN U4389 ( .A(n56036), .B(n3989), .Z(n3990) );
  AND U4390 ( .A(n56037), .B(n3990), .Z(n3991) );
  OR U4391 ( .A(n56038), .B(n3991), .Z(n3992) );
  NAND U4392 ( .A(n56039), .B(n3992), .Z(n3993) );
  NANDN U4393 ( .A(n56040), .B(n3993), .Z(n3994) );
  NAND U4394 ( .A(n56041), .B(n3994), .Z(n3995) );
  NANDN U4395 ( .A(n56042), .B(n3995), .Z(n3996) );
  AND U4396 ( .A(n56043), .B(n3996), .Z(n3997) );
  NANDN U4397 ( .A(n3997), .B(n56044), .Z(n3998) );
  AND U4398 ( .A(n56045), .B(n3998), .Z(n3999) );
  ANDN U4399 ( .B(n51797), .A(n3999), .Z(n4000) );
  NAND U4400 ( .A(n51798), .B(n4000), .Z(n4001) );
  AND U4401 ( .A(n56046), .B(n4001), .Z(n4002) );
  NANDN U4402 ( .A(n4002), .B(n56047), .Z(n4003) );
  ANDN U4403 ( .B(n4003), .A(n56048), .Z(n4004) );
  ANDN U4404 ( .B(n56049), .A(n4004), .Z(n4005) );
  OR U4405 ( .A(n56050), .B(n56051), .Z(n4006) );
  NAND U4406 ( .A(n4005), .B(n4006), .Z(n56052) );
  NAND U4407 ( .A(n56074), .B(n56073), .Z(n4007) );
  NAND U4408 ( .A(n56075), .B(n4007), .Z(n4008) );
  ANDN U4409 ( .B(n4008), .A(n51790), .Z(n4009) );
  NANDN U4410 ( .A(n4009), .B(n51789), .Z(n4010) );
  NANDN U4411 ( .A(n56076), .B(n4010), .Z(n4011) );
  NAND U4412 ( .A(n56077), .B(n4011), .Z(n4012) );
  AND U4413 ( .A(n51788), .B(n51787), .Z(n4013) );
  NAND U4414 ( .A(n4012), .B(n4013), .Z(n4014) );
  NAND U4415 ( .A(n56078), .B(n4014), .Z(n4015) );
  ANDN U4416 ( .B(n51786), .A(n51785), .Z(n4016) );
  NAND U4417 ( .A(n4015), .B(n4016), .Z(n4017) );
  NANDN U4418 ( .A(n56079), .B(n4017), .Z(n4018) );
  NAND U4419 ( .A(n56080), .B(n4018), .Z(n56083) );
  NAND U4420 ( .A(n56106), .B(n51779), .Z(n4019) );
  NANDN U4421 ( .A(n56107), .B(n4019), .Z(n4020) );
  AND U4422 ( .A(n56108), .B(n4020), .Z(n4021) );
  OR U4423 ( .A(n4021), .B(n56109), .Z(n4022) );
  NAND U4424 ( .A(n56110), .B(n4022), .Z(n4023) );
  NANDN U4425 ( .A(n56111), .B(n4023), .Z(n4024) );
  NAND U4426 ( .A(n56112), .B(n4024), .Z(n4025) );
  NAND U4427 ( .A(n51778), .B(n4025), .Z(n4026) );
  ANDN U4428 ( .B(n4026), .A(n56113), .Z(n4027) );
  NANDN U4429 ( .A(n4027), .B(n56114), .Z(n4028) );
  NANDN U4430 ( .A(n56115), .B(n4028), .Z(n4029) );
  NAND U4431 ( .A(n56116), .B(n4029), .Z(n4030) );
  NANDN U4432 ( .A(n51777), .B(n4030), .Z(n56117) );
  NAND U4433 ( .A(n56146), .B(n51770), .Z(n4031) );
  NANDN U4434 ( .A(n56147), .B(n4031), .Z(n4032) );
  AND U4435 ( .A(n56148), .B(n4032), .Z(n4033) );
  OR U4436 ( .A(n4033), .B(n56149), .Z(n4034) );
  NAND U4437 ( .A(n56150), .B(n4034), .Z(n4035) );
  NANDN U4438 ( .A(n56151), .B(n4035), .Z(n4036) );
  NAND U4439 ( .A(n56152), .B(n4036), .Z(n4037) );
  NANDN U4440 ( .A(n56153), .B(n4037), .Z(n4038) );
  AND U4441 ( .A(n56154), .B(n4038), .Z(n4039) );
  OR U4442 ( .A(n51769), .B(n4039), .Z(n4040) );
  AND U4443 ( .A(n51768), .B(n4040), .Z(n4041) );
  OR U4444 ( .A(n56155), .B(n4041), .Z(n4042) );
  NAND U4445 ( .A(n56156), .B(n4042), .Z(n4043) );
  NANDN U4446 ( .A(n51767), .B(n4043), .Z(n56157) );
  NAND U4447 ( .A(n56183), .B(n56182), .Z(n4044) );
  NAND U4448 ( .A(n51759), .B(n4044), .Z(n4045) );
  ANDN U4449 ( .B(n4045), .A(n56184), .Z(n4046) );
  NANDN U4450 ( .A(n4046), .B(n56185), .Z(n4047) );
  NAND U4451 ( .A(n56186), .B(n4047), .Z(n4048) );
  NANDN U4452 ( .A(n56187), .B(n4048), .Z(n4049) );
  NAND U4453 ( .A(n56188), .B(n4049), .Z(n4050) );
  NANDN U4454 ( .A(n56189), .B(n4050), .Z(n4051) );
  AND U4455 ( .A(n56190), .B(n4051), .Z(n4052) );
  OR U4456 ( .A(n51758), .B(n4052), .Z(n4053) );
  NAND U4457 ( .A(n51757), .B(n4053), .Z(n4054) );
  NANDN U4458 ( .A(n56191), .B(n4054), .Z(n4055) );
  NAND U4459 ( .A(n56192), .B(n4055), .Z(n56193) );
  NANDN U4460 ( .A(n56222), .B(n56221), .Z(n4056) );
  NANDN U4461 ( .A(n56223), .B(n4056), .Z(n4057) );
  AND U4462 ( .A(n56224), .B(n4057), .Z(n4058) );
  OR U4463 ( .A(n51748), .B(n4058), .Z(n4059) );
  NAND U4464 ( .A(n51747), .B(n4059), .Z(n4060) );
  NANDN U4465 ( .A(n56225), .B(n4060), .Z(n4061) );
  AND U4466 ( .A(n56227), .B(n56226), .Z(n4062) );
  NAND U4467 ( .A(n4061), .B(n4062), .Z(n4063) );
  NANDN U4468 ( .A(n56228), .B(n4063), .Z(n4064) );
  AND U4469 ( .A(n56229), .B(n4064), .Z(n4065) );
  AND U4470 ( .A(n51746), .B(n51745), .Z(n4066) );
  NANDN U4471 ( .A(n4065), .B(n56230), .Z(n4067) );
  AND U4472 ( .A(n4066), .B(n4067), .Z(n56231) );
  OR U4473 ( .A(n56260), .B(n56261), .Z(n4068) );
  NANDN U4474 ( .A(n51738), .B(n4068), .Z(n4069) );
  AND U4475 ( .A(n51737), .B(n4069), .Z(n4070) );
  NANDN U4476 ( .A(n4070), .B(n56262), .Z(n4071) );
  NANDN U4477 ( .A(n56263), .B(n4071), .Z(n4072) );
  NAND U4478 ( .A(n56264), .B(n4072), .Z(n4073) );
  NAND U4479 ( .A(n56265), .B(n4073), .Z(n4074) );
  NANDN U4480 ( .A(n51736), .B(n4074), .Z(n4075) );
  AND U4481 ( .A(n51735), .B(n4075), .Z(n4076) );
  OR U4482 ( .A(n56266), .B(n4076), .Z(n4077) );
  NAND U4483 ( .A(n56267), .B(n4077), .Z(n4078) );
  NANDN U4484 ( .A(n51734), .B(n4078), .Z(n56268) );
  NANDN U4485 ( .A(n56291), .B(n56290), .Z(n4079) );
  NAND U4486 ( .A(n56292), .B(n4079), .Z(n4080) );
  ANDN U4487 ( .B(n4080), .A(n56293), .Z(n4081) );
  NANDN U4488 ( .A(n4081), .B(n51724), .Z(n4082) );
  NANDN U4489 ( .A(n56294), .B(n4082), .Z(n4083) );
  NAND U4490 ( .A(n56295), .B(n4083), .Z(n4084) );
  NANDN U4491 ( .A(n51723), .B(n4084), .Z(n4085) );
  NAND U4492 ( .A(n51722), .B(n4085), .Z(n4086) );
  AND U4493 ( .A(n56296), .B(n4086), .Z(n4087) );
  OR U4494 ( .A(n56297), .B(n4087), .Z(n4088) );
  AND U4495 ( .A(n56298), .B(n4088), .Z(n4089) );
  OR U4496 ( .A(n4089), .B(n56299), .Z(n4090) );
  NAND U4497 ( .A(n56300), .B(n4090), .Z(n4091) );
  NANDN U4498 ( .A(n56301), .B(n4091), .Z(n56302) );
  NAND U4499 ( .A(n56324), .B(n51713), .Z(n4092) );
  NAND U4500 ( .A(n56325), .B(n4092), .Z(n4093) );
  ANDN U4501 ( .B(n4093), .A(n56326), .Z(n4094) );
  ANDN U4502 ( .B(n51712), .A(n4094), .Z(n4095) );
  NAND U4503 ( .A(n51711), .B(n4095), .Z(n4096) );
  ANDN U4504 ( .B(n4096), .A(n56327), .Z(n4097) );
  NANDN U4505 ( .A(n4097), .B(n56328), .Z(n4098) );
  NAND U4506 ( .A(n51710), .B(n4098), .Z(n4099) );
  NAND U4507 ( .A(n56329), .B(n4099), .Z(n4100) );
  NANDN U4508 ( .A(n4100), .B(n56330), .Z(n4101) );
  AND U4509 ( .A(n56331), .B(n4101), .Z(n4102) );
  OR U4510 ( .A(n56332), .B(n4102), .Z(n4103) );
  NAND U4511 ( .A(n56333), .B(n4103), .Z(n4104) );
  NANDN U4512 ( .A(n51709), .B(n4104), .Z(n56334) );
  NAND U4513 ( .A(n56360), .B(n56359), .Z(n4105) );
  NAND U4514 ( .A(n56361), .B(n4105), .Z(n4106) );
  ANDN U4515 ( .B(n4106), .A(n56362), .Z(n4107) );
  NANDN U4516 ( .A(n4107), .B(n56363), .Z(n4108) );
  ANDN U4517 ( .B(n4108), .A(n51702), .Z(n4109) );
  ANDN U4518 ( .B(n56364), .A(n56365), .Z(n4110) );
  NANDN U4519 ( .A(n4109), .B(n51701), .Z(n4111) );
  AND U4520 ( .A(n4110), .B(n4111), .Z(n4112) );
  NANDN U4521 ( .A(n4112), .B(n56366), .Z(n4113) );
  NANDN U4522 ( .A(n56367), .B(n4113), .Z(n4114) );
  NAND U4523 ( .A(n56368), .B(n4114), .Z(n56369) );
  NANDN U4524 ( .A(n56387), .B(n56386), .Z(n4115) );
  NANDN U4525 ( .A(n56388), .B(n4115), .Z(n4116) );
  AND U4526 ( .A(n56389), .B(n4116), .Z(n4117) );
  OR U4527 ( .A(n51688), .B(n4117), .Z(n4118) );
  NAND U4528 ( .A(n51687), .B(n4118), .Z(n4119) );
  NANDN U4529 ( .A(n51686), .B(n4119), .Z(n4120) );
  NAND U4530 ( .A(n56390), .B(n4120), .Z(n4121) );
  NANDN U4531 ( .A(n51685), .B(n4121), .Z(n4122) );
  AND U4532 ( .A(n56391), .B(n4122), .Z(n4123) );
  OR U4533 ( .A(n51684), .B(n4123), .Z(n4124) );
  NAND U4534 ( .A(n56392), .B(n4124), .Z(n4125) );
  NAND U4535 ( .A(n56393), .B(n4125), .Z(n4126) );
  NANDN U4536 ( .A(n56394), .B(n4126), .Z(n56395) );
  NAND U4537 ( .A(n56426), .B(n56425), .Z(n4127) );
  NAND U4538 ( .A(n56429), .B(n4127), .Z(n4128) );
  AND U4539 ( .A(n56430), .B(n4128), .Z(n4129) );
  OR U4540 ( .A(n4129), .B(n56431), .Z(n4130) );
  NAND U4541 ( .A(n56432), .B(n4130), .Z(n4131) );
  NANDN U4542 ( .A(n56433), .B(n4131), .Z(n4132) );
  NAND U4543 ( .A(n56434), .B(n4132), .Z(n4133) );
  NANDN U4544 ( .A(n56435), .B(n4133), .Z(n4134) );
  AND U4545 ( .A(n56436), .B(n4134), .Z(n4135) );
  NANDN U4546 ( .A(n4135), .B(n56437), .Z(n4136) );
  ANDN U4547 ( .B(n4136), .A(n56438), .Z(n4137) );
  NOR U4548 ( .A(n4137), .B(n51678), .Z(n4138) );
  NAND U4549 ( .A(n51679), .B(n4138), .Z(n4139) );
  NANDN U4550 ( .A(n56439), .B(n4139), .Z(n4140) );
  NAND U4551 ( .A(n56440), .B(n4140), .Z(n4141) );
  NANDN U4552 ( .A(n56441), .B(n4141), .Z(n4142) );
  AND U4553 ( .A(n56442), .B(n4142), .Z(n4143) );
  OR U4554 ( .A(n56443), .B(n4143), .Z(n4144) );
  AND U4555 ( .A(n56444), .B(n4144), .Z(n56445) );
  NAND U4556 ( .A(n56511), .B(n56512), .Z(n4145) );
  ANDN U4557 ( .B(n4145), .A(n56513), .Z(n4146) );
  ANDN U4558 ( .B(n51669), .A(n4146), .Z(n4147) );
  NAND U4559 ( .A(n51668), .B(n4147), .Z(n4148) );
  NAND U4560 ( .A(n56514), .B(n4148), .Z(n4149) );
  NANDN U4561 ( .A(n56515), .B(n4149), .Z(n4150) );
  NAND U4562 ( .A(n56516), .B(n4150), .Z(n4151) );
  AND U4563 ( .A(n56517), .B(n4151), .Z(n4152) );
  NAND U4564 ( .A(n4152), .B(n56518), .Z(n4153) );
  NANDN U4565 ( .A(n56519), .B(n4153), .Z(n4154) );
  AND U4566 ( .A(n56520), .B(n4154), .Z(n4155) );
  OR U4567 ( .A(n4155), .B(n56521), .Z(n4156) );
  AND U4568 ( .A(n56522), .B(n4156), .Z(n4157) );
  NANDN U4569 ( .A(n4157), .B(n56523), .Z(n4158) );
  NANDN U4570 ( .A(n56524), .B(n4158), .Z(n4159) );
  NAND U4571 ( .A(n56525), .B(n4159), .Z(n56528) );
  NAND U4572 ( .A(n51659), .B(n56552), .Z(n4160) );
  NANDN U4573 ( .A(n56553), .B(n4160), .Z(n4161) );
  AND U4574 ( .A(n56554), .B(n4161), .Z(n4162) );
  OR U4575 ( .A(n4162), .B(n56555), .Z(n4163) );
  NAND U4576 ( .A(n56556), .B(n4163), .Z(n4164) );
  NANDN U4577 ( .A(n56557), .B(n4164), .Z(n4165) );
  NAND U4578 ( .A(n56558), .B(n4165), .Z(n4166) );
  NANDN U4579 ( .A(n56559), .B(n4166), .Z(n4167) );
  AND U4580 ( .A(n56560), .B(n4167), .Z(n4168) );
  OR U4581 ( .A(n4168), .B(n56561), .Z(n4169) );
  NAND U4582 ( .A(n56562), .B(n4169), .Z(n4170) );
  ANDN U4583 ( .B(n4170), .A(n56563), .Z(n4171) );
  ANDN U4584 ( .B(n56564), .A(n4171), .Z(n4172) );
  NAND U4585 ( .A(n56565), .B(n4172), .Z(n4173) );
  ANDN U4586 ( .B(n4173), .A(n56566), .Z(n4174) );
  NANDN U4587 ( .A(n4174), .B(n56567), .Z(n4175) );
  NANDN U4588 ( .A(n56568), .B(n4175), .Z(n4176) );
  NAND U4589 ( .A(n56569), .B(n4176), .Z(n56570) );
  NAND U4590 ( .A(n56593), .B(n56592), .Z(n4177) );
  NANDN U4591 ( .A(n56595), .B(n4177), .Z(n4178) );
  NANDN U4592 ( .A(n56596), .B(n4178), .Z(n4179) );
  NAND U4593 ( .A(n56597), .B(n4179), .Z(n4180) );
  NANDN U4594 ( .A(n51650), .B(n4180), .Z(n4181) );
  AND U4595 ( .A(n51649), .B(n4181), .Z(n4182) );
  OR U4596 ( .A(n56598), .B(n4182), .Z(n4183) );
  NAND U4597 ( .A(n56599), .B(n4183), .Z(n4184) );
  NANDN U4598 ( .A(n51648), .B(n4184), .Z(n4185) );
  AND U4599 ( .A(n56601), .B(n56600), .Z(n4186) );
  NAND U4600 ( .A(n4185), .B(n4186), .Z(n4187) );
  NANDN U4601 ( .A(n56602), .B(n4187), .Z(n56603) );
  NANDN U4602 ( .A(n56626), .B(n56625), .Z(n4188) );
  NAND U4603 ( .A(n56627), .B(n4188), .Z(n4189) );
  NANDN U4604 ( .A(n56628), .B(n4189), .Z(n4190) );
  NAND U4605 ( .A(n56629), .B(n4190), .Z(n4191) );
  NANDN U4606 ( .A(n51638), .B(n4191), .Z(n4192) );
  AND U4607 ( .A(n51637), .B(n4192), .Z(n4193) );
  OR U4608 ( .A(n56630), .B(n4193), .Z(n4194) );
  AND U4609 ( .A(n56631), .B(n4194), .Z(n4195) );
  AND U4610 ( .A(n56634), .B(n56633), .Z(n4196) );
  OR U4611 ( .A(n4195), .B(n56632), .Z(n4197) );
  AND U4612 ( .A(n4196), .B(n4197), .Z(n4198) );
  OR U4613 ( .A(n4198), .B(n56635), .Z(n4199) );
  NAND U4614 ( .A(n56636), .B(n4199), .Z(n4200) );
  NANDN U4615 ( .A(n56637), .B(n4200), .Z(n56638) );
  NANDN U4616 ( .A(n51629), .B(n56662), .Z(n4201) );
  NAND U4617 ( .A(n51628), .B(n4201), .Z(n4202) );
  ANDN U4618 ( .B(n4202), .A(n56663), .Z(n4203) );
  NANDN U4619 ( .A(n4203), .B(n56664), .Z(n4204) );
  NANDN U4620 ( .A(n51627), .B(n4204), .Z(n4205) );
  NAND U4621 ( .A(n51626), .B(n4205), .Z(n4206) );
  ANDN U4622 ( .B(n56665), .A(n56666), .Z(n4207) );
  NAND U4623 ( .A(n4206), .B(n4207), .Z(n4208) );
  NAND U4624 ( .A(n56667), .B(n4208), .Z(n4209) );
  ANDN U4625 ( .B(n56669), .A(n56668), .Z(n4210) );
  NAND U4626 ( .A(n4209), .B(n4210), .Z(n4211) );
  NANDN U4627 ( .A(n56670), .B(n4211), .Z(n56671) );
  ANDN U4628 ( .B(n51619), .A(n51618), .Z(n4212) );
  NANDN U4629 ( .A(n56697), .B(n56696), .Z(n4213) );
  NAND U4630 ( .A(n4212), .B(n4213), .Z(n4214) );
  ANDN U4631 ( .B(n56699), .A(n56700), .Z(n4215) );
  NANDN U4632 ( .A(n56698), .B(n4214), .Z(n4216) );
  NAND U4633 ( .A(n4215), .B(n4216), .Z(n4217) );
  NANDN U4634 ( .A(n56701), .B(n4217), .Z(n4218) );
  NAND U4635 ( .A(n56702), .B(n4218), .Z(n4219) );
  ANDN U4636 ( .B(n4219), .A(n51616), .Z(n4220) );
  NANDN U4637 ( .A(n4220), .B(n56703), .Z(n4221) );
  ANDN U4638 ( .B(n4221), .A(n56704), .Z(n4222) );
  NANDN U4639 ( .A(n4222), .B(n56705), .Z(n4223) );
  NAND U4640 ( .A(n56706), .B(n4223), .Z(n4224) );
  NANDN U4641 ( .A(n56707), .B(n4224), .Z(n56708) );
  NAND U4642 ( .A(n56738), .B(n56737), .Z(n4225) );
  NAND U4643 ( .A(n56739), .B(n4225), .Z(n4226) );
  NANDN U4644 ( .A(n56740), .B(n4226), .Z(n4227) );
  NAND U4645 ( .A(n56741), .B(n4227), .Z(n4228) );
  NANDN U4646 ( .A(n56742), .B(n4228), .Z(n4229) );
  AND U4647 ( .A(n56743), .B(n4229), .Z(n4230) );
  OR U4648 ( .A(n4230), .B(n56744), .Z(n4231) );
  NAND U4649 ( .A(n56745), .B(n4231), .Z(n4232) );
  NANDN U4650 ( .A(n56746), .B(n4232), .Z(n4233) );
  NAND U4651 ( .A(n56747), .B(n4233), .Z(n4234) );
  NANDN U4652 ( .A(n56748), .B(n4234), .Z(n4235) );
  AND U4653 ( .A(n56749), .B(n4235), .Z(n4236) );
  NANDN U4654 ( .A(n4236), .B(n51609), .Z(n4237) );
  NANDN U4655 ( .A(n56750), .B(n4237), .Z(n4238) );
  NAND U4656 ( .A(n56751), .B(n4238), .Z(n4239) );
  NANDN U4657 ( .A(n51608), .B(n4239), .Z(n56752) );
  NAND U4658 ( .A(n56805), .B(n56806), .Z(n4240) );
  ANDN U4659 ( .B(n4240), .A(n56807), .Z(n4241) );
  ANDN U4660 ( .B(n56808), .A(n4241), .Z(n4242) );
  NAND U4661 ( .A(n56809), .B(n4242), .Z(n4243) );
  NANDN U4662 ( .A(n56810), .B(n4243), .Z(n4244) );
  ANDN U4663 ( .B(n56811), .A(n56812), .Z(n4245) );
  NAND U4664 ( .A(n4244), .B(n4245), .Z(n4246) );
  NAND U4665 ( .A(n56813), .B(n4246), .Z(n4247) );
  ANDN U4666 ( .B(n51604), .A(n51603), .Z(n4248) );
  NAND U4667 ( .A(n4247), .B(n4248), .Z(n4249) );
  NANDN U4668 ( .A(n56814), .B(n4249), .Z(n4250) );
  NAND U4669 ( .A(n56815), .B(n4250), .Z(n4251) );
  NANDN U4670 ( .A(n56816), .B(n4251), .Z(n4252) );
  AND U4671 ( .A(n56817), .B(n4252), .Z(n4253) );
  OR U4672 ( .A(n56818), .B(n4253), .Z(n4254) );
  NAND U4673 ( .A(n56819), .B(n4254), .Z(n4255) );
  NANDN U4674 ( .A(n56820), .B(n4255), .Z(n56821) );
  NAND U4675 ( .A(n56859), .B(n56860), .Z(n4256) );
  NANDN U4676 ( .A(n56861), .B(n4256), .Z(n4257) );
  AND U4677 ( .A(n56862), .B(n4257), .Z(n4258) );
  OR U4678 ( .A(n4258), .B(n56863), .Z(n4259) );
  NAND U4679 ( .A(n56864), .B(n4259), .Z(n4260) );
  NAND U4680 ( .A(n56865), .B(n4260), .Z(n4261) );
  NAND U4681 ( .A(n51600), .B(n4261), .Z(n4262) );
  NANDN U4682 ( .A(n56866), .B(n4262), .Z(n4263) );
  AND U4683 ( .A(n56867), .B(n4263), .Z(n4264) );
  OR U4684 ( .A(n51599), .B(n4264), .Z(n4265) );
  NAND U4685 ( .A(n51598), .B(n4265), .Z(n4266) );
  NANDN U4686 ( .A(n56868), .B(n4266), .Z(n4267) );
  NAND U4687 ( .A(n56869), .B(n4267), .Z(n56872) );
  OR U4688 ( .A(n56895), .B(n56896), .Z(n4268) );
  NANDN U4689 ( .A(n56897), .B(n4268), .Z(n4269) );
  NAND U4690 ( .A(n56898), .B(n4269), .Z(n4270) );
  NANDN U4691 ( .A(n51589), .B(n4270), .Z(n4271) );
  NAND U4692 ( .A(n51588), .B(n4271), .Z(n4272) );
  AND U4693 ( .A(n56899), .B(n4272), .Z(n4273) );
  OR U4694 ( .A(n56900), .B(n4273), .Z(n4274) );
  NAND U4695 ( .A(n56901), .B(n4274), .Z(n4275) );
  NANDN U4696 ( .A(n56902), .B(n4275), .Z(n4276) );
  NAND U4697 ( .A(n56903), .B(n4276), .Z(n4277) );
  NANDN U4698 ( .A(n56904), .B(n4277), .Z(n4278) );
  AND U4699 ( .A(n56905), .B(n4278), .Z(n4279) );
  NANDN U4700 ( .A(n4279), .B(n56906), .Z(n4280) );
  NANDN U4701 ( .A(n56907), .B(n4280), .Z(n4281) );
  NAND U4702 ( .A(n56908), .B(n4281), .Z(n56909) );
  NAND U4703 ( .A(n56937), .B(n56938), .Z(n4282) );
  NANDN U4704 ( .A(n56939), .B(n4282), .Z(n4283) );
  AND U4705 ( .A(n56940), .B(n4283), .Z(n4284) );
  OR U4706 ( .A(n56941), .B(n4284), .Z(n4285) );
  NAND U4707 ( .A(n56942), .B(n4285), .Z(n4286) );
  NANDN U4708 ( .A(n56943), .B(n4286), .Z(n4287) );
  NAND U4709 ( .A(n56944), .B(n4287), .Z(n4288) );
  NANDN U4710 ( .A(n56945), .B(n4288), .Z(n4289) );
  AND U4711 ( .A(n56946), .B(n4289), .Z(n4290) );
  OR U4712 ( .A(n56947), .B(n4290), .Z(n4291) );
  NAND U4713 ( .A(n56948), .B(n4291), .Z(n4292) );
  NANDN U4714 ( .A(n56949), .B(n4292), .Z(n4293) );
  AND U4715 ( .A(n51580), .B(n51579), .Z(n4294) );
  NAND U4716 ( .A(n4293), .B(n4294), .Z(n4295) );
  NANDN U4717 ( .A(n56950), .B(n4295), .Z(n4296) );
  NAND U4718 ( .A(n56951), .B(n4296), .Z(n4297) );
  NANDN U4719 ( .A(n56952), .B(n4297), .Z(n4298) );
  ANDN U4720 ( .B(n4298), .A(n56953), .Z(n56955) );
  ANDN U4721 ( .B(n56973), .A(n56974), .Z(n56975) );
  NAND U4722 ( .A(n57011), .B(n57010), .Z(n4299) );
  NAND U4723 ( .A(n57012), .B(n4299), .Z(n4300) );
  AND U4724 ( .A(n57013), .B(n4300), .Z(n4301) );
  NAND U4725 ( .A(n4301), .B(n57014), .Z(n4302) );
  NAND U4726 ( .A(n51570), .B(n4302), .Z(n4303) );
  AND U4727 ( .A(n57015), .B(n4303), .Z(n4304) );
  NAND U4728 ( .A(n4304), .B(n57016), .Z(n4305) );
  NANDN U4729 ( .A(n57017), .B(n4305), .Z(n4306) );
  AND U4730 ( .A(n57018), .B(n4306), .Z(n4307) );
  OR U4731 ( .A(n57019), .B(n4307), .Z(n4308) );
  NAND U4732 ( .A(n57020), .B(n4308), .Z(n4309) );
  NANDN U4733 ( .A(n57021), .B(n4309), .Z(n4310) );
  NAND U4734 ( .A(n57022), .B(n4310), .Z(n4311) );
  NANDN U4735 ( .A(n57023), .B(n4311), .Z(n4312) );
  AND U4736 ( .A(n57024), .B(n4312), .Z(n4313) );
  OR U4737 ( .A(n57025), .B(n4313), .Z(n4314) );
  NAND U4738 ( .A(n57026), .B(n4314), .Z(n4315) );
  NANDN U4739 ( .A(n57027), .B(n4315), .Z(n4316) );
  AND U4740 ( .A(n57028), .B(n4316), .Z(n57030) );
  NANDN U4741 ( .A(n57050), .B(n57049), .Z(n4317) );
  AND U4742 ( .A(n57052), .B(n4317), .Z(n4318) );
  NOR U4743 ( .A(n57054), .B(n4318), .Z(n4319) );
  NAND U4744 ( .A(n57055), .B(n4319), .Z(n4320) );
  NANDN U4745 ( .A(n57056), .B(n4320), .Z(n4321) );
  NAND U4746 ( .A(n57057), .B(n4321), .Z(n4322) );
  NANDN U4747 ( .A(n57058), .B(n4322), .Z(n4323) );
  AND U4748 ( .A(n57059), .B(n4323), .Z(n4324) );
  AND U4749 ( .A(n57061), .B(n57062), .Z(n4325) );
  OR U4750 ( .A(n57060), .B(n4324), .Z(n4326) );
  AND U4751 ( .A(n4325), .B(n4326), .Z(n4327) );
  AND U4752 ( .A(n57064), .B(n57063), .Z(n4328) );
  NANDN U4753 ( .A(n4327), .B(n51560), .Z(n4329) );
  AND U4754 ( .A(n4328), .B(n4329), .Z(n4330) );
  OR U4755 ( .A(n57065), .B(n4330), .Z(n4331) );
  NAND U4756 ( .A(n57066), .B(n4331), .Z(n4332) );
  NANDN U4757 ( .A(n57067), .B(n4332), .Z(n57068) );
  AND U4758 ( .A(n51553), .B(n57098), .Z(n4333) );
  NAND U4759 ( .A(n51554), .B(n4333), .Z(n4334) );
  AND U4760 ( .A(n57099), .B(n4334), .Z(n4335) );
  OR U4761 ( .A(n51551), .B(n4335), .Z(n4336) );
  NAND U4762 ( .A(n51550), .B(n4336), .Z(n4337) );
  NANDN U4763 ( .A(n57100), .B(n4337), .Z(n4338) );
  NAND U4764 ( .A(n57101), .B(n4338), .Z(n4339) );
  NAND U4765 ( .A(n57102), .B(n4339), .Z(n4340) );
  ANDN U4766 ( .B(n4340), .A(n57103), .Z(n4341) );
  NANDN U4767 ( .A(n4341), .B(n57104), .Z(n4342) );
  NANDN U4768 ( .A(n57105), .B(n4342), .Z(n4343) );
  NAND U4769 ( .A(n57106), .B(n4343), .Z(n4344) );
  AND U4770 ( .A(n51548), .B(n51549), .Z(n4345) );
  NANDN U4771 ( .A(n57107), .B(n4344), .Z(n4346) );
  NAND U4772 ( .A(n4345), .B(n4346), .Z(n57110) );
  AND U4773 ( .A(n57143), .B(n57142), .Z(n57144) );
  ANDN U4774 ( .B(n57173), .A(n57172), .Z(n4347) );
  NAND U4775 ( .A(n57170), .B(n57169), .Z(n4348) );
  AND U4776 ( .A(n4347), .B(n4348), .Z(n4349) );
  AND U4777 ( .A(n57176), .B(n57175), .Z(n4350) );
  OR U4778 ( .A(n4349), .B(n57174), .Z(n4351) );
  AND U4779 ( .A(n4350), .B(n4351), .Z(n4352) );
  AND U4780 ( .A(n57179), .B(n57178), .Z(n4353) );
  NANDN U4781 ( .A(n4352), .B(n57177), .Z(n4354) );
  AND U4782 ( .A(n4353), .B(n4354), .Z(n4355) );
  NANDN U4783 ( .A(n4355), .B(n57180), .Z(n4356) );
  ANDN U4784 ( .B(n4356), .A(n57181), .Z(n4357) );
  NANDN U4785 ( .A(n4357), .B(n57182), .Z(n4358) );
  NANDN U4786 ( .A(n51536), .B(n4358), .Z(n4359) );
  NAND U4787 ( .A(n51535), .B(n4359), .Z(n57183) );
  NAND U4788 ( .A(n57214), .B(n57215), .Z(n4360) );
  ANDN U4789 ( .B(n4360), .A(n57216), .Z(n4361) );
  ANDN U4790 ( .B(n57217), .A(n4361), .Z(n4362) );
  NAND U4791 ( .A(n57218), .B(n4362), .Z(n4363) );
  ANDN U4792 ( .B(n4363), .A(n57219), .Z(n4364) );
  ANDN U4793 ( .B(n57221), .A(n4364), .Z(n4365) );
  NAND U4794 ( .A(n57220), .B(n4365), .Z(n4366) );
  AND U4795 ( .A(n57222), .B(n4366), .Z(n4367) );
  ANDN U4796 ( .B(n51530), .A(n4367), .Z(n4368) );
  NAND U4797 ( .A(n57223), .B(n4368), .Z(n4369) );
  ANDN U4798 ( .B(n4369), .A(n51529), .Z(n4370) );
  NANDN U4799 ( .A(n4370), .B(n51528), .Z(n4371) );
  ANDN U4800 ( .B(n4371), .A(n57224), .Z(n57227) );
  ANDN U4801 ( .B(n57253), .A(n57255), .Z(n4372) );
  NAND U4802 ( .A(n57254), .B(n4372), .Z(n4373) );
  NAND U4803 ( .A(n57256), .B(n4373), .Z(n4374) );
  ANDN U4804 ( .B(n51522), .A(n51521), .Z(n4375) );
  NAND U4805 ( .A(n4374), .B(n4375), .Z(n4376) );
  NAND U4806 ( .A(n57257), .B(n4376), .Z(n4377) );
  ANDN U4807 ( .B(n57259), .A(n57258), .Z(n4378) );
  NAND U4808 ( .A(n4377), .B(n4378), .Z(n4379) );
  NANDN U4809 ( .A(n57260), .B(n4379), .Z(n4380) );
  ANDN U4810 ( .B(n51520), .A(n57261), .Z(n4381) );
  NAND U4811 ( .A(n4380), .B(n4381), .Z(n4382) );
  NAND U4812 ( .A(n57262), .B(n4382), .Z(n4383) );
  NANDN U4813 ( .A(n57263), .B(n4383), .Z(n4384) );
  NAND U4814 ( .A(n57264), .B(n4384), .Z(n4385) );
  AND U4815 ( .A(n57266), .B(n4385), .Z(n4386) );
  NANDN U4816 ( .A(n57265), .B(n4386), .Z(n57267) );
  NAND U4817 ( .A(n57297), .B(n57296), .Z(n4387) );
  AND U4818 ( .A(n57298), .B(n4387), .Z(n4388) );
  ANDN U4819 ( .B(n57300), .A(n4388), .Z(n4389) );
  NAND U4820 ( .A(n57301), .B(n4389), .Z(n4390) );
  NANDN U4821 ( .A(n57302), .B(n4390), .Z(n4391) );
  ANDN U4822 ( .B(n57303), .A(n57304), .Z(n4392) );
  NAND U4823 ( .A(n4391), .B(n4392), .Z(n4393) );
  NANDN U4824 ( .A(n57305), .B(n4393), .Z(n4394) );
  ANDN U4825 ( .B(n57307), .A(n57306), .Z(n4395) );
  NAND U4826 ( .A(n4394), .B(n4395), .Z(n4396) );
  NAND U4827 ( .A(n57308), .B(n4396), .Z(n4397) );
  ANDN U4828 ( .B(n57310), .A(n57309), .Z(n4398) );
  NAND U4829 ( .A(n4397), .B(n4398), .Z(n4399) );
  NAND U4830 ( .A(n51510), .B(n4399), .Z(n4400) );
  ANDN U4831 ( .B(n57312), .A(n57311), .Z(n4401) );
  NAND U4832 ( .A(n4400), .B(n4401), .Z(n4402) );
  NANDN U4833 ( .A(n57313), .B(n4402), .Z(n57315) );
  ANDN U4834 ( .B(n57350), .A(n57351), .Z(n4403) );
  NANDN U4835 ( .A(n57348), .B(n57347), .Z(n4404) );
  NAND U4836 ( .A(n4403), .B(n4404), .Z(n4405) );
  NANDN U4837 ( .A(n51505), .B(n4405), .Z(n4406) );
  NAND U4838 ( .A(n51504), .B(n4406), .Z(n4407) );
  ANDN U4839 ( .B(n4407), .A(n57352), .Z(n4408) );
  ANDN U4840 ( .B(n57354), .A(n4408), .Z(n4409) );
  NAND U4841 ( .A(n57353), .B(n4409), .Z(n4410) );
  ANDN U4842 ( .B(n4410), .A(n57355), .Z(n4411) );
  NOR U4843 ( .A(n57357), .B(n4411), .Z(n4412) );
  NAND U4844 ( .A(n57356), .B(n4412), .Z(n4413) );
  ANDN U4845 ( .B(n4413), .A(n51503), .Z(n4414) );
  NANDN U4846 ( .A(n4414), .B(n57358), .Z(n4415) );
  ANDN U4847 ( .B(n4415), .A(n57359), .Z(n57363) );
  ANDN U4848 ( .B(n57391), .A(n57390), .Z(n4416) );
  NAND U4849 ( .A(n57392), .B(n4416), .Z(n4417) );
  NANDN U4850 ( .A(n57393), .B(n4417), .Z(n4418) );
  NAND U4851 ( .A(n57394), .B(n4418), .Z(n4419) );
  NANDN U4852 ( .A(n57395), .B(n4419), .Z(n4420) );
  AND U4853 ( .A(n57396), .B(n4420), .Z(n4421) );
  ANDN U4854 ( .B(n57398), .A(n57399), .Z(n4422) );
  OR U4855 ( .A(n57397), .B(n4421), .Z(n4423) );
  AND U4856 ( .A(n4422), .B(n4423), .Z(n4424) );
  ANDN U4857 ( .B(n51495), .A(n51496), .Z(n4425) );
  NANDN U4858 ( .A(n4424), .B(n57400), .Z(n4426) );
  AND U4859 ( .A(n4425), .B(n4426), .Z(n4427) );
  ANDN U4860 ( .B(n57403), .A(n57402), .Z(n4428) );
  NANDN U4861 ( .A(n4427), .B(n57401), .Z(n4429) );
  AND U4862 ( .A(n4428), .B(n4429), .Z(n4430) );
  ANDN U4863 ( .B(n57406), .A(n57405), .Z(n4431) );
  OR U4864 ( .A(n4430), .B(n57404), .Z(n4432) );
  AND U4865 ( .A(n4431), .B(n4432), .Z(n57408) );
  NANDN U4866 ( .A(n57436), .B(n57435), .Z(n4433) );
  AND U4867 ( .A(n57437), .B(n4433), .Z(n4434) );
  OR U4868 ( .A(n4434), .B(n57438), .Z(n4435) );
  NAND U4869 ( .A(n57439), .B(n4435), .Z(n4436) );
  NANDN U4870 ( .A(n57440), .B(n4436), .Z(n4437) );
  AND U4871 ( .A(n57442), .B(n57441), .Z(n4438) );
  NAND U4872 ( .A(n4437), .B(n4438), .Z(n4439) );
  NAND U4873 ( .A(n57443), .B(n4439), .Z(n4440) );
  AND U4874 ( .A(n51489), .B(n51488), .Z(n4441) );
  NAND U4875 ( .A(n4440), .B(n4441), .Z(n4442) );
  NANDN U4876 ( .A(n57444), .B(n4442), .Z(n4443) );
  NAND U4877 ( .A(n57445), .B(n4443), .Z(n4444) );
  NANDN U4878 ( .A(n57446), .B(n4444), .Z(n4445) );
  AND U4879 ( .A(n57447), .B(n4445), .Z(n4446) );
  OR U4880 ( .A(n57448), .B(n4446), .Z(n4447) );
  AND U4881 ( .A(n57449), .B(n4447), .Z(n4448) );
  OR U4882 ( .A(n4448), .B(n57450), .Z(n4449) );
  NAND U4883 ( .A(n57451), .B(n4449), .Z(n4450) );
  NANDN U4884 ( .A(n57452), .B(n4450), .Z(n57453) );
  ANDN U4885 ( .B(n57484), .A(n57485), .Z(n4451) );
  NANDN U4886 ( .A(n57483), .B(n57482), .Z(n4452) );
  AND U4887 ( .A(n4451), .B(n4452), .Z(n4453) );
  ANDN U4888 ( .B(n57488), .A(n57487), .Z(n4454) );
  OR U4889 ( .A(n57486), .B(n4453), .Z(n4455) );
  AND U4890 ( .A(n4454), .B(n4455), .Z(n4456) );
  AND U4891 ( .A(n51477), .B(n51478), .Z(n4457) );
  NANDN U4892 ( .A(n4456), .B(n57489), .Z(n4458) );
  AND U4893 ( .A(n4457), .B(n4458), .Z(n4459) );
  ANDN U4894 ( .B(n57492), .A(n57491), .Z(n4460) );
  NANDN U4895 ( .A(n4459), .B(n57490), .Z(n4461) );
  AND U4896 ( .A(n4460), .B(n4461), .Z(n4462) );
  OR U4897 ( .A(n57493), .B(n4462), .Z(n4463) );
  NAND U4898 ( .A(n57494), .B(n4463), .Z(n4464) );
  NANDN U4899 ( .A(n51476), .B(n4464), .Z(n57495) );
  OR U4900 ( .A(n57524), .B(n57523), .Z(n4465) );
  NAND U4901 ( .A(n57525), .B(n4465), .Z(n4466) );
  ANDN U4902 ( .B(n4466), .A(n57526), .Z(n4467) );
  ANDN U4903 ( .B(n57528), .A(n4467), .Z(n4468) );
  NAND U4904 ( .A(n57527), .B(n4468), .Z(n4469) );
  ANDN U4905 ( .B(n4469), .A(n57529), .Z(n4470) );
  NOR U4906 ( .A(n51467), .B(n4470), .Z(n4471) );
  NAND U4907 ( .A(n51466), .B(n4471), .Z(n4472) );
  AND U4908 ( .A(n57530), .B(n4472), .Z(n4473) );
  NOR U4909 ( .A(n57532), .B(n4473), .Z(n4474) );
  NAND U4910 ( .A(n57531), .B(n4474), .Z(n4475) );
  ANDN U4911 ( .B(n4475), .A(n57533), .Z(n4476) );
  NOR U4912 ( .A(n57535), .B(n4476), .Z(n4477) );
  NAND U4913 ( .A(n57534), .B(n4477), .Z(n4478) );
  AND U4914 ( .A(n57536), .B(n4478), .Z(n4479) );
  OR U4915 ( .A(n57537), .B(n4479), .Z(n4480) );
  AND U4916 ( .A(n57538), .B(n4480), .Z(n57542) );
  NAND U4917 ( .A(n57565), .B(n57564), .Z(n4481) );
  AND U4918 ( .A(n57566), .B(n4481), .Z(n4482) );
  NOR U4919 ( .A(n51456), .B(n4482), .Z(n4483) );
  NAND U4920 ( .A(n51455), .B(n4483), .Z(n4484) );
  ANDN U4921 ( .B(n4484), .A(n57567), .Z(n4485) );
  NANDN U4922 ( .A(n4485), .B(n57568), .Z(n4486) );
  NANDN U4923 ( .A(n51454), .B(n4486), .Z(n4487) );
  NAND U4924 ( .A(n51453), .B(n4487), .Z(n4488) );
  ANDN U4925 ( .B(n57570), .A(n57571), .Z(n4489) );
  NANDN U4926 ( .A(n57569), .B(n4488), .Z(n4490) );
  NAND U4927 ( .A(n4489), .B(n4490), .Z(n4491) );
  NAND U4928 ( .A(n51452), .B(n4491), .Z(n57574) );
  OR U4929 ( .A(n57613), .B(n57614), .Z(n4492) );
  AND U4930 ( .A(n57615), .B(n4492), .Z(n4493) );
  AND U4931 ( .A(n57617), .B(n57618), .Z(n4494) );
  NANDN U4932 ( .A(n4493), .B(n57616), .Z(n4495) );
  AND U4933 ( .A(n4494), .B(n4495), .Z(n4496) );
  AND U4934 ( .A(n51440), .B(n57620), .Z(n4497) );
  OR U4935 ( .A(n57619), .B(n4496), .Z(n4498) );
  AND U4936 ( .A(n4497), .B(n4498), .Z(n4499) );
  NANDN U4937 ( .A(n4499), .B(n57621), .Z(n4500) );
  NANDN U4938 ( .A(n57622), .B(n4500), .Z(n4501) );
  NAND U4939 ( .A(n57623), .B(n4501), .Z(n4502) );
  AND U4940 ( .A(n57624), .B(n57625), .Z(n4503) );
  NAND U4941 ( .A(n4502), .B(n4503), .Z(n4504) );
  NAND U4942 ( .A(n51439), .B(n4504), .Z(n4505) );
  AND U4943 ( .A(n57626), .B(n57627), .Z(n4506) );
  NAND U4944 ( .A(n4505), .B(n4506), .Z(n4507) );
  NANDN U4945 ( .A(n57628), .B(n4507), .Z(n57630) );
  NANDN U4946 ( .A(n57657), .B(n57658), .Z(n57659) );
  AND U4947 ( .A(n57696), .B(n57697), .Z(n4508) );
  AND U4948 ( .A(n51419), .B(n51418), .Z(n4509) );
  NANDN U4949 ( .A(n4508), .B(n57698), .Z(n4510) );
  AND U4950 ( .A(n4509), .B(n4510), .Z(n4511) );
  OR U4951 ( .A(n57699), .B(n4511), .Z(n4512) );
  NAND U4952 ( .A(n57700), .B(n4512), .Z(n4513) );
  NAND U4953 ( .A(n51417), .B(n4513), .Z(n4514) );
  AND U4954 ( .A(n57702), .B(n57701), .Z(n4515) );
  NAND U4955 ( .A(n4514), .B(n4515), .Z(n4516) );
  NAND U4956 ( .A(n57703), .B(n4516), .Z(n4517) );
  ANDN U4957 ( .B(n51416), .A(n51415), .Z(n4518) );
  NAND U4958 ( .A(n4517), .B(n4518), .Z(n4519) );
  NAND U4959 ( .A(n57704), .B(n4519), .Z(n4520) );
  ANDN U4960 ( .B(n57705), .A(n57706), .Z(n4521) );
  NAND U4961 ( .A(n4520), .B(n4521), .Z(n4522) );
  NANDN U4962 ( .A(n57707), .B(n4522), .Z(n4523) );
  AND U4963 ( .A(n57708), .B(n4523), .Z(n57711) );
  NANDN U4964 ( .A(n57736), .B(n57735), .Z(n4524) );
  ANDN U4965 ( .B(n4524), .A(n57737), .Z(n4525) );
  NOR U4966 ( .A(n57739), .B(n4525), .Z(n4526) );
  NAND U4967 ( .A(n57738), .B(n4526), .Z(n4527) );
  NANDN U4968 ( .A(n57740), .B(n4527), .Z(n4528) );
  NAND U4969 ( .A(n57741), .B(n4528), .Z(n4529) );
  NANDN U4970 ( .A(n51407), .B(n4529), .Z(n4530) );
  AND U4971 ( .A(n51406), .B(n4530), .Z(n4531) );
  ANDN U4972 ( .B(n57742), .A(n57743), .Z(n4532) );
  OR U4973 ( .A(n51405), .B(n4531), .Z(n4533) );
  AND U4974 ( .A(n4532), .B(n4533), .Z(n4534) );
  NANDN U4975 ( .A(n4534), .B(n51404), .Z(n4535) );
  AND U4976 ( .A(n57744), .B(n4535), .Z(n57746) );
  NAND U4977 ( .A(n57768), .B(n57767), .Z(n4536) );
  AND U4978 ( .A(n57771), .B(n4536), .Z(n4537) );
  ANDN U4979 ( .B(n57773), .A(n57774), .Z(n4538) );
  OR U4980 ( .A(n57772), .B(n4537), .Z(n4539) );
  AND U4981 ( .A(n4538), .B(n4539), .Z(n4540) );
  OR U4982 ( .A(n51394), .B(n4540), .Z(n4541) );
  NAND U4983 ( .A(n57775), .B(n4541), .Z(n4542) );
  NAND U4984 ( .A(n57776), .B(n4542), .Z(n4543) );
  ANDN U4985 ( .B(n57778), .A(n57777), .Z(n4544) );
  NAND U4986 ( .A(n4543), .B(n4544), .Z(n4545) );
  NANDN U4987 ( .A(n57779), .B(n4545), .Z(n4546) );
  ANDN U4988 ( .B(n57781), .A(n57780), .Z(n4547) );
  NAND U4989 ( .A(n4546), .B(n4547), .Z(n4548) );
  NAND U4990 ( .A(n57782), .B(n4548), .Z(n4549) );
  AND U4991 ( .A(n57784), .B(n57783), .Z(n4550) );
  NAND U4992 ( .A(n4549), .B(n4550), .Z(n4551) );
  NAND U4993 ( .A(n57785), .B(n4551), .Z(n57786) );
  NAND U4994 ( .A(n57815), .B(n57816), .Z(n4552) );
  ANDN U4995 ( .B(n4552), .A(n57818), .Z(n4553) );
  NANDN U4996 ( .A(n57819), .B(n4553), .Z(n4554) );
  ANDN U4997 ( .B(n51387), .A(n51386), .Z(n4555) );
  NANDN U4998 ( .A(n57820), .B(n4554), .Z(n4556) );
  NAND U4999 ( .A(n4555), .B(n4556), .Z(n4557) );
  NAND U5000 ( .A(n57821), .B(n4557), .Z(n4558) );
  AND U5001 ( .A(n57823), .B(n4558), .Z(n4559) );
  NANDN U5002 ( .A(n57822), .B(n4559), .Z(n4560) );
  ANDN U5003 ( .B(n57826), .A(n57825), .Z(n4561) );
  NANDN U5004 ( .A(n57824), .B(n4560), .Z(n4562) );
  NAND U5005 ( .A(n4561), .B(n4562), .Z(n4563) );
  AND U5006 ( .A(n57828), .B(n57827), .Z(n4564) );
  NANDN U5007 ( .A(n51385), .B(n4563), .Z(n4565) );
  NAND U5008 ( .A(n4564), .B(n4565), .Z(n4566) );
  NANDN U5009 ( .A(n57829), .B(n4566), .Z(n57830) );
  OR U5010 ( .A(n57881), .B(n57882), .Z(n4567) );
  AND U5011 ( .A(n57883), .B(n4567), .Z(n4568) );
  AND U5012 ( .A(n57885), .B(n57884), .Z(n4569) );
  NANDN U5013 ( .A(n4568), .B(n51372), .Z(n4570) );
  AND U5014 ( .A(n4569), .B(n4570), .Z(n4571) );
  ANDN U5015 ( .B(n51371), .A(n51370), .Z(n4572) );
  OR U5016 ( .A(n4571), .B(n57886), .Z(n4573) );
  AND U5017 ( .A(n4572), .B(n4573), .Z(n4574) );
  ANDN U5018 ( .B(n57888), .A(n57889), .Z(n4575) );
  OR U5019 ( .A(n57887), .B(n4574), .Z(n4576) );
  AND U5020 ( .A(n4575), .B(n4576), .Z(n4577) );
  OR U5021 ( .A(n57890), .B(n4577), .Z(n4578) );
  NAND U5022 ( .A(n57891), .B(n4578), .Z(n4579) );
  NANDN U5023 ( .A(n51369), .B(n4579), .Z(n57892) );
  NANDN U5024 ( .A(n57921), .B(n57920), .Z(n4580) );
  NANDN U5025 ( .A(n57922), .B(n4580), .Z(n4581) );
  NAND U5026 ( .A(n57923), .B(n4581), .Z(n4582) );
  NANDN U5027 ( .A(n4582), .B(n51364), .Z(n4583) );
  NANDN U5028 ( .A(n51363), .B(n4583), .Z(n4584) );
  NAND U5029 ( .A(n51362), .B(n4584), .Z(n4585) );
  ANDN U5030 ( .B(n57926), .A(n57925), .Z(n4586) );
  NANDN U5031 ( .A(n57924), .B(n4585), .Z(n4587) );
  NAND U5032 ( .A(n4586), .B(n4587), .Z(n4588) );
  NAND U5033 ( .A(n51361), .B(n4588), .Z(n4589) );
  AND U5034 ( .A(n57928), .B(n4589), .Z(n4590) );
  NANDN U5035 ( .A(n57927), .B(n4590), .Z(n4591) );
  NAND U5036 ( .A(n57929), .B(n4591), .Z(n57930) );
  AND U5037 ( .A(n51352), .B(n51351), .Z(n4592) );
  NANDN U5038 ( .A(n57956), .B(n57955), .Z(n4593) );
  AND U5039 ( .A(n4592), .B(n4593), .Z(n4594) );
  AND U5040 ( .A(n57959), .B(n57958), .Z(n4595) );
  NANDN U5041 ( .A(n4594), .B(n57957), .Z(n4596) );
  AND U5042 ( .A(n4595), .B(n4596), .Z(n4597) );
  AND U5043 ( .A(n57962), .B(n57961), .Z(n4598) );
  OR U5044 ( .A(n57960), .B(n4597), .Z(n4599) );
  AND U5045 ( .A(n4598), .B(n4599), .Z(n4600) );
  ANDN U5046 ( .B(n57964), .A(n57965), .Z(n4601) );
  OR U5047 ( .A(n57963), .B(n4600), .Z(n4602) );
  AND U5048 ( .A(n4601), .B(n4602), .Z(n4603) );
  OR U5049 ( .A(n57966), .B(n4603), .Z(n4604) );
  NAND U5050 ( .A(n57967), .B(n4604), .Z(n4605) );
  NANDN U5051 ( .A(n57968), .B(n4605), .Z(n4606) );
  NAND U5052 ( .A(n57969), .B(n4606), .Z(n57970) );
  NOR U5053 ( .A(n57997), .B(n57998), .Z(n4607) );
  NAND U5054 ( .A(n57994), .B(n57995), .Z(n4608) );
  AND U5055 ( .A(n4607), .B(n4608), .Z(n4609) );
  ANDN U5056 ( .B(n58000), .A(n58001), .Z(n4610) );
  OR U5057 ( .A(n4609), .B(n57999), .Z(n4611) );
  NAND U5058 ( .A(n4610), .B(n4611), .Z(n4612) );
  NOR U5059 ( .A(n58003), .B(n58004), .Z(n4613) );
  NANDN U5060 ( .A(n58002), .B(n4612), .Z(n4614) );
  NAND U5061 ( .A(n4613), .B(n4614), .Z(n4615) );
  NANDN U5062 ( .A(n58005), .B(n4615), .Z(n4616) );
  NAND U5063 ( .A(n58006), .B(n4616), .Z(n4617) );
  ANDN U5064 ( .B(n4617), .A(n58007), .Z(n4618) );
  NANDN U5065 ( .A(n4618), .B(n58008), .Z(n4619) );
  NANDN U5066 ( .A(n58009), .B(n4619), .Z(n4620) );
  NAND U5067 ( .A(n58010), .B(n4620), .Z(n4621) );
  NAND U5068 ( .A(n58011), .B(n4621), .Z(n4622) );
  NANDN U5069 ( .A(n58012), .B(n4622), .Z(n4623) );
  AND U5070 ( .A(n58013), .B(n4623), .Z(n58014) );
  NAND U5071 ( .A(n58043), .B(n58044), .Z(n4624) );
  NAND U5072 ( .A(n58047), .B(n4624), .Z(n4625) );
  NANDN U5073 ( .A(n58048), .B(n4625), .Z(n4626) );
  AND U5074 ( .A(n58049), .B(n4626), .Z(n4627) );
  AND U5075 ( .A(n51336), .B(n51337), .Z(n4628) );
  OR U5076 ( .A(n4627), .B(n58050), .Z(n4629) );
  AND U5077 ( .A(n4628), .B(n4629), .Z(n4630) );
  OR U5078 ( .A(n4630), .B(n58051), .Z(n4631) );
  NAND U5079 ( .A(n58052), .B(n4631), .Z(n4632) );
  NAND U5080 ( .A(n58053), .B(n4632), .Z(n4633) );
  AND U5081 ( .A(n58054), .B(n58055), .Z(n4634) );
  NAND U5082 ( .A(n4633), .B(n4634), .Z(n4635) );
  NAND U5083 ( .A(n58056), .B(n4635), .Z(n4636) );
  AND U5084 ( .A(n51335), .B(n51334), .Z(n4637) );
  NAND U5085 ( .A(n4636), .B(n4637), .Z(n4638) );
  NAND U5086 ( .A(n58057), .B(n4638), .Z(n4639) );
  NANDN U5087 ( .A(n51333), .B(n4639), .Z(n58058) );
  NAND U5088 ( .A(n58091), .B(n58090), .Z(n4640) );
  AND U5089 ( .A(n58092), .B(n4640), .Z(n4641) );
  ANDN U5090 ( .B(n58094), .A(n4641), .Z(n4642) );
  NAND U5091 ( .A(n58093), .B(n4642), .Z(n4643) );
  NANDN U5092 ( .A(n58095), .B(n4643), .Z(n4644) );
  AND U5093 ( .A(n58097), .B(n58096), .Z(n4645) );
  NAND U5094 ( .A(n4644), .B(n4645), .Z(n4646) );
  NAND U5095 ( .A(n58098), .B(n4646), .Z(n4647) );
  AND U5096 ( .A(n58099), .B(n58100), .Z(n4648) );
  NAND U5097 ( .A(n4647), .B(n4648), .Z(n4649) );
  NAND U5098 ( .A(n58101), .B(n4649), .Z(n4650) );
  AND U5099 ( .A(n51323), .B(n51322), .Z(n4651) );
  NAND U5100 ( .A(n4650), .B(n4651), .Z(n4652) );
  NANDN U5101 ( .A(n58102), .B(n4652), .Z(n4653) );
  NAND U5102 ( .A(n58103), .B(n4653), .Z(n4654) );
  NANDN U5103 ( .A(n58104), .B(n4654), .Z(n4655) );
  AND U5104 ( .A(n58105), .B(n4655), .Z(n4656) );
  AND U5105 ( .A(n58106), .B(n4656), .Z(n58109) );
  NAND U5106 ( .A(n58132), .B(n58133), .Z(n4657) );
  NAND U5107 ( .A(n58136), .B(n4657), .Z(n4658) );
  NANDN U5108 ( .A(n58137), .B(n4658), .Z(n4659) );
  AND U5109 ( .A(n58139), .B(n58138), .Z(n4660) );
  NAND U5110 ( .A(n4659), .B(n4660), .Z(n4661) );
  NAND U5111 ( .A(n58140), .B(n4661), .Z(n4662) );
  ANDN U5112 ( .B(n58141), .A(n58142), .Z(n4663) );
  NAND U5113 ( .A(n4662), .B(n4663), .Z(n4664) );
  NAND U5114 ( .A(n58143), .B(n4664), .Z(n4665) );
  AND U5115 ( .A(n51310), .B(n51311), .Z(n4666) );
  NAND U5116 ( .A(n4665), .B(n4666), .Z(n4667) );
  NANDN U5117 ( .A(n58144), .B(n4667), .Z(n4668) );
  AND U5118 ( .A(n58145), .B(n58146), .Z(n4669) );
  NAND U5119 ( .A(n4668), .B(n4669), .Z(n4670) );
  NAND U5120 ( .A(n51309), .B(n4670), .Z(n58148) );
  AND U5121 ( .A(n51300), .B(n58178), .Z(n4671) );
  NANDN U5122 ( .A(n58177), .B(n58176), .Z(n4672) );
  AND U5123 ( .A(n4671), .B(n4672), .Z(n4673) );
  OR U5124 ( .A(n51299), .B(n4673), .Z(n4674) );
  NAND U5125 ( .A(n51298), .B(n4674), .Z(n4675) );
  NAND U5126 ( .A(n58179), .B(n4675), .Z(n4676) );
  AND U5127 ( .A(n58180), .B(n58181), .Z(n4677) );
  NAND U5128 ( .A(n4676), .B(n4677), .Z(n4678) );
  NAND U5129 ( .A(n51297), .B(n4678), .Z(n4679) );
  AND U5130 ( .A(n58183), .B(n58182), .Z(n4680) );
  NAND U5131 ( .A(n4679), .B(n4680), .Z(n4681) );
  NAND U5132 ( .A(n58184), .B(n4681), .Z(n4682) );
  AND U5133 ( .A(n58185), .B(n58186), .Z(n4683) );
  NAND U5134 ( .A(n4682), .B(n4683), .Z(n4684) );
  NANDN U5135 ( .A(n58187), .B(n4684), .Z(n58188) );
  NAND U5136 ( .A(n57661), .B(n17427), .Z(n4685) );
  NANDN U5137 ( .A(n51432), .B(n4685), .Z(n4686) );
  AND U5138 ( .A(n51431), .B(n4686), .Z(n4687) );
  AND U5139 ( .A(n43564), .B(n57664), .Z(n4688) );
  OR U5140 ( .A(n57662), .B(n4687), .Z(n4689) );
  AND U5141 ( .A(n4688), .B(n4689), .Z(n4690) );
  OR U5142 ( .A(n57665), .B(n4690), .Z(n4691) );
  NAND U5143 ( .A(n57666), .B(n4691), .Z(n4692) );
  NANDN U5144 ( .A(n51430), .B(n4692), .Z(n4693) );
  NAND U5145 ( .A(n51429), .B(n4693), .Z(n4694) );
  NANDN U5146 ( .A(n57669), .B(n4694), .Z(n4695) );
  AND U5147 ( .A(n57671), .B(n4695), .Z(n4696) );
  OR U5148 ( .A(n57672), .B(n4696), .Z(n4697) );
  AND U5149 ( .A(n57673), .B(n4697), .Z(n4698) );
  XNOR U5150 ( .A(x[5292]), .B(y[5292]), .Z(n4699) );
  AND U5151 ( .A(n4698), .B(n4699), .Z(n4700) );
  OR U5152 ( .A(n57675), .B(n4700), .Z(n4701) );
  NAND U5153 ( .A(n57676), .B(n4701), .Z(n4702) );
  NANDN U5154 ( .A(n57677), .B(n4702), .Z(n17429) );
  AND U5155 ( .A(n58212), .B(n58213), .Z(n4703) );
  AND U5156 ( .A(n51287), .B(n51288), .Z(n4704) );
  OR U5157 ( .A(n58214), .B(n4703), .Z(n4705) );
  AND U5158 ( .A(n4704), .B(n4705), .Z(n4706) );
  NANDN U5159 ( .A(n4706), .B(n58215), .Z(n4707) );
  NAND U5160 ( .A(n58216), .B(n4707), .Z(n4708) );
  NAND U5161 ( .A(n51286), .B(n4708), .Z(n4709) );
  AND U5162 ( .A(n58218), .B(n58217), .Z(n4710) );
  NAND U5163 ( .A(n4709), .B(n4710), .Z(n4711) );
  NAND U5164 ( .A(n58219), .B(n4711), .Z(n4712) );
  AND U5165 ( .A(n51285), .B(n51284), .Z(n4713) );
  NAND U5166 ( .A(n4712), .B(n4713), .Z(n4714) );
  NANDN U5167 ( .A(n58220), .B(n4714), .Z(n4715) );
  AND U5168 ( .A(n58222), .B(n58221), .Z(n4716) );
  NAND U5169 ( .A(n4715), .B(n4716), .Z(n4717) );
  NANDN U5170 ( .A(n58223), .B(n4717), .Z(n58224) );
  AND U5171 ( .A(n58249), .B(n58250), .Z(n4718) );
  NAND U5172 ( .A(n58251), .B(n4718), .Z(n4719) );
  NAND U5173 ( .A(n58252), .B(n4719), .Z(n4720) );
  AND U5174 ( .A(n51275), .B(n51276), .Z(n4721) );
  NAND U5175 ( .A(n4720), .B(n4721), .Z(n4722) );
  NAND U5176 ( .A(n58253), .B(n4722), .Z(n4723) );
  AND U5177 ( .A(n58255), .B(n58254), .Z(n4724) );
  NAND U5178 ( .A(n4723), .B(n4724), .Z(n4725) );
  NANDN U5179 ( .A(n58256), .B(n4725), .Z(n4726) );
  AND U5180 ( .A(n58258), .B(n58257), .Z(n4727) );
  NAND U5181 ( .A(n4726), .B(n4727), .Z(n4728) );
  NANDN U5182 ( .A(n58259), .B(n4728), .Z(n4729) );
  AND U5183 ( .A(n58261), .B(n58260), .Z(n4730) );
  NAND U5184 ( .A(n4729), .B(n4730), .Z(n4731) );
  NAND U5185 ( .A(n58262), .B(n4731), .Z(n4732) );
  AND U5186 ( .A(n51273), .B(n51274), .Z(n4733) );
  NAND U5187 ( .A(n4732), .B(n4733), .Z(n4734) );
  NAND U5188 ( .A(n58263), .B(n4734), .Z(n58264) );
  AND U5189 ( .A(n58351), .B(n58352), .Z(n4735) );
  NAND U5190 ( .A(n58350), .B(n51256), .Z(n4736) );
  AND U5191 ( .A(n4735), .B(n4736), .Z(n4737) );
  AND U5192 ( .A(n58355), .B(n58354), .Z(n4738) );
  OR U5193 ( .A(n58353), .B(n4737), .Z(n4739) );
  AND U5194 ( .A(n4738), .B(n4739), .Z(n4740) );
  AND U5195 ( .A(n51255), .B(n51254), .Z(n4741) );
  OR U5196 ( .A(n58356), .B(n4740), .Z(n4742) );
  AND U5197 ( .A(n4741), .B(n4742), .Z(n4743) );
  AND U5198 ( .A(n58359), .B(n58358), .Z(n4744) );
  NANDN U5199 ( .A(n4743), .B(n58357), .Z(n4745) );
  AND U5200 ( .A(n4744), .B(n4745), .Z(n4746) );
  AND U5201 ( .A(n58360), .B(n58361), .Z(n4747) );
  NANDN U5202 ( .A(n4746), .B(n51253), .Z(n4748) );
  AND U5203 ( .A(n4747), .B(n4748), .Z(n4749) );
  AND U5204 ( .A(n58363), .B(n58364), .Z(n4750) );
  OR U5205 ( .A(n58362), .B(n4749), .Z(n4751) );
  AND U5206 ( .A(n4750), .B(n4751), .Z(n58366) );
  ANDN U5207 ( .B(n58391), .A(n58390), .Z(n4752) );
  NANDN U5208 ( .A(n58389), .B(n58388), .Z(n4753) );
  NAND U5209 ( .A(n4752), .B(n4753), .Z(n4754) );
  NAND U5210 ( .A(n58392), .B(n4754), .Z(n4755) );
  AND U5211 ( .A(n58393), .B(n4755), .Z(n4756) );
  NAND U5212 ( .A(n4756), .B(n58394), .Z(n4757) );
  AND U5213 ( .A(n51243), .B(n51244), .Z(n4758) );
  NANDN U5214 ( .A(n58395), .B(n4757), .Z(n4759) );
  NAND U5215 ( .A(n4758), .B(n4759), .Z(n4760) );
  AND U5216 ( .A(n58397), .B(n58398), .Z(n4761) );
  NANDN U5217 ( .A(n58396), .B(n4760), .Z(n4762) );
  NAND U5218 ( .A(n4761), .B(n4762), .Z(n4763) );
  AND U5219 ( .A(n58401), .B(n58400), .Z(n4764) );
  NANDN U5220 ( .A(n58399), .B(n4763), .Z(n4765) );
  NAND U5221 ( .A(n4764), .B(n4765), .Z(n4766) );
  NAND U5222 ( .A(n58402), .B(n4766), .Z(n58404) );
  AND U5223 ( .A(n58440), .B(n58439), .Z(n4767) );
  OR U5224 ( .A(n58437), .B(n58438), .Z(n4768) );
  AND U5225 ( .A(n4767), .B(n4768), .Z(n4769) );
  AND U5226 ( .A(n51235), .B(n51236), .Z(n4770) );
  OR U5227 ( .A(n58441), .B(n4769), .Z(n4771) );
  AND U5228 ( .A(n4770), .B(n4771), .Z(n4772) );
  AND U5229 ( .A(n58444), .B(n58443), .Z(n4773) );
  OR U5230 ( .A(n58442), .B(n4772), .Z(n4774) );
  AND U5231 ( .A(n4773), .B(n4774), .Z(n4775) );
  OR U5232 ( .A(n58445), .B(n4775), .Z(n4776) );
  AND U5233 ( .A(n58446), .B(n4776), .Z(n4777) );
  OR U5234 ( .A(n51234), .B(n4777), .Z(n4778) );
  NAND U5235 ( .A(n51233), .B(n4778), .Z(n4779) );
  NAND U5236 ( .A(n58447), .B(n4779), .Z(n58449) );
  NAND U5237 ( .A(n58475), .B(n58474), .Z(n4780) );
  ANDN U5238 ( .B(n4780), .A(n58476), .Z(n4781) );
  NOR U5239 ( .A(n58478), .B(n4781), .Z(n4782) );
  NAND U5240 ( .A(n58479), .B(n4782), .Z(n4783) );
  NANDN U5241 ( .A(n58480), .B(n4783), .Z(n4784) );
  AND U5242 ( .A(n58482), .B(n58481), .Z(n4785) );
  NAND U5243 ( .A(n4784), .B(n4785), .Z(n4786) );
  NAND U5244 ( .A(n58483), .B(n4786), .Z(n4787) );
  AND U5245 ( .A(n58485), .B(n58484), .Z(n4788) );
  NAND U5246 ( .A(n4787), .B(n4788), .Z(n4789) );
  NAND U5247 ( .A(n58486), .B(n4789), .Z(n4790) );
  AND U5248 ( .A(n51225), .B(n51224), .Z(n4791) );
  NAND U5249 ( .A(n4790), .B(n4791), .Z(n4792) );
  NANDN U5250 ( .A(n58487), .B(n4792), .Z(n4793) );
  NAND U5251 ( .A(n58488), .B(n4793), .Z(n4794) );
  NANDN U5252 ( .A(n58489), .B(n4794), .Z(n4795) );
  AND U5253 ( .A(n58490), .B(n4795), .Z(n58492) );
  AND U5254 ( .A(n58508), .B(n58507), .Z(n58509) );
  AND U5255 ( .A(n51210), .B(n58538), .Z(n4796) );
  NAND U5256 ( .A(n51209), .B(n4796), .Z(n4797) );
  ANDN U5257 ( .B(n4797), .A(n58539), .Z(n4798) );
  ANDN U5258 ( .B(n58541), .A(n4798), .Z(n4799) );
  NAND U5259 ( .A(n58540), .B(n4799), .Z(n4800) );
  AND U5260 ( .A(n51208), .B(n4800), .Z(n4801) );
  ANDN U5261 ( .B(n58543), .A(n4801), .Z(n4802) );
  NAND U5262 ( .A(n58542), .B(n4802), .Z(n4803) );
  AND U5263 ( .A(n58544), .B(n4803), .Z(n4804) );
  ANDN U5264 ( .B(n58545), .A(n4804), .Z(n4805) );
  NAND U5265 ( .A(n58546), .B(n4805), .Z(n4806) );
  ANDN U5266 ( .B(n4806), .A(n58547), .Z(n4807) );
  ANDN U5267 ( .B(n51207), .A(n4807), .Z(n4808) );
  NAND U5268 ( .A(n51206), .B(n4808), .Z(n4809) );
  ANDN U5269 ( .B(n4809), .A(n58548), .Z(n58552) );
  NAND U5270 ( .A(n58577), .B(n58576), .Z(n4810) );
  AND U5271 ( .A(n58580), .B(n4810), .Z(n4811) );
  NANDN U5272 ( .A(n58579), .B(n4811), .Z(n4812) );
  AND U5273 ( .A(n58582), .B(n58583), .Z(n4813) );
  NANDN U5274 ( .A(n58581), .B(n4812), .Z(n4814) );
  NAND U5275 ( .A(n4813), .B(n4814), .Z(n4815) );
  AND U5276 ( .A(n58585), .B(n58586), .Z(n4816) );
  NANDN U5277 ( .A(n58584), .B(n4815), .Z(n4817) );
  NAND U5278 ( .A(n4816), .B(n4817), .Z(n4818) );
  NAND U5279 ( .A(n58587), .B(n4818), .Z(n4819) );
  AND U5280 ( .A(n51196), .B(n4819), .Z(n4820) );
  NAND U5281 ( .A(n4820), .B(n51197), .Z(n4821) );
  NAND U5282 ( .A(n58588), .B(n4821), .Z(n4822) );
  AND U5283 ( .A(n58589), .B(n4822), .Z(n4823) );
  NAND U5284 ( .A(n4823), .B(n58590), .Z(n4824) );
  AND U5285 ( .A(n51195), .B(n58592), .Z(n4825) );
  NANDN U5286 ( .A(n58591), .B(n4824), .Z(n4826) );
  NAND U5287 ( .A(n4825), .B(n4826), .Z(n58593) );
  NAND U5288 ( .A(n58627), .B(n58626), .Z(n4827) );
  NANDN U5289 ( .A(n58628), .B(n4827), .Z(n4828) );
  NAND U5290 ( .A(n58629), .B(n4828), .Z(n4829) );
  NAND U5291 ( .A(n58630), .B(n4829), .Z(n4830) );
  AND U5292 ( .A(n51187), .B(n4830), .Z(n4831) );
  NAND U5293 ( .A(n4831), .B(n51188), .Z(n4832) );
  NAND U5294 ( .A(n58631), .B(n4832), .Z(n4833) );
  AND U5295 ( .A(n58632), .B(n4833), .Z(n4834) );
  NAND U5296 ( .A(n4834), .B(n58633), .Z(n4835) );
  AND U5297 ( .A(n58635), .B(n58636), .Z(n4836) );
  NANDN U5298 ( .A(n58634), .B(n4835), .Z(n4837) );
  NAND U5299 ( .A(n4836), .B(n4837), .Z(n4838) );
  NAND U5300 ( .A(n58637), .B(n4838), .Z(n4839) );
  AND U5301 ( .A(n58639), .B(n4839), .Z(n4840) );
  NAND U5302 ( .A(n4840), .B(n58638), .Z(n4841) );
  NAND U5303 ( .A(n58640), .B(n4841), .Z(n58641) );
  NANDN U5304 ( .A(n58676), .B(n58675), .Z(n4842) );
  ANDN U5305 ( .B(n4842), .A(n58677), .Z(n4843) );
  ANDN U5306 ( .B(n58678), .A(n4843), .Z(n4844) );
  NAND U5307 ( .A(n58679), .B(n4844), .Z(n4845) );
  NANDN U5308 ( .A(n51175), .B(n4845), .Z(n4846) );
  AND U5309 ( .A(n58681), .B(n58680), .Z(n4847) );
  NAND U5310 ( .A(n4846), .B(n4847), .Z(n4848) );
  NAND U5311 ( .A(n58682), .B(n4848), .Z(n4849) );
  AND U5312 ( .A(n51174), .B(n51173), .Z(n4850) );
  NAND U5313 ( .A(n4849), .B(n4850), .Z(n4851) );
  NAND U5314 ( .A(n58683), .B(n4851), .Z(n4852) );
  AND U5315 ( .A(n58684), .B(n58685), .Z(n4853) );
  NAND U5316 ( .A(n4852), .B(n4853), .Z(n4854) );
  NANDN U5317 ( .A(n58686), .B(n4854), .Z(n4855) );
  AND U5318 ( .A(n58688), .B(n58687), .Z(n4856) );
  NAND U5319 ( .A(n4855), .B(n4856), .Z(n4857) );
  NANDN U5320 ( .A(n58689), .B(n4857), .Z(n58690) );
  NANDN U5321 ( .A(n58726), .B(n58725), .Z(n4858) );
  NANDN U5322 ( .A(n58727), .B(n4858), .Z(n4859) );
  ANDN U5323 ( .B(n4859), .A(n58728), .Z(n4860) );
  NAND U5324 ( .A(n4860), .B(n51166), .Z(n4861) );
  NAND U5325 ( .A(n58729), .B(n4861), .Z(n4862) );
  AND U5326 ( .A(n51165), .B(n4862), .Z(n4863) );
  ANDN U5327 ( .B(n58732), .A(n58731), .Z(n4864) );
  NANDN U5328 ( .A(n4863), .B(n58730), .Z(n4865) );
  AND U5329 ( .A(n4864), .B(n4865), .Z(n4866) );
  ANDN U5330 ( .B(n58734), .A(n58733), .Z(n4867) );
  NANDN U5331 ( .A(n4866), .B(n51164), .Z(n4868) );
  AND U5332 ( .A(n4867), .B(n4868), .Z(n4869) );
  ANDN U5333 ( .B(n58736), .A(n58737), .Z(n4870) );
  OR U5334 ( .A(n58735), .B(n4869), .Z(n4871) );
  AND U5335 ( .A(n4870), .B(n4871), .Z(n58738) );
  NAND U5336 ( .A(n51150), .B(n58780), .Z(n4872) );
  AND U5337 ( .A(n58781), .B(n4872), .Z(n4873) );
  NANDN U5338 ( .A(n58782), .B(n4873), .Z(n4874) );
  ANDN U5339 ( .B(n58785), .A(n58784), .Z(n4875) );
  NANDN U5340 ( .A(n58783), .B(n4874), .Z(n4876) );
  NAND U5341 ( .A(n4875), .B(n4876), .Z(n4877) );
  ANDN U5342 ( .B(n51149), .A(n51148), .Z(n4878) );
  NANDN U5343 ( .A(n58786), .B(n4877), .Z(n4879) );
  NAND U5344 ( .A(n4878), .B(n4879), .Z(n4880) );
  NAND U5345 ( .A(n58787), .B(n4880), .Z(n4881) );
  AND U5346 ( .A(n58788), .B(n4881), .Z(n4882) );
  NANDN U5347 ( .A(n58789), .B(n4882), .Z(n4883) );
  NAND U5348 ( .A(n51147), .B(n4883), .Z(n4884) );
  AND U5349 ( .A(n58790), .B(n4884), .Z(n4885) );
  NANDN U5350 ( .A(n58791), .B(n4885), .Z(n58792) );
  NAND U5351 ( .A(n58830), .B(n58831), .Z(n4886) );
  NAND U5352 ( .A(n58832), .B(n4886), .Z(n4887) );
  AND U5353 ( .A(n58834), .B(n4887), .Z(n4888) );
  NANDN U5354 ( .A(n58833), .B(n4888), .Z(n4889) );
  NAND U5355 ( .A(n51130), .B(n4889), .Z(n4890) );
  AND U5356 ( .A(n58836), .B(n4890), .Z(n4891) );
  NANDN U5357 ( .A(n58835), .B(n4891), .Z(n4892) );
  ANDN U5358 ( .B(n58838), .A(n58839), .Z(n4893) );
  NANDN U5359 ( .A(n58837), .B(n4892), .Z(n4894) );
  NAND U5360 ( .A(n4893), .B(n4894), .Z(n4895) );
  ANDN U5361 ( .B(n51129), .A(n51128), .Z(n4896) );
  NANDN U5362 ( .A(n58840), .B(n4895), .Z(n4897) );
  NAND U5363 ( .A(n4896), .B(n4897), .Z(n4898) );
  AND U5364 ( .A(n58843), .B(n58842), .Z(n4899) );
  NANDN U5365 ( .A(n58841), .B(n4898), .Z(n4900) );
  NAND U5366 ( .A(n4899), .B(n4900), .Z(n58844) );
  AND U5367 ( .A(n58870), .B(n58869), .Z(n58871) );
  ANDN U5368 ( .B(n58898), .A(n58897), .Z(n4901) );
  NAND U5369 ( .A(n58896), .B(n58895), .Z(n4902) );
  AND U5370 ( .A(n4901), .B(n4902), .Z(n4903) );
  ANDN U5371 ( .B(n58901), .A(n58900), .Z(n4904) );
  OR U5372 ( .A(n4903), .B(n58899), .Z(n4905) );
  AND U5373 ( .A(n4904), .B(n4905), .Z(n4906) );
  AND U5374 ( .A(n58903), .B(n58904), .Z(n4907) );
  OR U5375 ( .A(n58902), .B(n4906), .Z(n4908) );
  AND U5376 ( .A(n4907), .B(n4908), .Z(n4909) );
  AND U5377 ( .A(n51111), .B(n51112), .Z(n4910) );
  NANDN U5378 ( .A(n4909), .B(n58905), .Z(n4911) );
  AND U5379 ( .A(n4910), .B(n4911), .Z(n4912) );
  AND U5380 ( .A(n58908), .B(n58907), .Z(n4913) );
  NANDN U5381 ( .A(n4912), .B(n58906), .Z(n4914) );
  AND U5382 ( .A(n4913), .B(n4914), .Z(n4915) );
  AND U5383 ( .A(n58911), .B(n58910), .Z(n4916) );
  OR U5384 ( .A(n4915), .B(n58909), .Z(n4917) );
  AND U5385 ( .A(n4916), .B(n4917), .Z(n58913) );
  ANDN U5386 ( .B(n51108), .A(n51107), .Z(n58928) );
  NANDN U5387 ( .A(n58958), .B(n58957), .Z(n4918) );
  NAND U5388 ( .A(n58959), .B(n4918), .Z(n4919) );
  NANDN U5389 ( .A(n58960), .B(n4919), .Z(n4920) );
  NAND U5390 ( .A(n58961), .B(n4920), .Z(n4921) );
  NANDN U5391 ( .A(n58962), .B(n4921), .Z(n4922) );
  AND U5392 ( .A(n58963), .B(n4922), .Z(n4923) );
  OR U5393 ( .A(n4923), .B(n58964), .Z(n4924) );
  NAND U5394 ( .A(n58965), .B(n4924), .Z(n4925) );
  ANDN U5395 ( .B(n4925), .A(n58966), .Z(n4926) );
  ANDN U5396 ( .B(n51099), .A(n4926), .Z(n4927) );
  NAND U5397 ( .A(n51098), .B(n4927), .Z(n4928) );
  ANDN U5398 ( .B(n4928), .A(n58967), .Z(n4929) );
  NANDN U5399 ( .A(n4929), .B(n58968), .Z(n4930) );
  NANDN U5400 ( .A(n58969), .B(n4930), .Z(n4931) );
  NAND U5401 ( .A(n58970), .B(n4931), .Z(n4932) );
  NANDN U5402 ( .A(n51097), .B(n4932), .Z(n58971) );
  NAND U5403 ( .A(n59006), .B(n59005), .Z(n4933) );
  NAND U5404 ( .A(n59007), .B(n4933), .Z(n4934) );
  ANDN U5405 ( .B(n4934), .A(n51088), .Z(n4935) );
  AND U5406 ( .A(n59009), .B(n59008), .Z(n4936) );
  NANDN U5407 ( .A(n4935), .B(n51087), .Z(n4937) );
  AND U5408 ( .A(n4936), .B(n4937), .Z(n4938) );
  ANDN U5409 ( .B(n51086), .A(n51085), .Z(n4939) );
  OR U5410 ( .A(n4938), .B(n59010), .Z(n4940) );
  NAND U5411 ( .A(n4939), .B(n4940), .Z(n4941) );
  ANDN U5412 ( .B(n59012), .A(n59013), .Z(n4942) );
  NANDN U5413 ( .A(n59011), .B(n4941), .Z(n4943) );
  NAND U5414 ( .A(n4942), .B(n4943), .Z(n4944) );
  NAND U5415 ( .A(n51084), .B(n4944), .Z(n59016) );
  NAND U5416 ( .A(n59059), .B(n59058), .Z(n4945) );
  NANDN U5417 ( .A(n59061), .B(n4945), .Z(n4946) );
  AND U5418 ( .A(n59062), .B(n4946), .Z(n4947) );
  ANDN U5419 ( .B(n4947), .A(n59063), .Z(n4948) );
  ANDN U5420 ( .B(n51071), .A(n51070), .Z(n4949) );
  OR U5421 ( .A(n4948), .B(n59064), .Z(n4950) );
  AND U5422 ( .A(n4949), .B(n4950), .Z(n4951) );
  AND U5423 ( .A(n59067), .B(n59066), .Z(n4952) );
  OR U5424 ( .A(n59065), .B(n4951), .Z(n4953) );
  AND U5425 ( .A(n4952), .B(n4953), .Z(n4954) );
  AND U5426 ( .A(n59068), .B(n59069), .Z(n4955) );
  NANDN U5427 ( .A(n4954), .B(n51069), .Z(n4956) );
  AND U5428 ( .A(n4955), .B(n4956), .Z(n4957) );
  AND U5429 ( .A(n59071), .B(n59072), .Z(n4958) );
  NANDN U5430 ( .A(n4957), .B(n59070), .Z(n4959) );
  AND U5431 ( .A(n4958), .B(n4959), .Z(n59073) );
  NAND U5432 ( .A(n59101), .B(n59100), .Z(n4960) );
  ANDN U5433 ( .B(n4960), .A(n59102), .Z(n4961) );
  NOR U5434 ( .A(n59104), .B(n4961), .Z(n4962) );
  NAND U5435 ( .A(n59105), .B(n4962), .Z(n4963) );
  AND U5436 ( .A(n59106), .B(n4963), .Z(n4964) );
  OR U5437 ( .A(n59107), .B(n4964), .Z(n4965) );
  NAND U5438 ( .A(n59108), .B(n4965), .Z(n4966) );
  NANDN U5439 ( .A(n59109), .B(n4966), .Z(n4967) );
  NAND U5440 ( .A(n59110), .B(n4967), .Z(n4968) );
  AND U5441 ( .A(n59111), .B(n4968), .Z(n4969) );
  NAND U5442 ( .A(n4969), .B(n59112), .Z(n4970) );
  AND U5443 ( .A(n59114), .B(n59115), .Z(n4971) );
  NANDN U5444 ( .A(n59113), .B(n4970), .Z(n4972) );
  NAND U5445 ( .A(n4971), .B(n4972), .Z(n4973) );
  AND U5446 ( .A(n59118), .B(n59117), .Z(n4974) );
  NANDN U5447 ( .A(n59116), .B(n4973), .Z(n4975) );
  NAND U5448 ( .A(n4974), .B(n4975), .Z(n4976) );
  NAND U5449 ( .A(n59119), .B(n4976), .Z(n59120) );
  NAND U5450 ( .A(n59189), .B(n59188), .Z(n4977) );
  ANDN U5451 ( .B(n4977), .A(n59190), .Z(n4978) );
  ANDN U5452 ( .B(n59192), .A(n4978), .Z(n4979) );
  NAND U5453 ( .A(n59191), .B(n4979), .Z(n4980) );
  NAND U5454 ( .A(n59193), .B(n4980), .Z(n4981) );
  AND U5455 ( .A(n51049), .B(n51048), .Z(n4982) );
  NAND U5456 ( .A(n4981), .B(n4982), .Z(n4983) );
  NANDN U5457 ( .A(n59194), .B(n4983), .Z(n4984) );
  AND U5458 ( .A(n59195), .B(n59196), .Z(n4985) );
  NAND U5459 ( .A(n4984), .B(n4985), .Z(n4986) );
  NAND U5460 ( .A(n59197), .B(n4986), .Z(n4987) );
  AND U5461 ( .A(n59199), .B(n59198), .Z(n4988) );
  NAND U5462 ( .A(n4987), .B(n4988), .Z(n4989) );
  NAND U5463 ( .A(n59200), .B(n4989), .Z(n4990) );
  AND U5464 ( .A(n59202), .B(n59201), .Z(n4991) );
  NAND U5465 ( .A(n4990), .B(n4991), .Z(n4992) );
  NAND U5466 ( .A(n59203), .B(n4992), .Z(n59204) );
  NAND U5467 ( .A(n59235), .B(n51038), .Z(n4993) );
  AND U5468 ( .A(n59236), .B(n4993), .Z(n4994) );
  NAND U5469 ( .A(n4994), .B(n59237), .Z(n4995) );
  NAND U5470 ( .A(n59238), .B(n4995), .Z(n4996) );
  AND U5471 ( .A(n59240), .B(n4996), .Z(n4997) );
  NAND U5472 ( .A(n4997), .B(n59239), .Z(n4998) );
  AND U5473 ( .A(n51037), .B(n51036), .Z(n4999) );
  NANDN U5474 ( .A(n59241), .B(n4998), .Z(n5000) );
  NAND U5475 ( .A(n4999), .B(n5000), .Z(n5001) );
  ANDN U5476 ( .B(n59244), .A(n59243), .Z(n5002) );
  NANDN U5477 ( .A(n59242), .B(n5001), .Z(n5003) );
  NAND U5478 ( .A(n5002), .B(n5003), .Z(n5004) );
  NAND U5479 ( .A(n51035), .B(n5004), .Z(n5005) );
  AND U5480 ( .A(n51034), .B(n5005), .Z(n5006) );
  NAND U5481 ( .A(n5006), .B(n59245), .Z(n5007) );
  NAND U5482 ( .A(n59246), .B(n5007), .Z(n59247) );
  NAND U5483 ( .A(n59279), .B(n59278), .Z(n5008) );
  AND U5484 ( .A(n59280), .B(n5008), .Z(n5009) );
  ANDN U5485 ( .B(n59282), .A(n5009), .Z(n5010) );
  NAND U5486 ( .A(n59281), .B(n5010), .Z(n5011) );
  NAND U5487 ( .A(n59283), .B(n5011), .Z(n5012) );
  AND U5488 ( .A(n51027), .B(n51028), .Z(n5013) );
  NAND U5489 ( .A(n5012), .B(n5013), .Z(n5014) );
  NAND U5490 ( .A(n59284), .B(n5014), .Z(n5015) );
  AND U5491 ( .A(n59285), .B(n59286), .Z(n5016) );
  NAND U5492 ( .A(n5015), .B(n5016), .Z(n5017) );
  NANDN U5493 ( .A(n59287), .B(n5017), .Z(n5018) );
  AND U5494 ( .A(n59289), .B(n59288), .Z(n5019) );
  NAND U5495 ( .A(n5018), .B(n5019), .Z(n5020) );
  NAND U5496 ( .A(n59290), .B(n5020), .Z(n5021) );
  AND U5497 ( .A(n59292), .B(n59291), .Z(n5022) );
  NAND U5498 ( .A(n5021), .B(n5022), .Z(n5023) );
  NANDN U5499 ( .A(n59293), .B(n5023), .Z(n59294) );
  AND U5500 ( .A(n59327), .B(n59326), .Z(n5024) );
  NAND U5501 ( .A(n59328), .B(n5024), .Z(n5025) );
  AND U5502 ( .A(n59329), .B(n5025), .Z(n5026) );
  NOR U5503 ( .A(n5026), .B(n51018), .Z(n5027) );
  NAND U5504 ( .A(n51019), .B(n5027), .Z(n5028) );
  NAND U5505 ( .A(n59330), .B(n5028), .Z(n5029) );
  ANDN U5506 ( .B(n59331), .A(n59332), .Z(n5030) );
  NAND U5507 ( .A(n5029), .B(n5030), .Z(n5031) );
  NAND U5508 ( .A(n59333), .B(n5031), .Z(n5032) );
  ANDN U5509 ( .B(n51017), .A(n51016), .Z(n5033) );
  NAND U5510 ( .A(n5032), .B(n5033), .Z(n5034) );
  NAND U5511 ( .A(n51015), .B(n5034), .Z(n5035) );
  AND U5512 ( .A(n59335), .B(n59334), .Z(n5036) );
  NAND U5513 ( .A(n5035), .B(n5036), .Z(n5037) );
  NAND U5514 ( .A(n59336), .B(n5037), .Z(n5038) );
  ANDN U5515 ( .B(n5038), .A(n59337), .Z(n5039) );
  NAND U5516 ( .A(n59338), .B(n5039), .Z(n59339) );
  ANDN U5517 ( .B(n59371), .A(n59370), .Z(n5040) );
  NANDN U5518 ( .A(n59369), .B(n59368), .Z(n5041) );
  AND U5519 ( .A(n5040), .B(n5041), .Z(n5042) );
  ANDN U5520 ( .B(n51007), .A(n51006), .Z(n5043) );
  NANDN U5521 ( .A(n5042), .B(n59372), .Z(n5044) );
  AND U5522 ( .A(n5043), .B(n5044), .Z(n5045) );
  OR U5523 ( .A(n51005), .B(n5045), .Z(n5046) );
  NAND U5524 ( .A(n59373), .B(n5046), .Z(n5047) );
  NAND U5525 ( .A(n59374), .B(n5047), .Z(n5048) );
  NAND U5526 ( .A(n59375), .B(n5048), .Z(n5049) );
  NAND U5527 ( .A(n59376), .B(n5049), .Z(n5050) );
  AND U5528 ( .A(n59377), .B(n5050), .Z(n5051) );
  AND U5529 ( .A(n59380), .B(n59379), .Z(n5052) );
  OR U5530 ( .A(n59378), .B(n5051), .Z(n5053) );
  AND U5531 ( .A(n5052), .B(n5053), .Z(n5054) );
  ANDN U5532 ( .B(n59383), .A(n59382), .Z(n5055) );
  NANDN U5533 ( .A(n5054), .B(n59381), .Z(n5056) );
  AND U5534 ( .A(n5055), .B(n5056), .Z(n59386) );
  AND U5535 ( .A(n59424), .B(n59425), .Z(n5057) );
  AND U5536 ( .A(n59428), .B(n59427), .Z(n5058) );
  OR U5537 ( .A(n59426), .B(n5057), .Z(n5059) );
  AND U5538 ( .A(n5058), .B(n5059), .Z(n5060) );
  AND U5539 ( .A(n59429), .B(n59430), .Z(n5061) );
  NANDN U5540 ( .A(n5060), .B(n50984), .Z(n5062) );
  AND U5541 ( .A(n5061), .B(n5062), .Z(n5063) );
  ANDN U5542 ( .B(n59433), .A(n59432), .Z(n5064) );
  NANDN U5543 ( .A(n5063), .B(n59431), .Z(n5065) );
  AND U5544 ( .A(n5064), .B(n5065), .Z(n5066) );
  AND U5545 ( .A(n59436), .B(n59435), .Z(n5067) );
  NANDN U5546 ( .A(n5066), .B(n59434), .Z(n5068) );
  AND U5547 ( .A(n5067), .B(n5068), .Z(n5069) );
  ANDN U5548 ( .B(n59439), .A(n59438), .Z(n5070) );
  NANDN U5549 ( .A(n5069), .B(n59437), .Z(n5071) );
  AND U5550 ( .A(n5070), .B(n5071), .Z(n59441) );
  NOR U5551 ( .A(n50975), .B(n50974), .Z(n5072) );
  NAND U5552 ( .A(n59470), .B(n5072), .Z(n5073) );
  ANDN U5553 ( .B(n5073), .A(n50972), .Z(n5074) );
  NOR U5554 ( .A(n59471), .B(n5074), .Z(n5075) );
  NAND U5555 ( .A(n59472), .B(n5075), .Z(n5076) );
  AND U5556 ( .A(n59473), .B(n5076), .Z(n5077) );
  NANDN U5557 ( .A(n5077), .B(n59474), .Z(n5078) );
  ANDN U5558 ( .B(n5078), .A(n59475), .Z(n5079) );
  ANDN U5559 ( .B(n59477), .A(n5079), .Z(n5080) );
  NAND U5560 ( .A(n59476), .B(n5080), .Z(n5081) );
  NAND U5561 ( .A(n59478), .B(n5081), .Z(n5082) );
  AND U5562 ( .A(n59479), .B(n59480), .Z(n5083) );
  NAND U5563 ( .A(n5082), .B(n5083), .Z(n5084) );
  NANDN U5564 ( .A(n59481), .B(n5084), .Z(n5085) );
  ANDN U5565 ( .B(n50971), .A(n50970), .Z(n5086) );
  NAND U5566 ( .A(n5085), .B(n5086), .Z(n5087) );
  NAND U5567 ( .A(n59482), .B(n5087), .Z(n5088) );
  AND U5568 ( .A(n59483), .B(n5088), .Z(n59485) );
  ANDN U5569 ( .B(n59517), .A(n59518), .Z(n5089) );
  NAND U5570 ( .A(n59516), .B(n59515), .Z(n5090) );
  AND U5571 ( .A(n5089), .B(n5090), .Z(n5091) );
  ANDN U5572 ( .B(n50964), .A(n50963), .Z(n5092) );
  OR U5573 ( .A(n5091), .B(n59519), .Z(n5093) );
  NAND U5574 ( .A(n5092), .B(n5093), .Z(n5094) );
  AND U5575 ( .A(n59522), .B(n59521), .Z(n5095) );
  NANDN U5576 ( .A(n59520), .B(n5094), .Z(n5096) );
  NAND U5577 ( .A(n5095), .B(n5096), .Z(n5097) );
  NAND U5578 ( .A(n59523), .B(n5097), .Z(n5098) );
  AND U5579 ( .A(n59524), .B(n5098), .Z(n5099) );
  NAND U5580 ( .A(n5099), .B(n59525), .Z(n5100) );
  AND U5581 ( .A(n59527), .B(n59528), .Z(n5101) );
  NANDN U5582 ( .A(n59526), .B(n5100), .Z(n5102) );
  NAND U5583 ( .A(n5101), .B(n5102), .Z(n5103) );
  NAND U5584 ( .A(n59529), .B(n5103), .Z(n5104) );
  AND U5585 ( .A(n59531), .B(n5104), .Z(n5105) );
  NANDN U5586 ( .A(n59530), .B(n5105), .Z(n5106) );
  NAND U5587 ( .A(n59532), .B(n5106), .Z(n59533) );
  NAND U5588 ( .A(n59563), .B(n59562), .Z(n5107) );
  NANDN U5589 ( .A(n59564), .B(n5107), .Z(n5108) );
  AND U5590 ( .A(n59565), .B(n5108), .Z(n5109) );
  NAND U5591 ( .A(n5109), .B(n59566), .Z(n5110) );
  NAND U5592 ( .A(n59567), .B(n5110), .Z(n5111) );
  AND U5593 ( .A(n59568), .B(n5111), .Z(n5112) );
  NANDN U5594 ( .A(n5112), .B(n59569), .Z(n5113) );
  NAND U5595 ( .A(n59570), .B(n5113), .Z(n5114) );
  NANDN U5596 ( .A(n50953), .B(n5114), .Z(n5115) );
  ANDN U5597 ( .B(n59572), .A(n59571), .Z(n5116) );
  NAND U5598 ( .A(n5115), .B(n5116), .Z(n5117) );
  NAND U5599 ( .A(n59573), .B(n5117), .Z(n5118) );
  ANDN U5600 ( .B(n59574), .A(n59575), .Z(n5119) );
  NAND U5601 ( .A(n5118), .B(n5119), .Z(n5120) );
  NANDN U5602 ( .A(n59576), .B(n5120), .Z(n5121) );
  ANDN U5603 ( .B(n59578), .A(n59577), .Z(n5122) );
  NAND U5604 ( .A(n5121), .B(n5122), .Z(n5123) );
  NAND U5605 ( .A(n59579), .B(n5123), .Z(n59580) );
  OR U5606 ( .A(n59611), .B(n59612), .Z(n5124) );
  ANDN U5607 ( .B(n5124), .A(n50944), .Z(n5125) );
  NOR U5608 ( .A(n50943), .B(n5125), .Z(n5126) );
  NAND U5609 ( .A(n50942), .B(n5126), .Z(n5127) );
  NAND U5610 ( .A(n59613), .B(n5127), .Z(n5128) );
  AND U5611 ( .A(n59614), .B(n59615), .Z(n5129) );
  NAND U5612 ( .A(n5128), .B(n5129), .Z(n5130) );
  NANDN U5613 ( .A(n59616), .B(n5130), .Z(n5131) );
  AND U5614 ( .A(n50941), .B(n50940), .Z(n5132) );
  NAND U5615 ( .A(n5131), .B(n5132), .Z(n5133) );
  NAND U5616 ( .A(n50939), .B(n5133), .Z(n5134) );
  AND U5617 ( .A(n59618), .B(n59617), .Z(n5135) );
  NAND U5618 ( .A(n5134), .B(n5135), .Z(n5136) );
  NAND U5619 ( .A(n59619), .B(n5136), .Z(n5137) );
  ANDN U5620 ( .B(n59621), .A(n59620), .Z(n5138) );
  NAND U5621 ( .A(n5137), .B(n5138), .Z(n5139) );
  NAND U5622 ( .A(n59622), .B(n5139), .Z(n5140) );
  AND U5623 ( .A(n59623), .B(n5140), .Z(n59625) );
  NAND U5624 ( .A(n59654), .B(n59655), .Z(n5141) );
  AND U5625 ( .A(n59656), .B(n5141), .Z(n5142) );
  NAND U5626 ( .A(n5142), .B(n59657), .Z(n5143) );
  AND U5627 ( .A(n59660), .B(n59659), .Z(n5144) );
  NANDN U5628 ( .A(n59658), .B(n5143), .Z(n5145) );
  NAND U5629 ( .A(n5144), .B(n5145), .Z(n5146) );
  NAND U5630 ( .A(n59661), .B(n5146), .Z(n5147) );
  AND U5631 ( .A(n59663), .B(n5147), .Z(n5148) );
  NANDN U5632 ( .A(n59662), .B(n5148), .Z(n5149) );
  NOR U5633 ( .A(n50930), .B(n50929), .Z(n5150) );
  NANDN U5634 ( .A(n59664), .B(n5149), .Z(n5151) );
  NAND U5635 ( .A(n5150), .B(n5151), .Z(n5152) );
  NAND U5636 ( .A(n59665), .B(n5152), .Z(n5153) );
  AND U5637 ( .A(n59667), .B(n5153), .Z(n5154) );
  NANDN U5638 ( .A(n59666), .B(n5154), .Z(n5155) );
  NAND U5639 ( .A(n59668), .B(n5155), .Z(n5156) );
  AND U5640 ( .A(n50928), .B(n5156), .Z(n5157) );
  NAND U5641 ( .A(n5157), .B(n50927), .Z(n59669) );
  NAND U5642 ( .A(n59702), .B(n59701), .Z(n5158) );
  AND U5643 ( .A(n59703), .B(n5158), .Z(n5159) );
  NOR U5644 ( .A(n50918), .B(n5159), .Z(n5160) );
  NAND U5645 ( .A(n50919), .B(n5160), .Z(n5161) );
  NANDN U5646 ( .A(n59704), .B(n5161), .Z(n5162) );
  ANDN U5647 ( .B(n59705), .A(n59706), .Z(n5163) );
  NAND U5648 ( .A(n5162), .B(n5163), .Z(n5164) );
  NANDN U5649 ( .A(n59707), .B(n5164), .Z(n5165) );
  ANDN U5650 ( .B(n59709), .A(n59708), .Z(n5166) );
  NAND U5651 ( .A(n5165), .B(n5166), .Z(n5167) );
  NAND U5652 ( .A(n59710), .B(n5167), .Z(n5168) );
  AND U5653 ( .A(n59712), .B(n59711), .Z(n5169) );
  NAND U5654 ( .A(n5168), .B(n5169), .Z(n5170) );
  NAND U5655 ( .A(n59713), .B(n5170), .Z(n5171) );
  ANDN U5656 ( .B(n59715), .A(n59714), .Z(n5172) );
  NAND U5657 ( .A(n5171), .B(n5172), .Z(n5173) );
  NAND U5658 ( .A(n59716), .B(n5173), .Z(n59717) );
  NAND U5659 ( .A(n59749), .B(n59748), .Z(n5174) );
  AND U5660 ( .A(n59750), .B(n5174), .Z(n5175) );
  NOR U5661 ( .A(n59751), .B(n5175), .Z(n5176) );
  NAND U5662 ( .A(n59752), .B(n5176), .Z(n5177) );
  NAND U5663 ( .A(n59753), .B(n5177), .Z(n5178) );
  ANDN U5664 ( .B(n50907), .A(n50908), .Z(n5179) );
  NAND U5665 ( .A(n5178), .B(n5179), .Z(n5180) );
  NAND U5666 ( .A(n59754), .B(n5180), .Z(n5181) );
  ANDN U5667 ( .B(n59756), .A(n59755), .Z(n5182) );
  NAND U5668 ( .A(n5181), .B(n5182), .Z(n5183) );
  NAND U5669 ( .A(n59757), .B(n5183), .Z(n5184) );
  NAND U5670 ( .A(n59758), .B(n5184), .Z(n5185) );
  NANDN U5671 ( .A(n59759), .B(n5185), .Z(n5186) );
  ANDN U5672 ( .B(n5186), .A(n59760), .Z(n5187) );
  NAND U5673 ( .A(n59761), .B(n5187), .Z(n5188) );
  NAND U5674 ( .A(n59762), .B(n5188), .Z(n5189) );
  AND U5675 ( .A(n50906), .B(n5189), .Z(n5190) );
  NANDN U5676 ( .A(n50905), .B(n5190), .Z(n59763) );
  NAND U5677 ( .A(n59792), .B(n59791), .Z(n5191) );
  ANDN U5678 ( .B(n5191), .A(n59793), .Z(n5192) );
  NOR U5679 ( .A(n59794), .B(n5192), .Z(n5193) );
  NAND U5680 ( .A(n59795), .B(n5193), .Z(n5194) );
  NAND U5681 ( .A(n59796), .B(n5194), .Z(n5195) );
  AND U5682 ( .A(n59798), .B(n59797), .Z(n5196) );
  NAND U5683 ( .A(n5195), .B(n5196), .Z(n5197) );
  NAND U5684 ( .A(n59799), .B(n5197), .Z(n5198) );
  ANDN U5685 ( .B(n50894), .A(n50893), .Z(n5199) );
  NAND U5686 ( .A(n5198), .B(n5199), .Z(n5200) );
  NAND U5687 ( .A(n59800), .B(n5200), .Z(n5201) );
  ANDN U5688 ( .B(n59801), .A(n59802), .Z(n5202) );
  NAND U5689 ( .A(n5201), .B(n5202), .Z(n5203) );
  NANDN U5690 ( .A(n59803), .B(n5203), .Z(n5204) );
  ANDN U5691 ( .B(n50892), .A(n50891), .Z(n5205) );
  NAND U5692 ( .A(n5204), .B(n5205), .Z(n5206) );
  NANDN U5693 ( .A(n59804), .B(n5206), .Z(n59805) );
  ANDN U5694 ( .B(n50878), .A(n50877), .Z(n5207) );
  AND U5695 ( .A(n50883), .B(n50884), .Z(n5208) );
  NAND U5696 ( .A(n59838), .B(n5208), .Z(n5209) );
  NAND U5697 ( .A(n50881), .B(n5209), .Z(n5210) );
  ANDN U5698 ( .B(n59840), .A(n59839), .Z(n5211) );
  NAND U5699 ( .A(n5210), .B(n5211), .Z(n5212) );
  NAND U5700 ( .A(n59841), .B(n5212), .Z(n5213) );
  ANDN U5701 ( .B(n59842), .A(n50880), .Z(n5214) );
  NAND U5702 ( .A(n5213), .B(n5214), .Z(n5215) );
  NAND U5703 ( .A(n50879), .B(n5215), .Z(n5216) );
  ANDN U5704 ( .B(n59844), .A(n59843), .Z(n5217) );
  NAND U5705 ( .A(n5216), .B(n5217), .Z(n5218) );
  NAND U5706 ( .A(n59845), .B(n5218), .Z(n5219) );
  AND U5707 ( .A(n59847), .B(n59846), .Z(n5220) );
  NAND U5708 ( .A(n5219), .B(n5220), .Z(n5221) );
  NAND U5709 ( .A(n59848), .B(n5221), .Z(n5222) );
  NAND U5710 ( .A(n5207), .B(n5222), .Z(n59849) );
  ANDN U5711 ( .B(n59878), .A(n59877), .Z(n5223) );
  NAND U5712 ( .A(n59876), .B(n50869), .Z(n5224) );
  AND U5713 ( .A(n5223), .B(n5224), .Z(n5225) );
  AND U5714 ( .A(n59881), .B(n59880), .Z(n5226) );
  NANDN U5715 ( .A(n5225), .B(n59879), .Z(n5227) );
  AND U5716 ( .A(n5226), .B(n5227), .Z(n5228) );
  NANDN U5717 ( .A(n5228), .B(n59882), .Z(n5229) );
  AND U5718 ( .A(n59883), .B(n5229), .Z(n5230) );
  AND U5719 ( .A(n59886), .B(n59885), .Z(n5231) );
  NANDN U5720 ( .A(n5230), .B(n59884), .Z(n5232) );
  AND U5721 ( .A(n5231), .B(n5232), .Z(n5233) );
  AND U5722 ( .A(n50868), .B(n50867), .Z(n5234) );
  NANDN U5723 ( .A(n5233), .B(n59887), .Z(n5235) );
  AND U5724 ( .A(n5234), .B(n5235), .Z(n5236) );
  AND U5725 ( .A(n59889), .B(n59890), .Z(n5237) );
  OR U5726 ( .A(n5236), .B(n59888), .Z(n5238) );
  NAND U5727 ( .A(n5237), .B(n5238), .Z(n59891) );
  AND U5728 ( .A(n59919), .B(n59920), .Z(n5239) );
  NAND U5729 ( .A(n59921), .B(n5239), .Z(n5240) );
  NAND U5730 ( .A(n59922), .B(n5240), .Z(n5241) );
  ANDN U5731 ( .B(n59924), .A(n59923), .Z(n5242) );
  NAND U5732 ( .A(n5241), .B(n5242), .Z(n5243) );
  NANDN U5733 ( .A(n50858), .B(n5243), .Z(n5244) );
  AND U5734 ( .A(n59926), .B(n59925), .Z(n5245) );
  NAND U5735 ( .A(n5244), .B(n5245), .Z(n5246) );
  NAND U5736 ( .A(n59927), .B(n5246), .Z(n5247) );
  AND U5737 ( .A(n59928), .B(n5247), .Z(n5248) );
  ANDN U5738 ( .B(n50857), .A(n50856), .Z(n5249) );
  NANDN U5739 ( .A(n5248), .B(n59929), .Z(n5250) );
  AND U5740 ( .A(n5249), .B(n5250), .Z(n5251) );
  ANDN U5741 ( .B(n59932), .A(n59931), .Z(n5252) );
  NANDN U5742 ( .A(n5251), .B(n59930), .Z(n5253) );
  AND U5743 ( .A(n5252), .B(n5253), .Z(n59935) );
  NOR U5744 ( .A(n50845), .B(n50846), .Z(n5254) );
  NANDN U5745 ( .A(n59966), .B(n59965), .Z(n5255) );
  AND U5746 ( .A(n5254), .B(n5255), .Z(n5256) );
  ANDN U5747 ( .B(n59969), .A(n59968), .Z(n5257) );
  NANDN U5748 ( .A(n5256), .B(n59967), .Z(n5258) );
  AND U5749 ( .A(n5257), .B(n5258), .Z(n5259) );
  ANDN U5750 ( .B(n59972), .A(n59971), .Z(n5260) );
  NANDN U5751 ( .A(n5259), .B(n59970), .Z(n5261) );
  AND U5752 ( .A(n5260), .B(n5261), .Z(n5262) );
  ANDN U5753 ( .B(n59974), .A(n59973), .Z(n5263) );
  NANDN U5754 ( .A(n5262), .B(n50843), .Z(n5264) );
  AND U5755 ( .A(n5263), .B(n5264), .Z(n5265) );
  ANDN U5756 ( .B(n59976), .A(n50842), .Z(n5266) );
  NANDN U5757 ( .A(n5265), .B(n59975), .Z(n5267) );
  AND U5758 ( .A(n5266), .B(n5267), .Z(n5268) );
  OR U5759 ( .A(n5268), .B(n59977), .Z(n5269) );
  ANDN U5760 ( .B(n5269), .A(n59978), .Z(n59980) );
  AND U5761 ( .A(n50828), .B(n50827), .Z(n5270) );
  NANDN U5762 ( .A(n50829), .B(n60002), .Z(n5271) );
  AND U5763 ( .A(n5270), .B(n5271), .Z(n5272) );
  NANDN U5764 ( .A(n5272), .B(n60003), .Z(n5273) );
  AND U5765 ( .A(n60004), .B(n5273), .Z(n5274) );
  AND U5766 ( .A(n60007), .B(n60006), .Z(n5275) );
  NANDN U5767 ( .A(n5274), .B(n60005), .Z(n5276) );
  NAND U5768 ( .A(n5275), .B(n5276), .Z(n5277) );
  NAND U5769 ( .A(n50826), .B(n5277), .Z(n5278) );
  AND U5770 ( .A(n60008), .B(n5278), .Z(n5279) );
  NAND U5771 ( .A(n5279), .B(n60009), .Z(n5280) );
  NAND U5772 ( .A(n60010), .B(n5280), .Z(n5281) );
  AND U5773 ( .A(n60012), .B(n5281), .Z(n5282) );
  NANDN U5774 ( .A(n60011), .B(n5282), .Z(n5283) );
  NAND U5775 ( .A(n60013), .B(n5283), .Z(n5284) );
  AND U5776 ( .A(n60014), .B(n5284), .Z(n5285) );
  NAND U5777 ( .A(n5285), .B(n60015), .Z(n60016) );
  AND U5778 ( .A(n60047), .B(n60048), .Z(n5286) );
  ANDN U5779 ( .B(n50816), .A(n50817), .Z(n5287) );
  NANDN U5780 ( .A(n5286), .B(n60049), .Z(n5288) );
  AND U5781 ( .A(n5287), .B(n5288), .Z(n5289) );
  ANDN U5782 ( .B(n60052), .A(n60051), .Z(n5290) );
  NANDN U5783 ( .A(n5289), .B(n60050), .Z(n5291) );
  AND U5784 ( .A(n5290), .B(n5291), .Z(n5292) );
  ANDN U5785 ( .B(n50815), .A(n50814), .Z(n5293) );
  OR U5786 ( .A(n60053), .B(n5292), .Z(n5294) );
  AND U5787 ( .A(n5293), .B(n5294), .Z(n5295) );
  NANDN U5788 ( .A(n5295), .B(n50813), .Z(n5296) );
  NAND U5789 ( .A(n60054), .B(n5296), .Z(n5297) );
  NAND U5790 ( .A(n60055), .B(n5297), .Z(n5298) );
  AND U5791 ( .A(n60056), .B(n50812), .Z(n5299) );
  NAND U5792 ( .A(n5298), .B(n5299), .Z(n5300) );
  NAND U5793 ( .A(n60057), .B(n5300), .Z(n60058) );
  ANDN U5794 ( .B(n60088), .A(n60087), .Z(n5301) );
  NAND U5795 ( .A(n60086), .B(n50804), .Z(n5302) );
  AND U5796 ( .A(n5301), .B(n5302), .Z(n5303) );
  AND U5797 ( .A(n60091), .B(n60090), .Z(n5304) );
  NANDN U5798 ( .A(n5303), .B(n60089), .Z(n5305) );
  AND U5799 ( .A(n5304), .B(n5305), .Z(n5306) );
  ANDN U5800 ( .B(n50803), .A(n50802), .Z(n5307) );
  OR U5801 ( .A(n60092), .B(n5306), .Z(n5308) );
  AND U5802 ( .A(n5307), .B(n5308), .Z(n5309) );
  AND U5803 ( .A(n60095), .B(n60094), .Z(n5310) );
  NANDN U5804 ( .A(n5309), .B(n60093), .Z(n5311) );
  AND U5805 ( .A(n5310), .B(n5311), .Z(n5312) );
  AND U5806 ( .A(n50800), .B(n50801), .Z(n5313) );
  NANDN U5807 ( .A(n5312), .B(n60096), .Z(n5314) );
  AND U5808 ( .A(n5313), .B(n5314), .Z(n5315) );
  NANDN U5809 ( .A(n5315), .B(n60097), .Z(n5316) );
  AND U5810 ( .A(n60098), .B(n5316), .Z(n60100) );
  NAND U5811 ( .A(n60132), .B(n60131), .Z(n5317) );
  AND U5812 ( .A(n60134), .B(n5317), .Z(n5318) );
  NOR U5813 ( .A(n50794), .B(n5318), .Z(n5319) );
  NAND U5814 ( .A(n50793), .B(n5319), .Z(n5320) );
  NAND U5815 ( .A(n60135), .B(n5320), .Z(n5321) );
  AND U5816 ( .A(n50792), .B(n50791), .Z(n5322) );
  NAND U5817 ( .A(n5321), .B(n5322), .Z(n5323) );
  NAND U5818 ( .A(n60136), .B(n5323), .Z(n5324) );
  ANDN U5819 ( .B(n60138), .A(n60137), .Z(n5325) );
  NAND U5820 ( .A(n5324), .B(n5325), .Z(n5326) );
  NAND U5821 ( .A(n60139), .B(n5326), .Z(n5327) );
  ANDN U5822 ( .B(n50790), .A(n50789), .Z(n5328) );
  NAND U5823 ( .A(n5327), .B(n5328), .Z(n5329) );
  NANDN U5824 ( .A(n60140), .B(n5329), .Z(n5330) );
  ANDN U5825 ( .B(n60142), .A(n60141), .Z(n5331) );
  NAND U5826 ( .A(n5330), .B(n5331), .Z(n5332) );
  NAND U5827 ( .A(n60143), .B(n5332), .Z(n5333) );
  AND U5828 ( .A(n60144), .B(n5333), .Z(n60145) );
  ANDN U5829 ( .B(n60172), .A(n50779), .Z(n5334) );
  NAND U5830 ( .A(n50778), .B(n5334), .Z(n5335) );
  NAND U5831 ( .A(n60173), .B(n5335), .Z(n5336) );
  ANDN U5832 ( .B(n60174), .A(n60175), .Z(n5337) );
  NAND U5833 ( .A(n5336), .B(n5337), .Z(n5338) );
  NAND U5834 ( .A(n60176), .B(n5338), .Z(n5339) );
  ANDN U5835 ( .B(n50777), .A(n50776), .Z(n5340) );
  NAND U5836 ( .A(n5339), .B(n5340), .Z(n5341) );
  NANDN U5837 ( .A(n60177), .B(n5341), .Z(n5342) );
  AND U5838 ( .A(n60179), .B(n60178), .Z(n5343) );
  NAND U5839 ( .A(n5342), .B(n5343), .Z(n5344) );
  NAND U5840 ( .A(n60180), .B(n5344), .Z(n5345) );
  AND U5841 ( .A(n60182), .B(n60181), .Z(n5346) );
  NAND U5842 ( .A(n5345), .B(n5346), .Z(n5347) );
  NAND U5843 ( .A(n60183), .B(n5347), .Z(n5348) );
  AND U5844 ( .A(n60185), .B(n60184), .Z(n5349) );
  NAND U5845 ( .A(n5348), .B(n5349), .Z(n5350) );
  NAND U5846 ( .A(n60186), .B(n5350), .Z(n5351) );
  AND U5847 ( .A(n60187), .B(n5351), .Z(n60189) );
  ANDN U5848 ( .B(n60216), .A(n60215), .Z(n5352) );
  NAND U5849 ( .A(n60217), .B(n5352), .Z(n5353) );
  NANDN U5850 ( .A(n60218), .B(n5353), .Z(n5354) );
  AND U5851 ( .A(n60220), .B(n60219), .Z(n5355) );
  NAND U5852 ( .A(n5354), .B(n5355), .Z(n5356) );
  NAND U5853 ( .A(n60221), .B(n5356), .Z(n5357) );
  AND U5854 ( .A(n60222), .B(n60223), .Z(n5358) );
  NAND U5855 ( .A(n5357), .B(n5358), .Z(n5359) );
  NANDN U5856 ( .A(n60224), .B(n5359), .Z(n5360) );
  ANDN U5857 ( .B(n50764), .A(n50765), .Z(n5361) );
  NAND U5858 ( .A(n5360), .B(n5361), .Z(n5362) );
  NAND U5859 ( .A(n60225), .B(n5362), .Z(n5363) );
  ANDN U5860 ( .B(n60227), .A(n60226), .Z(n5364) );
  NAND U5861 ( .A(n5363), .B(n5364), .Z(n5365) );
  NAND U5862 ( .A(n60228), .B(n5365), .Z(n5366) );
  NANDN U5863 ( .A(n50763), .B(n5366), .Z(n60229) );
  NAND U5864 ( .A(n60256), .B(n60257), .Z(n5367) );
  AND U5865 ( .A(n50756), .B(n50755), .Z(n5368) );
  NANDN U5866 ( .A(n60259), .B(n5367), .Z(n5369) );
  NAND U5867 ( .A(n5368), .B(n5369), .Z(n5370) );
  NAND U5868 ( .A(n60260), .B(n5370), .Z(n5371) );
  AND U5869 ( .A(n50754), .B(n5371), .Z(n5372) );
  NANDN U5870 ( .A(n50753), .B(n5372), .Z(n5373) );
  AND U5871 ( .A(n50752), .B(n50751), .Z(n5374) );
  NANDN U5872 ( .A(n60261), .B(n5373), .Z(n5375) );
  NAND U5873 ( .A(n5374), .B(n5375), .Z(n5376) );
  NAND U5874 ( .A(n60262), .B(n5376), .Z(n5377) );
  AND U5875 ( .A(n60264), .B(n5377), .Z(n5378) );
  NANDN U5876 ( .A(n60263), .B(n5378), .Z(n5379) );
  AND U5877 ( .A(n60266), .B(n60265), .Z(n5380) );
  NANDN U5878 ( .A(n50750), .B(n5379), .Z(n5381) );
  NAND U5879 ( .A(n5380), .B(n5381), .Z(n60267) );
  AND U5880 ( .A(n60292), .B(n60295), .Z(n5382) );
  NAND U5881 ( .A(n60293), .B(n5382), .Z(n5383) );
  NANDN U5882 ( .A(n60296), .B(n5383), .Z(n5384) );
  ANDN U5883 ( .B(n60298), .A(n60297), .Z(n5385) );
  NAND U5884 ( .A(n5384), .B(n5385), .Z(n5386) );
  NAND U5885 ( .A(n60299), .B(n5386), .Z(n5387) );
  AND U5886 ( .A(n50740), .B(n50741), .Z(n5388) );
  NAND U5887 ( .A(n5387), .B(n5388), .Z(n5389) );
  NAND U5888 ( .A(n60300), .B(n5389), .Z(n5390) );
  ANDN U5889 ( .B(n60302), .A(n60301), .Z(n5391) );
  NAND U5890 ( .A(n5390), .B(n5391), .Z(n5392) );
  NAND U5891 ( .A(n60303), .B(n5392), .Z(n5393) );
  ANDN U5892 ( .B(n60304), .A(n60305), .Z(n5394) );
  NAND U5893 ( .A(n5393), .B(n5394), .Z(n5395) );
  NANDN U5894 ( .A(n60306), .B(n5395), .Z(n5396) );
  ANDN U5895 ( .B(n5396), .A(n60307), .Z(n5397) );
  NAND U5896 ( .A(n60308), .B(n5397), .Z(n60309) );
  NAND U5897 ( .A(n60338), .B(n60339), .Z(n5398) );
  AND U5898 ( .A(n60340), .B(n5398), .Z(n5399) );
  NANDN U5899 ( .A(n60341), .B(n5399), .Z(n5400) );
  NAND U5900 ( .A(n60342), .B(n5400), .Z(n5401) );
  AND U5901 ( .A(n50728), .B(n5401), .Z(n5402) );
  NANDN U5902 ( .A(n50729), .B(n5402), .Z(n5403) );
  NAND U5903 ( .A(n60343), .B(n5403), .Z(n5404) );
  AND U5904 ( .A(n60344), .B(n5404), .Z(n5405) );
  NANDN U5905 ( .A(n60345), .B(n5405), .Z(n5406) );
  ANDN U5906 ( .B(n50727), .A(n50726), .Z(n5407) );
  NANDN U5907 ( .A(n60346), .B(n5406), .Z(n5408) );
  NAND U5908 ( .A(n5407), .B(n5408), .Z(n5409) );
  NAND U5909 ( .A(n50725), .B(n5409), .Z(n5410) );
  AND U5910 ( .A(n60348), .B(n5410), .Z(n5411) );
  NAND U5911 ( .A(n5411), .B(n60347), .Z(n5412) );
  AND U5912 ( .A(n60349), .B(n5412), .Z(n60351) );
  ANDN U5913 ( .B(n50719), .A(n50718), .Z(n5413) );
  OR U5914 ( .A(n60384), .B(n60383), .Z(n5414) );
  NAND U5915 ( .A(n5413), .B(n5414), .Z(n5415) );
  NAND U5916 ( .A(n50717), .B(n5415), .Z(n5416) );
  NAND U5917 ( .A(n60385), .B(n5416), .Z(n5417) );
  ANDN U5918 ( .B(n5417), .A(n60386), .Z(n5418) );
  ANDN U5919 ( .B(n50716), .A(n5418), .Z(n5419) );
  NAND U5920 ( .A(n50715), .B(n5419), .Z(n5420) );
  ANDN U5921 ( .B(n5420), .A(n50714), .Z(n5421) );
  NOR U5922 ( .A(n50712), .B(n5421), .Z(n5422) );
  NAND U5923 ( .A(n50713), .B(n5422), .Z(n5423) );
  AND U5924 ( .A(n60387), .B(n5423), .Z(n5424) );
  NANDN U5925 ( .A(n5424), .B(n60388), .Z(n5425) );
  NANDN U5926 ( .A(n60389), .B(n5425), .Z(n5426) );
  NAND U5927 ( .A(n60390), .B(n5426), .Z(n60391) );
  NAND U5928 ( .A(n60420), .B(n50704), .Z(n5427) );
  AND U5929 ( .A(n60422), .B(n5427), .Z(n5428) );
  NANDN U5930 ( .A(n60421), .B(n5428), .Z(n5429) );
  ANDN U5931 ( .B(n60424), .A(n60425), .Z(n5430) );
  NANDN U5932 ( .A(n60423), .B(n5429), .Z(n5431) );
  NAND U5933 ( .A(n5430), .B(n5431), .Z(n5432) );
  NAND U5934 ( .A(n60426), .B(n5432), .Z(n5433) );
  AND U5935 ( .A(n50703), .B(n5433), .Z(n5434) );
  NANDN U5936 ( .A(n50702), .B(n5434), .Z(n5435) );
  NAND U5937 ( .A(n60427), .B(n5435), .Z(n5436) );
  AND U5938 ( .A(n60429), .B(n5436), .Z(n5437) );
  NANDN U5939 ( .A(n60428), .B(n5437), .Z(n5438) );
  NAND U5940 ( .A(n60430), .B(n5438), .Z(n5439) );
  AND U5941 ( .A(n60432), .B(n5439), .Z(n5440) );
  NANDN U5942 ( .A(n60431), .B(n5440), .Z(n5441) );
  AND U5943 ( .A(n60435), .B(n60434), .Z(n5442) );
  NANDN U5944 ( .A(n60433), .B(n5441), .Z(n5443) );
  NAND U5945 ( .A(n5442), .B(n5443), .Z(n60436) );
  NAND U5946 ( .A(n60463), .B(n60462), .Z(n5444) );
  ANDN U5947 ( .B(n5444), .A(n60464), .Z(n5445) );
  ANDN U5948 ( .B(n60466), .A(n5445), .Z(n5446) );
  NAND U5949 ( .A(n60465), .B(n5446), .Z(n5447) );
  NAND U5950 ( .A(n60467), .B(n5447), .Z(n5448) );
  ANDN U5951 ( .B(n60469), .A(n60468), .Z(n5449) );
  NAND U5952 ( .A(n5448), .B(n5449), .Z(n5450) );
  NAND U5953 ( .A(n50692), .B(n5450), .Z(n5451) );
  AND U5954 ( .A(n60471), .B(n60470), .Z(n5452) );
  NAND U5955 ( .A(n5451), .B(n5452), .Z(n5453) );
  NAND U5956 ( .A(n60472), .B(n5453), .Z(n5454) );
  ANDN U5957 ( .B(n60474), .A(n60473), .Z(n5455) );
  NAND U5958 ( .A(n5454), .B(n5455), .Z(n5456) );
  NANDN U5959 ( .A(n60475), .B(n5456), .Z(n5457) );
  ANDN U5960 ( .B(n50691), .A(n50690), .Z(n5458) );
  NAND U5961 ( .A(n5457), .B(n5458), .Z(n5459) );
  NAND U5962 ( .A(n60476), .B(n5459), .Z(n5460) );
  ANDN U5963 ( .B(n5460), .A(n60477), .Z(n60479) );
  AND U5964 ( .A(n60509), .B(n60510), .Z(n5461) );
  NAND U5965 ( .A(n60511), .B(n5461), .Z(n5462) );
  NANDN U5966 ( .A(n60512), .B(n5462), .Z(n5463) );
  ANDN U5967 ( .B(n50684), .A(n50683), .Z(n5464) );
  NAND U5968 ( .A(n5463), .B(n5464), .Z(n5465) );
  NAND U5969 ( .A(n60513), .B(n5465), .Z(n5466) );
  ANDN U5970 ( .B(n50681), .A(n50682), .Z(n5467) );
  NAND U5971 ( .A(n5466), .B(n5467), .Z(n5468) );
  NAND U5972 ( .A(n60514), .B(n5468), .Z(n5469) );
  ANDN U5973 ( .B(n60515), .A(n60516), .Z(n5470) );
  NAND U5974 ( .A(n5469), .B(n5470), .Z(n5471) );
  NAND U5975 ( .A(n60517), .B(n5471), .Z(n5472) );
  ANDN U5976 ( .B(n50680), .A(n50679), .Z(n5473) );
  NAND U5977 ( .A(n5472), .B(n5473), .Z(n5474) );
  NAND U5978 ( .A(n50678), .B(n5474), .Z(n5475) );
  AND U5979 ( .A(n60518), .B(n5475), .Z(n60520) );
  ANDN U5980 ( .B(n50675), .A(n50674), .Z(n60536) );
  AND U5981 ( .A(n60562), .B(n60563), .Z(n5476) );
  NANDN U5982 ( .A(n60561), .B(n60560), .Z(n5477) );
  AND U5983 ( .A(n5476), .B(n5477), .Z(n5478) );
  ANDN U5984 ( .B(n60565), .A(n50659), .Z(n5479) );
  NANDN U5985 ( .A(n5478), .B(n60564), .Z(n5480) );
  AND U5986 ( .A(n5479), .B(n5480), .Z(n5481) );
  NOR U5987 ( .A(n60566), .B(n50657), .Z(n5482) );
  NANDN U5988 ( .A(n5481), .B(n50658), .Z(n5483) );
  AND U5989 ( .A(n5482), .B(n5483), .Z(n5484) );
  AND U5990 ( .A(n60569), .B(n60568), .Z(n5485) );
  NANDN U5991 ( .A(n5484), .B(n60567), .Z(n5486) );
  AND U5992 ( .A(n5485), .B(n5486), .Z(n5487) );
  ANDN U5993 ( .B(n50656), .A(n50655), .Z(n5488) );
  OR U5994 ( .A(n60570), .B(n5487), .Z(n5489) );
  AND U5995 ( .A(n5488), .B(n5489), .Z(n5490) );
  OR U5996 ( .A(n60571), .B(n5490), .Z(n5491) );
  AND U5997 ( .A(n60572), .B(n5491), .Z(n60574) );
  NANDN U5998 ( .A(n60605), .B(n60604), .Z(n5492) );
  ANDN U5999 ( .B(n5492), .A(n60606), .Z(n5493) );
  ANDN U6000 ( .B(n60608), .A(n5493), .Z(n5494) );
  NAND U6001 ( .A(n60607), .B(n5494), .Z(n5495) );
  NAND U6002 ( .A(n60609), .B(n5495), .Z(n5496) );
  ANDN U6003 ( .B(n50647), .A(n50648), .Z(n5497) );
  NAND U6004 ( .A(n5496), .B(n5497), .Z(n5498) );
  NANDN U6005 ( .A(n50646), .B(n5498), .Z(n5499) );
  ANDN U6006 ( .B(n50645), .A(n50644), .Z(n5500) );
  NAND U6007 ( .A(n5499), .B(n5500), .Z(n5501) );
  NAND U6008 ( .A(n60610), .B(n5501), .Z(n5502) );
  NAND U6009 ( .A(n60611), .B(n5502), .Z(n5503) );
  NANDN U6010 ( .A(n60612), .B(n5503), .Z(n5504) );
  AND U6011 ( .A(n60613), .B(n5504), .Z(n5505) );
  NANDN U6012 ( .A(n5505), .B(n60614), .Z(n5506) );
  NAND U6013 ( .A(n60615), .B(n5506), .Z(n5507) );
  NAND U6014 ( .A(n60616), .B(n5507), .Z(n5508) );
  AND U6015 ( .A(n60617), .B(n5508), .Z(n60619) );
  AND U6016 ( .A(n60641), .B(n60640), .Z(n5509) );
  NAND U6017 ( .A(n60643), .B(n5509), .Z(n5510) );
  NANDN U6018 ( .A(n60644), .B(n5510), .Z(n5511) );
  ANDN U6019 ( .B(n50629), .A(n50628), .Z(n5512) );
  NAND U6020 ( .A(n5511), .B(n5512), .Z(n5513) );
  NAND U6021 ( .A(n50627), .B(n5513), .Z(n5514) );
  AND U6022 ( .A(n60646), .B(n60645), .Z(n5515) );
  NAND U6023 ( .A(n5514), .B(n5515), .Z(n5516) );
  NAND U6024 ( .A(n60647), .B(n5516), .Z(n5517) );
  ANDN U6025 ( .B(n60649), .A(n60648), .Z(n5518) );
  NAND U6026 ( .A(n5517), .B(n5518), .Z(n5519) );
  NAND U6027 ( .A(n60650), .B(n5519), .Z(n5520) );
  AND U6028 ( .A(n60652), .B(n60651), .Z(n5521) );
  NAND U6029 ( .A(n5520), .B(n5521), .Z(n5522) );
  NAND U6030 ( .A(n60653), .B(n5522), .Z(n5523) );
  ANDN U6031 ( .B(n60655), .A(n60654), .Z(n5524) );
  NAND U6032 ( .A(n5523), .B(n5524), .Z(n5525) );
  NAND U6033 ( .A(n60656), .B(n5525), .Z(n60657) );
  AND U6034 ( .A(n60733), .B(n60734), .Z(n5526) );
  NAND U6035 ( .A(n60732), .B(n5526), .Z(n5527) );
  AND U6036 ( .A(n60735), .B(n5527), .Z(n5528) );
  NOR U6037 ( .A(n60736), .B(n5528), .Z(n5529) );
  NAND U6038 ( .A(n60737), .B(n5529), .Z(n5530) );
  ANDN U6039 ( .B(n5530), .A(n60738), .Z(n5531) );
  ANDN U6040 ( .B(n60740), .A(n5531), .Z(n5532) );
  NAND U6041 ( .A(n60739), .B(n5532), .Z(n5533) );
  AND U6042 ( .A(n60741), .B(n5533), .Z(n5534) );
  NANDN U6043 ( .A(n5534), .B(n60742), .Z(n5535) );
  AND U6044 ( .A(n60743), .B(n5535), .Z(n5536) );
  ANDN U6045 ( .B(n50605), .A(n5536), .Z(n5537) );
  NAND U6046 ( .A(n50604), .B(n5537), .Z(n5538) );
  AND U6047 ( .A(n60744), .B(n5538), .Z(n5539) );
  NANDN U6048 ( .A(n5539), .B(n60745), .Z(n5540) );
  NAND U6049 ( .A(n60746), .B(n5540), .Z(n5541) );
  NANDN U6050 ( .A(n50603), .B(n5541), .Z(n60747) );
  NAND U6051 ( .A(n60771), .B(n60770), .Z(n5542) );
  NAND U6052 ( .A(n60772), .B(n5542), .Z(n5543) );
  AND U6053 ( .A(n60773), .B(n5543), .Z(n5544) );
  NAND U6054 ( .A(n5544), .B(n60774), .Z(n5545) );
  NAND U6055 ( .A(n50591), .B(n5545), .Z(n5546) );
  ANDN U6056 ( .B(n5546), .A(n60775), .Z(n5547) );
  NAND U6057 ( .A(n60776), .B(n5547), .Z(n5548) );
  NAND U6058 ( .A(n60777), .B(n5548), .Z(n5549) );
  AND U6059 ( .A(n50590), .B(n5549), .Z(n5550) );
  NANDN U6060 ( .A(n50589), .B(n5550), .Z(n5551) );
  ANDN U6061 ( .B(n50586), .A(n50587), .Z(n5552) );
  NANDN U6062 ( .A(n50588), .B(n5551), .Z(n5553) );
  NAND U6063 ( .A(n5552), .B(n5553), .Z(n5554) );
  NAND U6064 ( .A(n60778), .B(n5554), .Z(n5555) );
  AND U6065 ( .A(n60779), .B(n5555), .Z(n5556) );
  NAND U6066 ( .A(n5556), .B(n60780), .Z(n60783) );
  AND U6067 ( .A(n50572), .B(n50573), .Z(n5557) );
  OR U6068 ( .A(n60853), .B(n60854), .Z(n5558) );
  AND U6069 ( .A(n5557), .B(n5558), .Z(n5559) );
  ANDN U6070 ( .B(n60857), .A(n60856), .Z(n5560) );
  NANDN U6071 ( .A(n5559), .B(n60855), .Z(n5561) );
  AND U6072 ( .A(n5560), .B(n5561), .Z(n5562) );
  ANDN U6073 ( .B(n60859), .A(n50571), .Z(n5563) );
  NANDN U6074 ( .A(n5562), .B(n60858), .Z(n5564) );
  AND U6075 ( .A(n5563), .B(n5564), .Z(n5565) );
  ANDN U6076 ( .B(n60862), .A(n60861), .Z(n5566) );
  NANDN U6077 ( .A(n5565), .B(n60860), .Z(n5567) );
  AND U6078 ( .A(n5566), .B(n5567), .Z(n5568) );
  ANDN U6079 ( .B(n60864), .A(n60865), .Z(n5569) );
  NANDN U6080 ( .A(n5568), .B(n60863), .Z(n5570) );
  AND U6081 ( .A(n5569), .B(n5570), .Z(n5571) );
  ANDN U6082 ( .B(n50570), .A(n50569), .Z(n5572) );
  OR U6083 ( .A(n60866), .B(n5571), .Z(n5573) );
  AND U6084 ( .A(n5572), .B(n5573), .Z(n60869) );
  NAND U6085 ( .A(n60898), .B(n60897), .Z(n5574) );
  NAND U6086 ( .A(n50561), .B(n5574), .Z(n5575) );
  NAND U6087 ( .A(n60899), .B(n5575), .Z(n5576) );
  NAND U6088 ( .A(n60900), .B(n5576), .Z(n5577) );
  AND U6089 ( .A(n60901), .B(n5577), .Z(n5578) );
  NANDN U6090 ( .A(n60902), .B(n5578), .Z(n5579) );
  NAND U6091 ( .A(n60903), .B(n5579), .Z(n5580) );
  AND U6092 ( .A(n50559), .B(n5580), .Z(n5581) );
  NANDN U6093 ( .A(n50560), .B(n5581), .Z(n5582) );
  NAND U6094 ( .A(n60904), .B(n5582), .Z(n5583) );
  AND U6095 ( .A(n60905), .B(n5583), .Z(n5584) );
  NANDN U6096 ( .A(n60906), .B(n5584), .Z(n5585) );
  NAND U6097 ( .A(n60907), .B(n5585), .Z(n5586) );
  AND U6098 ( .A(n50558), .B(n5586), .Z(n5587) );
  NANDN U6099 ( .A(n50557), .B(n5587), .Z(n5588) );
  NANDN U6100 ( .A(n60908), .B(n5588), .Z(n60909) );
  NAND U6101 ( .A(n60939), .B(n60938), .Z(n5589) );
  AND U6102 ( .A(n60940), .B(n5589), .Z(n5590) );
  NOR U6103 ( .A(n60942), .B(n5590), .Z(n5591) );
  NAND U6104 ( .A(n60941), .B(n5591), .Z(n5592) );
  NAND U6105 ( .A(n60943), .B(n5592), .Z(n5593) );
  ANDN U6106 ( .B(n50547), .A(n50546), .Z(n5594) );
  NAND U6107 ( .A(n5593), .B(n5594), .Z(n5595) );
  NANDN U6108 ( .A(n60944), .B(n5595), .Z(n5596) );
  AND U6109 ( .A(n60946), .B(n60945), .Z(n5597) );
  NAND U6110 ( .A(n5596), .B(n5597), .Z(n5598) );
  NAND U6111 ( .A(n60947), .B(n5598), .Z(n5599) );
  ANDN U6112 ( .B(n60949), .A(n60948), .Z(n5600) );
  NAND U6113 ( .A(n5599), .B(n5600), .Z(n5601) );
  NAND U6114 ( .A(n50545), .B(n5601), .Z(n5602) );
  AND U6115 ( .A(n60951), .B(n60950), .Z(n5603) );
  NAND U6116 ( .A(n5602), .B(n5603), .Z(n5604) );
  NAND U6117 ( .A(n60952), .B(n5604), .Z(n60954) );
  AND U6118 ( .A(n60978), .B(n60977), .Z(n5605) );
  NAND U6119 ( .A(n60979), .B(n5605), .Z(n5606) );
  AND U6120 ( .A(n60980), .B(n5606), .Z(n5607) );
  NOR U6121 ( .A(n60981), .B(n50533), .Z(n5608) );
  NANDN U6122 ( .A(n5607), .B(n5608), .Z(n5609) );
  AND U6123 ( .A(n50532), .B(n5609), .Z(n5610) );
  ANDN U6124 ( .B(n60983), .A(n5610), .Z(n5611) );
  NAND U6125 ( .A(n60982), .B(n5611), .Z(n5612) );
  AND U6126 ( .A(n60984), .B(n5612), .Z(n5613) );
  NOR U6127 ( .A(n60985), .B(n5613), .Z(n5614) );
  NAND U6128 ( .A(n60986), .B(n5614), .Z(n5615) );
  AND U6129 ( .A(n60987), .B(n5615), .Z(n5616) );
  NOR U6130 ( .A(n50531), .B(n5616), .Z(n5617) );
  NAND U6131 ( .A(n50530), .B(n5617), .Z(n5618) );
  AND U6132 ( .A(n60988), .B(n5618), .Z(n5619) );
  NANDN U6133 ( .A(n5619), .B(n60989), .Z(n5620) );
  AND U6134 ( .A(n60990), .B(n5620), .Z(n60994) );
  ANDN U6135 ( .B(n61025), .A(n61024), .Z(n5621) );
  NANDN U6136 ( .A(n61023), .B(n61022), .Z(n5622) );
  AND U6137 ( .A(n5621), .B(n5622), .Z(n5623) );
  ANDN U6138 ( .B(n61027), .A(n50520), .Z(n5624) );
  NANDN U6139 ( .A(n5623), .B(n61026), .Z(n5625) );
  AND U6140 ( .A(n5624), .B(n5625), .Z(n5626) );
  ANDN U6141 ( .B(n61030), .A(n61029), .Z(n5627) );
  OR U6142 ( .A(n5626), .B(n61028), .Z(n5628) );
  NAND U6143 ( .A(n5627), .B(n5628), .Z(n5629) );
  NAND U6144 ( .A(n61031), .B(n5629), .Z(n5630) );
  AND U6145 ( .A(n61032), .B(n5630), .Z(n5631) );
  NAND U6146 ( .A(n5631), .B(n61033), .Z(n5632) );
  AND U6147 ( .A(n50519), .B(n50518), .Z(n5633) );
  NANDN U6148 ( .A(n61034), .B(n5632), .Z(n5634) );
  NAND U6149 ( .A(n5633), .B(n5634), .Z(n5635) );
  NAND U6150 ( .A(n61035), .B(n5635), .Z(n61036) );
  NAND U6151 ( .A(n61068), .B(n61069), .Z(n5636) );
  AND U6152 ( .A(n61070), .B(n5636), .Z(n5637) );
  NAND U6153 ( .A(n5637), .B(n61071), .Z(n5638) );
  ANDN U6154 ( .B(n50510), .A(n50509), .Z(n5639) );
  NANDN U6155 ( .A(n61072), .B(n5638), .Z(n5640) );
  NAND U6156 ( .A(n5639), .B(n5640), .Z(n5641) );
  NAND U6157 ( .A(n61073), .B(n5641), .Z(n5642) );
  AND U6158 ( .A(n61074), .B(n5642), .Z(n5643) );
  NANDN U6159 ( .A(n61075), .B(n5643), .Z(n5644) );
  NAND U6160 ( .A(n61076), .B(n5644), .Z(n5645) );
  AND U6161 ( .A(n50508), .B(n5645), .Z(n5646) );
  NANDN U6162 ( .A(n50507), .B(n5646), .Z(n5647) );
  AND U6163 ( .A(n61078), .B(n61079), .Z(n5648) );
  NANDN U6164 ( .A(n61077), .B(n5647), .Z(n5649) );
  NAND U6165 ( .A(n5648), .B(n5649), .Z(n5650) );
  NAND U6166 ( .A(n61080), .B(n5650), .Z(n5651) );
  AND U6167 ( .A(n61082), .B(n5651), .Z(n5652) );
  NANDN U6168 ( .A(n61081), .B(n5652), .Z(n61083) );
  OR U6169 ( .A(n61110), .B(n61111), .Z(n5653) );
  ANDN U6170 ( .B(n5653), .A(n50497), .Z(n5654) );
  AND U6171 ( .A(n61113), .B(n61112), .Z(n5655) );
  NANDN U6172 ( .A(n5654), .B(n50496), .Z(n5656) );
  AND U6173 ( .A(n5655), .B(n5656), .Z(n5657) );
  AND U6174 ( .A(n61116), .B(n61115), .Z(n5658) );
  NANDN U6175 ( .A(n5657), .B(n61114), .Z(n5659) );
  AND U6176 ( .A(n5658), .B(n5659), .Z(n5660) );
  OR U6177 ( .A(n50495), .B(n5660), .Z(n5661) );
  NAND U6178 ( .A(n50494), .B(n5661), .Z(n5662) );
  NAND U6179 ( .A(n61117), .B(n5662), .Z(n5663) );
  AND U6180 ( .A(n61119), .B(n61118), .Z(n5664) );
  NAND U6181 ( .A(n5663), .B(n5664), .Z(n5665) );
  NAND U6182 ( .A(n61120), .B(n5665), .Z(n61121) );
  NAND U6183 ( .A(n61142), .B(n61141), .Z(n5666) );
  AND U6184 ( .A(n61143), .B(n5666), .Z(n5667) );
  ANDN U6185 ( .B(n61144), .A(n5667), .Z(n5668) );
  NAND U6186 ( .A(n61145), .B(n5668), .Z(n5669) );
  NANDN U6187 ( .A(n61146), .B(n5669), .Z(n5670) );
  ANDN U6188 ( .B(n50479), .A(n50478), .Z(n5671) );
  NAND U6189 ( .A(n5670), .B(n5671), .Z(n5672) );
  NAND U6190 ( .A(n61147), .B(n5672), .Z(n5673) );
  ANDN U6191 ( .B(n61148), .A(n61149), .Z(n5674) );
  NAND U6192 ( .A(n5673), .B(n5674), .Z(n5675) );
  NANDN U6193 ( .A(n61150), .B(n5675), .Z(n5676) );
  ANDN U6194 ( .B(n50477), .A(n50476), .Z(n5677) );
  NAND U6195 ( .A(n5676), .B(n5677), .Z(n5678) );
  NANDN U6196 ( .A(n61151), .B(n5678), .Z(n5679) );
  AND U6197 ( .A(n61153), .B(n61152), .Z(n5680) );
  NAND U6198 ( .A(n5679), .B(n5680), .Z(n5681) );
  NAND U6199 ( .A(n61154), .B(n5681), .Z(n5682) );
  ANDN U6200 ( .B(n5682), .A(n61155), .Z(n61157) );
  ANDN U6201 ( .B(n61188), .A(n61187), .Z(n5683) );
  OR U6202 ( .A(n61185), .B(n61186), .Z(n5684) );
  NAND U6203 ( .A(n5683), .B(n5684), .Z(n5685) );
  NAND U6204 ( .A(n61189), .B(n5685), .Z(n5686) );
  AND U6205 ( .A(n50468), .B(n5686), .Z(n5687) );
  NANDN U6206 ( .A(n50467), .B(n5687), .Z(n5688) );
  AND U6207 ( .A(n61191), .B(n61192), .Z(n5689) );
  NANDN U6208 ( .A(n61190), .B(n5688), .Z(n5690) );
  NAND U6209 ( .A(n5689), .B(n5690), .Z(n5691) );
  AND U6210 ( .A(n61194), .B(n61195), .Z(n5692) );
  NANDN U6211 ( .A(n61193), .B(n5691), .Z(n5693) );
  NAND U6212 ( .A(n5692), .B(n5693), .Z(n5694) );
  NAND U6213 ( .A(n61196), .B(n5694), .Z(n5695) );
  AND U6214 ( .A(n61198), .B(n5695), .Z(n5696) );
  NAND U6215 ( .A(n5696), .B(n61197), .Z(n5697) );
  NAND U6216 ( .A(n61199), .B(n5697), .Z(n61200) );
  AND U6217 ( .A(n61283), .B(e), .Z(n5698) );
  ANDN U6218 ( .B(n61274), .A(n50444), .Z(n5699) );
  NAND U6219 ( .A(n50445), .B(n5699), .Z(n5700) );
  AND U6220 ( .A(n61275), .B(n5700), .Z(n5701) );
  NANDN U6221 ( .A(n5701), .B(n61276), .Z(n5702) );
  NAND U6222 ( .A(n61277), .B(n5702), .Z(n5703) );
  NAND U6223 ( .A(n61278), .B(n5703), .Z(n5704) );
  NAND U6224 ( .A(n61279), .B(n5704), .Z(n5705) );
  NANDN U6225 ( .A(n61280), .B(n61281), .Z(n5706) );
  NAND U6226 ( .A(n5705), .B(n5706), .Z(n5707) );
  NANDN U6227 ( .A(n5707), .B(n61282), .Z(n5708) );
  AND U6228 ( .A(n50443), .B(n5708), .Z(n5709) );
  XOR U6229 ( .A(n5709), .B(y[8191]), .Z(n5710) );
  NANDN U6230 ( .A(x[8191]), .B(n5710), .Z(n5711) );
  NAND U6231 ( .A(n5709), .B(y[8191]), .Z(n5712) );
  AND U6232 ( .A(n5711), .B(n5712), .Z(n5713) );
  NAND U6233 ( .A(n5713), .B(n5698), .Z(n5714) );
  NANDN U6234 ( .A(n5698), .B(g), .Z(n5715) );
  NAND U6235 ( .A(n5714), .B(n5715), .Z(n4) );
  ANDN U6236 ( .B(n34411), .A(n34410), .Z(n5716) );
  AND U6237 ( .A(n34414), .B(n34413), .Z(n5717) );
  NANDN U6238 ( .A(n34412), .B(n5716), .Z(n5718) );
  NAND U6239 ( .A(n5717), .B(n5718), .Z(n5719) );
  NAND U6240 ( .A(n27407), .B(n27408), .Z(n5720) );
  NOR U6241 ( .A(n34416), .B(n34415), .Z(n5721) );
  NAND U6242 ( .A(n5719), .B(n5721), .Z(n5722) );
  NANDN U6243 ( .A(n5720), .B(n5722), .Z(n5723) );
  ANDN U6244 ( .B(n5723), .A(n34417), .Z(n5724) );
  XNOR U6245 ( .A(y[1966]), .B(x[1966]), .Z(n5725) );
  AND U6246 ( .A(n5724), .B(n5725), .Z(n5726) );
  NOR U6247 ( .A(n5726), .B(n34418), .Z(n5727) );
  NANDN U6248 ( .A(x[1966]), .B(y[1966]), .Z(n5728) );
  AND U6249 ( .A(n5727), .B(n5728), .Z(n5729) );
  NANDN U6250 ( .A(n5729), .B(n52170), .Z(n5730) );
  ANDN U6251 ( .B(n5730), .A(n52169), .Z(n5731) );
  ANDN U6252 ( .B(n34420), .A(n52171), .Z(n5732) );
  NANDN U6253 ( .A(n34419), .B(n5731), .Z(n5733) );
  NAND U6254 ( .A(n5732), .B(n5733), .Z(n34421) );
  NANDN U6255 ( .A(n52443), .B(n52442), .Z(n5734) );
  NAND U6256 ( .A(n52444), .B(n5734), .Z(n5735) );
  NAND U6257 ( .A(n52445), .B(n5735), .Z(n5736) );
  NANDN U6258 ( .A(n52446), .B(n5736), .Z(n5737) );
  NAND U6259 ( .A(n52447), .B(n5737), .Z(n5738) );
  ANDN U6260 ( .B(n5738), .A(n52448), .Z(n5739) );
  NANDN U6261 ( .A(n5739), .B(n52449), .Z(n5740) );
  NANDN U6262 ( .A(n52450), .B(n5740), .Z(n5741) );
  NAND U6263 ( .A(n52451), .B(n5741), .Z(n5742) );
  NAND U6264 ( .A(n52452), .B(n5742), .Z(n5743) );
  NAND U6265 ( .A(n52453), .B(n5743), .Z(n5744) );
  ANDN U6266 ( .B(n5744), .A(n52454), .Z(n5745) );
  NANDN U6267 ( .A(n5745), .B(n52455), .Z(n5746) );
  NANDN U6268 ( .A(n52437), .B(n5746), .Z(n5747) );
  NAND U6269 ( .A(n52456), .B(n5747), .Z(n5748) );
  NANDN U6270 ( .A(n52457), .B(n5748), .Z(n5749) );
  NAND U6271 ( .A(n52458), .B(n5749), .Z(n5750) );
  AND U6272 ( .A(n52459), .B(n5750), .Z(n52461) );
  NAND U6273 ( .A(n52491), .B(n52492), .Z(n5751) );
  NANDN U6274 ( .A(n52493), .B(n5751), .Z(n5752) );
  AND U6275 ( .A(n52494), .B(n5752), .Z(n5753) );
  NANDN U6276 ( .A(n5753), .B(n52495), .Z(n5754) );
  NAND U6277 ( .A(n52496), .B(n5754), .Z(n5755) );
  NANDN U6278 ( .A(n52497), .B(n5755), .Z(n5756) );
  NAND U6279 ( .A(n52498), .B(n5756), .Z(n5757) );
  NANDN U6280 ( .A(n52499), .B(n5757), .Z(n5758) );
  AND U6281 ( .A(n52500), .B(n5758), .Z(n5759) );
  OR U6282 ( .A(n52501), .B(n5759), .Z(n5760) );
  NAND U6283 ( .A(n52502), .B(n5760), .Z(n5761) );
  NAND U6284 ( .A(n52503), .B(n5761), .Z(n5762) );
  NAND U6285 ( .A(n52504), .B(n5762), .Z(n5763) );
  NANDN U6286 ( .A(n52505), .B(n5763), .Z(n5764) );
  AND U6287 ( .A(n52506), .B(n5764), .Z(n5765) );
  OR U6288 ( .A(n52430), .B(n5765), .Z(n5766) );
  NAND U6289 ( .A(n52507), .B(n5766), .Z(n5767) );
  NANDN U6290 ( .A(n52508), .B(n5767), .Z(n52509) );
  OR U6291 ( .A(n52568), .B(n52567), .Z(n5768) );
  NAND U6292 ( .A(n52569), .B(n5768), .Z(n5769) );
  NANDN U6293 ( .A(n52570), .B(n5769), .Z(n5770) );
  NANDN U6294 ( .A(n52571), .B(n5770), .Z(n5771) );
  NAND U6295 ( .A(n52572), .B(n5771), .Z(n5772) );
  ANDN U6296 ( .B(n5772), .A(n52428), .Z(n5773) );
  NANDN U6297 ( .A(n5773), .B(n52427), .Z(n5774) );
  NANDN U6298 ( .A(n52573), .B(n5774), .Z(n5775) );
  NANDN U6299 ( .A(n52574), .B(n5775), .Z(n5776) );
  NAND U6300 ( .A(n52575), .B(n5776), .Z(n5777) );
  NANDN U6301 ( .A(n52576), .B(n5777), .Z(n5778) );
  AND U6302 ( .A(n52577), .B(n5778), .Z(n5779) );
  OR U6303 ( .A(n52578), .B(n5779), .Z(n5780) );
  AND U6304 ( .A(n52579), .B(n5780), .Z(n5781) );
  OR U6305 ( .A(n52580), .B(n5781), .Z(n5782) );
  NAND U6306 ( .A(n52581), .B(n5782), .Z(n5783) );
  NANDN U6307 ( .A(n52582), .B(n5783), .Z(n52583) );
  NAND U6308 ( .A(n52415), .B(n52599), .Z(n5784) );
  NANDN U6309 ( .A(n52414), .B(n5784), .Z(n5785) );
  AND U6310 ( .A(n52413), .B(n5785), .Z(n5786) );
  OR U6311 ( .A(n52600), .B(n5786), .Z(n5787) );
  NAND U6312 ( .A(n52601), .B(n5787), .Z(n5788) );
  NANDN U6313 ( .A(n52412), .B(n5788), .Z(n5789) );
  NAND U6314 ( .A(n52602), .B(n5789), .Z(n5790) );
  NAND U6315 ( .A(n52603), .B(n5790), .Z(n5791) );
  AND U6316 ( .A(n52604), .B(n5791), .Z(n5792) );
  NANDN U6317 ( .A(n5792), .B(n52605), .Z(n5793) );
  AND U6318 ( .A(n52606), .B(n5793), .Z(n5794) );
  NANDN U6319 ( .A(n5794), .B(n52607), .Z(n5795) );
  NANDN U6320 ( .A(n52608), .B(n5795), .Z(n5796) );
  NAND U6321 ( .A(n52609), .B(n5796), .Z(n52610) );
  NANDN U6322 ( .A(n52411), .B(n52670), .Z(n5797) );
  NAND U6323 ( .A(n52410), .B(n5797), .Z(n5798) );
  AND U6324 ( .A(n52671), .B(n5798), .Z(n5799) );
  OR U6325 ( .A(n52672), .B(n5799), .Z(n5800) );
  NAND U6326 ( .A(n52673), .B(n5800), .Z(n5801) );
  NANDN U6327 ( .A(n52674), .B(n5801), .Z(n5802) );
  NAND U6328 ( .A(n52675), .B(n5802), .Z(n5803) );
  NANDN U6329 ( .A(n52676), .B(n5803), .Z(n5804) );
  AND U6330 ( .A(n52677), .B(n5804), .Z(n5805) );
  OR U6331 ( .A(n52678), .B(n5805), .Z(n5806) );
  NAND U6332 ( .A(n52679), .B(n5806), .Z(n5807) );
  NANDN U6333 ( .A(n52680), .B(n5807), .Z(n5808) );
  NAND U6334 ( .A(n52681), .B(n5808), .Z(n5809) );
  NAND U6335 ( .A(n52682), .B(n5809), .Z(n5810) );
  AND U6336 ( .A(n52683), .B(n5810), .Z(n5811) );
  OR U6337 ( .A(n52684), .B(n5811), .Z(n5812) );
  NAND U6338 ( .A(n52685), .B(n5812), .Z(n5813) );
  NANDN U6339 ( .A(n52686), .B(n5813), .Z(n52687) );
  NAND U6340 ( .A(n52751), .B(n52752), .Z(n5814) );
  NANDN U6341 ( .A(n52753), .B(n5814), .Z(n5815) );
  NAND U6342 ( .A(n52754), .B(n5815), .Z(n5816) );
  NAND U6343 ( .A(n52400), .B(n5816), .Z(n5817) );
  NAND U6344 ( .A(n52755), .B(n5817), .Z(n5818) );
  ANDN U6345 ( .B(n5818), .A(n52756), .Z(n5819) );
  NANDN U6346 ( .A(n5819), .B(n52757), .Z(n5820) );
  NANDN U6347 ( .A(n52758), .B(n5820), .Z(n5821) );
  NAND U6348 ( .A(n52759), .B(n5821), .Z(n5822) );
  NANDN U6349 ( .A(n52760), .B(n5822), .Z(n5823) );
  NAND U6350 ( .A(n52761), .B(n5823), .Z(n5824) );
  ANDN U6351 ( .B(n5824), .A(n52762), .Z(n5825) );
  OR U6352 ( .A(n52763), .B(n5825), .Z(n5826) );
  NAND U6353 ( .A(n52764), .B(n5826), .Z(n5827) );
  NANDN U6354 ( .A(n52399), .B(n5827), .Z(n5828) );
  NAND U6355 ( .A(n52398), .B(n5828), .Z(n52765) );
  NANDN U6356 ( .A(n52847), .B(n52846), .Z(n5829) );
  NAND U6357 ( .A(n52848), .B(n5829), .Z(n5830) );
  NANDN U6358 ( .A(n52397), .B(n5830), .Z(n5831) );
  NAND U6359 ( .A(n52849), .B(n5831), .Z(n5832) );
  NANDN U6360 ( .A(n52850), .B(n5832), .Z(n5833) );
  ANDN U6361 ( .B(n5833), .A(n52851), .Z(n5834) );
  OR U6362 ( .A(n52852), .B(n5834), .Z(n5835) );
  NANDN U6363 ( .A(n52853), .B(n5835), .Z(n5836) );
  NAND U6364 ( .A(n52854), .B(n5836), .Z(n5837) );
  NANDN U6365 ( .A(n52855), .B(n5837), .Z(n5838) );
  NAND U6366 ( .A(n52856), .B(n5838), .Z(n5839) );
  ANDN U6367 ( .B(n5839), .A(n52857), .Z(n5840) );
  OR U6368 ( .A(n52858), .B(n5840), .Z(n5841) );
  AND U6369 ( .A(n52859), .B(n5841), .Z(n5842) );
  OR U6370 ( .A(n52860), .B(n5842), .Z(n5843) );
  NANDN U6371 ( .A(n52861), .B(n5843), .Z(n5844) );
  NANDN U6372 ( .A(n52396), .B(n5844), .Z(n52862) );
  NANDN U6373 ( .A(n52875), .B(n52874), .Z(n5845) );
  NANDN U6374 ( .A(n52381), .B(n5845), .Z(n5846) );
  AND U6375 ( .A(n52876), .B(n5846), .Z(n5847) );
  OR U6376 ( .A(n52877), .B(n5847), .Z(n5848) );
  NAND U6377 ( .A(n52878), .B(n5848), .Z(n5849) );
  NANDN U6378 ( .A(n52380), .B(n5849), .Z(n5850) );
  NAND U6379 ( .A(n52879), .B(n5850), .Z(n5851) );
  NAND U6380 ( .A(n52880), .B(n5851), .Z(n5852) );
  AND U6381 ( .A(n52881), .B(n5852), .Z(n5853) );
  NANDN U6382 ( .A(n5853), .B(n52882), .Z(n5854) );
  AND U6383 ( .A(n52883), .B(n5854), .Z(n5855) );
  OR U6384 ( .A(n52884), .B(n5855), .Z(n5856) );
  NAND U6385 ( .A(n52379), .B(n5856), .Z(n5857) );
  NANDN U6386 ( .A(n52378), .B(n5857), .Z(n52885) );
  NAND U6387 ( .A(n52902), .B(n52903), .Z(n5858) );
  NAND U6388 ( .A(n52904), .B(n5858), .Z(n5859) );
  NANDN U6389 ( .A(n52365), .B(n5859), .Z(n5860) );
  NAND U6390 ( .A(n52905), .B(n5860), .Z(n5861) );
  NANDN U6391 ( .A(n52364), .B(n5861), .Z(n5862) );
  AND U6392 ( .A(n52906), .B(n5862), .Z(n5863) );
  OR U6393 ( .A(n52907), .B(n5863), .Z(n5864) );
  NAND U6394 ( .A(n52908), .B(n5864), .Z(n5865) );
  NANDN U6395 ( .A(n52363), .B(n5865), .Z(n5866) );
  NAND U6396 ( .A(n52909), .B(n5866), .Z(n5867) );
  NANDN U6397 ( .A(n52910), .B(n5867), .Z(n5868) );
  AND U6398 ( .A(n52911), .B(n5868), .Z(n5869) );
  NANDN U6399 ( .A(n5869), .B(n52912), .Z(n5870) );
  NANDN U6400 ( .A(n52913), .B(n5870), .Z(n5871) );
  NAND U6401 ( .A(n52914), .B(n5871), .Z(n52915) );
  NANDN U6402 ( .A(n52943), .B(n52944), .Z(n5872) );
  NANDN U6403 ( .A(n52946), .B(n5872), .Z(n5873) );
  ANDN U6404 ( .B(n5873), .A(n52357), .Z(n5874) );
  NANDN U6405 ( .A(n5874), .B(n52356), .Z(n5875) );
  NANDN U6406 ( .A(n52947), .B(n5875), .Z(n5876) );
  NANDN U6407 ( .A(n52948), .B(n5876), .Z(n5877) );
  NAND U6408 ( .A(n52949), .B(n5877), .Z(n5878) );
  NANDN U6409 ( .A(n52950), .B(n5878), .Z(n5879) );
  AND U6410 ( .A(n52951), .B(n5879), .Z(n5880) );
  OR U6411 ( .A(n52952), .B(n5880), .Z(n5881) );
  NAND U6412 ( .A(n52953), .B(n5881), .Z(n5882) );
  NANDN U6413 ( .A(n52954), .B(n5882), .Z(n5883) );
  NAND U6414 ( .A(n52955), .B(n5883), .Z(n5884) );
  NANDN U6415 ( .A(n52956), .B(n5884), .Z(n5885) );
  AND U6416 ( .A(n52957), .B(n5885), .Z(n5886) );
  OR U6417 ( .A(n52958), .B(n5886), .Z(n5887) );
  NAND U6418 ( .A(n52959), .B(n5887), .Z(n5888) );
  NANDN U6419 ( .A(n52960), .B(n5888), .Z(n52961) );
  NANDN U6420 ( .A(n53000), .B(n52999), .Z(n5889) );
  NAND U6421 ( .A(n53001), .B(n5889), .Z(n5890) );
  NANDN U6422 ( .A(n53002), .B(n5890), .Z(n5891) );
  NANDN U6423 ( .A(n53003), .B(n5891), .Z(n5892) );
  NAND U6424 ( .A(n53004), .B(n5892), .Z(n5893) );
  ANDN U6425 ( .B(n5893), .A(n52354), .Z(n5894) );
  NANDN U6426 ( .A(n5894), .B(n52353), .Z(n5895) );
  NAND U6427 ( .A(n53005), .B(n5895), .Z(n5896) );
  NANDN U6428 ( .A(n53006), .B(n5896), .Z(n5897) );
  NAND U6429 ( .A(n53007), .B(n5897), .Z(n5898) );
  NANDN U6430 ( .A(n53008), .B(n5898), .Z(n5899) );
  AND U6431 ( .A(n53009), .B(n5899), .Z(n5900) );
  OR U6432 ( .A(n53010), .B(n5900), .Z(n5901) );
  AND U6433 ( .A(n53011), .B(n5901), .Z(n5902) );
  OR U6434 ( .A(n53012), .B(n5902), .Z(n5903) );
  NAND U6435 ( .A(n53013), .B(n5903), .Z(n5904) );
  NANDN U6436 ( .A(n53014), .B(n5904), .Z(n53015) );
  NAND U6437 ( .A(n53054), .B(n53055), .Z(n5905) );
  NANDN U6438 ( .A(n53056), .B(n5905), .Z(n5906) );
  NAND U6439 ( .A(n53057), .B(n5906), .Z(n5907) );
  NANDN U6440 ( .A(n53058), .B(n5907), .Z(n5908) );
  NAND U6441 ( .A(n53059), .B(n5908), .Z(n5909) );
  ANDN U6442 ( .B(n5909), .A(n53060), .Z(n5910) );
  NANDN U6443 ( .A(n5910), .B(n53061), .Z(n5911) );
  NANDN U6444 ( .A(n53062), .B(n5911), .Z(n5912) );
  NAND U6445 ( .A(n53063), .B(n5912), .Z(n5913) );
  NAND U6446 ( .A(n53064), .B(n5913), .Z(n5914) );
  NAND U6447 ( .A(n53065), .B(n5914), .Z(n5915) );
  AND U6448 ( .A(n52351), .B(n5915), .Z(n5916) );
  OR U6449 ( .A(n53066), .B(n5916), .Z(n5917) );
  ANDN U6450 ( .B(n5917), .A(n53067), .Z(n5918) );
  NANDN U6451 ( .A(n5918), .B(n53068), .Z(n5919) );
  NAND U6452 ( .A(n53069), .B(n5919), .Z(n5920) );
  NANDN U6453 ( .A(n52350), .B(n5920), .Z(n53070) );
  NAND U6454 ( .A(n53103), .B(n53104), .Z(n5921) );
  NANDN U6455 ( .A(n53105), .B(n5921), .Z(n5922) );
  AND U6456 ( .A(n53106), .B(n5922), .Z(n5923) );
  OR U6457 ( .A(n53107), .B(n5923), .Z(n5924) );
  NAND U6458 ( .A(n53108), .B(n5924), .Z(n5925) );
  NANDN U6459 ( .A(n53109), .B(n5925), .Z(n5926) );
  NAND U6460 ( .A(n53110), .B(n5926), .Z(n5927) );
  NANDN U6461 ( .A(n53111), .B(n5927), .Z(n5928) );
  AND U6462 ( .A(n53112), .B(n5928), .Z(n5929) );
  NANDN U6463 ( .A(n5929), .B(n53113), .Z(n5930) );
  NANDN U6464 ( .A(n53114), .B(n5930), .Z(n5931) );
  NAND U6465 ( .A(n53115), .B(n5931), .Z(n5932) );
  NAND U6466 ( .A(n53116), .B(n5932), .Z(n5933) );
  NANDN U6467 ( .A(n53117), .B(n5933), .Z(n5934) );
  AND U6468 ( .A(n52346), .B(n5934), .Z(n5935) );
  OR U6469 ( .A(n53118), .B(n5935), .Z(n5936) );
  NAND U6470 ( .A(n53119), .B(n5936), .Z(n5937) );
  NAND U6471 ( .A(n53120), .B(n5937), .Z(n53121) );
  NAND U6472 ( .A(n53171), .B(n53170), .Z(n5938) );
  NANDN U6473 ( .A(n53173), .B(n5938), .Z(n5939) );
  ANDN U6474 ( .B(n5939), .A(n52339), .Z(n5940) );
  NANDN U6475 ( .A(n5940), .B(n52338), .Z(n5941) );
  NANDN U6476 ( .A(n52337), .B(n5941), .Z(n5942) );
  NAND U6477 ( .A(n52336), .B(n5942), .Z(n5943) );
  NANDN U6478 ( .A(n53174), .B(n5943), .Z(n5944) );
  NAND U6479 ( .A(n53175), .B(n5944), .Z(n5945) );
  ANDN U6480 ( .B(n5945), .A(n52335), .Z(n5946) );
  NANDN U6481 ( .A(n5946), .B(n53176), .Z(n5947) );
  NANDN U6482 ( .A(n52334), .B(n5947), .Z(n5948) );
  NAND U6483 ( .A(n53177), .B(n5948), .Z(n53180) );
  NAND U6484 ( .A(n53209), .B(n53208), .Z(n5949) );
  NAND U6485 ( .A(n53210), .B(n5949), .Z(n5950) );
  ANDN U6486 ( .B(n5950), .A(n52327), .Z(n5951) );
  NANDN U6487 ( .A(n5951), .B(n53211), .Z(n5952) );
  NAND U6488 ( .A(n53212), .B(n5952), .Z(n5953) );
  NANDN U6489 ( .A(n53213), .B(n5953), .Z(n5954) );
  NANDN U6490 ( .A(n53214), .B(n5954), .Z(n5955) );
  NAND U6491 ( .A(n53215), .B(n5955), .Z(n5956) );
  ANDN U6492 ( .B(n5956), .A(n53216), .Z(n5957) );
  NANDN U6493 ( .A(n5957), .B(n53217), .Z(n5958) );
  NANDN U6494 ( .A(n53218), .B(n5958), .Z(n5959) );
  NANDN U6495 ( .A(n53219), .B(n5959), .Z(n5960) );
  NAND U6496 ( .A(n53220), .B(n5960), .Z(n5961) );
  NANDN U6497 ( .A(n53221), .B(n5961), .Z(n5962) );
  AND U6498 ( .A(n53222), .B(n5962), .Z(n5963) );
  OR U6499 ( .A(n53223), .B(n5963), .Z(n5964) );
  NAND U6500 ( .A(n53224), .B(n5964), .Z(n5965) );
  NANDN U6501 ( .A(n53225), .B(n5965), .Z(n53226) );
  NAND U6502 ( .A(n53253), .B(n53252), .Z(n5966) );
  NAND U6503 ( .A(n53254), .B(n5966), .Z(n5967) );
  ANDN U6504 ( .B(n5967), .A(n52318), .Z(n5968) );
  NANDN U6505 ( .A(n5968), .B(n53255), .Z(n5969) );
  NANDN U6506 ( .A(n53256), .B(n5969), .Z(n5970) );
  NANDN U6507 ( .A(n53257), .B(n5970), .Z(n5971) );
  NAND U6508 ( .A(n53258), .B(n5971), .Z(n5972) );
  NANDN U6509 ( .A(n53259), .B(n5972), .Z(n5973) );
  AND U6510 ( .A(n53260), .B(n5973), .Z(n5974) );
  OR U6511 ( .A(n53261), .B(n5974), .Z(n5975) );
  NAND U6512 ( .A(n53262), .B(n5975), .Z(n5976) );
  NANDN U6513 ( .A(n53263), .B(n5976), .Z(n5977) );
  NAND U6514 ( .A(n53264), .B(n5977), .Z(n5978) );
  NANDN U6515 ( .A(n53265), .B(n5978), .Z(n5979) );
  AND U6516 ( .A(n53266), .B(n5979), .Z(n5980) );
  OR U6517 ( .A(n53267), .B(n5980), .Z(n5981) );
  NAND U6518 ( .A(n53268), .B(n5981), .Z(n5982) );
  NANDN U6519 ( .A(n53269), .B(n5982), .Z(n53271) );
  OR U6520 ( .A(n53302), .B(n53301), .Z(n5983) );
  NANDN U6521 ( .A(n52313), .B(n5983), .Z(n5984) );
  NAND U6522 ( .A(n53303), .B(n5984), .Z(n5985) );
  NANDN U6523 ( .A(n52312), .B(n5985), .Z(n5986) );
  NAND U6524 ( .A(n53304), .B(n5986), .Z(n5987) );
  ANDN U6525 ( .B(n5987), .A(n53305), .Z(n5988) );
  NANDN U6526 ( .A(n5988), .B(n53306), .Z(n5989) );
  NANDN U6527 ( .A(n53307), .B(n5989), .Z(n5990) );
  NAND U6528 ( .A(n53308), .B(n5990), .Z(n5991) );
  NANDN U6529 ( .A(n53309), .B(n5991), .Z(n5992) );
  NAND U6530 ( .A(n53310), .B(n5992), .Z(n5993) );
  ANDN U6531 ( .B(n5993), .A(n53311), .Z(n5994) );
  NANDN U6532 ( .A(n5994), .B(n53312), .Z(n5995) );
  NAND U6533 ( .A(n53313), .B(n5995), .Z(n5996) );
  NANDN U6534 ( .A(n53314), .B(n5996), .Z(n5997) );
  NAND U6535 ( .A(n53315), .B(n5997), .Z(n5998) );
  NANDN U6536 ( .A(n53316), .B(n5998), .Z(n5999) );
  AND U6537 ( .A(n53317), .B(n5999), .Z(n53319) );
  NANDN U6538 ( .A(n53350), .B(n53349), .Z(n6000) );
  NAND U6539 ( .A(n52307), .B(n6000), .Z(n6001) );
  NANDN U6540 ( .A(n53351), .B(n6001), .Z(n6002) );
  NAND U6541 ( .A(n53352), .B(n6002), .Z(n6003) );
  NANDN U6542 ( .A(n52306), .B(n6003), .Z(n6004) );
  ANDN U6543 ( .B(n6004), .A(n53353), .Z(n6005) );
  NANDN U6544 ( .A(n6005), .B(n53354), .Z(n6006) );
  AND U6545 ( .A(n53355), .B(n6006), .Z(n6007) );
  NANDN U6546 ( .A(n6007), .B(n53356), .Z(n6008) );
  NAND U6547 ( .A(n53357), .B(n6008), .Z(n6009) );
  NAND U6548 ( .A(n53358), .B(n6009), .Z(n6010) );
  NAND U6549 ( .A(n53359), .B(n6010), .Z(n6011) );
  AND U6550 ( .A(n52304), .B(n6011), .Z(n6012) );
  NAND U6551 ( .A(n6012), .B(n52305), .Z(n6013) );
  AND U6552 ( .A(n53361), .B(n53360), .Z(n6014) );
  NAND U6553 ( .A(n6013), .B(n6014), .Z(n6015) );
  NANDN U6554 ( .A(n53362), .B(n6015), .Z(n53363) );
  NAND U6555 ( .A(n53418), .B(n53419), .Z(n6016) );
  ANDN U6556 ( .B(n6016), .A(n53420), .Z(n6017) );
  NANDN U6557 ( .A(n6017), .B(n53421), .Z(n6018) );
  NANDN U6558 ( .A(n53422), .B(n6018), .Z(n6019) );
  NANDN U6559 ( .A(n53423), .B(n6019), .Z(n6020) );
  AND U6560 ( .A(n52301), .B(n52300), .Z(n6021) );
  NANDN U6561 ( .A(n6020), .B(n53424), .Z(n6022) );
  AND U6562 ( .A(n6021), .B(n6022), .Z(n6023) );
  NOR U6563 ( .A(n53425), .B(n6023), .Z(n6024) );
  NAND U6564 ( .A(n53426), .B(n6024), .Z(n6025) );
  ANDN U6565 ( .B(n6025), .A(n53427), .Z(n6026) );
  NANDN U6566 ( .A(n6026), .B(n53428), .Z(n6027) );
  ANDN U6567 ( .B(n6027), .A(n52299), .Z(n6028) );
  NANDN U6568 ( .A(n6028), .B(n53429), .Z(n6029) );
  NANDN U6569 ( .A(n52298), .B(n6029), .Z(n6030) );
  NAND U6570 ( .A(n52297), .B(n6030), .Z(n53432) );
  ANDN U6571 ( .B(n27880), .A(n27879), .Z(n53455) );
  NAND U6572 ( .A(n53482), .B(n53481), .Z(n6031) );
  NANDN U6573 ( .A(n53484), .B(n6031), .Z(n6032) );
  ANDN U6574 ( .B(n6032), .A(n52281), .Z(n6033) );
  OR U6575 ( .A(n6033), .B(n53485), .Z(n6034) );
  NAND U6576 ( .A(n53486), .B(n6034), .Z(n6035) );
  ANDN U6577 ( .B(n6035), .A(n53487), .Z(n6036) );
  NANDN U6578 ( .A(n6036), .B(n53488), .Z(n6037) );
  NANDN U6579 ( .A(n53489), .B(n6037), .Z(n6038) );
  NANDN U6580 ( .A(n53490), .B(n6038), .Z(n6039) );
  NAND U6581 ( .A(n53491), .B(n6039), .Z(n6040) );
  NANDN U6582 ( .A(n53492), .B(n6040), .Z(n6041) );
  AND U6583 ( .A(n53493), .B(n6041), .Z(n6042) );
  OR U6584 ( .A(n52280), .B(n6042), .Z(n6043) );
  NAND U6585 ( .A(n53494), .B(n6043), .Z(n6044) );
  NAND U6586 ( .A(n53495), .B(n6044), .Z(n53496) );
  NANDN U6587 ( .A(n52272), .B(n53521), .Z(n6045) );
  NAND U6588 ( .A(n53522), .B(n6045), .Z(n6046) );
  ANDN U6589 ( .B(n6046), .A(n53523), .Z(n6047) );
  NANDN U6590 ( .A(n6047), .B(n53524), .Z(n6048) );
  NANDN U6591 ( .A(n52271), .B(n6048), .Z(n6049) );
  NAND U6592 ( .A(n52270), .B(n6049), .Z(n6050) );
  NANDN U6593 ( .A(n52269), .B(n6050), .Z(n6051) );
  NAND U6594 ( .A(n53525), .B(n6051), .Z(n6052) );
  ANDN U6595 ( .B(n6052), .A(n53526), .Z(n6053) );
  NANDN U6596 ( .A(n6053), .B(n53527), .Z(n6054) );
  NANDN U6597 ( .A(n52268), .B(n6054), .Z(n6055) );
  NAND U6598 ( .A(n53528), .B(n6055), .Z(n53530) );
  OR U6599 ( .A(n53561), .B(n53562), .Z(n6056) );
  NAND U6600 ( .A(n53563), .B(n6056), .Z(n6057) );
  ANDN U6601 ( .B(n6057), .A(n53564), .Z(n6058) );
  NANDN U6602 ( .A(n6058), .B(n53565), .Z(n6059) );
  NANDN U6603 ( .A(n52263), .B(n6059), .Z(n6060) );
  NANDN U6604 ( .A(n53566), .B(n6060), .Z(n6061) );
  NANDN U6605 ( .A(n52262), .B(n6061), .Z(n6062) );
  NAND U6606 ( .A(n53567), .B(n6062), .Z(n6063) );
  AND U6607 ( .A(n53568), .B(n6063), .Z(n6064) );
  NANDN U6608 ( .A(n6064), .B(n53569), .Z(n6065) );
  NAND U6609 ( .A(n53570), .B(n6065), .Z(n6066) );
  NAND U6610 ( .A(n53571), .B(n6066), .Z(n6067) );
  NANDN U6611 ( .A(n53572), .B(n6067), .Z(n6068) );
  NAND U6612 ( .A(n53573), .B(n6068), .Z(n6069) );
  ANDN U6613 ( .B(n6069), .A(n53574), .Z(n6070) );
  NANDN U6614 ( .A(n6070), .B(n53575), .Z(n6071) );
  NANDN U6615 ( .A(n53576), .B(n6071), .Z(n6072) );
  NAND U6616 ( .A(n53577), .B(n6072), .Z(n53578) );
  NAND U6617 ( .A(n53606), .B(n53607), .Z(n6073) );
  NANDN U6618 ( .A(n53608), .B(n6073), .Z(n6074) );
  ANDN U6619 ( .B(n6074), .A(n53609), .Z(n6075) );
  NANDN U6620 ( .A(n6075), .B(n53610), .Z(n6076) );
  NANDN U6621 ( .A(n53611), .B(n6076), .Z(n6077) );
  NAND U6622 ( .A(n53612), .B(n6077), .Z(n6078) );
  NANDN U6623 ( .A(n53613), .B(n6078), .Z(n6079) );
  NAND U6624 ( .A(n53614), .B(n6079), .Z(n6080) );
  ANDN U6625 ( .B(n6080), .A(n53615), .Z(n6081) );
  NANDN U6626 ( .A(n6081), .B(n53616), .Z(n6082) );
  NANDN U6627 ( .A(n53617), .B(n6082), .Z(n6083) );
  NANDN U6628 ( .A(n52256), .B(n6083), .Z(n6084) );
  NAND U6629 ( .A(n53618), .B(n6084), .Z(n6085) );
  NANDN U6630 ( .A(n52255), .B(n6085), .Z(n6086) );
  ANDN U6631 ( .B(n6086), .A(n53619), .Z(n6087) );
  ANDN U6632 ( .B(n53620), .A(n6087), .Z(n6088) );
  NANDN U6633 ( .A(n53622), .B(n53621), .Z(n6089) );
  NAND U6634 ( .A(n6088), .B(n6089), .Z(n53623) );
  OR U6635 ( .A(n53675), .B(n53674), .Z(n6090) );
  NAND U6636 ( .A(n53676), .B(n6090), .Z(n6091) );
  ANDN U6637 ( .B(n6091), .A(n53677), .Z(n6092) );
  NANDN U6638 ( .A(n6092), .B(n53678), .Z(n6093) );
  NAND U6639 ( .A(n53679), .B(n6093), .Z(n6094) );
  NAND U6640 ( .A(n53680), .B(n6094), .Z(n6095) );
  AND U6641 ( .A(n6095), .B(n53681), .Z(n6096) );
  OR U6642 ( .A(n53682), .B(n53683), .Z(n6097) );
  AND U6643 ( .A(n6096), .B(n6097), .Z(n6098) );
  OR U6644 ( .A(n53684), .B(n6098), .Z(n6099) );
  ANDN U6645 ( .B(n6099), .A(n52249), .Z(n6100) );
  NANDN U6646 ( .A(n6100), .B(n53685), .Z(n6101) );
  NAND U6647 ( .A(n53686), .B(n6101), .Z(n6102) );
  NAND U6648 ( .A(n52248), .B(n6102), .Z(n6103) );
  ANDN U6649 ( .B(n53687), .A(n52247), .Z(n6104) );
  NAND U6650 ( .A(n6103), .B(n6104), .Z(n6105) );
  NAND U6651 ( .A(n53688), .B(n6105), .Z(n53689) );
  ANDN U6652 ( .B(n27699), .A(n27698), .Z(n53711) );
  NAND U6653 ( .A(n53744), .B(n53743), .Z(n6106) );
  NAND U6654 ( .A(n53745), .B(n6106), .Z(n6107) );
  NAND U6655 ( .A(n53746), .B(n6107), .Z(n6108) );
  NAND U6656 ( .A(n52242), .B(n6108), .Z(n6109) );
  NAND U6657 ( .A(n53747), .B(n6109), .Z(n6110) );
  AND U6658 ( .A(n52241), .B(n6110), .Z(n6111) );
  OR U6659 ( .A(n53748), .B(n6111), .Z(n6112) );
  NAND U6660 ( .A(n53749), .B(n6112), .Z(n6113) );
  NANDN U6661 ( .A(n52240), .B(n6113), .Z(n6114) );
  NAND U6662 ( .A(n52239), .B(n6114), .Z(n6115) );
  NANDN U6663 ( .A(n52238), .B(n6115), .Z(n6116) );
  ANDN U6664 ( .B(n6116), .A(n53750), .Z(n53751) );
  ANDN U6665 ( .B(n27648), .A(n27647), .Z(n53799) );
  NAND U6666 ( .A(n53824), .B(n53823), .Z(n6117) );
  NAND U6667 ( .A(n52230), .B(n6117), .Z(n6118) );
  ANDN U6668 ( .B(n6118), .A(n52229), .Z(n6119) );
  NANDN U6669 ( .A(n6119), .B(n52228), .Z(n6120) );
  NANDN U6670 ( .A(n53825), .B(n6120), .Z(n6121) );
  NAND U6671 ( .A(n53826), .B(n6121), .Z(n6122) );
  NANDN U6672 ( .A(n52227), .B(n6122), .Z(n6123) );
  NAND U6673 ( .A(n52226), .B(n6123), .Z(n6124) );
  ANDN U6674 ( .B(n6124), .A(n52225), .Z(n6125) );
  NANDN U6675 ( .A(n6125), .B(n53827), .Z(n6126) );
  ANDN U6676 ( .B(n6126), .A(n53828), .Z(n53831) );
  NAND U6677 ( .A(n53858), .B(n53859), .Z(n6127) );
  NANDN U6678 ( .A(n53860), .B(n6127), .Z(n6128) );
  AND U6679 ( .A(n53861), .B(n6128), .Z(n6129) );
  OR U6680 ( .A(n53862), .B(n6129), .Z(n6130) );
  NAND U6681 ( .A(n53863), .B(n6130), .Z(n6131) );
  NANDN U6682 ( .A(n52219), .B(n6131), .Z(n6132) );
  NAND U6683 ( .A(n52218), .B(n6132), .Z(n6133) );
  NANDN U6684 ( .A(n52217), .B(n6133), .Z(n6134) );
  AND U6685 ( .A(n52216), .B(n6134), .Z(n6135) );
  OR U6686 ( .A(n53864), .B(n6135), .Z(n6136) );
  NAND U6687 ( .A(n53865), .B(n6136), .Z(n6137) );
  NANDN U6688 ( .A(n52215), .B(n6137), .Z(n53866) );
  NAND U6689 ( .A(n53897), .B(n53896), .Z(n6138) );
  NANDN U6690 ( .A(n53898), .B(n6138), .Z(n6139) );
  AND U6691 ( .A(n53899), .B(n6139), .Z(n6140) );
  NANDN U6692 ( .A(n6140), .B(n53900), .Z(n6141) );
  NAND U6693 ( .A(n53901), .B(n6141), .Z(n6142) );
  NAND U6694 ( .A(n53902), .B(n6142), .Z(n6143) );
  NANDN U6695 ( .A(n53903), .B(n6143), .Z(n6144) );
  NANDN U6696 ( .A(n53904), .B(n6144), .Z(n6145) );
  ANDN U6697 ( .B(n6145), .A(n53905), .Z(n6146) );
  NANDN U6698 ( .A(n6146), .B(n53906), .Z(n6147) );
  NANDN U6699 ( .A(n53907), .B(n6147), .Z(n6148) );
  NAND U6700 ( .A(n53908), .B(n6148), .Z(n6149) );
  NANDN U6701 ( .A(n53909), .B(n6149), .Z(n6150) );
  NAND U6702 ( .A(n53910), .B(n6150), .Z(n6151) );
  ANDN U6703 ( .B(n6151), .A(n53911), .Z(n6152) );
  NANDN U6704 ( .A(n6152), .B(n52208), .Z(n6153) );
  ANDN U6705 ( .B(n6153), .A(n53912), .Z(n53915) );
  NANDN U6706 ( .A(n53944), .B(n53943), .Z(n6154) );
  NAND U6707 ( .A(n53945), .B(n6154), .Z(n6155) );
  NANDN U6708 ( .A(n53946), .B(n6155), .Z(n6156) );
  NANDN U6709 ( .A(n52202), .B(n6156), .Z(n6157) );
  NAND U6710 ( .A(n52201), .B(n6157), .Z(n6158) );
  ANDN U6711 ( .B(n6158), .A(n52200), .Z(n6159) );
  NANDN U6712 ( .A(n6159), .B(n53947), .Z(n6160) );
  NAND U6713 ( .A(n53948), .B(n6160), .Z(n6161) );
  NANDN U6714 ( .A(n53949), .B(n6161), .Z(n6162) );
  NAND U6715 ( .A(n53950), .B(n6162), .Z(n6163) );
  NANDN U6716 ( .A(n53951), .B(n6163), .Z(n6164) );
  AND U6717 ( .A(n53952), .B(n6164), .Z(n6165) );
  NANDN U6718 ( .A(n6165), .B(n52199), .Z(n6166) );
  NAND U6719 ( .A(n53953), .B(n6166), .Z(n6167) );
  NANDN U6720 ( .A(n53954), .B(n6167), .Z(n6168) );
  NAND U6721 ( .A(n53955), .B(n6168), .Z(n53956) );
  OR U6722 ( .A(n53993), .B(n53994), .Z(n6169) );
  NAND U6723 ( .A(n53995), .B(n6169), .Z(n6170) );
  NANDN U6724 ( .A(n53996), .B(n6170), .Z(n6171) );
  NANDN U6725 ( .A(n52197), .B(n6171), .Z(n6172) );
  NANDN U6726 ( .A(n53997), .B(n6172), .Z(n6173) );
  AND U6727 ( .A(n53998), .B(n6173), .Z(n6174) );
  OR U6728 ( .A(n53999), .B(n6174), .Z(n6175) );
  NAND U6729 ( .A(n54000), .B(n6175), .Z(n6176) );
  NANDN U6730 ( .A(n54001), .B(n6176), .Z(n6177) );
  NAND U6731 ( .A(n54002), .B(n6177), .Z(n6178) );
  NAND U6732 ( .A(n52196), .B(n6178), .Z(n6179) );
  ANDN U6733 ( .B(n6179), .A(n54003), .Z(n6180) );
  NANDN U6734 ( .A(n6180), .B(n54004), .Z(n6181) );
  NAND U6735 ( .A(n54005), .B(n6181), .Z(n6182) );
  NANDN U6736 ( .A(n54006), .B(n6182), .Z(n6183) );
  NAND U6737 ( .A(n54007), .B(n6183), .Z(n54008) );
  NAND U6738 ( .A(n52189), .B(n54036), .Z(n6184) );
  NANDN U6739 ( .A(n52188), .B(n6184), .Z(n6185) );
  NAND U6740 ( .A(n52187), .B(n6185), .Z(n6186) );
  NANDN U6741 ( .A(n54037), .B(n6186), .Z(n6187) );
  NAND U6742 ( .A(n54038), .B(n6187), .Z(n6188) );
  ANDN U6743 ( .B(n6188), .A(n54039), .Z(n6189) );
  NANDN U6744 ( .A(n6189), .B(n54040), .Z(n6190) );
  ANDN U6745 ( .B(n6190), .A(n52186), .Z(n6191) );
  NANDN U6746 ( .A(n6191), .B(n54041), .Z(n6192) );
  NAND U6747 ( .A(n54042), .B(n6192), .Z(n6193) );
  NAND U6748 ( .A(n52185), .B(n6193), .Z(n54044) );
  NANDN U6749 ( .A(n54074), .B(n54073), .Z(n6194) );
  NANDN U6750 ( .A(n54075), .B(n6194), .Z(n6195) );
  AND U6751 ( .A(n54076), .B(n6195), .Z(n6196) );
  OR U6752 ( .A(n52179), .B(n6196), .Z(n6197) );
  NAND U6753 ( .A(n52178), .B(n6197), .Z(n6198) );
  NANDN U6754 ( .A(n54077), .B(n6198), .Z(n6199) );
  NAND U6755 ( .A(n54078), .B(n6199), .Z(n6200) );
  NANDN U6756 ( .A(n54079), .B(n6200), .Z(n6201) );
  AND U6757 ( .A(n54080), .B(n6201), .Z(n6202) );
  OR U6758 ( .A(n6202), .B(n54081), .Z(n6203) );
  NAND U6759 ( .A(n52177), .B(n6203), .Z(n6204) );
  NANDN U6760 ( .A(n54082), .B(n6204), .Z(n6205) );
  NAND U6761 ( .A(n54083), .B(n6205), .Z(n54084) );
  XNOR U6762 ( .A(y[1975]), .B(x[1975]), .Z(n6206) );
  NAND U6763 ( .A(n54104), .B(n6206), .Z(n6207) );
  NAND U6764 ( .A(n54105), .B(n6207), .Z(n6208) );
  NAND U6765 ( .A(n54106), .B(n6208), .Z(n6209) );
  NAND U6766 ( .A(n54107), .B(n6209), .Z(n6210) );
  AND U6767 ( .A(n54108), .B(n6210), .Z(n6211) );
  OR U6768 ( .A(n54109), .B(n6211), .Z(n6212) );
  NAND U6769 ( .A(n52164), .B(n6212), .Z(n6213) );
  NANDN U6770 ( .A(n54110), .B(n6213), .Z(n6214) );
  NAND U6771 ( .A(n54111), .B(n6214), .Z(n6215) );
  NANDN U6772 ( .A(n52163), .B(n6215), .Z(n6216) );
  ANDN U6773 ( .B(n6216), .A(n54112), .Z(n6217) );
  NANDN U6774 ( .A(n6217), .B(n52162), .Z(n6218) );
  ANDN U6775 ( .B(n6218), .A(n54113), .Z(n54116) );
  OR U6776 ( .A(n54144), .B(n54145), .Z(n6219) );
  NANDN U6777 ( .A(n54146), .B(n6219), .Z(n6220) );
  AND U6778 ( .A(n54147), .B(n6220), .Z(n6221) );
  OR U6779 ( .A(n52155), .B(n6221), .Z(n6222) );
  NANDN U6780 ( .A(n54148), .B(n6222), .Z(n6223) );
  NAND U6781 ( .A(n54149), .B(n6223), .Z(n6224) );
  NANDN U6782 ( .A(n54150), .B(n6224), .Z(n6225) );
  NAND U6783 ( .A(n54151), .B(n6225), .Z(n6226) );
  ANDN U6784 ( .B(n6226), .A(n54152), .Z(n6227) );
  NANDN U6785 ( .A(n6227), .B(n54153), .Z(n6228) );
  NANDN U6786 ( .A(n54154), .B(n6228), .Z(n6229) );
  NAND U6787 ( .A(n54155), .B(n6229), .Z(n6230) );
  NANDN U6788 ( .A(n54156), .B(n6230), .Z(n6231) );
  NAND U6789 ( .A(n54157), .B(n6231), .Z(n6232) );
  ANDN U6790 ( .B(n6232), .A(n54158), .Z(n6233) );
  NANDN U6791 ( .A(n6233), .B(n54159), .Z(n6234) );
  NANDN U6792 ( .A(n54160), .B(n6234), .Z(n6235) );
  NAND U6793 ( .A(n54161), .B(n6235), .Z(n54162) );
  OR U6794 ( .A(n54197), .B(n54198), .Z(n6236) );
  NANDN U6795 ( .A(n54199), .B(n6236), .Z(n6237) );
  AND U6796 ( .A(n54200), .B(n6237), .Z(n6238) );
  OR U6797 ( .A(n6238), .B(n54201), .Z(n6239) );
  NAND U6798 ( .A(n54202), .B(n6239), .Z(n6240) );
  NAND U6799 ( .A(n54203), .B(n6240), .Z(n6241) );
  NANDN U6800 ( .A(n52152), .B(n6241), .Z(n6242) );
  NAND U6801 ( .A(n54204), .B(n6242), .Z(n6243) );
  ANDN U6802 ( .B(n6243), .A(n54205), .Z(n6244) );
  OR U6803 ( .A(n54206), .B(n6244), .Z(n6245) );
  NAND U6804 ( .A(n54207), .B(n6245), .Z(n6246) );
  NANDN U6805 ( .A(n52151), .B(n6246), .Z(n6247) );
  NAND U6806 ( .A(n54208), .B(n6247), .Z(n6248) );
  NANDN U6807 ( .A(n54209), .B(n6248), .Z(n6249) );
  ANDN U6808 ( .B(n6249), .A(n54210), .Z(n54212) );
  NANDN U6809 ( .A(n52147), .B(n54266), .Z(n6250) );
  NAND U6810 ( .A(n54267), .B(n6250), .Z(n6251) );
  NANDN U6811 ( .A(n52146), .B(n6251), .Z(n6252) );
  NAND U6812 ( .A(n54268), .B(n6252), .Z(n6253) );
  NAND U6813 ( .A(n54269), .B(n6253), .Z(n6254) );
  ANDN U6814 ( .B(n6254), .A(n54270), .Z(n6255) );
  NANDN U6815 ( .A(n6255), .B(n54271), .Z(n6256) );
  NANDN U6816 ( .A(n54272), .B(n6256), .Z(n6257) );
  NAND U6817 ( .A(n54273), .B(n6257), .Z(n6258) );
  NANDN U6818 ( .A(n54274), .B(n6258), .Z(n6259) );
  NAND U6819 ( .A(n54275), .B(n6259), .Z(n6260) );
  ANDN U6820 ( .B(n6260), .A(n54276), .Z(n6261) );
  NANDN U6821 ( .A(n6261), .B(n54277), .Z(n6262) );
  ANDN U6822 ( .B(n6262), .A(n54278), .Z(n6263) );
  OR U6823 ( .A(n6263), .B(n54279), .Z(n6264) );
  NAND U6824 ( .A(n54280), .B(n6264), .Z(n6265) );
  NANDN U6825 ( .A(n54281), .B(n6265), .Z(n54282) );
  NANDN U6826 ( .A(n54318), .B(n54317), .Z(n6266) );
  NAND U6827 ( .A(n54319), .B(n6266), .Z(n6267) );
  NANDN U6828 ( .A(n54320), .B(n6267), .Z(n6268) );
  NAND U6829 ( .A(n54321), .B(n6268), .Z(n6269) );
  NAND U6830 ( .A(n54322), .B(n6269), .Z(n6270) );
  ANDN U6831 ( .B(n6270), .A(n54323), .Z(n6271) );
  NANDN U6832 ( .A(n6271), .B(n54324), .Z(n6272) );
  NANDN U6833 ( .A(n54325), .B(n6272), .Z(n6273) );
  NAND U6834 ( .A(n54326), .B(n6273), .Z(n6274) );
  NANDN U6835 ( .A(n54327), .B(n6274), .Z(n6275) );
  NAND U6836 ( .A(n54328), .B(n6275), .Z(n6276) );
  ANDN U6837 ( .B(n6276), .A(n54329), .Z(n6277) );
  NANDN U6838 ( .A(n6277), .B(n54330), .Z(n6278) );
  ANDN U6839 ( .B(n6278), .A(n54331), .Z(n6279) );
  NANDN U6840 ( .A(n6279), .B(n54332), .Z(n6280) );
  NANDN U6841 ( .A(n54333), .B(n6280), .Z(n6281) );
  NAND U6842 ( .A(n54334), .B(n6281), .Z(n54335) );
  OR U6843 ( .A(n54358), .B(n54359), .Z(n6282) );
  NAND U6844 ( .A(n54360), .B(n6282), .Z(n6283) );
  ANDN U6845 ( .B(n6283), .A(n54361), .Z(n6284) );
  NANDN U6846 ( .A(n6284), .B(n54362), .Z(n6285) );
  NANDN U6847 ( .A(n54363), .B(n6285), .Z(n6286) );
  NAND U6848 ( .A(n52134), .B(n6286), .Z(n6287) );
  NANDN U6849 ( .A(n54364), .B(n6287), .Z(n6288) );
  NAND U6850 ( .A(n54365), .B(n6288), .Z(n6289) );
  ANDN U6851 ( .B(n6289), .A(n54366), .Z(n6290) );
  NANDN U6852 ( .A(n6290), .B(n54367), .Z(n6291) );
  NANDN U6853 ( .A(n52133), .B(n6291), .Z(n6292) );
  NANDN U6854 ( .A(n54368), .B(n6292), .Z(n6293) );
  NAND U6855 ( .A(n52132), .B(n6293), .Z(n54371) );
  NANDN U6856 ( .A(n54396), .B(n54395), .Z(n6294) );
  NAND U6857 ( .A(n54398), .B(n6294), .Z(n6295) );
  NAND U6858 ( .A(n54399), .B(n6295), .Z(n6296) );
  NANDN U6859 ( .A(n52124), .B(n6296), .Z(n6297) );
  NAND U6860 ( .A(n54400), .B(n6297), .Z(n6298) );
  AND U6861 ( .A(n54401), .B(n6298), .Z(n6299) );
  ANDN U6862 ( .B(n54403), .A(n54404), .Z(n6300) );
  NAND U6863 ( .A(n54402), .B(n6299), .Z(n6301) );
  AND U6864 ( .A(n6300), .B(n6301), .Z(n6302) );
  ANDN U6865 ( .B(n52122), .A(n6302), .Z(n6303) );
  NAND U6866 ( .A(n52123), .B(n6303), .Z(n6304) );
  AND U6867 ( .A(n54405), .B(n6304), .Z(n6305) );
  NAND U6868 ( .A(n6305), .B(n52121), .Z(n6306) );
  AND U6869 ( .A(n52120), .B(n6306), .Z(n6307) );
  NAND U6870 ( .A(n6307), .B(n52119), .Z(n6308) );
  ANDN U6871 ( .B(n6308), .A(n54406), .Z(n54407) );
  OR U6872 ( .A(n54436), .B(n54437), .Z(n6309) );
  NAND U6873 ( .A(n54438), .B(n6309), .Z(n6310) );
  NANDN U6874 ( .A(n54439), .B(n6310), .Z(n6311) );
  NAND U6875 ( .A(n54440), .B(n6311), .Z(n6312) );
  NANDN U6876 ( .A(n54441), .B(n6312), .Z(n6313) );
  ANDN U6877 ( .B(n6313), .A(n54442), .Z(n6314) );
  NANDN U6878 ( .A(n6314), .B(n54443), .Z(n6315) );
  NANDN U6879 ( .A(n52114), .B(n6315), .Z(n6316) );
  NAND U6880 ( .A(n52113), .B(n6316), .Z(n6317) );
  NANDN U6881 ( .A(n54444), .B(n6317), .Z(n6318) );
  NAND U6882 ( .A(n54445), .B(n6318), .Z(n6319) );
  ANDN U6883 ( .B(n6319), .A(n54446), .Z(n6320) );
  OR U6884 ( .A(n54447), .B(n6320), .Z(n6321) );
  NAND U6885 ( .A(n54448), .B(n6321), .Z(n6322) );
  NANDN U6886 ( .A(n54449), .B(n6322), .Z(n6323) );
  NAND U6887 ( .A(n54450), .B(n6323), .Z(n54451) );
  NAND U6888 ( .A(n54478), .B(n54479), .Z(n6324) );
  NANDN U6889 ( .A(n54480), .B(n6324), .Z(n6325) );
  NAND U6890 ( .A(n54481), .B(n6325), .Z(n6326) );
  AND U6891 ( .A(n6326), .B(n54484), .Z(n6327) );
  NANDN U6892 ( .A(n54483), .B(n54482), .Z(n6328) );
  AND U6893 ( .A(n6327), .B(n6328), .Z(n6329) );
  NAND U6894 ( .A(n54487), .B(n54486), .Z(n6330) );
  AND U6895 ( .A(n54485), .B(n6330), .Z(n6331) );
  NANDN U6896 ( .A(n6329), .B(n6331), .Z(n6332) );
  NANDN U6897 ( .A(n54488), .B(n6332), .Z(n6333) );
  NAND U6898 ( .A(n54489), .B(n6333), .Z(n6334) );
  AND U6899 ( .A(n52104), .B(n6334), .Z(n6335) );
  OR U6900 ( .A(n54490), .B(n6335), .Z(n6336) );
  NAND U6901 ( .A(n54491), .B(n6336), .Z(n6337) );
  NANDN U6902 ( .A(n52103), .B(n6337), .Z(n54492) );
  NANDN U6903 ( .A(n52094), .B(n54516), .Z(n6338) );
  NAND U6904 ( .A(n52093), .B(n6338), .Z(n6339) );
  NANDN U6905 ( .A(n54517), .B(n6339), .Z(n6340) );
  NAND U6906 ( .A(n54518), .B(n6340), .Z(n6341) );
  NANDN U6907 ( .A(n54519), .B(n6341), .Z(n6342) );
  AND U6908 ( .A(n54520), .B(n6342), .Z(n6343) );
  OR U6909 ( .A(n6343), .B(n54521), .Z(n6344) );
  NAND U6910 ( .A(n54522), .B(n6344), .Z(n6345) );
  AND U6911 ( .A(n54523), .B(n6345), .Z(n6346) );
  OR U6912 ( .A(n54524), .B(n6346), .Z(n6347) );
  NAND U6913 ( .A(n54525), .B(n6347), .Z(n6348) );
  NANDN U6914 ( .A(n54526), .B(n6348), .Z(n6349) );
  NAND U6915 ( .A(n54527), .B(n6349), .Z(n6350) );
  NANDN U6916 ( .A(n54528), .B(n6350), .Z(n6351) );
  AND U6917 ( .A(n54529), .B(n6351), .Z(n6352) );
  NANDN U6918 ( .A(n6352), .B(n54530), .Z(n6353) );
  NANDN U6919 ( .A(n54531), .B(n6353), .Z(n6354) );
  NAND U6920 ( .A(n54532), .B(n6354), .Z(n54533) );
  NAND U6921 ( .A(n54568), .B(n54567), .Z(n6355) );
  NANDN U6922 ( .A(n54569), .B(n6355), .Z(n6356) );
  ANDN U6923 ( .B(n6356), .A(n54570), .Z(n6357) );
  NANDN U6924 ( .A(n6357), .B(n54571), .Z(n6358) );
  NAND U6925 ( .A(n54572), .B(n6358), .Z(n6359) );
  NAND U6926 ( .A(n54573), .B(n6359), .Z(n6360) );
  NAND U6927 ( .A(n54574), .B(n6360), .Z(n6361) );
  NAND U6928 ( .A(n54575), .B(n6361), .Z(n6362) );
  ANDN U6929 ( .B(n6362), .A(n54576), .Z(n6363) );
  NANDN U6930 ( .A(n6363), .B(n52089), .Z(n6364) );
  NANDN U6931 ( .A(n54577), .B(n6364), .Z(n6365) );
  NAND U6932 ( .A(n54578), .B(n6365), .Z(n6366) );
  NANDN U6933 ( .A(n52088), .B(n6366), .Z(n54579) );
  NAND U6934 ( .A(n54616), .B(n54615), .Z(n6367) );
  NANDN U6935 ( .A(n54618), .B(n6367), .Z(n6368) );
  ANDN U6936 ( .B(n6368), .A(n52084), .Z(n6369) );
  AND U6937 ( .A(n54620), .B(n54621), .Z(n6370) );
  NANDN U6938 ( .A(n6369), .B(n54619), .Z(n6371) );
  AND U6939 ( .A(n6370), .B(n6371), .Z(n6372) );
  OR U6940 ( .A(n54622), .B(n6372), .Z(n6373) );
  NAND U6941 ( .A(n54623), .B(n6373), .Z(n6374) );
  NANDN U6942 ( .A(n52083), .B(n6374), .Z(n6375) );
  NAND U6943 ( .A(n52082), .B(n6375), .Z(n6376) );
  NAND U6944 ( .A(n54624), .B(n6376), .Z(n6377) );
  AND U6945 ( .A(n54625), .B(n6377), .Z(n6378) );
  OR U6946 ( .A(n54626), .B(n6378), .Z(n6379) );
  NAND U6947 ( .A(n54627), .B(n6379), .Z(n6380) );
  NANDN U6948 ( .A(n52081), .B(n6380), .Z(n54628) );
  NANDN U6949 ( .A(n54658), .B(n54657), .Z(n6381) );
  NANDN U6950 ( .A(n52073), .B(n6381), .Z(n6382) );
  NAND U6951 ( .A(n52072), .B(n6382), .Z(n6383) );
  NANDN U6952 ( .A(n54659), .B(n6383), .Z(n6384) );
  NANDN U6953 ( .A(n54660), .B(n6384), .Z(n6385) );
  AND U6954 ( .A(n54661), .B(n6385), .Z(n6386) );
  OR U6955 ( .A(n6386), .B(n54662), .Z(n6387) );
  NAND U6956 ( .A(n54663), .B(n6387), .Z(n6388) );
  ANDN U6957 ( .B(n6388), .A(n54664), .Z(n6389) );
  OR U6958 ( .A(n6389), .B(n54665), .Z(n6390) );
  NAND U6959 ( .A(n54666), .B(n6390), .Z(n6391) );
  NANDN U6960 ( .A(n54667), .B(n6391), .Z(n6392) );
  NAND U6961 ( .A(n54668), .B(n6392), .Z(n6393) );
  AND U6962 ( .A(n52071), .B(n6393), .Z(n6394) );
  NAND U6963 ( .A(n6394), .B(n52070), .Z(n6395) );
  NANDN U6964 ( .A(n54669), .B(n6395), .Z(n54670) );
  NAND U6965 ( .A(n54700), .B(n52067), .Z(n6396) );
  NANDN U6966 ( .A(n52066), .B(n6396), .Z(n6397) );
  AND U6967 ( .A(n52065), .B(n6397), .Z(n6398) );
  NANDN U6968 ( .A(n6398), .B(n54701), .Z(n6399) );
  NAND U6969 ( .A(n54702), .B(n6399), .Z(n6400) );
  NANDN U6970 ( .A(n54703), .B(n6400), .Z(n6401) );
  NAND U6971 ( .A(n54704), .B(n6401), .Z(n6402) );
  NANDN U6972 ( .A(n52064), .B(n6402), .Z(n6403) );
  ANDN U6973 ( .B(n6403), .A(n54705), .Z(n6404) );
  NANDN U6974 ( .A(n6404), .B(n54706), .Z(n6405) );
  NAND U6975 ( .A(n54707), .B(n6405), .Z(n6406) );
  NAND U6976 ( .A(n54708), .B(n6406), .Z(n54709) );
  NAND U6977 ( .A(n54733), .B(n54734), .Z(n6407) );
  NANDN U6978 ( .A(n54735), .B(n6407), .Z(n6408) );
  NAND U6979 ( .A(n54736), .B(n6408), .Z(n6409) );
  NAND U6980 ( .A(n52057), .B(n6409), .Z(n6410) );
  NANDN U6981 ( .A(n54737), .B(n6410), .Z(n6411) );
  AND U6982 ( .A(n54738), .B(n6411), .Z(n6412) );
  NANDN U6983 ( .A(n6412), .B(n54739), .Z(n6413) );
  NAND U6984 ( .A(n54740), .B(n6413), .Z(n6414) );
  NAND U6985 ( .A(n54741), .B(n6414), .Z(n6415) );
  NANDN U6986 ( .A(n54742), .B(n6415), .Z(n6416) );
  NAND U6987 ( .A(n54743), .B(n6416), .Z(n6417) );
  ANDN U6988 ( .B(n6417), .A(n54744), .Z(n6418) );
  OR U6989 ( .A(n52056), .B(n6418), .Z(n6419) );
  AND U6990 ( .A(n52055), .B(n6419), .Z(n6420) );
  OR U6991 ( .A(n54745), .B(n6420), .Z(n6421) );
  NAND U6992 ( .A(n54746), .B(n6421), .Z(n6422) );
  NANDN U6993 ( .A(n54747), .B(n6422), .Z(n54749) );
  NANDN U6994 ( .A(n54784), .B(n54783), .Z(n6423) );
  NAND U6995 ( .A(n54785), .B(n6423), .Z(n6424) );
  NAND U6996 ( .A(n54786), .B(n6424), .Z(n6425) );
  NANDN U6997 ( .A(n52051), .B(n6425), .Z(n6426) );
  NAND U6998 ( .A(n54787), .B(n6426), .Z(n6427) );
  ANDN U6999 ( .B(n6427), .A(n54788), .Z(n6428) );
  ANDN U7000 ( .B(n54790), .A(n6428), .Z(n6429) );
  NAND U7001 ( .A(n54789), .B(n6429), .Z(n6430) );
  ANDN U7002 ( .B(n6430), .A(n54791), .Z(n6431) );
  NOR U7003 ( .A(n52050), .B(n6431), .Z(n6432) );
  NAND U7004 ( .A(n54792), .B(n6432), .Z(n6433) );
  ANDN U7005 ( .B(n6433), .A(n54793), .Z(n6434) );
  NANDN U7006 ( .A(n6434), .B(n54794), .Z(n6435) );
  NANDN U7007 ( .A(n54795), .B(n6435), .Z(n6436) );
  NAND U7008 ( .A(n54796), .B(n6436), .Z(n54797) );
  NAND U7009 ( .A(n54819), .B(n54818), .Z(n6437) );
  NANDN U7010 ( .A(n54821), .B(n6437), .Z(n6438) );
  ANDN U7011 ( .B(n6438), .A(n52040), .Z(n6439) );
  OR U7012 ( .A(n6439), .B(n54822), .Z(n6440) );
  NAND U7013 ( .A(n52039), .B(n6440), .Z(n6441) );
  NANDN U7014 ( .A(n54823), .B(n6441), .Z(n6442) );
  NAND U7015 ( .A(n54824), .B(n6442), .Z(n6443) );
  NANDN U7016 ( .A(n52038), .B(n6443), .Z(n6444) );
  AND U7017 ( .A(n52037), .B(n6444), .Z(n6445) );
  OR U7018 ( .A(n6445), .B(n54825), .Z(n6446) );
  NANDN U7019 ( .A(n54826), .B(n6446), .Z(n6447) );
  NAND U7020 ( .A(n54827), .B(n6447), .Z(n54828) );
  NANDN U7021 ( .A(n52025), .B(n54850), .Z(n6448) );
  NANDN U7022 ( .A(n54851), .B(n6448), .Z(n6449) );
  AND U7023 ( .A(n54852), .B(n6449), .Z(n6450) );
  OR U7024 ( .A(n6450), .B(n54853), .Z(n6451) );
  NAND U7025 ( .A(n54854), .B(n6451), .Z(n6452) );
  ANDN U7026 ( .B(n6452), .A(n54855), .Z(n6453) );
  NANDN U7027 ( .A(n6453), .B(n54856), .Z(n6454) );
  NANDN U7028 ( .A(n54857), .B(n6454), .Z(n6455) );
  NANDN U7029 ( .A(n54858), .B(n6455), .Z(n6456) );
  NAND U7030 ( .A(n54859), .B(n6456), .Z(n6457) );
  NANDN U7031 ( .A(n54860), .B(n6457), .Z(n6458) );
  AND U7032 ( .A(n54861), .B(n6458), .Z(n6459) );
  OR U7033 ( .A(n6459), .B(n54862), .Z(n6460) );
  NANDN U7034 ( .A(n54863), .B(n6460), .Z(n6461) );
  NAND U7035 ( .A(n54864), .B(n6461), .Z(n6462) );
  NAND U7036 ( .A(n54865), .B(n6462), .Z(n54866) );
  NANDN U7037 ( .A(n53434), .B(n12512), .Z(n6463) );
  NAND U7038 ( .A(n53435), .B(n6463), .Z(n6464) );
  NANDN U7039 ( .A(n52292), .B(n6464), .Z(n6465) );
  NAND U7040 ( .A(n52291), .B(n6465), .Z(n6466) );
  NANDN U7041 ( .A(n52290), .B(n6466), .Z(n6467) );
  AND U7042 ( .A(n52289), .B(n6467), .Z(n6468) );
  OR U7043 ( .A(n53438), .B(n6468), .Z(n6469) );
  NAND U7044 ( .A(n53440), .B(n6469), .Z(n6470) );
  NANDN U7045 ( .A(n52288), .B(n6470), .Z(n6471) );
  NAND U7046 ( .A(n52287), .B(n6471), .Z(n6472) );
  NANDN U7047 ( .A(n53441), .B(n6472), .Z(n6473) );
  AND U7048 ( .A(n53442), .B(n6473), .Z(n6474) );
  NANDN U7049 ( .A(n6474), .B(n53443), .Z(n6475) );
  NANDN U7050 ( .A(n52286), .B(n6475), .Z(n6476) );
  NAND U7051 ( .A(n27890), .B(n6476), .Z(n6477) );
  NANDN U7052 ( .A(n6477), .B(n32973), .Z(n6478) );
  NAND U7053 ( .A(n53445), .B(n6478), .Z(n6479) );
  NAND U7054 ( .A(n27892), .B(n6479), .Z(n6480) );
  NANDN U7055 ( .A(n53447), .B(n6480), .Z(n12516) );
  NANDN U7056 ( .A(n54926), .B(n54925), .Z(n6481) );
  NAND U7057 ( .A(n54927), .B(n6481), .Z(n6482) );
  ANDN U7058 ( .B(n6482), .A(n54928), .Z(n6483) );
  NANDN U7059 ( .A(n6483), .B(n54929), .Z(n6484) );
  NANDN U7060 ( .A(n54930), .B(n6484), .Z(n6485) );
  NANDN U7061 ( .A(n52021), .B(n6485), .Z(n6486) );
  NAND U7062 ( .A(n54931), .B(n6486), .Z(n6487) );
  NANDN U7063 ( .A(n54932), .B(n6487), .Z(n6488) );
  AND U7064 ( .A(n54933), .B(n6488), .Z(n6489) );
  NANDN U7065 ( .A(n6489), .B(n54934), .Z(n6490) );
  NANDN U7066 ( .A(n54935), .B(n6490), .Z(n6491) );
  NAND U7067 ( .A(n54936), .B(n6491), .Z(n6492) );
  NANDN U7068 ( .A(n54937), .B(n6492), .Z(n6493) );
  NAND U7069 ( .A(n54938), .B(n6493), .Z(n6494) );
  ANDN U7070 ( .B(n6494), .A(n54939), .Z(n6495) );
  AND U7071 ( .A(n52019), .B(n52020), .Z(n6496) );
  NANDN U7072 ( .A(n6495), .B(n54940), .Z(n6497) );
  AND U7073 ( .A(n6496), .B(n6497), .Z(n54941) );
  OR U7074 ( .A(n54999), .B(n55000), .Z(n6498) );
  NAND U7075 ( .A(n55001), .B(n6498), .Z(n6499) );
  NANDN U7076 ( .A(n55002), .B(n6499), .Z(n6500) );
  NANDN U7077 ( .A(n52017), .B(n6500), .Z(n6501) );
  NAND U7078 ( .A(n52016), .B(n6501), .Z(n6502) );
  AND U7079 ( .A(n55003), .B(n6502), .Z(n6503) );
  NANDN U7080 ( .A(n52015), .B(n6503), .Z(n6504) );
  NANDN U7081 ( .A(n55004), .B(n6504), .Z(n6505) );
  AND U7082 ( .A(n55005), .B(n6505), .Z(n6506) );
  OR U7083 ( .A(n6506), .B(n55006), .Z(n6507) );
  NAND U7084 ( .A(n55007), .B(n6507), .Z(n6508) );
  ANDN U7085 ( .B(n6508), .A(n55008), .Z(n6509) );
  OR U7086 ( .A(n6509), .B(n55009), .Z(n6510) );
  ANDN U7087 ( .B(n6510), .A(n55010), .Z(n6511) );
  OR U7088 ( .A(n6511), .B(n55011), .Z(n6512) );
  NAND U7089 ( .A(n55012), .B(n6512), .Z(n6513) );
  NANDN U7090 ( .A(n55013), .B(n6513), .Z(n55014) );
  NANDN U7091 ( .A(n55047), .B(n55046), .Z(n6514) );
  NANDN U7092 ( .A(n55048), .B(n6514), .Z(n6515) );
  AND U7093 ( .A(n55049), .B(n6515), .Z(n6516) );
  OR U7094 ( .A(n6516), .B(n55050), .Z(n6517) );
  NAND U7095 ( .A(n55051), .B(n6517), .Z(n6518) );
  NAND U7096 ( .A(n55052), .B(n6518), .Z(n6519) );
  NANDN U7097 ( .A(n6519), .B(n55053), .Z(n6520) );
  NAND U7098 ( .A(n52011), .B(n6520), .Z(n6521) );
  NANDN U7099 ( .A(n55054), .B(n6521), .Z(n6522) );
  NAND U7100 ( .A(n55055), .B(n6522), .Z(n6523) );
  NANDN U7101 ( .A(n52010), .B(n6523), .Z(n6524) );
  AND U7102 ( .A(n52009), .B(n6524), .Z(n6525) );
  OR U7103 ( .A(n6525), .B(n55056), .Z(n6526) );
  AND U7104 ( .A(n55057), .B(n6526), .Z(n55059) );
  NANDN U7105 ( .A(n55079), .B(n55078), .Z(n6527) );
  NAND U7106 ( .A(n55081), .B(n6527), .Z(n6528) );
  AND U7107 ( .A(n55082), .B(n6528), .Z(n6529) );
  OR U7108 ( .A(n52000), .B(n6529), .Z(n6530) );
  NAND U7109 ( .A(n51999), .B(n6530), .Z(n6531) );
  NANDN U7110 ( .A(n55083), .B(n6531), .Z(n6532) );
  NANDN U7111 ( .A(n55084), .B(n6532), .Z(n6533) );
  NAND U7112 ( .A(n55085), .B(n6533), .Z(n6534) );
  ANDN U7113 ( .B(n6534), .A(n51998), .Z(n6535) );
  NANDN U7114 ( .A(n6535), .B(n51997), .Z(n6536) );
  NANDN U7115 ( .A(n55086), .B(n6536), .Z(n6537) );
  NAND U7116 ( .A(n55087), .B(n6537), .Z(n6538) );
  NANDN U7117 ( .A(n55088), .B(n6538), .Z(n55089) );
  NAND U7118 ( .A(n55113), .B(n51990), .Z(n6539) );
  NANDN U7119 ( .A(n55114), .B(n6539), .Z(n6540) );
  ANDN U7120 ( .B(n6540), .A(n55115), .Z(n6541) );
  NANDN U7121 ( .A(n6541), .B(n55116), .Z(n6542) );
  NANDN U7122 ( .A(n55117), .B(n6542), .Z(n6543) );
  NAND U7123 ( .A(n55118), .B(n6543), .Z(n6544) );
  NANDN U7124 ( .A(n55119), .B(n6544), .Z(n6545) );
  NANDN U7125 ( .A(n55120), .B(n6545), .Z(n6546) );
  AND U7126 ( .A(n55121), .B(n6546), .Z(n6547) );
  OR U7127 ( .A(n6547), .B(n55122), .Z(n6548) );
  NAND U7128 ( .A(n55123), .B(n6548), .Z(n6549) );
  ANDN U7129 ( .B(n6549), .A(n55124), .Z(n6550) );
  OR U7130 ( .A(n6550), .B(n55125), .Z(n6551) );
  AND U7131 ( .A(n55126), .B(n6551), .Z(n6552) );
  OR U7132 ( .A(n6552), .B(n55127), .Z(n6553) );
  NAND U7133 ( .A(n55128), .B(n6553), .Z(n6554) );
  NANDN U7134 ( .A(n55129), .B(n6554), .Z(n55130) );
  OR U7135 ( .A(n55195), .B(n55194), .Z(n6555) );
  NAND U7136 ( .A(n55196), .B(n6555), .Z(n6556) );
  ANDN U7137 ( .B(n6556), .A(n55197), .Z(n6557) );
  OR U7138 ( .A(n6557), .B(n55198), .Z(n6558) );
  NAND U7139 ( .A(n55199), .B(n6558), .Z(n6559) );
  AND U7140 ( .A(n55200), .B(n6559), .Z(n6560) );
  OR U7141 ( .A(n51980), .B(n6560), .Z(n6561) );
  NAND U7142 ( .A(n51979), .B(n6561), .Z(n6562) );
  NANDN U7143 ( .A(n55201), .B(n6562), .Z(n6563) );
  NAND U7144 ( .A(n55202), .B(n6563), .Z(n6564) );
  NANDN U7145 ( .A(n55203), .B(n6564), .Z(n6565) );
  AND U7146 ( .A(n55204), .B(n6565), .Z(n6566) );
  OR U7147 ( .A(n6566), .B(n55205), .Z(n6567) );
  ANDN U7148 ( .B(n6567), .A(n55206), .Z(n6568) );
  NANDN U7149 ( .A(n6568), .B(n55207), .Z(n6569) );
  NANDN U7150 ( .A(n55208), .B(n6569), .Z(n6570) );
  NAND U7151 ( .A(n55209), .B(n6570), .Z(n55210) );
  OR U7152 ( .A(n55269), .B(n55270), .Z(n6571) );
  AND U7153 ( .A(n55271), .B(n6571), .Z(n6572) );
  ANDN U7154 ( .B(n55275), .A(n6572), .Z(n6573) );
  NAND U7155 ( .A(n55274), .B(n6573), .Z(n6574) );
  ANDN U7156 ( .B(n6574), .A(n55276), .Z(n6575) );
  NANDN U7157 ( .A(n6575), .B(n55277), .Z(n6576) );
  ANDN U7158 ( .B(n6576), .A(n55278), .Z(n6577) );
  ANDN U7159 ( .B(n55280), .A(n6577), .Z(n6578) );
  NAND U7160 ( .A(n55279), .B(n6578), .Z(n6579) );
  ANDN U7161 ( .B(n6579), .A(n55281), .Z(n6580) );
  NANDN U7162 ( .A(n6580), .B(n55282), .Z(n6581) );
  NANDN U7163 ( .A(n55283), .B(n6581), .Z(n6582) );
  NAND U7164 ( .A(n55284), .B(n6582), .Z(n6583) );
  OR U7165 ( .A(n6583), .B(n55285), .Z(n6584) );
  NANDN U7166 ( .A(n55286), .B(n6584), .Z(n6585) );
  NAND U7167 ( .A(n55287), .B(n6585), .Z(n55288) );
  NAND U7168 ( .A(n51968), .B(n55308), .Z(n6586) );
  NANDN U7169 ( .A(n55309), .B(n6586), .Z(n6587) );
  AND U7170 ( .A(n55310), .B(n6587), .Z(n6588) );
  NOR U7171 ( .A(n55311), .B(n6588), .Z(n6589) );
  NAND U7172 ( .A(n51967), .B(n6589), .Z(n6590) );
  AND U7173 ( .A(n55312), .B(n6590), .Z(n6591) );
  OR U7174 ( .A(n55313), .B(n6591), .Z(n6592) );
  AND U7175 ( .A(n55314), .B(n6592), .Z(n6593) );
  OR U7176 ( .A(n55315), .B(n6593), .Z(n6594) );
  NAND U7177 ( .A(n55316), .B(n6594), .Z(n6595) );
  NANDN U7178 ( .A(n55317), .B(n6595), .Z(n6596) );
  NAND U7179 ( .A(n55318), .B(n6596), .Z(n6597) );
  AND U7180 ( .A(n55320), .B(n6597), .Z(n6598) );
  NAND U7181 ( .A(n6598), .B(n55319), .Z(n55321) );
  NANDN U7182 ( .A(n55399), .B(n55398), .Z(n6599) );
  NANDN U7183 ( .A(n55400), .B(n6599), .Z(n6600) );
  AND U7184 ( .A(n55401), .B(n6600), .Z(n6601) );
  OR U7185 ( .A(n6601), .B(n55402), .Z(n6602) );
  NAND U7186 ( .A(n55403), .B(n6602), .Z(n6603) );
  ANDN U7187 ( .B(n6603), .A(n55404), .Z(n6604) );
  OR U7188 ( .A(n6604), .B(n55405), .Z(n6605) );
  NAND U7189 ( .A(n55406), .B(n6605), .Z(n6606) );
  ANDN U7190 ( .B(n6606), .A(n55407), .Z(n6607) );
  NANDN U7191 ( .A(n6607), .B(n55408), .Z(n6608) );
  NANDN U7192 ( .A(n55409), .B(n6608), .Z(n6609) );
  NANDN U7193 ( .A(n55410), .B(n6609), .Z(n6610) );
  AND U7194 ( .A(n55411), .B(n6610), .Z(n6611) );
  AND U7195 ( .A(n51962), .B(n51963), .Z(n6612) );
  OR U7196 ( .A(n6611), .B(n55412), .Z(n6613) );
  AND U7197 ( .A(n6612), .B(n6613), .Z(n6614) );
  OR U7198 ( .A(n6614), .B(n55413), .Z(n6615) );
  NAND U7199 ( .A(n55414), .B(n6615), .Z(n6616) );
  NAND U7200 ( .A(n55415), .B(n6616), .Z(n55417) );
  NAND U7201 ( .A(n55447), .B(n55446), .Z(n6617) );
  AND U7202 ( .A(n51954), .B(n6617), .Z(n6618) );
  NAND U7203 ( .A(n6618), .B(n51955), .Z(n6619) );
  NANDN U7204 ( .A(n55448), .B(n6619), .Z(n6620) );
  NAND U7205 ( .A(n55449), .B(n6620), .Z(n6621) );
  ANDN U7206 ( .B(n6621), .A(n55450), .Z(n6622) );
  OR U7207 ( .A(n51953), .B(n6622), .Z(n6623) );
  AND U7208 ( .A(n51952), .B(n6623), .Z(n6624) );
  AND U7209 ( .A(n51950), .B(n51951), .Z(n6625) );
  NANDN U7210 ( .A(n6624), .B(n55451), .Z(n6626) );
  AND U7211 ( .A(n6625), .B(n6626), .Z(n6627) );
  NANDN U7212 ( .A(n6627), .B(n55452), .Z(n6628) );
  NANDN U7213 ( .A(n51949), .B(n6628), .Z(n6629) );
  NAND U7214 ( .A(n51948), .B(n6629), .Z(n55453) );
  NANDN U7215 ( .A(x[1920]), .B(y[1920]), .Z(n6630) );
  ANDN U7216 ( .B(n6630), .A(n13276), .Z(n34305) );
  NANDN U7217 ( .A(n55475), .B(n55474), .Z(n6631) );
  NAND U7218 ( .A(n55477), .B(n6631), .Z(n6632) );
  AND U7219 ( .A(n55478), .B(n6632), .Z(n6633) );
  NOR U7220 ( .A(n6633), .B(n55480), .Z(n6634) );
  NAND U7221 ( .A(n55479), .B(n6634), .Z(n6635) );
  ANDN U7222 ( .B(n6635), .A(n55481), .Z(n6636) );
  NANDN U7223 ( .A(n6636), .B(n55482), .Z(n6637) );
  NANDN U7224 ( .A(n51939), .B(n6637), .Z(n6638) );
  NANDN U7225 ( .A(n55483), .B(n6638), .Z(n6639) );
  NAND U7226 ( .A(n55484), .B(n6639), .Z(n6640) );
  NANDN U7227 ( .A(n55485), .B(n6640), .Z(n6641) );
  AND U7228 ( .A(n55486), .B(n6641), .Z(n6642) );
  OR U7229 ( .A(n6642), .B(n55487), .Z(n6643) );
  NANDN U7230 ( .A(n51938), .B(n6643), .Z(n6644) );
  NAND U7231 ( .A(n51937), .B(n6644), .Z(n55490) );
  AND U7232 ( .A(n51928), .B(n51929), .Z(n6645) );
  NAND U7233 ( .A(n55508), .B(n55509), .Z(n6646) );
  AND U7234 ( .A(n6645), .B(n6646), .Z(n6647) );
  OR U7235 ( .A(n6647), .B(n55510), .Z(n6648) );
  NAND U7236 ( .A(n55511), .B(n6648), .Z(n6649) );
  ANDN U7237 ( .B(n6649), .A(n55512), .Z(n6650) );
  NANDN U7238 ( .A(n6650), .B(n51927), .Z(n6651) );
  NANDN U7239 ( .A(n55513), .B(n6651), .Z(n6652) );
  NANDN U7240 ( .A(n55514), .B(n6652), .Z(n6653) );
  NAND U7241 ( .A(n55515), .B(n6653), .Z(n6654) );
  NANDN U7242 ( .A(n55516), .B(n6654), .Z(n6655) );
  AND U7243 ( .A(n51926), .B(n6655), .Z(n6656) );
  OR U7244 ( .A(n55517), .B(n6656), .Z(n6657) );
  NANDN U7245 ( .A(n55518), .B(n6657), .Z(n6658) );
  NAND U7246 ( .A(n55519), .B(n6658), .Z(n6659) );
  NANDN U7247 ( .A(n55520), .B(n6659), .Z(n55521) );
  NAND U7248 ( .A(n55545), .B(n55544), .Z(n6660) );
  NANDN U7249 ( .A(n55546), .B(n6660), .Z(n6661) );
  NAND U7250 ( .A(n51918), .B(n6661), .Z(n6662) );
  NANDN U7251 ( .A(n55547), .B(n6662), .Z(n6663) );
  NAND U7252 ( .A(n55548), .B(n6663), .Z(n6664) );
  ANDN U7253 ( .B(n6664), .A(n51917), .Z(n6665) );
  OR U7254 ( .A(n6665), .B(n55549), .Z(n6666) );
  NAND U7255 ( .A(n51916), .B(n6666), .Z(n6667) );
  ANDN U7256 ( .B(n6667), .A(n55550), .Z(n6668) );
  NANDN U7257 ( .A(n6668), .B(n55551), .Z(n6669) );
  NANDN U7258 ( .A(n51915), .B(n6669), .Z(n6670) );
  NANDN U7259 ( .A(n55552), .B(n6670), .Z(n55553) );
  NANDN U7260 ( .A(n55572), .B(n55571), .Z(n6671) );
  NAND U7261 ( .A(n55573), .B(n6671), .Z(n6672) );
  NAND U7262 ( .A(n51905), .B(n6672), .Z(n6673) );
  NANDN U7263 ( .A(n55574), .B(n6673), .Z(n6674) );
  NANDN U7264 ( .A(n55575), .B(n6674), .Z(n6675) );
  AND U7265 ( .A(n55576), .B(n6675), .Z(n6676) );
  OR U7266 ( .A(n6676), .B(n55577), .Z(n6677) );
  NANDN U7267 ( .A(n55578), .B(n6677), .Z(n6678) );
  AND U7268 ( .A(n55579), .B(n6678), .Z(n6679) );
  OR U7269 ( .A(n51904), .B(n6679), .Z(n6680) );
  AND U7270 ( .A(n51903), .B(n6680), .Z(n6681) );
  AND U7271 ( .A(n51900), .B(n51901), .Z(n6682) );
  OR U7272 ( .A(n51902), .B(n6681), .Z(n6683) );
  AND U7273 ( .A(n6682), .B(n6683), .Z(n55582) );
  OR U7274 ( .A(n55601), .B(n55602), .Z(n6684) );
  NAND U7275 ( .A(n55603), .B(n6684), .Z(n6685) );
  AND U7276 ( .A(n55604), .B(n6685), .Z(n6686) );
  NANDN U7277 ( .A(n55605), .B(n6686), .Z(n6687) );
  NAND U7278 ( .A(n51891), .B(n6687), .Z(n6688) );
  ANDN U7279 ( .B(n6688), .A(n55606), .Z(n6689) );
  NANDN U7280 ( .A(n6689), .B(n55607), .Z(n6690) );
  ANDN U7281 ( .B(n6690), .A(n51890), .Z(n6691) );
  OR U7282 ( .A(n6691), .B(n55608), .Z(n6692) );
  NAND U7283 ( .A(n51889), .B(n6692), .Z(n6693) );
  NAND U7284 ( .A(n55609), .B(n6693), .Z(n6694) );
  AND U7285 ( .A(n55610), .B(n55611), .Z(n6695) );
  NAND U7286 ( .A(n6694), .B(n6695), .Z(n6696) );
  NAND U7287 ( .A(n51888), .B(n6696), .Z(n55614) );
  OR U7288 ( .A(n55646), .B(n55645), .Z(n6697) );
  NAND U7289 ( .A(n55647), .B(n6697), .Z(n6698) );
  NANDN U7290 ( .A(n55648), .B(n6698), .Z(n6699) );
  AND U7291 ( .A(n55650), .B(n55649), .Z(n6700) );
  NAND U7292 ( .A(n6699), .B(n6700), .Z(n6701) );
  NAND U7293 ( .A(n55651), .B(n6701), .Z(n6702) );
  NANDN U7294 ( .A(n55652), .B(n6702), .Z(n6703) );
  NAND U7295 ( .A(n55653), .B(n6703), .Z(n6704) );
  ANDN U7296 ( .B(n6704), .A(n55654), .Z(n6705) );
  OR U7297 ( .A(n55655), .B(n6705), .Z(n6706) );
  AND U7298 ( .A(n55656), .B(n6706), .Z(n6707) );
  AND U7299 ( .A(n55659), .B(n55658), .Z(n6708) );
  NANDN U7300 ( .A(n6707), .B(n55657), .Z(n6709) );
  AND U7301 ( .A(n6708), .B(n6709), .Z(n6710) );
  NANDN U7302 ( .A(n6710), .B(n55660), .Z(n6711) );
  NANDN U7303 ( .A(n55661), .B(n6711), .Z(n6712) );
  NAND U7304 ( .A(n55662), .B(n6712), .Z(n55663) );
  NANDN U7305 ( .A(y[2211]), .B(x[2211]), .Z(n6713) );
  ANDN U7306 ( .B(n6713), .A(n13659), .Z(n27242) );
  NANDN U7307 ( .A(n55761), .B(n55760), .Z(n6714) );
  ANDN U7308 ( .B(n6714), .A(n55762), .Z(n6715) );
  NANDN U7309 ( .A(n6715), .B(n55763), .Z(n6716) );
  NAND U7310 ( .A(n55764), .B(n6716), .Z(n6717) );
  NAND U7311 ( .A(n55765), .B(n6717), .Z(n6718) );
  AND U7312 ( .A(n6718), .B(n55766), .Z(n6719) );
  NANDN U7313 ( .A(n51877), .B(n51878), .Z(n6720) );
  AND U7314 ( .A(n6719), .B(n6720), .Z(n6721) );
  NANDN U7315 ( .A(n6721), .B(n55767), .Z(n6722) );
  NANDN U7316 ( .A(n55768), .B(n6722), .Z(n6723) );
  NAND U7317 ( .A(n55769), .B(n6723), .Z(n6724) );
  NANDN U7318 ( .A(n55770), .B(n6724), .Z(n6725) );
  NAND U7319 ( .A(n55771), .B(n6725), .Z(n6726) );
  ANDN U7320 ( .B(n6726), .A(n55772), .Z(n6727) );
  NANDN U7321 ( .A(n6727), .B(n55773), .Z(n6728) );
  AND U7322 ( .A(n55774), .B(n6728), .Z(n6729) );
  NAND U7323 ( .A(n55775), .B(n6729), .Z(n6730) );
  NAND U7324 ( .A(n55776), .B(n6730), .Z(n6731) );
  NANDN U7325 ( .A(n55777), .B(n6731), .Z(n55778) );
  AND U7326 ( .A(n55801), .B(n55800), .Z(n6732) );
  NAND U7327 ( .A(n51867), .B(n55799), .Z(n6733) );
  AND U7328 ( .A(n6732), .B(n6733), .Z(n6734) );
  NANDN U7329 ( .A(n6734), .B(n55802), .Z(n6735) );
  ANDN U7330 ( .B(n6735), .A(n55803), .Z(n6736) );
  NANDN U7331 ( .A(n6736), .B(n55804), .Z(n6737) );
  NANDN U7332 ( .A(n55805), .B(n6737), .Z(n6738) );
  NAND U7333 ( .A(n55806), .B(n6738), .Z(n6739) );
  AND U7334 ( .A(n51866), .B(n51865), .Z(n6740) );
  NAND U7335 ( .A(n6739), .B(n6740), .Z(n6741) );
  NAND U7336 ( .A(n55807), .B(n6741), .Z(n6742) );
  NANDN U7337 ( .A(n51864), .B(n6742), .Z(n6743) );
  NAND U7338 ( .A(n55808), .B(n6743), .Z(n6744) );
  ANDN U7339 ( .B(n6744), .A(n55809), .Z(n6745) );
  NANDN U7340 ( .A(n6745), .B(n55810), .Z(n6746) );
  NANDN U7341 ( .A(n55811), .B(n6746), .Z(n6747) );
  NAND U7342 ( .A(n55812), .B(n6747), .Z(n55813) );
  NANDN U7343 ( .A(n55844), .B(n55843), .Z(n6748) );
  ANDN U7344 ( .B(n6748), .A(n51858), .Z(n6749) );
  NANDN U7345 ( .A(n6749), .B(n55845), .Z(n6750) );
  NANDN U7346 ( .A(n55846), .B(n6750), .Z(n6751) );
  NAND U7347 ( .A(n55847), .B(n6751), .Z(n6752) );
  AND U7348 ( .A(n55848), .B(n55849), .Z(n6753) );
  NAND U7349 ( .A(n6752), .B(n6753), .Z(n6754) );
  NANDN U7350 ( .A(n55850), .B(n6754), .Z(n6755) );
  NAND U7351 ( .A(n55851), .B(n6755), .Z(n6756) );
  NANDN U7352 ( .A(n55852), .B(n6756), .Z(n6757) );
  AND U7353 ( .A(n55853), .B(n6757), .Z(n6758) );
  OR U7354 ( .A(n6758), .B(n55854), .Z(n6759) );
  NAND U7355 ( .A(n55855), .B(n6759), .Z(n6760) );
  AND U7356 ( .A(n55856), .B(n6760), .Z(n6761) );
  OR U7357 ( .A(n6761), .B(n55857), .Z(n6762) );
  NAND U7358 ( .A(n55858), .B(n6762), .Z(n6763) );
  NANDN U7359 ( .A(n55859), .B(n6763), .Z(n6764) );
  NAND U7360 ( .A(n51857), .B(n6764), .Z(n55862) );
  NAND U7361 ( .A(n55884), .B(n51848), .Z(n6765) );
  NANDN U7362 ( .A(n55885), .B(n6765), .Z(n6766) );
  AND U7363 ( .A(n55886), .B(n6766), .Z(n6767) );
  OR U7364 ( .A(n51847), .B(n6767), .Z(n6768) );
  NAND U7365 ( .A(n51846), .B(n6768), .Z(n6769) );
  NANDN U7366 ( .A(n55887), .B(n6769), .Z(n6770) );
  NAND U7367 ( .A(n55888), .B(n6770), .Z(n6771) );
  AND U7368 ( .A(n51845), .B(n6771), .Z(n6772) );
  NAND U7369 ( .A(n6772), .B(n51844), .Z(n6773) );
  NAND U7370 ( .A(n55889), .B(n6773), .Z(n6774) );
  NANDN U7371 ( .A(n51843), .B(n6774), .Z(n55890) );
  NAND U7372 ( .A(n55912), .B(n55911), .Z(n6775) );
  ANDN U7373 ( .B(n6775), .A(n55913), .Z(n6776) );
  ANDN U7374 ( .B(n55915), .A(n6776), .Z(n6777) );
  NAND U7375 ( .A(n55914), .B(n6777), .Z(n6778) );
  ANDN U7376 ( .B(n6778), .A(n55916), .Z(n6779) );
  NANDN U7377 ( .A(n6779), .B(n55917), .Z(n6780) );
  NANDN U7378 ( .A(n51834), .B(n6780), .Z(n6781) );
  NAND U7379 ( .A(n51833), .B(n6781), .Z(n6782) );
  ANDN U7380 ( .B(n55920), .A(n55919), .Z(n6783) );
  NANDN U7381 ( .A(n55918), .B(n6782), .Z(n6784) );
  NAND U7382 ( .A(n6783), .B(n6784), .Z(n6785) );
  ANDN U7383 ( .B(n6785), .A(n55921), .Z(n55923) );
  NAND U7384 ( .A(n51824), .B(n55942), .Z(n6786) );
  NANDN U7385 ( .A(n55943), .B(n6786), .Z(n6787) );
  AND U7386 ( .A(n55944), .B(n6787), .Z(n6788) );
  OR U7387 ( .A(n51823), .B(n6788), .Z(n6789) );
  AND U7388 ( .A(n51822), .B(n6789), .Z(n6790) );
  AND U7389 ( .A(n55947), .B(n55946), .Z(n6791) );
  OR U7390 ( .A(n55945), .B(n6790), .Z(n6792) );
  AND U7391 ( .A(n6791), .B(n6792), .Z(n6793) );
  OR U7392 ( .A(n55948), .B(n6793), .Z(n6794) );
  NAND U7393 ( .A(n55949), .B(n6794), .Z(n6795) );
  NANDN U7394 ( .A(n51821), .B(n6795), .Z(n55950) );
  NANDN U7395 ( .A(n55977), .B(n55976), .Z(n6796) );
  NANDN U7396 ( .A(n55978), .B(n6796), .Z(n6797) );
  AND U7397 ( .A(n55979), .B(n6797), .Z(n6798) );
  OR U7398 ( .A(n6798), .B(n55980), .Z(n6799) );
  NAND U7399 ( .A(n55981), .B(n6799), .Z(n6800) );
  NANDN U7400 ( .A(n55982), .B(n6800), .Z(n6801) );
  AND U7401 ( .A(n55984), .B(n55983), .Z(n6802) );
  NAND U7402 ( .A(n6801), .B(n6802), .Z(n6803) );
  NAND U7403 ( .A(n55985), .B(n6803), .Z(n6804) );
  AND U7404 ( .A(n51814), .B(n51813), .Z(n6805) );
  NAND U7405 ( .A(n6804), .B(n6805), .Z(n6806) );
  NAND U7406 ( .A(n55986), .B(n6806), .Z(n6807) );
  NANDN U7407 ( .A(n51812), .B(n6807), .Z(n6808) );
  NAND U7408 ( .A(n51811), .B(n6808), .Z(n6809) );
  ANDN U7409 ( .B(n6809), .A(n55987), .Z(n55989) );
  NAND U7410 ( .A(n56010), .B(n56009), .Z(n6810) );
  NANDN U7411 ( .A(n56011), .B(n6810), .Z(n6811) );
  AND U7412 ( .A(n56012), .B(n6811), .Z(n6812) );
  OR U7413 ( .A(n6812), .B(n56013), .Z(n6813) );
  NAND U7414 ( .A(n51803), .B(n6813), .Z(n6814) );
  ANDN U7415 ( .B(n6814), .A(n56014), .Z(n6815) );
  NANDN U7416 ( .A(n6815), .B(n56015), .Z(n6816) );
  NANDN U7417 ( .A(n51802), .B(n6816), .Z(n6817) );
  NAND U7418 ( .A(n51801), .B(n6817), .Z(n6818) );
  AND U7419 ( .A(n56017), .B(n56016), .Z(n6819) );
  NAND U7420 ( .A(n6818), .B(n6819), .Z(n6820) );
  NANDN U7421 ( .A(n51800), .B(n6820), .Z(n56018) );
  NANDN U7422 ( .A(n56053), .B(n56052), .Z(n6821) );
  NAND U7423 ( .A(n56054), .B(n6821), .Z(n6822) );
  ANDN U7424 ( .B(n6822), .A(n56055), .Z(n6823) );
  NANDN U7425 ( .A(n6823), .B(n51796), .Z(n6824) );
  NANDN U7426 ( .A(n56056), .B(n6824), .Z(n6825) );
  NAND U7427 ( .A(n56057), .B(n6825), .Z(n6826) );
  NANDN U7428 ( .A(n51795), .B(n6826), .Z(n6827) );
  NAND U7429 ( .A(n51794), .B(n6827), .Z(n6828) );
  ANDN U7430 ( .B(n6828), .A(n56058), .Z(n6829) );
  NANDN U7431 ( .A(n6829), .B(n56059), .Z(n6830) );
  ANDN U7432 ( .B(n6830), .A(n56060), .Z(n56063) );
  OR U7433 ( .A(n56082), .B(n56083), .Z(n6831) );
  NAND U7434 ( .A(n56084), .B(n6831), .Z(n6832) );
  ANDN U7435 ( .B(n6832), .A(n56085), .Z(n6833) );
  AND U7436 ( .A(n56088), .B(n56087), .Z(n6834) );
  NANDN U7437 ( .A(n6833), .B(n56086), .Z(n6835) );
  AND U7438 ( .A(n6834), .B(n6835), .Z(n6836) );
  AND U7439 ( .A(n56091), .B(n56090), .Z(n6837) );
  OR U7440 ( .A(n56089), .B(n6836), .Z(n6838) );
  AND U7441 ( .A(n6837), .B(n6838), .Z(n6839) );
  NANDN U7442 ( .A(n6839), .B(n51784), .Z(n6840) );
  ANDN U7443 ( .B(n6840), .A(n56092), .Z(n6841) );
  NANDN U7444 ( .A(n6841), .B(n56093), .Z(n6842) );
  NANDN U7445 ( .A(n51783), .B(n6842), .Z(n6843) );
  NAND U7446 ( .A(n51782), .B(n6843), .Z(n56096) );
  NANDN U7447 ( .A(n56118), .B(n56117), .Z(n6844) );
  NAND U7448 ( .A(n56119), .B(n6844), .Z(n6845) );
  AND U7449 ( .A(n56120), .B(n6845), .Z(n6846) );
  NAND U7450 ( .A(n6846), .B(n56121), .Z(n6847) );
  NANDN U7451 ( .A(n56122), .B(n6847), .Z(n6848) );
  AND U7452 ( .A(n56123), .B(n6848), .Z(n6849) );
  AND U7453 ( .A(n51775), .B(n51774), .Z(n6850) );
  OR U7454 ( .A(n56124), .B(n6849), .Z(n6851) );
  AND U7455 ( .A(n6850), .B(n6851), .Z(n6852) );
  ANDN U7456 ( .B(n56126), .A(n56127), .Z(n6853) );
  NANDN U7457 ( .A(n6852), .B(n56125), .Z(n6854) );
  AND U7458 ( .A(n6853), .B(n6854), .Z(n6855) );
  AND U7459 ( .A(n56129), .B(n56128), .Z(n6856) );
  NANDN U7460 ( .A(n6855), .B(n51773), .Z(n6857) );
  AND U7461 ( .A(n6856), .B(n6857), .Z(n6858) );
  OR U7462 ( .A(n56130), .B(n6858), .Z(n6859) );
  NAND U7463 ( .A(n56131), .B(n6859), .Z(n6860) );
  NANDN U7464 ( .A(n56132), .B(n6860), .Z(n56133) );
  NANDN U7465 ( .A(n56158), .B(n56157), .Z(n6861) );
  NANDN U7466 ( .A(n56159), .B(n6861), .Z(n6862) );
  NAND U7467 ( .A(n56160), .B(n6862), .Z(n6863) );
  NAND U7468 ( .A(n56161), .B(n6863), .Z(n6864) );
  NANDN U7469 ( .A(n56162), .B(n6864), .Z(n6865) );
  AND U7470 ( .A(n56163), .B(n6865), .Z(n6866) );
  OR U7471 ( .A(n6866), .B(n56164), .Z(n6867) );
  NAND U7472 ( .A(n56165), .B(n6867), .Z(n6868) );
  ANDN U7473 ( .B(n6868), .A(n56166), .Z(n6869) );
  NANDN U7474 ( .A(n6869), .B(n51765), .Z(n6870) );
  NANDN U7475 ( .A(n56167), .B(n6870), .Z(n6871) );
  NAND U7476 ( .A(n56168), .B(n6871), .Z(n6872) );
  NANDN U7477 ( .A(n51764), .B(n6872), .Z(n56169) );
  NANDN U7478 ( .A(n51756), .B(n56193), .Z(n6873) );
  NAND U7479 ( .A(n51755), .B(n6873), .Z(n6874) );
  AND U7480 ( .A(n56194), .B(n6874), .Z(n6875) );
  NANDN U7481 ( .A(n51753), .B(n51752), .Z(n6876) );
  AND U7482 ( .A(n51754), .B(n6876), .Z(n6877) );
  NANDN U7483 ( .A(n6875), .B(n56195), .Z(n6878) );
  NAND U7484 ( .A(n6877), .B(n6878), .Z(n6879) );
  NANDN U7485 ( .A(n56196), .B(n6879), .Z(n6880) );
  NAND U7486 ( .A(n56197), .B(n6880), .Z(n6881) );
  NANDN U7487 ( .A(n56198), .B(n6881), .Z(n6882) );
  AND U7488 ( .A(n56199), .B(n6882), .Z(n6883) );
  NAND U7489 ( .A(n6883), .B(n56200), .Z(n6884) );
  NANDN U7490 ( .A(n56201), .B(n6884), .Z(n6885) );
  AND U7491 ( .A(n56202), .B(n6885), .Z(n6886) );
  OR U7492 ( .A(n56203), .B(n6886), .Z(n6887) );
  NAND U7493 ( .A(n56204), .B(n6887), .Z(n6888) );
  NANDN U7494 ( .A(n56205), .B(n6888), .Z(n6889) );
  AND U7495 ( .A(n56206), .B(n6889), .Z(n56209) );
  OR U7496 ( .A(n56231), .B(n56232), .Z(n6890) );
  NAND U7497 ( .A(n56233), .B(n6890), .Z(n6891) );
  ANDN U7498 ( .B(n6891), .A(n56234), .Z(n6892) );
  ANDN U7499 ( .B(n56236), .A(n6892), .Z(n6893) );
  NAND U7500 ( .A(n56235), .B(n6893), .Z(n6894) );
  ANDN U7501 ( .B(n6894), .A(n56237), .Z(n6895) );
  ANDN U7502 ( .B(n51744), .A(n6895), .Z(n6896) );
  NAND U7503 ( .A(n51743), .B(n6896), .Z(n6897) );
  ANDN U7504 ( .B(n6897), .A(n56238), .Z(n6898) );
  NANDN U7505 ( .A(n6898), .B(n56239), .Z(n6899) );
  NANDN U7506 ( .A(n56240), .B(n6899), .Z(n6900) );
  NAND U7507 ( .A(n56241), .B(n6900), .Z(n6901) );
  NANDN U7508 ( .A(n6901), .B(n56242), .Z(n6902) );
  ANDN U7509 ( .B(n6902), .A(n56243), .Z(n6903) );
  ANDN U7510 ( .B(n51741), .A(n6903), .Z(n6904) );
  NAND U7511 ( .A(n51742), .B(n6904), .Z(n6905) );
  ANDN U7512 ( .B(n6905), .A(n56244), .Z(n56248) );
  ANDN U7513 ( .B(n56268), .A(n56269), .Z(n6906) );
  ANDN U7514 ( .B(n56273), .A(n56272), .Z(n6907) );
  NANDN U7515 ( .A(n6906), .B(n56270), .Z(n6908) );
  AND U7516 ( .A(n6907), .B(n6908), .Z(n6909) );
  OR U7517 ( .A(n56274), .B(n6909), .Z(n6910) );
  NAND U7518 ( .A(n56275), .B(n6910), .Z(n6911) );
  NANDN U7519 ( .A(n51732), .B(n6911), .Z(n6912) );
  AND U7520 ( .A(n56276), .B(n51731), .Z(n6913) );
  NAND U7521 ( .A(n6912), .B(n6913), .Z(n6914) );
  NANDN U7522 ( .A(n56277), .B(n6914), .Z(n6915) );
  AND U7523 ( .A(n56278), .B(n56279), .Z(n6916) );
  NAND U7524 ( .A(n6915), .B(n6916), .Z(n6917) );
  NANDN U7525 ( .A(n56280), .B(n6917), .Z(n6918) );
  NAND U7526 ( .A(n56281), .B(n6918), .Z(n56282) );
  NANDN U7527 ( .A(n26596), .B(n9939), .Z(n6919) );
  AND U7528 ( .A(n26594), .B(n6919), .Z(n55160) );
  NAND U7529 ( .A(n56302), .B(n56303), .Z(n6920) );
  NAND U7530 ( .A(n56305), .B(n6920), .Z(n6921) );
  NAND U7531 ( .A(n51721), .B(n6921), .Z(n6922) );
  NANDN U7532 ( .A(n56306), .B(n6922), .Z(n6923) );
  NAND U7533 ( .A(n56307), .B(n6923), .Z(n6924) );
  ANDN U7534 ( .B(n6924), .A(n51720), .Z(n6925) );
  NANDN U7535 ( .A(n6925), .B(n51719), .Z(n6926) );
  NAND U7536 ( .A(n56308), .B(n6926), .Z(n6927) );
  NANDN U7537 ( .A(n56309), .B(n6927), .Z(n6928) );
  NAND U7538 ( .A(n56310), .B(n6928), .Z(n6929) );
  NANDN U7539 ( .A(n56311), .B(n6929), .Z(n6930) );
  AND U7540 ( .A(n56312), .B(n6930), .Z(n6931) );
  OR U7541 ( .A(n6931), .B(n56313), .Z(n6932) );
  NAND U7542 ( .A(n56314), .B(n6932), .Z(n6933) );
  NANDN U7543 ( .A(n56315), .B(n6933), .Z(n56316) );
  NANDN U7544 ( .A(n56335), .B(n56334), .Z(n6934) );
  NANDN U7545 ( .A(n56336), .B(n6934), .Z(n6935) );
  AND U7546 ( .A(n56337), .B(n6935), .Z(n6936) );
  OR U7547 ( .A(n56338), .B(n6936), .Z(n6937) );
  NAND U7548 ( .A(n56339), .B(n6937), .Z(n6938) );
  NANDN U7549 ( .A(n51707), .B(n6938), .Z(n6939) );
  NAND U7550 ( .A(n51706), .B(n6939), .Z(n6940) );
  NANDN U7551 ( .A(n56340), .B(n6940), .Z(n6941) );
  AND U7552 ( .A(n56341), .B(n6941), .Z(n6942) );
  OR U7553 ( .A(n6942), .B(n56342), .Z(n6943) );
  NAND U7554 ( .A(n56343), .B(n6943), .Z(n6944) );
  NANDN U7555 ( .A(n56344), .B(n6944), .Z(n6945) );
  NAND U7556 ( .A(n56345), .B(n6945), .Z(n56346) );
  NANDN U7557 ( .A(n51700), .B(n56369), .Z(n6946) );
  NAND U7558 ( .A(n51699), .B(n6946), .Z(n6947) );
  NANDN U7559 ( .A(n56370), .B(n6947), .Z(n6948) );
  NAND U7560 ( .A(n56371), .B(n6948), .Z(n6949) );
  NANDN U7561 ( .A(n56372), .B(n6949), .Z(n6950) );
  AND U7562 ( .A(n56373), .B(n6950), .Z(n6951) );
  OR U7563 ( .A(n51698), .B(n6951), .Z(n6952) );
  NAND U7564 ( .A(n51697), .B(n6952), .Z(n6953) );
  NANDN U7565 ( .A(n56374), .B(n6953), .Z(n6954) );
  NAND U7566 ( .A(n56375), .B(n6954), .Z(n56376) );
  NAND U7567 ( .A(n56395), .B(n56396), .Z(n6955) );
  NANDN U7568 ( .A(n56397), .B(n6955), .Z(n6956) );
  AND U7569 ( .A(n56398), .B(n6956), .Z(n6957) );
  OR U7570 ( .A(n6957), .B(n56399), .Z(n6958) );
  NAND U7571 ( .A(n56400), .B(n6958), .Z(n6959) );
  ANDN U7572 ( .B(n6959), .A(n56401), .Z(n6960) );
  NANDN U7573 ( .A(n6960), .B(n51683), .Z(n6961) );
  NANDN U7574 ( .A(n56402), .B(n6961), .Z(n6962) );
  NAND U7575 ( .A(n56403), .B(n6962), .Z(n6963) );
  NAND U7576 ( .A(n56404), .B(n6963), .Z(n6964) );
  NANDN U7577 ( .A(n56405), .B(n6964), .Z(n6965) );
  AND U7578 ( .A(n56406), .B(n6965), .Z(n6966) );
  OR U7579 ( .A(n56407), .B(n6966), .Z(n6967) );
  NAND U7580 ( .A(n56408), .B(n6967), .Z(n6968) );
  NANDN U7581 ( .A(n56409), .B(n6968), .Z(n6969) );
  NAND U7582 ( .A(n56410), .B(n6969), .Z(n56411) );
  AND U7583 ( .A(n56428), .B(n56427), .Z(n56429) );
  NANDN U7584 ( .A(n56484), .B(n56483), .Z(n6970) );
  NAND U7585 ( .A(n56485), .B(n6970), .Z(n6971) );
  NANDN U7586 ( .A(n56486), .B(n6971), .Z(n6972) );
  NAND U7587 ( .A(n56487), .B(n6972), .Z(n6973) );
  NANDN U7588 ( .A(n56488), .B(n6973), .Z(n6974) );
  AND U7589 ( .A(n56489), .B(n6974), .Z(n6975) );
  OR U7590 ( .A(n6975), .B(n56490), .Z(n6976) );
  NAND U7591 ( .A(n56491), .B(n6976), .Z(n6977) );
  ANDN U7592 ( .B(n6977), .A(n56492), .Z(n6978) );
  ANDN U7593 ( .B(n51675), .A(n6978), .Z(n6979) );
  NAND U7594 ( .A(n51674), .B(n6979), .Z(n6980) );
  ANDN U7595 ( .B(n6980), .A(n56493), .Z(n6981) );
  NANDN U7596 ( .A(n6981), .B(n56494), .Z(n6982) );
  NANDN U7597 ( .A(n56495), .B(n6982), .Z(n6983) );
  NAND U7598 ( .A(n56496), .B(n6983), .Z(n6984) );
  NANDN U7599 ( .A(n51673), .B(n6984), .Z(n56497) );
  NAND U7600 ( .A(n56527), .B(n56528), .Z(n6985) );
  NAND U7601 ( .A(n56529), .B(n6985), .Z(n6986) );
  NANDN U7602 ( .A(n51667), .B(n6986), .Z(n6987) );
  NAND U7603 ( .A(n51666), .B(n6987), .Z(n6988) );
  NANDN U7604 ( .A(n51665), .B(n6988), .Z(n6989) );
  AND U7605 ( .A(n56530), .B(n6989), .Z(n6990) );
  OR U7606 ( .A(n6990), .B(n56531), .Z(n6991) );
  NAND U7607 ( .A(n56532), .B(n6991), .Z(n6992) );
  ANDN U7608 ( .B(n6992), .A(n56533), .Z(n6993) );
  NANDN U7609 ( .A(n6993), .B(n56534), .Z(n6994) );
  NAND U7610 ( .A(n51664), .B(n6994), .Z(n6995) );
  NANDN U7611 ( .A(n56535), .B(n6995), .Z(n6996) );
  NAND U7612 ( .A(n56536), .B(n6996), .Z(n56539) );
  NANDN U7613 ( .A(n56571), .B(n56570), .Z(n6997) );
  NAND U7614 ( .A(n56572), .B(n6997), .Z(n6998) );
  NANDN U7615 ( .A(n56573), .B(n6998), .Z(n6999) );
  NAND U7616 ( .A(n56574), .B(n6999), .Z(n7000) );
  NANDN U7617 ( .A(n56575), .B(n7000), .Z(n7001) );
  AND U7618 ( .A(n56576), .B(n7001), .Z(n7002) );
  OR U7619 ( .A(n7002), .B(n56577), .Z(n7003) );
  AND U7620 ( .A(n56578), .B(n7003), .Z(n7004) );
  AND U7621 ( .A(n51657), .B(n56579), .Z(n7005) );
  OR U7622 ( .A(n51658), .B(n7004), .Z(n7006) );
  AND U7623 ( .A(n7005), .B(n7006), .Z(n7007) );
  OR U7624 ( .A(n56580), .B(n7007), .Z(n7008) );
  NAND U7625 ( .A(n56581), .B(n7008), .Z(n7009) );
  NANDN U7626 ( .A(n51656), .B(n7009), .Z(n56582) );
  NAND U7627 ( .A(n56604), .B(n56603), .Z(n7010) );
  ANDN U7628 ( .B(n7010), .A(n56605), .Z(n7011) );
  NOR U7629 ( .A(n56607), .B(n7011), .Z(n7012) );
  NAND U7630 ( .A(n56608), .B(n7012), .Z(n7013) );
  NAND U7631 ( .A(n51647), .B(n7013), .Z(n7014) );
  ANDN U7632 ( .B(n56609), .A(n51646), .Z(n7015) );
  NAND U7633 ( .A(n7014), .B(n7015), .Z(n7016) );
  NAND U7634 ( .A(n56610), .B(n7016), .Z(n7017) );
  NANDN U7635 ( .A(n56611), .B(n7017), .Z(n7018) );
  NAND U7636 ( .A(n56612), .B(n7018), .Z(n7019) );
  ANDN U7637 ( .B(n7019), .A(n51645), .Z(n7020) );
  NANDN U7638 ( .A(n7020), .B(n56613), .Z(n7021) );
  NANDN U7639 ( .A(n56614), .B(n7021), .Z(n7022) );
  NAND U7640 ( .A(n56615), .B(n7022), .Z(n56616) );
  NAND U7641 ( .A(n56639), .B(n56638), .Z(n7023) );
  NANDN U7642 ( .A(n56640), .B(n7023), .Z(n7024) );
  AND U7643 ( .A(n56641), .B(n7024), .Z(n7025) );
  OR U7644 ( .A(n56642), .B(n7025), .Z(n7026) );
  AND U7645 ( .A(n56643), .B(n7026), .Z(n7027) );
  OR U7646 ( .A(n7027), .B(n56644), .Z(n7028) );
  NAND U7647 ( .A(n56645), .B(n7028), .Z(n7029) );
  NAND U7648 ( .A(n51636), .B(n7029), .Z(n7030) );
  ANDN U7649 ( .B(n56646), .A(n56647), .Z(n7031) );
  NAND U7650 ( .A(n7030), .B(n7031), .Z(n7032) );
  NAND U7651 ( .A(n56648), .B(n7032), .Z(n7033) );
  ANDN U7652 ( .B(n51635), .A(n51634), .Z(n7034) );
  NAND U7653 ( .A(n7033), .B(n7034), .Z(n7035) );
  NAND U7654 ( .A(n56649), .B(n7035), .Z(n7036) );
  NANDN U7655 ( .A(n51633), .B(n7036), .Z(n56650) );
  NAND U7656 ( .A(n56671), .B(n56672), .Z(n7037) );
  NANDN U7657 ( .A(n56673), .B(n7037), .Z(n7038) );
  AND U7658 ( .A(n56674), .B(n7038), .Z(n7039) );
  OR U7659 ( .A(n7039), .B(n56675), .Z(n7040) );
  NAND U7660 ( .A(n56676), .B(n7040), .Z(n7041) );
  ANDN U7661 ( .B(n7041), .A(n56677), .Z(n7042) );
  NANDN U7662 ( .A(n7042), .B(n51625), .Z(n7043) );
  NANDN U7663 ( .A(n56678), .B(n7043), .Z(n7044) );
  NAND U7664 ( .A(n56679), .B(n7044), .Z(n7045) );
  NAND U7665 ( .A(n56680), .B(n7045), .Z(n7046) );
  NANDN U7666 ( .A(n56681), .B(n7046), .Z(n7047) );
  AND U7667 ( .A(n56682), .B(n7047), .Z(n7048) );
  OR U7668 ( .A(n56683), .B(n7048), .Z(n7049) );
  NAND U7669 ( .A(n56684), .B(n7049), .Z(n7050) );
  NANDN U7670 ( .A(n56685), .B(n7050), .Z(n7051) );
  NAND U7671 ( .A(n56686), .B(n7051), .Z(n56687) );
  NAND U7672 ( .A(n56708), .B(n56709), .Z(n7052) );
  NAND U7673 ( .A(n56711), .B(n7052), .Z(n7053) );
  NAND U7674 ( .A(n56712), .B(n7053), .Z(n7054) );
  NANDN U7675 ( .A(n51615), .B(n7054), .Z(n7055) );
  NAND U7676 ( .A(n51614), .B(n7055), .Z(n7056) );
  AND U7677 ( .A(n56713), .B(n7056), .Z(n7057) );
  AND U7678 ( .A(n51612), .B(n51613), .Z(n7058) );
  OR U7679 ( .A(n56714), .B(n7057), .Z(n7059) );
  AND U7680 ( .A(n7058), .B(n7059), .Z(n7060) );
  OR U7681 ( .A(n7060), .B(n56715), .Z(n7061) );
  NAND U7682 ( .A(n56716), .B(n7061), .Z(n7062) );
  ANDN U7683 ( .B(n7062), .A(n56717), .Z(n7063) );
  NANDN U7684 ( .A(n7063), .B(n56718), .Z(n7064) );
  NANDN U7685 ( .A(n56719), .B(n7064), .Z(n7065) );
  NAND U7686 ( .A(n56720), .B(n7065), .Z(n7066) );
  ANDN U7687 ( .B(n7066), .A(n56721), .Z(n56725) );
  NANDN U7688 ( .A(n56753), .B(n56752), .Z(n7067) );
  ANDN U7689 ( .B(n7067), .A(n56754), .Z(n7068) );
  NOR U7690 ( .A(n56756), .B(n7068), .Z(n7069) );
  NAND U7691 ( .A(n56755), .B(n7069), .Z(n7070) );
  ANDN U7692 ( .B(n7070), .A(n56757), .Z(n7071) );
  NANDN U7693 ( .A(n7071), .B(n56758), .Z(n7072) );
  NANDN U7694 ( .A(n51606), .B(n7072), .Z(n7073) );
  NAND U7695 ( .A(n51605), .B(n7073), .Z(n7074) );
  NANDN U7696 ( .A(n56759), .B(n7074), .Z(n7075) );
  NAND U7697 ( .A(n56760), .B(n7075), .Z(n7076) );
  AND U7698 ( .A(n56761), .B(n7076), .Z(n7077) );
  OR U7699 ( .A(n7077), .B(n56762), .Z(n7078) );
  NAND U7700 ( .A(n56763), .B(n7078), .Z(n7079) );
  NANDN U7701 ( .A(n56764), .B(n7079), .Z(n56765) );
  NANDN U7702 ( .A(n56841), .B(n56840), .Z(n7080) );
  NAND U7703 ( .A(n56842), .B(n7080), .Z(n7081) );
  ANDN U7704 ( .B(n7081), .A(n56843), .Z(n7082) );
  NANDN U7705 ( .A(n7082), .B(n56844), .Z(n7083) );
  NANDN U7706 ( .A(n56845), .B(n7083), .Z(n7084) );
  NAND U7707 ( .A(n56846), .B(n7084), .Z(n7085) );
  NAND U7708 ( .A(n56847), .B(n7085), .Z(n7086) );
  NAND U7709 ( .A(n56848), .B(n7086), .Z(n7087) );
  ANDN U7710 ( .B(n7087), .A(n56849), .Z(n7088) );
  NANDN U7711 ( .A(n7088), .B(n56850), .Z(n7089) );
  NANDN U7712 ( .A(n56851), .B(n7089), .Z(n7090) );
  NAND U7713 ( .A(n56852), .B(n7090), .Z(n7091) );
  ANDN U7714 ( .B(n56854), .A(n56853), .Z(n7092) );
  NAND U7715 ( .A(n7091), .B(n7092), .Z(n7093) );
  NANDN U7716 ( .A(n56855), .B(n7093), .Z(n7094) );
  NOR U7717 ( .A(n56856), .B(n56857), .Z(n7095) );
  NAND U7718 ( .A(n7094), .B(n7095), .Z(n7096) );
  NANDN U7719 ( .A(n56858), .B(n7096), .Z(n56859) );
  NAND U7720 ( .A(n56884), .B(n56885), .Z(n7097) );
  AND U7721 ( .A(n56887), .B(n7097), .Z(n7098) );
  ANDN U7722 ( .B(n51593), .A(n7098), .Z(n7099) );
  NAND U7723 ( .A(n51592), .B(n7099), .Z(n7100) );
  ANDN U7724 ( .B(n7100), .A(n56888), .Z(n7101) );
  ANDN U7725 ( .B(n56890), .A(n7101), .Z(n7102) );
  NAND U7726 ( .A(n56889), .B(n7102), .Z(n7103) );
  ANDN U7727 ( .B(n7103), .A(n56891), .Z(n7104) );
  NANDN U7728 ( .A(n7104), .B(n56892), .Z(n7105) );
  NANDN U7729 ( .A(n51591), .B(n7105), .Z(n7106) );
  NAND U7730 ( .A(n51590), .B(n7106), .Z(n7107) );
  ANDN U7731 ( .B(n7107), .A(n56893), .Z(n56896) );
  NANDN U7732 ( .A(n56920), .B(n56921), .Z(n7108) );
  NANDN U7733 ( .A(n56923), .B(n7108), .Z(n7109) );
  NANDN U7734 ( .A(n51582), .B(n7109), .Z(n7110) );
  AND U7735 ( .A(n56925), .B(n56924), .Z(n7111) );
  NAND U7736 ( .A(n7110), .B(n7111), .Z(n7112) );
  NANDN U7737 ( .A(n56926), .B(n7112), .Z(n7113) );
  NAND U7738 ( .A(n56927), .B(n7113), .Z(n7114) );
  NANDN U7739 ( .A(n56928), .B(n7114), .Z(n7115) );
  AND U7740 ( .A(n56929), .B(n7115), .Z(n7116) );
  OR U7741 ( .A(n56930), .B(n7116), .Z(n7117) );
  AND U7742 ( .A(n56931), .B(n7117), .Z(n7118) );
  OR U7743 ( .A(n56932), .B(n7118), .Z(n7119) );
  NAND U7744 ( .A(n56933), .B(n7119), .Z(n7120) );
  NANDN U7745 ( .A(n56934), .B(n7120), .Z(n7121) );
  NOR U7746 ( .A(n56935), .B(n51581), .Z(n7122) );
  NAND U7747 ( .A(n7121), .B(n7122), .Z(n7123) );
  NANDN U7748 ( .A(n56936), .B(n7123), .Z(n56937) );
  NAND U7749 ( .A(n56971), .B(n56972), .Z(n7124) );
  NAND U7750 ( .A(n56975), .B(n7124), .Z(n7125) );
  NAND U7751 ( .A(n56976), .B(n7125), .Z(n7126) );
  NANDN U7752 ( .A(n56977), .B(n7126), .Z(n7127) );
  NAND U7753 ( .A(n56978), .B(n7127), .Z(n7128) );
  ANDN U7754 ( .B(n7128), .A(n56979), .Z(n7129) );
  NANDN U7755 ( .A(n7129), .B(n56980), .Z(n7130) );
  NANDN U7756 ( .A(n56981), .B(n7130), .Z(n7131) );
  NAND U7757 ( .A(n56982), .B(n7131), .Z(n7132) );
  NANDN U7758 ( .A(n56983), .B(n7132), .Z(n7133) );
  NAND U7759 ( .A(n56984), .B(n7133), .Z(n7134) );
  ANDN U7760 ( .B(n7134), .A(n56985), .Z(n7135) );
  ANDN U7761 ( .B(n56988), .A(n56987), .Z(n7136) );
  NANDN U7762 ( .A(n7135), .B(n56986), .Z(n7137) );
  AND U7763 ( .A(n7136), .B(n7137), .Z(n7138) );
  ANDN U7764 ( .B(n56990), .A(n56989), .Z(n7139) );
  NANDN U7765 ( .A(n7138), .B(n51574), .Z(n7140) );
  AND U7766 ( .A(n7139), .B(n7140), .Z(n56992) );
  NAND U7767 ( .A(n57030), .B(n57029), .Z(n7141) );
  NANDN U7768 ( .A(n57031), .B(n7141), .Z(n7142) );
  AND U7769 ( .A(n57032), .B(n7142), .Z(n7143) );
  AND U7770 ( .A(n57035), .B(n57034), .Z(n7144) );
  OR U7771 ( .A(n57033), .B(n7143), .Z(n7145) );
  AND U7772 ( .A(n7144), .B(n7145), .Z(n7146) );
  OR U7773 ( .A(n7146), .B(n51569), .Z(n7147) );
  NAND U7774 ( .A(n57036), .B(n7147), .Z(n7148) );
  ANDN U7775 ( .B(n7148), .A(n51568), .Z(n7149) );
  NANDN U7776 ( .A(n7149), .B(n51567), .Z(n7150) );
  ANDN U7777 ( .B(n7150), .A(n57037), .Z(n7151) );
  NANDN U7778 ( .A(n7151), .B(n57038), .Z(n7152) );
  NAND U7779 ( .A(n57039), .B(n7152), .Z(n7153) );
  NANDN U7780 ( .A(n57040), .B(n7153), .Z(n57041) );
  NAND U7781 ( .A(n57069), .B(n57068), .Z(n7154) );
  NAND U7782 ( .A(n51559), .B(n7154), .Z(n7155) );
  ANDN U7783 ( .B(n7155), .A(n57070), .Z(n7156) );
  NANDN U7784 ( .A(n7156), .B(n57071), .Z(n7157) );
  NAND U7785 ( .A(n57072), .B(n7157), .Z(n7158) );
  NANDN U7786 ( .A(n57073), .B(n7158), .Z(n7159) );
  NAND U7787 ( .A(n57074), .B(n7159), .Z(n7160) );
  NANDN U7788 ( .A(n57075), .B(n7160), .Z(n7161) );
  AND U7789 ( .A(n57076), .B(n7161), .Z(n7162) );
  OR U7790 ( .A(n7162), .B(n57077), .Z(n7163) );
  AND U7791 ( .A(n57078), .B(n7163), .Z(n7164) );
  NANDN U7792 ( .A(n7164), .B(n51558), .Z(n7165) );
  NANDN U7793 ( .A(n57079), .B(n7165), .Z(n7166) );
  NAND U7794 ( .A(n57080), .B(n7166), .Z(n57083) );
  NAND U7795 ( .A(n57110), .B(n57109), .Z(n7167) );
  AND U7796 ( .A(n57111), .B(n7167), .Z(n7168) );
  NANDN U7797 ( .A(n7168), .B(n57112), .Z(n7169) );
  NAND U7798 ( .A(n57113), .B(n7169), .Z(n7170) );
  NANDN U7799 ( .A(n57114), .B(n7170), .Z(n7171) );
  AND U7800 ( .A(n51547), .B(n51546), .Z(n7172) );
  NAND U7801 ( .A(n7171), .B(n7172), .Z(n7173) );
  NANDN U7802 ( .A(n57115), .B(n7173), .Z(n7174) );
  NAND U7803 ( .A(n57116), .B(n7174), .Z(n7175) );
  NANDN U7804 ( .A(n57117), .B(n7175), .Z(n7176) );
  AND U7805 ( .A(n57118), .B(n7176), .Z(n7177) );
  OR U7806 ( .A(n57119), .B(n7177), .Z(n7178) );
  NAND U7807 ( .A(n57120), .B(n7178), .Z(n7179) );
  NANDN U7808 ( .A(n57121), .B(n7179), .Z(n7180) );
  AND U7809 ( .A(n57122), .B(n57123), .Z(n7181) );
  NAND U7810 ( .A(n7180), .B(n7181), .Z(n7182) );
  NANDN U7811 ( .A(n57124), .B(n7182), .Z(n57125) );
  NAND U7812 ( .A(n57156), .B(n57157), .Z(n7183) );
  AND U7813 ( .A(n51541), .B(n51540), .Z(n7184) );
  NANDN U7814 ( .A(n57158), .B(n7183), .Z(n7185) );
  NAND U7815 ( .A(n7184), .B(n7185), .Z(n7186) );
  AND U7816 ( .A(n57160), .B(n57161), .Z(n7187) );
  NANDN U7817 ( .A(n57159), .B(n7186), .Z(n7188) );
  NAND U7818 ( .A(n7187), .B(n7188), .Z(n7189) );
  NAND U7819 ( .A(n51539), .B(n7189), .Z(n7190) );
  AND U7820 ( .A(n57162), .B(n7190), .Z(n7191) );
  NANDN U7821 ( .A(n57163), .B(n7191), .Z(n7192) );
  NAND U7822 ( .A(n57164), .B(n7192), .Z(n7193) );
  AND U7823 ( .A(n57166), .B(n7193), .Z(n7194) );
  NAND U7824 ( .A(n7194), .B(n57165), .Z(n7195) );
  AND U7825 ( .A(n51538), .B(n51537), .Z(n7196) );
  NANDN U7826 ( .A(n57167), .B(n7195), .Z(n7197) );
  NAND U7827 ( .A(n7196), .B(n7197), .Z(n57170) );
  NAND U7828 ( .A(n57203), .B(n57204), .Z(n7198) );
  NANDN U7829 ( .A(n57205), .B(n7198), .Z(n7199) );
  NAND U7830 ( .A(n57206), .B(n7199), .Z(n7200) );
  NANDN U7831 ( .A(n57207), .B(n7200), .Z(n7201) );
  NAND U7832 ( .A(n57208), .B(n7201), .Z(n7202) );
  ANDN U7833 ( .B(n7202), .A(n57209), .Z(n7203) );
  AND U7834 ( .A(n51533), .B(n51534), .Z(n7204) );
  NANDN U7835 ( .A(n7203), .B(n57210), .Z(n7205) );
  AND U7836 ( .A(n7204), .B(n7205), .Z(n7206) );
  NANDN U7837 ( .A(n7206), .B(n57211), .Z(n7207) );
  ANDN U7838 ( .B(n7207), .A(n51532), .Z(n7208) );
  NANDN U7839 ( .A(n7208), .B(n51531), .Z(n7209) );
  NANDN U7840 ( .A(n57212), .B(n7209), .Z(n7210) );
  NAND U7841 ( .A(n57213), .B(n7210), .Z(n57214) );
  AND U7842 ( .A(n57238), .B(n57237), .Z(n7211) );
  AND U7843 ( .A(n57240), .B(n57241), .Z(n7212) );
  OR U7844 ( .A(n57239), .B(n7211), .Z(n7213) );
  AND U7845 ( .A(n7212), .B(n7213), .Z(n7214) );
  AND U7846 ( .A(n51523), .B(n57243), .Z(n7215) );
  OR U7847 ( .A(n57242), .B(n7214), .Z(n7216) );
  AND U7848 ( .A(n7215), .B(n7216), .Z(n7217) );
  NANDN U7849 ( .A(n7217), .B(n57244), .Z(n7218) );
  NANDN U7850 ( .A(n57245), .B(n7218), .Z(n7219) );
  NAND U7851 ( .A(n57246), .B(n7219), .Z(n7220) );
  AND U7852 ( .A(n57247), .B(n57248), .Z(n7221) );
  NAND U7853 ( .A(n7220), .B(n7221), .Z(n7222) );
  NANDN U7854 ( .A(n57249), .B(n7222), .Z(n7223) );
  AND U7855 ( .A(n57250), .B(n57251), .Z(n7224) );
  NAND U7856 ( .A(n7223), .B(n7224), .Z(n7225) );
  NANDN U7857 ( .A(n57252), .B(n7225), .Z(n57253) );
  ANDN U7858 ( .B(n57315), .A(n57316), .Z(n7226) );
  NAND U7859 ( .A(n57314), .B(n7226), .Z(n7227) );
  NAND U7860 ( .A(n57317), .B(n7227), .Z(n7228) );
  AND U7861 ( .A(n57321), .B(n57320), .Z(n7229) );
  NANDN U7862 ( .A(n57318), .B(n7228), .Z(n7230) );
  NAND U7863 ( .A(n57319), .B(n7230), .Z(n7231) );
  AND U7864 ( .A(n7229), .B(n7231), .Z(n7232) );
  AND U7865 ( .A(n57324), .B(n57323), .Z(n7233) );
  OR U7866 ( .A(n57322), .B(n7232), .Z(n7234) );
  AND U7867 ( .A(n7233), .B(n7234), .Z(n7235) );
  NANDN U7868 ( .A(n7235), .B(n57325), .Z(n7236) );
  NAND U7869 ( .A(n57326), .B(n7236), .Z(n7237) );
  NAND U7870 ( .A(n57327), .B(n7237), .Z(n7238) );
  AND U7871 ( .A(n57328), .B(n57329), .Z(n7239) );
  NAND U7872 ( .A(n7238), .B(n7239), .Z(n7240) );
  NAND U7873 ( .A(n51509), .B(n7240), .Z(n7241) );
  AND U7874 ( .A(n57330), .B(n7241), .Z(n57331) );
  NANDN U7875 ( .A(n57363), .B(n57362), .Z(n7242) );
  NANDN U7876 ( .A(n57364), .B(n7242), .Z(n7243) );
  ANDN U7877 ( .B(n7243), .A(n57365), .Z(n7244) );
  NAND U7878 ( .A(n7244), .B(n57366), .Z(n7245) );
  NANDN U7879 ( .A(n57367), .B(n7245), .Z(n7246) );
  AND U7880 ( .A(n57368), .B(n7246), .Z(n7247) );
  OR U7881 ( .A(n57369), .B(n7247), .Z(n7248) );
  NAND U7882 ( .A(n57370), .B(n7248), .Z(n7249) );
  NANDN U7883 ( .A(n57371), .B(n7249), .Z(n7250) );
  AND U7884 ( .A(n57372), .B(n7250), .Z(n7251) );
  AND U7885 ( .A(n51502), .B(n51501), .Z(n7252) );
  OR U7886 ( .A(n57373), .B(n7251), .Z(n7253) );
  AND U7887 ( .A(n7252), .B(n7253), .Z(n7254) );
  OR U7888 ( .A(n57374), .B(n7254), .Z(n7255) );
  NAND U7889 ( .A(n57375), .B(n7255), .Z(n7256) );
  NANDN U7890 ( .A(n57376), .B(n7256), .Z(n7257) );
  ANDN U7891 ( .B(n57377), .A(n57378), .Z(n7258) );
  NAND U7892 ( .A(n7257), .B(n7258), .Z(n7259) );
  NANDN U7893 ( .A(n51500), .B(n7259), .Z(n57379) );
  ANDN U7894 ( .B(n57409), .A(n57410), .Z(n7260) );
  OR U7895 ( .A(n57407), .B(n57408), .Z(n7261) );
  AND U7896 ( .A(n7260), .B(n7261), .Z(n7262) );
  OR U7897 ( .A(n57411), .B(n7262), .Z(n7263) );
  AND U7898 ( .A(n57412), .B(n7263), .Z(n7264) );
  AND U7899 ( .A(n57415), .B(n57414), .Z(n7265) );
  OR U7900 ( .A(n57413), .B(n7264), .Z(n7266) );
  AND U7901 ( .A(n7265), .B(n7266), .Z(n7267) );
  OR U7902 ( .A(n57416), .B(n7267), .Z(n7268) );
  NAND U7903 ( .A(n57417), .B(n7268), .Z(n7269) );
  NANDN U7904 ( .A(n57418), .B(n7269), .Z(n7270) );
  ANDN U7905 ( .B(n51494), .A(n51493), .Z(n7271) );
  NAND U7906 ( .A(n7270), .B(n7271), .Z(n7272) );
  NANDN U7907 ( .A(n57419), .B(n7272), .Z(n7273) );
  NAND U7908 ( .A(n57420), .B(n7273), .Z(n57421) );
  AND U7909 ( .A(n51482), .B(n51483), .Z(n7274) );
  AND U7910 ( .A(n57453), .B(n57455), .Z(n7275) );
  NAND U7911 ( .A(n57454), .B(n7275), .Z(n7276) );
  NANDN U7912 ( .A(n57456), .B(n7276), .Z(n7277) );
  AND U7913 ( .A(n51487), .B(n51486), .Z(n7278) );
  NAND U7914 ( .A(n7277), .B(n7278), .Z(n7279) );
  NANDN U7915 ( .A(n57457), .B(n7279), .Z(n7280) );
  AND U7916 ( .A(n51485), .B(n51484), .Z(n7281) );
  NAND U7917 ( .A(n7280), .B(n7281), .Z(n7282) );
  NAND U7918 ( .A(n57458), .B(n7282), .Z(n7283) );
  ANDN U7919 ( .B(n57459), .A(n57460), .Z(n7284) );
  NAND U7920 ( .A(n7283), .B(n7284), .Z(n7285) );
  NANDN U7921 ( .A(n57461), .B(n7285), .Z(n7286) );
  ANDN U7922 ( .B(n57463), .A(n57462), .Z(n7287) );
  NAND U7923 ( .A(n7286), .B(n7287), .Z(n7288) );
  NANDN U7924 ( .A(n57464), .B(n7288), .Z(n7289) );
  NAND U7925 ( .A(n7274), .B(n7289), .Z(n57465) );
  NOR U7926 ( .A(n16258), .B(n25144), .Z(n7290) );
  XNOR U7927 ( .A(y[4412]), .B(x[4412]), .Z(n7291) );
  NAND U7928 ( .A(n7290), .B(n7291), .Z(n7292) );
  NAND U7929 ( .A(n56654), .B(n7292), .Z(n7293) );
  AND U7930 ( .A(n41295), .B(n7293), .Z(n7294) );
  NAND U7931 ( .A(n7294), .B(n56655), .Z(n7295) );
  NAND U7932 ( .A(n56657), .B(n7295), .Z(n7296) );
  NANDN U7933 ( .A(n51631), .B(n7296), .Z(n7297) );
  AND U7934 ( .A(n51630), .B(n7297), .Z(n7298) );
  OR U7935 ( .A(n56658), .B(n7298), .Z(n7299) );
  NAND U7936 ( .A(n56659), .B(n7299), .Z(n7300) );
  NANDN U7937 ( .A(n56660), .B(n7300), .Z(n7301) );
  NAND U7938 ( .A(n56661), .B(n7301), .Z(n7302) );
  NANDN U7939 ( .A(n51629), .B(n7302), .Z(n7303) );
  AND U7940 ( .A(n51628), .B(n7303), .Z(n7304) );
  OR U7941 ( .A(n56663), .B(n7304), .Z(n7305) );
  NAND U7942 ( .A(n56664), .B(n7305), .Z(n7306) );
  NANDN U7943 ( .A(n51627), .B(n7306), .Z(n7307) );
  NAND U7944 ( .A(n51626), .B(n7307), .Z(n16261) );
  NANDN U7945 ( .A(n57496), .B(n57495), .Z(n7308) );
  NANDN U7946 ( .A(n57497), .B(n7308), .Z(n7309) );
  AND U7947 ( .A(n57498), .B(n7309), .Z(n7310) );
  AND U7948 ( .A(n57500), .B(n57501), .Z(n7311) );
  OR U7949 ( .A(n57499), .B(n7310), .Z(n7312) );
  AND U7950 ( .A(n7311), .B(n7312), .Z(n7313) );
  AND U7951 ( .A(n51474), .B(n51473), .Z(n7314) );
  OR U7952 ( .A(n57502), .B(n7313), .Z(n7315) );
  AND U7953 ( .A(n7314), .B(n7315), .Z(n7316) );
  NANDN U7954 ( .A(n7316), .B(n57503), .Z(n7317) );
  NANDN U7955 ( .A(n51472), .B(n7317), .Z(n7318) );
  NAND U7956 ( .A(n57504), .B(n7318), .Z(n7319) );
  AND U7957 ( .A(n57506), .B(n57505), .Z(n7320) );
  NAND U7958 ( .A(n7319), .B(n7320), .Z(n7321) );
  NANDN U7959 ( .A(n51471), .B(n7321), .Z(n57507) );
  NANDN U7960 ( .A(n57542), .B(n57541), .Z(n7322) );
  NAND U7961 ( .A(n51465), .B(n7322), .Z(n7323) );
  ANDN U7962 ( .B(n7323), .A(n57543), .Z(n7324) );
  NANDN U7963 ( .A(n57544), .B(n7324), .Z(n7325) );
  NANDN U7964 ( .A(n57545), .B(n7325), .Z(n7326) );
  AND U7965 ( .A(n57546), .B(n7326), .Z(n7327) );
  NAND U7966 ( .A(n57547), .B(n7327), .Z(n7328) );
  NAND U7967 ( .A(n57548), .B(n7328), .Z(n7329) );
  NANDN U7968 ( .A(n57549), .B(n7329), .Z(n7330) );
  NAND U7969 ( .A(n57550), .B(n7330), .Z(n7331) );
  AND U7970 ( .A(n51464), .B(n7331), .Z(n7332) );
  NAND U7971 ( .A(n7332), .B(n51463), .Z(n7333) );
  NANDN U7972 ( .A(n51462), .B(n7333), .Z(n57551) );
  AND U7973 ( .A(n57574), .B(n57575), .Z(n7334) );
  NAND U7974 ( .A(n57573), .B(n7334), .Z(n7335) );
  NANDN U7975 ( .A(n57576), .B(n7335), .Z(n7336) );
  ANDN U7976 ( .B(n51450), .A(n51451), .Z(n7337) );
  NAND U7977 ( .A(n7336), .B(n7337), .Z(n7338) );
  NANDN U7978 ( .A(n57577), .B(n7338), .Z(n7339) );
  AND U7979 ( .A(n57578), .B(n57579), .Z(n7340) );
  NAND U7980 ( .A(n7339), .B(n7340), .Z(n7341) );
  NANDN U7981 ( .A(n57580), .B(n7341), .Z(n7342) );
  AND U7982 ( .A(n51449), .B(n57581), .Z(n7343) );
  NAND U7983 ( .A(n7342), .B(n7343), .Z(n7344) );
  NANDN U7984 ( .A(n51448), .B(n7344), .Z(n7345) );
  NAND U7985 ( .A(n51447), .B(n7345), .Z(n57584) );
  XNOR U7986 ( .A(x[4586]), .B(y[4586]), .Z(n16467) );
  AND U7987 ( .A(n51442), .B(n51441), .Z(n57595) );
  ANDN U7988 ( .B(n57630), .A(n57631), .Z(n7346) );
  NAND U7989 ( .A(n57629), .B(n7346), .Z(n7347) );
  NAND U7990 ( .A(n57632), .B(n7347), .Z(n7348) );
  NANDN U7991 ( .A(n57633), .B(n7348), .Z(n7349) );
  NAND U7992 ( .A(n57634), .B(n7349), .Z(n7350) );
  AND U7993 ( .A(n57635), .B(n7350), .Z(n7351) );
  NAND U7994 ( .A(n57636), .B(n7351), .Z(n7352) );
  NANDN U7995 ( .A(n57637), .B(n7352), .Z(n7353) );
  NANDN U7996 ( .A(n57638), .B(n7353), .Z(n7354) );
  NANDN U7997 ( .A(n7354), .B(n57639), .Z(n7355) );
  AND U7998 ( .A(n57640), .B(n7355), .Z(n7356) );
  ANDN U7999 ( .B(n51438), .A(n7356), .Z(n7357) );
  NAND U8000 ( .A(n51437), .B(n7357), .Z(n7358) );
  AND U8001 ( .A(n57641), .B(n7358), .Z(n57645) );
  NANDN U8002 ( .A(n57668), .B(n57667), .Z(n7359) );
  NAND U8003 ( .A(n57670), .B(n7359), .Z(n7360) );
  AND U8004 ( .A(n57671), .B(n7360), .Z(n7361) );
  AND U8005 ( .A(n57674), .B(n57673), .Z(n7362) );
  OR U8006 ( .A(n7361), .B(n57672), .Z(n7363) );
  AND U8007 ( .A(n7362), .B(n7363), .Z(n7364) );
  OR U8008 ( .A(n57675), .B(n7364), .Z(n7365) );
  NAND U8009 ( .A(n57676), .B(n7365), .Z(n7366) );
  NANDN U8010 ( .A(n57677), .B(n7366), .Z(n7367) );
  NAND U8011 ( .A(n57678), .B(n7367), .Z(n7368) );
  NANDN U8012 ( .A(n57679), .B(n7368), .Z(n7369) );
  AND U8013 ( .A(n57680), .B(n7369), .Z(n7370) );
  AND U8014 ( .A(n51427), .B(n51428), .Z(n7371) );
  OR U8015 ( .A(n7370), .B(n57681), .Z(n7372) );
  AND U8016 ( .A(n7371), .B(n7372), .Z(n7373) );
  NANDN U8017 ( .A(n7373), .B(n57682), .Z(n7374) );
  NANDN U8018 ( .A(n57683), .B(n7374), .Z(n7375) );
  NAND U8019 ( .A(n51426), .B(n7375), .Z(n57685) );
  NAND U8020 ( .A(n57711), .B(n57710), .Z(n7376) );
  NANDN U8021 ( .A(n57712), .B(n7376), .Z(n7377) );
  ANDN U8022 ( .B(n7377), .A(n57713), .Z(n7378) );
  NANDN U8023 ( .A(n57714), .B(n7378), .Z(n7379) );
  NAND U8024 ( .A(n57715), .B(n7379), .Z(n7380) );
  AND U8025 ( .A(n57716), .B(n7380), .Z(n7381) );
  AND U8026 ( .A(n57719), .B(n57718), .Z(n7382) );
  NANDN U8027 ( .A(n7381), .B(n57717), .Z(n7383) );
  AND U8028 ( .A(n7382), .B(n7383), .Z(n7384) );
  NANDN U8029 ( .A(n7384), .B(n51414), .Z(n7385) );
  AND U8030 ( .A(n57720), .B(n7385), .Z(n7386) );
  NAND U8031 ( .A(n7386), .B(n51413), .Z(n7387) );
  NAND U8032 ( .A(n57721), .B(n7387), .Z(n7388) );
  NAND U8033 ( .A(n51412), .B(n7388), .Z(n57724) );
  NAND U8034 ( .A(n57746), .B(n57745), .Z(n7389) );
  AND U8035 ( .A(n57748), .B(n7389), .Z(n7390) );
  NOR U8036 ( .A(n7390), .B(n51402), .Z(n7391) );
  NAND U8037 ( .A(n51403), .B(n7391), .Z(n7392) );
  NANDN U8038 ( .A(n57749), .B(n7392), .Z(n7393) );
  ANDN U8039 ( .B(n57750), .A(n57751), .Z(n7394) );
  NAND U8040 ( .A(n7393), .B(n7394), .Z(n7395) );
  NANDN U8041 ( .A(n57752), .B(n7395), .Z(n7396) );
  NAND U8042 ( .A(n57753), .B(n7396), .Z(n7397) );
  NANDN U8043 ( .A(n51401), .B(n7397), .Z(n7398) );
  AND U8044 ( .A(n51400), .B(n7398), .Z(n7399) );
  OR U8045 ( .A(n57754), .B(n7399), .Z(n7400) );
  NAND U8046 ( .A(n57755), .B(n7400), .Z(n7401) );
  NANDN U8047 ( .A(n57756), .B(n7401), .Z(n57757) );
  AND U8048 ( .A(n51392), .B(n57786), .Z(n7402) );
  NAND U8049 ( .A(n51393), .B(n7402), .Z(n7403) );
  AND U8050 ( .A(n57787), .B(n7403), .Z(n7404) );
  ANDN U8051 ( .B(n57788), .A(n7404), .Z(n7405) );
  NAND U8052 ( .A(n57789), .B(n7405), .Z(n7406) );
  ANDN U8053 ( .B(n7406), .A(n57790), .Z(n7407) );
  ANDN U8054 ( .B(n57792), .A(n7407), .Z(n7408) );
  NAND U8055 ( .A(n57791), .B(n7408), .Z(n7409) );
  ANDN U8056 ( .B(n7409), .A(n57793), .Z(n7410) );
  ANDN U8057 ( .B(n57795), .A(n7410), .Z(n7411) );
  NAND U8058 ( .A(n57794), .B(n7411), .Z(n7412) );
  ANDN U8059 ( .B(n7412), .A(n57796), .Z(n7413) );
  NANDN U8060 ( .A(n7413), .B(n57797), .Z(n7414) );
  ANDN U8061 ( .B(n7414), .A(n57798), .Z(n7415) );
  NOR U8062 ( .A(n57800), .B(n7415), .Z(n7416) );
  NAND U8063 ( .A(n57799), .B(n7416), .Z(n7417) );
  NANDN U8064 ( .A(n57801), .B(n7417), .Z(n57803) );
  NAND U8065 ( .A(n57831), .B(n57830), .Z(n7418) );
  NAND U8066 ( .A(n57832), .B(n7418), .Z(n7419) );
  AND U8067 ( .A(n57833), .B(n7419), .Z(n7420) );
  NAND U8068 ( .A(n7420), .B(n57834), .Z(n7421) );
  NANDN U8069 ( .A(n57835), .B(n7421), .Z(n7422) );
  AND U8070 ( .A(n57836), .B(n7422), .Z(n7423) );
  NAND U8071 ( .A(n7423), .B(n57837), .Z(n7424) );
  NANDN U8072 ( .A(n57838), .B(n7424), .Z(n7425) );
  AND U8073 ( .A(n57839), .B(n7425), .Z(n7426) );
  ANDN U8074 ( .B(n7426), .A(n57840), .Z(n7427) );
  ANDN U8075 ( .B(n51382), .A(n51381), .Z(n7428) );
  OR U8076 ( .A(n57841), .B(n7427), .Z(n7429) );
  AND U8077 ( .A(n7428), .B(n7429), .Z(n7430) );
  ANDN U8078 ( .B(n57844), .A(n57843), .Z(n7431) );
  NANDN U8079 ( .A(n7430), .B(n57842), .Z(n7432) );
  AND U8080 ( .A(n7431), .B(n7432), .Z(n7433) );
  ANDN U8081 ( .B(n57847), .A(n57846), .Z(n7434) );
  OR U8082 ( .A(n7433), .B(n57845), .Z(n7435) );
  AND U8083 ( .A(n7434), .B(n7435), .Z(n57849) );
  AND U8084 ( .A(n57866), .B(n57865), .Z(n57867) );
  NANDN U8085 ( .A(n57893), .B(n57892), .Z(n7436) );
  ANDN U8086 ( .B(n7436), .A(n57894), .Z(n7437) );
  NOR U8087 ( .A(n57896), .B(n7437), .Z(n7438) );
  NAND U8088 ( .A(n57895), .B(n7438), .Z(n7439) );
  NANDN U8089 ( .A(n57897), .B(n7439), .Z(n7440) );
  NAND U8090 ( .A(n57898), .B(n7440), .Z(n7441) );
  NANDN U8091 ( .A(n51367), .B(n7441), .Z(n7442) );
  AND U8092 ( .A(n51366), .B(n7442), .Z(n7443) );
  OR U8093 ( .A(n57899), .B(n7443), .Z(n7444) );
  NAND U8094 ( .A(n57900), .B(n7444), .Z(n7445) );
  NANDN U8095 ( .A(n57901), .B(n7445), .Z(n7446) );
  AND U8096 ( .A(n57903), .B(n57902), .Z(n7447) );
  NAND U8097 ( .A(n7446), .B(n7447), .Z(n7448) );
  NANDN U8098 ( .A(n57904), .B(n7448), .Z(n57905) );
  ANDN U8099 ( .B(n24655), .A(n57261), .Z(n7449) );
  NANDN U8100 ( .A(n57260), .B(n16961), .Z(n7450) );
  AND U8101 ( .A(n7449), .B(n7450), .Z(n7451) );
  NANDN U8102 ( .A(n7451), .B(n57262), .Z(n7452) );
  NANDN U8103 ( .A(n57263), .B(n7452), .Z(n7453) );
  NAND U8104 ( .A(n57264), .B(n7453), .Z(n7454) );
  AND U8105 ( .A(n57266), .B(n7454), .Z(n7455) );
  XNOR U8106 ( .A(y[4954]), .B(x[4954]), .Z(n7456) );
  AND U8107 ( .A(n7455), .B(n7456), .Z(n7457) );
  ANDN U8108 ( .B(n42783), .A(n42779), .Z(n7458) );
  NANDN U8109 ( .A(n7457), .B(n51519), .Z(n7459) );
  AND U8110 ( .A(n7458), .B(n7459), .Z(n7460) );
  ANDN U8111 ( .B(n24647), .A(n57272), .Z(n7461) );
  OR U8112 ( .A(n57271), .B(n7460), .Z(n7462) );
  AND U8113 ( .A(n7461), .B(n7462), .Z(n7463) );
  AND U8114 ( .A(n24645), .B(n51517), .Z(n7464) );
  OR U8115 ( .A(n7463), .B(n57274), .Z(n7465) );
  NAND U8116 ( .A(n7464), .B(n7465), .Z(n7466) );
  NAND U8117 ( .A(n57275), .B(n7466), .Z(n16964) );
  ANDN U8118 ( .B(n57930), .A(n57932), .Z(n7467) );
  NAND U8119 ( .A(n57931), .B(n7467), .Z(n7468) );
  ANDN U8120 ( .B(n7468), .A(n57933), .Z(n7469) );
  NANDN U8121 ( .A(n7469), .B(n57934), .Z(n7470) );
  ANDN U8122 ( .B(n7470), .A(n57935), .Z(n7471) );
  ANDN U8123 ( .B(n51360), .A(n7471), .Z(n7472) );
  NAND U8124 ( .A(n51359), .B(n7472), .Z(n7473) );
  AND U8125 ( .A(n57936), .B(n7473), .Z(n7474) );
  ANDN U8126 ( .B(n51358), .A(n7474), .Z(n7475) );
  NAND U8127 ( .A(n57937), .B(n7475), .Z(n7476) );
  ANDN U8128 ( .B(n7476), .A(n51357), .Z(n7477) );
  NANDN U8129 ( .A(n7477), .B(n51356), .Z(n7478) );
  NANDN U8130 ( .A(n57938), .B(n7478), .Z(n7479) );
  NAND U8131 ( .A(n57939), .B(n7479), .Z(n57940) );
  ANDN U8132 ( .B(n57973), .A(n57972), .Z(n7480) );
  NANDN U8133 ( .A(n57971), .B(n57970), .Z(n7481) );
  AND U8134 ( .A(n7480), .B(n7481), .Z(n7482) );
  NANDN U8135 ( .A(n7482), .B(n57974), .Z(n7483) );
  NANDN U8136 ( .A(n57975), .B(n7483), .Z(n7484) );
  NAND U8137 ( .A(n57976), .B(n7484), .Z(n7485) );
  AND U8138 ( .A(n51349), .B(n51350), .Z(n7486) );
  NAND U8139 ( .A(n7485), .B(n7486), .Z(n7487) );
  NANDN U8140 ( .A(n51348), .B(n7487), .Z(n7488) );
  ANDN U8141 ( .B(n57977), .A(n57978), .Z(n7489) );
  NAND U8142 ( .A(n7488), .B(n7489), .Z(n7490) );
  NAND U8143 ( .A(n57979), .B(n7490), .Z(n7491) );
  ANDN U8144 ( .B(n7491), .A(n57980), .Z(n57982) );
  OR U8145 ( .A(n58015), .B(n58014), .Z(n7492) );
  NAND U8146 ( .A(n58016), .B(n7492), .Z(n7493) );
  ANDN U8147 ( .B(n7493), .A(n58017), .Z(n7494) );
  AND U8148 ( .A(n58019), .B(n58020), .Z(n7495) );
  NANDN U8149 ( .A(n7494), .B(n58018), .Z(n7496) );
  AND U8150 ( .A(n7495), .B(n7496), .Z(n7497) );
  OR U8151 ( .A(n58021), .B(n7497), .Z(n7498) );
  AND U8152 ( .A(n58022), .B(n7498), .Z(n7499) );
  AND U8153 ( .A(n51343), .B(n51342), .Z(n7500) );
  NANDN U8154 ( .A(n7499), .B(n58023), .Z(n7501) );
  AND U8155 ( .A(n7500), .B(n7501), .Z(n7502) );
  AND U8156 ( .A(n58026), .B(n58025), .Z(n7503) );
  NANDN U8157 ( .A(n7502), .B(n58024), .Z(n7504) );
  AND U8158 ( .A(n7503), .B(n7504), .Z(n7505) );
  OR U8159 ( .A(n58027), .B(n7505), .Z(n7506) );
  NAND U8160 ( .A(n58028), .B(n7506), .Z(n7507) );
  NAND U8161 ( .A(n58029), .B(n7507), .Z(n58030) );
  NANDN U8162 ( .A(n58059), .B(n58058), .Z(n7508) );
  ANDN U8163 ( .B(n7508), .A(n58060), .Z(n7509) );
  AND U8164 ( .A(n51331), .B(n51330), .Z(n7510) );
  NANDN U8165 ( .A(n7509), .B(n58061), .Z(n7511) );
  AND U8166 ( .A(n7510), .B(n7511), .Z(n7512) );
  OR U8167 ( .A(n58062), .B(n7512), .Z(n7513) );
  NAND U8168 ( .A(n58063), .B(n7513), .Z(n7514) );
  NANDN U8169 ( .A(n58064), .B(n7514), .Z(n7515) );
  AND U8170 ( .A(n58065), .B(n58066), .Z(n7516) );
  NAND U8171 ( .A(n7515), .B(n7516), .Z(n7517) );
  NANDN U8172 ( .A(n58067), .B(n7517), .Z(n7518) );
  AND U8173 ( .A(n51329), .B(n51328), .Z(n7519) );
  NAND U8174 ( .A(n7518), .B(n7519), .Z(n7520) );
  NAND U8175 ( .A(n58068), .B(n7520), .Z(n7521) );
  AND U8176 ( .A(n58070), .B(n58069), .Z(n7522) );
  NAND U8177 ( .A(n7521), .B(n7522), .Z(n7523) );
  NANDN U8178 ( .A(n58071), .B(n7523), .Z(n58072) );
  XNOR U8179 ( .A(x[5146]), .B(y[5146]), .Z(n17231) );
  AND U8180 ( .A(n51320), .B(n51321), .Z(n7524) );
  NANDN U8181 ( .A(n58109), .B(n58108), .Z(n7525) );
  NAND U8182 ( .A(n7524), .B(n7525), .Z(n7526) );
  AND U8183 ( .A(n58112), .B(n58111), .Z(n7527) );
  NANDN U8184 ( .A(n58110), .B(n7526), .Z(n7528) );
  NAND U8185 ( .A(n7527), .B(n7528), .Z(n7529) );
  NAND U8186 ( .A(n51319), .B(n7529), .Z(n7530) );
  AND U8187 ( .A(n58113), .B(n7530), .Z(n7531) );
  NAND U8188 ( .A(n7531), .B(n58114), .Z(n7532) );
  AND U8189 ( .A(n58116), .B(n58117), .Z(n7533) );
  NANDN U8190 ( .A(n58115), .B(n7532), .Z(n7534) );
  NAND U8191 ( .A(n7533), .B(n7534), .Z(n7535) );
  AND U8192 ( .A(n51318), .B(n51317), .Z(n7536) );
  NANDN U8193 ( .A(n58118), .B(n7535), .Z(n7537) );
  NAND U8194 ( .A(n7536), .B(n7537), .Z(n7538) );
  NANDN U8195 ( .A(n58119), .B(n7538), .Z(n58120) );
  AND U8196 ( .A(n58148), .B(n58149), .Z(n7539) );
  NAND U8197 ( .A(n58147), .B(n7539), .Z(n7540) );
  AND U8198 ( .A(n58150), .B(n7540), .Z(n7541) );
  ANDN U8199 ( .B(n58152), .A(n7541), .Z(n7542) );
  NAND U8200 ( .A(n58151), .B(n7542), .Z(n7543) );
  ANDN U8201 ( .B(n7543), .A(n58153), .Z(n7544) );
  NANDN U8202 ( .A(n7544), .B(n58154), .Z(n7545) );
  ANDN U8203 ( .B(n7545), .A(n58155), .Z(n7546) );
  ANDN U8204 ( .B(n51308), .A(n7546), .Z(n7547) );
  NAND U8205 ( .A(n51307), .B(n7547), .Z(n7548) );
  NAND U8206 ( .A(n51306), .B(n7548), .Z(n7549) );
  AND U8207 ( .A(n58156), .B(n58157), .Z(n7550) );
  NAND U8208 ( .A(n7549), .B(n7550), .Z(n7551) );
  NAND U8209 ( .A(n58158), .B(n7551), .Z(n7552) );
  AND U8210 ( .A(n51304), .B(n51305), .Z(n7553) );
  NAND U8211 ( .A(n7552), .B(n7553), .Z(n7554) );
  NANDN U8212 ( .A(n58159), .B(n7554), .Z(n58160) );
  AND U8213 ( .A(n58188), .B(n51296), .Z(n7555) );
  NAND U8214 ( .A(n51295), .B(n7555), .Z(n7556) );
  NANDN U8215 ( .A(n58189), .B(n7556), .Z(n7557) );
  AND U8216 ( .A(n58191), .B(n58190), .Z(n7558) );
  NAND U8217 ( .A(n7557), .B(n7558), .Z(n7559) );
  NAND U8218 ( .A(n51294), .B(n7559), .Z(n7560) );
  AND U8219 ( .A(n58193), .B(n58192), .Z(n7561) );
  NAND U8220 ( .A(n7560), .B(n7561), .Z(n7562) );
  NAND U8221 ( .A(n58194), .B(n7562), .Z(n7563) );
  AND U8222 ( .A(n58196), .B(n58195), .Z(n7564) );
  NAND U8223 ( .A(n7563), .B(n7564), .Z(n7565) );
  NANDN U8224 ( .A(n51293), .B(n7565), .Z(n7566) );
  NAND U8225 ( .A(n51292), .B(n7566), .Z(n7567) );
  NAND U8226 ( .A(n58197), .B(n7567), .Z(n58199) );
  AND U8227 ( .A(n58224), .B(n58226), .Z(n7568) );
  NAND U8228 ( .A(n58225), .B(n7568), .Z(n7569) );
  AND U8229 ( .A(n58227), .B(n7569), .Z(n7570) );
  ANDN U8230 ( .B(n58228), .A(n7570), .Z(n7571) );
  NAND U8231 ( .A(n58229), .B(n7571), .Z(n7572) );
  AND U8232 ( .A(n58230), .B(n7572), .Z(n7573) );
  ANDN U8233 ( .B(n51283), .A(n7573), .Z(n7574) );
  NAND U8234 ( .A(n51282), .B(n7574), .Z(n7575) );
  AND U8235 ( .A(n58231), .B(n7575), .Z(n7576) );
  OR U8236 ( .A(n51281), .B(n7576), .Z(n7577) );
  NAND U8237 ( .A(n51280), .B(n7577), .Z(n7578) );
  NANDN U8238 ( .A(n58232), .B(n7578), .Z(n7579) );
  NAND U8239 ( .A(n58233), .B(n7579), .Z(n58236) );
  ANDN U8240 ( .B(n51421), .A(n43630), .Z(n7580) );
  NAND U8241 ( .A(n17451), .B(n7580), .Z(n7581) );
  ANDN U8242 ( .B(n7581), .A(n57693), .Z(n7582) );
  NANDN U8243 ( .A(n7582), .B(n57694), .Z(n7583) );
  AND U8244 ( .A(n51420), .B(n7583), .Z(n7584) );
  NOR U8245 ( .A(n7584), .B(n24263), .Z(n7585) );
  NAND U8246 ( .A(n24262), .B(n7585), .Z(n7586) );
  AND U8247 ( .A(n57698), .B(n7586), .Z(n7587) );
  NOR U8248 ( .A(n24260), .B(n7587), .Z(n7588) );
  NAND U8249 ( .A(n24259), .B(n7588), .Z(n7589) );
  ANDN U8250 ( .B(n7589), .A(n57699), .Z(n7590) );
  NANDN U8251 ( .A(n7590), .B(n57700), .Z(n7591) );
  AND U8252 ( .A(n51417), .B(n7591), .Z(n7592) );
  NOR U8253 ( .A(n24255), .B(n7592), .Z(n7593) );
  NAND U8254 ( .A(n24254), .B(n7593), .Z(n7594) );
  AND U8255 ( .A(n57703), .B(n7594), .Z(n7595) );
  ANDN U8256 ( .B(n51416), .A(n7595), .Z(n7596) );
  XNOR U8257 ( .A(x[5324]), .B(y[5324]), .Z(n7597) );
  NAND U8258 ( .A(n7596), .B(n7597), .Z(n17453) );
  NAND U8259 ( .A(n58265), .B(n58264), .Z(n7598) );
  ANDN U8260 ( .B(n7598), .A(n51270), .Z(n7599) );
  ANDN U8261 ( .B(n58267), .A(n7599), .Z(n7600) );
  NAND U8262 ( .A(n58266), .B(n7600), .Z(n7601) );
  NANDN U8263 ( .A(n58268), .B(n7601), .Z(n7602) );
  AND U8264 ( .A(n58270), .B(n58269), .Z(n7603) );
  NAND U8265 ( .A(n7602), .B(n7603), .Z(n7604) );
  NAND U8266 ( .A(n58271), .B(n7604), .Z(n7605) );
  AND U8267 ( .A(n58273), .B(n58272), .Z(n7606) );
  NAND U8268 ( .A(n7605), .B(n7606), .Z(n7607) );
  NAND U8269 ( .A(n58274), .B(n7607), .Z(n7608) );
  AND U8270 ( .A(n58275), .B(n58276), .Z(n7609) );
  NAND U8271 ( .A(n7608), .B(n7609), .Z(n7610) );
  NANDN U8272 ( .A(n58277), .B(n7610), .Z(n7611) );
  AND U8273 ( .A(n58279), .B(n58278), .Z(n7612) );
  NAND U8274 ( .A(n7611), .B(n7612), .Z(n7613) );
  NANDN U8275 ( .A(n58280), .B(n7613), .Z(n7614) );
  AND U8276 ( .A(n58281), .B(n7614), .Z(n58283) );
  AND U8277 ( .A(n58380), .B(n51249), .Z(n7615) );
  NAND U8278 ( .A(n51250), .B(n7615), .Z(n7616) );
  NAND U8279 ( .A(n58381), .B(n7616), .Z(n7617) );
  NANDN U8280 ( .A(n51248), .B(n7617), .Z(n7618) );
  NAND U8281 ( .A(n51247), .B(n7618), .Z(n7619) );
  AND U8282 ( .A(n58382), .B(n7619), .Z(n7620) );
  NAND U8283 ( .A(n58383), .B(n7620), .Z(n7621) );
  AND U8284 ( .A(n51245), .B(n51246), .Z(n7622) );
  NANDN U8285 ( .A(n58384), .B(n7621), .Z(n7623) );
  NAND U8286 ( .A(n7622), .B(n7623), .Z(n7624) );
  ANDN U8287 ( .B(n58386), .A(n58387), .Z(n7625) );
  NANDN U8288 ( .A(n58385), .B(n7624), .Z(n7626) );
  NAND U8289 ( .A(n7625), .B(n7626), .Z(n58388) );
  ANDN U8290 ( .B(n58422), .A(n58421), .Z(n7627) );
  NAND U8291 ( .A(n58419), .B(n58418), .Z(n7628) );
  AND U8292 ( .A(n7627), .B(n7628), .Z(n7629) );
  AND U8293 ( .A(n58425), .B(n58424), .Z(n7630) );
  OR U8294 ( .A(n58423), .B(n7629), .Z(n7631) );
  AND U8295 ( .A(n7630), .B(n7631), .Z(n7632) );
  AND U8296 ( .A(n58427), .B(n58428), .Z(n7633) );
  NANDN U8297 ( .A(n7632), .B(n58426), .Z(n7634) );
  AND U8298 ( .A(n7633), .B(n7634), .Z(n7635) );
  AND U8299 ( .A(n51238), .B(n51237), .Z(n7636) );
  OR U8300 ( .A(n58429), .B(n7635), .Z(n7637) );
  AND U8301 ( .A(n7636), .B(n7637), .Z(n7638) );
  AND U8302 ( .A(n58431), .B(n58432), .Z(n7639) );
  OR U8303 ( .A(n58430), .B(n7638), .Z(n7640) );
  AND U8304 ( .A(n7639), .B(n7640), .Z(n7641) );
  AND U8305 ( .A(n58435), .B(n58434), .Z(n7642) );
  OR U8306 ( .A(n58433), .B(n7641), .Z(n7643) );
  AND U8307 ( .A(n7642), .B(n7643), .Z(n58438) );
  NAND U8308 ( .A(n58463), .B(n51230), .Z(n7644) );
  NANDN U8309 ( .A(n51229), .B(n7644), .Z(n7645) );
  NAND U8310 ( .A(n51228), .B(n7645), .Z(n7646) );
  AND U8311 ( .A(n58466), .B(n58465), .Z(n7647) );
  NANDN U8312 ( .A(n58464), .B(n7646), .Z(n7648) );
  NAND U8313 ( .A(n7647), .B(n7648), .Z(n7649) );
  AND U8314 ( .A(n58468), .B(n58469), .Z(n7650) );
  NANDN U8315 ( .A(n58467), .B(n7649), .Z(n7651) );
  NAND U8316 ( .A(n7650), .B(n7651), .Z(n7652) );
  NAND U8317 ( .A(n58470), .B(n7652), .Z(n7653) );
  AND U8318 ( .A(n58472), .B(n7653), .Z(n7654) );
  NAND U8319 ( .A(n7654), .B(n58471), .Z(n7655) );
  NAND U8320 ( .A(n58473), .B(n7655), .Z(n58474) );
  NAND U8321 ( .A(n58506), .B(n58505), .Z(n7656) );
  AND U8322 ( .A(n58509), .B(n7656), .Z(n7657) );
  AND U8323 ( .A(n58512), .B(n58511), .Z(n7658) );
  OR U8324 ( .A(n7657), .B(n58510), .Z(n7659) );
  AND U8325 ( .A(n7658), .B(n7659), .Z(n7660) );
  AND U8326 ( .A(n58515), .B(n58514), .Z(n7661) );
  NANDN U8327 ( .A(n7660), .B(n58513), .Z(n7662) );
  AND U8328 ( .A(n7661), .B(n7662), .Z(n7663) );
  AND U8329 ( .A(n51216), .B(n51215), .Z(n7664) );
  OR U8330 ( .A(n58516), .B(n7663), .Z(n7665) );
  AND U8331 ( .A(n7664), .B(n7665), .Z(n7666) );
  ANDN U8332 ( .B(n58519), .A(n58518), .Z(n7667) );
  NANDN U8333 ( .A(n7666), .B(n58517), .Z(n7668) );
  AND U8334 ( .A(n7667), .B(n7668), .Z(n7669) );
  ANDN U8335 ( .B(n58520), .A(n58521), .Z(n7670) );
  NANDN U8336 ( .A(n7669), .B(n51214), .Z(n7671) );
  AND U8337 ( .A(n7670), .B(n7671), .Z(n58524) );
  NANDN U8338 ( .A(n58552), .B(n58551), .Z(n7672) );
  AND U8339 ( .A(n51205), .B(n7672), .Z(n7673) );
  ANDN U8340 ( .B(n58553), .A(n7673), .Z(n7674) );
  NAND U8341 ( .A(n58554), .B(n7674), .Z(n7675) );
  NAND U8342 ( .A(n58555), .B(n7675), .Z(n7676) );
  AND U8343 ( .A(n58557), .B(n58556), .Z(n7677) );
  NAND U8344 ( .A(n7676), .B(n7677), .Z(n7678) );
  NANDN U8345 ( .A(n58558), .B(n7678), .Z(n7679) );
  AND U8346 ( .A(n51204), .B(n51203), .Z(n7680) );
  NAND U8347 ( .A(n7679), .B(n7680), .Z(n7681) );
  NANDN U8348 ( .A(n58559), .B(n7681), .Z(n7682) );
  AND U8349 ( .A(n58561), .B(n58560), .Z(n7683) );
  NAND U8350 ( .A(n7682), .B(n7683), .Z(n7684) );
  NAND U8351 ( .A(n51202), .B(n7684), .Z(n7685) );
  AND U8352 ( .A(n58562), .B(n7685), .Z(n58564) );
  NAND U8353 ( .A(n58593), .B(n58594), .Z(n7686) );
  NANDN U8354 ( .A(n58595), .B(n7686), .Z(n7687) );
  NAND U8355 ( .A(n58596), .B(n7687), .Z(n7688) );
  AND U8356 ( .A(n58597), .B(n58598), .Z(n7689) );
  NAND U8357 ( .A(n7688), .B(n7689), .Z(n7690) );
  NANDN U8358 ( .A(n58599), .B(n7690), .Z(n7691) );
  AND U8359 ( .A(n58600), .B(n58601), .Z(n7692) );
  NAND U8360 ( .A(n7691), .B(n7692), .Z(n7693) );
  NANDN U8361 ( .A(n58602), .B(n7693), .Z(n7694) );
  AND U8362 ( .A(n58604), .B(n58603), .Z(n7695) );
  NAND U8363 ( .A(n7694), .B(n7695), .Z(n7696) );
  NANDN U8364 ( .A(n58605), .B(n7696), .Z(n7697) );
  AND U8365 ( .A(n51194), .B(n51193), .Z(n7698) );
  NAND U8366 ( .A(n7697), .B(n7698), .Z(n7699) );
  NAND U8367 ( .A(n58606), .B(n7699), .Z(n7700) );
  AND U8368 ( .A(n58607), .B(n58608), .Z(n7701) );
  NAND U8369 ( .A(n7700), .B(n7701), .Z(n7702) );
  NAND U8370 ( .A(n58609), .B(n7702), .Z(n7703) );
  NANDN U8371 ( .A(n58610), .B(n7703), .Z(n58611) );
  AND U8372 ( .A(n58641), .B(n58642), .Z(n7704) );
  ANDN U8373 ( .B(n58646), .A(n58645), .Z(n7705) );
  OR U8374 ( .A(n58643), .B(n7704), .Z(n7706) );
  AND U8375 ( .A(n7705), .B(n7706), .Z(n7707) );
  AND U8376 ( .A(n58649), .B(n58648), .Z(n7708) );
  OR U8377 ( .A(n58647), .B(n7707), .Z(n7709) );
  AND U8378 ( .A(n7708), .B(n7709), .Z(n7710) );
  AND U8379 ( .A(n58651), .B(n58652), .Z(n7711) );
  OR U8380 ( .A(n58650), .B(n7710), .Z(n7712) );
  AND U8381 ( .A(n7711), .B(n7712), .Z(n7713) );
  AND U8382 ( .A(n51184), .B(n51183), .Z(n7714) );
  OR U8383 ( .A(n58653), .B(n7713), .Z(n7715) );
  AND U8384 ( .A(n7714), .B(n7715), .Z(n7716) );
  AND U8385 ( .A(n58656), .B(n58655), .Z(n7717) );
  NANDN U8386 ( .A(n7716), .B(n58654), .Z(n7718) );
  AND U8387 ( .A(n7717), .B(n7718), .Z(n7719) );
  AND U8388 ( .A(n58659), .B(n58658), .Z(n7720) );
  OR U8389 ( .A(n7719), .B(n58657), .Z(n7721) );
  AND U8390 ( .A(n7720), .B(n7721), .Z(n58661) );
  AND U8391 ( .A(n58690), .B(n58691), .Z(n7722) );
  NAND U8392 ( .A(n58692), .B(n7722), .Z(n7723) );
  NANDN U8393 ( .A(n58693), .B(n7723), .Z(n7724) );
  AND U8394 ( .A(n51172), .B(n51171), .Z(n7725) );
  NAND U8395 ( .A(n7724), .B(n7725), .Z(n7726) );
  NAND U8396 ( .A(n58694), .B(n7726), .Z(n7727) );
  AND U8397 ( .A(n58695), .B(n58696), .Z(n7728) );
  NAND U8398 ( .A(n7727), .B(n7728), .Z(n7729) );
  NANDN U8399 ( .A(n58697), .B(n7729), .Z(n7730) );
  ANDN U8400 ( .B(n58698), .A(n58699), .Z(n7731) );
  NAND U8401 ( .A(n7730), .B(n7731), .Z(n7732) );
  NAND U8402 ( .A(n58700), .B(n7732), .Z(n7733) );
  AND U8403 ( .A(n58701), .B(n7733), .Z(n7734) );
  AND U8404 ( .A(n58704), .B(n58703), .Z(n7735) );
  NANDN U8405 ( .A(n7734), .B(n58702), .Z(n7736) );
  AND U8406 ( .A(n7735), .B(n7736), .Z(n7737) );
  AND U8407 ( .A(n58706), .B(n58705), .Z(n7738) );
  NANDN U8408 ( .A(n7737), .B(n51170), .Z(n7739) );
  AND U8409 ( .A(n7738), .B(n7739), .Z(n58708) );
  ANDN U8410 ( .B(n51163), .A(n51162), .Z(n7740) );
  OR U8411 ( .A(n58739), .B(n58738), .Z(n7741) );
  NAND U8412 ( .A(n7740), .B(n7741), .Z(n7742) );
  NAND U8413 ( .A(n58740), .B(n7742), .Z(n7743) );
  AND U8414 ( .A(n58742), .B(n7743), .Z(n7744) );
  NANDN U8415 ( .A(n58741), .B(n7744), .Z(n7745) );
  NAND U8416 ( .A(n51161), .B(n7745), .Z(n7746) );
  AND U8417 ( .A(n58744), .B(n7746), .Z(n7747) );
  NANDN U8418 ( .A(n58743), .B(n7747), .Z(n7748) );
  ANDN U8419 ( .B(n58746), .A(n58747), .Z(n7749) );
  NANDN U8420 ( .A(n58745), .B(n7748), .Z(n7750) );
  NAND U8421 ( .A(n7749), .B(n7750), .Z(n7751) );
  ANDN U8422 ( .B(n51160), .A(n51159), .Z(n7752) );
  NANDN U8423 ( .A(n58748), .B(n7751), .Z(n7753) );
  NAND U8424 ( .A(n7752), .B(n7753), .Z(n7754) );
  NANDN U8425 ( .A(n58749), .B(n7754), .Z(n7755) );
  NAND U8426 ( .A(n58750), .B(n7755), .Z(n58751) );
  ANDN U8427 ( .B(n51155), .A(n51154), .Z(n58765) );
  AND U8428 ( .A(n23757), .B(n18215), .Z(n7756) );
  NAND U8429 ( .A(n51262), .B(n7756), .Z(n7757) );
  AND U8430 ( .A(n58327), .B(n7757), .Z(n7758) );
  ANDN U8431 ( .B(n58329), .A(n7758), .Z(n7759) );
  XNOR U8432 ( .A(x[5828]), .B(y[5828]), .Z(n7760) );
  NAND U8433 ( .A(n7759), .B(n7760), .Z(n7761) );
  NAND U8434 ( .A(n51260), .B(n7761), .Z(n7762) );
  AND U8435 ( .A(n23755), .B(n7762), .Z(n7763) );
  NANDN U8436 ( .A(n44845), .B(n7763), .Z(n7764) );
  ANDN U8437 ( .B(n23752), .A(n23753), .Z(n7765) );
  NANDN U8438 ( .A(n58332), .B(n7764), .Z(n7766) );
  NAND U8439 ( .A(n7765), .B(n7766), .Z(n7767) );
  NAND U8440 ( .A(n58336), .B(n7767), .Z(n7768) );
  NAND U8441 ( .A(n58337), .B(n7768), .Z(n7769) );
  AND U8442 ( .A(n58338), .B(n7769), .Z(n7770) );
  ANDN U8443 ( .B(n58340), .A(n7770), .Z(n7771) );
  XNOR U8444 ( .A(x[5836]), .B(y[5836]), .Z(n7772) );
  NAND U8445 ( .A(n7771), .B(n7772), .Z(n18218) );
  ANDN U8446 ( .B(n58794), .A(n58793), .Z(n7773) );
  NANDN U8447 ( .A(n51146), .B(n58792), .Z(n7774) );
  AND U8448 ( .A(n7773), .B(n7774), .Z(n7775) );
  ANDN U8449 ( .B(n51145), .A(n51144), .Z(n7776) );
  OR U8450 ( .A(n58795), .B(n7775), .Z(n7777) );
  AND U8451 ( .A(n7776), .B(n7777), .Z(n7778) );
  ANDN U8452 ( .B(n58797), .A(n58798), .Z(n7779) );
  NANDN U8453 ( .A(n7778), .B(n58796), .Z(n7780) );
  AND U8454 ( .A(n7779), .B(n7780), .Z(n7781) );
  ANDN U8455 ( .B(n58799), .A(n58800), .Z(n7782) );
  NANDN U8456 ( .A(n7781), .B(n51143), .Z(n7783) );
  AND U8457 ( .A(n7782), .B(n7783), .Z(n7784) );
  ANDN U8458 ( .B(n58802), .A(n58801), .Z(n7785) );
  OR U8459 ( .A(n51142), .B(n7784), .Z(n7786) );
  AND U8460 ( .A(n7785), .B(n7786), .Z(n58804) );
  ANDN U8461 ( .B(n58815), .A(n58816), .Z(n58817) );
  NAND U8462 ( .A(n58844), .B(n58845), .Z(n7787) );
  AND U8463 ( .A(n58846), .B(n7787), .Z(n7788) );
  OR U8464 ( .A(n51127), .B(n7788), .Z(n7789) );
  NAND U8465 ( .A(n51126), .B(n7789), .Z(n7790) );
  NANDN U8466 ( .A(n58847), .B(n7790), .Z(n7791) );
  AND U8467 ( .A(n58849), .B(n58848), .Z(n7792) );
  NAND U8468 ( .A(n7791), .B(n7792), .Z(n7793) );
  NAND U8469 ( .A(n58850), .B(n7793), .Z(n7794) );
  AND U8470 ( .A(n51125), .B(n51124), .Z(n7795) );
  NAND U8471 ( .A(n7794), .B(n7795), .Z(n7796) );
  NAND U8472 ( .A(n58851), .B(n7796), .Z(n7797) );
  AND U8473 ( .A(n58853), .B(n58852), .Z(n7798) );
  NAND U8474 ( .A(n7797), .B(n7798), .Z(n7799) );
  NAND U8475 ( .A(n58854), .B(n7799), .Z(n58855) );
  NAND U8476 ( .A(n58882), .B(n58883), .Z(n7800) );
  NAND U8477 ( .A(n58884), .B(n7800), .Z(n7801) );
  AND U8478 ( .A(n51116), .B(n7801), .Z(n7802) );
  NANDN U8479 ( .A(n51115), .B(n7802), .Z(n7803) );
  NAND U8480 ( .A(n58885), .B(n7803), .Z(n7804) );
  AND U8481 ( .A(n58887), .B(n7804), .Z(n7805) );
  NANDN U8482 ( .A(n58886), .B(n7805), .Z(n7806) );
  ANDN U8483 ( .B(n58890), .A(n58889), .Z(n7807) );
  NANDN U8484 ( .A(n58888), .B(n7806), .Z(n7808) );
  NAND U8485 ( .A(n7807), .B(n7808), .Z(n7809) );
  NAND U8486 ( .A(n58891), .B(n7809), .Z(n7810) );
  AND U8487 ( .A(n58892), .B(n7810), .Z(n7811) );
  NAND U8488 ( .A(n7811), .B(n58893), .Z(n7812) );
  NAND U8489 ( .A(n58894), .B(n7812), .Z(n7813) );
  AND U8490 ( .A(n51113), .B(n7813), .Z(n7814) );
  NAND U8491 ( .A(n7814), .B(n51114), .Z(n58895) );
  NAND U8492 ( .A(n58928), .B(n58927), .Z(n7815) );
  AND U8493 ( .A(n58929), .B(n7815), .Z(n7816) );
  NOR U8494 ( .A(n51105), .B(n7816), .Z(n7817) );
  NAND U8495 ( .A(n51106), .B(n7817), .Z(n7818) );
  NANDN U8496 ( .A(n51104), .B(n7818), .Z(n7819) );
  ANDN U8497 ( .B(n58931), .A(n58930), .Z(n7820) );
  NAND U8498 ( .A(n7819), .B(n7820), .Z(n7821) );
  NANDN U8499 ( .A(n58932), .B(n7821), .Z(n7822) );
  AND U8500 ( .A(n58933), .B(n58934), .Z(n7823) );
  NAND U8501 ( .A(n7822), .B(n7823), .Z(n7824) );
  NAND U8502 ( .A(n58935), .B(n7824), .Z(n7825) );
  ANDN U8503 ( .B(n51103), .A(n51102), .Z(n7826) );
  NAND U8504 ( .A(n7825), .B(n7826), .Z(n7827) );
  NAND U8505 ( .A(n58936), .B(n7827), .Z(n7828) );
  ANDN U8506 ( .B(n58938), .A(n58937), .Z(n7829) );
  NAND U8507 ( .A(n7828), .B(n7829), .Z(n7830) );
  NANDN U8508 ( .A(n58939), .B(n7830), .Z(n58941) );
  NAND U8509 ( .A(n58972), .B(n58971), .Z(n7831) );
  AND U8510 ( .A(n58974), .B(n7831), .Z(n7832) );
  ANDN U8511 ( .B(n58977), .A(n7832), .Z(n7833) );
  NAND U8512 ( .A(n58976), .B(n7833), .Z(n7834) );
  ANDN U8513 ( .B(n7834), .A(n58978), .Z(n7835) );
  NOR U8514 ( .A(n58979), .B(n7835), .Z(n7836) );
  NAND U8515 ( .A(n58980), .B(n7836), .Z(n7837) );
  ANDN U8516 ( .B(n7837), .A(n58981), .Z(n7838) );
  NOR U8517 ( .A(n7838), .B(n51095), .Z(n7839) );
  NAND U8518 ( .A(n51096), .B(n7839), .Z(n7840) );
  AND U8519 ( .A(n58982), .B(n7840), .Z(n7841) );
  NOR U8520 ( .A(n58984), .B(n7841), .Z(n7842) );
  NAND U8521 ( .A(n58983), .B(n7842), .Z(n7843) );
  ANDN U8522 ( .B(n7843), .A(n58985), .Z(n7844) );
  NOR U8523 ( .A(n7844), .B(n58987), .Z(n7845) );
  NAND U8524 ( .A(n58986), .B(n7845), .Z(n7846) );
  NAND U8525 ( .A(n58988), .B(n7846), .Z(n7847) );
  ANDN U8526 ( .B(n7847), .A(n58989), .Z(n58991) );
  AND U8527 ( .A(n59016), .B(n59015), .Z(n7848) );
  NAND U8528 ( .A(n59017), .B(n7848), .Z(n7849) );
  NAND U8529 ( .A(n59018), .B(n7849), .Z(n7850) );
  ANDN U8530 ( .B(n59019), .A(n59020), .Z(n7851) );
  NAND U8531 ( .A(n7850), .B(n7851), .Z(n7852) );
  NANDN U8532 ( .A(n59021), .B(n7852), .Z(n7853) );
  ANDN U8533 ( .B(n51083), .A(n51082), .Z(n7854) );
  NAND U8534 ( .A(n7853), .B(n7854), .Z(n7855) );
  NANDN U8535 ( .A(n59022), .B(n7855), .Z(n7856) );
  ANDN U8536 ( .B(n59023), .A(n59024), .Z(n7857) );
  NAND U8537 ( .A(n7856), .B(n7857), .Z(n7858) );
  NANDN U8538 ( .A(n59025), .B(n7858), .Z(n7859) );
  ANDN U8539 ( .B(n59027), .A(n59026), .Z(n7860) );
  NAND U8540 ( .A(n7859), .B(n7860), .Z(n7861) );
  NAND U8541 ( .A(n59028), .B(n7861), .Z(n7862) );
  AND U8542 ( .A(n59029), .B(n7862), .Z(n59032) );
  ANDN U8543 ( .B(n59044), .A(n59045), .Z(n59046) );
  AND U8544 ( .A(n51068), .B(n51067), .Z(n7863) );
  OR U8545 ( .A(n59073), .B(n59074), .Z(n7864) );
  AND U8546 ( .A(n7863), .B(n7864), .Z(n7865) );
  AND U8547 ( .A(n59077), .B(n59076), .Z(n7866) );
  OR U8548 ( .A(n59075), .B(n7865), .Z(n7867) );
  AND U8549 ( .A(n7866), .B(n7867), .Z(n7868) );
  OR U8550 ( .A(n59078), .B(n7868), .Z(n7869) );
  AND U8551 ( .A(n59079), .B(n7869), .Z(n7870) );
  AND U8552 ( .A(n51065), .B(n51066), .Z(n7871) );
  NANDN U8553 ( .A(n7870), .B(n59080), .Z(n7872) );
  AND U8554 ( .A(n7871), .B(n7872), .Z(n7873) );
  NANDN U8555 ( .A(n7873), .B(n59081), .Z(n7874) );
  NANDN U8556 ( .A(n51064), .B(n7874), .Z(n7875) );
  NAND U8557 ( .A(n51063), .B(n7875), .Z(n59084) );
  AND U8558 ( .A(n59120), .B(n51058), .Z(n7876) );
  NAND U8559 ( .A(n51059), .B(n7876), .Z(n7877) );
  NAND U8560 ( .A(n59121), .B(n7877), .Z(n7878) );
  AND U8561 ( .A(n59123), .B(n59122), .Z(n7879) );
  NAND U8562 ( .A(n7878), .B(n7879), .Z(n7880) );
  NANDN U8563 ( .A(n59124), .B(n7880), .Z(n7881) );
  AND U8564 ( .A(n59125), .B(n59126), .Z(n7882) );
  NAND U8565 ( .A(n7881), .B(n7882), .Z(n7883) );
  NANDN U8566 ( .A(n59127), .B(n7883), .Z(n7884) );
  AND U8567 ( .A(n59129), .B(n59128), .Z(n7885) );
  NAND U8568 ( .A(n7884), .B(n7885), .Z(n7886) );
  NAND U8569 ( .A(n59130), .B(n7886), .Z(n7887) );
  AND U8570 ( .A(n51056), .B(n51057), .Z(n7888) );
  NAND U8571 ( .A(n7887), .B(n7888), .Z(n7889) );
  NAND U8572 ( .A(n59131), .B(n7889), .Z(n7890) );
  AND U8573 ( .A(n59133), .B(n59132), .Z(n7891) );
  NAND U8574 ( .A(n7890), .B(n7891), .Z(n7892) );
  NANDN U8575 ( .A(n59134), .B(n7892), .Z(n59135) );
  NAND U8576 ( .A(n59205), .B(n59204), .Z(n7893) );
  ANDN U8577 ( .B(n7893), .A(n59206), .Z(n7894) );
  NOR U8578 ( .A(n59208), .B(n7894), .Z(n7895) );
  NAND U8579 ( .A(n59209), .B(n7895), .Z(n7896) );
  NAND U8580 ( .A(n51045), .B(n7896), .Z(n7897) );
  AND U8581 ( .A(n59211), .B(n59210), .Z(n7898) );
  NAND U8582 ( .A(n7897), .B(n7898), .Z(n7899) );
  NAND U8583 ( .A(n59212), .B(n7899), .Z(n7900) );
  AND U8584 ( .A(n59214), .B(n59213), .Z(n7901) );
  NAND U8585 ( .A(n7900), .B(n7901), .Z(n7902) );
  NANDN U8586 ( .A(n59215), .B(n7902), .Z(n7903) );
  AND U8587 ( .A(n51044), .B(n51043), .Z(n7904) );
  NAND U8588 ( .A(n7903), .B(n7904), .Z(n7905) );
  NAND U8589 ( .A(n59216), .B(n7905), .Z(n7906) );
  AND U8590 ( .A(n59218), .B(n59217), .Z(n7907) );
  NAND U8591 ( .A(n7906), .B(n7907), .Z(n7908) );
  NANDN U8592 ( .A(n59219), .B(n7908), .Z(n59220) );
  NAND U8593 ( .A(n18900), .B(n58860), .Z(n7909) );
  AND U8594 ( .A(n58862), .B(n7909), .Z(n7910) );
  NOR U8595 ( .A(n58863), .B(n7910), .Z(n7911) );
  NAND U8596 ( .A(n23339), .B(n7911), .Z(n7912) );
  AND U8597 ( .A(n58865), .B(n7912), .Z(n7913) );
  NOR U8598 ( .A(n45822), .B(n7913), .Z(n7914) );
  NAND U8599 ( .A(n23337), .B(n7914), .Z(n7915) );
  ANDN U8600 ( .B(n7915), .A(n58866), .Z(n7916) );
  ANDN U8601 ( .B(n23335), .A(n7916), .Z(n7917) );
  NAND U8602 ( .A(n58870), .B(n7917), .Z(n7918) );
  ANDN U8603 ( .B(n7918), .A(n58872), .Z(n7919) );
  ANDN U8604 ( .B(n23333), .A(n7919), .Z(n7920) );
  NAND U8605 ( .A(n58873), .B(n7920), .Z(n7921) );
  ANDN U8606 ( .B(n7921), .A(n51118), .Z(n7922) );
  NANDN U8607 ( .A(n7922), .B(n51117), .Z(n7923) );
  NANDN U8608 ( .A(n58874), .B(n7923), .Z(n7924) );
  NAND U8609 ( .A(n58875), .B(n7924), .Z(n7925) );
  XNOR U8610 ( .A(x[6268]), .B(y[6268]), .Z(n7926) );
  NANDN U8611 ( .A(n7925), .B(n7926), .Z(n18905) );
  NANDN U8612 ( .A(n59248), .B(n59247), .Z(n7927) );
  AND U8613 ( .A(n59249), .B(n7927), .Z(n7928) );
  ANDN U8614 ( .B(n59251), .A(n7928), .Z(n7929) );
  NAND U8615 ( .A(n59250), .B(n7929), .Z(n7930) );
  NANDN U8616 ( .A(n59252), .B(n7930), .Z(n7931) );
  AND U8617 ( .A(n59254), .B(n59253), .Z(n7932) );
  NAND U8618 ( .A(n7931), .B(n7932), .Z(n7933) );
  NAND U8619 ( .A(n59255), .B(n7933), .Z(n7934) );
  AND U8620 ( .A(n59257), .B(n59256), .Z(n7935) );
  NAND U8621 ( .A(n7934), .B(n7935), .Z(n7936) );
  NANDN U8622 ( .A(n59258), .B(n7936), .Z(n7937) );
  AND U8623 ( .A(n51032), .B(n51033), .Z(n7938) );
  NAND U8624 ( .A(n7937), .B(n7938), .Z(n7939) );
  NANDN U8625 ( .A(n59259), .B(n7939), .Z(n7940) );
  AND U8626 ( .A(n59261), .B(n59260), .Z(n7941) );
  NAND U8627 ( .A(n7940), .B(n7941), .Z(n7942) );
  NANDN U8628 ( .A(n59262), .B(n7942), .Z(n59263) );
  NAND U8629 ( .A(n59295), .B(n59294), .Z(n7943) );
  NANDN U8630 ( .A(n59296), .B(n7943), .Z(n7944) );
  AND U8631 ( .A(n59297), .B(n7944), .Z(n7945) );
  NAND U8632 ( .A(n7945), .B(n59298), .Z(n7946) );
  NAND U8633 ( .A(n51024), .B(n7946), .Z(n7947) );
  AND U8634 ( .A(n59299), .B(n7947), .Z(n7948) );
  NAND U8635 ( .A(n59300), .B(n7948), .Z(n7949) );
  NANDN U8636 ( .A(n59301), .B(n7949), .Z(n7950) );
  AND U8637 ( .A(n59302), .B(n7950), .Z(n7951) );
  NAND U8638 ( .A(n59303), .B(n7951), .Z(n7952) );
  NAND U8639 ( .A(n59304), .B(n7952), .Z(n7953) );
  AND U8640 ( .A(n51022), .B(n7953), .Z(n7954) );
  NAND U8641 ( .A(n7954), .B(n51023), .Z(n7955) );
  NAND U8642 ( .A(n59305), .B(n7955), .Z(n7956) );
  AND U8643 ( .A(n59306), .B(n7956), .Z(n7957) );
  NAND U8644 ( .A(n7957), .B(n59307), .Z(n59308) );
  AND U8645 ( .A(n59342), .B(n59341), .Z(n7958) );
  NAND U8646 ( .A(n59339), .B(n59340), .Z(n7959) );
  AND U8647 ( .A(n7958), .B(n7959), .Z(n7960) );
  NANDN U8648 ( .A(n7960), .B(n59343), .Z(n7961) );
  NANDN U8649 ( .A(n51014), .B(n7961), .Z(n7962) );
  NAND U8650 ( .A(n59344), .B(n7962), .Z(n7963) );
  NAND U8651 ( .A(n59345), .B(n7963), .Z(n7964) );
  NAND U8652 ( .A(n59346), .B(n7964), .Z(n7965) );
  AND U8653 ( .A(n59347), .B(n7965), .Z(n7966) );
  NAND U8654 ( .A(n59348), .B(n7966), .Z(n7967) );
  NAND U8655 ( .A(n59349), .B(n7967), .Z(n7968) );
  AND U8656 ( .A(n59350), .B(n7968), .Z(n7969) );
  AND U8657 ( .A(n51012), .B(n51013), .Z(n7970) );
  OR U8658 ( .A(n7969), .B(n59351), .Z(n7971) );
  AND U8659 ( .A(n7970), .B(n7971), .Z(n7972) );
  NANDN U8660 ( .A(n7972), .B(n59352), .Z(n7973) );
  AND U8661 ( .A(n59353), .B(n7973), .Z(n59354) );
  NOR U8662 ( .A(n51003), .B(n51004), .Z(n7974) );
  NANDN U8663 ( .A(n59386), .B(n59385), .Z(n7975) );
  NAND U8664 ( .A(n7974), .B(n7975), .Z(n7976) );
  NAND U8665 ( .A(n59387), .B(n7976), .Z(n7977) );
  AND U8666 ( .A(n59389), .B(n7977), .Z(n7978) );
  NANDN U8667 ( .A(n59388), .B(n7978), .Z(n7979) );
  NAND U8668 ( .A(n59390), .B(n7979), .Z(n7980) );
  AND U8669 ( .A(n51001), .B(n7980), .Z(n7981) );
  NAND U8670 ( .A(n7981), .B(n51000), .Z(n7982) );
  NAND U8671 ( .A(n50999), .B(n7982), .Z(n7983) );
  AND U8672 ( .A(n59392), .B(n7983), .Z(n7984) );
  NANDN U8673 ( .A(n59391), .B(n7984), .Z(n7985) );
  NAND U8674 ( .A(n59393), .B(n7985), .Z(n7986) );
  AND U8675 ( .A(n50998), .B(n7986), .Z(n7987) );
  NANDN U8676 ( .A(n50997), .B(n7987), .Z(n7988) );
  NANDN U8677 ( .A(n59394), .B(n7988), .Z(n59395) );
  ANDN U8678 ( .B(n50992), .A(n50991), .Z(n59412) );
  ANDN U8679 ( .B(n50982), .A(n50983), .Z(n7989) );
  NANDN U8680 ( .A(n59441), .B(n59440), .Z(n7990) );
  NAND U8681 ( .A(n7989), .B(n7990), .Z(n7991) );
  NAND U8682 ( .A(n59442), .B(n7991), .Z(n7992) );
  AND U8683 ( .A(n59444), .B(n7992), .Z(n7993) );
  NANDN U8684 ( .A(n59443), .B(n7993), .Z(n7994) );
  NAND U8685 ( .A(n59445), .B(n7994), .Z(n7995) );
  AND U8686 ( .A(n50981), .B(n7995), .Z(n7996) );
  NANDN U8687 ( .A(n50980), .B(n7996), .Z(n7997) );
  ANDN U8688 ( .B(n59448), .A(n59447), .Z(n7998) );
  NANDN U8689 ( .A(n59446), .B(n7997), .Z(n7999) );
  NAND U8690 ( .A(n7998), .B(n7999), .Z(n8000) );
  AND U8691 ( .A(n50979), .B(n50978), .Z(n8001) );
  NANDN U8692 ( .A(n59449), .B(n8000), .Z(n8002) );
  NAND U8693 ( .A(n8001), .B(n8002), .Z(n8003) );
  NAND U8694 ( .A(n59450), .B(n8003), .Z(n8004) );
  NANDN U8695 ( .A(n59451), .B(n8004), .Z(n59452) );
  NAND U8696 ( .A(n59485), .B(n59484), .Z(n8005) );
  ANDN U8697 ( .B(n8005), .A(n59486), .Z(n8006) );
  ANDN U8698 ( .B(n59487), .A(n8006), .Z(n8007) );
  NAND U8699 ( .A(n59488), .B(n8007), .Z(n8008) );
  NANDN U8700 ( .A(n59489), .B(n8008), .Z(n8009) );
  AND U8701 ( .A(n59491), .B(n59490), .Z(n8010) );
  NAND U8702 ( .A(n8009), .B(n8010), .Z(n8011) );
  NAND U8703 ( .A(n59492), .B(n8011), .Z(n8012) );
  ANDN U8704 ( .B(n59494), .A(n59493), .Z(n8013) );
  NAND U8705 ( .A(n8012), .B(n8013), .Z(n8014) );
  NAND U8706 ( .A(n59495), .B(n8014), .Z(n8015) );
  NAND U8707 ( .A(n59496), .B(n8015), .Z(n8016) );
  NAND U8708 ( .A(n59497), .B(n8016), .Z(n8017) );
  AND U8709 ( .A(n59498), .B(n8017), .Z(n8018) );
  AND U8710 ( .A(n59499), .B(n8018), .Z(n59502) );
  AND U8711 ( .A(n23124), .B(n51050), .Z(n8019) );
  NAND U8712 ( .A(n59182), .B(n19256), .Z(n8020) );
  AND U8713 ( .A(n8019), .B(n8020), .Z(n8021) );
  AND U8714 ( .A(n59185), .B(n23122), .Z(n8022) );
  NANDN U8715 ( .A(n8021), .B(n59183), .Z(n8023) );
  AND U8716 ( .A(n8022), .B(n8023), .Z(n8024) );
  AND U8717 ( .A(n59187), .B(n23120), .Z(n8025) );
  NANDN U8718 ( .A(n8024), .B(n59186), .Z(n8026) );
  AND U8719 ( .A(n8025), .B(n8026), .Z(n8027) );
  AND U8720 ( .A(n23118), .B(n59191), .Z(n8028) );
  OR U8721 ( .A(n59190), .B(n8027), .Z(n8029) );
  AND U8722 ( .A(n8028), .B(n8029), .Z(n8030) );
  AND U8723 ( .A(n51048), .B(n46396), .Z(n8031) );
  NANDN U8724 ( .A(n8030), .B(n59193), .Z(n8032) );
  AND U8725 ( .A(n8031), .B(n8032), .Z(n8033) );
  AND U8726 ( .A(n23116), .B(n59196), .Z(n8034) );
  OR U8727 ( .A(n8033), .B(n59194), .Z(n8035) );
  NAND U8728 ( .A(n8034), .B(n8035), .Z(n8036) );
  NAND U8729 ( .A(n59197), .B(n8036), .Z(n19257) );
  NAND U8730 ( .A(n59534), .B(n59533), .Z(n8037) );
  AND U8731 ( .A(n59535), .B(n8037), .Z(n8038) );
  NOR U8732 ( .A(n59536), .B(n8038), .Z(n8039) );
  NAND U8733 ( .A(n59537), .B(n8039), .Z(n8040) );
  NANDN U8734 ( .A(n59538), .B(n8040), .Z(n8041) );
  ANDN U8735 ( .B(n50960), .A(n50959), .Z(n8042) );
  NAND U8736 ( .A(n8041), .B(n8042), .Z(n8043) );
  NAND U8737 ( .A(n59539), .B(n8043), .Z(n8044) );
  ANDN U8738 ( .B(n59541), .A(n59540), .Z(n8045) );
  NAND U8739 ( .A(n8044), .B(n8045), .Z(n8046) );
  NAND U8740 ( .A(n59542), .B(n8046), .Z(n8047) );
  ANDN U8741 ( .B(n59543), .A(n50958), .Z(n8048) );
  NAND U8742 ( .A(n8047), .B(n8048), .Z(n8049) );
  NANDN U8743 ( .A(n59544), .B(n8049), .Z(n8050) );
  ANDN U8744 ( .B(n59546), .A(n59545), .Z(n8051) );
  NAND U8745 ( .A(n8050), .B(n8051), .Z(n8052) );
  NAND U8746 ( .A(n59547), .B(n8052), .Z(n8053) );
  AND U8747 ( .A(n59548), .B(n8053), .Z(n59551) );
  AND U8748 ( .A(n59580), .B(n59582), .Z(n8054) );
  NAND U8749 ( .A(n59581), .B(n8054), .Z(n8055) );
  NANDN U8750 ( .A(n59583), .B(n8055), .Z(n8056) );
  AND U8751 ( .A(n59585), .B(n59584), .Z(n8057) );
  NAND U8752 ( .A(n8056), .B(n8057), .Z(n8058) );
  NAND U8753 ( .A(n59586), .B(n8058), .Z(n8059) );
  AND U8754 ( .A(n59587), .B(n59588), .Z(n8060) );
  NAND U8755 ( .A(n8059), .B(n8060), .Z(n8061) );
  NANDN U8756 ( .A(n59589), .B(n8061), .Z(n8062) );
  ANDN U8757 ( .B(n50952), .A(n50951), .Z(n8063) );
  NAND U8758 ( .A(n8062), .B(n8063), .Z(n8064) );
  NAND U8759 ( .A(n59590), .B(n8064), .Z(n8065) );
  ANDN U8760 ( .B(n59591), .A(n59592), .Z(n8066) );
  NAND U8761 ( .A(n8065), .B(n8066), .Z(n8067) );
  NANDN U8762 ( .A(n59593), .B(n8067), .Z(n8068) );
  ANDN U8763 ( .B(n59595), .A(n59594), .Z(n8069) );
  NAND U8764 ( .A(n8068), .B(n8069), .Z(n8070) );
  NANDN U8765 ( .A(n59596), .B(n8070), .Z(n59597) );
  NANDN U8766 ( .A(n50945), .B(n50946), .Z(n59612) );
  AND U8767 ( .A(n59640), .B(n59642), .Z(n8071) );
  NAND U8768 ( .A(n59641), .B(n8071), .Z(n8072) );
  AND U8769 ( .A(n59643), .B(n8072), .Z(n8073) );
  NOR U8770 ( .A(n59645), .B(n8073), .Z(n8074) );
  NAND U8771 ( .A(n59644), .B(n8074), .Z(n8075) );
  ANDN U8772 ( .B(n8075), .A(n59646), .Z(n8076) );
  NOR U8773 ( .A(n8076), .B(n50933), .Z(n8077) );
  NAND U8774 ( .A(n50934), .B(n8077), .Z(n8078) );
  NAND U8775 ( .A(n59647), .B(n8078), .Z(n8079) );
  AND U8776 ( .A(n59649), .B(n59648), .Z(n8080) );
  NAND U8777 ( .A(n8079), .B(n8080), .Z(n8081) );
  NAND U8778 ( .A(n59650), .B(n8081), .Z(n8082) );
  AND U8779 ( .A(n50932), .B(n50931), .Z(n8083) );
  NAND U8780 ( .A(n8082), .B(n8083), .Z(n8084) );
  NAND U8781 ( .A(n59651), .B(n8084), .Z(n8085) );
  AND U8782 ( .A(n59652), .B(n8085), .Z(n8086) );
  NAND U8783 ( .A(n59653), .B(n8086), .Z(n59654) );
  NAND U8784 ( .A(n59686), .B(n59685), .Z(n8087) );
  NANDN U8785 ( .A(n59687), .B(n8087), .Z(n8088) );
  AND U8786 ( .A(n59688), .B(n8088), .Z(n8089) );
  AND U8787 ( .A(n59690), .B(n59691), .Z(n8090) );
  OR U8788 ( .A(n59689), .B(n8089), .Z(n8091) );
  AND U8789 ( .A(n8090), .B(n8091), .Z(n8092) );
  ANDN U8790 ( .B(n50922), .A(n50921), .Z(n8093) );
  NANDN U8791 ( .A(n8092), .B(n59692), .Z(n8094) );
  AND U8792 ( .A(n8093), .B(n8094), .Z(n8095) );
  NOR U8793 ( .A(n59695), .B(n59694), .Z(n8096) );
  OR U8794 ( .A(n59693), .B(n8095), .Z(n8097) );
  AND U8795 ( .A(n8096), .B(n8097), .Z(n8098) );
  ANDN U8796 ( .B(n59697), .A(n59696), .Z(n8099) );
  NANDN U8797 ( .A(n8098), .B(n50920), .Z(n8100) );
  AND U8798 ( .A(n8099), .B(n8100), .Z(n8101) );
  NANDN U8799 ( .A(n8101), .B(n59698), .Z(n8102) );
  AND U8800 ( .A(n59699), .B(n8102), .Z(n59702) );
  AND U8801 ( .A(n59730), .B(n59733), .Z(n8103) );
  NAND U8802 ( .A(n59731), .B(n8103), .Z(n8104) );
  AND U8803 ( .A(n59734), .B(n8104), .Z(n8105) );
  NOR U8804 ( .A(n50910), .B(n8105), .Z(n8106) );
  NAND U8805 ( .A(n50909), .B(n8106), .Z(n8107) );
  AND U8806 ( .A(n59735), .B(n8107), .Z(n8108) );
  NANDN U8807 ( .A(n8108), .B(n59736), .Z(n8109) );
  AND U8808 ( .A(n59737), .B(n8109), .Z(n8110) );
  ANDN U8809 ( .B(n59738), .A(n8110), .Z(n8111) );
  NAND U8810 ( .A(n59739), .B(n8111), .Z(n8112) );
  NANDN U8811 ( .A(n59740), .B(n8112), .Z(n8113) );
  AND U8812 ( .A(n59742), .B(n59741), .Z(n8114) );
  NAND U8813 ( .A(n8113), .B(n8114), .Z(n8115) );
  NAND U8814 ( .A(n59743), .B(n8115), .Z(n8116) );
  ANDN U8815 ( .B(n59745), .A(n59744), .Z(n8117) );
  NAND U8816 ( .A(n8116), .B(n8117), .Z(n8118) );
  NANDN U8817 ( .A(n59746), .B(n8118), .Z(n8119) );
  AND U8818 ( .A(n59747), .B(n8119), .Z(n59749) );
  ANDN U8819 ( .B(n59780), .A(n59779), .Z(n8120) );
  NAND U8820 ( .A(n59778), .B(n59777), .Z(n8121) );
  AND U8821 ( .A(n8120), .B(n8121), .Z(n8122) );
  AND U8822 ( .A(n50899), .B(n50898), .Z(n8123) );
  OR U8823 ( .A(n8122), .B(n59781), .Z(n8124) );
  AND U8824 ( .A(n8123), .B(n8124), .Z(n8125) );
  AND U8825 ( .A(n59784), .B(n59783), .Z(n8126) );
  NANDN U8826 ( .A(n8125), .B(n59782), .Z(n8127) );
  AND U8827 ( .A(n8126), .B(n8127), .Z(n8128) );
  ANDN U8828 ( .B(n50897), .A(n50896), .Z(n8129) );
  OR U8829 ( .A(n59785), .B(n8128), .Z(n8130) );
  AND U8830 ( .A(n8129), .B(n8130), .Z(n8131) );
  ANDN U8831 ( .B(n59788), .A(n59787), .Z(n8132) );
  OR U8832 ( .A(n59786), .B(n8131), .Z(n8133) );
  AND U8833 ( .A(n8132), .B(n8133), .Z(n8134) );
  NANDN U8834 ( .A(n8134), .B(n59789), .Z(n8135) );
  AND U8835 ( .A(n59790), .B(n8135), .Z(n59791) );
  ANDN U8836 ( .B(n50873), .A(n50872), .Z(n8136) );
  NANDN U8837 ( .A(n59865), .B(n59864), .Z(n8137) );
  NAND U8838 ( .A(n8136), .B(n8137), .Z(n8138) );
  NAND U8839 ( .A(n59866), .B(n8138), .Z(n8139) );
  AND U8840 ( .A(n59868), .B(n8139), .Z(n8140) );
  NANDN U8841 ( .A(n59867), .B(n8140), .Z(n8141) );
  NAND U8842 ( .A(n59869), .B(n8141), .Z(n8142) );
  AND U8843 ( .A(n59870), .B(n8142), .Z(n8143) );
  NANDN U8844 ( .A(n59871), .B(n8143), .Z(n8144) );
  NAND U8845 ( .A(n50871), .B(n8144), .Z(n8145) );
  AND U8846 ( .A(n59873), .B(n8145), .Z(n8146) );
  NANDN U8847 ( .A(n59872), .B(n8146), .Z(n8147) );
  NAND U8848 ( .A(n59874), .B(n8147), .Z(n8148) );
  AND U8849 ( .A(n59875), .B(n8148), .Z(n8149) );
  NANDN U8850 ( .A(n50870), .B(n8149), .Z(n59876) );
  ANDN U8851 ( .B(n59909), .A(n59908), .Z(n8150) );
  NANDN U8852 ( .A(n59907), .B(n59906), .Z(n8151) );
  NAND U8853 ( .A(n8150), .B(n8151), .Z(n8152) );
  NAND U8854 ( .A(n59910), .B(n8152), .Z(n8153) );
  AND U8855 ( .A(n59911), .B(n8153), .Z(n8154) );
  NAND U8856 ( .A(n8154), .B(n59912), .Z(n8155) );
  NAND U8857 ( .A(n50862), .B(n8155), .Z(n8156) );
  AND U8858 ( .A(n59913), .B(n8156), .Z(n8157) );
  NAND U8859 ( .A(n8157), .B(n59914), .Z(n8158) );
  ANDN U8860 ( .B(n50861), .A(n50860), .Z(n8159) );
  NANDN U8861 ( .A(n59915), .B(n8158), .Z(n8160) );
  NAND U8862 ( .A(n8159), .B(n8160), .Z(n8161) );
  NAND U8863 ( .A(n59916), .B(n8161), .Z(n8162) );
  AND U8864 ( .A(n59918), .B(n8162), .Z(n8163) );
  NAND U8865 ( .A(n8163), .B(n59917), .Z(n8164) );
  NAND U8866 ( .A(n50859), .B(n8164), .Z(n59919) );
  AND U8867 ( .A(n59950), .B(n59949), .Z(n8165) );
  NAND U8868 ( .A(n59948), .B(n59947), .Z(n8166) );
  AND U8869 ( .A(n8165), .B(n8166), .Z(n8167) );
  AND U8870 ( .A(n59953), .B(n59952), .Z(n8168) );
  NANDN U8871 ( .A(n8167), .B(n59951), .Z(n8169) );
  AND U8872 ( .A(n8168), .B(n8169), .Z(n8170) );
  AND U8873 ( .A(n59954), .B(n59955), .Z(n8171) );
  NANDN U8874 ( .A(n8170), .B(n50847), .Z(n8172) );
  AND U8875 ( .A(n8171), .B(n8172), .Z(n8173) );
  ANDN U8876 ( .B(n59958), .A(n59957), .Z(n8174) );
  NANDN U8877 ( .A(n8173), .B(n59956), .Z(n8175) );
  AND U8878 ( .A(n8174), .B(n8175), .Z(n8176) );
  AND U8879 ( .A(n59960), .B(n59961), .Z(n8177) );
  OR U8880 ( .A(n59959), .B(n8176), .Z(n8178) );
  AND U8881 ( .A(n8177), .B(n8178), .Z(n8179) );
  ANDN U8882 ( .B(n59964), .A(n59963), .Z(n8180) );
  NANDN U8883 ( .A(n8179), .B(n59962), .Z(n8181) );
  AND U8884 ( .A(n8180), .B(n8181), .Z(n59966) );
  ANDN U8885 ( .B(n50835), .A(n50834), .Z(n8182) );
  NANDN U8886 ( .A(n50836), .B(n59993), .Z(n8183) );
  NAND U8887 ( .A(n8182), .B(n8183), .Z(n8184) );
  NAND U8888 ( .A(n59994), .B(n8184), .Z(n8185) );
  AND U8889 ( .A(n59996), .B(n8185), .Z(n8186) );
  NANDN U8890 ( .A(n59995), .B(n8186), .Z(n8187) );
  NAND U8891 ( .A(n59997), .B(n8187), .Z(n8188) );
  AND U8892 ( .A(n50833), .B(n8188), .Z(n8189) );
  NANDN U8893 ( .A(n50832), .B(n8189), .Z(n8190) );
  NAND U8894 ( .A(n59998), .B(n8190), .Z(n8191) );
  AND U8895 ( .A(n60000), .B(n8191), .Z(n8192) );
  NANDN U8896 ( .A(n59999), .B(n8192), .Z(n8193) );
  AND U8897 ( .A(n50831), .B(n50830), .Z(n8194) );
  NANDN U8898 ( .A(n60001), .B(n8193), .Z(n8195) );
  NAND U8899 ( .A(n8194), .B(n8195), .Z(n60002) );
  NANDN U8900 ( .A(n50891), .B(n20020), .Z(n8196) );
  NANDN U8901 ( .A(n59804), .B(n8196), .Z(n8197) );
  NAND U8902 ( .A(n22737), .B(n8197), .Z(n8198) );
  NANDN U8903 ( .A(n8198), .B(n59806), .Z(n8199) );
  NAND U8904 ( .A(n59807), .B(n8199), .Z(n8200) );
  NAND U8905 ( .A(n50889), .B(n8200), .Z(n8201) );
  ANDN U8906 ( .B(n59810), .A(n47569), .Z(n8202) );
  NANDN U8907 ( .A(n59808), .B(n8201), .Z(n8203) );
  NAND U8908 ( .A(n8202), .B(n8203), .Z(n8204) );
  NAND U8909 ( .A(n59811), .B(n8204), .Z(n8205) );
  AND U8910 ( .A(n59812), .B(n8205), .Z(n8206) );
  NAND U8911 ( .A(n8206), .B(n22731), .Z(n8207) );
  AND U8912 ( .A(n59815), .B(n22729), .Z(n8208) );
  NANDN U8913 ( .A(n59814), .B(n8207), .Z(n8209) );
  NAND U8914 ( .A(n8208), .B(n8209), .Z(n8210) );
  NAND U8915 ( .A(n59817), .B(n8210), .Z(n8211) );
  AND U8916 ( .A(n50887), .B(n8211), .Z(n8212) );
  NAND U8917 ( .A(n8212), .B(n22727), .Z(n8213) );
  NANDN U8918 ( .A(n59818), .B(n8213), .Z(n20023) );
  AND U8919 ( .A(n60033), .B(n60032), .Z(n8214) );
  NANDN U8920 ( .A(n60031), .B(n60030), .Z(n8215) );
  AND U8921 ( .A(n8214), .B(n8215), .Z(n8216) );
  AND U8922 ( .A(n60036), .B(n60035), .Z(n8217) );
  NANDN U8923 ( .A(n8216), .B(n60034), .Z(n8218) );
  AND U8924 ( .A(n8217), .B(n8218), .Z(n8219) );
  ANDN U8925 ( .B(n50819), .A(n50818), .Z(n8220) );
  NANDN U8926 ( .A(n8219), .B(n60037), .Z(n8221) );
  AND U8927 ( .A(n8220), .B(n8221), .Z(n8222) );
  ANDN U8928 ( .B(n60039), .A(n60040), .Z(n8223) );
  NANDN U8929 ( .A(n8222), .B(n60038), .Z(n8224) );
  AND U8930 ( .A(n8223), .B(n8224), .Z(n8225) );
  OR U8931 ( .A(n60041), .B(n8225), .Z(n8226) );
  NAND U8932 ( .A(n60042), .B(n8226), .Z(n8227) );
  NAND U8933 ( .A(n60043), .B(n8227), .Z(n8228) );
  NAND U8934 ( .A(n60044), .B(n8228), .Z(n8229) );
  NAND U8935 ( .A(n60045), .B(n8229), .Z(n8230) );
  ANDN U8936 ( .B(n8230), .A(n60046), .Z(n60048) );
  NAND U8937 ( .A(n60075), .B(n60076), .Z(n8231) );
  NOR U8938 ( .A(n50809), .B(n50810), .Z(n8232) );
  NANDN U8939 ( .A(n60077), .B(n8231), .Z(n8233) );
  NAND U8940 ( .A(n8232), .B(n8233), .Z(n8234) );
  NAND U8941 ( .A(n60078), .B(n8234), .Z(n8235) );
  AND U8942 ( .A(n60080), .B(n8235), .Z(n8236) );
  NANDN U8943 ( .A(n60079), .B(n8236), .Z(n8237) );
  ANDN U8944 ( .B(n50808), .A(n50807), .Z(n8238) );
  NANDN U8945 ( .A(n60081), .B(n8237), .Z(n8239) );
  NAND U8946 ( .A(n8238), .B(n8239), .Z(n8240) );
  NAND U8947 ( .A(n50806), .B(n8240), .Z(n8241) );
  AND U8948 ( .A(n60083), .B(n8241), .Z(n8242) );
  NANDN U8949 ( .A(n60082), .B(n8242), .Z(n8243) );
  NAND U8950 ( .A(n60084), .B(n8243), .Z(n8244) );
  AND U8951 ( .A(n60085), .B(n8244), .Z(n8245) );
  NANDN U8952 ( .A(n50805), .B(n8245), .Z(n60086) );
  NAND U8953 ( .A(n60114), .B(n60113), .Z(n8246) );
  AND U8954 ( .A(n60115), .B(n8246), .Z(n8247) );
  NOR U8955 ( .A(n60116), .B(n8247), .Z(n8248) );
  NAND U8956 ( .A(n60117), .B(n8248), .Z(n8249) );
  NANDN U8957 ( .A(n60118), .B(n8249), .Z(n8250) );
  ANDN U8958 ( .B(n60120), .A(n60119), .Z(n8251) );
  NAND U8959 ( .A(n8250), .B(n8251), .Z(n8252) );
  NAND U8960 ( .A(n60121), .B(n8252), .Z(n8253) );
  ANDN U8961 ( .B(n60123), .A(n60122), .Z(n8254) );
  NAND U8962 ( .A(n8253), .B(n8254), .Z(n8255) );
  NAND U8963 ( .A(n60124), .B(n8255), .Z(n8256) );
  ANDN U8964 ( .B(n60125), .A(n60126), .Z(n8257) );
  NAND U8965 ( .A(n8256), .B(n8257), .Z(n8258) );
  NANDN U8966 ( .A(n60127), .B(n8258), .Z(n8259) );
  NAND U8967 ( .A(n60128), .B(n8259), .Z(n8260) );
  NAND U8968 ( .A(n60129), .B(n8260), .Z(n8261) );
  AND U8969 ( .A(n60130), .B(n8261), .Z(n60132) );
  NAND U8970 ( .A(n60163), .B(n60162), .Z(n8262) );
  AND U8971 ( .A(n60164), .B(n8262), .Z(n8263) );
  NOR U8972 ( .A(n8263), .B(n50785), .Z(n8264) );
  NAND U8973 ( .A(n50784), .B(n8264), .Z(n8265) );
  AND U8974 ( .A(n60165), .B(n8265), .Z(n8266) );
  NOR U8975 ( .A(n60166), .B(n8266), .Z(n8267) );
  NAND U8976 ( .A(n50783), .B(n8267), .Z(n8268) );
  AND U8977 ( .A(n60167), .B(n8268), .Z(n8269) );
  NANDN U8978 ( .A(n8269), .B(n50782), .Z(n8270) );
  NAND U8979 ( .A(n60168), .B(n8270), .Z(n8271) );
  NAND U8980 ( .A(n60169), .B(n8271), .Z(n8272) );
  ANDN U8981 ( .B(n50781), .A(n50780), .Z(n8273) );
  NANDN U8982 ( .A(n60170), .B(n8272), .Z(n8274) );
  NAND U8983 ( .A(n8273), .B(n8274), .Z(n8275) );
  NAND U8984 ( .A(n60171), .B(n8275), .Z(n60172) );
  NAND U8985 ( .A(n20226), .B(n20225), .Z(n8276) );
  AND U8986 ( .A(n59981), .B(n8276), .Z(n8277) );
  ANDN U8987 ( .B(n59982), .A(n8277), .Z(n8278) );
  NAND U8988 ( .A(n47898), .B(n8278), .Z(n8279) );
  NANDN U8989 ( .A(n50841), .B(n8279), .Z(n8280) );
  AND U8990 ( .A(n22643), .B(n22642), .Z(n8281) );
  NAND U8991 ( .A(n8280), .B(n8281), .Z(n8282) );
  NAND U8992 ( .A(n59986), .B(n8282), .Z(n8283) );
  AND U8993 ( .A(n47908), .B(n59987), .Z(n8284) );
  NAND U8994 ( .A(n8283), .B(n8284), .Z(n8285) );
  NAND U8995 ( .A(n59989), .B(n8285), .Z(n8286) );
  ANDN U8996 ( .B(n8286), .A(n50839), .Z(n8287) );
  XNOR U8997 ( .A(y[7142]), .B(x[7142]), .Z(n8288) );
  AND U8998 ( .A(n8287), .B(n8288), .Z(n8289) );
  OR U8999 ( .A(n59990), .B(n8289), .Z(n8290) );
  AND U9000 ( .A(n59991), .B(n8290), .Z(n8291) );
  AND U9001 ( .A(n50837), .B(n22634), .Z(n8292) );
  NANDN U9002 ( .A(n8291), .B(n59992), .Z(n8293) );
  AND U9003 ( .A(n8292), .B(n8293), .Z(n20229) );
  ANDN U9004 ( .B(n60202), .A(n60201), .Z(n8294) );
  NAND U9005 ( .A(n60203), .B(n8294), .Z(n8295) );
  NAND U9006 ( .A(n60204), .B(n8295), .Z(n8296) );
  AND U9007 ( .A(n60206), .B(n60205), .Z(n8297) );
  NAND U9008 ( .A(n8296), .B(n8297), .Z(n8298) );
  NAND U9009 ( .A(n60207), .B(n8298), .Z(n8299) );
  ANDN U9010 ( .B(n50770), .A(n50769), .Z(n8300) );
  NAND U9011 ( .A(n8299), .B(n8300), .Z(n8301) );
  NAND U9012 ( .A(n60208), .B(n8301), .Z(n8302) );
  ANDN U9013 ( .B(n60209), .A(n60210), .Z(n8303) );
  NAND U9014 ( .A(n8302), .B(n8303), .Z(n8304) );
  NAND U9015 ( .A(n60211), .B(n8304), .Z(n8305) );
  ANDN U9016 ( .B(n50768), .A(n50767), .Z(n8306) );
  NAND U9017 ( .A(n8305), .B(n8306), .Z(n8307) );
  NAND U9018 ( .A(n50766), .B(n8307), .Z(n8308) );
  AND U9019 ( .A(n60213), .B(n60212), .Z(n8309) );
  NAND U9020 ( .A(n8308), .B(n8309), .Z(n8310) );
  NAND U9021 ( .A(n60214), .B(n8310), .Z(n60216) );
  AND U9022 ( .A(n60245), .B(n60244), .Z(n8311) );
  NAND U9023 ( .A(n60242), .B(n60243), .Z(n8312) );
  AND U9024 ( .A(n8311), .B(n8312), .Z(n8313) );
  AND U9025 ( .A(n60248), .B(n60247), .Z(n8314) );
  OR U9026 ( .A(n60246), .B(n8313), .Z(n8315) );
  AND U9027 ( .A(n8314), .B(n8315), .Z(n8316) );
  OR U9028 ( .A(n50759), .B(n8316), .Z(n8317) );
  NAND U9029 ( .A(n60249), .B(n8317), .Z(n8318) );
  NAND U9030 ( .A(n60250), .B(n8318), .Z(n8319) );
  ANDN U9031 ( .B(n60252), .A(n60251), .Z(n8320) );
  NAND U9032 ( .A(n8319), .B(n8320), .Z(n8321) );
  NANDN U9033 ( .A(n60253), .B(n8321), .Z(n8322) );
  ANDN U9034 ( .B(n50758), .A(n50757), .Z(n8323) );
  NAND U9035 ( .A(n8322), .B(n8323), .Z(n8324) );
  NAND U9036 ( .A(n60254), .B(n8324), .Z(n8325) );
  ANDN U9037 ( .B(n8325), .A(n60255), .Z(n60257) );
  AND U9038 ( .A(n60280), .B(n50743), .Z(n8326) );
  NANDN U9039 ( .A(n50744), .B(n60279), .Z(n8327) );
  AND U9040 ( .A(n8326), .B(n8327), .Z(n8328) );
  NANDN U9041 ( .A(n8328), .B(n60281), .Z(n8329) );
  NAND U9042 ( .A(n60282), .B(n8329), .Z(n8330) );
  NAND U9043 ( .A(n60283), .B(n8330), .Z(n8331) );
  AND U9044 ( .A(n60284), .B(n60285), .Z(n8332) );
  NAND U9045 ( .A(n8331), .B(n8332), .Z(n8333) );
  NAND U9046 ( .A(n50742), .B(n8333), .Z(n8334) );
  AND U9047 ( .A(n60287), .B(n60286), .Z(n8335) );
  NAND U9048 ( .A(n8334), .B(n8335), .Z(n8336) );
  NAND U9049 ( .A(n60288), .B(n8336), .Z(n8337) );
  ANDN U9050 ( .B(n60290), .A(n60289), .Z(n8338) );
  NAND U9051 ( .A(n8337), .B(n8338), .Z(n8339) );
  NANDN U9052 ( .A(n60291), .B(n8339), .Z(n60292) );
  NOR U9053 ( .A(n60322), .B(n60323), .Z(n8340) );
  AND U9054 ( .A(n50732), .B(n50733), .Z(n8341) );
  NANDN U9055 ( .A(n8340), .B(n60324), .Z(n8342) );
  AND U9056 ( .A(n8341), .B(n8342), .Z(n8343) );
  AND U9057 ( .A(n60326), .B(n60327), .Z(n8344) );
  NANDN U9058 ( .A(n8343), .B(n60325), .Z(n8345) );
  AND U9059 ( .A(n8344), .B(n8345), .Z(n8346) );
  ANDN U9060 ( .B(n50731), .A(n50730), .Z(n8347) );
  OR U9061 ( .A(n8346), .B(n60328), .Z(n8348) );
  AND U9062 ( .A(n8347), .B(n8348), .Z(n8349) );
  ANDN U9063 ( .B(n60331), .A(n60330), .Z(n8350) );
  OR U9064 ( .A(n60329), .B(n8349), .Z(n8351) );
  AND U9065 ( .A(n8350), .B(n8351), .Z(n8352) );
  AND U9066 ( .A(n60334), .B(n60333), .Z(n8353) );
  NANDN U9067 ( .A(n8352), .B(n60332), .Z(n8354) );
  AND U9068 ( .A(n8353), .B(n8354), .Z(n8355) );
  AND U9069 ( .A(n60336), .B(n60337), .Z(n8356) );
  OR U9070 ( .A(n8355), .B(n60335), .Z(n8357) );
  NAND U9071 ( .A(n8356), .B(n8357), .Z(n60338) );
  NAND U9072 ( .A(n60368), .B(n60369), .Z(n8358) );
  NAND U9073 ( .A(n60370), .B(n8358), .Z(n8359) );
  AND U9074 ( .A(n60371), .B(n8359), .Z(n8360) );
  NAND U9075 ( .A(n8360), .B(n60372), .Z(n8361) );
  NAND U9076 ( .A(n60373), .B(n8361), .Z(n8362) );
  ANDN U9077 ( .B(n8362), .A(n50722), .Z(n8363) );
  NANDN U9078 ( .A(n8363), .B(n60374), .Z(n8364) );
  AND U9079 ( .A(n60375), .B(n8364), .Z(n8365) );
  AND U9080 ( .A(n60378), .B(n60377), .Z(n8366) );
  NANDN U9081 ( .A(n8365), .B(n60376), .Z(n8367) );
  AND U9082 ( .A(n8366), .B(n8367), .Z(n8368) );
  NOR U9083 ( .A(n50720), .B(n50721), .Z(n8369) );
  OR U9084 ( .A(n8368), .B(n60379), .Z(n8370) );
  AND U9085 ( .A(n8369), .B(n8370), .Z(n8371) );
  ANDN U9086 ( .B(n60382), .A(n60381), .Z(n8372) );
  NANDN U9087 ( .A(n8371), .B(n60380), .Z(n8373) );
  AND U9088 ( .A(n8372), .B(n8373), .Z(n60383) );
  NOR U9089 ( .A(n60419), .B(n60418), .Z(n8374) );
  ANDN U9090 ( .B(n50709), .A(n50708), .Z(n8375) );
  NAND U9091 ( .A(n60407), .B(n8375), .Z(n8376) );
  NAND U9092 ( .A(n50707), .B(n8376), .Z(n8377) );
  AND U9093 ( .A(n60409), .B(n60408), .Z(n8378) );
  NAND U9094 ( .A(n8377), .B(n8378), .Z(n8379) );
  NAND U9095 ( .A(n60410), .B(n8379), .Z(n8380) );
  ANDN U9096 ( .B(n60412), .A(n60411), .Z(n8381) );
  NAND U9097 ( .A(n8380), .B(n8381), .Z(n8382) );
  NAND U9098 ( .A(n60413), .B(n8382), .Z(n8383) );
  ANDN U9099 ( .B(n60414), .A(n60415), .Z(n8384) );
  NAND U9100 ( .A(n8383), .B(n8384), .Z(n8385) );
  NANDN U9101 ( .A(n60416), .B(n8385), .Z(n8386) );
  ANDN U9102 ( .B(n50706), .A(n50705), .Z(n8387) );
  NAND U9103 ( .A(n8386), .B(n8387), .Z(n8388) );
  NANDN U9104 ( .A(n60417), .B(n8388), .Z(n8389) );
  NAND U9105 ( .A(n8374), .B(n8389), .Z(n60420) );
  AND U9106 ( .A(n60449), .B(n60450), .Z(n8390) );
  NAND U9107 ( .A(n60451), .B(n8390), .Z(n8391) );
  NAND U9108 ( .A(n50697), .B(n8391), .Z(n8392) );
  ANDN U9109 ( .B(n60453), .A(n60452), .Z(n8393) );
  NAND U9110 ( .A(n8392), .B(n8393), .Z(n8394) );
  NAND U9111 ( .A(n60454), .B(n8394), .Z(n8395) );
  AND U9112 ( .A(n60455), .B(n60456), .Z(n8396) );
  NAND U9113 ( .A(n8395), .B(n8396), .Z(n8397) );
  NANDN U9114 ( .A(n60457), .B(n8397), .Z(n8398) );
  ANDN U9115 ( .B(n50696), .A(n50695), .Z(n8399) );
  NAND U9116 ( .A(n8398), .B(n8399), .Z(n8400) );
  NAND U9117 ( .A(n60458), .B(n8400), .Z(n8401) );
  ANDN U9118 ( .B(n60459), .A(n60460), .Z(n8402) );
  NAND U9119 ( .A(n8401), .B(n8402), .Z(n8403) );
  NAND U9120 ( .A(n60461), .B(n8403), .Z(n60462) );
  ANDN U9121 ( .B(n60495), .A(n60496), .Z(n8404) );
  NAND U9122 ( .A(n60494), .B(n8404), .Z(n8405) );
  NANDN U9123 ( .A(n60497), .B(n8405), .Z(n8406) );
  AND U9124 ( .A(n60498), .B(n60499), .Z(n8407) );
  NAND U9125 ( .A(n8406), .B(n8407), .Z(n8408) );
  NANDN U9126 ( .A(n60500), .B(n8408), .Z(n8409) );
  NAND U9127 ( .A(n60501), .B(n8409), .Z(n8410) );
  NANDN U9128 ( .A(n50686), .B(n8410), .Z(n8411) );
  AND U9129 ( .A(n50685), .B(n8411), .Z(n8412) );
  NAND U9130 ( .A(n60502), .B(n8412), .Z(n8413) );
  NAND U9131 ( .A(n60503), .B(n8413), .Z(n8414) );
  NANDN U9132 ( .A(n60504), .B(n8414), .Z(n8415) );
  OR U9133 ( .A(n8415), .B(n60505), .Z(n8416) );
  NANDN U9134 ( .A(n60506), .B(n8416), .Z(n8417) );
  NAND U9135 ( .A(n60507), .B(n8417), .Z(n8418) );
  NANDN U9136 ( .A(n60508), .B(n8418), .Z(n60509) );
  NAND U9137 ( .A(n60536), .B(n60535), .Z(n8419) );
  NANDN U9138 ( .A(n60537), .B(n8419), .Z(n8420) );
  ANDN U9139 ( .B(n8420), .A(n60538), .Z(n8421) );
  NAND U9140 ( .A(n8421), .B(n60539), .Z(n8422) );
  NAND U9141 ( .A(n60540), .B(n8422), .Z(n8423) );
  AND U9142 ( .A(n60541), .B(n8423), .Z(n8424) );
  NANDN U9143 ( .A(n50673), .B(n8424), .Z(n8425) );
  NANDN U9144 ( .A(n60542), .B(n8425), .Z(n8426) );
  ANDN U9145 ( .B(n8426), .A(n60543), .Z(n8427) );
  NAND U9146 ( .A(n8427), .B(n60544), .Z(n8428) );
  NAND U9147 ( .A(n60545), .B(n8428), .Z(n8429) );
  AND U9148 ( .A(n60546), .B(n8429), .Z(n8430) );
  AND U9149 ( .A(n60547), .B(n8430), .Z(n8431) );
  ANDN U9150 ( .B(n50672), .A(n50671), .Z(n8432) );
  NANDN U9151 ( .A(n8431), .B(n60548), .Z(n8433) );
  AND U9152 ( .A(n8432), .B(n8433), .Z(n8434) );
  AND U9153 ( .A(n60550), .B(n60551), .Z(n8435) );
  NANDN U9154 ( .A(n8434), .B(n60549), .Z(n8436) );
  AND U9155 ( .A(n8435), .B(n8436), .Z(n60553) );
  NAND U9156 ( .A(n60574), .B(n60573), .Z(n8437) );
  AND U9157 ( .A(n60575), .B(n8437), .Z(n8438) );
  NOR U9158 ( .A(n60576), .B(n8438), .Z(n8439) );
  NAND U9159 ( .A(n60577), .B(n8439), .Z(n8440) );
  NANDN U9160 ( .A(n60578), .B(n8440), .Z(n8441) );
  NOR U9161 ( .A(n60580), .B(n60579), .Z(n8442) );
  NAND U9162 ( .A(n8441), .B(n8442), .Z(n8443) );
  NAND U9163 ( .A(n50654), .B(n8443), .Z(n8444) );
  ANDN U9164 ( .B(n60582), .A(n60581), .Z(n8445) );
  NAND U9165 ( .A(n8444), .B(n8445), .Z(n8446) );
  NAND U9166 ( .A(n60583), .B(n8446), .Z(n8447) );
  ANDN U9167 ( .B(n50653), .A(n50652), .Z(n8448) );
  NAND U9168 ( .A(n8447), .B(n8448), .Z(n8449) );
  NAND U9169 ( .A(n60584), .B(n8449), .Z(n8450) );
  ANDN U9170 ( .B(n8450), .A(n60585), .Z(n60587) );
  XNOR U9171 ( .A(x[7582]), .B(y[7582]), .Z(n20909) );
  AND U9172 ( .A(n60618), .B(n60619), .Z(n8451) );
  AND U9173 ( .A(n50643), .B(n50642), .Z(n8452) );
  OR U9174 ( .A(n60620), .B(n8451), .Z(n8453) );
  AND U9175 ( .A(n8452), .B(n8453), .Z(n8454) );
  ANDN U9176 ( .B(n60622), .A(n60623), .Z(n8455) );
  NANDN U9177 ( .A(n8454), .B(n60621), .Z(n8456) );
  AND U9178 ( .A(n8455), .B(n8456), .Z(n8457) );
  ANDN U9179 ( .B(n50641), .A(n50640), .Z(n8458) );
  OR U9180 ( .A(n60624), .B(n8457), .Z(n8459) );
  AND U9181 ( .A(n8458), .B(n8459), .Z(n8460) );
  NANDN U9182 ( .A(n8460), .B(n50639), .Z(n8461) );
  NAND U9183 ( .A(n60625), .B(n8461), .Z(n8462) );
  NANDN U9184 ( .A(n60626), .B(n8462), .Z(n8463) );
  AND U9185 ( .A(n50638), .B(n50637), .Z(n8464) );
  NAND U9186 ( .A(n8463), .B(n8464), .Z(n8465) );
  NANDN U9187 ( .A(n50636), .B(n8465), .Z(n60627) );
  NOR U9188 ( .A(n50625), .B(n50626), .Z(n8466) );
  NAND U9189 ( .A(n60657), .B(n8466), .Z(n8467) );
  NAND U9190 ( .A(n60658), .B(n8467), .Z(n8468) );
  ANDN U9191 ( .B(n60660), .A(n60659), .Z(n8469) );
  NAND U9192 ( .A(n8468), .B(n8469), .Z(n8470) );
  NAND U9193 ( .A(n60661), .B(n8470), .Z(n8471) );
  AND U9194 ( .A(n50623), .B(n50622), .Z(n8472) );
  NAND U9195 ( .A(n8471), .B(n8472), .Z(n8473) );
  NANDN U9196 ( .A(n60662), .B(n8473), .Z(n8474) );
  AND U9197 ( .A(n60664), .B(n60663), .Z(n8475) );
  NAND U9198 ( .A(n8474), .B(n8475), .Z(n8476) );
  NAND U9199 ( .A(n60665), .B(n8476), .Z(n8477) );
  ANDN U9200 ( .B(n60666), .A(n50621), .Z(n8478) );
  NAND U9201 ( .A(n8477), .B(n8478), .Z(n8479) );
  NANDN U9202 ( .A(n60667), .B(n8479), .Z(n8480) );
  ANDN U9203 ( .B(n60669), .A(n60668), .Z(n8481) );
  NAND U9204 ( .A(n8480), .B(n8481), .Z(n8482) );
  NAND U9205 ( .A(n60670), .B(n8482), .Z(n8483) );
  AND U9206 ( .A(n60671), .B(n8483), .Z(n60673) );
  NANDN U9207 ( .A(n50611), .B(n60720), .Z(n8484) );
  ANDN U9208 ( .B(n8484), .A(n60721), .Z(n8485) );
  NOR U9209 ( .A(n60722), .B(n8485), .Z(n8486) );
  NAND U9210 ( .A(n60723), .B(n8486), .Z(n8487) );
  NAND U9211 ( .A(n60724), .B(n8487), .Z(n8488) );
  AND U9212 ( .A(n60726), .B(n60725), .Z(n8489) );
  NAND U9213 ( .A(n8488), .B(n8489), .Z(n8490) );
  NAND U9214 ( .A(n60727), .B(n8490), .Z(n8491) );
  ANDN U9215 ( .B(n50610), .A(n50609), .Z(n8492) );
  NAND U9216 ( .A(n8491), .B(n8492), .Z(n8493) );
  NAND U9217 ( .A(n60728), .B(n8493), .Z(n8494) );
  ANDN U9218 ( .B(n60729), .A(n60730), .Z(n8495) );
  NAND U9219 ( .A(n8494), .B(n8495), .Z(n8496) );
  NAND U9220 ( .A(n60731), .B(n8496), .Z(n8497) );
  ANDN U9221 ( .B(n50608), .A(n50607), .Z(n8498) );
  NAND U9222 ( .A(n8497), .B(n8498), .Z(n8499) );
  NAND U9223 ( .A(n50606), .B(n8499), .Z(n60733) );
  ANDN U9224 ( .B(n60759), .A(n60761), .Z(n8500) );
  NAND U9225 ( .A(n60760), .B(n8500), .Z(n8501) );
  NAND U9226 ( .A(n60762), .B(n8501), .Z(n8502) );
  ANDN U9227 ( .B(n50597), .A(n50596), .Z(n8503) );
  NAND U9228 ( .A(n8502), .B(n8503), .Z(n8504) );
  NAND U9229 ( .A(n60763), .B(n8504), .Z(n8505) );
  AND U9230 ( .A(n50595), .B(n50594), .Z(n8506) );
  NAND U9231 ( .A(n8505), .B(n8506), .Z(n8507) );
  NAND U9232 ( .A(n60764), .B(n8507), .Z(n8508) );
  ANDN U9233 ( .B(n60766), .A(n60765), .Z(n8509) );
  NAND U9234 ( .A(n8508), .B(n8509), .Z(n8510) );
  NANDN U9235 ( .A(n60767), .B(n8510), .Z(n8511) );
  ANDN U9236 ( .B(n50593), .A(n50592), .Z(n8512) );
  NAND U9237 ( .A(n8511), .B(n8512), .Z(n8513) );
  NANDN U9238 ( .A(n60768), .B(n8513), .Z(n8514) );
  ANDN U9239 ( .B(n8514), .A(n60769), .Z(n60771) );
  AND U9240 ( .A(n60785), .B(n60784), .Z(n60786) );
  AND U9241 ( .A(n60840), .B(n60839), .Z(n8515) );
  NAND U9242 ( .A(n60836), .B(n60837), .Z(n8516) );
  AND U9243 ( .A(n8515), .B(n8516), .Z(n8517) );
  ANDN U9244 ( .B(n50577), .A(n50576), .Z(n8518) );
  OR U9245 ( .A(n60841), .B(n8517), .Z(n8519) );
  AND U9246 ( .A(n8518), .B(n8519), .Z(n8520) );
  AND U9247 ( .A(n60843), .B(n60844), .Z(n8521) );
  OR U9248 ( .A(n60842), .B(n8520), .Z(n8522) );
  AND U9249 ( .A(n8521), .B(n8522), .Z(n8523) );
  AND U9250 ( .A(n60847), .B(n60846), .Z(n8524) );
  NANDN U9251 ( .A(n8523), .B(n60845), .Z(n8525) );
  AND U9252 ( .A(n8524), .B(n8525), .Z(n8526) );
  NOR U9253 ( .A(n50575), .B(n50574), .Z(n8527) );
  OR U9254 ( .A(n60848), .B(n8526), .Z(n8528) );
  AND U9255 ( .A(n8527), .B(n8528), .Z(n8529) );
  NOR U9256 ( .A(n60850), .B(n60851), .Z(n8530) );
  NANDN U9257 ( .A(n8529), .B(n60849), .Z(n8531) );
  AND U9258 ( .A(n8530), .B(n8531), .Z(n60854) );
  NANDN U9259 ( .A(n60884), .B(n60883), .Z(n8532) );
  NAND U9260 ( .A(n60885), .B(n8532), .Z(n8533) );
  AND U9261 ( .A(n60886), .B(n8533), .Z(n8534) );
  ANDN U9262 ( .B(n50564), .A(n8534), .Z(n8535) );
  NAND U9263 ( .A(n50565), .B(n8535), .Z(n8536) );
  AND U9264 ( .A(n60887), .B(n8536), .Z(n8537) );
  OR U9265 ( .A(n50563), .B(n8537), .Z(n8538) );
  NAND U9266 ( .A(n60888), .B(n8538), .Z(n8539) );
  NAND U9267 ( .A(n60889), .B(n8539), .Z(n8540) );
  OR U9268 ( .A(n8540), .B(n60890), .Z(n8541) );
  NANDN U9269 ( .A(n60891), .B(n8541), .Z(n8542) );
  NAND U9270 ( .A(n60892), .B(n8542), .Z(n8543) );
  NAND U9271 ( .A(n60893), .B(n8543), .Z(n8544) );
  AND U9272 ( .A(n60894), .B(n8544), .Z(n8545) );
  NAND U9273 ( .A(n8545), .B(n60895), .Z(n8546) );
  NAND U9274 ( .A(n60896), .B(n8546), .Z(n60897) );
  ANDN U9275 ( .B(n50553), .A(n50552), .Z(n8547) );
  OR U9276 ( .A(n60925), .B(n60926), .Z(n8548) );
  NAND U9277 ( .A(n8547), .B(n8548), .Z(n8549) );
  ANDN U9278 ( .B(n60929), .A(n60928), .Z(n8550) );
  NANDN U9279 ( .A(n60927), .B(n8549), .Z(n8551) );
  NAND U9280 ( .A(n8550), .B(n8551), .Z(n8552) );
  NAND U9281 ( .A(n60930), .B(n8552), .Z(n8553) );
  AND U9282 ( .A(n60931), .B(n8553), .Z(n8554) );
  NANDN U9283 ( .A(n50551), .B(n8554), .Z(n8555) );
  NAND U9284 ( .A(n50550), .B(n8555), .Z(n8556) );
  AND U9285 ( .A(n60933), .B(n8556), .Z(n8557) );
  NANDN U9286 ( .A(n60932), .B(n8557), .Z(n8558) );
  NAND U9287 ( .A(n60934), .B(n8558), .Z(n8559) );
  AND U9288 ( .A(n60936), .B(n8559), .Z(n8560) );
  NAND U9289 ( .A(n8560), .B(n60935), .Z(n8561) );
  NANDN U9290 ( .A(n60937), .B(n8561), .Z(n60938) );
  ANDN U9291 ( .B(n60964), .A(n50539), .Z(n8562) );
  NAND U9292 ( .A(n60965), .B(n8562), .Z(n8563) );
  NANDN U9293 ( .A(n60966), .B(n8563), .Z(n8564) );
  ANDN U9294 ( .B(n60968), .A(n60967), .Z(n8565) );
  NAND U9295 ( .A(n8564), .B(n8565), .Z(n8566) );
  NAND U9296 ( .A(n60969), .B(n8566), .Z(n8567) );
  AND U9297 ( .A(n60971), .B(n60970), .Z(n8568) );
  NAND U9298 ( .A(n8567), .B(n8568), .Z(n8569) );
  NAND U9299 ( .A(n60972), .B(n8569), .Z(n8570) );
  ANDN U9300 ( .B(n50538), .A(n50537), .Z(n8571) );
  NAND U9301 ( .A(n8570), .B(n8571), .Z(n8572) );
  NAND U9302 ( .A(n60973), .B(n8572), .Z(n8573) );
  AND U9303 ( .A(n60975), .B(n60974), .Z(n8574) );
  NAND U9304 ( .A(n8573), .B(n8574), .Z(n8575) );
  NAND U9305 ( .A(n60976), .B(n8575), .Z(n8576) );
  AND U9306 ( .A(n50536), .B(n50535), .Z(n8577) );
  NAND U9307 ( .A(n8576), .B(n8577), .Z(n8578) );
  NAND U9308 ( .A(n50534), .B(n8578), .Z(n60978) );
  NAND U9309 ( .A(n61007), .B(n61006), .Z(n8579) );
  NAND U9310 ( .A(n61008), .B(n8579), .Z(n8580) );
  ANDN U9311 ( .B(n8580), .A(n61009), .Z(n8581) );
  NAND U9312 ( .A(n8581), .B(n61010), .Z(n8582) );
  NANDN U9313 ( .A(n61011), .B(n8582), .Z(n8583) );
  AND U9314 ( .A(n61012), .B(n8583), .Z(n8584) );
  NAND U9315 ( .A(n8584), .B(n61013), .Z(n8585) );
  NAND U9316 ( .A(n61014), .B(n8585), .Z(n8586) );
  ANDN U9317 ( .B(n8586), .A(n61015), .Z(n8587) );
  NAND U9318 ( .A(n61016), .B(n8587), .Z(n8588) );
  NAND U9319 ( .A(n61017), .B(n8588), .Z(n8589) );
  AND U9320 ( .A(n50524), .B(n8589), .Z(n8590) );
  NAND U9321 ( .A(n8590), .B(n50525), .Z(n8591) );
  NAND U9322 ( .A(n61018), .B(n8591), .Z(n8592) );
  AND U9323 ( .A(n61020), .B(n8592), .Z(n8593) );
  NAND U9324 ( .A(n8593), .B(n61019), .Z(n8594) );
  NAND U9325 ( .A(n61021), .B(n8594), .Z(n8595) );
  AND U9326 ( .A(n50522), .B(n8595), .Z(n8596) );
  NAND U9327 ( .A(n8596), .B(n50523), .Z(n61022) );
  NAND U9328 ( .A(n61055), .B(n61054), .Z(n8597) );
  NAND U9329 ( .A(n61056), .B(n8597), .Z(n8598) );
  ANDN U9330 ( .B(n8598), .A(n61057), .Z(n8599) );
  NAND U9331 ( .A(n61058), .B(n8599), .Z(n8600) );
  NAND U9332 ( .A(n61059), .B(n8600), .Z(n8601) );
  AND U9333 ( .A(n50513), .B(n8601), .Z(n8602) );
  NANDN U9334 ( .A(n50512), .B(n8602), .Z(n8603) );
  ANDN U9335 ( .B(n61062), .A(n61061), .Z(n8604) );
  NANDN U9336 ( .A(n61060), .B(n8603), .Z(n8605) );
  NAND U9337 ( .A(n8604), .B(n8605), .Z(n8606) );
  NAND U9338 ( .A(n61063), .B(n8606), .Z(n8607) );
  AND U9339 ( .A(n61064), .B(n8607), .Z(n8608) );
  NAND U9340 ( .A(n8608), .B(n61065), .Z(n8609) );
  NAND U9341 ( .A(n50511), .B(n8609), .Z(n8610) );
  AND U9342 ( .A(n61067), .B(n8610), .Z(n8611) );
  NANDN U9343 ( .A(n61066), .B(n8611), .Z(n61068) );
  ANDN U9344 ( .B(n61096), .A(n61095), .Z(n8612) );
  NAND U9345 ( .A(n61097), .B(n8612), .Z(n8613) );
  NAND U9346 ( .A(n61098), .B(n8613), .Z(n8614) );
  ANDN U9347 ( .B(n61099), .A(n50501), .Z(n8615) );
  NAND U9348 ( .A(n8614), .B(n8615), .Z(n8616) );
  NAND U9349 ( .A(n50500), .B(n8616), .Z(n8617) );
  ANDN U9350 ( .B(n61101), .A(n61100), .Z(n8618) );
  NAND U9351 ( .A(n8617), .B(n8618), .Z(n8619) );
  NAND U9352 ( .A(n61102), .B(n8619), .Z(n8620) );
  AND U9353 ( .A(n61103), .B(n61104), .Z(n8621) );
  NAND U9354 ( .A(n8620), .B(n8621), .Z(n8622) );
  NANDN U9355 ( .A(n61105), .B(n8622), .Z(n8623) );
  ANDN U9356 ( .B(n50499), .A(n50498), .Z(n8624) );
  NAND U9357 ( .A(n8623), .B(n8624), .Z(n8625) );
  NAND U9358 ( .A(n61106), .B(n8625), .Z(n8626) );
  AND U9359 ( .A(n61107), .B(n8626), .Z(n8627) );
  AND U9360 ( .A(n61108), .B(n8627), .Z(n61111) );
  AND U9361 ( .A(n61133), .B(n61132), .Z(n8628) );
  NANDN U9362 ( .A(n61131), .B(n61130), .Z(n8629) );
  AND U9363 ( .A(n8628), .B(n8629), .Z(n8630) );
  NANDN U9364 ( .A(n8630), .B(n61134), .Z(n8631) );
  AND U9365 ( .A(n61135), .B(n8631), .Z(n8632) );
  OR U9366 ( .A(n50484), .B(n8632), .Z(n8633) );
  NAND U9367 ( .A(n50483), .B(n8633), .Z(n8634) );
  NAND U9368 ( .A(n61136), .B(n8634), .Z(n8635) );
  AND U9369 ( .A(n61138), .B(n61137), .Z(n8636) );
  NAND U9370 ( .A(n8635), .B(n8636), .Z(n8637) );
  NAND U9371 ( .A(n61139), .B(n8637), .Z(n8638) );
  ANDN U9372 ( .B(n50481), .A(n50482), .Z(n8639) );
  NAND U9373 ( .A(n8638), .B(n8639), .Z(n8640) );
  NAND U9374 ( .A(n50480), .B(n8640), .Z(n8641) );
  ANDN U9375 ( .B(n8641), .A(n61140), .Z(n61142) );
  NAND U9376 ( .A(n61173), .B(n61172), .Z(n8642) );
  NAND U9377 ( .A(n61174), .B(n8642), .Z(n8643) );
  AND U9378 ( .A(n61175), .B(n8643), .Z(n8644) );
  NANDN U9379 ( .A(n50472), .B(n8644), .Z(n8645) );
  NANDN U9380 ( .A(n61176), .B(n8645), .Z(n8646) );
  ANDN U9381 ( .B(n8646), .A(n61177), .Z(n8647) );
  AND U9382 ( .A(n61178), .B(n8647), .Z(n8648) );
  ANDN U9383 ( .B(n50470), .A(n50471), .Z(n8649) );
  NANDN U9384 ( .A(n8648), .B(n61179), .Z(n8650) );
  AND U9385 ( .A(n8649), .B(n8650), .Z(n8651) );
  ANDN U9386 ( .B(n61181), .A(n61182), .Z(n8652) );
  NANDN U9387 ( .A(n8651), .B(n61180), .Z(n8653) );
  AND U9388 ( .A(n8652), .B(n8653), .Z(n8654) );
  ANDN U9389 ( .B(n61183), .A(n61184), .Z(n8655) );
  NANDN U9390 ( .A(n8654), .B(n50469), .Z(n8656) );
  AND U9391 ( .A(n8655), .B(n8656), .Z(n61186) );
  ANDN U9392 ( .B(n61239), .A(n61238), .Z(n8657) );
  NAND U9393 ( .A(n61236), .B(n61237), .Z(n8658) );
  AND U9394 ( .A(n8657), .B(n8658), .Z(n8659) );
  ANDN U9395 ( .B(n50461), .A(n50462), .Z(n8660) );
  NANDN U9396 ( .A(n8659), .B(n61240), .Z(n8661) );
  AND U9397 ( .A(n8660), .B(n8661), .Z(n8662) );
  NANDN U9398 ( .A(n8662), .B(n61241), .Z(n8663) );
  NAND U9399 ( .A(n61242), .B(n8663), .Z(n8664) );
  NANDN U9400 ( .A(n61243), .B(n8664), .Z(n8665) );
  NAND U9401 ( .A(n61244), .B(n8665), .Z(n8666) );
  NAND U9402 ( .A(n50460), .B(n8666), .Z(n8667) );
  AND U9403 ( .A(n61245), .B(n8667), .Z(n8668) );
  NANDN U9404 ( .A(n8668), .B(n61246), .Z(n8669) );
  ANDN U9405 ( .B(n8669), .A(n61247), .Z(n8670) );
  ANDN U9406 ( .B(n50459), .A(n50458), .Z(n8671) );
  NANDN U9407 ( .A(n8670), .B(n61248), .Z(n8672) );
  AND U9408 ( .A(n8671), .B(n8672), .Z(n61250) );
  IV U9409 ( .A(ebreg), .Z(e) );
  NANDN U9410 ( .A(x[8190]), .B(y[8190]), .Z(n8674) );
  NANDN U9411 ( .A(x[8189]), .B(y[8189]), .Z(n8673) );
  AND U9412 ( .A(n8674), .B(n8673), .Z(n61282) );
  NANDN U9413 ( .A(y[8190]), .B(x[8190]), .Z(n50443) );
  NANDN U9414 ( .A(x[8182]), .B(y[8182]), .Z(n50445) );
  AND U9415 ( .A(n50443), .B(n50445), .Z(n8676) );
  XNOR U9416 ( .A(y[8191]), .B(x[8191]), .Z(n8675) );
  AND U9417 ( .A(n8676), .B(n8675), .Z(n8679) );
  NANDN U9418 ( .A(x[8187]), .B(y[8187]), .Z(n8678) );
  NANDN U9419 ( .A(x[8188]), .B(y[8188]), .Z(n8677) );
  AND U9420 ( .A(n8678), .B(n8677), .Z(n61280) );
  AND U9421 ( .A(n8679), .B(n61280), .Z(n8680) );
  AND U9422 ( .A(n61282), .B(n8680), .Z(n8682) );
  NANDN U9423 ( .A(x[8183]), .B(y[8183]), .Z(n21861) );
  NANDN U9424 ( .A(x[8184]), .B(y[8184]), .Z(n8681) );
  AND U9425 ( .A(n21861), .B(n8681), .Z(n61276) );
  AND U9426 ( .A(n8682), .B(n61276), .Z(n8690) );
  NANDN U9427 ( .A(x[8186]), .B(y[8186]), .Z(n8684) );
  NANDN U9428 ( .A(x[8185]), .B(y[8185]), .Z(n8683) );
  AND U9429 ( .A(n8684), .B(n8683), .Z(n61278) );
  NANDN U9430 ( .A(y[8186]), .B(x[8186]), .Z(n21866) );
  NANDN U9431 ( .A(y[8188]), .B(x[8188]), .Z(n8686) );
  NANDN U9432 ( .A(y[8189]), .B(x[8189]), .Z(n8685) );
  AND U9433 ( .A(n8686), .B(n8685), .Z(n61281) );
  AND U9434 ( .A(n21866), .B(n61281), .Z(n8688) );
  NANDN U9435 ( .A(y[8187]), .B(x[8187]), .Z(n8687) );
  AND U9436 ( .A(n8688), .B(n8687), .Z(n61279) );
  AND U9437 ( .A(n61278), .B(n61279), .Z(n8689) );
  AND U9438 ( .A(n8690), .B(n8689), .Z(n21868) );
  NANDN U9439 ( .A(y[8182]), .B(x[8182]), .Z(n8692) );
  NANDN U9440 ( .A(y[8183]), .B(x[8183]), .Z(n8691) );
  AND U9441 ( .A(n8692), .B(n8691), .Z(n61275) );
  ANDN U9442 ( .B(y[8181]), .A(x[8181]), .Z(n50444) );
  XNOR U9443 ( .A(x[8182]), .B(y[8182]), .Z(n21870) );
  NANDN U9444 ( .A(y[8180]), .B(x[8180]), .Z(n8693) );
  NANDN U9445 ( .A(y[8181]), .B(x[8181]), .Z(n21869) );
  NAND U9446 ( .A(n8693), .B(n21869), .Z(n61273) );
  NANDN U9447 ( .A(y[8178]), .B(x[8178]), .Z(n8694) );
  NANDN U9448 ( .A(y[8179]), .B(x[8179]), .Z(n50433) );
  AND U9449 ( .A(n8694), .B(n50433), .Z(n61270) );
  XNOR U9450 ( .A(x[8178]), .B(y[8178]), .Z(n21872) );
  NANDN U9451 ( .A(y[8176]), .B(x[8176]), .Z(n8695) );
  NANDN U9452 ( .A(y[8177]), .B(x[8177]), .Z(n21871) );
  AND U9453 ( .A(n8695), .B(n21871), .Z(n61269) );
  XNOR U9454 ( .A(x[8176]), .B(y[8176]), .Z(n50424) );
  ANDN U9455 ( .B(y[8175]), .A(x[8175]), .Z(n50420) );
  ANDN U9456 ( .B(n50424), .A(n50420), .Z(n21850) );
  XNOR U9457 ( .A(x[8174]), .B(y[8174]), .Z(n21874) );
  XNOR U9458 ( .A(x[8172]), .B(y[8172]), .Z(n21876) );
  NANDN U9459 ( .A(y[8170]), .B(x[8170]), .Z(n8696) );
  NANDN U9460 ( .A(y[8171]), .B(x[8171]), .Z(n21875) );
  NAND U9461 ( .A(n8696), .B(n21875), .Z(n50448) );
  XNOR U9462 ( .A(x[8170]), .B(y[8170]), .Z(n21878) );
  NANDN U9463 ( .A(x[8169]), .B(y[8169]), .Z(n61258) );
  AND U9464 ( .A(n21878), .B(n61258), .Z(n21839) );
  NANDN U9465 ( .A(y[8168]), .B(x[8168]), .Z(n8697) );
  NANDN U9466 ( .A(y[8169]), .B(x[8169]), .Z(n21877) );
  NAND U9467 ( .A(n8697), .B(n21877), .Z(n61257) );
  XNOR U9468 ( .A(x[8168]), .B(y[8168]), .Z(n21880) );
  NANDN U9469 ( .A(y[8166]), .B(x[8166]), .Z(n8698) );
  NANDN U9470 ( .A(y[8167]), .B(x[8167]), .Z(n21879) );
  AND U9471 ( .A(n8698), .B(n21879), .Z(n61256) );
  ANDN U9472 ( .B(y[8165]), .A(x[8165]), .Z(n61254) );
  XNOR U9473 ( .A(x[8166]), .B(y[8166]), .Z(n21882) );
  NANDN U9474 ( .A(n61254), .B(n21882), .Z(n21833) );
  NANDN U9475 ( .A(y[8164]), .B(x[8164]), .Z(n8699) );
  NANDN U9476 ( .A(y[8165]), .B(x[8165]), .Z(n21881) );
  AND U9477 ( .A(n8699), .B(n21881), .Z(n61253) );
  NANDN U9478 ( .A(y[8162]), .B(x[8162]), .Z(n8700) );
  NANDN U9479 ( .A(y[8163]), .B(x[8163]), .Z(n50397) );
  AND U9480 ( .A(n8700), .B(n50397), .Z(n61252) );
  ANDN U9481 ( .B(y[8161]), .A(x[8161]), .Z(n50454) );
  XNOR U9482 ( .A(x[8162]), .B(y[8162]), .Z(n21884) );
  NANDN U9483 ( .A(y[8160]), .B(x[8160]), .Z(n8701) );
  NANDN U9484 ( .A(y[8161]), .B(x[8161]), .Z(n21883) );
  NAND U9485 ( .A(n8701), .B(n21883), .Z(n61251) );
  NANDN U9486 ( .A(x[8159]), .B(y[8159]), .Z(n50455) );
  XNOR U9487 ( .A(x[8160]), .B(y[8160]), .Z(n50387) );
  NANDN U9488 ( .A(y[8158]), .B(x[8158]), .Z(n8702) );
  NANDN U9489 ( .A(y[8159]), .B(x[8159]), .Z(n50386) );
  AND U9490 ( .A(n8702), .B(n50386), .Z(n61249) );
  ANDN U9491 ( .B(y[8157]), .A(x[8157]), .Z(n50458) );
  XNOR U9492 ( .A(x[8158]), .B(y[8158]), .Z(n21886) );
  NANDN U9493 ( .A(y[8156]), .B(x[8156]), .Z(n21887) );
  NANDN U9494 ( .A(y[8157]), .B(x[8157]), .Z(n21885) );
  AND U9495 ( .A(n21887), .B(n21885), .Z(n61248) );
  NANDN U9496 ( .A(x[8155]), .B(y[8155]), .Z(n21889) );
  NANDN U9497 ( .A(x[8156]), .B(y[8156]), .Z(n50380) );
  NAND U9498 ( .A(n21889), .B(n50380), .Z(n61247) );
  NANDN U9499 ( .A(y[8154]), .B(x[8154]), .Z(n21891) );
  NANDN U9500 ( .A(y[8155]), .B(x[8155]), .Z(n21888) );
  AND U9501 ( .A(n21891), .B(n21888), .Z(n61246) );
  NANDN U9502 ( .A(x[8151]), .B(y[8151]), .Z(n21895) );
  NANDN U9503 ( .A(x[8152]), .B(y[8152]), .Z(n50371) );
  AND U9504 ( .A(n21895), .B(n50371), .Z(n61244) );
  NANDN U9505 ( .A(y[8150]), .B(x[8150]), .Z(n21897) );
  NANDN U9506 ( .A(y[8151]), .B(x[8151]), .Z(n21894) );
  NAND U9507 ( .A(n21897), .B(n21894), .Z(n61243) );
  NANDN U9508 ( .A(x[8150]), .B(y[8150]), .Z(n21896) );
  ANDN U9509 ( .B(y[8149]), .A(x[8149]), .Z(n21899) );
  ANDN U9510 ( .B(n21896), .A(n21899), .Z(n61242) );
  XNOR U9511 ( .A(x[8148]), .B(y[8148]), .Z(n50358) );
  NANDN U9512 ( .A(y[8146]), .B(x[8146]), .Z(n8703) );
  NANDN U9513 ( .A(y[8147]), .B(x[8147]), .Z(n50357) );
  AND U9514 ( .A(n8703), .B(n50357), .Z(n61240) );
  ANDN U9515 ( .B(y[8145]), .A(x[8145]), .Z(n61238) );
  NANDN U9516 ( .A(y[8144]), .B(x[8144]), .Z(n8704) );
  NANDN U9517 ( .A(y[8145]), .B(x[8145]), .Z(n21901) );
  AND U9518 ( .A(n8704), .B(n21901), .Z(n61237) );
  XNOR U9519 ( .A(x[8144]), .B(y[8144]), .Z(n50348) );
  NANDN U9520 ( .A(y[8142]), .B(x[8142]), .Z(n8705) );
  NANDN U9521 ( .A(y[8143]), .B(x[8143]), .Z(n50347) );
  NAND U9522 ( .A(n8705), .B(n50347), .Z(n61231) );
  NANDN U9523 ( .A(y[8140]), .B(x[8140]), .Z(n8706) );
  NANDN U9524 ( .A(y[8141]), .B(x[8141]), .Z(n21902) );
  AND U9525 ( .A(n8706), .B(n21902), .Z(n61225) );
  XNOR U9526 ( .A(x[8140]), .B(y[8140]), .Z(n50338) );
  NANDN U9527 ( .A(x[8139]), .B(y[8139]), .Z(n61221) );
  AND U9528 ( .A(n50338), .B(n61221), .Z(n21799) );
  XNOR U9529 ( .A(x[8138]), .B(y[8138]), .Z(n21905) );
  NANDN U9530 ( .A(y[8136]), .B(x[8136]), .Z(n8707) );
  NANDN U9531 ( .A(y[8137]), .B(x[8137]), .Z(n21904) );
  AND U9532 ( .A(n8707), .B(n21904), .Z(n61214) );
  XNOR U9533 ( .A(x[8136]), .B(y[8136]), .Z(n21907) );
  ANDN U9534 ( .B(y[8135]), .A(x[8135]), .Z(n50326) );
  ANDN U9535 ( .B(n21907), .A(n50326), .Z(n21792) );
  XNOR U9536 ( .A(x[8134]), .B(y[8134]), .Z(n21909) );
  NANDN U9537 ( .A(y[8132]), .B(x[8132]), .Z(n8708) );
  NANDN U9538 ( .A(y[8133]), .B(x[8133]), .Z(n21908) );
  AND U9539 ( .A(n8708), .B(n21908), .Z(n61204) );
  XNOR U9540 ( .A(x[8132]), .B(y[8132]), .Z(n50319) );
  NANDN U9541 ( .A(y[8130]), .B(x[8130]), .Z(n8709) );
  NANDN U9542 ( .A(y[8131]), .B(x[8131]), .Z(n50318) );
  AND U9543 ( .A(n8709), .B(n50318), .Z(n61199) );
  XNOR U9544 ( .A(x[8128]), .B(y[8128]), .Z(n21914) );
  NANDN U9545 ( .A(y[8126]), .B(x[8126]), .Z(n8710) );
  NANDN U9546 ( .A(y[8127]), .B(x[8127]), .Z(n21913) );
  NAND U9547 ( .A(n8710), .B(n21913), .Z(n61193) );
  XNOR U9548 ( .A(x[8126]), .B(y[8126]), .Z(n21916) );
  NANDN U9549 ( .A(x[8125]), .B(y[8125]), .Z(n61192) );
  AND U9550 ( .A(n21916), .B(n61192), .Z(n21775) );
  XNOR U9551 ( .A(x[8124]), .B(y[8124]), .Z(n50301) );
  NANDN U9552 ( .A(y[8122]), .B(x[8122]), .Z(n8711) );
  NANDN U9553 ( .A(y[8123]), .B(x[8123]), .Z(n50300) );
  AND U9554 ( .A(n8711), .B(n50300), .Z(n61189) );
  ANDN U9555 ( .B(y[8121]), .A(x[8121]), .Z(n61187) );
  XNOR U9556 ( .A(x[8122]), .B(y[8122]), .Z(n21918) );
  NANDN U9557 ( .A(y[8120]), .B(x[8120]), .Z(n8712) );
  NANDN U9558 ( .A(y[8121]), .B(x[8121]), .Z(n21917) );
  NAND U9559 ( .A(n8712), .B(n21917), .Z(n61185) );
  XNOR U9560 ( .A(x[8120]), .B(y[8120]), .Z(n50291) );
  ANDN U9561 ( .B(y[8119]), .A(x[8119]), .Z(n50287) );
  ANDN U9562 ( .B(y[8117]), .A(x[8117]), .Z(n61182) );
  XNOR U9563 ( .A(x[8118]), .B(y[8118]), .Z(n21920) );
  NANDN U9564 ( .A(y[8116]), .B(x[8116]), .Z(n8713) );
  NANDN U9565 ( .A(y[8117]), .B(x[8117]), .Z(n21919) );
  AND U9566 ( .A(n8713), .B(n21919), .Z(n61180) );
  NANDN U9567 ( .A(y[8114]), .B(x[8114]), .Z(n8714) );
  NANDN U9568 ( .A(y[8115]), .B(x[8115]), .Z(n50279) );
  AND U9569 ( .A(n8714), .B(n50279), .Z(n61179) );
  ANDN U9570 ( .B(y[8113]), .A(x[8113]), .Z(n61177) );
  XNOR U9571 ( .A(x[8114]), .B(y[8114]), .Z(n21922) );
  NANDN U9572 ( .A(y[8112]), .B(x[8112]), .Z(n8715) );
  NANDN U9573 ( .A(y[8113]), .B(x[8113]), .Z(n21921) );
  NAND U9574 ( .A(n8715), .B(n21921), .Z(n61176) );
  XNOR U9575 ( .A(x[8112]), .B(y[8112]), .Z(n50270) );
  NANDN U9576 ( .A(x[8111]), .B(y[8111]), .Z(n61175) );
  AND U9577 ( .A(n50270), .B(n61175), .Z(n21752) );
  XNOR U9578 ( .A(x[8110]), .B(y[8110]), .Z(n21924) );
  NANDN U9579 ( .A(y[8108]), .B(x[8108]), .Z(n8716) );
  NANDN U9580 ( .A(y[8109]), .B(x[8109]), .Z(n21923) );
  AND U9581 ( .A(n8716), .B(n21923), .Z(n61170) );
  XNOR U9582 ( .A(x[8108]), .B(y[8108]), .Z(n21926) );
  NANDN U9583 ( .A(x[8107]), .B(y[8107]), .Z(n61169) );
  AND U9584 ( .A(n21926), .B(n61169), .Z(n21745) );
  XNOR U9585 ( .A(x[8106]), .B(y[8106]), .Z(n21928) );
  NANDN U9586 ( .A(y[8104]), .B(x[8104]), .Z(n8717) );
  NANDN U9587 ( .A(y[8105]), .B(x[8105]), .Z(n21927) );
  AND U9588 ( .A(n8717), .B(n21927), .Z(n61164) );
  XNOR U9589 ( .A(x[8104]), .B(y[8104]), .Z(n50252) );
  ANDN U9590 ( .B(y[8103]), .A(x[8103]), .Z(n50248) );
  ANDN U9591 ( .B(n50252), .A(n50248), .Z(n21738) );
  XNOR U9592 ( .A(x[8102]), .B(y[8102]), .Z(n21930) );
  NANDN U9593 ( .A(y[8100]), .B(x[8100]), .Z(n8718) );
  NANDN U9594 ( .A(y[8101]), .B(x[8101]), .Z(n21929) );
  AND U9595 ( .A(n8718), .B(n21929), .Z(n61160) );
  XNOR U9596 ( .A(x[8100]), .B(y[8100]), .Z(n50241) );
  NANDN U9597 ( .A(y[8098]), .B(x[8098]), .Z(n8719) );
  NANDN U9598 ( .A(y[8099]), .B(x[8099]), .Z(n50240) );
  NAND U9599 ( .A(n8719), .B(n50240), .Z(n61158) );
  NANDN U9600 ( .A(y[8096]), .B(x[8096]), .Z(n8720) );
  NANDN U9601 ( .A(y[8097]), .B(x[8097]), .Z(n21931) );
  AND U9602 ( .A(n8720), .B(n21931), .Z(n61154) );
  XNOR U9603 ( .A(x[8096]), .B(y[8096]), .Z(n50231) );
  NANDN U9604 ( .A(y[8094]), .B(x[8094]), .Z(n8721) );
  NANDN U9605 ( .A(y[8095]), .B(x[8095]), .Z(n50230) );
  NAND U9606 ( .A(n8721), .B(n50230), .Z(n61151) );
  XNOR U9607 ( .A(x[8094]), .B(y[8094]), .Z(n21934) );
  ANDN U9608 ( .B(y[8093]), .A(x[8093]), .Z(n50476) );
  ANDN U9609 ( .B(n21934), .A(n50476), .Z(n21722) );
  NANDN U9610 ( .A(y[8092]), .B(x[8092]), .Z(n8722) );
  NANDN U9611 ( .A(y[8093]), .B(x[8093]), .Z(n21933) );
  NAND U9612 ( .A(n8722), .B(n21933), .Z(n61150) );
  XNOR U9613 ( .A(x[8092]), .B(y[8092]), .Z(n50221) );
  NANDN U9614 ( .A(y[8090]), .B(x[8090]), .Z(n8723) );
  NANDN U9615 ( .A(y[8091]), .B(x[8091]), .Z(n50220) );
  AND U9616 ( .A(n8723), .B(n50220), .Z(n61147) );
  XNOR U9617 ( .A(x[8090]), .B(y[8090]), .Z(n21936) );
  NANDN U9618 ( .A(x[8089]), .B(y[8089]), .Z(n21937) );
  AND U9619 ( .A(n21936), .B(n21937), .Z(n21716) );
  XNOR U9620 ( .A(x[8088]), .B(y[8088]), .Z(n50211) );
  NANDN U9621 ( .A(y[8086]), .B(x[8086]), .Z(n8724) );
  NANDN U9622 ( .A(y[8087]), .B(x[8087]), .Z(n50210) );
  AND U9623 ( .A(n8724), .B(n50210), .Z(n61143) );
  ANDN U9624 ( .B(y[8085]), .A(x[8085]), .Z(n61140) );
  XNOR U9625 ( .A(x[8086]), .B(y[8086]), .Z(n21939) );
  NANDN U9626 ( .A(n61140), .B(n21939), .Z(n21709) );
  NANDN U9627 ( .A(y[8084]), .B(x[8084]), .Z(n8725) );
  NANDN U9628 ( .A(y[8085]), .B(x[8085]), .Z(n21938) );
  AND U9629 ( .A(n8725), .B(n21938), .Z(n50480) );
  NANDN U9630 ( .A(x[8083]), .B(y[8083]), .Z(n50481) );
  XNOR U9631 ( .A(x[8084]), .B(y[8084]), .Z(n50201) );
  NAND U9632 ( .A(n50481), .B(n50201), .Z(n21706) );
  NANDN U9633 ( .A(y[8082]), .B(x[8082]), .Z(n8726) );
  NANDN U9634 ( .A(y[8083]), .B(x[8083]), .Z(n50200) );
  AND U9635 ( .A(n8726), .B(n50200), .Z(n61139) );
  XNOR U9636 ( .A(x[8082]), .B(y[8082]), .Z(n21941) );
  NANDN U9637 ( .A(y[8081]), .B(x[8081]), .Z(n21940) );
  ANDN U9638 ( .B(x[8080]), .A(y[8080]), .Z(n50191) );
  ANDN U9639 ( .B(n21940), .A(n50191), .Z(n61136) );
  NANDN U9640 ( .A(x[8079]), .B(y[8079]), .Z(n21943) );
  NANDN U9641 ( .A(x[8080]), .B(y[8080]), .Z(n21942) );
  AND U9642 ( .A(n21943), .B(n21942), .Z(n50483) );
  NANDN U9643 ( .A(y[8076]), .B(x[8076]), .Z(n8727) );
  NANDN U9644 ( .A(y[8077]), .B(x[8077]), .Z(n21946) );
  AND U9645 ( .A(n8727), .B(n21946), .Z(n61134) );
  XNOR U9646 ( .A(x[8076]), .B(y[8076]), .Z(n21949) );
  NANDN U9647 ( .A(x[8075]), .B(y[8075]), .Z(n61132) );
  NANDN U9648 ( .A(y[8074]), .B(x[8074]), .Z(n8728) );
  NANDN U9649 ( .A(y[8075]), .B(x[8075]), .Z(n21948) );
  NAND U9650 ( .A(n8728), .B(n21948), .Z(n61131) );
  XNOR U9651 ( .A(x[8072]), .B(y[8072]), .Z(n50173) );
  NANDN U9652 ( .A(y[8070]), .B(x[8070]), .Z(n8729) );
  NANDN U9653 ( .A(y[8071]), .B(x[8071]), .Z(n50172) );
  AND U9654 ( .A(n8729), .B(n50172), .Z(n61126) );
  NANDN U9655 ( .A(y[8068]), .B(x[8068]), .Z(n8730) );
  NANDN U9656 ( .A(y[8069]), .B(x[8069]), .Z(n21952) );
  AND U9657 ( .A(n8730), .B(n21952), .Z(n61125) );
  XNOR U9658 ( .A(x[8068]), .B(y[8068]), .Z(n50163) );
  NANDN U9659 ( .A(y[8066]), .B(x[8066]), .Z(n21955) );
  NANDN U9660 ( .A(y[8067]), .B(x[8067]), .Z(n50162) );
  NAND U9661 ( .A(n21955), .B(n50162), .Z(n61124) );
  NANDN U9662 ( .A(x[8066]), .B(y[8066]), .Z(n21954) );
  ANDN U9663 ( .B(y[8065]), .A(x[8065]), .Z(n21957) );
  ANDN U9664 ( .B(n21954), .A(n21957), .Z(n61123) );
  NANDN U9665 ( .A(y[8064]), .B(x[8064]), .Z(n8731) );
  NANDN U9666 ( .A(y[8065]), .B(x[8065]), .Z(n21956) );
  AND U9667 ( .A(n8731), .B(n21956), .Z(n50491) );
  XNOR U9668 ( .A(x[8064]), .B(y[8064]), .Z(n50153) );
  ANDN U9669 ( .B(y[8063]), .A(x[8063]), .Z(n50149) );
  ANDN U9670 ( .B(n50153), .A(n50149), .Z(n21678) );
  XNOR U9671 ( .A(x[8062]), .B(y[8062]), .Z(n21959) );
  NANDN U9672 ( .A(y[8060]), .B(x[8060]), .Z(n21961) );
  NANDN U9673 ( .A(y[8061]), .B(x[8061]), .Z(n21958) );
  AND U9674 ( .A(n21961), .B(n21958), .Z(n61117) );
  NANDN U9675 ( .A(x[8059]), .B(y[8059]), .Z(n21963) );
  NANDN U9676 ( .A(x[8060]), .B(y[8060]), .Z(n21960) );
  AND U9677 ( .A(n21963), .B(n21960), .Z(n50494) );
  XNOR U9678 ( .A(x[8058]), .B(y[8058]), .Z(n21965) );
  NANDN U9679 ( .A(y[8056]), .B(x[8056]), .Z(n8732) );
  NANDN U9680 ( .A(y[8057]), .B(x[8057]), .Z(n21964) );
  AND U9681 ( .A(n8732), .B(n21964), .Z(n61114) );
  ANDN U9682 ( .B(y[8055]), .A(x[8055]), .Z(n50131) );
  NANDN U9683 ( .A(y[8054]), .B(x[8054]), .Z(n21968) );
  NANDN U9684 ( .A(y[8055]), .B(x[8055]), .Z(n21966) );
  AND U9685 ( .A(n21968), .B(n21966), .Z(n50496) );
  XNOR U9686 ( .A(x[8052]), .B(y[8052]), .Z(n21971) );
  NANDN U9687 ( .A(y[8050]), .B(x[8050]), .Z(n8733) );
  NANDN U9688 ( .A(y[8051]), .B(x[8051]), .Z(n21970) );
  AND U9689 ( .A(n8733), .B(n21970), .Z(n61106) );
  XNOR U9690 ( .A(x[8050]), .B(y[8050]), .Z(n21973) );
  NANDN U9691 ( .A(x[8049]), .B(y[8049]), .Z(n21974) );
  AND U9692 ( .A(n21973), .B(n21974), .Z(n21656) );
  XNOR U9693 ( .A(x[8048]), .B(y[8048]), .Z(n50115) );
  NANDN U9694 ( .A(y[8046]), .B(x[8046]), .Z(n8734) );
  NANDN U9695 ( .A(y[8047]), .B(x[8047]), .Z(n50114) );
  AND U9696 ( .A(n8734), .B(n50114), .Z(n61102) );
  ANDN U9697 ( .B(y[8045]), .A(x[8045]), .Z(n61100) );
  XNOR U9698 ( .A(x[8046]), .B(y[8046]), .Z(n21976) );
  NANDN U9699 ( .A(n61100), .B(n21976), .Z(n21649) );
  NANDN U9700 ( .A(y[8044]), .B(x[8044]), .Z(n8735) );
  NANDN U9701 ( .A(y[8045]), .B(x[8045]), .Z(n21975) );
  AND U9702 ( .A(n8735), .B(n21975), .Z(n50500) );
  XNOR U9703 ( .A(x[8044]), .B(y[8044]), .Z(n50105) );
  NANDN U9704 ( .A(x[8043]), .B(y[8043]), .Z(n61099) );
  NAND U9705 ( .A(n50105), .B(n61099), .Z(n21646) );
  NANDN U9706 ( .A(y[8042]), .B(x[8042]), .Z(n8736) );
  NANDN U9707 ( .A(y[8043]), .B(x[8043]), .Z(n50104) );
  AND U9708 ( .A(n8736), .B(n50104), .Z(n61098) );
  ANDN U9709 ( .B(y[8041]), .A(x[8041]), .Z(n61095) );
  XNOR U9710 ( .A(x[8042]), .B(y[8042]), .Z(n21978) );
  NANDN U9711 ( .A(y[8040]), .B(x[8040]), .Z(n8737) );
  NANDN U9712 ( .A(y[8041]), .B(x[8041]), .Z(n21977) );
  NAND U9713 ( .A(n8737), .B(n21977), .Z(n61094) );
  XNOR U9714 ( .A(x[8040]), .B(y[8040]), .Z(n50095) );
  ANDN U9715 ( .B(y[8039]), .A(x[8039]), .Z(n50091) );
  ANDN U9716 ( .B(y[8037]), .A(x[8037]), .Z(n61091) );
  XNOR U9717 ( .A(x[8038]), .B(y[8038]), .Z(n21980) );
  NANDN U9718 ( .A(y[8036]), .B(x[8036]), .Z(n8738) );
  NANDN U9719 ( .A(y[8037]), .B(x[8037]), .Z(n21979) );
  AND U9720 ( .A(n8738), .B(n21979), .Z(n61090) );
  XNOR U9721 ( .A(x[8036]), .B(y[8036]), .Z(n50084) );
  NANDN U9722 ( .A(x[8035]), .B(y[8035]), .Z(n50504) );
  AND U9723 ( .A(n50084), .B(n50504), .Z(n21633) );
  XNOR U9724 ( .A(x[8034]), .B(y[8034]), .Z(n21982) );
  NANDN U9725 ( .A(y[8032]), .B(x[8032]), .Z(n8739) );
  NANDN U9726 ( .A(y[8033]), .B(x[8033]), .Z(n21981) );
  AND U9727 ( .A(n8739), .B(n21981), .Z(n61086) );
  XNOR U9728 ( .A(x[8032]), .B(y[8032]), .Z(n50074) );
  NANDN U9729 ( .A(x[8031]), .B(y[8031]), .Z(n61084) );
  NAND U9730 ( .A(n50074), .B(n61084), .Z(n21626) );
  NANDN U9731 ( .A(y[8030]), .B(x[8030]), .Z(n8740) );
  NANDN U9732 ( .A(y[8031]), .B(x[8031]), .Z(n50073) );
  AND U9733 ( .A(n8740), .B(n50073), .Z(n50506) );
  NANDN U9734 ( .A(y[8028]), .B(x[8028]), .Z(n8741) );
  NANDN U9735 ( .A(y[8029]), .B(x[8029]), .Z(n21983) );
  AND U9736 ( .A(n8741), .B(n21983), .Z(n61080) );
  XNOR U9737 ( .A(x[8028]), .B(y[8028]), .Z(n50064) );
  NANDN U9738 ( .A(y[8026]), .B(x[8026]), .Z(n8742) );
  NANDN U9739 ( .A(y[8027]), .B(x[8027]), .Z(n50063) );
  NAND U9740 ( .A(n8742), .B(n50063), .Z(n61077) );
  XNOR U9741 ( .A(x[8026]), .B(y[8026]), .Z(n21986) );
  NANDN U9742 ( .A(y[8024]), .B(x[8024]), .Z(n8743) );
  NANDN U9743 ( .A(y[8025]), .B(x[8025]), .Z(n21985) );
  AND U9744 ( .A(n8743), .B(n21985), .Z(n61076) );
  XNOR U9745 ( .A(x[8024]), .B(y[8024]), .Z(n50054) );
  ANDN U9746 ( .B(y[8023]), .A(x[8023]), .Z(n50050) );
  ANDN U9747 ( .B(n50054), .A(n50050), .Z(n21614) );
  XNOR U9748 ( .A(x[8022]), .B(y[8022]), .Z(n21988) );
  NANDN U9749 ( .A(x[8021]), .B(y[8021]), .Z(n21989) );
  AND U9750 ( .A(n21988), .B(n21989), .Z(n21610) );
  XNOR U9751 ( .A(x[8020]), .B(y[8020]), .Z(n50043) );
  NANDN U9752 ( .A(y[8018]), .B(x[8018]), .Z(n8744) );
  NANDN U9753 ( .A(y[8019]), .B(x[8019]), .Z(n50042) );
  AND U9754 ( .A(n8744), .B(n50042), .Z(n61069) );
  XNOR U9755 ( .A(x[8018]), .B(y[8018]), .Z(n21991) );
  ANDN U9756 ( .B(y[8017]), .A(x[8017]), .Z(n61066) );
  ANDN U9757 ( .B(n21991), .A(n61066), .Z(n21603) );
  XNOR U9758 ( .A(x[8016]), .B(y[8016]), .Z(n50033) );
  NANDN U9759 ( .A(y[8014]), .B(x[8014]), .Z(n8745) );
  NANDN U9760 ( .A(y[8015]), .B(x[8015]), .Z(n50032) );
  AND U9761 ( .A(n8745), .B(n50032), .Z(n61063) );
  ANDN U9762 ( .B(y[8013]), .A(x[8013]), .Z(n61061) );
  XNOR U9763 ( .A(x[8014]), .B(y[8014]), .Z(n21993) );
  NANDN U9764 ( .A(y[8012]), .B(x[8012]), .Z(n8746) );
  NANDN U9765 ( .A(y[8013]), .B(x[8013]), .Z(n21992) );
  NAND U9766 ( .A(n8746), .B(n21992), .Z(n61060) );
  ANDN U9767 ( .B(y[8009]), .A(x[8009]), .Z(n61057) );
  XNOR U9768 ( .A(x[8010]), .B(y[8010]), .Z(n21995) );
  NANDN U9769 ( .A(y[8008]), .B(x[8008]), .Z(n8747) );
  NANDN U9770 ( .A(y[8009]), .B(x[8009]), .Z(n21994) );
  AND U9771 ( .A(n8747), .B(n21994), .Z(n61056) );
  XNOR U9772 ( .A(x[8008]), .B(y[8008]), .Z(n50013) );
  NANDN U9773 ( .A(x[8007]), .B(y[8007]), .Z(n50514) );
  AND U9774 ( .A(n50013), .B(n50514), .Z(n21586) );
  XNOR U9775 ( .A(x[8006]), .B(y[8006]), .Z(n21997) );
  NANDN U9776 ( .A(y[8004]), .B(x[8004]), .Z(n8748) );
  NANDN U9777 ( .A(y[8005]), .B(x[8005]), .Z(n21996) );
  AND U9778 ( .A(n8748), .B(n21996), .Z(n61050) );
  XNOR U9779 ( .A(x[8004]), .B(y[8004]), .Z(n21999) );
  NANDN U9780 ( .A(x[8003]), .B(y[8003]), .Z(n61048) );
  AND U9781 ( .A(n21999), .B(n61048), .Z(n21579) );
  XNOR U9782 ( .A(x[8002]), .B(y[8002]), .Z(n22001) );
  ANDN U9783 ( .B(x[7999]), .A(y[7999]), .Z(n49995) );
  NANDN U9784 ( .A(y[7998]), .B(x[7998]), .Z(n8749) );
  NANDN U9785 ( .A(n49995), .B(n8749), .Z(n61041) );
  XNOR U9786 ( .A(x[7996]), .B(y[7996]), .Z(n49985) );
  NANDN U9787 ( .A(y[7994]), .B(x[7994]), .Z(n8750) );
  NANDN U9788 ( .A(y[7995]), .B(x[7995]), .Z(n49984) );
  AND U9789 ( .A(n8750), .B(n49984), .Z(n61035) );
  XNOR U9790 ( .A(x[7994]), .B(y[7994]), .Z(n22005) );
  NANDN U9791 ( .A(x[7993]), .B(y[7993]), .Z(n50518) );
  AND U9792 ( .A(n22005), .B(n50518), .Z(n21561) );
  XNOR U9793 ( .A(x[7992]), .B(y[7992]), .Z(n22007) );
  NANDN U9794 ( .A(y[7990]), .B(x[7990]), .Z(n8751) );
  NANDN U9795 ( .A(y[7991]), .B(x[7991]), .Z(n22006) );
  AND U9796 ( .A(n8751), .B(n22006), .Z(n61031) );
  XNOR U9797 ( .A(x[7990]), .B(y[7990]), .Z(n22009) );
  ANDN U9798 ( .B(y[7989]), .A(x[7989]), .Z(n61029) );
  ANDN U9799 ( .B(n22009), .A(n61029), .Z(n21554) );
  XNOR U9800 ( .A(x[7988]), .B(y[7988]), .Z(n49967) );
  NANDN U9801 ( .A(y[7986]), .B(x[7986]), .Z(n8752) );
  NANDN U9802 ( .A(y[7987]), .B(x[7987]), .Z(n49966) );
  AND U9803 ( .A(n8752), .B(n49966), .Z(n61026) );
  XNOR U9804 ( .A(x[7986]), .B(y[7986]), .Z(n22011) );
  ANDN U9805 ( .B(y[7985]), .A(x[7985]), .Z(n61024) );
  ANDN U9806 ( .B(n22011), .A(n61024), .Z(n21547) );
  XNOR U9807 ( .A(x[7984]), .B(y[7984]), .Z(n49957) );
  NANDN U9808 ( .A(y[7982]), .B(x[7982]), .Z(n8753) );
  NANDN U9809 ( .A(y[7983]), .B(x[7983]), .Z(n49956) );
  AND U9810 ( .A(n8753), .B(n49956), .Z(n61021) );
  XNOR U9811 ( .A(x[7982]), .B(y[7982]), .Z(n22013) );
  XNOR U9812 ( .A(x[7980]), .B(y[7980]), .Z(n22015) );
  XNOR U9813 ( .A(x[7978]), .B(y[7978]), .Z(n22017) );
  NANDN U9814 ( .A(y[7976]), .B(x[7976]), .Z(n8754) );
  NANDN U9815 ( .A(y[7977]), .B(x[7977]), .Z(n22016) );
  AND U9816 ( .A(n8754), .B(n22016), .Z(n61014) );
  XNOR U9817 ( .A(x[7976]), .B(y[7976]), .Z(n49939) );
  NANDN U9818 ( .A(x[7975]), .B(y[7975]), .Z(n61012) );
  AND U9819 ( .A(n49939), .B(n61012), .Z(n21529) );
  NANDN U9820 ( .A(y[7974]), .B(x[7974]), .Z(n8755) );
  NANDN U9821 ( .A(y[7975]), .B(x[7975]), .Z(n49938) );
  NAND U9822 ( .A(n8755), .B(n49938), .Z(n61011) );
  XNOR U9823 ( .A(x[7974]), .B(y[7974]), .Z(n22019) );
  NANDN U9824 ( .A(y[7972]), .B(x[7972]), .Z(n8756) );
  NANDN U9825 ( .A(y[7973]), .B(x[7973]), .Z(n22018) );
  AND U9826 ( .A(n8756), .B(n22018), .Z(n61008) );
  XNOR U9827 ( .A(x[7972]), .B(y[7972]), .Z(n49929) );
  ANDN U9828 ( .B(y[7971]), .A(x[7971]), .Z(n49925) );
  ANDN U9829 ( .B(n49929), .A(n49925), .Z(n21523) );
  XNOR U9830 ( .A(x[7970]), .B(y[7970]), .Z(n22021) );
  NANDN U9831 ( .A(y[7968]), .B(x[7968]), .Z(n22022) );
  NANDN U9832 ( .A(y[7969]), .B(x[7969]), .Z(n22020) );
  AND U9833 ( .A(n22022), .B(n22020), .Z(n61002) );
  NANDN U9834 ( .A(x[7967]), .B(y[7967]), .Z(n22024) );
  ANDN U9835 ( .B(y[7968]), .A(x[7968]), .Z(n49921) );
  ANDN U9836 ( .B(n22024), .A(n49921), .Z(n61001) );
  NANDN U9837 ( .A(y[7966]), .B(x[7966]), .Z(n22026) );
  NANDN U9838 ( .A(y[7967]), .B(x[7967]), .Z(n22023) );
  AND U9839 ( .A(n22026), .B(n22023), .Z(n61000) );
  NANDN U9840 ( .A(x[7966]), .B(y[7966]), .Z(n22025) );
  ANDN U9841 ( .B(y[7965]), .A(x[7965]), .Z(n22028) );
  ANDN U9842 ( .B(n22025), .A(n22028), .Z(n60999) );
  XNOR U9843 ( .A(x[7964]), .B(y[7964]), .Z(n49909) );
  NANDN U9844 ( .A(y[7962]), .B(x[7962]), .Z(n8757) );
  NANDN U9845 ( .A(y[7963]), .B(x[7963]), .Z(n49908) );
  AND U9846 ( .A(n8757), .B(n49908), .Z(n60998) );
  XNOR U9847 ( .A(x[7962]), .B(y[7962]), .Z(n22030) );
  ANDN U9848 ( .B(y[7961]), .A(x[7961]), .Z(n60996) );
  ANDN U9849 ( .B(n22030), .A(n60996), .Z(n21508) );
  NANDN U9850 ( .A(y[7960]), .B(x[7960]), .Z(n8758) );
  NANDN U9851 ( .A(y[7961]), .B(x[7961]), .Z(n22029) );
  NAND U9852 ( .A(n8758), .B(n22029), .Z(n60995) );
  XNOR U9853 ( .A(x[7960]), .B(y[7960]), .Z(n22032) );
  NANDN U9854 ( .A(y[7958]), .B(x[7958]), .Z(n22034) );
  NANDN U9855 ( .A(y[7959]), .B(x[7959]), .Z(n22031) );
  AND U9856 ( .A(n22034), .B(n22031), .Z(n60990) );
  NANDN U9857 ( .A(x[7958]), .B(y[7958]), .Z(n22033) );
  ANDN U9858 ( .B(y[7957]), .A(x[7957]), .Z(n22036) );
  ANDN U9859 ( .B(n22033), .A(n22036), .Z(n60989) );
  NANDN U9860 ( .A(y[7956]), .B(x[7956]), .Z(n8759) );
  NANDN U9861 ( .A(y[7957]), .B(x[7957]), .Z(n22035) );
  AND U9862 ( .A(n8759), .B(n22035), .Z(n60988) );
  NANDN U9863 ( .A(x[7955]), .B(y[7955]), .Z(n50530) );
  XNOR U9864 ( .A(x[7956]), .B(y[7956]), .Z(n49891) );
  NAND U9865 ( .A(n50530), .B(n49891), .Z(n21500) );
  NANDN U9866 ( .A(y[7954]), .B(x[7954]), .Z(n8760) );
  NANDN U9867 ( .A(y[7955]), .B(x[7955]), .Z(n49890) );
  AND U9868 ( .A(n8760), .B(n49890), .Z(n60987) );
  ANDN U9869 ( .B(y[7953]), .A(x[7953]), .Z(n60985) );
  XNOR U9870 ( .A(x[7954]), .B(y[7954]), .Z(n22038) );
  NANDN U9871 ( .A(y[7952]), .B(x[7952]), .Z(n8761) );
  NANDN U9872 ( .A(y[7953]), .B(x[7953]), .Z(n22037) );
  AND U9873 ( .A(n8761), .B(n22037), .Z(n60984) );
  XNOR U9874 ( .A(x[7952]), .B(y[7952]), .Z(n22040) );
  ANDN U9875 ( .B(y[7951]), .A(x[7951]), .Z(n49879) );
  NANDN U9876 ( .A(y[7948]), .B(x[7948]), .Z(n8762) );
  NANDN U9877 ( .A(y[7949]), .B(x[7949]), .Z(n22041) );
  AND U9878 ( .A(n8762), .B(n22041), .Z(n60980) );
  XNOR U9879 ( .A(x[7948]), .B(y[7948]), .Z(n49872) );
  ANDN U9880 ( .B(y[7947]), .A(x[7947]), .Z(n49868) );
  ANDN U9881 ( .B(n49872), .A(n49868), .Z(n21487) );
  XNOR U9882 ( .A(x[7946]), .B(y[7946]), .Z(n22044) );
  NANDN U9883 ( .A(y[7944]), .B(x[7944]), .Z(n8763) );
  NANDN U9884 ( .A(y[7945]), .B(x[7945]), .Z(n22043) );
  AND U9885 ( .A(n8763), .B(n22043), .Z(n60976) );
  XNOR U9886 ( .A(x[7944]), .B(y[7944]), .Z(n22046) );
  NANDN U9887 ( .A(y[7942]), .B(x[7942]), .Z(n8764) );
  NANDN U9888 ( .A(y[7943]), .B(x[7943]), .Z(n22045) );
  AND U9889 ( .A(n8764), .B(n22045), .Z(n60973) );
  NANDN U9890 ( .A(y[7940]), .B(x[7940]), .Z(n8765) );
  NANDN U9891 ( .A(y[7941]), .B(x[7941]), .Z(n22047) );
  AND U9892 ( .A(n8765), .B(n22047), .Z(n60972) );
  XNOR U9893 ( .A(x[7940]), .B(y[7940]), .Z(n49853) );
  NANDN U9894 ( .A(y[7938]), .B(x[7938]), .Z(n8766) );
  NANDN U9895 ( .A(y[7939]), .B(x[7939]), .Z(n49852) );
  AND U9896 ( .A(n8766), .B(n49852), .Z(n60969) );
  XNOR U9897 ( .A(x[7938]), .B(y[7938]), .Z(n22051) );
  ANDN U9898 ( .B(y[7937]), .A(x[7937]), .Z(n60967) );
  ANDN U9899 ( .B(n22051), .A(n60967), .Z(n21471) );
  NANDN U9900 ( .A(y[7936]), .B(x[7936]), .Z(n8767) );
  NANDN U9901 ( .A(y[7937]), .B(x[7937]), .Z(n22050) );
  NAND U9902 ( .A(n8767), .B(n22050), .Z(n60966) );
  XNOR U9903 ( .A(x[7936]), .B(y[7936]), .Z(n49843) );
  NANDN U9904 ( .A(y[7934]), .B(x[7934]), .Z(n8768) );
  NANDN U9905 ( .A(y[7935]), .B(x[7935]), .Z(n49842) );
  AND U9906 ( .A(n8768), .B(n49842), .Z(n60963) );
  ANDN U9907 ( .B(y[7933]), .A(x[7933]), .Z(n60961) );
  XNOR U9908 ( .A(x[7934]), .B(y[7934]), .Z(n22053) );
  NANDN U9909 ( .A(n60961), .B(n22053), .Z(n21465) );
  NANDN U9910 ( .A(y[7932]), .B(x[7932]), .Z(n8769) );
  NANDN U9911 ( .A(y[7933]), .B(x[7933]), .Z(n22052) );
  AND U9912 ( .A(n8769), .B(n22052), .Z(n50540) );
  XNOR U9913 ( .A(x[7932]), .B(y[7932]), .Z(n49833) );
  NANDN U9914 ( .A(x[7931]), .B(y[7931]), .Z(n50542) );
  NAND U9915 ( .A(n49833), .B(n50542), .Z(n21462) );
  ANDN U9916 ( .B(y[7929]), .A(x[7929]), .Z(n60958) );
  XNOR U9917 ( .A(x[7930]), .B(y[7930]), .Z(n22055) );
  NANDN U9918 ( .A(y[7928]), .B(x[7928]), .Z(n8770) );
  NANDN U9919 ( .A(y[7929]), .B(x[7929]), .Z(n22054) );
  AND U9920 ( .A(n8770), .B(n22054), .Z(n60957) );
  NANDN U9921 ( .A(x[7927]), .B(y[7927]), .Z(n50543) );
  XNOR U9922 ( .A(x[7928]), .B(y[7928]), .Z(n49823) );
  NANDN U9923 ( .A(y[7926]), .B(x[7926]), .Z(n8771) );
  NANDN U9924 ( .A(y[7927]), .B(x[7927]), .Z(n49822) );
  NAND U9925 ( .A(n8771), .B(n49822), .Z(n60956) );
  NANDN U9926 ( .A(y[7924]), .B(x[7924]), .Z(n8772) );
  NANDN U9927 ( .A(y[7925]), .B(x[7925]), .Z(n22056) );
  AND U9928 ( .A(n8772), .B(n22056), .Z(n60952) );
  XNOR U9929 ( .A(x[7924]), .B(y[7924]), .Z(n49813) );
  ANDN U9930 ( .B(y[7923]), .A(x[7923]), .Z(n49809) );
  ANDN U9931 ( .B(n49813), .A(n49809), .Z(n21449) );
  XNOR U9932 ( .A(x[7922]), .B(y[7922]), .Z(n22059) );
  NANDN U9933 ( .A(y[7920]), .B(x[7920]), .Z(n8773) );
  NANDN U9934 ( .A(y[7921]), .B(x[7921]), .Z(n22058) );
  AND U9935 ( .A(n8773), .B(n22058), .Z(n60947) );
  XNOR U9936 ( .A(x[7920]), .B(y[7920]), .Z(n49802) );
  NANDN U9937 ( .A(y[7918]), .B(x[7918]), .Z(n8774) );
  NANDN U9938 ( .A(y[7919]), .B(x[7919]), .Z(n49801) );
  NAND U9939 ( .A(n8774), .B(n49801), .Z(n60944) );
  XNOR U9940 ( .A(x[7916]), .B(y[7916]), .Z(n49792) );
  NANDN U9941 ( .A(y[7914]), .B(x[7914]), .Z(n8775) );
  NANDN U9942 ( .A(y[7915]), .B(x[7915]), .Z(n49791) );
  AND U9943 ( .A(n8775), .B(n49791), .Z(n60940) );
  XNOR U9944 ( .A(x[7914]), .B(y[7914]), .Z(n22063) );
  NANDN U9945 ( .A(x[7913]), .B(y[7913]), .Z(n22064) );
  AND U9946 ( .A(n22063), .B(n22064), .Z(n21432) );
  XNOR U9947 ( .A(x[7912]), .B(y[7912]), .Z(n49782) );
  NANDN U9948 ( .A(y[7910]), .B(x[7910]), .Z(n8776) );
  NANDN U9949 ( .A(y[7911]), .B(x[7911]), .Z(n49781) );
  AND U9950 ( .A(n8776), .B(n49781), .Z(n60934) );
  ANDN U9951 ( .B(y[7909]), .A(x[7909]), .Z(n60932) );
  XNOR U9952 ( .A(x[7910]), .B(y[7910]), .Z(n22066) );
  NANDN U9953 ( .A(n60932), .B(n22066), .Z(n21425) );
  NANDN U9954 ( .A(y[7908]), .B(x[7908]), .Z(n8777) );
  NANDN U9955 ( .A(y[7909]), .B(x[7909]), .Z(n22065) );
  AND U9956 ( .A(n8777), .B(n22065), .Z(n50550) );
  XNOR U9957 ( .A(x[7908]), .B(y[7908]), .Z(n49772) );
  NANDN U9958 ( .A(x[7907]), .B(y[7907]), .Z(n60931) );
  NAND U9959 ( .A(n49772), .B(n60931), .Z(n21422) );
  NANDN U9960 ( .A(y[7906]), .B(x[7906]), .Z(n8778) );
  NANDN U9961 ( .A(y[7907]), .B(x[7907]), .Z(n49771) );
  AND U9962 ( .A(n8778), .B(n49771), .Z(n60930) );
  ANDN U9963 ( .B(y[7905]), .A(x[7905]), .Z(n60928) );
  XNOR U9964 ( .A(x[7906]), .B(y[7906]), .Z(n22068) );
  NANDN U9965 ( .A(y[7904]), .B(x[7904]), .Z(n8779) );
  NANDN U9966 ( .A(y[7905]), .B(x[7905]), .Z(n22067) );
  NAND U9967 ( .A(n8779), .B(n22067), .Z(n60927) );
  ANDN U9968 ( .B(y[7901]), .A(x[7901]), .Z(n60922) );
  XNOR U9969 ( .A(x[7902]), .B(y[7902]), .Z(n22070) );
  NANDN U9970 ( .A(y[7900]), .B(x[7900]), .Z(n8780) );
  NANDN U9971 ( .A(y[7901]), .B(x[7901]), .Z(n22069) );
  AND U9972 ( .A(n8780), .B(n22069), .Z(n60921) );
  XNOR U9973 ( .A(x[7900]), .B(y[7900]), .Z(n49752) );
  NANDN U9974 ( .A(x[7899]), .B(y[7899]), .Z(n50554) );
  AND U9975 ( .A(n49752), .B(n50554), .Z(n21409) );
  XNOR U9976 ( .A(x[7898]), .B(y[7898]), .Z(n22072) );
  NANDN U9977 ( .A(y[7896]), .B(x[7896]), .Z(n8781) );
  NANDN U9978 ( .A(y[7897]), .B(x[7897]), .Z(n22071) );
  AND U9979 ( .A(n8781), .B(n22071), .Z(n60917) );
  XNOR U9980 ( .A(x[7896]), .B(y[7896]), .Z(n49742) );
  ANDN U9981 ( .B(y[7895]), .A(x[7895]), .Z(n49738) );
  ANDN U9982 ( .B(n49742), .A(n49738), .Z(n21402) );
  XNOR U9983 ( .A(x[7894]), .B(y[7894]), .Z(n22074) );
  NANDN U9984 ( .A(y[7892]), .B(x[7892]), .Z(n8782) );
  NANDN U9985 ( .A(y[7893]), .B(x[7893]), .Z(n22073) );
  AND U9986 ( .A(n8782), .B(n22073), .Z(n60912) );
  XNOR U9987 ( .A(x[7892]), .B(y[7892]), .Z(n22076) );
  NANDN U9988 ( .A(y[7890]), .B(x[7890]), .Z(n8783) );
  NANDN U9989 ( .A(y[7891]), .B(x[7891]), .Z(n22075) );
  NAND U9990 ( .A(n8783), .B(n22075), .Z(n60908) );
  ANDN U9991 ( .B(y[7889]), .A(x[7889]), .Z(n50557) );
  XNOR U9992 ( .A(x[7890]), .B(y[7890]), .Z(n22078) );
  NANDN U9993 ( .A(y[7888]), .B(x[7888]), .Z(n8784) );
  NANDN U9994 ( .A(y[7889]), .B(x[7889]), .Z(n22077) );
  AND U9995 ( .A(n8784), .B(n22077), .Z(n60907) );
  XNOR U9996 ( .A(x[7888]), .B(y[7888]), .Z(n49723) );
  NANDN U9997 ( .A(y[7886]), .B(x[7886]), .Z(n8785) );
  NANDN U9998 ( .A(y[7887]), .B(x[7887]), .Z(n49722) );
  AND U9999 ( .A(n8785), .B(n49722), .Z(n60904) );
  XNOR U10000 ( .A(x[7886]), .B(y[7886]), .Z(n22080) );
  ANDN U10001 ( .B(y[7885]), .A(x[7885]), .Z(n50560) );
  NANDN U10002 ( .A(y[7884]), .B(x[7884]), .Z(n8786) );
  NANDN U10003 ( .A(y[7885]), .B(x[7885]), .Z(n22079) );
  AND U10004 ( .A(n8786), .B(n22079), .Z(n60903) );
  XNOR U10005 ( .A(x[7884]), .B(y[7884]), .Z(n49713) );
  NANDN U10006 ( .A(y[7882]), .B(x[7882]), .Z(n22082) );
  NANDN U10007 ( .A(y[7883]), .B(x[7883]), .Z(n49712) );
  AND U10008 ( .A(n22082), .B(n49712), .Z(n60900) );
  NANDN U10009 ( .A(x[7881]), .B(y[7881]), .Z(n22084) );
  NANDN U10010 ( .A(x[7882]), .B(y[7882]), .Z(n22081) );
  AND U10011 ( .A(n22084), .B(n22081), .Z(n60899) );
  NANDN U10012 ( .A(y[7880]), .B(x[7880]), .Z(n22086) );
  NANDN U10013 ( .A(y[7881]), .B(x[7881]), .Z(n22083) );
  AND U10014 ( .A(n22086), .B(n22083), .Z(n50561) );
  XNOR U10015 ( .A(x[7878]), .B(y[7878]), .Z(n22090) );
  NANDN U10016 ( .A(y[7876]), .B(x[7876]), .Z(n22092) );
  NANDN U10017 ( .A(y[7877]), .B(x[7877]), .Z(n22089) );
  AND U10018 ( .A(n22092), .B(n22089), .Z(n60893) );
  NANDN U10019 ( .A(x[7875]), .B(y[7875]), .Z(n49693) );
  NANDN U10020 ( .A(x[7876]), .B(y[7876]), .Z(n22091) );
  AND U10021 ( .A(n49693), .B(n22091), .Z(n60892) );
  NANDN U10022 ( .A(y[7874]), .B(x[7874]), .Z(n8787) );
  NANDN U10023 ( .A(y[7875]), .B(x[7875]), .Z(n22093) );
  NAND U10024 ( .A(n8787), .B(n22093), .Z(n60891) );
  XNOR U10025 ( .A(x[7874]), .B(y[7874]), .Z(n22095) );
  NANDN U10026 ( .A(y[7872]), .B(x[7872]), .Z(n22097) );
  NANDN U10027 ( .A(y[7873]), .B(x[7873]), .Z(n22094) );
  AND U10028 ( .A(n22097), .B(n22094), .Z(n60888) );
  NANDN U10029 ( .A(x[7871]), .B(y[7871]), .Z(n49684) );
  NANDN U10030 ( .A(x[7872]), .B(y[7872]), .Z(n22096) );
  NAND U10031 ( .A(n49684), .B(n22096), .Z(n50563) );
  NANDN U10032 ( .A(y[7870]), .B(x[7870]), .Z(n8788) );
  NANDN U10033 ( .A(y[7871]), .B(x[7871]), .Z(n22098) );
  AND U10034 ( .A(n8788), .B(n22098), .Z(n60887) );
  ANDN U10035 ( .B(y[7869]), .A(x[7869]), .Z(n22101) );
  XNOR U10036 ( .A(x[7870]), .B(y[7870]), .Z(n22100) );
  NANDN U10037 ( .A(y[7868]), .B(x[7868]), .Z(n22103) );
  NANDN U10038 ( .A(y[7869]), .B(x[7869]), .Z(n22099) );
  AND U10039 ( .A(n22103), .B(n22099), .Z(n60886) );
  NANDN U10040 ( .A(x[7867]), .B(y[7867]), .Z(n22105) );
  NANDN U10041 ( .A(x[7868]), .B(y[7868]), .Z(n22102) );
  AND U10042 ( .A(n22105), .B(n22102), .Z(n60885) );
  NANDN U10043 ( .A(y[7866]), .B(x[7866]), .Z(n22107) );
  NANDN U10044 ( .A(y[7867]), .B(x[7867]), .Z(n22104) );
  NAND U10045 ( .A(n22107), .B(n22104), .Z(n60882) );
  NANDN U10046 ( .A(x[7865]), .B(y[7865]), .Z(n22109) );
  NANDN U10047 ( .A(x[7866]), .B(y[7866]), .Z(n22106) );
  AND U10048 ( .A(n22109), .B(n22106), .Z(n60881) );
  NANDN U10049 ( .A(y[7864]), .B(x[7864]), .Z(n8789) );
  NANDN U10050 ( .A(y[7865]), .B(x[7865]), .Z(n22108) );
  NAND U10051 ( .A(n8789), .B(n22108), .Z(n60880) );
  NANDN U10052 ( .A(y[7862]), .B(x[7862]), .Z(n22111) );
  ANDN U10053 ( .B(x[7863]), .A(y[7863]), .Z(n49671) );
  ANDN U10054 ( .B(n22111), .A(n49671), .Z(n60879) );
  NANDN U10055 ( .A(x[7861]), .B(y[7861]), .Z(n22113) );
  NANDN U10056 ( .A(x[7862]), .B(y[7862]), .Z(n22110) );
  NAND U10057 ( .A(n22113), .B(n22110), .Z(n60878) );
  NANDN U10058 ( .A(y[7860]), .B(x[7860]), .Z(n8790) );
  NANDN U10059 ( .A(y[7861]), .B(x[7861]), .Z(n22112) );
  AND U10060 ( .A(n8790), .B(n22112), .Z(n50568) );
  XNOR U10061 ( .A(x[7860]), .B(y[7860]), .Z(n22115) );
  NANDN U10062 ( .A(y[7858]), .B(x[7858]), .Z(n8791) );
  NANDN U10063 ( .A(y[7859]), .B(x[7859]), .Z(n22114) );
  AND U10064 ( .A(n8791), .B(n22114), .Z(n60875) );
  ANDN U10065 ( .B(y[7857]), .A(x[7857]), .Z(n60874) );
  XNOR U10066 ( .A(x[7858]), .B(y[7858]), .Z(n22117) );
  NANDN U10067 ( .A(y[7856]), .B(x[7856]), .Z(n8792) );
  NANDN U10068 ( .A(y[7857]), .B(x[7857]), .Z(n22116) );
  NAND U10069 ( .A(n8792), .B(n22116), .Z(n60872) );
  ANDN U10070 ( .B(y[7853]), .A(x[7853]), .Z(n50569) );
  XNOR U10071 ( .A(x[7854]), .B(y[7854]), .Z(n22119) );
  NANDN U10072 ( .A(y[7852]), .B(x[7852]), .Z(n8793) );
  NANDN U10073 ( .A(y[7853]), .B(x[7853]), .Z(n22118) );
  NAND U10074 ( .A(n8793), .B(n22118), .Z(n60866) );
  XNOR U10075 ( .A(x[7852]), .B(y[7852]), .Z(n49641) );
  NANDN U10076 ( .A(x[7851]), .B(y[7851]), .Z(n60864) );
  AND U10077 ( .A(n49641), .B(n60864), .Z(n21340) );
  XNOR U10078 ( .A(x[7850]), .B(y[7850]), .Z(n22121) );
  NANDN U10079 ( .A(y[7848]), .B(x[7848]), .Z(n8794) );
  NANDN U10080 ( .A(y[7849]), .B(x[7849]), .Z(n22120) );
  AND U10081 ( .A(n8794), .B(n22120), .Z(n60860) );
  XNOR U10082 ( .A(x[7848]), .B(y[7848]), .Z(n49631) );
  NANDN U10083 ( .A(x[7847]), .B(y[7847]), .Z(n60859) );
  AND U10084 ( .A(n49631), .B(n60859), .Z(n21333) );
  XNOR U10085 ( .A(x[7846]), .B(y[7846]), .Z(n22123) );
  NANDN U10086 ( .A(y[7844]), .B(x[7844]), .Z(n8795) );
  NANDN U10087 ( .A(y[7845]), .B(x[7845]), .Z(n22122) );
  AND U10088 ( .A(n8795), .B(n22122), .Z(n60855) );
  XNOR U10089 ( .A(x[7844]), .B(y[7844]), .Z(n22125) );
  ANDN U10090 ( .B(y[7843]), .A(x[7843]), .Z(n49619) );
  ANDN U10091 ( .B(n22125), .A(n49619), .Z(n21326) );
  XNOR U10092 ( .A(x[7842]), .B(y[7842]), .Z(n22127) );
  NANDN U10093 ( .A(y[7840]), .B(x[7840]), .Z(n8796) );
  NANDN U10094 ( .A(y[7841]), .B(x[7841]), .Z(n22126) );
  AND U10095 ( .A(n8796), .B(n22126), .Z(n60849) );
  NANDN U10096 ( .A(x[7839]), .B(y[7839]), .Z(n49608) );
  IV U10097 ( .A(n49608), .Z(n50575) );
  XNOR U10098 ( .A(x[7840]), .B(y[7840]), .Z(n49612) );
  NANDN U10099 ( .A(y[7838]), .B(x[7838]), .Z(n8797) );
  NANDN U10100 ( .A(y[7839]), .B(x[7839]), .Z(n49611) );
  NAND U10101 ( .A(n8797), .B(n49611), .Z(n60848) );
  NANDN U10102 ( .A(y[7836]), .B(x[7836]), .Z(n8798) );
  NANDN U10103 ( .A(y[7837]), .B(x[7837]), .Z(n22128) );
  AND U10104 ( .A(n8798), .B(n22128), .Z(n60845) );
  NANDN U10105 ( .A(x[7835]), .B(y[7835]), .Z(n60843) );
  XNOR U10106 ( .A(x[7836]), .B(y[7836]), .Z(n22131) );
  AND U10107 ( .A(n60843), .B(n22131), .Z(n21313) );
  NANDN U10108 ( .A(y[7834]), .B(x[7834]), .Z(n8799) );
  NANDN U10109 ( .A(y[7835]), .B(x[7835]), .Z(n22130) );
  NAND U10110 ( .A(n8799), .B(n22130), .Z(n60842) );
  XNOR U10111 ( .A(x[7834]), .B(y[7834]), .Z(n22133) );
  ANDN U10112 ( .B(y[7833]), .A(x[7833]), .Z(n50576) );
  ANDN U10113 ( .B(n22133), .A(n50576), .Z(n21310) );
  XNOR U10114 ( .A(x[7832]), .B(y[7832]), .Z(n49593) );
  NANDN U10115 ( .A(y[7830]), .B(x[7830]), .Z(n8800) );
  NANDN U10116 ( .A(y[7831]), .B(x[7831]), .Z(n49592) );
  AND U10117 ( .A(n8800), .B(n49592), .Z(n60837) );
  XNOR U10118 ( .A(x[7830]), .B(y[7830]), .Z(n22135) );
  NANDN U10119 ( .A(x[7829]), .B(y[7829]), .Z(n22136) );
  AND U10120 ( .A(n22135), .B(n22136), .Z(n21303) );
  XNOR U10121 ( .A(x[7828]), .B(y[7828]), .Z(n49583) );
  NANDN U10122 ( .A(y[7826]), .B(x[7826]), .Z(n8801) );
  NANDN U10123 ( .A(y[7827]), .B(x[7827]), .Z(n49582) );
  AND U10124 ( .A(n8801), .B(n49582), .Z(n60832) );
  ANDN U10125 ( .B(y[7825]), .A(x[7825]), .Z(n60830) );
  XNOR U10126 ( .A(x[7826]), .B(y[7826]), .Z(n22138) );
  NANDN U10127 ( .A(y[7824]), .B(x[7824]), .Z(n8802) );
  NANDN U10128 ( .A(y[7825]), .B(x[7825]), .Z(n22137) );
  NAND U10129 ( .A(n8802), .B(n22137), .Z(n60829) );
  XNOR U10130 ( .A(x[7824]), .B(y[7824]), .Z(n49573) );
  NANDN U10131 ( .A(x[7823]), .B(y[7823]), .Z(n60828) );
  AND U10132 ( .A(n49573), .B(n60828), .Z(n21293) );
  XNOR U10133 ( .A(x[7822]), .B(y[7822]), .Z(n22140) );
  NANDN U10134 ( .A(y[7820]), .B(x[7820]), .Z(n8803) );
  NANDN U10135 ( .A(y[7821]), .B(x[7821]), .Z(n22139) );
  NAND U10136 ( .A(n8803), .B(n22139), .Z(n60824) );
  XNOR U10137 ( .A(x[7820]), .B(y[7820]), .Z(n49563) );
  NANDN U10138 ( .A(x[7819]), .B(y[7819]), .Z(n50583) );
  AND U10139 ( .A(n49563), .B(n50583), .Z(n21286) );
  NANDN U10140 ( .A(y[7818]), .B(x[7818]), .Z(n8804) );
  NANDN U10141 ( .A(y[7819]), .B(x[7819]), .Z(n49562) );
  NAND U10142 ( .A(n8804), .B(n49562), .Z(n60823) );
  XNOR U10143 ( .A(x[7818]), .B(y[7818]), .Z(n22142) );
  NANDN U10144 ( .A(y[7816]), .B(x[7816]), .Z(n8805) );
  NANDN U10145 ( .A(y[7817]), .B(x[7817]), .Z(n22141) );
  AND U10146 ( .A(n8805), .B(n22141), .Z(n60817) );
  NANDN U10147 ( .A(x[7815]), .B(y[7815]), .Z(n50584) );
  XNOR U10148 ( .A(x[7816]), .B(y[7816]), .Z(n22144) );
  AND U10149 ( .A(n50584), .B(n22144), .Z(n21280) );
  XNOR U10150 ( .A(x[7814]), .B(y[7814]), .Z(n22146) );
  NANDN U10151 ( .A(y[7812]), .B(x[7812]), .Z(n8806) );
  NANDN U10152 ( .A(y[7813]), .B(x[7813]), .Z(n22145) );
  AND U10153 ( .A(n8806), .B(n22145), .Z(n60807) );
  XNOR U10154 ( .A(x[7812]), .B(y[7812]), .Z(n49545) );
  NANDN U10155 ( .A(y[7810]), .B(x[7810]), .Z(n8807) );
  NANDN U10156 ( .A(y[7811]), .B(x[7811]), .Z(n49544) );
  NAND U10157 ( .A(n8807), .B(n49544), .Z(n60801) );
  NANDN U10158 ( .A(y[7808]), .B(x[7808]), .Z(n8808) );
  NANDN U10159 ( .A(y[7809]), .B(x[7809]), .Z(n22147) );
  AND U10160 ( .A(n8808), .B(n22147), .Z(n60795) );
  XNOR U10161 ( .A(x[7808]), .B(y[7808]), .Z(n49535) );
  NANDN U10162 ( .A(y[7806]), .B(x[7806]), .Z(n8809) );
  NANDN U10163 ( .A(y[7807]), .B(x[7807]), .Z(n49534) );
  NAND U10164 ( .A(n8809), .B(n49534), .Z(n60789) );
  XNOR U10165 ( .A(x[7806]), .B(y[7806]), .Z(n22150) );
  NANDN U10166 ( .A(x[7805]), .B(y[7805]), .Z(n60785) );
  AND U10167 ( .A(n22150), .B(n60785), .Z(n21264) );
  XNOR U10168 ( .A(x[7804]), .B(y[7804]), .Z(n49525) );
  NANDN U10169 ( .A(y[7802]), .B(x[7802]), .Z(n8810) );
  NANDN U10170 ( .A(y[7803]), .B(x[7803]), .Z(n49524) );
  AND U10171 ( .A(n8810), .B(n49524), .Z(n60778) );
  XNOR U10172 ( .A(x[7802]), .B(y[7802]), .Z(n22152) );
  ANDN U10173 ( .B(y[7801]), .A(x[7801]), .Z(n50587) );
  ANDN U10174 ( .B(n22152), .A(n50587), .Z(n21257) );
  XNOR U10175 ( .A(x[7800]), .B(y[7800]), .Z(n49515) );
  NANDN U10176 ( .A(y[7798]), .B(x[7798]), .Z(n8811) );
  NANDN U10177 ( .A(y[7799]), .B(x[7799]), .Z(n49514) );
  AND U10178 ( .A(n8811), .B(n49514), .Z(n60777) );
  XNOR U10179 ( .A(x[7798]), .B(y[7798]), .Z(n22154) );
  ANDN U10180 ( .B(y[7797]), .A(x[7797]), .Z(n60775) );
  ANDN U10181 ( .B(n22154), .A(n60775), .Z(n21250) );
  XNOR U10182 ( .A(x[7796]), .B(y[7796]), .Z(n49505) );
  NANDN U10183 ( .A(y[7794]), .B(x[7794]), .Z(n8812) );
  NANDN U10184 ( .A(y[7795]), .B(x[7795]), .Z(n49504) );
  AND U10185 ( .A(n8812), .B(n49504), .Z(n60772) );
  ANDN U10186 ( .B(y[7793]), .A(x[7793]), .Z(n60769) );
  XNOR U10187 ( .A(x[7794]), .B(y[7794]), .Z(n22156) );
  NANDN U10188 ( .A(y[7792]), .B(x[7792]), .Z(n8813) );
  NANDN U10189 ( .A(y[7793]), .B(x[7793]), .Z(n22155) );
  NAND U10190 ( .A(n8813), .B(n22155), .Z(n60768) );
  XNOR U10191 ( .A(x[7792]), .B(y[7792]), .Z(n49495) );
  NANDN U10192 ( .A(y[7790]), .B(x[7790]), .Z(n8814) );
  NANDN U10193 ( .A(y[7791]), .B(x[7791]), .Z(n49494) );
  NAND U10194 ( .A(n8814), .B(n49494), .Z(n60767) );
  XNOR U10195 ( .A(x[7790]), .B(y[7790]), .Z(n22158) );
  ANDN U10196 ( .B(y[7789]), .A(x[7789]), .Z(n60765) );
  NANDN U10197 ( .A(y[7788]), .B(x[7788]), .Z(n8815) );
  NANDN U10198 ( .A(y[7789]), .B(x[7789]), .Z(n22157) );
  AND U10199 ( .A(n8815), .B(n22157), .Z(n60764) );
  XNOR U10200 ( .A(x[7788]), .B(y[7788]), .Z(n49485) );
  ANDN U10201 ( .B(y[7787]), .A(x[7787]), .Z(n49481) );
  ANDN U10202 ( .B(n49485), .A(n49481), .Z(n21234) );
  XNOR U10203 ( .A(x[7786]), .B(y[7786]), .Z(n22160) );
  NANDN U10204 ( .A(y[7784]), .B(x[7784]), .Z(n8816) );
  NANDN U10205 ( .A(y[7785]), .B(x[7785]), .Z(n22159) );
  AND U10206 ( .A(n8816), .B(n22159), .Z(n60762) );
  XNOR U10207 ( .A(x[7784]), .B(y[7784]), .Z(n49474) );
  NANDN U10208 ( .A(y[7782]), .B(x[7782]), .Z(n8817) );
  NANDN U10209 ( .A(y[7783]), .B(x[7783]), .Z(n49473) );
  NAND U10210 ( .A(n8817), .B(n49473), .Z(n60758) );
  XNOR U10211 ( .A(x[7780]), .B(y[7780]), .Z(n49464) );
  NANDN U10212 ( .A(y[7778]), .B(x[7778]), .Z(n8818) );
  NANDN U10213 ( .A(y[7779]), .B(x[7779]), .Z(n49463) );
  AND U10214 ( .A(n8818), .B(n49463), .Z(n60754) );
  XNOR U10215 ( .A(x[7778]), .B(y[7778]), .Z(n22164) );
  NANDN U10216 ( .A(x[7777]), .B(y[7777]), .Z(n22165) );
  AND U10217 ( .A(n22164), .B(n22165), .Z(n21217) );
  XNOR U10218 ( .A(x[7776]), .B(y[7776]), .Z(n49454) );
  NANDN U10219 ( .A(y[7774]), .B(x[7774]), .Z(n8819) );
  NANDN U10220 ( .A(y[7775]), .B(x[7775]), .Z(n49453) );
  AND U10221 ( .A(n8819), .B(n49453), .Z(n60750) );
  XNOR U10222 ( .A(x[7774]), .B(y[7774]), .Z(n22167) );
  NANDN U10223 ( .A(x[7773]), .B(y[7773]), .Z(n60748) );
  NAND U10224 ( .A(n22167), .B(n60748), .Z(n21210) );
  NANDN U10225 ( .A(y[7772]), .B(x[7772]), .Z(n22168) );
  NANDN U10226 ( .A(y[7773]), .B(x[7773]), .Z(n22166) );
  AND U10227 ( .A(n22168), .B(n22166), .Z(n50602) );
  NANDN U10228 ( .A(x[7770]), .B(y[7770]), .Z(n22171) );
  ANDN U10229 ( .B(y[7769]), .A(x[7769]), .Z(n49438) );
  ANDN U10230 ( .B(n22171), .A(n49438), .Z(n60745) );
  NANDN U10231 ( .A(y[7768]), .B(x[7768]), .Z(n8820) );
  NANDN U10232 ( .A(y[7769]), .B(x[7769]), .Z(n22173) );
  AND U10233 ( .A(n8820), .B(n22173), .Z(n60744) );
  XNOR U10234 ( .A(x[7768]), .B(y[7768]), .Z(n22175) );
  ANDN U10235 ( .B(y[7767]), .A(x[7767]), .Z(n22176) );
  ANDN U10236 ( .B(n22175), .A(n22176), .Z(n21203) );
  NANDN U10237 ( .A(x[7766]), .B(y[7766]), .Z(n22177) );
  ANDN U10238 ( .B(y[7765]), .A(x[7765]), .Z(n22180) );
  ANDN U10239 ( .B(n22177), .A(n22180), .Z(n60742) );
  NANDN U10240 ( .A(y[7764]), .B(x[7764]), .Z(n8821) );
  NANDN U10241 ( .A(y[7765]), .B(x[7765]), .Z(n22179) );
  AND U10242 ( .A(n8821), .B(n22179), .Z(n60741) );
  XNOR U10243 ( .A(x[7764]), .B(y[7764]), .Z(n49426) );
  NANDN U10244 ( .A(x[7763]), .B(y[7763]), .Z(n60739) );
  AND U10245 ( .A(n49426), .B(n60739), .Z(n21198) );
  XNOR U10246 ( .A(x[7762]), .B(y[7762]), .Z(n22182) );
  NANDN U10247 ( .A(y[7760]), .B(x[7760]), .Z(n8822) );
  NANDN U10248 ( .A(y[7761]), .B(x[7761]), .Z(n22181) );
  AND U10249 ( .A(n8822), .B(n22181), .Z(n60735) );
  XNOR U10250 ( .A(x[7760]), .B(y[7760]), .Z(n49416) );
  ANDN U10251 ( .B(y[7759]), .A(x[7759]), .Z(n49412) );
  ANDN U10252 ( .B(n49416), .A(n49412), .Z(n21191) );
  XNOR U10253 ( .A(x[7758]), .B(y[7758]), .Z(n22184) );
  NANDN U10254 ( .A(y[7756]), .B(x[7756]), .Z(n8823) );
  NANDN U10255 ( .A(y[7757]), .B(x[7757]), .Z(n22183) );
  AND U10256 ( .A(n8823), .B(n22183), .Z(n60731) );
  XNOR U10257 ( .A(x[7756]), .B(y[7756]), .Z(n49405) );
  NANDN U10258 ( .A(y[7754]), .B(x[7754]), .Z(n8824) );
  NANDN U10259 ( .A(y[7755]), .B(x[7755]), .Z(n49404) );
  AND U10260 ( .A(n8824), .B(n49404), .Z(n60728) );
  NANDN U10261 ( .A(y[7752]), .B(x[7752]), .Z(n8825) );
  NANDN U10262 ( .A(y[7753]), .B(x[7753]), .Z(n22185) );
  AND U10263 ( .A(n8825), .B(n22185), .Z(n60727) );
  XNOR U10264 ( .A(x[7752]), .B(y[7752]), .Z(n49395) );
  NANDN U10265 ( .A(y[7750]), .B(x[7750]), .Z(n8826) );
  NANDN U10266 ( .A(y[7751]), .B(x[7751]), .Z(n49394) );
  AND U10267 ( .A(n8826), .B(n49394), .Z(n60724) );
  XNOR U10268 ( .A(x[7750]), .B(y[7750]), .Z(n22189) );
  ANDN U10269 ( .B(y[7749]), .A(x[7749]), .Z(n60722) );
  ANDN U10270 ( .B(n22189), .A(n60722), .Z(n21175) );
  NANDN U10271 ( .A(y[7748]), .B(x[7748]), .Z(n8827) );
  NANDN U10272 ( .A(y[7749]), .B(x[7749]), .Z(n22188) );
  NAND U10273 ( .A(n8827), .B(n22188), .Z(n60721) );
  XNOR U10274 ( .A(x[7748]), .B(y[7748]), .Z(n49385) );
  NANDN U10275 ( .A(y[7746]), .B(x[7746]), .Z(n8828) );
  NANDN U10276 ( .A(y[7747]), .B(x[7747]), .Z(n49384) );
  AND U10277 ( .A(n8828), .B(n49384), .Z(n60718) );
  ANDN U10278 ( .B(y[7745]), .A(x[7745]), .Z(n60716) );
  XNOR U10279 ( .A(x[7746]), .B(y[7746]), .Z(n22191) );
  NANDN U10280 ( .A(n60716), .B(n22191), .Z(n21169) );
  NANDN U10281 ( .A(y[7744]), .B(x[7744]), .Z(n8829) );
  NANDN U10282 ( .A(y[7745]), .B(x[7745]), .Z(n22190) );
  AND U10283 ( .A(n8829), .B(n22190), .Z(n50612) );
  XNOR U10284 ( .A(x[7744]), .B(y[7744]), .Z(n49375) );
  NANDN U10285 ( .A(x[7743]), .B(y[7743]), .Z(n50614) );
  NAND U10286 ( .A(n49375), .B(n50614), .Z(n21166) );
  ANDN U10287 ( .B(y[7741]), .A(x[7741]), .Z(n60713) );
  XNOR U10288 ( .A(x[7742]), .B(y[7742]), .Z(n22193) );
  NANDN U10289 ( .A(y[7740]), .B(x[7740]), .Z(n8830) );
  NANDN U10290 ( .A(y[7741]), .B(x[7741]), .Z(n22192) );
  AND U10291 ( .A(n8830), .B(n22192), .Z(n60712) );
  NANDN U10292 ( .A(y[7738]), .B(x[7738]), .Z(n8831) );
  NANDN U10293 ( .A(y[7739]), .B(x[7739]), .Z(n49364) );
  AND U10294 ( .A(n8831), .B(n49364), .Z(n60711) );
  ANDN U10295 ( .B(y[7737]), .A(x[7737]), .Z(n60708) );
  XNOR U10296 ( .A(x[7738]), .B(y[7738]), .Z(n22195) );
  NANDN U10297 ( .A(y[7736]), .B(x[7736]), .Z(n8832) );
  NANDN U10298 ( .A(y[7737]), .B(x[7737]), .Z(n22194) );
  AND U10299 ( .A(n8832), .B(n22194), .Z(n60707) );
  NANDN U10300 ( .A(x[7735]), .B(y[7735]), .Z(n60703) );
  XNOR U10301 ( .A(x[7736]), .B(y[7736]), .Z(n49355) );
  NANDN U10302 ( .A(y[7734]), .B(x[7734]), .Z(n8833) );
  NANDN U10303 ( .A(y[7735]), .B(x[7735]), .Z(n49354) );
  AND U10304 ( .A(n8833), .B(n49354), .Z(n60701) );
  NANDN U10305 ( .A(y[7732]), .B(x[7732]), .Z(n8834) );
  NANDN U10306 ( .A(y[7733]), .B(x[7733]), .Z(n22196) );
  AND U10307 ( .A(n8834), .B(n22196), .Z(n60695) );
  XNOR U10308 ( .A(x[7732]), .B(y[7732]), .Z(n49345) );
  NANDN U10309 ( .A(x[7731]), .B(y[7731]), .Z(n60691) );
  AND U10310 ( .A(n49345), .B(n60691), .Z(n21147) );
  XNOR U10311 ( .A(x[7730]), .B(y[7730]), .Z(n22199) );
  NANDN U10312 ( .A(y[7728]), .B(x[7728]), .Z(n8835) );
  NANDN U10313 ( .A(y[7729]), .B(x[7729]), .Z(n22198) );
  AND U10314 ( .A(n8835), .B(n22198), .Z(n60684) );
  NANDN U10315 ( .A(x[7727]), .B(y[7727]), .Z(n60681) );
  XNOR U10316 ( .A(x[7728]), .B(y[7728]), .Z(n22201) );
  AND U10317 ( .A(n60681), .B(n22201), .Z(n21140) );
  XNOR U10318 ( .A(x[7726]), .B(y[7726]), .Z(n22203) );
  NANDN U10319 ( .A(y[7724]), .B(x[7724]), .Z(n8836) );
  NANDN U10320 ( .A(y[7725]), .B(x[7725]), .Z(n22202) );
  AND U10321 ( .A(n8836), .B(n22202), .Z(n60674) );
  XNOR U10322 ( .A(x[7724]), .B(y[7724]), .Z(n49327) );
  NANDN U10323 ( .A(y[7722]), .B(x[7722]), .Z(n8837) );
  NANDN U10324 ( .A(y[7723]), .B(x[7723]), .Z(n49326) );
  AND U10325 ( .A(n8837), .B(n49326), .Z(n60670) );
  XNOR U10326 ( .A(x[7722]), .B(y[7722]), .Z(n22206) );
  ANDN U10327 ( .B(y[7721]), .A(x[7721]), .Z(n60668) );
  ANDN U10328 ( .B(n22206), .A(n60668), .Z(n21130) );
  NANDN U10329 ( .A(y[7720]), .B(x[7720]), .Z(n8838) );
  NANDN U10330 ( .A(y[7721]), .B(x[7721]), .Z(n22205) );
  NAND U10331 ( .A(n8838), .B(n22205), .Z(n60667) );
  XNOR U10332 ( .A(x[7720]), .B(y[7720]), .Z(n49317) );
  NANDN U10333 ( .A(y[7718]), .B(x[7718]), .Z(n8839) );
  NANDN U10334 ( .A(y[7719]), .B(x[7719]), .Z(n49316) );
  AND U10335 ( .A(n8839), .B(n49316), .Z(n60665) );
  XNOR U10336 ( .A(x[7718]), .B(y[7718]), .Z(n22208) );
  NANDN U10337 ( .A(x[7717]), .B(y[7717]), .Z(n60663) );
  AND U10338 ( .A(n22208), .B(n60663), .Z(n21124) );
  NANDN U10339 ( .A(y[7716]), .B(x[7716]), .Z(n8840) );
  NANDN U10340 ( .A(y[7717]), .B(x[7717]), .Z(n22207) );
  NAND U10341 ( .A(n8840), .B(n22207), .Z(n60662) );
  XNOR U10342 ( .A(x[7716]), .B(y[7716]), .Z(n22210) );
  NANDN U10343 ( .A(y[7714]), .B(x[7714]), .Z(n8841) );
  NANDN U10344 ( .A(y[7715]), .B(x[7715]), .Z(n22209) );
  AND U10345 ( .A(n8841), .B(n22209), .Z(n60661) );
  XNOR U10346 ( .A(x[7714]), .B(y[7714]), .Z(n22212) );
  ANDN U10347 ( .B(y[7713]), .A(x[7713]), .Z(n60659) );
  ANDN U10348 ( .B(n22212), .A(n60659), .Z(n21118) );
  XNOR U10349 ( .A(x[7712]), .B(y[7712]), .Z(n49299) );
  NANDN U10350 ( .A(y[7710]), .B(x[7710]), .Z(n8842) );
  NANDN U10351 ( .A(y[7711]), .B(x[7711]), .Z(n49298) );
  AND U10352 ( .A(n8842), .B(n49298), .Z(n60656) );
  XNOR U10353 ( .A(x[7710]), .B(y[7710]), .Z(n22214) );
  ANDN U10354 ( .B(y[7709]), .A(x[7709]), .Z(n60654) );
  ANDN U10355 ( .B(n22214), .A(n60654), .Z(n21111) );
  XNOR U10356 ( .A(x[7708]), .B(y[7708]), .Z(n49289) );
  NANDN U10357 ( .A(y[7706]), .B(x[7706]), .Z(n8843) );
  NANDN U10358 ( .A(y[7707]), .B(x[7707]), .Z(n49288) );
  AND U10359 ( .A(n8843), .B(n49288), .Z(n60650) );
  ANDN U10360 ( .B(y[7705]), .A(x[7705]), .Z(n60648) );
  XNOR U10361 ( .A(x[7706]), .B(y[7706]), .Z(n22216) );
  NANDN U10362 ( .A(y[7704]), .B(x[7704]), .Z(n8844) );
  NANDN U10363 ( .A(y[7705]), .B(x[7705]), .Z(n22215) );
  AND U10364 ( .A(n8844), .B(n22215), .Z(n60647) );
  ANDN U10365 ( .B(y[7701]), .A(x[7701]), .Z(n50628) );
  XNOR U10366 ( .A(x[7702]), .B(y[7702]), .Z(n22218) );
  NANDN U10367 ( .A(y[7700]), .B(x[7700]), .Z(n8845) );
  NANDN U10368 ( .A(y[7701]), .B(x[7701]), .Z(n22217) );
  NAND U10369 ( .A(n8845), .B(n22217), .Z(n60644) );
  XNOR U10370 ( .A(x[7700]), .B(y[7700]), .Z(n49269) );
  ANDN U10371 ( .B(y[7699]), .A(x[7699]), .Z(n22219) );
  NANDN U10372 ( .A(y[7698]), .B(x[7698]), .Z(n22221) );
  NANDN U10373 ( .A(y[7699]), .B(x[7699]), .Z(n49268) );
  AND U10374 ( .A(n22221), .B(n49268), .Z(n60639) );
  NANDN U10375 ( .A(x[7698]), .B(y[7698]), .Z(n22220) );
  ANDN U10376 ( .B(y[7697]), .A(x[7697]), .Z(n22223) );
  ANDN U10377 ( .B(n22220), .A(n22223), .Z(n60638) );
  NANDN U10378 ( .A(y[7696]), .B(x[7696]), .Z(n8846) );
  NANDN U10379 ( .A(y[7697]), .B(x[7697]), .Z(n22222) );
  AND U10380 ( .A(n8846), .B(n22222), .Z(n60637) );
  XNOR U10381 ( .A(x[7696]), .B(y[7696]), .Z(n49259) );
  NANDN U10382 ( .A(x[7695]), .B(y[7695]), .Z(n50631) );
  NAND U10383 ( .A(n49259), .B(n50631), .Z(n21089) );
  NANDN U10384 ( .A(y[7694]), .B(x[7694]), .Z(n8847) );
  NANDN U10385 ( .A(y[7695]), .B(x[7695]), .Z(n49258) );
  AND U10386 ( .A(n8847), .B(n49258), .Z(n60636) );
  ANDN U10387 ( .B(y[7693]), .A(x[7693]), .Z(n60634) );
  XNOR U10388 ( .A(x[7694]), .B(y[7694]), .Z(n22225) );
  NANDN U10389 ( .A(n60634), .B(n22225), .Z(n21086) );
  NANDN U10390 ( .A(x[7691]), .B(y[7691]), .Z(n49245) );
  IV U10391 ( .A(n49245), .Z(n60633) );
  XNOR U10392 ( .A(x[7692]), .B(y[7692]), .Z(n49249) );
  XNOR U10393 ( .A(x[7690]), .B(y[7690]), .Z(n22227) );
  XNOR U10394 ( .A(x[7688]), .B(y[7688]), .Z(n49238) );
  NANDN U10395 ( .A(y[7686]), .B(x[7686]), .Z(n8848) );
  NANDN U10396 ( .A(y[7687]), .B(x[7687]), .Z(n49237) );
  NAND U10397 ( .A(n8848), .B(n49237), .Z(n50636) );
  XNOR U10398 ( .A(x[7686]), .B(y[7686]), .Z(n22229) );
  NANDN U10399 ( .A(x[7685]), .B(y[7685]), .Z(n50637) );
  AND U10400 ( .A(n22229), .B(n50637), .Z(n21071) );
  NANDN U10401 ( .A(x[7683]), .B(y[7683]), .Z(n22233) );
  NANDN U10402 ( .A(x[7684]), .B(y[7684]), .Z(n22230) );
  AND U10403 ( .A(n22233), .B(n22230), .Z(n60625) );
  XNOR U10404 ( .A(x[7682]), .B(y[7682]), .Z(n22235) );
  NANDN U10405 ( .A(y[7680]), .B(x[7680]), .Z(n8849) );
  NANDN U10406 ( .A(y[7681]), .B(x[7681]), .Z(n22234) );
  NAND U10407 ( .A(n8849), .B(n22234), .Z(n60624) );
  NANDN U10408 ( .A(y[7678]), .B(x[7678]), .Z(n8850) );
  NANDN U10409 ( .A(y[7679]), .B(x[7679]), .Z(n49219) );
  AND U10410 ( .A(n8850), .B(n49219), .Z(n60621) );
  XNOR U10411 ( .A(x[7678]), .B(y[7678]), .Z(n22237) );
  NANDN U10412 ( .A(y[7676]), .B(x[7676]), .Z(n8851) );
  NANDN U10413 ( .A(y[7677]), .B(x[7677]), .Z(n22236) );
  NAND U10414 ( .A(n8851), .B(n22236), .Z(n60620) );
  XNOR U10415 ( .A(x[7676]), .B(y[7676]), .Z(n22239) );
  ANDN U10416 ( .B(y[7675]), .A(x[7675]), .Z(n22240) );
  NANDN U10417 ( .A(y[7674]), .B(x[7674]), .Z(n22242) );
  NANDN U10418 ( .A(y[7675]), .B(x[7675]), .Z(n22238) );
  AND U10419 ( .A(n22242), .B(n22238), .Z(n60616) );
  NANDN U10420 ( .A(x[7674]), .B(y[7674]), .Z(n22241) );
  ANDN U10421 ( .B(y[7673]), .A(x[7673]), .Z(n49204) );
  ANDN U10422 ( .B(n22241), .A(n49204), .Z(n60615) );
  NANDN U10423 ( .A(y[7672]), .B(x[7672]), .Z(n22244) );
  NANDN U10424 ( .A(y[7673]), .B(x[7673]), .Z(n22243) );
  AND U10425 ( .A(n22244), .B(n22243), .Z(n60614) );
  NANDN U10426 ( .A(x[7671]), .B(y[7671]), .Z(n22246) );
  NANDN U10427 ( .A(x[7672]), .B(y[7672]), .Z(n49205) );
  AND U10428 ( .A(n22246), .B(n49205), .Z(n60613) );
  NANDN U10429 ( .A(x[7670]), .B(y[7670]), .Z(n22247) );
  ANDN U10430 ( .B(y[7669]), .A(x[7669]), .Z(n22250) );
  ANDN U10431 ( .B(n22247), .A(n22250), .Z(n60611) );
  NANDN U10432 ( .A(y[7668]), .B(x[7668]), .Z(n8852) );
  NANDN U10433 ( .A(y[7669]), .B(x[7669]), .Z(n22249) );
  AND U10434 ( .A(n8852), .B(n22249), .Z(n60610) );
  XNOR U10435 ( .A(x[7668]), .B(y[7668]), .Z(n49192) );
  NANDN U10436 ( .A(y[7666]), .B(x[7666]), .Z(n8853) );
  NANDN U10437 ( .A(y[7667]), .B(x[7667]), .Z(n49191) );
  NAND U10438 ( .A(n8853), .B(n49191), .Z(n50646) );
  NANDN U10439 ( .A(y[7664]), .B(x[7664]), .Z(n8854) );
  NANDN U10440 ( .A(y[7665]), .B(x[7665]), .Z(n22251) );
  AND U10441 ( .A(n8854), .B(n22251), .Z(n60609) );
  XNOR U10442 ( .A(x[7664]), .B(y[7664]), .Z(n49182) );
  NANDN U10443 ( .A(y[7662]), .B(x[7662]), .Z(n8855) );
  NANDN U10444 ( .A(y[7663]), .B(x[7663]), .Z(n49181) );
  NAND U10445 ( .A(n8855), .B(n49181), .Z(n60606) );
  ANDN U10446 ( .B(y[7661]), .A(x[7661]), .Z(n60605) );
  XNOR U10447 ( .A(x[7662]), .B(y[7662]), .Z(n22254) );
  NANDN U10448 ( .A(y[7660]), .B(x[7660]), .Z(n8856) );
  NANDN U10449 ( .A(y[7661]), .B(x[7661]), .Z(n22253) );
  AND U10450 ( .A(n8856), .B(n22253), .Z(n60602) );
  XNOR U10451 ( .A(x[7660]), .B(y[7660]), .Z(n49172) );
  ANDN U10452 ( .B(y[7659]), .A(x[7659]), .Z(n49168) );
  ANDN U10453 ( .B(n49172), .A(n49168), .Z(n21035) );
  XNOR U10454 ( .A(x[7658]), .B(y[7658]), .Z(n22256) );
  NANDN U10455 ( .A(y[7656]), .B(x[7656]), .Z(n8857) );
  NANDN U10456 ( .A(y[7657]), .B(x[7657]), .Z(n22255) );
  NAND U10457 ( .A(n8857), .B(n22255), .Z(n50651) );
  NANDN U10458 ( .A(y[7654]), .B(x[7654]), .Z(n8858) );
  NANDN U10459 ( .A(y[7655]), .B(x[7655]), .Z(n49160) );
  AND U10460 ( .A(n8858), .B(n49160), .Z(n60596) );
  ANDN U10461 ( .B(y[7653]), .A(x[7653]), .Z(n60594) );
  XNOR U10462 ( .A(x[7654]), .B(y[7654]), .Z(n22259) );
  NANDN U10463 ( .A(y[7652]), .B(x[7652]), .Z(n8859) );
  NANDN U10464 ( .A(y[7653]), .B(x[7653]), .Z(n22258) );
  NAND U10465 ( .A(n8859), .B(n22258), .Z(n60593) );
  XNOR U10466 ( .A(x[7652]), .B(y[7652]), .Z(n49151) );
  NANDN U10467 ( .A(x[7651]), .B(y[7651]), .Z(n60590) );
  AND U10468 ( .A(n49151), .B(n60590), .Z(n21022) );
  XNOR U10469 ( .A(x[7650]), .B(y[7650]), .Z(n22261) );
  NANDN U10470 ( .A(y[7648]), .B(x[7648]), .Z(n8860) );
  NANDN U10471 ( .A(y[7649]), .B(x[7649]), .Z(n22260) );
  AND U10472 ( .A(n8860), .B(n22260), .Z(n60584) );
  XNOR U10473 ( .A(x[7648]), .B(y[7648]), .Z(n49141) );
  NANDN U10474 ( .A(x[7647]), .B(y[7647]), .Z(n50653) );
  NAND U10475 ( .A(n49141), .B(n50653), .Z(n21015) );
  NANDN U10476 ( .A(y[7646]), .B(x[7646]), .Z(n8861) );
  NANDN U10477 ( .A(y[7647]), .B(x[7647]), .Z(n49140) );
  AND U10478 ( .A(n8861), .B(n49140), .Z(n60583) );
  ANDN U10479 ( .B(y[7645]), .A(x[7645]), .Z(n60581) );
  XNOR U10480 ( .A(x[7646]), .B(y[7646]), .Z(n22263) );
  NANDN U10481 ( .A(n60581), .B(n22263), .Z(n21012) );
  NANDN U10482 ( .A(x[7643]), .B(y[7643]), .Z(n49127) );
  IV U10483 ( .A(n49127), .Z(n60580) );
  XNOR U10484 ( .A(x[7644]), .B(y[7644]), .Z(n49131) );
  NANDN U10485 ( .A(y[7642]), .B(x[7642]), .Z(n8862) );
  NANDN U10486 ( .A(y[7643]), .B(x[7643]), .Z(n49130) );
  NAND U10487 ( .A(n8862), .B(n49130), .Z(n60578) );
  XNOR U10488 ( .A(x[7642]), .B(y[7642]), .Z(n22265) );
  ANDN U10489 ( .B(y[7641]), .A(x[7641]), .Z(n60576) );
  NANDN U10490 ( .A(y[7640]), .B(x[7640]), .Z(n8863) );
  NANDN U10491 ( .A(y[7641]), .B(x[7641]), .Z(n22264) );
  AND U10492 ( .A(n8863), .B(n22264), .Z(n60575) );
  XNOR U10493 ( .A(x[7640]), .B(y[7640]), .Z(n49120) );
  NANDN U10494 ( .A(y[7638]), .B(x[7638]), .Z(n8864) );
  NANDN U10495 ( .A(y[7639]), .B(x[7639]), .Z(n49119) );
  NAND U10496 ( .A(n8864), .B(n49119), .Z(n60571) );
  XNOR U10497 ( .A(x[7638]), .B(y[7638]), .Z(n22267) );
  ANDN U10498 ( .B(y[7637]), .A(x[7637]), .Z(n50655) );
  ANDN U10499 ( .B(n22267), .A(n50655), .Z(n20999) );
  NANDN U10500 ( .A(y[7636]), .B(x[7636]), .Z(n8865) );
  NANDN U10501 ( .A(y[7637]), .B(x[7637]), .Z(n22266) );
  NAND U10502 ( .A(n8865), .B(n22266), .Z(n60570) );
  XNOR U10503 ( .A(x[7636]), .B(y[7636]), .Z(n22269) );
  NANDN U10504 ( .A(y[7634]), .B(x[7634]), .Z(n8866) );
  NANDN U10505 ( .A(y[7635]), .B(x[7635]), .Z(n22268) );
  AND U10506 ( .A(n8866), .B(n22268), .Z(n60567) );
  ANDN U10507 ( .B(y[7633]), .A(x[7633]), .Z(n60566) );
  XNOR U10508 ( .A(x[7634]), .B(y[7634]), .Z(n22271) );
  NANDN U10509 ( .A(n60566), .B(n22271), .Z(n20993) );
  NANDN U10510 ( .A(y[7632]), .B(x[7632]), .Z(n8867) );
  NANDN U10511 ( .A(y[7633]), .B(x[7633]), .Z(n22270) );
  AND U10512 ( .A(n8867), .B(n22270), .Z(n50658) );
  NANDN U10513 ( .A(y[7630]), .B(x[7630]), .Z(n8868) );
  NANDN U10514 ( .A(y[7631]), .B(x[7631]), .Z(n49101) );
  AND U10515 ( .A(n8868), .B(n49101), .Z(n60564) );
  XNOR U10516 ( .A(x[7630]), .B(y[7630]), .Z(n22273) );
  NANDN U10517 ( .A(y[7628]), .B(x[7628]), .Z(n8869) );
  NANDN U10518 ( .A(y[7629]), .B(x[7629]), .Z(n22272) );
  NAND U10519 ( .A(n8869), .B(n22272), .Z(n60561) );
  XNOR U10520 ( .A(x[7628]), .B(y[7628]), .Z(n22275) );
  NANDN U10521 ( .A(y[7626]), .B(x[7626]), .Z(n8870) );
  NANDN U10522 ( .A(y[7627]), .B(x[7627]), .Z(n22274) );
  AND U10523 ( .A(n8870), .B(n22274), .Z(n60559) );
  XNOR U10524 ( .A(x[7626]), .B(y[7626]), .Z(n22277) );
  ANDN U10525 ( .B(y[7625]), .A(x[7625]), .Z(n60557) );
  ANDN U10526 ( .B(n22277), .A(n60557), .Z(n20981) );
  XNOR U10527 ( .A(x[7624]), .B(y[7624]), .Z(n49084) );
  NANDN U10528 ( .A(x[7623]), .B(y[7623]), .Z(n50662) );
  AND U10529 ( .A(n49084), .B(n50662), .Z(n20977) );
  XNOR U10530 ( .A(x[7622]), .B(y[7622]), .Z(n22279) );
  NANDN U10531 ( .A(y[7620]), .B(x[7620]), .Z(n22281) );
  NANDN U10532 ( .A(y[7621]), .B(x[7621]), .Z(n22278) );
  AND U10533 ( .A(n22281), .B(n22278), .Z(n60555) );
  NANDN U10534 ( .A(x[7619]), .B(y[7619]), .Z(n22283) );
  NANDN U10535 ( .A(x[7620]), .B(y[7620]), .Z(n22280) );
  AND U10536 ( .A(n22283), .B(n22280), .Z(n60554) );
  NANDN U10537 ( .A(y[7618]), .B(x[7618]), .Z(n8871) );
  NANDN U10538 ( .A(y[7619]), .B(x[7619]), .Z(n22282) );
  AND U10539 ( .A(n8871), .B(n22282), .Z(n50667) );
  XNOR U10540 ( .A(x[7618]), .B(y[7618]), .Z(n22285) );
  NANDN U10541 ( .A(y[7616]), .B(x[7616]), .Z(n8872) );
  NANDN U10542 ( .A(y[7617]), .B(x[7617]), .Z(n22284) );
  AND U10543 ( .A(n8872), .B(n22284), .Z(n60552) );
  XNOR U10544 ( .A(x[7616]), .B(y[7616]), .Z(n49066) );
  NANDN U10545 ( .A(y[7614]), .B(x[7614]), .Z(n8873) );
  NANDN U10546 ( .A(y[7615]), .B(x[7615]), .Z(n49065) );
  AND U10547 ( .A(n8873), .B(n49065), .Z(n60549) );
  NANDN U10548 ( .A(y[7612]), .B(x[7612]), .Z(n8874) );
  NANDN U10549 ( .A(y[7613]), .B(x[7613]), .Z(n22286) );
  AND U10550 ( .A(n8874), .B(n22286), .Z(n60548) );
  XNOR U10551 ( .A(x[7612]), .B(y[7612]), .Z(n49056) );
  NANDN U10552 ( .A(y[7610]), .B(x[7610]), .Z(n8875) );
  NANDN U10553 ( .A(y[7611]), .B(x[7611]), .Z(n49055) );
  AND U10554 ( .A(n8875), .B(n49055), .Z(n60545) );
  ANDN U10555 ( .B(y[7609]), .A(x[7609]), .Z(n60543) );
  XNOR U10556 ( .A(x[7610]), .B(y[7610]), .Z(n22290) );
  NANDN U10557 ( .A(y[7608]), .B(x[7608]), .Z(n8876) );
  NANDN U10558 ( .A(y[7609]), .B(x[7609]), .Z(n22289) );
  NAND U10559 ( .A(n8876), .B(n22289), .Z(n60542) );
  XNOR U10560 ( .A(x[7608]), .B(y[7608]), .Z(n49046) );
  ANDN U10561 ( .B(y[7607]), .A(x[7607]), .Z(n49042) );
  NANDN U10562 ( .A(y[7606]), .B(x[7606]), .Z(n8877) );
  NANDN U10563 ( .A(y[7607]), .B(x[7607]), .Z(n49045) );
  AND U10564 ( .A(n8877), .B(n49045), .Z(n60540) );
  ANDN U10565 ( .B(y[7605]), .A(x[7605]), .Z(n60538) );
  XNOR U10566 ( .A(x[7606]), .B(y[7606]), .Z(n22292) );
  NANDN U10567 ( .A(y[7604]), .B(x[7604]), .Z(n8878) );
  NANDN U10568 ( .A(y[7605]), .B(x[7605]), .Z(n22291) );
  NAND U10569 ( .A(n8878), .B(n22291), .Z(n60537) );
  ANDN U10570 ( .B(y[7601]), .A(x[7601]), .Z(n60532) );
  XNOR U10571 ( .A(x[7602]), .B(y[7602]), .Z(n22294) );
  NANDN U10572 ( .A(y[7600]), .B(x[7600]), .Z(n8879) );
  NANDN U10573 ( .A(y[7601]), .B(x[7601]), .Z(n22293) );
  AND U10574 ( .A(n8879), .B(n22293), .Z(n60531) );
  XNOR U10575 ( .A(x[7600]), .B(y[7600]), .Z(n49025) );
  NANDN U10576 ( .A(x[7599]), .B(y[7599]), .Z(n50676) );
  AND U10577 ( .A(n49025), .B(n50676), .Z(n20940) );
  XNOR U10578 ( .A(x[7598]), .B(y[7598]), .Z(n22296) );
  NANDN U10579 ( .A(y[7596]), .B(x[7596]), .Z(n8880) );
  NANDN U10580 ( .A(y[7597]), .B(x[7597]), .Z(n22295) );
  AND U10581 ( .A(n8880), .B(n22295), .Z(n60527) );
  XNOR U10582 ( .A(x[7596]), .B(y[7596]), .Z(n49015) );
  NANDN U10583 ( .A(x[7595]), .B(y[7595]), .Z(n60525) );
  AND U10584 ( .A(n49015), .B(n60525), .Z(n20933) );
  XNOR U10585 ( .A(x[7594]), .B(y[7594]), .Z(n22298) );
  NANDN U10586 ( .A(y[7592]), .B(x[7592]), .Z(n8881) );
  NANDN U10587 ( .A(y[7593]), .B(x[7593]), .Z(n22297) );
  AND U10588 ( .A(n8881), .B(n22297), .Z(n60521) );
  XNOR U10589 ( .A(x[7592]), .B(y[7592]), .Z(n49005) );
  ANDN U10590 ( .B(y[7591]), .A(x[7591]), .Z(n49001) );
  ANDN U10591 ( .B(n49005), .A(n49001), .Z(n20926) );
  XNOR U10592 ( .A(x[7590]), .B(y[7590]), .Z(n22300) );
  NANDN U10593 ( .A(y[7588]), .B(x[7588]), .Z(n8882) );
  NANDN U10594 ( .A(y[7589]), .B(x[7589]), .Z(n22299) );
  AND U10595 ( .A(n8882), .B(n22299), .Z(n60517) );
  XNOR U10596 ( .A(x[7588]), .B(y[7588]), .Z(n48994) );
  NANDN U10597 ( .A(y[7586]), .B(x[7586]), .Z(n8883) );
  NANDN U10598 ( .A(y[7587]), .B(x[7587]), .Z(n48993) );
  AND U10599 ( .A(n8883), .B(n48993), .Z(n60514) );
  NANDN U10600 ( .A(y[7584]), .B(x[7584]), .Z(n8884) );
  NANDN U10601 ( .A(y[7585]), .B(x[7585]), .Z(n22301) );
  AND U10602 ( .A(n8884), .B(n22301), .Z(n60513) );
  XNOR U10603 ( .A(x[7584]), .B(y[7584]), .Z(n48984) );
  NANDN U10604 ( .A(y[7582]), .B(x[7582]), .Z(n8885) );
  NANDN U10605 ( .A(y[7583]), .B(x[7583]), .Z(n48983) );
  NAND U10606 ( .A(n8885), .B(n48983), .Z(n60512) );
  NANDN U10607 ( .A(x[7581]), .B(y[7581]), .Z(n60510) );
  NANDN U10608 ( .A(y[7580]), .B(x[7580]), .Z(n22306) );
  NANDN U10609 ( .A(y[7581]), .B(x[7581]), .Z(n22303) );
  NAND U10610 ( .A(n22306), .B(n22303), .Z(n60508) );
  NANDN U10611 ( .A(x[7579]), .B(y[7579]), .Z(n48972) );
  NANDN U10612 ( .A(x[7580]), .B(y[7580]), .Z(n22305) );
  AND U10613 ( .A(n48972), .B(n22305), .Z(n60507) );
  NANDN U10614 ( .A(y[7578]), .B(x[7578]), .Z(n8886) );
  NANDN U10615 ( .A(y[7579]), .B(x[7579]), .Z(n22307) );
  NAND U10616 ( .A(n8886), .B(n22307), .Z(n60506) );
  XNOR U10617 ( .A(x[7578]), .B(y[7578]), .Z(n22309) );
  NANDN U10618 ( .A(y[7576]), .B(x[7576]), .Z(n8887) );
  NANDN U10619 ( .A(y[7577]), .B(x[7577]), .Z(n22308) );
  AND U10620 ( .A(n8887), .B(n22308), .Z(n60503) );
  NANDN U10621 ( .A(x[7575]), .B(y[7575]), .Z(n50685) );
  XNOR U10622 ( .A(x[7576]), .B(y[7576]), .Z(n22311) );
  NANDN U10623 ( .A(y[7574]), .B(x[7574]), .Z(n22313) );
  NANDN U10624 ( .A(y[7575]), .B(x[7575]), .Z(n22310) );
  NAND U10625 ( .A(n22313), .B(n22310), .Z(n50686) );
  NANDN U10626 ( .A(x[7574]), .B(y[7574]), .Z(n22312) );
  ANDN U10627 ( .B(y[7573]), .A(x[7573]), .Z(n22315) );
  ANDN U10628 ( .B(n22312), .A(n22315), .Z(n60501) );
  XNOR U10629 ( .A(x[7572]), .B(y[7572]), .Z(n48957) );
  NANDN U10630 ( .A(y[7570]), .B(x[7570]), .Z(n8888) );
  NANDN U10631 ( .A(y[7571]), .B(x[7571]), .Z(n48956) );
  NAND U10632 ( .A(n8888), .B(n48956), .Z(n60497) );
  ANDN U10633 ( .B(y[7569]), .A(x[7569]), .Z(n60496) );
  XNOR U10634 ( .A(x[7570]), .B(y[7570]), .Z(n22317) );
  NANDN U10635 ( .A(y[7568]), .B(x[7568]), .Z(n8889) );
  NANDN U10636 ( .A(y[7569]), .B(x[7569]), .Z(n22316) );
  NAND U10637 ( .A(n8889), .B(n22316), .Z(n60493) );
  XNOR U10638 ( .A(x[7568]), .B(y[7568]), .Z(n48947) );
  NANDN U10639 ( .A(x[7567]), .B(y[7567]), .Z(n60492) );
  NANDN U10640 ( .A(y[7566]), .B(x[7566]), .Z(n8890) );
  NANDN U10641 ( .A(y[7567]), .B(x[7567]), .Z(n48946) );
  AND U10642 ( .A(n8890), .B(n48946), .Z(n60490) );
  XNOR U10643 ( .A(x[7566]), .B(y[7566]), .Z(n22319) );
  ANDN U10644 ( .B(y[7565]), .A(x[7565]), .Z(n60488) );
  ANDN U10645 ( .B(n22319), .A(n60488), .Z(n20886) );
  XNOR U10646 ( .A(x[7564]), .B(y[7564]), .Z(n48937) );
  NANDN U10647 ( .A(y[7562]), .B(x[7562]), .Z(n8891) );
  NANDN U10648 ( .A(y[7563]), .B(x[7563]), .Z(n48936) );
  AND U10649 ( .A(n8891), .B(n48936), .Z(n60485) );
  ANDN U10650 ( .B(y[7561]), .A(x[7561]), .Z(n60483) );
  XNOR U10651 ( .A(x[7562]), .B(y[7562]), .Z(n22321) );
  NANDN U10652 ( .A(y[7560]), .B(x[7560]), .Z(n8892) );
  NANDN U10653 ( .A(y[7561]), .B(x[7561]), .Z(n22320) );
  NAND U10654 ( .A(n8892), .B(n22320), .Z(n60482) );
  ANDN U10655 ( .B(y[7557]), .A(x[7557]), .Z(n60477) );
  XNOR U10656 ( .A(x[7558]), .B(y[7558]), .Z(n22323) );
  NANDN U10657 ( .A(y[7556]), .B(x[7556]), .Z(n8893) );
  NANDN U10658 ( .A(y[7557]), .B(x[7557]), .Z(n22322) );
  AND U10659 ( .A(n8893), .B(n22322), .Z(n60476) );
  XNOR U10660 ( .A(x[7556]), .B(y[7556]), .Z(n48917) );
  NANDN U10661 ( .A(x[7555]), .B(y[7555]), .Z(n50691) );
  AND U10662 ( .A(n48917), .B(n50691), .Z(n20869) );
  NANDN U10663 ( .A(y[7554]), .B(x[7554]), .Z(n8894) );
  NANDN U10664 ( .A(y[7555]), .B(x[7555]), .Z(n48916) );
  NAND U10665 ( .A(n8894), .B(n48916), .Z(n60475) );
  XNOR U10666 ( .A(x[7554]), .B(y[7554]), .Z(n22325) );
  NANDN U10667 ( .A(y[7552]), .B(x[7552]), .Z(n8895) );
  NANDN U10668 ( .A(y[7553]), .B(x[7553]), .Z(n22324) );
  AND U10669 ( .A(n8895), .B(n22324), .Z(n60472) );
  XNOR U10670 ( .A(x[7552]), .B(y[7552]), .Z(n48907) );
  NANDN U10671 ( .A(x[7551]), .B(y[7551]), .Z(n60470) );
  NAND U10672 ( .A(n48907), .B(n60470), .Z(n20863) );
  NANDN U10673 ( .A(y[7550]), .B(x[7550]), .Z(n8896) );
  NANDN U10674 ( .A(y[7551]), .B(x[7551]), .Z(n48906) );
  AND U10675 ( .A(n8896), .B(n48906), .Z(n50692) );
  ANDN U10676 ( .B(y[7549]), .A(x[7549]), .Z(n60468) );
  XNOR U10677 ( .A(x[7550]), .B(y[7550]), .Z(n22327) );
  NANDN U10678 ( .A(n60468), .B(n22327), .Z(n20860) );
  NANDN U10679 ( .A(y[7548]), .B(x[7548]), .Z(n8897) );
  NANDN U10680 ( .A(y[7549]), .B(x[7549]), .Z(n22326) );
  AND U10681 ( .A(n8897), .B(n22326), .Z(n60467) );
  XNOR U10682 ( .A(x[7548]), .B(y[7548]), .Z(n48897) );
  NANDN U10683 ( .A(y[7546]), .B(x[7546]), .Z(n8898) );
  NANDN U10684 ( .A(y[7547]), .B(x[7547]), .Z(n48896) );
  NAND U10685 ( .A(n8898), .B(n48896), .Z(n60464) );
  XNOR U10686 ( .A(x[7544]), .B(y[7544]), .Z(n48887) );
  NANDN U10687 ( .A(y[7542]), .B(x[7542]), .Z(n8899) );
  NANDN U10688 ( .A(y[7543]), .B(x[7543]), .Z(n48886) );
  AND U10689 ( .A(n8899), .B(n48886), .Z(n60458) );
  XNOR U10690 ( .A(x[7542]), .B(y[7542]), .Z(n22331) );
  NANDN U10691 ( .A(x[7541]), .B(y[7541]), .Z(n22332) );
  AND U10692 ( .A(n22331), .B(n22332), .Z(n20847) );
  XNOR U10693 ( .A(x[7540]), .B(y[7540]), .Z(n48877) );
  NANDN U10694 ( .A(y[7538]), .B(x[7538]), .Z(n8900) );
  NANDN U10695 ( .A(y[7539]), .B(x[7539]), .Z(n48876) );
  AND U10696 ( .A(n8900), .B(n48876), .Z(n60454) );
  XNOR U10697 ( .A(x[7538]), .B(y[7538]), .Z(n22334) );
  ANDN U10698 ( .B(y[7537]), .A(x[7537]), .Z(n60452) );
  ANDN U10699 ( .B(n22334), .A(n60452), .Z(n20840) );
  XNOR U10700 ( .A(x[7536]), .B(y[7536]), .Z(n48867) );
  NANDN U10701 ( .A(y[7534]), .B(x[7534]), .Z(n8901) );
  NANDN U10702 ( .A(y[7535]), .B(x[7535]), .Z(n48866) );
  AND U10703 ( .A(n8901), .B(n48866), .Z(n60448) );
  ANDN U10704 ( .B(y[7533]), .A(x[7533]), .Z(n60446) );
  XNOR U10705 ( .A(x[7534]), .B(y[7534]), .Z(n22336) );
  NANDN U10706 ( .A(y[7532]), .B(x[7532]), .Z(n8902) );
  NANDN U10707 ( .A(y[7533]), .B(x[7533]), .Z(n22335) );
  NAND U10708 ( .A(n8902), .B(n22335), .Z(n60445) );
  ANDN U10709 ( .B(y[7529]), .A(x[7529]), .Z(n60442) );
  XNOR U10710 ( .A(x[7530]), .B(y[7530]), .Z(n22338) );
  NANDN U10711 ( .A(y[7528]), .B(x[7528]), .Z(n8903) );
  NANDN U10712 ( .A(y[7529]), .B(x[7529]), .Z(n22337) );
  AND U10713 ( .A(n8903), .B(n22337), .Z(n60441) );
  XNOR U10714 ( .A(x[7528]), .B(y[7528]), .Z(n48847) );
  NANDN U10715 ( .A(x[7527]), .B(y[7527]), .Z(n50700) );
  AND U10716 ( .A(n48847), .B(n50700), .Z(n20823) );
  XNOR U10717 ( .A(x[7526]), .B(y[7526]), .Z(n22340) );
  NANDN U10718 ( .A(y[7524]), .B(x[7524]), .Z(n8904) );
  NANDN U10719 ( .A(y[7525]), .B(x[7525]), .Z(n22339) );
  AND U10720 ( .A(n8904), .B(n22339), .Z(n60437) );
  XNOR U10721 ( .A(x[7524]), .B(y[7524]), .Z(n48837) );
  NANDN U10722 ( .A(x[7523]), .B(y[7523]), .Z(n60434) );
  AND U10723 ( .A(n48837), .B(n60434), .Z(n20816) );
  XNOR U10724 ( .A(x[7522]), .B(y[7522]), .Z(n22342) );
  NANDN U10725 ( .A(y[7520]), .B(x[7520]), .Z(n8905) );
  NANDN U10726 ( .A(y[7521]), .B(x[7521]), .Z(n22341) );
  AND U10727 ( .A(n8905), .B(n22341), .Z(n60430) );
  XNOR U10728 ( .A(x[7520]), .B(y[7520]), .Z(n48827) );
  NANDN U10729 ( .A(y[7518]), .B(x[7518]), .Z(n8906) );
  NANDN U10730 ( .A(y[7519]), .B(x[7519]), .Z(n48826) );
  AND U10731 ( .A(n8906), .B(n48826), .Z(n60427) );
  ANDN U10732 ( .B(y[7517]), .A(x[7517]), .Z(n50702) );
  XNOR U10733 ( .A(x[7518]), .B(y[7518]), .Z(n22344) );
  NANDN U10734 ( .A(y[7516]), .B(x[7516]), .Z(n8907) );
  NANDN U10735 ( .A(y[7517]), .B(x[7517]), .Z(n22343) );
  AND U10736 ( .A(n8907), .B(n22343), .Z(n60426) );
  XNOR U10737 ( .A(x[7516]), .B(y[7516]), .Z(n48817) );
  NANDN U10738 ( .A(y[7514]), .B(x[7514]), .Z(n8908) );
  NANDN U10739 ( .A(y[7515]), .B(x[7515]), .Z(n48816) );
  NAND U10740 ( .A(n8908), .B(n48816), .Z(n60423) );
  NANDN U10741 ( .A(x[7511]), .B(y[7511]), .Z(n48803) );
  IV U10742 ( .A(n48803), .Z(n60419) );
  XNOR U10743 ( .A(x[7512]), .B(y[7512]), .Z(n48807) );
  NANDN U10744 ( .A(y[7510]), .B(x[7510]), .Z(n8909) );
  NANDN U10745 ( .A(y[7511]), .B(x[7511]), .Z(n48806) );
  NAND U10746 ( .A(n8909), .B(n48806), .Z(n60417) );
  XNOR U10747 ( .A(x[7510]), .B(y[7510]), .Z(n22348) );
  ANDN U10748 ( .B(y[7509]), .A(x[7509]), .Z(n50705) );
  ANDN U10749 ( .B(n22348), .A(n50705), .Z(n20793) );
  NANDN U10750 ( .A(y[7508]), .B(x[7508]), .Z(n8910) );
  NANDN U10751 ( .A(y[7509]), .B(x[7509]), .Z(n22347) );
  NAND U10752 ( .A(n8910), .B(n22347), .Z(n60416) );
  XNOR U10753 ( .A(x[7508]), .B(y[7508]), .Z(n48796) );
  NANDN U10754 ( .A(y[7506]), .B(x[7506]), .Z(n8911) );
  NANDN U10755 ( .A(y[7507]), .B(x[7507]), .Z(n48795) );
  AND U10756 ( .A(n8911), .B(n48795), .Z(n60413) );
  ANDN U10757 ( .B(y[7505]), .A(x[7505]), .Z(n60411) );
  XNOR U10758 ( .A(x[7506]), .B(y[7506]), .Z(n22350) );
  NANDN U10759 ( .A(n60411), .B(n22350), .Z(n20787) );
  NANDN U10760 ( .A(y[7504]), .B(x[7504]), .Z(n8912) );
  NANDN U10761 ( .A(y[7505]), .B(x[7505]), .Z(n22349) );
  AND U10762 ( .A(n8912), .B(n22349), .Z(n60410) );
  XNOR U10763 ( .A(x[7504]), .B(y[7504]), .Z(n48786) );
  NANDN U10764 ( .A(x[7503]), .B(y[7503]), .Z(n60408) );
  NAND U10765 ( .A(n48786), .B(n60408), .Z(n20784) );
  ANDN U10766 ( .B(y[7501]), .A(x[7501]), .Z(n50708) );
  XNOR U10767 ( .A(x[7502]), .B(y[7502]), .Z(n22352) );
  NANDN U10768 ( .A(y[7500]), .B(x[7500]), .Z(n8913) );
  NANDN U10769 ( .A(y[7501]), .B(x[7501]), .Z(n22351) );
  NAND U10770 ( .A(n8913), .B(n22351), .Z(n60406) );
  NANDN U10771 ( .A(y[7498]), .B(x[7498]), .Z(n8914) );
  NANDN U10772 ( .A(y[7499]), .B(x[7499]), .Z(n48775) );
  AND U10773 ( .A(n8914), .B(n48775), .Z(n60403) );
  XNOR U10774 ( .A(x[7498]), .B(y[7498]), .Z(n22354) );
  NANDN U10775 ( .A(y[7496]), .B(x[7496]), .Z(n22355) );
  NANDN U10776 ( .A(y[7497]), .B(x[7497]), .Z(n22353) );
  NAND U10777 ( .A(n22355), .B(n22353), .Z(n60402) );
  NANDN U10778 ( .A(x[7495]), .B(y[7495]), .Z(n22357) );
  NANDN U10779 ( .A(x[7496]), .B(y[7496]), .Z(n48769) );
  AND U10780 ( .A(n22357), .B(n48769), .Z(n60401) );
  NANDN U10781 ( .A(x[7493]), .B(y[7493]), .Z(n22361) );
  NANDN U10782 ( .A(x[7494]), .B(y[7494]), .Z(n22358) );
  AND U10783 ( .A(n22361), .B(n22358), .Z(n60399) );
  NANDN U10784 ( .A(y[7492]), .B(x[7492]), .Z(n22363) );
  NANDN U10785 ( .A(y[7493]), .B(x[7493]), .Z(n22360) );
  AND U10786 ( .A(n22363), .B(n22360), .Z(n60398) );
  NANDN U10787 ( .A(x[7491]), .B(y[7491]), .Z(n22365) );
  NANDN U10788 ( .A(x[7492]), .B(y[7492]), .Z(n22362) );
  AND U10789 ( .A(n22365), .B(n22362), .Z(n60397) );
  NANDN U10790 ( .A(y[7490]), .B(x[7490]), .Z(n22367) );
  NANDN U10791 ( .A(y[7491]), .B(x[7491]), .Z(n22364) );
  NAND U10792 ( .A(n22367), .B(n22364), .Z(n60396) );
  NANDN U10793 ( .A(x[7490]), .B(y[7490]), .Z(n22366) );
  ANDN U10794 ( .B(y[7489]), .A(x[7489]), .Z(n48751) );
  ANDN U10795 ( .B(n22366), .A(n48751), .Z(n60395) );
  NANDN U10796 ( .A(x[7487]), .B(y[7487]), .Z(n22371) );
  NANDN U10797 ( .A(x[7488]), .B(y[7488]), .Z(n48752) );
  AND U10798 ( .A(n22371), .B(n48752), .Z(n60393) );
  NANDN U10799 ( .A(y[7486]), .B(x[7486]), .Z(n22373) );
  NANDN U10800 ( .A(y[7487]), .B(x[7487]), .Z(n22370) );
  AND U10801 ( .A(n22373), .B(n22370), .Z(n60392) );
  NANDN U10802 ( .A(x[7485]), .B(y[7485]), .Z(n22375) );
  NANDN U10803 ( .A(x[7486]), .B(y[7486]), .Z(n22372) );
  AND U10804 ( .A(n22375), .B(n22372), .Z(n60390) );
  NANDN U10805 ( .A(x[7483]), .B(y[7483]), .Z(n48737) );
  NANDN U10806 ( .A(x[7484]), .B(y[7484]), .Z(n22376) );
  AND U10807 ( .A(n48737), .B(n22376), .Z(n60388) );
  XNOR U10808 ( .A(x[7482]), .B(y[7482]), .Z(n22380) );
  NANDN U10809 ( .A(y[7480]), .B(x[7480]), .Z(n8915) );
  NANDN U10810 ( .A(y[7481]), .B(x[7481]), .Z(n22379) );
  NAND U10811 ( .A(n8915), .B(n22379), .Z(n50714) );
  XNOR U10812 ( .A(x[7480]), .B(y[7480]), .Z(n22382) );
  NANDN U10813 ( .A(x[7479]), .B(y[7479]), .Z(n50715) );
  AND U10814 ( .A(n22382), .B(n50715), .Z(n20753) );
  NANDN U10815 ( .A(x[7478]), .B(y[7478]), .Z(n22383) );
  ANDN U10816 ( .B(y[7477]), .A(x[7477]), .Z(n22386) );
  ANDN U10817 ( .B(n22383), .A(n22386), .Z(n60385) );
  XNOR U10818 ( .A(x[7476]), .B(y[7476]), .Z(n48722) );
  NANDN U10819 ( .A(y[7474]), .B(x[7474]), .Z(n8916) );
  NANDN U10820 ( .A(y[7475]), .B(x[7475]), .Z(n48721) );
  NAND U10821 ( .A(n8916), .B(n48721), .Z(n60384) );
  NANDN U10822 ( .A(y[7472]), .B(x[7472]), .Z(n8917) );
  NANDN U10823 ( .A(y[7473]), .B(x[7473]), .Z(n22387) );
  AND U10824 ( .A(n8917), .B(n22387), .Z(n60380) );
  NANDN U10825 ( .A(x[7471]), .B(y[7471]), .Z(n48708) );
  IV U10826 ( .A(n48708), .Z(n50721) );
  XNOR U10827 ( .A(x[7472]), .B(y[7472]), .Z(n48712) );
  NANDN U10828 ( .A(y[7470]), .B(x[7470]), .Z(n8918) );
  NANDN U10829 ( .A(y[7471]), .B(x[7471]), .Z(n48711) );
  NAND U10830 ( .A(n8918), .B(n48711), .Z(n60379) );
  XNOR U10831 ( .A(x[7470]), .B(y[7470]), .Z(n22390) );
  ANDN U10832 ( .B(y[7469]), .A(x[7469]), .Z(n22391) );
  NANDN U10833 ( .A(y[7469]), .B(x[7469]), .Z(n22389) );
  ANDN U10834 ( .B(x[7468]), .A(y[7468]), .Z(n48701) );
  ANDN U10835 ( .B(n22389), .A(n48701), .Z(n60376) );
  NANDN U10836 ( .A(x[7467]), .B(y[7467]), .Z(n48699) );
  NANDN U10837 ( .A(x[7468]), .B(y[7468]), .Z(n22392) );
  AND U10838 ( .A(n48699), .B(n22392), .Z(n60375) );
  NANDN U10839 ( .A(y[7466]), .B(x[7466]), .Z(n8919) );
  ANDN U10840 ( .B(x[7467]), .A(y[7467]), .Z(n48703) );
  ANDN U10841 ( .B(n8919), .A(n48703), .Z(n60374) );
  XNOR U10842 ( .A(y[7466]), .B(x[7466]), .Z(n22394) );
  NANDN U10843 ( .A(x[7465]), .B(y[7465]), .Z(n22395) );
  NAND U10844 ( .A(n22394), .B(n22395), .Z(n50722) );
  NANDN U10845 ( .A(y[7464]), .B(x[7464]), .Z(n8920) );
  NANDN U10846 ( .A(y[7465]), .B(x[7465]), .Z(n22393) );
  AND U10847 ( .A(n8920), .B(n22393), .Z(n60373) );
  XNOR U10848 ( .A(x[7464]), .B(y[7464]), .Z(n22397) );
  NANDN U10849 ( .A(y[7462]), .B(x[7462]), .Z(n8921) );
  NANDN U10850 ( .A(y[7463]), .B(x[7463]), .Z(n22396) );
  AND U10851 ( .A(n8921), .B(n22396), .Z(n60370) );
  XNOR U10852 ( .A(x[7462]), .B(y[7462]), .Z(n22400) );
  NANDN U10853 ( .A(y[7460]), .B(x[7460]), .Z(n8922) );
  NANDN U10854 ( .A(y[7461]), .B(x[7461]), .Z(n22399) );
  NAND U10855 ( .A(n8922), .B(n22399), .Z(n60367) );
  NANDN U10856 ( .A(y[7458]), .B(x[7458]), .Z(n8923) );
  NANDN U10857 ( .A(y[7459]), .B(x[7459]), .Z(n48680) );
  AND U10858 ( .A(n8923), .B(n48680), .Z(n60364) );
  ANDN U10859 ( .B(y[7457]), .A(x[7457]), .Z(n60362) );
  XNOR U10860 ( .A(x[7458]), .B(y[7458]), .Z(n22402) );
  NANDN U10861 ( .A(y[7456]), .B(x[7456]), .Z(n8924) );
  NANDN U10862 ( .A(y[7457]), .B(x[7457]), .Z(n22401) );
  NAND U10863 ( .A(n8924), .B(n22401), .Z(n60361) );
  XNOR U10864 ( .A(x[7456]), .B(y[7456]), .Z(n48671) );
  NANDN U10865 ( .A(x[7455]), .B(y[7455]), .Z(n60360) );
  NANDN U10866 ( .A(y[7454]), .B(x[7454]), .Z(n8925) );
  NANDN U10867 ( .A(y[7455]), .B(x[7455]), .Z(n48670) );
  AND U10868 ( .A(n8925), .B(n48670), .Z(n60358) );
  NANDN U10869 ( .A(y[7452]), .B(x[7452]), .Z(n8926) );
  NANDN U10870 ( .A(y[7453]), .B(x[7453]), .Z(n22403) );
  AND U10871 ( .A(n8926), .B(n22403), .Z(n60355) );
  NANDN U10872 ( .A(x[7451]), .B(y[7451]), .Z(n60353) );
  XNOR U10873 ( .A(x[7452]), .B(y[7452]), .Z(n48661) );
  AND U10874 ( .A(n60353), .B(n48661), .Z(n20713) );
  XNOR U10875 ( .A(y[7450]), .B(x[7450]), .Z(n22406) );
  ANDN U10876 ( .B(y[7449]), .A(x[7449]), .Z(n22407) );
  ANDN U10877 ( .B(n22406), .A(n22407), .Z(n60350) );
  NANDN U10878 ( .A(y[7448]), .B(x[7448]), .Z(n8927) );
  NANDN U10879 ( .A(y[7449]), .B(x[7449]), .Z(n22405) );
  AND U10880 ( .A(n8927), .B(n22405), .Z(n60349) );
  XNOR U10881 ( .A(x[7448]), .B(y[7448]), .Z(n48650) );
  ANDN U10882 ( .B(y[7447]), .A(x[7447]), .Z(n48646) );
  ANDN U10883 ( .B(n48650), .A(n48646), .Z(n20707) );
  XNOR U10884 ( .A(x[7446]), .B(y[7446]), .Z(n22409) );
  ANDN U10885 ( .B(y[7445]), .A(x[7445]), .Z(n50726) );
  ANDN U10886 ( .B(n22409), .A(n50726), .Z(n20703) );
  XNOR U10887 ( .A(x[7444]), .B(y[7444]), .Z(n48639) );
  NANDN U10888 ( .A(y[7442]), .B(x[7442]), .Z(n8928) );
  NANDN U10889 ( .A(y[7443]), .B(x[7443]), .Z(n48638) );
  AND U10890 ( .A(n8928), .B(n48638), .Z(n60343) );
  XNOR U10891 ( .A(x[7442]), .B(y[7442]), .Z(n22411) );
  ANDN U10892 ( .B(y[7441]), .A(x[7441]), .Z(n50729) );
  ANDN U10893 ( .B(n22411), .A(n50729), .Z(n20696) );
  XNOR U10894 ( .A(x[7440]), .B(y[7440]), .Z(n48629) );
  NANDN U10895 ( .A(y[7438]), .B(x[7438]), .Z(n8929) );
  NANDN U10896 ( .A(y[7439]), .B(x[7439]), .Z(n48628) );
  AND U10897 ( .A(n8929), .B(n48628), .Z(n60339) );
  XNOR U10898 ( .A(x[7438]), .B(y[7438]), .Z(n22413) );
  NANDN U10899 ( .A(y[7436]), .B(x[7436]), .Z(n8930) );
  NANDN U10900 ( .A(y[7437]), .B(x[7437]), .Z(n22412) );
  NAND U10901 ( .A(n8930), .B(n22412), .Z(n60335) );
  NANDN U10902 ( .A(y[7434]), .B(x[7434]), .Z(n8931) );
  NANDN U10903 ( .A(y[7435]), .B(x[7435]), .Z(n22414) );
  AND U10904 ( .A(n8931), .B(n22414), .Z(n60332) );
  ANDN U10905 ( .B(y[7433]), .A(x[7433]), .Z(n60330) );
  XNOR U10906 ( .A(x[7434]), .B(y[7434]), .Z(n22417) );
  NANDN U10907 ( .A(y[7432]), .B(x[7432]), .Z(n8932) );
  NANDN U10908 ( .A(y[7433]), .B(x[7433]), .Z(n22416) );
  NAND U10909 ( .A(n8932), .B(n22416), .Z(n60329) );
  XNOR U10910 ( .A(x[7432]), .B(y[7432]), .Z(n48611) );
  NANDN U10911 ( .A(x[7431]), .B(y[7431]), .Z(n50731) );
  AND U10912 ( .A(n48611), .B(n50731), .Z(n20680) );
  NANDN U10913 ( .A(y[7430]), .B(x[7430]), .Z(n8933) );
  NANDN U10914 ( .A(y[7431]), .B(x[7431]), .Z(n48610) );
  NAND U10915 ( .A(n8933), .B(n48610), .Z(n60328) );
  XNOR U10916 ( .A(x[7430]), .B(y[7430]), .Z(n22419) );
  NANDN U10917 ( .A(y[7428]), .B(x[7428]), .Z(n8934) );
  NANDN U10918 ( .A(y[7429]), .B(x[7429]), .Z(n22418) );
  AND U10919 ( .A(n8934), .B(n22418), .Z(n60325) );
  XNOR U10920 ( .A(x[7428]), .B(y[7428]), .Z(n22421) );
  ANDN U10921 ( .B(y[7427]), .A(x[7427]), .Z(n48599) );
  ANDN U10922 ( .B(n22421), .A(n48599), .Z(n20674) );
  XNOR U10923 ( .A(x[7426]), .B(y[7426]), .Z(n22423) );
  NANDN U10924 ( .A(y[7424]), .B(x[7424]), .Z(n8935) );
  NANDN U10925 ( .A(y[7425]), .B(x[7425]), .Z(n22422) );
  AND U10926 ( .A(n8935), .B(n22422), .Z(n60321) );
  XNOR U10927 ( .A(x[7424]), .B(y[7424]), .Z(n22425) );
  NANDN U10928 ( .A(y[7422]), .B(x[7422]), .Z(n8936) );
  NANDN U10929 ( .A(y[7423]), .B(x[7423]), .Z(n22424) );
  NAND U10930 ( .A(n8936), .B(n22424), .Z(n60318) );
  XNOR U10931 ( .A(x[7420]), .B(y[7420]), .Z(n48584) );
  NANDN U10932 ( .A(y[7418]), .B(x[7418]), .Z(n8937) );
  NANDN U10933 ( .A(y[7419]), .B(x[7419]), .Z(n48583) );
  NAND U10934 ( .A(n8937), .B(n48583), .Z(n60315) );
  XNOR U10935 ( .A(x[7418]), .B(y[7418]), .Z(n22429) );
  NANDN U10936 ( .A(x[7417]), .B(y[7417]), .Z(n60313) );
  AND U10937 ( .A(n22429), .B(n60313), .Z(n20657) );
  XNOR U10938 ( .A(y[7416]), .B(x[7416]), .Z(n48574) );
  NANDN U10939 ( .A(y[7414]), .B(x[7414]), .Z(n8938) );
  ANDN U10940 ( .B(x[7415]), .A(y[7415]), .Z(n48576) );
  ANDN U10941 ( .B(n8938), .A(n48576), .Z(n60310) );
  XNOR U10942 ( .A(x[7414]), .B(y[7414]), .Z(n22431) );
  ANDN U10943 ( .B(y[7413]), .A(x[7413]), .Z(n60307) );
  ANDN U10944 ( .B(n22431), .A(n60307), .Z(n20650) );
  XNOR U10945 ( .A(x[7412]), .B(y[7412]), .Z(n48564) );
  NANDN U10946 ( .A(y[7410]), .B(x[7410]), .Z(n8939) );
  NANDN U10947 ( .A(y[7411]), .B(x[7411]), .Z(n48563) );
  AND U10948 ( .A(n8939), .B(n48563), .Z(n60303) );
  XNOR U10949 ( .A(x[7410]), .B(y[7410]), .Z(n22433) );
  ANDN U10950 ( .B(y[7409]), .A(x[7409]), .Z(n60301) );
  ANDN U10951 ( .B(n22433), .A(n60301), .Z(n20643) );
  XNOR U10952 ( .A(x[7408]), .B(y[7408]), .Z(n48554) );
  NANDN U10953 ( .A(y[7406]), .B(x[7406]), .Z(n8940) );
  NANDN U10954 ( .A(y[7407]), .B(x[7407]), .Z(n48553) );
  AND U10955 ( .A(n8940), .B(n48553), .Z(n60299) );
  ANDN U10956 ( .B(y[7405]), .A(x[7405]), .Z(n60297) );
  XNOR U10957 ( .A(x[7406]), .B(y[7406]), .Z(n22435) );
  NANDN U10958 ( .A(y[7404]), .B(x[7404]), .Z(n8941) );
  NANDN U10959 ( .A(y[7405]), .B(x[7405]), .Z(n22434) );
  NAND U10960 ( .A(n8941), .B(n22434), .Z(n60296) );
  XNOR U10961 ( .A(x[7404]), .B(y[7404]), .Z(n48544) );
  NANDN U10962 ( .A(y[7402]), .B(x[7402]), .Z(n8942) );
  NANDN U10963 ( .A(y[7403]), .B(x[7403]), .Z(n48543) );
  NAND U10964 ( .A(n8942), .B(n48543), .Z(n60291) );
  XNOR U10965 ( .A(x[7402]), .B(y[7402]), .Z(n22437) );
  ANDN U10966 ( .B(y[7401]), .A(x[7401]), .Z(n60289) );
  NANDN U10967 ( .A(y[7400]), .B(x[7400]), .Z(n8943) );
  NANDN U10968 ( .A(y[7401]), .B(x[7401]), .Z(n22436) );
  AND U10969 ( .A(n8943), .B(n22436), .Z(n60288) );
  XNOR U10970 ( .A(x[7400]), .B(y[7400]), .Z(n48534) );
  NANDN U10971 ( .A(x[7399]), .B(y[7399]), .Z(n60286) );
  NAND U10972 ( .A(n48534), .B(n60286), .Z(n20627) );
  NANDN U10973 ( .A(y[7398]), .B(x[7398]), .Z(n8944) );
  NANDN U10974 ( .A(y[7399]), .B(x[7399]), .Z(n48533) );
  AND U10975 ( .A(n8944), .B(n48533), .Z(n50742) );
  NANDN U10976 ( .A(x[7397]), .B(y[7397]), .Z(n60285) );
  XNOR U10977 ( .A(x[7398]), .B(y[7398]), .Z(n22439) );
  NAND U10978 ( .A(n60285), .B(n22439), .Z(n20624) );
  NANDN U10979 ( .A(y[7396]), .B(x[7396]), .Z(n22441) );
  NANDN U10980 ( .A(y[7397]), .B(x[7397]), .Z(n22438) );
  AND U10981 ( .A(n22441), .B(n22438), .Z(n60283) );
  NANDN U10982 ( .A(x[7395]), .B(y[7395]), .Z(n22443) );
  NANDN U10983 ( .A(x[7396]), .B(y[7396]), .Z(n22440) );
  AND U10984 ( .A(n22443), .B(n22440), .Z(n60282) );
  NANDN U10985 ( .A(y[7394]), .B(x[7394]), .Z(n8945) );
  NANDN U10986 ( .A(y[7395]), .B(x[7395]), .Z(n22442) );
  AND U10987 ( .A(n8945), .B(n22442), .Z(n60281) );
  XNOR U10988 ( .A(x[7394]), .B(y[7394]), .Z(n22445) );
  NANDN U10989 ( .A(x[7393]), .B(y[7393]), .Z(n50743) );
  AND U10990 ( .A(n22445), .B(n50743), .Z(n20619) );
  NANDN U10991 ( .A(y[7390]), .B(x[7390]), .Z(n8946) );
  NANDN U10992 ( .A(y[7391]), .B(x[7391]), .Z(n22448) );
  AND U10993 ( .A(n8946), .B(n22448), .Z(n60277) );
  XNOR U10994 ( .A(x[7390]), .B(y[7390]), .Z(n22450) );
  ANDN U10995 ( .B(y[7389]), .A(x[7389]), .Z(n60275) );
  ANDN U10996 ( .B(n22450), .A(n60275), .Z(n20614) );
  XNOR U10997 ( .A(x[7388]), .B(y[7388]), .Z(n48507) );
  NANDN U10998 ( .A(y[7386]), .B(x[7386]), .Z(n8947) );
  NANDN U10999 ( .A(y[7387]), .B(x[7387]), .Z(n48506) );
  AND U11000 ( .A(n8947), .B(n48506), .Z(n60274) );
  ANDN U11001 ( .B(y[7385]), .A(x[7385]), .Z(n60272) );
  XNOR U11002 ( .A(x[7386]), .B(y[7386]), .Z(n22452) );
  NANDN U11003 ( .A(y[7384]), .B(x[7384]), .Z(n8948) );
  NANDN U11004 ( .A(y[7385]), .B(x[7385]), .Z(n22451) );
  AND U11005 ( .A(n8948), .B(n22451), .Z(n60271) );
  XNOR U11006 ( .A(x[7384]), .B(y[7384]), .Z(n48497) );
  NANDN U11007 ( .A(y[7382]), .B(x[7382]), .Z(n22454) );
  NANDN U11008 ( .A(y[7383]), .B(x[7383]), .Z(n48496) );
  AND U11009 ( .A(n22454), .B(n48496), .Z(n60270) );
  NANDN U11010 ( .A(x[7381]), .B(y[7381]), .Z(n22456) );
  NANDN U11011 ( .A(x[7382]), .B(y[7382]), .Z(n22453) );
  AND U11012 ( .A(n22456), .B(n22453), .Z(n60269) );
  NANDN U11013 ( .A(y[7380]), .B(x[7380]), .Z(n8949) );
  NANDN U11014 ( .A(y[7381]), .B(x[7381]), .Z(n22455) );
  AND U11015 ( .A(n8949), .B(n22455), .Z(n60268) );
  XNOR U11016 ( .A(x[7380]), .B(y[7380]), .Z(n22458) );
  NANDN U11017 ( .A(x[7379]), .B(y[7379]), .Z(n60265) );
  AND U11018 ( .A(n22458), .B(n60265), .Z(n20599) );
  XNOR U11019 ( .A(x[7378]), .B(y[7378]), .Z(n22460) );
  NANDN U11020 ( .A(y[7376]), .B(x[7376]), .Z(n8950) );
  NANDN U11021 ( .A(y[7377]), .B(x[7377]), .Z(n22459) );
  AND U11022 ( .A(n8950), .B(n22459), .Z(n60262) );
  XNOR U11023 ( .A(x[7376]), .B(y[7376]), .Z(n48479) );
  NANDN U11024 ( .A(x[7375]), .B(y[7375]), .Z(n50751) );
  AND U11025 ( .A(n48479), .B(n50751), .Z(n20592) );
  XNOR U11026 ( .A(x[7374]), .B(y[7374]), .Z(n22463) );
  NANDN U11027 ( .A(y[7372]), .B(x[7372]), .Z(n8951) );
  NANDN U11028 ( .A(y[7373]), .B(x[7373]), .Z(n22462) );
  AND U11029 ( .A(n8951), .B(n22462), .Z(n60260) );
  XNOR U11030 ( .A(x[7372]), .B(y[7372]), .Z(n48469) );
  ANDN U11031 ( .B(y[7371]), .A(x[7371]), .Z(n48465) );
  ANDN U11032 ( .B(n48469), .A(n48465), .Z(n20585) );
  XNOR U11033 ( .A(x[7370]), .B(y[7370]), .Z(n22465) );
  NANDN U11034 ( .A(y[7368]), .B(x[7368]), .Z(n8952) );
  NANDN U11035 ( .A(y[7369]), .B(x[7369]), .Z(n22464) );
  AND U11036 ( .A(n8952), .B(n22464), .Z(n60254) );
  XNOR U11037 ( .A(x[7368]), .B(y[7368]), .Z(n48458) );
  NANDN U11038 ( .A(y[7366]), .B(x[7366]), .Z(n8953) );
  NANDN U11039 ( .A(y[7367]), .B(x[7367]), .Z(n48457) );
  NAND U11040 ( .A(n8953), .B(n48457), .Z(n60253) );
  ANDN U11041 ( .B(y[7365]), .A(x[7365]), .Z(n60251) );
  XNOR U11042 ( .A(x[7366]), .B(y[7366]), .Z(n22467) );
  NANDN U11043 ( .A(y[7364]), .B(x[7364]), .Z(n8954) );
  NANDN U11044 ( .A(y[7365]), .B(x[7365]), .Z(n22466) );
  AND U11045 ( .A(n8954), .B(n22466), .Z(n60250) );
  XNOR U11046 ( .A(y[7364]), .B(x[7364]), .Z(n48448) );
  NANDN U11047 ( .A(x[7363]), .B(y[7363]), .Z(n48444) );
  AND U11048 ( .A(n48448), .B(n48444), .Z(n60249) );
  NANDN U11049 ( .A(y[7362]), .B(x[7362]), .Z(n8955) );
  NANDN U11050 ( .A(y[7363]), .B(x[7363]), .Z(n48447) );
  NAND U11051 ( .A(n8955), .B(n48447), .Z(n50759) );
  XNOR U11052 ( .A(x[7362]), .B(y[7362]), .Z(n22470) );
  NANDN U11053 ( .A(x[7361]), .B(y[7361]), .Z(n60247) );
  AND U11054 ( .A(n22470), .B(n60247), .Z(n20570) );
  XNOR U11055 ( .A(x[7360]), .B(y[7360]), .Z(n22472) );
  NANDN U11056 ( .A(y[7358]), .B(x[7358]), .Z(n8956) );
  NANDN U11057 ( .A(y[7359]), .B(x[7359]), .Z(n22471) );
  AND U11058 ( .A(n8956), .B(n22471), .Z(n60243) );
  XNOR U11059 ( .A(x[7358]), .B(y[7358]), .Z(n22474) );
  NANDN U11060 ( .A(x[7357]), .B(y[7357]), .Z(n60241) );
  AND U11061 ( .A(n22474), .B(n60241), .Z(n20563) );
  XNOR U11062 ( .A(x[7356]), .B(y[7356]), .Z(n48429) );
  NANDN U11063 ( .A(y[7354]), .B(x[7354]), .Z(n8957) );
  NANDN U11064 ( .A(y[7355]), .B(x[7355]), .Z(n48428) );
  AND U11065 ( .A(n8957), .B(n48428), .Z(n60236) );
  XNOR U11066 ( .A(x[7354]), .B(y[7354]), .Z(n22476) );
  ANDN U11067 ( .B(y[7353]), .A(x[7353]), .Z(n50761) );
  ANDN U11068 ( .B(n22476), .A(n50761), .Z(n20556) );
  XNOR U11069 ( .A(x[7352]), .B(y[7352]), .Z(n48419) );
  NANDN U11070 ( .A(y[7350]), .B(x[7350]), .Z(n8958) );
  NANDN U11071 ( .A(y[7351]), .B(x[7351]), .Z(n48418) );
  AND U11072 ( .A(n8958), .B(n48418), .Z(n60232) );
  XNOR U11073 ( .A(x[7350]), .B(y[7350]), .Z(n22478) );
  NANDN U11074 ( .A(y[7348]), .B(x[7348]), .Z(n8959) );
  NANDN U11075 ( .A(y[7349]), .B(x[7349]), .Z(n22477) );
  AND U11076 ( .A(n8959), .B(n22477), .Z(n50762) );
  ANDN U11077 ( .B(y[7345]), .A(x[7345]), .Z(n60226) );
  XNOR U11078 ( .A(x[7346]), .B(y[7346]), .Z(n22484) );
  NANDN U11079 ( .A(y[7344]), .B(x[7344]), .Z(n8960) );
  NANDN U11080 ( .A(y[7345]), .B(x[7345]), .Z(n22483) );
  AND U11081 ( .A(n8960), .B(n22483), .Z(n60225) );
  XNOR U11082 ( .A(x[7344]), .B(y[7344]), .Z(n48401) );
  NANDN U11083 ( .A(x[7343]), .B(y[7343]), .Z(n50764) );
  AND U11084 ( .A(n48401), .B(n50764), .Z(n20540) );
  XNOR U11085 ( .A(x[7342]), .B(y[7342]), .Z(n22486) );
  NANDN U11086 ( .A(y[7340]), .B(x[7340]), .Z(n8961) );
  NANDN U11087 ( .A(y[7341]), .B(x[7341]), .Z(n22485) );
  AND U11088 ( .A(n8961), .B(n22485), .Z(n60221) );
  XNOR U11089 ( .A(x[7340]), .B(y[7340]), .Z(n22488) );
  NANDN U11090 ( .A(x[7339]), .B(y[7339]), .Z(n60219) );
  AND U11091 ( .A(n22488), .B(n60219), .Z(n20533) );
  XNOR U11092 ( .A(x[7338]), .B(y[7338]), .Z(n22490) );
  NANDN U11093 ( .A(y[7336]), .B(x[7336]), .Z(n8962) );
  NANDN U11094 ( .A(y[7337]), .B(x[7337]), .Z(n22489) );
  AND U11095 ( .A(n8962), .B(n22489), .Z(n60214) );
  XNOR U11096 ( .A(x[7336]), .B(y[7336]), .Z(n48383) );
  ANDN U11097 ( .B(y[7335]), .A(x[7335]), .Z(n48379) );
  ANDN U11098 ( .B(n48383), .A(n48379), .Z(n20526) );
  XNOR U11099 ( .A(x[7334]), .B(y[7334]), .Z(n22492) );
  NANDN U11100 ( .A(y[7332]), .B(x[7332]), .Z(n8963) );
  NANDN U11101 ( .A(y[7333]), .B(x[7333]), .Z(n22491) );
  AND U11102 ( .A(n8963), .B(n22491), .Z(n60211) );
  XNOR U11103 ( .A(x[7332]), .B(y[7332]), .Z(n48372) );
  XNOR U11104 ( .A(x[7330]), .B(y[7330]), .Z(n22494) );
  XNOR U11105 ( .A(x[7328]), .B(y[7328]), .Z(n48362) );
  NANDN U11106 ( .A(y[7326]), .B(x[7326]), .Z(n8964) );
  NANDN U11107 ( .A(y[7327]), .B(x[7327]), .Z(n48361) );
  AND U11108 ( .A(n8964), .B(n48361), .Z(n60204) );
  NANDN U11109 ( .A(y[7324]), .B(x[7324]), .Z(n8965) );
  NANDN U11110 ( .A(y[7325]), .B(x[7325]), .Z(n22496) );
  AND U11111 ( .A(n8965), .B(n22496), .Z(n60200) );
  XNOR U11112 ( .A(x[7324]), .B(y[7324]), .Z(n48352) );
  XNOR U11113 ( .A(x[7322]), .B(y[7322]), .Z(n22499) );
  ANDN U11114 ( .B(y[7321]), .A(x[7321]), .Z(n60196) );
  ANDN U11115 ( .B(n22499), .A(n60196), .Z(n20501) );
  XNOR U11116 ( .A(x[7320]), .B(y[7320]), .Z(n48342) );
  NANDN U11117 ( .A(y[7318]), .B(x[7318]), .Z(n8966) );
  NANDN U11118 ( .A(y[7319]), .B(x[7319]), .Z(n48341) );
  AND U11119 ( .A(n8966), .B(n48341), .Z(n60194) );
  XNOR U11120 ( .A(x[7318]), .B(y[7318]), .Z(n22501) );
  ANDN U11121 ( .B(y[7317]), .A(x[7317]), .Z(n22502) );
  ANDN U11122 ( .B(n22501), .A(n22502), .Z(n20494) );
  XNOR U11123 ( .A(x[7316]), .B(y[7316]), .Z(n22504) );
  NANDN U11124 ( .A(y[7314]), .B(x[7314]), .Z(n8967) );
  NANDN U11125 ( .A(y[7315]), .B(x[7315]), .Z(n22503) );
  AND U11126 ( .A(n8967), .B(n22503), .Z(n60190) );
  XNOR U11127 ( .A(x[7314]), .B(y[7314]), .Z(n22506) );
  NANDN U11128 ( .A(y[7312]), .B(x[7312]), .Z(n8968) );
  NANDN U11129 ( .A(y[7313]), .B(x[7313]), .Z(n22505) );
  AND U11130 ( .A(n8968), .B(n22505), .Z(n60186) );
  NANDN U11131 ( .A(y[7310]), .B(x[7310]), .Z(n8969) );
  ANDN U11132 ( .B(x[7311]), .A(y[7311]), .Z(n48326) );
  ANDN U11133 ( .B(n8969), .A(n48326), .Z(n60183) );
  XNOR U11134 ( .A(x[7310]), .B(y[7310]), .Z(n22508) );
  NANDN U11135 ( .A(y[7308]), .B(x[7308]), .Z(n8970) );
  NANDN U11136 ( .A(y[7309]), .B(x[7309]), .Z(n22507) );
  AND U11137 ( .A(n8970), .B(n22507), .Z(n60180) );
  XNOR U11138 ( .A(x[7308]), .B(y[7308]), .Z(n48314) );
  NANDN U11139 ( .A(x[7307]), .B(y[7307]), .Z(n60178) );
  AND U11140 ( .A(n48314), .B(n60178), .Z(n20478) );
  NANDN U11141 ( .A(y[7306]), .B(x[7306]), .Z(n8971) );
  NANDN U11142 ( .A(y[7307]), .B(x[7307]), .Z(n48313) );
  NAND U11143 ( .A(n8971), .B(n48313), .Z(n60177) );
  XNOR U11144 ( .A(x[7306]), .B(y[7306]), .Z(n22510) );
  NANDN U11145 ( .A(y[7304]), .B(x[7304]), .Z(n8972) );
  NANDN U11146 ( .A(y[7305]), .B(x[7305]), .Z(n22509) );
  AND U11147 ( .A(n8972), .B(n22509), .Z(n60176) );
  XNOR U11148 ( .A(x[7304]), .B(y[7304]), .Z(n48304) );
  NANDN U11149 ( .A(x[7303]), .B(y[7303]), .Z(n60174) );
  NAND U11150 ( .A(n48304), .B(n60174), .Z(n20472) );
  NANDN U11151 ( .A(y[7302]), .B(x[7302]), .Z(n8973) );
  NANDN U11152 ( .A(y[7303]), .B(x[7303]), .Z(n48303) );
  AND U11153 ( .A(n8973), .B(n48303), .Z(n60173) );
  ANDN U11154 ( .B(y[7301]), .A(x[7301]), .Z(n50779) );
  XNOR U11155 ( .A(x[7302]), .B(y[7302]), .Z(n22512) );
  NANDN U11156 ( .A(n50779), .B(n22512), .Z(n20469) );
  NANDN U11157 ( .A(y[7300]), .B(x[7300]), .Z(n8974) );
  NANDN U11158 ( .A(y[7301]), .B(x[7301]), .Z(n22511) );
  AND U11159 ( .A(n8974), .B(n22511), .Z(n60171) );
  XNOR U11160 ( .A(x[7300]), .B(y[7300]), .Z(n48294) );
  NANDN U11161 ( .A(y[7298]), .B(x[7298]), .Z(n22514) );
  NANDN U11162 ( .A(y[7299]), .B(x[7299]), .Z(n48293) );
  NAND U11163 ( .A(n22514), .B(n48293), .Z(n60170) );
  NANDN U11164 ( .A(x[7297]), .B(y[7297]), .Z(n22516) );
  NANDN U11165 ( .A(x[7298]), .B(y[7298]), .Z(n22513) );
  AND U11166 ( .A(n22516), .B(n22513), .Z(n60169) );
  NANDN U11167 ( .A(y[7294]), .B(x[7294]), .Z(n8975) );
  NANDN U11168 ( .A(y[7295]), .B(x[7295]), .Z(n22519) );
  AND U11169 ( .A(n8975), .B(n22519), .Z(n60167) );
  ANDN U11170 ( .B(y[7293]), .A(x[7293]), .Z(n60166) );
  XNOR U11171 ( .A(x[7294]), .B(y[7294]), .Z(n22522) );
  NANDN U11172 ( .A(n60166), .B(n22522), .Z(n20459) );
  NANDN U11173 ( .A(y[7292]), .B(x[7292]), .Z(n8976) );
  NANDN U11174 ( .A(y[7293]), .B(x[7293]), .Z(n22521) );
  AND U11175 ( .A(n8976), .B(n22521), .Z(n60165) );
  NANDN U11176 ( .A(x[7291]), .B(y[7291]), .Z(n50784) );
  XNOR U11177 ( .A(x[7292]), .B(y[7292]), .Z(n48276) );
  NAND U11178 ( .A(n50784), .B(n48276), .Z(n20456) );
  NANDN U11179 ( .A(y[7290]), .B(x[7290]), .Z(n8977) );
  NANDN U11180 ( .A(y[7291]), .B(x[7291]), .Z(n48275) );
  AND U11181 ( .A(n8977), .B(n48275), .Z(n60164) );
  XNOR U11182 ( .A(x[7290]), .B(y[7290]), .Z(n22524) );
  NANDN U11183 ( .A(y[7288]), .B(x[7288]), .Z(n22526) );
  NANDN U11184 ( .A(y[7289]), .B(x[7289]), .Z(n22523) );
  AND U11185 ( .A(n22526), .B(n22523), .Z(n60160) );
  NANDN U11186 ( .A(x[7287]), .B(y[7287]), .Z(n22528) );
  NANDN U11187 ( .A(x[7288]), .B(y[7288]), .Z(n22525) );
  AND U11188 ( .A(n22528), .B(n22525), .Z(n60159) );
  NANDN U11189 ( .A(y[7286]), .B(x[7286]), .Z(n22530) );
  NANDN U11190 ( .A(y[7287]), .B(x[7287]), .Z(n22527) );
  NAND U11191 ( .A(n22530), .B(n22527), .Z(n60158) );
  NANDN U11192 ( .A(x[7285]), .B(y[7285]), .Z(n22532) );
  NANDN U11193 ( .A(x[7286]), .B(y[7286]), .Z(n22529) );
  AND U11194 ( .A(n22532), .B(n22529), .Z(n60157) );
  NANDN U11195 ( .A(y[7284]), .B(x[7284]), .Z(n8978) );
  NANDN U11196 ( .A(y[7285]), .B(x[7285]), .Z(n22531) );
  AND U11197 ( .A(n8978), .B(n22531), .Z(n60156) );
  XNOR U11198 ( .A(x[7284]), .B(y[7284]), .Z(n22534) );
  ANDN U11199 ( .B(y[7283]), .A(x[7283]), .Z(n48256) );
  ANDN U11200 ( .B(n22534), .A(n48256), .Z(n20446) );
  XNOR U11201 ( .A(x[7282]), .B(y[7282]), .Z(n22536) );
  NANDN U11202 ( .A(y[7280]), .B(x[7280]), .Z(n8979) );
  NANDN U11203 ( .A(y[7281]), .B(x[7281]), .Z(n22535) );
  AND U11204 ( .A(n8979), .B(n22535), .Z(n60152) );
  XNOR U11205 ( .A(x[7280]), .B(y[7280]), .Z(n48249) );
  NANDN U11206 ( .A(y[7278]), .B(x[7278]), .Z(n8980) );
  NANDN U11207 ( .A(y[7279]), .B(x[7279]), .Z(n48248) );
  AND U11208 ( .A(n8980), .B(n48248), .Z(n60149) );
  ANDN U11209 ( .B(y[7277]), .A(x[7277]), .Z(n60147) );
  XNOR U11210 ( .A(x[7278]), .B(y[7278]), .Z(n22539) );
  NANDN U11211 ( .A(y[7276]), .B(x[7276]), .Z(n8981) );
  NANDN U11212 ( .A(y[7277]), .B(x[7277]), .Z(n22538) );
  NAND U11213 ( .A(n8981), .B(n22538), .Z(n60146) );
  NANDN U11214 ( .A(y[7274]), .B(x[7274]), .Z(n8982) );
  NANDN U11215 ( .A(y[7275]), .B(x[7275]), .Z(n48238) );
  AND U11216 ( .A(n8982), .B(n48238), .Z(n60143) );
  XNOR U11217 ( .A(x[7274]), .B(y[7274]), .Z(n22541) );
  ANDN U11218 ( .B(y[7273]), .A(x[7273]), .Z(n60141) );
  ANDN U11219 ( .B(n22541), .A(n60141), .Z(n20430) );
  XNOR U11220 ( .A(x[7272]), .B(y[7272]), .Z(n48229) );
  NANDN U11221 ( .A(y[7270]), .B(x[7270]), .Z(n8983) );
  NANDN U11222 ( .A(y[7271]), .B(x[7271]), .Z(n48228) );
  AND U11223 ( .A(n8983), .B(n48228), .Z(n60139) );
  XNOR U11224 ( .A(x[7270]), .B(y[7270]), .Z(n22543) );
  ANDN U11225 ( .B(y[7269]), .A(x[7269]), .Z(n60137) );
  ANDN U11226 ( .B(n22543), .A(n60137), .Z(n20423) );
  XNOR U11227 ( .A(x[7268]), .B(y[7268]), .Z(n48219) );
  NANDN U11228 ( .A(y[7266]), .B(x[7266]), .Z(n8984) );
  NANDN U11229 ( .A(y[7267]), .B(x[7267]), .Z(n48218) );
  AND U11230 ( .A(n8984), .B(n48218), .Z(n60135) );
  ANDN U11231 ( .B(y[7265]), .A(x[7265]), .Z(n50794) );
  XNOR U11232 ( .A(x[7266]), .B(y[7266]), .Z(n22545) );
  NANDN U11233 ( .A(y[7264]), .B(x[7264]), .Z(n8985) );
  NANDN U11234 ( .A(y[7265]), .B(x[7265]), .Z(n22544) );
  NAND U11235 ( .A(n8985), .B(n22544), .Z(n60133) );
  XNOR U11236 ( .A(x[7264]), .B(y[7264]), .Z(n22547) );
  NANDN U11237 ( .A(y[7262]), .B(x[7262]), .Z(n8986) );
  NANDN U11238 ( .A(y[7263]), .B(x[7263]), .Z(n22546) );
  AND U11239 ( .A(n8986), .B(n22546), .Z(n60129) );
  XNOR U11240 ( .A(y[7262]), .B(x[7262]), .Z(n22549) );
  ANDN U11241 ( .B(y[7261]), .A(x[7261]), .Z(n22550) );
  ANDN U11242 ( .B(n22549), .A(n22550), .Z(n60128) );
  NANDN U11243 ( .A(y[7260]), .B(x[7260]), .Z(n8987) );
  NANDN U11244 ( .A(y[7261]), .B(x[7261]), .Z(n22548) );
  NAND U11245 ( .A(n8987), .B(n22548), .Z(n60127) );
  XNOR U11246 ( .A(x[7260]), .B(y[7260]), .Z(n48200) );
  NANDN U11247 ( .A(x[7259]), .B(y[7259]), .Z(n60125) );
  AND U11248 ( .A(n48200), .B(n60125), .Z(n20408) );
  XNOR U11249 ( .A(x[7258]), .B(y[7258]), .Z(n22552) );
  NANDN U11250 ( .A(y[7256]), .B(x[7256]), .Z(n8988) );
  NANDN U11251 ( .A(y[7257]), .B(x[7257]), .Z(n22551) );
  AND U11252 ( .A(n8988), .B(n22551), .Z(n60121) );
  XNOR U11253 ( .A(x[7256]), .B(y[7256]), .Z(n48190) );
  NANDN U11254 ( .A(x[7255]), .B(y[7255]), .Z(n60120) );
  AND U11255 ( .A(n48190), .B(n60120), .Z(n20401) );
  XNOR U11256 ( .A(x[7254]), .B(y[7254]), .Z(n22554) );
  NANDN U11257 ( .A(y[7252]), .B(x[7252]), .Z(n8989) );
  NANDN U11258 ( .A(y[7253]), .B(x[7253]), .Z(n22553) );
  AND U11259 ( .A(n8989), .B(n22553), .Z(n60115) );
  XNOR U11260 ( .A(x[7252]), .B(y[7252]), .Z(n48180) );
  ANDN U11261 ( .B(y[7251]), .A(x[7251]), .Z(n48176) );
  ANDN U11262 ( .B(n48180), .A(n48176), .Z(n20394) );
  XNOR U11263 ( .A(x[7250]), .B(y[7250]), .Z(n22556) );
  NANDN U11264 ( .A(y[7248]), .B(x[7248]), .Z(n8990) );
  NANDN U11265 ( .A(y[7249]), .B(x[7249]), .Z(n22555) );
  AND U11266 ( .A(n8990), .B(n22555), .Z(n60110) );
  XNOR U11267 ( .A(x[7248]), .B(y[7248]), .Z(n48169) );
  NANDN U11268 ( .A(y[7246]), .B(x[7246]), .Z(n8991) );
  NANDN U11269 ( .A(y[7247]), .B(x[7247]), .Z(n48168) );
  AND U11270 ( .A(n8991), .B(n48168), .Z(n60109) );
  NANDN U11271 ( .A(y[7244]), .B(x[7244]), .Z(n8992) );
  NANDN U11272 ( .A(y[7245]), .B(x[7245]), .Z(n22557) );
  AND U11273 ( .A(n8992), .B(n22557), .Z(n60107) );
  XNOR U11274 ( .A(x[7244]), .B(y[7244]), .Z(n22561) );
  NANDN U11275 ( .A(y[7242]), .B(x[7242]), .Z(n8993) );
  NANDN U11276 ( .A(y[7243]), .B(x[7243]), .Z(n22560) );
  NAND U11277 ( .A(n8993), .B(n22560), .Z(n60104) );
  XNOR U11278 ( .A(x[7242]), .B(y[7242]), .Z(n22563) );
  ANDN U11279 ( .B(y[7241]), .A(x[7241]), .Z(n60102) );
  ANDN U11280 ( .B(n22563), .A(n60102), .Z(n20379) );
  XNOR U11281 ( .A(x[7240]), .B(y[7240]), .Z(n48150) );
  NANDN U11282 ( .A(y[7238]), .B(x[7238]), .Z(n8994) );
  NANDN U11283 ( .A(y[7239]), .B(x[7239]), .Z(n48149) );
  AND U11284 ( .A(n8994), .B(n48149), .Z(n60097) );
  XNOR U11285 ( .A(x[7238]), .B(y[7238]), .Z(n22565) );
  NANDN U11286 ( .A(x[7237]), .B(y[7237]), .Z(n50800) );
  NAND U11287 ( .A(n22565), .B(n50800), .Z(n20372) );
  NANDN U11288 ( .A(y[7236]), .B(x[7236]), .Z(n8995) );
  NANDN U11289 ( .A(y[7237]), .B(x[7237]), .Z(n22564) );
  AND U11290 ( .A(n8995), .B(n22564), .Z(n60096) );
  XNOR U11291 ( .A(x[7236]), .B(y[7236]), .Z(n22567) );
  NANDN U11292 ( .A(x[7235]), .B(y[7235]), .Z(n60094) );
  NAND U11293 ( .A(n22567), .B(n60094), .Z(n20369) );
  NANDN U11294 ( .A(y[7234]), .B(x[7234]), .Z(n8996) );
  NANDN U11295 ( .A(y[7235]), .B(x[7235]), .Z(n22566) );
  AND U11296 ( .A(n8996), .B(n22566), .Z(n60093) );
  NANDN U11297 ( .A(x[7233]), .B(y[7233]), .Z(n22570) );
  IV U11298 ( .A(n22570), .Z(n50802) );
  XNOR U11299 ( .A(x[7234]), .B(y[7234]), .Z(n22569) );
  XNOR U11300 ( .A(y[7232]), .B(x[7232]), .Z(n48132) );
  NANDN U11301 ( .A(x[7231]), .B(y[7231]), .Z(n60090) );
  AND U11302 ( .A(n48132), .B(n60090), .Z(n20362) );
  NANDN U11303 ( .A(y[7230]), .B(x[7230]), .Z(n8997) );
  ANDN U11304 ( .B(x[7231]), .A(y[7231]), .Z(n48134) );
  ANDN U11305 ( .B(n8997), .A(n48134), .Z(n60089) );
  XNOR U11306 ( .A(x[7228]), .B(y[7228]), .Z(n48122) );
  NANDN U11307 ( .A(x[7227]), .B(y[7227]), .Z(n60085) );
  NAND U11308 ( .A(n48122), .B(n60085), .Z(n20355) );
  NANDN U11309 ( .A(y[7226]), .B(x[7226]), .Z(n8998) );
  NANDN U11310 ( .A(y[7227]), .B(x[7227]), .Z(n48121) );
  AND U11311 ( .A(n8998), .B(n48121), .Z(n60084) );
  ANDN U11312 ( .B(y[7225]), .A(x[7225]), .Z(n60082) );
  XNOR U11313 ( .A(x[7226]), .B(y[7226]), .Z(n22574) );
  NANDN U11314 ( .A(n60082), .B(n22574), .Z(n20352) );
  XNOR U11315 ( .A(x[7224]), .B(y[7224]), .Z(n48112) );
  NANDN U11316 ( .A(y[7222]), .B(x[7222]), .Z(n8999) );
  NANDN U11317 ( .A(y[7223]), .B(x[7223]), .Z(n48111) );
  NAND U11318 ( .A(n8999), .B(n48111), .Z(n60081) );
  NANDN U11319 ( .A(y[7220]), .B(x[7220]), .Z(n9000) );
  NANDN U11320 ( .A(y[7221]), .B(x[7221]), .Z(n22575) );
  AND U11321 ( .A(n9000), .B(n22575), .Z(n60078) );
  NANDN U11322 ( .A(x[7219]), .B(y[7219]), .Z(n48098) );
  IV U11323 ( .A(n48098), .Z(n50810) );
  XNOR U11324 ( .A(x[7220]), .B(y[7220]), .Z(n48102) );
  NANDN U11325 ( .A(y[7218]), .B(x[7218]), .Z(n9001) );
  NANDN U11326 ( .A(y[7219]), .B(x[7219]), .Z(n48101) );
  NAND U11327 ( .A(n9001), .B(n48101), .Z(n60077) );
  XNOR U11328 ( .A(x[7218]), .B(y[7218]), .Z(n22578) );
  ANDN U11329 ( .B(y[7217]), .A(x[7217]), .Z(n60074) );
  NANDN U11330 ( .A(y[7216]), .B(x[7216]), .Z(n9002) );
  NANDN U11331 ( .A(y[7217]), .B(x[7217]), .Z(n22577) );
  AND U11332 ( .A(n9002), .B(n22577), .Z(n60073) );
  XNOR U11333 ( .A(x[7216]), .B(y[7216]), .Z(n48091) );
  NANDN U11334 ( .A(y[7214]), .B(x[7214]), .Z(n9003) );
  NANDN U11335 ( .A(y[7215]), .B(x[7215]), .Z(n48090) );
  AND U11336 ( .A(n9003), .B(n48090), .Z(n50811) );
  XNOR U11337 ( .A(x[7214]), .B(y[7214]), .Z(n22580) );
  ANDN U11338 ( .B(y[7213]), .A(x[7213]), .Z(n60069) );
  ANDN U11339 ( .B(n22580), .A(n60069), .Z(n20333) );
  XNOR U11340 ( .A(x[7212]), .B(y[7212]), .Z(n48081) );
  NANDN U11341 ( .A(y[7210]), .B(x[7210]), .Z(n9004) );
  NANDN U11342 ( .A(y[7211]), .B(x[7211]), .Z(n48080) );
  AND U11343 ( .A(n9004), .B(n48080), .Z(n60065) );
  NANDN U11344 ( .A(x[7209]), .B(y[7209]), .Z(n60064) );
  NANDN U11345 ( .A(y[7208]), .B(x[7208]), .Z(n22583) );
  NANDN U11346 ( .A(y[7209]), .B(x[7209]), .Z(n22581) );
  AND U11347 ( .A(n22583), .B(n22581), .Z(n60062) );
  NANDN U11348 ( .A(y[7206]), .B(x[7206]), .Z(n22587) );
  NANDN U11349 ( .A(y[7207]), .B(x[7207]), .Z(n22584) );
  AND U11350 ( .A(n22587), .B(n22584), .Z(n60060) );
  NANDN U11351 ( .A(x[7206]), .B(y[7206]), .Z(n22586) );
  ANDN U11352 ( .B(y[7205]), .A(x[7205]), .Z(n48065) );
  ANDN U11353 ( .B(n22586), .A(n48065), .Z(n60059) );
  NANDN U11354 ( .A(y[7204]), .B(x[7204]), .Z(n9005) );
  NANDN U11355 ( .A(y[7205]), .B(x[7205]), .Z(n22588) );
  AND U11356 ( .A(n9005), .B(n22588), .Z(n60057) );
  XNOR U11357 ( .A(x[7204]), .B(y[7204]), .Z(n22590) );
  NANDN U11358 ( .A(y[7202]), .B(x[7202]), .Z(n22593) );
  NANDN U11359 ( .A(y[7203]), .B(x[7203]), .Z(n22589) );
  AND U11360 ( .A(n22593), .B(n22589), .Z(n60055) );
  XNOR U11361 ( .A(x[7200]), .B(y[7200]), .Z(n48053) );
  NANDN U11362 ( .A(y[7198]), .B(x[7198]), .Z(n9006) );
  NANDN U11363 ( .A(y[7199]), .B(x[7199]), .Z(n48052) );
  NAND U11364 ( .A(n9006), .B(n48052), .Z(n60053) );
  XNOR U11365 ( .A(x[7198]), .B(y[7198]), .Z(n22597) );
  NANDN U11366 ( .A(y[7196]), .B(x[7196]), .Z(n9007) );
  NANDN U11367 ( .A(y[7197]), .B(x[7197]), .Z(n22596) );
  AND U11368 ( .A(n9007), .B(n22596), .Z(n60050) );
  NANDN U11369 ( .A(y[7194]), .B(x[7194]), .Z(n9008) );
  NANDN U11370 ( .A(y[7195]), .B(x[7195]), .Z(n48042) );
  AND U11371 ( .A(n9008), .B(n48042), .Z(n60049) );
  XNOR U11372 ( .A(x[7194]), .B(y[7194]), .Z(n22599) );
  ANDN U11373 ( .B(y[7193]), .A(x[7193]), .Z(n60046) );
  ANDN U11374 ( .B(n22599), .A(n60046), .Z(n20304) );
  NANDN U11375 ( .A(x[7191]), .B(y[7191]), .Z(n22602) );
  NANDN U11376 ( .A(x[7192]), .B(y[7192]), .Z(n48036) );
  AND U11377 ( .A(n22602), .B(n48036), .Z(n60044) );
  NANDN U11378 ( .A(y[7190]), .B(x[7190]), .Z(n22604) );
  NANDN U11379 ( .A(y[7191]), .B(x[7191]), .Z(n22601) );
  AND U11380 ( .A(n22604), .B(n22601), .Z(n60043) );
  NANDN U11381 ( .A(x[7190]), .B(y[7190]), .Z(n22603) );
  ANDN U11382 ( .B(y[7189]), .A(x[7189]), .Z(n22606) );
  ANDN U11383 ( .B(n22603), .A(n22606), .Z(n60042) );
  NANDN U11384 ( .A(y[7188]), .B(x[7188]), .Z(n9009) );
  NANDN U11385 ( .A(y[7189]), .B(x[7189]), .Z(n22605) );
  NAND U11386 ( .A(n9009), .B(n22605), .Z(n60041) );
  XNOR U11387 ( .A(x[7188]), .B(y[7188]), .Z(n48024) );
  NANDN U11388 ( .A(x[7187]), .B(y[7187]), .Z(n60039) );
  AND U11389 ( .A(n48024), .B(n60039), .Z(n20297) );
  XNOR U11390 ( .A(x[7186]), .B(y[7186]), .Z(n22608) );
  NANDN U11391 ( .A(y[7184]), .B(x[7184]), .Z(n9010) );
  NANDN U11392 ( .A(y[7185]), .B(x[7185]), .Z(n22607) );
  AND U11393 ( .A(n9010), .B(n22607), .Z(n60037) );
  XNOR U11394 ( .A(x[7184]), .B(y[7184]), .Z(n48014) );
  NANDN U11395 ( .A(x[7183]), .B(y[7183]), .Z(n60035) );
  NAND U11396 ( .A(n48014), .B(n60035), .Z(n20290) );
  NANDN U11397 ( .A(y[7182]), .B(x[7182]), .Z(n9011) );
  NANDN U11398 ( .A(y[7183]), .B(x[7183]), .Z(n48013) );
  AND U11399 ( .A(n9011), .B(n48013), .Z(n60034) );
  XNOR U11400 ( .A(x[7182]), .B(y[7182]), .Z(n22611) );
  NANDN U11401 ( .A(x[7181]), .B(y[7181]), .Z(n60032) );
  NAND U11402 ( .A(n22611), .B(n60032), .Z(n20287) );
  XNOR U11403 ( .A(x[7180]), .B(y[7180]), .Z(n22613) );
  NANDN U11404 ( .A(y[7178]), .B(x[7178]), .Z(n9012) );
  NANDN U11405 ( .A(y[7179]), .B(x[7179]), .Z(n22612) );
  AND U11406 ( .A(n9012), .B(n22612), .Z(n60027) );
  ANDN U11407 ( .B(x[7175]), .A(y[7175]), .Z(n47998) );
  NANDN U11408 ( .A(y[7174]), .B(x[7174]), .Z(n9013) );
  NANDN U11409 ( .A(n47998), .B(n9013), .Z(n60024) );
  XNOR U11410 ( .A(x[7174]), .B(y[7174]), .Z(n22617) );
  ANDN U11411 ( .B(y[7173]), .A(x[7173]), .Z(n60022) );
  NANDN U11412 ( .A(y[7172]), .B(x[7172]), .Z(n9014) );
  NANDN U11413 ( .A(y[7173]), .B(x[7173]), .Z(n22616) );
  AND U11414 ( .A(n9014), .B(n22616), .Z(n60021) );
  NANDN U11415 ( .A(x[7171]), .B(y[7171]), .Z(n47982) );
  IV U11416 ( .A(n47982), .Z(n50825) );
  XNOR U11417 ( .A(x[7172]), .B(y[7172]), .Z(n47986) );
  NANDN U11418 ( .A(y[7170]), .B(x[7170]), .Z(n9015) );
  NANDN U11419 ( .A(y[7171]), .B(x[7171]), .Z(n47985) );
  AND U11420 ( .A(n9015), .B(n47985), .Z(n60020) );
  XNOR U11421 ( .A(x[7170]), .B(y[7170]), .Z(n22619) );
  ANDN U11422 ( .B(y[7169]), .A(x[7169]), .Z(n60018) );
  ANDN U11423 ( .B(n22619), .A(n60018), .Z(n20267) );
  XNOR U11424 ( .A(x[7168]), .B(y[7168]), .Z(n47975) );
  NANDN U11425 ( .A(y[7166]), .B(x[7166]), .Z(n9016) );
  NANDN U11426 ( .A(y[7167]), .B(x[7167]), .Z(n47974) );
  AND U11427 ( .A(n9016), .B(n47974), .Z(n60013) );
  XNOR U11428 ( .A(x[7166]), .B(y[7166]), .Z(n22621) );
  ANDN U11429 ( .B(y[7165]), .A(x[7165]), .Z(n60011) );
  ANDN U11430 ( .B(n22621), .A(n60011), .Z(n20260) );
  XNOR U11431 ( .A(x[7164]), .B(y[7164]), .Z(n47965) );
  XNOR U11432 ( .A(x[7162]), .B(y[7162]), .Z(n22623) );
  NANDN U11433 ( .A(y[7160]), .B(x[7160]), .Z(n9017) );
  NANDN U11434 ( .A(y[7161]), .B(x[7161]), .Z(n22622) );
  AND U11435 ( .A(n9017), .B(n22622), .Z(n60005) );
  NANDN U11436 ( .A(y[7158]), .B(x[7158]), .Z(n9018) );
  NANDN U11437 ( .A(y[7159]), .B(x[7159]), .Z(n47954) );
  AND U11438 ( .A(n9018), .B(n47954), .Z(n60003) );
  XNOR U11439 ( .A(x[7158]), .B(y[7158]), .Z(n22626) );
  NANDN U11440 ( .A(y[7156]), .B(x[7156]), .Z(n9019) );
  NANDN U11441 ( .A(y[7157]), .B(x[7157]), .Z(n22625) );
  NAND U11442 ( .A(n9019), .B(n22625), .Z(n50829) );
  XNOR U11443 ( .A(x[7156]), .B(y[7156]), .Z(n22628) );
  NANDN U11444 ( .A(x[7155]), .B(y[7155]), .Z(n50830) );
  AND U11445 ( .A(n22628), .B(n50830), .Z(n20244) );
  XNOR U11446 ( .A(x[7154]), .B(y[7154]), .Z(n22630) );
  NANDN U11447 ( .A(y[7152]), .B(x[7152]), .Z(n9020) );
  NANDN U11448 ( .A(y[7153]), .B(x[7153]), .Z(n22629) );
  AND U11449 ( .A(n9020), .B(n22629), .Z(n59998) );
  XNOR U11450 ( .A(x[7152]), .B(y[7152]), .Z(n47936) );
  NANDN U11451 ( .A(x[7151]), .B(y[7151]), .Z(n50833) );
  NAND U11452 ( .A(n47936), .B(n50833), .Z(n20237) );
  NANDN U11453 ( .A(y[7150]), .B(x[7150]), .Z(n9021) );
  NANDN U11454 ( .A(y[7151]), .B(x[7151]), .Z(n47935) );
  AND U11455 ( .A(n9021), .B(n47935), .Z(n59997) );
  ANDN U11456 ( .B(y[7149]), .A(x[7149]), .Z(n59995) );
  XNOR U11457 ( .A(x[7150]), .B(y[7150]), .Z(n22632) );
  NANDN U11458 ( .A(n59995), .B(n22632), .Z(n20234) );
  NANDN U11459 ( .A(y[7148]), .B(x[7148]), .Z(n9022) );
  NANDN U11460 ( .A(y[7149]), .B(x[7149]), .Z(n22631) );
  AND U11461 ( .A(n9022), .B(n22631), .Z(n59994) );
  XNOR U11462 ( .A(x[7148]), .B(y[7148]), .Z(n47926) );
  XNOR U11463 ( .A(x[7146]), .B(y[7146]), .Z(n22634) );
  NANDN U11464 ( .A(y[7144]), .B(x[7144]), .Z(n9023) );
  NANDN U11465 ( .A(y[7145]), .B(x[7145]), .Z(n22633) );
  AND U11466 ( .A(n9023), .B(n22633), .Z(n59992) );
  XNOR U11467 ( .A(y[7144]), .B(x[7144]), .Z(n22637) );
  NANDN U11468 ( .A(x[7143]), .B(y[7143]), .Z(n22638) );
  AND U11469 ( .A(n22637), .B(n22638), .Z(n59991) );
  NANDN U11470 ( .A(y[7142]), .B(x[7142]), .Z(n9024) );
  NANDN U11471 ( .A(y[7143]), .B(x[7143]), .Z(n22636) );
  NAND U11472 ( .A(n9024), .B(n22636), .Z(n59990) );
  NANDN U11473 ( .A(y[7140]), .B(x[7140]), .Z(n9025) );
  NANDN U11474 ( .A(y[7141]), .B(x[7141]), .Z(n22639) );
  AND U11475 ( .A(n9025), .B(n22639), .Z(n59989) );
  XNOR U11476 ( .A(x[7140]), .B(y[7140]), .Z(n47908) );
  NANDN U11477 ( .A(y[7138]), .B(x[7138]), .Z(n9026) );
  NANDN U11478 ( .A(y[7139]), .B(x[7139]), .Z(n47907) );
  AND U11479 ( .A(n9026), .B(n47907), .Z(n59986) );
  XNOR U11480 ( .A(x[7138]), .B(y[7138]), .Z(n22642) );
  NANDN U11481 ( .A(x[7137]), .B(y[7137]), .Z(n22643) );
  XNOR U11482 ( .A(x[7136]), .B(y[7136]), .Z(n47898) );
  NANDN U11483 ( .A(y[7134]), .B(x[7134]), .Z(n9027) );
  NANDN U11484 ( .A(y[7135]), .B(x[7135]), .Z(n47897) );
  AND U11485 ( .A(n9027), .B(n47897), .Z(n59981) );
  XNOR U11486 ( .A(x[7134]), .B(y[7134]), .Z(n22645) );
  ANDN U11487 ( .B(y[7133]), .A(x[7133]), .Z(n59978) );
  ANDN U11488 ( .B(n22645), .A(n59978), .Z(n20226) );
  XNOR U11489 ( .A(x[7132]), .B(y[7132]), .Z(n47888) );
  NANDN U11490 ( .A(y[7130]), .B(x[7130]), .Z(n9028) );
  NANDN U11491 ( .A(y[7131]), .B(x[7131]), .Z(n47887) );
  AND U11492 ( .A(n9028), .B(n47887), .Z(n59975) );
  XNOR U11493 ( .A(x[7130]), .B(y[7130]), .Z(n22647) );
  NANDN U11494 ( .A(y[7128]), .B(x[7128]), .Z(n9029) );
  NANDN U11495 ( .A(y[7129]), .B(x[7129]), .Z(n22646) );
  AND U11496 ( .A(n9029), .B(n22646), .Z(n50843) );
  ANDN U11497 ( .B(y[7127]), .A(x[7127]), .Z(n47874) );
  XNOR U11498 ( .A(x[7128]), .B(y[7128]), .Z(n47878) );
  NANDN U11499 ( .A(y[7126]), .B(x[7126]), .Z(n9030) );
  NANDN U11500 ( .A(y[7127]), .B(x[7127]), .Z(n47877) );
  AND U11501 ( .A(n9030), .B(n47877), .Z(n59970) );
  ANDN U11502 ( .B(y[7125]), .A(x[7125]), .Z(n59968) );
  XNOR U11503 ( .A(x[7126]), .B(y[7126]), .Z(n22649) );
  NANDN U11504 ( .A(y[7124]), .B(x[7124]), .Z(n9031) );
  NANDN U11505 ( .A(y[7125]), .B(x[7125]), .Z(n22648) );
  AND U11506 ( .A(n9031), .B(n22648), .Z(n59967) );
  NANDN U11507 ( .A(y[7122]), .B(x[7122]), .Z(n9032) );
  NANDN U11508 ( .A(y[7123]), .B(x[7123]), .Z(n22650) );
  AND U11509 ( .A(n9032), .B(n22650), .Z(n59965) );
  ANDN U11510 ( .B(y[7121]), .A(x[7121]), .Z(n59963) );
  XNOR U11511 ( .A(x[7122]), .B(y[7122]), .Z(n22653) );
  NANDN U11512 ( .A(y[7120]), .B(x[7120]), .Z(n9033) );
  NANDN U11513 ( .A(y[7121]), .B(x[7121]), .Z(n22652) );
  AND U11514 ( .A(n9033), .B(n22652), .Z(n59962) );
  XNOR U11515 ( .A(x[7120]), .B(y[7120]), .Z(n47859) );
  NANDN U11516 ( .A(x[7119]), .B(y[7119]), .Z(n59960) );
  AND U11517 ( .A(n47859), .B(n59960), .Z(n20204) );
  NANDN U11518 ( .A(y[7118]), .B(x[7118]), .Z(n9034) );
  NANDN U11519 ( .A(y[7119]), .B(x[7119]), .Z(n47858) );
  NAND U11520 ( .A(n9034), .B(n47858), .Z(n59959) );
  XNOR U11521 ( .A(x[7118]), .B(y[7118]), .Z(n22655) );
  NANDN U11522 ( .A(y[7116]), .B(x[7116]), .Z(n9035) );
  NANDN U11523 ( .A(y[7117]), .B(x[7117]), .Z(n22654) );
  AND U11524 ( .A(n9035), .B(n22654), .Z(n59956) );
  XNOR U11525 ( .A(x[7116]), .B(y[7116]), .Z(n47849) );
  NANDN U11526 ( .A(x[7115]), .B(y[7115]), .Z(n59954) );
  NAND U11527 ( .A(n47849), .B(n59954), .Z(n20198) );
  NANDN U11528 ( .A(y[7114]), .B(x[7114]), .Z(n9036) );
  NANDN U11529 ( .A(y[7115]), .B(x[7115]), .Z(n47848) );
  AND U11530 ( .A(n9036), .B(n47848), .Z(n50847) );
  NANDN U11531 ( .A(x[7113]), .B(y[7113]), .Z(n59953) );
  XNOR U11532 ( .A(x[7114]), .B(y[7114]), .Z(n22657) );
  NAND U11533 ( .A(n59953), .B(n22657), .Z(n20195) );
  NANDN U11534 ( .A(y[7112]), .B(x[7112]), .Z(n9037) );
  NANDN U11535 ( .A(y[7113]), .B(x[7113]), .Z(n22656) );
  AND U11536 ( .A(n9037), .B(n22656), .Z(n59951) );
  XNOR U11537 ( .A(x[7112]), .B(y[7112]), .Z(n47839) );
  NANDN U11538 ( .A(y[7110]), .B(x[7110]), .Z(n9038) );
  NANDN U11539 ( .A(y[7111]), .B(x[7111]), .Z(n47838) );
  NAND U11540 ( .A(n9038), .B(n47838), .Z(n50848) );
  NANDN U11541 ( .A(y[7108]), .B(x[7108]), .Z(n9039) );
  NANDN U11542 ( .A(y[7109]), .B(x[7109]), .Z(n22658) );
  AND U11543 ( .A(n9039), .B(n22658), .Z(n59946) );
  XNOR U11544 ( .A(x[7108]), .B(y[7108]), .Z(n47829) );
  NANDN U11545 ( .A(y[7106]), .B(x[7106]), .Z(n9040) );
  NANDN U11546 ( .A(y[7107]), .B(x[7107]), .Z(n47828) );
  AND U11547 ( .A(n9040), .B(n47828), .Z(n59943) );
  XNOR U11548 ( .A(x[7106]), .B(y[7106]), .Z(n22662) );
  ANDN U11549 ( .B(y[7105]), .A(x[7105]), .Z(n59941) );
  ANDN U11550 ( .B(n22662), .A(n59941), .Z(n20183) );
  NANDN U11551 ( .A(y[7104]), .B(x[7104]), .Z(n9041) );
  NANDN U11552 ( .A(y[7105]), .B(x[7105]), .Z(n22661) );
  NAND U11553 ( .A(n9041), .B(n22661), .Z(n59940) );
  XNOR U11554 ( .A(x[7104]), .B(y[7104]), .Z(n47819) );
  NANDN U11555 ( .A(y[7102]), .B(x[7102]), .Z(n9042) );
  NANDN U11556 ( .A(y[7103]), .B(x[7103]), .Z(n47818) );
  AND U11557 ( .A(n9042), .B(n47818), .Z(n59938) );
  ANDN U11558 ( .B(y[7101]), .A(x[7101]), .Z(n59936) );
  XNOR U11559 ( .A(x[7102]), .B(y[7102]), .Z(n22664) );
  NANDN U11560 ( .A(n59936), .B(n22664), .Z(n20177) );
  NANDN U11561 ( .A(y[7100]), .B(x[7100]), .Z(n9043) );
  NANDN U11562 ( .A(y[7101]), .B(x[7101]), .Z(n22663) );
  AND U11563 ( .A(n9043), .B(n22663), .Z(n50852) );
  XNOR U11564 ( .A(x[7100]), .B(y[7100]), .Z(n47809) );
  NANDN U11565 ( .A(x[7099]), .B(y[7099]), .Z(n50855) );
  NAND U11566 ( .A(n47809), .B(n50855), .Z(n20174) );
  ANDN U11567 ( .B(y[7097]), .A(x[7097]), .Z(n59931) );
  XNOR U11568 ( .A(x[7098]), .B(y[7098]), .Z(n22666) );
  XNOR U11569 ( .A(x[7096]), .B(y[7096]), .Z(n47799) );
  NANDN U11570 ( .A(y[7094]), .B(x[7094]), .Z(n22668) );
  NANDN U11571 ( .A(y[7095]), .B(x[7095]), .Z(n47798) );
  AND U11572 ( .A(n22668), .B(n47798), .Z(n59929) );
  NANDN U11573 ( .A(x[7093]), .B(y[7093]), .Z(n22670) );
  NANDN U11574 ( .A(x[7094]), .B(y[7094]), .Z(n22667) );
  AND U11575 ( .A(n22670), .B(n22667), .Z(n59928) );
  NANDN U11576 ( .A(y[7092]), .B(x[7092]), .Z(n9044) );
  NANDN U11577 ( .A(y[7093]), .B(x[7093]), .Z(n22669) );
  AND U11578 ( .A(n9044), .B(n22669), .Z(n59927) );
  XNOR U11579 ( .A(x[7092]), .B(y[7092]), .Z(n22672) );
  NANDN U11580 ( .A(x[7091]), .B(y[7091]), .Z(n59925) );
  AND U11581 ( .A(n22672), .B(n59925), .Z(n20161) );
  XNOR U11582 ( .A(x[7090]), .B(y[7090]), .Z(n22674) );
  NANDN U11583 ( .A(y[7088]), .B(x[7088]), .Z(n9045) );
  NANDN U11584 ( .A(y[7089]), .B(x[7089]), .Z(n22673) );
  AND U11585 ( .A(n9045), .B(n22673), .Z(n59922) );
  XNOR U11586 ( .A(x[7088]), .B(y[7088]), .Z(n47781) );
  NANDN U11587 ( .A(x[7087]), .B(y[7087]), .Z(n59920) );
  NAND U11588 ( .A(n47781), .B(n59920), .Z(n20154) );
  NANDN U11589 ( .A(y[7086]), .B(x[7086]), .Z(n9046) );
  NANDN U11590 ( .A(y[7087]), .B(x[7087]), .Z(n47780) );
  AND U11591 ( .A(n9046), .B(n47780), .Z(n50859) );
  NANDN U11592 ( .A(x[7085]), .B(y[7085]), .Z(n59918) );
  XNOR U11593 ( .A(x[7086]), .B(y[7086]), .Z(n22676) );
  NAND U11594 ( .A(n59918), .B(n22676), .Z(n20151) );
  NANDN U11595 ( .A(y[7084]), .B(x[7084]), .Z(n9047) );
  NANDN U11596 ( .A(y[7085]), .B(x[7085]), .Z(n22675) );
  AND U11597 ( .A(n9047), .B(n22675), .Z(n59916) );
  XNOR U11598 ( .A(x[7084]), .B(y[7084]), .Z(n47771) );
  NANDN U11599 ( .A(y[7082]), .B(x[7082]), .Z(n9048) );
  NANDN U11600 ( .A(y[7083]), .B(x[7083]), .Z(n47770) );
  NAND U11601 ( .A(n9048), .B(n47770), .Z(n59915) );
  XNOR U11602 ( .A(x[7080]), .B(y[7080]), .Z(n22680) );
  NANDN U11603 ( .A(y[7078]), .B(x[7078]), .Z(n9049) );
  NANDN U11604 ( .A(y[7079]), .B(x[7079]), .Z(n22679) );
  AND U11605 ( .A(n9049), .B(n22679), .Z(n59910) );
  XNOR U11606 ( .A(x[7078]), .B(y[7078]), .Z(n22682) );
  ANDN U11607 ( .B(y[7077]), .A(x[7077]), .Z(n59908) );
  ANDN U11608 ( .B(n22682), .A(n59908), .Z(n20138) );
  NANDN U11609 ( .A(y[7076]), .B(x[7076]), .Z(n9050) );
  NANDN U11610 ( .A(y[7077]), .B(x[7077]), .Z(n22681) );
  NAND U11611 ( .A(n9050), .B(n22681), .Z(n59907) );
  XNOR U11612 ( .A(x[7076]), .B(y[7076]), .Z(n47753) );
  NANDN U11613 ( .A(y[7074]), .B(x[7074]), .Z(n9051) );
  NANDN U11614 ( .A(y[7075]), .B(x[7075]), .Z(n47752) );
  AND U11615 ( .A(n9051), .B(n47752), .Z(n59905) );
  ANDN U11616 ( .B(y[7073]), .A(x[7073]), .Z(n59903) );
  XNOR U11617 ( .A(x[7074]), .B(y[7074]), .Z(n22684) );
  NANDN U11618 ( .A(n59903), .B(n22684), .Z(n20132) );
  NANDN U11619 ( .A(y[7072]), .B(x[7072]), .Z(n9052) );
  NANDN U11620 ( .A(y[7073]), .B(x[7073]), .Z(n22683) );
  AND U11621 ( .A(n9052), .B(n22683), .Z(n59902) );
  NANDN U11622 ( .A(x[7071]), .B(y[7071]), .Z(n50865) );
  XNOR U11623 ( .A(x[7072]), .B(y[7072]), .Z(n47743) );
  NAND U11624 ( .A(n50865), .B(n47743), .Z(n20129) );
  NANDN U11625 ( .A(y[7070]), .B(x[7070]), .Z(n9053) );
  NANDN U11626 ( .A(y[7071]), .B(x[7071]), .Z(n47742) );
  AND U11627 ( .A(n9053), .B(n47742), .Z(n59901) );
  ANDN U11628 ( .B(y[7069]), .A(x[7069]), .Z(n59899) );
  XNOR U11629 ( .A(x[7070]), .B(y[7070]), .Z(n22686) );
  NANDN U11630 ( .A(y[7068]), .B(x[7068]), .Z(n9054) );
  NANDN U11631 ( .A(y[7069]), .B(x[7069]), .Z(n22685) );
  AND U11632 ( .A(n9054), .B(n22685), .Z(n59898) );
  XNOR U11633 ( .A(x[7068]), .B(y[7068]), .Z(n47733) );
  NANDN U11634 ( .A(y[7066]), .B(x[7066]), .Z(n9055) );
  NANDN U11635 ( .A(y[7067]), .B(x[7067]), .Z(n47732) );
  AND U11636 ( .A(n9055), .B(n47732), .Z(n59895) );
  ANDN U11637 ( .B(y[7065]), .A(x[7065]), .Z(n59893) );
  XNOR U11638 ( .A(x[7066]), .B(y[7066]), .Z(n22688) );
  NANDN U11639 ( .A(y[7064]), .B(x[7064]), .Z(n9056) );
  NANDN U11640 ( .A(y[7065]), .B(x[7065]), .Z(n22687) );
  AND U11641 ( .A(n9056), .B(n22687), .Z(n59892) );
  XNOR U11642 ( .A(x[7064]), .B(y[7064]), .Z(n47723) );
  NANDN U11643 ( .A(x[7063]), .B(y[7063]), .Z(n59889) );
  AND U11644 ( .A(n47723), .B(n59889), .Z(n20117) );
  NANDN U11645 ( .A(y[7062]), .B(x[7062]), .Z(n9057) );
  NANDN U11646 ( .A(y[7063]), .B(x[7063]), .Z(n47722) );
  NAND U11647 ( .A(n9057), .B(n47722), .Z(n59888) );
  XNOR U11648 ( .A(x[7062]), .B(y[7062]), .Z(n22690) );
  NANDN U11649 ( .A(x[7059]), .B(y[7059]), .Z(n59885) );
  XNOR U11650 ( .A(x[7060]), .B(y[7060]), .Z(n22692) );
  AND U11651 ( .A(n59885), .B(n22692), .Z(n20110) );
  XNOR U11652 ( .A(y[7058]), .B(x[7058]), .Z(n22695) );
  ANDN U11653 ( .B(y[7057]), .A(x[7057]), .Z(n47708) );
  ANDN U11654 ( .B(n22695), .A(n47708), .Z(n59883) );
  NANDN U11655 ( .A(y[7056]), .B(x[7056]), .Z(n9058) );
  NANDN U11656 ( .A(y[7057]), .B(x[7057]), .Z(n22694) );
  AND U11657 ( .A(n9058), .B(n22694), .Z(n59882) );
  XNOR U11658 ( .A(x[7056]), .B(y[7056]), .Z(n22697) );
  NANDN U11659 ( .A(y[7054]), .B(x[7054]), .Z(n9059) );
  NANDN U11660 ( .A(y[7055]), .B(x[7055]), .Z(n22696) );
  AND U11661 ( .A(n9059), .B(n22696), .Z(n59879) );
  XNOR U11662 ( .A(x[7052]), .B(y[7052]), .Z(n47696) );
  NANDN U11663 ( .A(y[7050]), .B(x[7050]), .Z(n9060) );
  NANDN U11664 ( .A(y[7051]), .B(x[7051]), .Z(n47695) );
  AND U11665 ( .A(n9060), .B(n47695), .Z(n59874) );
  XNOR U11666 ( .A(x[7050]), .B(y[7050]), .Z(n22701) );
  ANDN U11667 ( .B(y[7049]), .A(x[7049]), .Z(n59872) );
  ANDN U11668 ( .B(n22701), .A(n59872), .Z(n20094) );
  XNOR U11669 ( .A(x[7048]), .B(y[7048]), .Z(n22703) );
  NANDN U11670 ( .A(y[7046]), .B(x[7046]), .Z(n9061) );
  NANDN U11671 ( .A(y[7047]), .B(x[7047]), .Z(n22702) );
  AND U11672 ( .A(n9061), .B(n22702), .Z(n59869) );
  XNOR U11673 ( .A(x[7046]), .B(y[7046]), .Z(n22705) );
  ANDN U11674 ( .B(y[7045]), .A(x[7045]), .Z(n59867) );
  ANDN U11675 ( .B(n22705), .A(n59867), .Z(n20087) );
  XNOR U11676 ( .A(x[7044]), .B(y[7044]), .Z(n47678) );
  NANDN U11677 ( .A(y[7042]), .B(x[7042]), .Z(n9062) );
  NANDN U11678 ( .A(y[7043]), .B(x[7043]), .Z(n47677) );
  AND U11679 ( .A(n9062), .B(n47677), .Z(n59864) );
  ANDN U11680 ( .B(y[7041]), .A(x[7041]), .Z(n22708) );
  XNOR U11681 ( .A(y[7042]), .B(x[7042]), .Z(n22707) );
  NANDN U11682 ( .A(n22708), .B(n22707), .Z(n59863) );
  NANDN U11683 ( .A(y[7040]), .B(x[7040]), .Z(n9063) );
  NANDN U11684 ( .A(y[7041]), .B(x[7041]), .Z(n22706) );
  AND U11685 ( .A(n9063), .B(n22706), .Z(n59862) );
  XNOR U11686 ( .A(x[7040]), .B(y[7040]), .Z(n47667) );
  NANDN U11687 ( .A(y[7038]), .B(x[7038]), .Z(n9064) );
  NANDN U11688 ( .A(y[7039]), .B(x[7039]), .Z(n47666) );
  AND U11689 ( .A(n9064), .B(n47666), .Z(n59859) );
  ANDN U11690 ( .B(y[7037]), .A(x[7037]), .Z(n59857) );
  XNOR U11691 ( .A(x[7038]), .B(y[7038]), .Z(n22710) );
  NANDN U11692 ( .A(y[7036]), .B(x[7036]), .Z(n9065) );
  NANDN U11693 ( .A(y[7037]), .B(x[7037]), .Z(n22709) );
  AND U11694 ( .A(n9065), .B(n22709), .Z(n59856) );
  ANDN U11695 ( .B(y[7033]), .A(x[7033]), .Z(n50875) );
  XNOR U11696 ( .A(x[7034]), .B(y[7034]), .Z(n22712) );
  NANDN U11697 ( .A(y[7032]), .B(x[7032]), .Z(n9066) );
  NANDN U11698 ( .A(y[7033]), .B(x[7033]), .Z(n22711) );
  NAND U11699 ( .A(n9066), .B(n22711), .Z(n59853) );
  XNOR U11700 ( .A(x[7032]), .B(y[7032]), .Z(n47646) );
  NANDN U11701 ( .A(x[7031]), .B(y[7031]), .Z(n59851) );
  AND U11702 ( .A(n47646), .B(n59851), .Z(n20065) );
  XNOR U11703 ( .A(x[7030]), .B(y[7030]), .Z(n22714) );
  NANDN U11704 ( .A(y[7028]), .B(x[7028]), .Z(n9067) );
  NANDN U11705 ( .A(y[7029]), .B(x[7029]), .Z(n22713) );
  AND U11706 ( .A(n9067), .B(n22713), .Z(n59848) );
  XNOR U11707 ( .A(x[7028]), .B(y[7028]), .Z(n47636) );
  NANDN U11708 ( .A(x[7027]), .B(y[7027]), .Z(n59846) );
  NAND U11709 ( .A(n47636), .B(n59846), .Z(n20058) );
  NANDN U11710 ( .A(y[7026]), .B(x[7026]), .Z(n9068) );
  NANDN U11711 ( .A(y[7027]), .B(x[7027]), .Z(n47635) );
  AND U11712 ( .A(n9068), .B(n47635), .Z(n59845) );
  ANDN U11713 ( .B(y[7025]), .A(x[7025]), .Z(n59843) );
  XNOR U11714 ( .A(x[7026]), .B(y[7026]), .Z(n22717) );
  NANDN U11715 ( .A(n59843), .B(n22717), .Z(n20055) );
  XNOR U11716 ( .A(x[7024]), .B(y[7024]), .Z(n47626) );
  NANDN U11717 ( .A(y[7022]), .B(x[7022]), .Z(n9069) );
  NANDN U11718 ( .A(y[7023]), .B(x[7023]), .Z(n47625) );
  AND U11719 ( .A(n9069), .B(n47625), .Z(n59841) );
  XNOR U11720 ( .A(x[7020]), .B(y[7020]), .Z(n47616) );
  NANDN U11721 ( .A(y[7018]), .B(x[7018]), .Z(n9070) );
  NANDN U11722 ( .A(y[7019]), .B(x[7019]), .Z(n47615) );
  NAND U11723 ( .A(n9070), .B(n47615), .Z(n59837) );
  ANDN U11724 ( .B(y[7017]), .A(x[7017]), .Z(n59835) );
  XNOR U11725 ( .A(x[7018]), .B(y[7018]), .Z(n22721) );
  NANDN U11726 ( .A(y[7016]), .B(x[7016]), .Z(n9071) );
  NANDN U11727 ( .A(y[7017]), .B(x[7017]), .Z(n22720) );
  AND U11728 ( .A(n9071), .B(n22720), .Z(n59834) );
  NANDN U11729 ( .A(x[7015]), .B(y[7015]), .Z(n50886) );
  XNOR U11730 ( .A(x[7016]), .B(y[7016]), .Z(n47606) );
  AND U11731 ( .A(n50886), .B(n47606), .Z(n20038) );
  XNOR U11732 ( .A(x[7014]), .B(y[7014]), .Z(n22723) );
  NANDN U11733 ( .A(y[7012]), .B(x[7012]), .Z(n9072) );
  NANDN U11734 ( .A(y[7013]), .B(x[7013]), .Z(n22722) );
  AND U11735 ( .A(n9072), .B(n22722), .Z(n59830) );
  ANDN U11736 ( .B(y[7009]), .A(x[7009]), .Z(n59825) );
  XNOR U11737 ( .A(x[7010]), .B(y[7010]), .Z(n22725) );
  NANDN U11738 ( .A(y[7008]), .B(x[7008]), .Z(n9073) );
  NANDN U11739 ( .A(y[7009]), .B(x[7009]), .Z(n22724) );
  NAND U11740 ( .A(n9073), .B(n22724), .Z(n59824) );
  XNOR U11741 ( .A(x[7008]), .B(y[7008]), .Z(n47586) );
  NANDN U11742 ( .A(x[7007]), .B(y[7007]), .Z(n59821) );
  AND U11743 ( .A(n47586), .B(n59821), .Z(n20024) );
  XNOR U11744 ( .A(x[7006]), .B(y[7006]), .Z(n22727) );
  NANDN U11745 ( .A(y[7004]), .B(x[7004]), .Z(n9074) );
  NANDN U11746 ( .A(y[7005]), .B(x[7005]), .Z(n22726) );
  AND U11747 ( .A(n9074), .B(n22726), .Z(n59817) );
  XNOR U11748 ( .A(x[7004]), .B(y[7004]), .Z(n22729) );
  NANDN U11749 ( .A(x[7003]), .B(y[7003]), .Z(n59815) );
  XNOR U11750 ( .A(x[7002]), .B(y[7002]), .Z(n22731) );
  NANDN U11751 ( .A(y[7000]), .B(x[7000]), .Z(n9075) );
  NANDN U11752 ( .A(y[7001]), .B(x[7001]), .Z(n22730) );
  AND U11753 ( .A(n9075), .B(n22730), .Z(n59811) );
  NANDN U11754 ( .A(x[6999]), .B(y[6999]), .Z(n59810) );
  XOR U11755 ( .A(x[7000]), .B(y[7000]), .Z(n47569) );
  NANDN U11756 ( .A(y[6996]), .B(x[6996]), .Z(n9076) );
  NANDN U11757 ( .A(y[6997]), .B(x[6997]), .Z(n22734) );
  AND U11758 ( .A(n9076), .B(n22734), .Z(n59807) );
  XNOR U11759 ( .A(x[6996]), .B(y[6996]), .Z(n22737) );
  NANDN U11760 ( .A(y[6994]), .B(x[6994]), .Z(n9077) );
  NANDN U11761 ( .A(y[6995]), .B(x[6995]), .Z(n22736) );
  NAND U11762 ( .A(n9077), .B(n22736), .Z(n59804) );
  ANDN U11763 ( .B(y[6993]), .A(x[6993]), .Z(n50891) );
  XNOR U11764 ( .A(x[6994]), .B(y[6994]), .Z(n22739) );
  NANDN U11765 ( .A(y[6992]), .B(x[6992]), .Z(n9078) );
  NANDN U11766 ( .A(y[6993]), .B(x[6993]), .Z(n22738) );
  NAND U11767 ( .A(n9078), .B(n22738), .Z(n59803) );
  NANDN U11768 ( .A(y[6990]), .B(x[6990]), .Z(n9079) );
  NANDN U11769 ( .A(y[6991]), .B(x[6991]), .Z(n47549) );
  AND U11770 ( .A(n9079), .B(n47549), .Z(n59800) );
  XNOR U11771 ( .A(x[6990]), .B(y[6990]), .Z(n22741) );
  ANDN U11772 ( .B(y[6989]), .A(x[6989]), .Z(n50893) );
  ANDN U11773 ( .B(n22741), .A(n50893), .Z(n20014) );
  XNOR U11774 ( .A(x[6988]), .B(y[6988]), .Z(n47540) );
  NANDN U11775 ( .A(y[6986]), .B(x[6986]), .Z(n9080) );
  NANDN U11776 ( .A(y[6987]), .B(x[6987]), .Z(n47539) );
  AND U11777 ( .A(n9080), .B(n47539), .Z(n59796) );
  ANDN U11778 ( .B(y[6985]), .A(x[6985]), .Z(n59794) );
  XNOR U11779 ( .A(x[6986]), .B(y[6986]), .Z(n22743) );
  NANDN U11780 ( .A(y[6984]), .B(x[6984]), .Z(n9081) );
  NANDN U11781 ( .A(y[6985]), .B(x[6985]), .Z(n22742) );
  NAND U11782 ( .A(n9081), .B(n22742), .Z(n59793) );
  NANDN U11783 ( .A(y[6982]), .B(x[6982]), .Z(n9082) );
  NANDN U11784 ( .A(y[6983]), .B(x[6983]), .Z(n47529) );
  AND U11785 ( .A(n9082), .B(n47529), .Z(n59789) );
  XNOR U11786 ( .A(x[6982]), .B(y[6982]), .Z(n22745) );
  ANDN U11787 ( .B(y[6981]), .A(x[6981]), .Z(n59787) );
  ANDN U11788 ( .B(n22745), .A(n59787), .Z(n20001) );
  NANDN U11789 ( .A(y[6980]), .B(x[6980]), .Z(n9083) );
  NANDN U11790 ( .A(y[6981]), .B(x[6981]), .Z(n22744) );
  NAND U11791 ( .A(n9083), .B(n22744), .Z(n59786) );
  XNOR U11792 ( .A(x[6980]), .B(y[6980]), .Z(n47520) );
  NANDN U11793 ( .A(x[6979]), .B(y[6979]), .Z(n50897) );
  AND U11794 ( .A(n47520), .B(n50897), .Z(n19998) );
  XNOR U11795 ( .A(x[6978]), .B(y[6978]), .Z(n22747) );
  NANDN U11796 ( .A(y[6976]), .B(x[6976]), .Z(n9084) );
  NANDN U11797 ( .A(y[6977]), .B(x[6977]), .Z(n22746) );
  AND U11798 ( .A(n9084), .B(n22746), .Z(n59782) );
  XNOR U11799 ( .A(x[6976]), .B(y[6976]), .Z(n22749) );
  NANDN U11800 ( .A(x[6975]), .B(y[6975]), .Z(n50898) );
  AND U11801 ( .A(n22749), .B(n50898), .Z(n19991) );
  XNOR U11802 ( .A(x[6974]), .B(y[6974]), .Z(n22751) );
  NANDN U11803 ( .A(y[6972]), .B(x[6972]), .Z(n9085) );
  NANDN U11804 ( .A(y[6973]), .B(x[6973]), .Z(n22750) );
  AND U11805 ( .A(n9085), .B(n22750), .Z(n59778) );
  XNOR U11806 ( .A(x[6972]), .B(y[6972]), .Z(n47502) );
  NANDN U11807 ( .A(y[6970]), .B(x[6970]), .Z(n9086) );
  NANDN U11808 ( .A(y[6971]), .B(x[6971]), .Z(n47501) );
  NAND U11809 ( .A(n9086), .B(n47501), .Z(n59774) );
  XNOR U11810 ( .A(x[6970]), .B(y[6970]), .Z(n22753) );
  ANDN U11811 ( .B(y[6969]), .A(x[6969]), .Z(n59772) );
  ANDN U11812 ( .B(n22753), .A(n59772), .Z(n19981) );
  XNOR U11813 ( .A(x[6968]), .B(y[6968]), .Z(n47492) );
  NANDN U11814 ( .A(y[6966]), .B(x[6966]), .Z(n9087) );
  NANDN U11815 ( .A(y[6967]), .B(x[6967]), .Z(n47491) );
  NAND U11816 ( .A(n9087), .B(n47491), .Z(n59768) );
  XNOR U11817 ( .A(x[6966]), .B(y[6966]), .Z(n22755) );
  ANDN U11818 ( .B(y[6965]), .A(x[6965]), .Z(n50900) );
  ANDN U11819 ( .B(n22755), .A(n50900), .Z(n19974) );
  NANDN U11820 ( .A(y[6964]), .B(x[6964]), .Z(n9088) );
  NANDN U11821 ( .A(y[6965]), .B(x[6965]), .Z(n22754) );
  NAND U11822 ( .A(n9088), .B(n22754), .Z(n59767) );
  XNOR U11823 ( .A(x[6964]), .B(y[6964]), .Z(n47482) );
  NANDN U11824 ( .A(y[6962]), .B(x[6962]), .Z(n9089) );
  NANDN U11825 ( .A(y[6963]), .B(x[6963]), .Z(n47481) );
  AND U11826 ( .A(n9089), .B(n47481), .Z(n59764) );
  XNOR U11827 ( .A(x[6962]), .B(y[6962]), .Z(n22757) );
  ANDN U11828 ( .B(y[6961]), .A(x[6961]), .Z(n50903) );
  ANDN U11829 ( .B(n22757), .A(n50903), .Z(n19968) );
  XNOR U11830 ( .A(x[6960]), .B(y[6960]), .Z(n47472) );
  NANDN U11831 ( .A(y[6958]), .B(x[6958]), .Z(n9090) );
  NANDN U11832 ( .A(y[6959]), .B(x[6959]), .Z(n47471) );
  AND U11833 ( .A(n9090), .B(n47471), .Z(n59762) );
  XNOR U11834 ( .A(x[6958]), .B(y[6958]), .Z(n22759) );
  ANDN U11835 ( .B(y[6957]), .A(x[6957]), .Z(n59760) );
  ANDN U11836 ( .B(n22759), .A(n59760), .Z(n19961) );
  NANDN U11837 ( .A(y[6956]), .B(x[6956]), .Z(n9091) );
  NANDN U11838 ( .A(y[6957]), .B(x[6957]), .Z(n22758) );
  NAND U11839 ( .A(n9091), .B(n22758), .Z(n59759) );
  XNOR U11840 ( .A(y[6956]), .B(x[6956]), .Z(n47462) );
  NANDN U11841 ( .A(x[6955]), .B(y[6955]), .Z(n47458) );
  AND U11842 ( .A(n47462), .B(n47458), .Z(n59758) );
  NANDN U11843 ( .A(y[6954]), .B(x[6954]), .Z(n9092) );
  NANDN U11844 ( .A(y[6955]), .B(x[6955]), .Z(n47461) );
  AND U11845 ( .A(n9092), .B(n47461), .Z(n59757) );
  ANDN U11846 ( .B(y[6953]), .A(x[6953]), .Z(n59755) );
  XNOR U11847 ( .A(x[6954]), .B(y[6954]), .Z(n22762) );
  NANDN U11848 ( .A(y[6952]), .B(x[6952]), .Z(n9093) );
  NANDN U11849 ( .A(y[6953]), .B(x[6953]), .Z(n22761) );
  AND U11850 ( .A(n9093), .B(n22761), .Z(n59754) );
  NANDN U11851 ( .A(y[6950]), .B(x[6950]), .Z(n9094) );
  NANDN U11852 ( .A(y[6951]), .B(x[6951]), .Z(n47450) );
  AND U11853 ( .A(n9094), .B(n47450), .Z(n59753) );
  ANDN U11854 ( .B(y[6949]), .A(x[6949]), .Z(n59751) );
  XNOR U11855 ( .A(x[6950]), .B(y[6950]), .Z(n22764) );
  NANDN U11856 ( .A(y[6948]), .B(x[6948]), .Z(n9095) );
  NANDN U11857 ( .A(y[6949]), .B(x[6949]), .Z(n22763) );
  AND U11858 ( .A(n9095), .B(n22763), .Z(n59750) );
  XNOR U11859 ( .A(x[6948]), .B(y[6948]), .Z(n47441) );
  NANDN U11860 ( .A(x[6947]), .B(y[6947]), .Z(n59747) );
  AND U11861 ( .A(n47441), .B(n59747), .Z(n19947) );
  NANDN U11862 ( .A(y[6946]), .B(x[6946]), .Z(n9096) );
  NANDN U11863 ( .A(y[6947]), .B(x[6947]), .Z(n47440) );
  NAND U11864 ( .A(n9096), .B(n47440), .Z(n59746) );
  XNOR U11865 ( .A(x[6946]), .B(y[6946]), .Z(n22766) );
  NANDN U11866 ( .A(y[6944]), .B(x[6944]), .Z(n9097) );
  NANDN U11867 ( .A(y[6945]), .B(x[6945]), .Z(n22765) );
  AND U11868 ( .A(n9097), .B(n22765), .Z(n59743) );
  XNOR U11869 ( .A(x[6944]), .B(y[6944]), .Z(n47431) );
  NANDN U11870 ( .A(x[6943]), .B(y[6943]), .Z(n59741) );
  AND U11871 ( .A(n47431), .B(n59741), .Z(n19941) );
  XNOR U11872 ( .A(x[6942]), .B(y[6942]), .Z(n22768) );
  NANDN U11873 ( .A(y[6940]), .B(x[6940]), .Z(n9098) );
  NANDN U11874 ( .A(y[6941]), .B(x[6941]), .Z(n22767) );
  AND U11875 ( .A(n9098), .B(n22767), .Z(n59737) );
  XNOR U11876 ( .A(y[6940]), .B(x[6940]), .Z(n47421) );
  NANDN U11877 ( .A(x[6939]), .B(y[6939]), .Z(n47417) );
  AND U11878 ( .A(n47421), .B(n47417), .Z(n59736) );
  NANDN U11879 ( .A(y[6938]), .B(x[6938]), .Z(n9099) );
  NANDN U11880 ( .A(y[6939]), .B(x[6939]), .Z(n47420) );
  AND U11881 ( .A(n9099), .B(n47420), .Z(n59735) );
  XNOR U11882 ( .A(x[6938]), .B(y[6938]), .Z(n22771) );
  NANDN U11883 ( .A(y[6936]), .B(x[6936]), .Z(n9100) );
  NANDN U11884 ( .A(y[6937]), .B(x[6937]), .Z(n22770) );
  AND U11885 ( .A(n9100), .B(n22770), .Z(n59734) );
  XNOR U11886 ( .A(x[6936]), .B(y[6936]), .Z(n47410) );
  NANDN U11887 ( .A(y[6934]), .B(x[6934]), .Z(n9101) );
  NANDN U11888 ( .A(y[6935]), .B(x[6935]), .Z(n47409) );
  AND U11889 ( .A(n9101), .B(n47409), .Z(n59729) );
  XNOR U11890 ( .A(x[6932]), .B(y[6932]), .Z(n47400) );
  NANDN U11891 ( .A(y[6930]), .B(x[6930]), .Z(n9102) );
  NANDN U11892 ( .A(y[6931]), .B(x[6931]), .Z(n47399) );
  AND U11893 ( .A(n9102), .B(n47399), .Z(n59725) );
  XNOR U11894 ( .A(x[6930]), .B(y[6930]), .Z(n22775) );
  NANDN U11895 ( .A(x[6929]), .B(y[6929]), .Z(n59723) );
  AND U11896 ( .A(n22775), .B(n59723), .Z(n19919) );
  NANDN U11897 ( .A(y[6928]), .B(x[6928]), .Z(n9103) );
  NANDN U11898 ( .A(y[6929]), .B(x[6929]), .Z(n22774) );
  NAND U11899 ( .A(n9103), .B(n22774), .Z(n59722) );
  XNOR U11900 ( .A(x[6928]), .B(y[6928]), .Z(n22777) );
  NANDN U11901 ( .A(y[6926]), .B(x[6926]), .Z(n9104) );
  NANDN U11902 ( .A(y[6927]), .B(x[6927]), .Z(n22776) );
  AND U11903 ( .A(n9104), .B(n22776), .Z(n59721) );
  XNOR U11904 ( .A(x[6926]), .B(y[6926]), .Z(n22779) );
  NANDN U11905 ( .A(y[6924]), .B(x[6924]), .Z(n9105) );
  NANDN U11906 ( .A(y[6925]), .B(x[6925]), .Z(n22778) );
  AND U11907 ( .A(n9105), .B(n22778), .Z(n59718) );
  NANDN U11908 ( .A(y[6922]), .B(x[6922]), .Z(n9106) );
  NANDN U11909 ( .A(y[6923]), .B(x[6923]), .Z(n47381) );
  AND U11910 ( .A(n9106), .B(n47381), .Z(n59716) );
  ANDN U11911 ( .B(y[6921]), .A(x[6921]), .Z(n59714) );
  XNOR U11912 ( .A(x[6922]), .B(y[6922]), .Z(n22781) );
  NANDN U11913 ( .A(y[6920]), .B(x[6920]), .Z(n9107) );
  NANDN U11914 ( .A(y[6921]), .B(x[6921]), .Z(n22780) );
  AND U11915 ( .A(n9107), .B(n22780), .Z(n59713) );
  ANDN U11916 ( .B(y[6917]), .A(x[6917]), .Z(n59708) );
  XNOR U11917 ( .A(x[6918]), .B(y[6918]), .Z(n22783) );
  NANDN U11918 ( .A(y[6916]), .B(x[6916]), .Z(n9108) );
  NANDN U11919 ( .A(y[6917]), .B(x[6917]), .Z(n22782) );
  NAND U11920 ( .A(n9108), .B(n22782), .Z(n59707) );
  XNOR U11921 ( .A(x[6916]), .B(y[6916]), .Z(n47362) );
  NANDN U11922 ( .A(x[6915]), .B(y[6915]), .Z(n59705) );
  AND U11923 ( .A(n47362), .B(n59705), .Z(n19897) );
  XNOR U11924 ( .A(x[6914]), .B(y[6914]), .Z(n22785) );
  NANDN U11925 ( .A(y[6912]), .B(x[6912]), .Z(n9109) );
  NANDN U11926 ( .A(y[6913]), .B(x[6913]), .Z(n22784) );
  AND U11927 ( .A(n9109), .B(n22784), .Z(n59703) );
  XNOR U11928 ( .A(x[6912]), .B(y[6912]), .Z(n47352) );
  NANDN U11929 ( .A(x[6911]), .B(y[6911]), .Z(n59699) );
  NAND U11930 ( .A(n47352), .B(n59699), .Z(n19890) );
  NANDN U11931 ( .A(y[6910]), .B(x[6910]), .Z(n9110) );
  NANDN U11932 ( .A(y[6911]), .B(x[6911]), .Z(n47351) );
  AND U11933 ( .A(n9110), .B(n47351), .Z(n59698) );
  ANDN U11934 ( .B(y[6909]), .A(x[6909]), .Z(n59696) );
  XNOR U11935 ( .A(x[6910]), .B(y[6910]), .Z(n22787) );
  NANDN U11936 ( .A(n59696), .B(n22787), .Z(n19887) );
  NANDN U11937 ( .A(x[6907]), .B(y[6907]), .Z(n47338) );
  IV U11938 ( .A(n47338), .Z(n59695) );
  XNOR U11939 ( .A(x[6908]), .B(y[6908]), .Z(n47342) );
  XNOR U11940 ( .A(x[6906]), .B(y[6906]), .Z(n22789) );
  NANDN U11941 ( .A(y[6904]), .B(x[6904]), .Z(n9111) );
  NANDN U11942 ( .A(y[6905]), .B(x[6905]), .Z(n22788) );
  AND U11943 ( .A(n9111), .B(n22788), .Z(n59692) );
  XNOR U11944 ( .A(x[6904]), .B(y[6904]), .Z(n47331) );
  NANDN U11945 ( .A(y[6902]), .B(x[6902]), .Z(n22792) );
  NANDN U11946 ( .A(y[6903]), .B(x[6903]), .Z(n47330) );
  NAND U11947 ( .A(n22792), .B(n47330), .Z(n59689) );
  NANDN U11948 ( .A(x[6902]), .B(y[6902]), .Z(n22791) );
  ANDN U11949 ( .B(y[6901]), .A(x[6901]), .Z(n22794) );
  ANDN U11950 ( .B(n22791), .A(n22794), .Z(n59688) );
  NANDN U11951 ( .A(y[6900]), .B(x[6900]), .Z(n9112) );
  NANDN U11952 ( .A(y[6901]), .B(x[6901]), .Z(n22793) );
  NAND U11953 ( .A(n9112), .B(n22793), .Z(n59687) );
  XNOR U11954 ( .A(x[6900]), .B(y[6900]), .Z(n47321) );
  NANDN U11955 ( .A(y[6898]), .B(x[6898]), .Z(n9113) );
  NANDN U11956 ( .A(y[6899]), .B(x[6899]), .Z(n47320) );
  AND U11957 ( .A(n9113), .B(n47320), .Z(n59682) );
  ANDN U11958 ( .B(y[6897]), .A(x[6897]), .Z(n50923) );
  XNOR U11959 ( .A(x[6898]), .B(y[6898]), .Z(n22796) );
  NANDN U11960 ( .A(n50923), .B(n22796), .Z(n19868) );
  NANDN U11961 ( .A(y[6896]), .B(x[6896]), .Z(n9114) );
  NANDN U11962 ( .A(y[6897]), .B(x[6897]), .Z(n22795) );
  AND U11963 ( .A(n9114), .B(n22795), .Z(n59681) );
  XNOR U11964 ( .A(x[6896]), .B(y[6896]), .Z(n47311) );
  NANDN U11965 ( .A(x[6895]), .B(y[6895]), .Z(n59679) );
  NAND U11966 ( .A(n47311), .B(n59679), .Z(n19865) );
  NANDN U11967 ( .A(y[6894]), .B(x[6894]), .Z(n9115) );
  NANDN U11968 ( .A(y[6895]), .B(x[6895]), .Z(n47310) );
  AND U11969 ( .A(n9115), .B(n47310), .Z(n59678) );
  ANDN U11970 ( .B(y[6893]), .A(x[6893]), .Z(n59676) );
  XNOR U11971 ( .A(x[6894]), .B(y[6894]), .Z(n22798) );
  NANDN U11972 ( .A(y[6892]), .B(x[6892]), .Z(n9116) );
  NANDN U11973 ( .A(y[6893]), .B(x[6893]), .Z(n22797) );
  NAND U11974 ( .A(n9116), .B(n22797), .Z(n59675) );
  XNOR U11975 ( .A(x[6892]), .B(y[6892]), .Z(n47301) );
  NANDN U11976 ( .A(y[6890]), .B(x[6890]), .Z(n9117) );
  NANDN U11977 ( .A(y[6891]), .B(x[6891]), .Z(n47300) );
  AND U11978 ( .A(n9117), .B(n47300), .Z(n59673) );
  XNOR U11979 ( .A(x[6888]), .B(y[6888]), .Z(n47291) );
  ANDN U11980 ( .B(y[6887]), .A(x[6887]), .Z(n47287) );
  ANDN U11981 ( .B(n47291), .A(n47287), .Z(n19852) );
  XNOR U11982 ( .A(x[6886]), .B(y[6886]), .Z(n22802) );
  NANDN U11983 ( .A(y[6884]), .B(x[6884]), .Z(n9118) );
  NANDN U11984 ( .A(y[6885]), .B(x[6885]), .Z(n22801) );
  AND U11985 ( .A(n9118), .B(n22801), .Z(n59665) );
  NANDN U11986 ( .A(x[6883]), .B(y[6883]), .Z(n47276) );
  IV U11987 ( .A(n47276), .Z(n50930) );
  XNOR U11988 ( .A(x[6884]), .B(y[6884]), .Z(n47280) );
  NANDN U11989 ( .A(y[6882]), .B(x[6882]), .Z(n9119) );
  NANDN U11990 ( .A(y[6883]), .B(x[6883]), .Z(n47279) );
  NAND U11991 ( .A(n9119), .B(n47279), .Z(n59664) );
  NANDN U11992 ( .A(y[6880]), .B(x[6880]), .Z(n9120) );
  NANDN U11993 ( .A(y[6881]), .B(x[6881]), .Z(n22803) );
  AND U11994 ( .A(n9120), .B(n22803), .Z(n59661) );
  XNOR U11995 ( .A(x[6880]), .B(y[6880]), .Z(n47269) );
  NANDN U11996 ( .A(y[6878]), .B(x[6878]), .Z(n9121) );
  NANDN U11997 ( .A(y[6879]), .B(x[6879]), .Z(n47268) );
  NAND U11998 ( .A(n9121), .B(n47268), .Z(n59658) );
  XNOR U11999 ( .A(x[6878]), .B(y[6878]), .Z(n22806) );
  NANDN U12000 ( .A(x[6877]), .B(y[6877]), .Z(n59656) );
  AND U12001 ( .A(n22806), .B(n59656), .Z(n19836) );
  XNOR U12002 ( .A(x[6876]), .B(y[6876]), .Z(n22808) );
  NANDN U12003 ( .A(y[6874]), .B(x[6874]), .Z(n9122) );
  NANDN U12004 ( .A(y[6875]), .B(x[6875]), .Z(n22807) );
  AND U12005 ( .A(n9122), .B(n22807), .Z(n59651) );
  XNOR U12006 ( .A(x[6874]), .B(y[6874]), .Z(n22810) );
  NANDN U12007 ( .A(x[6873]), .B(y[6873]), .Z(n50931) );
  NAND U12008 ( .A(n22810), .B(n50931), .Z(n19829) );
  NANDN U12009 ( .A(y[6872]), .B(x[6872]), .Z(n9123) );
  NANDN U12010 ( .A(y[6873]), .B(x[6873]), .Z(n22809) );
  AND U12011 ( .A(n9123), .B(n22809), .Z(n59650) );
  XOR U12012 ( .A(x[6872]), .B(y[6872]), .Z(n47253) );
  NANDN U12013 ( .A(x[6871]), .B(y[6871]), .Z(n59648) );
  NANDN U12014 ( .A(n47253), .B(n59648), .Z(n19826) );
  NANDN U12015 ( .A(y[6870]), .B(x[6870]), .Z(n9124) );
  ANDN U12016 ( .B(x[6871]), .A(y[6871]), .Z(n47251) );
  ANDN U12017 ( .B(n9124), .A(n47251), .Z(n59647) );
  XNOR U12018 ( .A(x[6870]), .B(y[6870]), .Z(n22812) );
  NANDN U12019 ( .A(y[6868]), .B(x[6868]), .Z(n9125) );
  NANDN U12020 ( .A(y[6869]), .B(x[6869]), .Z(n22811) );
  NAND U12021 ( .A(n9125), .B(n22811), .Z(n59646) );
  NANDN U12022 ( .A(y[6866]), .B(x[6866]), .Z(n9126) );
  NANDN U12023 ( .A(y[6867]), .B(x[6867]), .Z(n47240) );
  AND U12024 ( .A(n9126), .B(n47240), .Z(n59643) );
  XNOR U12025 ( .A(x[6866]), .B(y[6866]), .Z(n22814) );
  NANDN U12026 ( .A(y[6864]), .B(x[6864]), .Z(n9127) );
  NANDN U12027 ( .A(y[6865]), .B(x[6865]), .Z(n22813) );
  NAND U12028 ( .A(n9127), .B(n22813), .Z(n59639) );
  XNOR U12029 ( .A(x[6864]), .B(y[6864]), .Z(n22816) );
  NANDN U12030 ( .A(x[6863]), .B(y[6863]), .Z(n59637) );
  AND U12031 ( .A(n22816), .B(n59637), .Z(n19814) );
  XNOR U12032 ( .A(x[6862]), .B(y[6862]), .Z(n22818) );
  NANDN U12033 ( .A(y[6860]), .B(x[6860]), .Z(n9128) );
  NANDN U12034 ( .A(y[6861]), .B(x[6861]), .Z(n22817) );
  AND U12035 ( .A(n9128), .B(n22817), .Z(n59633) );
  XNOR U12036 ( .A(x[6860]), .B(y[6860]), .Z(n47223) );
  NANDN U12037 ( .A(x[6859]), .B(y[6859]), .Z(n50936) );
  AND U12038 ( .A(n47223), .B(n50936), .Z(n19807) );
  NANDN U12039 ( .A(y[6858]), .B(x[6858]), .Z(n9129) );
  NANDN U12040 ( .A(y[6859]), .B(x[6859]), .Z(n47222) );
  NAND U12041 ( .A(n9129), .B(n47222), .Z(n59632) );
  XNOR U12042 ( .A(x[6858]), .B(y[6858]), .Z(n22820) );
  NANDN U12043 ( .A(x[6857]), .B(y[6857]), .Z(n59630) );
  XNOR U12044 ( .A(x[6856]), .B(y[6856]), .Z(n22822) );
  NANDN U12045 ( .A(y[6854]), .B(x[6854]), .Z(n9130) );
  NANDN U12046 ( .A(y[6855]), .B(x[6855]), .Z(n22821) );
  NAND U12047 ( .A(n9130), .B(n22821), .Z(n59628) );
  XNOR U12048 ( .A(y[6854]), .B(x[6854]), .Z(n22825) );
  NANDN U12049 ( .A(x[6853]), .B(y[6853]), .Z(n47208) );
  AND U12050 ( .A(n22825), .B(n47208), .Z(n59627) );
  XNOR U12051 ( .A(x[6852]), .B(y[6852]), .Z(n22827) );
  NANDN U12052 ( .A(y[6850]), .B(x[6850]), .Z(n9131) );
  NANDN U12053 ( .A(y[6851]), .B(x[6851]), .Z(n22826) );
  AND U12054 ( .A(n9131), .B(n22826), .Z(n59622) );
  ANDN U12055 ( .B(y[6849]), .A(x[6849]), .Z(n59620) );
  XNOR U12056 ( .A(x[6850]), .B(y[6850]), .Z(n22829) );
  NANDN U12057 ( .A(n59620), .B(n22829), .Z(n19791) );
  NANDN U12058 ( .A(y[6848]), .B(x[6848]), .Z(n9132) );
  NANDN U12059 ( .A(y[6849]), .B(x[6849]), .Z(n22828) );
  AND U12060 ( .A(n9132), .B(n22828), .Z(n59619) );
  XNOR U12061 ( .A(x[6848]), .B(y[6848]), .Z(n47196) );
  NANDN U12062 ( .A(x[6847]), .B(y[6847]), .Z(n59617) );
  NAND U12063 ( .A(n47196), .B(n59617), .Z(n19788) );
  XNOR U12064 ( .A(x[6846]), .B(y[6846]), .Z(n22831) );
  NANDN U12065 ( .A(y[6844]), .B(x[6844]), .Z(n9133) );
  NANDN U12066 ( .A(y[6845]), .B(x[6845]), .Z(n22830) );
  NAND U12067 ( .A(n9133), .B(n22830), .Z(n59616) );
  XNOR U12068 ( .A(x[6844]), .B(y[6844]), .Z(n22833) );
  NANDN U12069 ( .A(y[6842]), .B(x[6842]), .Z(n9134) );
  NANDN U12070 ( .A(y[6843]), .B(x[6843]), .Z(n22832) );
  AND U12071 ( .A(n9134), .B(n22832), .Z(n59613) );
  ANDN U12072 ( .B(y[6841]), .A(x[6841]), .Z(n50943) );
  XNOR U12073 ( .A(x[6842]), .B(y[6842]), .Z(n22835) );
  NANDN U12074 ( .A(y[6840]), .B(x[6840]), .Z(n9135) );
  NANDN U12075 ( .A(y[6841]), .B(x[6841]), .Z(n22834) );
  NAND U12076 ( .A(n9135), .B(n22834), .Z(n50944) );
  XNOR U12077 ( .A(x[6840]), .B(y[6840]), .Z(n47178) );
  NANDN U12078 ( .A(x[6839]), .B(y[6839]), .Z(n50946) );
  AND U12079 ( .A(n47178), .B(n50946), .Z(n19775) );
  XNOR U12080 ( .A(y[6838]), .B(x[6838]), .Z(n22837) );
  ANDN U12081 ( .B(y[6837]), .A(x[6837]), .Z(n22838) );
  ANDN U12082 ( .B(n22837), .A(n22838), .Z(n59609) );
  NANDN U12083 ( .A(y[6836]), .B(x[6836]), .Z(n9136) );
  NANDN U12084 ( .A(y[6837]), .B(x[6837]), .Z(n22836) );
  AND U12085 ( .A(n9136), .B(n22836), .Z(n59608) );
  XNOR U12086 ( .A(x[6836]), .B(y[6836]), .Z(n47167) );
  ANDN U12087 ( .B(y[6835]), .A(x[6835]), .Z(n47163) );
  ANDN U12088 ( .B(n47167), .A(n47163), .Z(n19769) );
  XNOR U12089 ( .A(x[6834]), .B(y[6834]), .Z(n22840) );
  NANDN U12090 ( .A(y[6832]), .B(x[6832]), .Z(n9137) );
  NANDN U12091 ( .A(y[6833]), .B(x[6833]), .Z(n22839) );
  AND U12092 ( .A(n9137), .B(n22839), .Z(n59604) );
  NANDN U12093 ( .A(x[6831]), .B(y[6831]), .Z(n47152) );
  IV U12094 ( .A(n47152), .Z(n50950) );
  XNOR U12095 ( .A(x[6832]), .B(y[6832]), .Z(n47156) );
  NANDN U12096 ( .A(y[6830]), .B(x[6830]), .Z(n9138) );
  NANDN U12097 ( .A(y[6831]), .B(x[6831]), .Z(n47155) );
  NAND U12098 ( .A(n9138), .B(n47155), .Z(n59603) );
  NANDN U12099 ( .A(y[6828]), .B(x[6828]), .Z(n9139) );
  NANDN U12100 ( .A(y[6829]), .B(x[6829]), .Z(n22841) );
  AND U12101 ( .A(n9139), .B(n22841), .Z(n59600) );
  XNOR U12102 ( .A(x[6828]), .B(y[6828]), .Z(n47145) );
  NANDN U12103 ( .A(y[6826]), .B(x[6826]), .Z(n9140) );
  NANDN U12104 ( .A(y[6827]), .B(x[6827]), .Z(n47144) );
  NAND U12105 ( .A(n9140), .B(n47144), .Z(n59596) );
  XNOR U12106 ( .A(x[6826]), .B(y[6826]), .Z(n22844) );
  ANDN U12107 ( .B(y[6825]), .A(x[6825]), .Z(n59594) );
  ANDN U12108 ( .B(n22844), .A(n59594), .Z(n19753) );
  NANDN U12109 ( .A(y[6824]), .B(x[6824]), .Z(n9141) );
  NANDN U12110 ( .A(y[6825]), .B(x[6825]), .Z(n22843) );
  NAND U12111 ( .A(n9141), .B(n22843), .Z(n59593) );
  XNOR U12112 ( .A(x[6824]), .B(y[6824]), .Z(n47135) );
  NANDN U12113 ( .A(y[6822]), .B(x[6822]), .Z(n9142) );
  NANDN U12114 ( .A(y[6823]), .B(x[6823]), .Z(n47134) );
  AND U12115 ( .A(n9142), .B(n47134), .Z(n59590) );
  XNOR U12116 ( .A(x[6822]), .B(y[6822]), .Z(n22846) );
  NANDN U12117 ( .A(x[6821]), .B(y[6821]), .Z(n22847) );
  AND U12118 ( .A(n22846), .B(n22847), .Z(n19747) );
  XNOR U12119 ( .A(x[6820]), .B(y[6820]), .Z(n47125) );
  NANDN U12120 ( .A(y[6818]), .B(x[6818]), .Z(n9143) );
  NANDN U12121 ( .A(y[6819]), .B(x[6819]), .Z(n47124) );
  AND U12122 ( .A(n9143), .B(n47124), .Z(n59586) );
  XNOR U12123 ( .A(x[6818]), .B(y[6818]), .Z(n22849) );
  NANDN U12124 ( .A(x[6817]), .B(y[6817]), .Z(n59584) );
  NANDN U12125 ( .A(y[6816]), .B(x[6816]), .Z(n9144) );
  NANDN U12126 ( .A(y[6817]), .B(x[6817]), .Z(n22848) );
  NAND U12127 ( .A(n9144), .B(n22848), .Z(n59583) );
  NANDN U12128 ( .A(y[6814]), .B(x[6814]), .Z(n9145) );
  NANDN U12129 ( .A(y[6815]), .B(x[6815]), .Z(n22850) );
  AND U12130 ( .A(n9145), .B(n22850), .Z(n59579) );
  ANDN U12131 ( .B(y[6813]), .A(x[6813]), .Z(n59577) );
  XNOR U12132 ( .A(x[6814]), .B(y[6814]), .Z(n22853) );
  NANDN U12133 ( .A(y[6812]), .B(x[6812]), .Z(n9146) );
  NANDN U12134 ( .A(y[6813]), .B(x[6813]), .Z(n22852) );
  NAND U12135 ( .A(n9146), .B(n22852), .Z(n59576) );
  NANDN U12136 ( .A(y[6810]), .B(x[6810]), .Z(n9147) );
  NANDN U12137 ( .A(y[6811]), .B(x[6811]), .Z(n47106) );
  AND U12138 ( .A(n9147), .B(n47106), .Z(n59573) );
  ANDN U12139 ( .B(y[6809]), .A(x[6809]), .Z(n59571) );
  XNOR U12140 ( .A(x[6810]), .B(y[6810]), .Z(n22855) );
  NANDN U12141 ( .A(y[6808]), .B(x[6808]), .Z(n9148) );
  NANDN U12142 ( .A(y[6809]), .B(x[6809]), .Z(n22854) );
  NAND U12143 ( .A(n9148), .B(n22854), .Z(n50953) );
  NANDN U12144 ( .A(x[6807]), .B(y[6807]), .Z(n47097) );
  NANDN U12145 ( .A(x[6808]), .B(y[6808]), .Z(n22856) );
  AND U12146 ( .A(n47097), .B(n22856), .Z(n59570) );
  NANDN U12147 ( .A(x[6806]), .B(y[6806]), .Z(n47094) );
  ANDN U12148 ( .B(y[6805]), .A(x[6805]), .Z(n22857) );
  ANDN U12149 ( .B(n47094), .A(n22857), .Z(n59568) );
  XNOR U12150 ( .A(x[6804]), .B(y[6804]), .Z(n47086) );
  NANDN U12151 ( .A(y[6802]), .B(x[6802]), .Z(n9149) );
  NANDN U12152 ( .A(y[6803]), .B(x[6803]), .Z(n47085) );
  NAND U12153 ( .A(n9149), .B(n47085), .Z(n59564) );
  XNOR U12154 ( .A(x[6802]), .B(y[6802]), .Z(n22859) );
  ANDN U12155 ( .B(y[6801]), .A(x[6801]), .Z(n59561) );
  NANDN U12156 ( .A(y[6800]), .B(x[6800]), .Z(n9150) );
  NANDN U12157 ( .A(y[6801]), .B(x[6801]), .Z(n22858) );
  AND U12158 ( .A(n9150), .B(n22858), .Z(n59560) );
  XNOR U12159 ( .A(x[6800]), .B(y[6800]), .Z(n47076) );
  NANDN U12160 ( .A(y[6798]), .B(x[6798]), .Z(n9151) );
  NANDN U12161 ( .A(y[6799]), .B(x[6799]), .Z(n47075) );
  AND U12162 ( .A(n9151), .B(n47075), .Z(n59557) );
  ANDN U12163 ( .B(y[6797]), .A(x[6797]), .Z(n50954) );
  XNOR U12164 ( .A(x[6798]), .B(y[6798]), .Z(n22861) );
  NANDN U12165 ( .A(n50954), .B(n22861), .Z(n19709) );
  NANDN U12166 ( .A(y[6796]), .B(x[6796]), .Z(n9152) );
  NANDN U12167 ( .A(y[6797]), .B(x[6797]), .Z(n22860) );
  AND U12168 ( .A(n9152), .B(n22860), .Z(n59556) );
  XNOR U12169 ( .A(x[6796]), .B(y[6796]), .Z(n47066) );
  NANDN U12170 ( .A(x[6795]), .B(y[6795]), .Z(n59554) );
  NAND U12171 ( .A(n47066), .B(n59554), .Z(n19706) );
  NANDN U12172 ( .A(y[6794]), .B(x[6794]), .Z(n9153) );
  NANDN U12173 ( .A(y[6795]), .B(x[6795]), .Z(n47065) );
  AND U12174 ( .A(n9153), .B(n47065), .Z(n59553) );
  XNOR U12175 ( .A(x[6794]), .B(y[6794]), .Z(n22863) );
  NANDN U12176 ( .A(y[6792]), .B(x[6792]), .Z(n9154) );
  NANDN U12177 ( .A(y[6793]), .B(x[6793]), .Z(n22862) );
  NAND U12178 ( .A(n9154), .B(n22862), .Z(n59552) );
  NANDN U12179 ( .A(y[6790]), .B(x[6790]), .Z(n9155) );
  NANDN U12180 ( .A(y[6791]), .B(x[6791]), .Z(n22864) );
  AND U12181 ( .A(n9155), .B(n22864), .Z(n59547) );
  ANDN U12182 ( .B(y[6789]), .A(x[6789]), .Z(n59545) );
  XNOR U12183 ( .A(x[6790]), .B(y[6790]), .Z(n22867) );
  NANDN U12184 ( .A(y[6788]), .B(x[6788]), .Z(n9156) );
  NANDN U12185 ( .A(y[6789]), .B(x[6789]), .Z(n22866) );
  NAND U12186 ( .A(n9156), .B(n22866), .Z(n59544) );
  XNOR U12187 ( .A(x[6788]), .B(y[6788]), .Z(n47048) );
  NANDN U12188 ( .A(x[6787]), .B(y[6787]), .Z(n59543) );
  AND U12189 ( .A(n47048), .B(n59543), .Z(n19694) );
  XNOR U12190 ( .A(x[6786]), .B(y[6786]), .Z(n22869) );
  NANDN U12191 ( .A(y[6784]), .B(x[6784]), .Z(n9157) );
  NANDN U12192 ( .A(y[6785]), .B(x[6785]), .Z(n22868) );
  AND U12193 ( .A(n9157), .B(n22868), .Z(n59539) );
  XNOR U12194 ( .A(x[6784]), .B(y[6784]), .Z(n47038) );
  NANDN U12195 ( .A(x[6783]), .B(y[6783]), .Z(n50960) );
  AND U12196 ( .A(n47038), .B(n50960), .Z(n19687) );
  XNOR U12197 ( .A(x[6782]), .B(y[6782]), .Z(n22871) );
  NANDN U12198 ( .A(y[6780]), .B(x[6780]), .Z(n9158) );
  NANDN U12199 ( .A(y[6781]), .B(x[6781]), .Z(n22870) );
  AND U12200 ( .A(n9158), .B(n22870), .Z(n59535) );
  NANDN U12201 ( .A(x[6779]), .B(y[6779]), .Z(n50962) );
  XNOR U12202 ( .A(x[6780]), .B(y[6780]), .Z(n47028) );
  AND U12203 ( .A(n50962), .B(n47028), .Z(n19680) );
  XNOR U12204 ( .A(x[6778]), .B(y[6778]), .Z(n22873) );
  NANDN U12205 ( .A(y[6776]), .B(x[6776]), .Z(n9159) );
  NANDN U12206 ( .A(y[6777]), .B(x[6777]), .Z(n22872) );
  AND U12207 ( .A(n9159), .B(n22872), .Z(n59529) );
  XNOR U12208 ( .A(x[6776]), .B(y[6776]), .Z(n47018) );
  NANDN U12209 ( .A(y[6774]), .B(x[6774]), .Z(n9160) );
  NANDN U12210 ( .A(y[6775]), .B(x[6775]), .Z(n47017) );
  NAND U12211 ( .A(n9160), .B(n47017), .Z(n59526) );
  NANDN U12212 ( .A(y[6772]), .B(x[6772]), .Z(n9161) );
  NANDN U12213 ( .A(y[6773]), .B(x[6773]), .Z(n22874) );
  AND U12214 ( .A(n9161), .B(n22874), .Z(n59523) );
  XNOR U12215 ( .A(x[6772]), .B(y[6772]), .Z(n22877) );
  NANDN U12216 ( .A(y[6770]), .B(x[6770]), .Z(n9162) );
  NANDN U12217 ( .A(y[6771]), .B(x[6771]), .Z(n22876) );
  NAND U12218 ( .A(n9162), .B(n22876), .Z(n59520) );
  XNOR U12219 ( .A(x[6770]), .B(y[6770]), .Z(n22879) );
  ANDN U12220 ( .B(y[6769]), .A(x[6769]), .Z(n50963) );
  ANDN U12221 ( .B(n22879), .A(n50963), .Z(n19664) );
  NANDN U12222 ( .A(y[6768]), .B(x[6768]), .Z(n9163) );
  NANDN U12223 ( .A(y[6769]), .B(x[6769]), .Z(n22878) );
  NAND U12224 ( .A(n9163), .B(n22878), .Z(n59519) );
  XNOR U12225 ( .A(x[6768]), .B(y[6768]), .Z(n47000) );
  NANDN U12226 ( .A(y[6766]), .B(x[6766]), .Z(n9164) );
  NANDN U12227 ( .A(y[6767]), .B(x[6767]), .Z(n46999) );
  AND U12228 ( .A(n9164), .B(n46999), .Z(n59516) );
  NANDN U12229 ( .A(x[6765]), .B(y[6765]), .Z(n22882) );
  XNOR U12230 ( .A(x[6766]), .B(y[6766]), .Z(n22881) );
  NAND U12231 ( .A(n22882), .B(n22881), .Z(n19658) );
  NANDN U12232 ( .A(y[6764]), .B(x[6764]), .Z(n9165) );
  NANDN U12233 ( .A(y[6765]), .B(x[6765]), .Z(n22880) );
  AND U12234 ( .A(n9165), .B(n22880), .Z(n59514) );
  XNOR U12235 ( .A(x[6764]), .B(y[6764]), .Z(n46990) );
  NANDN U12236 ( .A(x[6763]), .B(y[6763]), .Z(n59512) );
  NAND U12237 ( .A(n46990), .B(n59512), .Z(n19655) );
  NANDN U12238 ( .A(y[6762]), .B(x[6762]), .Z(n9166) );
  NANDN U12239 ( .A(y[6763]), .B(x[6763]), .Z(n46989) );
  AND U12240 ( .A(n9166), .B(n46989), .Z(n59511) );
  ANDN U12241 ( .B(y[6761]), .A(x[6761]), .Z(n59509) );
  XNOR U12242 ( .A(x[6762]), .B(y[6762]), .Z(n22884) );
  NANDN U12243 ( .A(y[6760]), .B(x[6760]), .Z(n9167) );
  NANDN U12244 ( .A(y[6761]), .B(x[6761]), .Z(n22883) );
  NAND U12245 ( .A(n9167), .B(n22883), .Z(n59508) );
  NANDN U12246 ( .A(y[6758]), .B(x[6758]), .Z(n9168) );
  NANDN U12247 ( .A(y[6759]), .B(x[6759]), .Z(n46979) );
  AND U12248 ( .A(n9168), .B(n46979), .Z(n59506) );
  ANDN U12249 ( .B(y[6757]), .A(x[6757]), .Z(n59504) );
  XNOR U12250 ( .A(x[6758]), .B(y[6758]), .Z(n22886) );
  NANDN U12251 ( .A(y[6756]), .B(x[6756]), .Z(n9169) );
  NANDN U12252 ( .A(y[6757]), .B(x[6757]), .Z(n22885) );
  NAND U12253 ( .A(n9169), .B(n22885), .Z(n59503) );
  NANDN U12254 ( .A(x[6755]), .B(y[6755]), .Z(n50969) );
  XNOR U12255 ( .A(x[6756]), .B(y[6756]), .Z(n46970) );
  XNOR U12256 ( .A(x[6754]), .B(y[6754]), .Z(n22888) );
  NANDN U12257 ( .A(y[6752]), .B(x[6752]), .Z(n9170) );
  NANDN U12258 ( .A(y[6753]), .B(x[6753]), .Z(n22887) );
  AND U12259 ( .A(n9170), .B(n22887), .Z(n59497) );
  XNOR U12260 ( .A(y[6752]), .B(x[6752]), .Z(n22891) );
  NANDN U12261 ( .A(x[6751]), .B(y[6751]), .Z(n22892) );
  AND U12262 ( .A(n22891), .B(n22892), .Z(n59496) );
  NANDN U12263 ( .A(y[6750]), .B(x[6750]), .Z(n9171) );
  NANDN U12264 ( .A(y[6751]), .B(x[6751]), .Z(n22890) );
  AND U12265 ( .A(n9171), .B(n22890), .Z(n59495) );
  ANDN U12266 ( .B(y[6749]), .A(x[6749]), .Z(n59493) );
  XNOR U12267 ( .A(x[6750]), .B(y[6750]), .Z(n22894) );
  XNOR U12268 ( .A(x[6748]), .B(y[6748]), .Z(n46952) );
  NANDN U12269 ( .A(y[6746]), .B(x[6746]), .Z(n9172) );
  NANDN U12270 ( .A(y[6747]), .B(x[6747]), .Z(n46951) );
  NAND U12271 ( .A(n9172), .B(n46951), .Z(n59489) );
  XNOR U12272 ( .A(x[6746]), .B(y[6746]), .Z(n22896) );
  NANDN U12273 ( .A(x[6745]), .B(y[6745]), .Z(n59488) );
  AND U12274 ( .A(n22896), .B(n59488), .Z(n19627) );
  XNOR U12275 ( .A(y[6744]), .B(x[6744]), .Z(n46942) );
  NANDN U12276 ( .A(y[6742]), .B(x[6742]), .Z(n9173) );
  ANDN U12277 ( .B(x[6743]), .A(y[6743]), .Z(n46944) );
  ANDN U12278 ( .B(n9173), .A(n46944), .Z(n59482) );
  XNOR U12279 ( .A(x[6742]), .B(y[6742]), .Z(n22898) );
  NANDN U12280 ( .A(x[6741]), .B(y[6741]), .Z(n22899) );
  AND U12281 ( .A(n22898), .B(n22899), .Z(n19620) );
  XNOR U12282 ( .A(x[6740]), .B(y[6740]), .Z(n46932) );
  NANDN U12283 ( .A(y[6738]), .B(x[6738]), .Z(n9174) );
  NANDN U12284 ( .A(y[6739]), .B(x[6739]), .Z(n46931) );
  AND U12285 ( .A(n9174), .B(n46931), .Z(n59478) );
  NANDN U12286 ( .A(x[6737]), .B(y[6737]), .Z(n59476) );
  XNOR U12287 ( .A(x[6738]), .B(y[6738]), .Z(n22901) );
  AND U12288 ( .A(n59476), .B(n22901), .Z(n19613) );
  NANDN U12289 ( .A(y[6736]), .B(x[6736]), .Z(n9175) );
  NANDN U12290 ( .A(y[6737]), .B(x[6737]), .Z(n22900) );
  NAND U12291 ( .A(n9175), .B(n22900), .Z(n59475) );
  XNOR U12292 ( .A(y[6736]), .B(x[6736]), .Z(n22904) );
  NANDN U12293 ( .A(x[6735]), .B(y[6735]), .Z(n46920) );
  AND U12294 ( .A(n22904), .B(n46920), .Z(n59474) );
  NANDN U12295 ( .A(y[6734]), .B(x[6734]), .Z(n9176) );
  NANDN U12296 ( .A(y[6735]), .B(x[6735]), .Z(n22903) );
  AND U12297 ( .A(n9176), .B(n22903), .Z(n59473) );
  ANDN U12298 ( .B(y[6733]), .A(x[6733]), .Z(n59471) );
  XNOR U12299 ( .A(x[6734]), .B(y[6734]), .Z(n22906) );
  NANDN U12300 ( .A(y[6732]), .B(x[6732]), .Z(n9177) );
  NANDN U12301 ( .A(y[6733]), .B(x[6733]), .Z(n22905) );
  NAND U12302 ( .A(n9177), .B(n22905), .Z(n50972) );
  NANDN U12303 ( .A(y[6730]), .B(x[6730]), .Z(n9178) );
  NANDN U12304 ( .A(y[6731]), .B(x[6731]), .Z(n46912) );
  AND U12305 ( .A(n9178), .B(n46912), .Z(n59469) );
  ANDN U12306 ( .B(y[6729]), .A(x[6729]), .Z(n59467) );
  XNOR U12307 ( .A(x[6730]), .B(y[6730]), .Z(n22908) );
  NANDN U12308 ( .A(y[6728]), .B(x[6728]), .Z(n9179) );
  NANDN U12309 ( .A(y[6729]), .B(x[6729]), .Z(n22907) );
  AND U12310 ( .A(n9179), .B(n22907), .Z(n59466) );
  XNOR U12311 ( .A(x[6728]), .B(y[6728]), .Z(n46903) );
  NANDN U12312 ( .A(x[6727]), .B(y[6727]), .Z(n59464) );
  AND U12313 ( .A(n46903), .B(n59464), .Z(n19599) );
  NANDN U12314 ( .A(y[6726]), .B(x[6726]), .Z(n9180) );
  NANDN U12315 ( .A(y[6727]), .B(x[6727]), .Z(n46902) );
  NAND U12316 ( .A(n9180), .B(n46902), .Z(n59463) );
  XNOR U12317 ( .A(x[6726]), .B(y[6726]), .Z(n22910) );
  NANDN U12318 ( .A(y[6724]), .B(x[6724]), .Z(n9181) );
  NANDN U12319 ( .A(y[6725]), .B(x[6725]), .Z(n22909) );
  AND U12320 ( .A(n9181), .B(n22909), .Z(n59460) );
  XNOR U12321 ( .A(x[6724]), .B(y[6724]), .Z(n22912) );
  NANDN U12322 ( .A(x[6723]), .B(y[6723]), .Z(n59458) );
  AND U12323 ( .A(n22912), .B(n59458), .Z(n19593) );
  XNOR U12324 ( .A(x[6722]), .B(y[6722]), .Z(n22914) );
  NANDN U12325 ( .A(y[6720]), .B(x[6720]), .Z(n9182) );
  NANDN U12326 ( .A(y[6721]), .B(x[6721]), .Z(n22913) );
  AND U12327 ( .A(n9182), .B(n22913), .Z(n59456) );
  ANDN U12328 ( .B(y[6719]), .A(x[6719]), .Z(n22915) );
  NANDN U12329 ( .A(y[6718]), .B(x[6718]), .Z(n22917) );
  NANDN U12330 ( .A(y[6719]), .B(x[6719]), .Z(n46884) );
  AND U12331 ( .A(n22917), .B(n46884), .Z(n59453) );
  NANDN U12332 ( .A(x[6717]), .B(y[6717]), .Z(n22919) );
  NANDN U12333 ( .A(x[6718]), .B(y[6718]), .Z(n22916) );
  NAND U12334 ( .A(n22919), .B(n22916), .Z(n59451) );
  NANDN U12335 ( .A(y[6716]), .B(x[6716]), .Z(n9183) );
  NANDN U12336 ( .A(y[6717]), .B(x[6717]), .Z(n22918) );
  AND U12337 ( .A(n9183), .B(n22918), .Z(n59450) );
  XNOR U12338 ( .A(x[6716]), .B(y[6716]), .Z(n22921) );
  NANDN U12339 ( .A(y[6714]), .B(x[6714]), .Z(n9184) );
  NANDN U12340 ( .A(y[6715]), .B(x[6715]), .Z(n22920) );
  NAND U12341 ( .A(n9184), .B(n22920), .Z(n59449) );
  XNOR U12342 ( .A(x[6714]), .B(y[6714]), .Z(n22923) );
  ANDN U12343 ( .B(y[6713]), .A(x[6713]), .Z(n59447) );
  ANDN U12344 ( .B(n22923), .A(n59447), .Z(n19578) );
  NANDN U12345 ( .A(y[6712]), .B(x[6712]), .Z(n9185) );
  NANDN U12346 ( .A(y[6713]), .B(x[6713]), .Z(n22922) );
  NAND U12347 ( .A(n9185), .B(n22922), .Z(n59446) );
  XNOR U12348 ( .A(x[6712]), .B(y[6712]), .Z(n46867) );
  NANDN U12349 ( .A(y[6710]), .B(x[6710]), .Z(n9186) );
  NANDN U12350 ( .A(y[6711]), .B(x[6711]), .Z(n46866) );
  AND U12351 ( .A(n9186), .B(n46866), .Z(n59445) );
  XNOR U12352 ( .A(x[6710]), .B(y[6710]), .Z(n22925) );
  ANDN U12353 ( .B(y[6709]), .A(x[6709]), .Z(n59443) );
  ANDN U12354 ( .B(n22925), .A(n59443), .Z(n19572) );
  XNOR U12355 ( .A(x[6708]), .B(y[6708]), .Z(n46857) );
  NANDN U12356 ( .A(y[6706]), .B(x[6706]), .Z(n9187) );
  NANDN U12357 ( .A(y[6707]), .B(x[6707]), .Z(n46856) );
  AND U12358 ( .A(n9187), .B(n46856), .Z(n59440) );
  XNOR U12359 ( .A(x[6706]), .B(y[6706]), .Z(n22927) );
  ANDN U12360 ( .B(y[6705]), .A(x[6705]), .Z(n59438) );
  ANDN U12361 ( .B(n22927), .A(n59438), .Z(n19565) );
  XNOR U12362 ( .A(x[6704]), .B(y[6704]), .Z(n46847) );
  NANDN U12363 ( .A(y[6702]), .B(x[6702]), .Z(n9188) );
  NANDN U12364 ( .A(y[6703]), .B(x[6703]), .Z(n46846) );
  AND U12365 ( .A(n9188), .B(n46846), .Z(n59434) );
  ANDN U12366 ( .B(y[6701]), .A(x[6701]), .Z(n59432) );
  XNOR U12367 ( .A(x[6702]), .B(y[6702]), .Z(n22929) );
  NANDN U12368 ( .A(y[6700]), .B(x[6700]), .Z(n9189) );
  NANDN U12369 ( .A(y[6701]), .B(x[6701]), .Z(n22928) );
  AND U12370 ( .A(n9189), .B(n22928), .Z(n59431) );
  XNOR U12371 ( .A(x[6698]), .B(y[6698]), .Z(n22931) );
  NANDN U12372 ( .A(x[6697]), .B(y[6697]), .Z(n59428) );
  AND U12373 ( .A(n22931), .B(n59428), .Z(n19551) );
  XNOR U12374 ( .A(x[6696]), .B(y[6696]), .Z(n46827) );
  NANDN U12375 ( .A(x[6695]), .B(y[6695]), .Z(n59423) );
  AND U12376 ( .A(n46827), .B(n59423), .Z(n19547) );
  XNOR U12377 ( .A(x[6694]), .B(y[6694]), .Z(n22933) );
  NANDN U12378 ( .A(y[6692]), .B(x[6692]), .Z(n9190) );
  NANDN U12379 ( .A(y[6693]), .B(x[6693]), .Z(n22932) );
  AND U12380 ( .A(n9190), .B(n22932), .Z(n59421) );
  NANDN U12381 ( .A(x[6691]), .B(y[6691]), .Z(n59419) );
  XNOR U12382 ( .A(x[6692]), .B(y[6692]), .Z(n46817) );
  AND U12383 ( .A(n59419), .B(n46817), .Z(n19540) );
  XNOR U12384 ( .A(x[6690]), .B(y[6690]), .Z(n22935) );
  NANDN U12385 ( .A(y[6688]), .B(x[6688]), .Z(n9191) );
  NANDN U12386 ( .A(y[6689]), .B(x[6689]), .Z(n22934) );
  AND U12387 ( .A(n9191), .B(n22934), .Z(n59417) );
  XNOR U12388 ( .A(x[6688]), .B(y[6688]), .Z(n22937) );
  NANDN U12389 ( .A(y[6686]), .B(x[6686]), .Z(n9192) );
  NANDN U12390 ( .A(y[6687]), .B(x[6687]), .Z(n22936) );
  NAND U12391 ( .A(n9192), .B(n22936), .Z(n59416) );
  XNOR U12392 ( .A(x[6686]), .B(y[6686]), .Z(n22939) );
  ANDN U12393 ( .B(y[6685]), .A(x[6685]), .Z(n59414) );
  ANDN U12394 ( .B(n22939), .A(n59414), .Z(n19530) );
  NANDN U12395 ( .A(y[6684]), .B(x[6684]), .Z(n9193) );
  NANDN U12396 ( .A(y[6685]), .B(x[6685]), .Z(n22938) );
  NAND U12397 ( .A(n9193), .B(n22938), .Z(n59413) );
  XNOR U12398 ( .A(x[6684]), .B(y[6684]), .Z(n46799) );
  NANDN U12399 ( .A(y[6682]), .B(x[6682]), .Z(n9194) );
  NANDN U12400 ( .A(y[6683]), .B(x[6683]), .Z(n46798) );
  NAND U12401 ( .A(n9194), .B(n46798), .Z(n59410) );
  XNOR U12402 ( .A(x[6682]), .B(y[6682]), .Z(n22941) );
  NANDN U12403 ( .A(x[6681]), .B(y[6681]), .Z(n59408) );
  AND U12404 ( .A(n22941), .B(n59408), .Z(n19524) );
  XNOR U12405 ( .A(x[6680]), .B(y[6680]), .Z(n22943) );
  NANDN U12406 ( .A(y[6678]), .B(x[6678]), .Z(n9195) );
  NANDN U12407 ( .A(y[6679]), .B(x[6679]), .Z(n22942) );
  AND U12408 ( .A(n9195), .B(n22942), .Z(n59406) );
  XNOR U12409 ( .A(x[6678]), .B(y[6678]), .Z(n22945) );
  NANDN U12410 ( .A(x[6677]), .B(y[6677]), .Z(n59404) );
  AND U12411 ( .A(n22945), .B(n59404), .Z(n19517) );
  XNOR U12412 ( .A(x[6676]), .B(y[6676]), .Z(n22947) );
  NANDN U12413 ( .A(y[6674]), .B(x[6674]), .Z(n22949) );
  NANDN U12414 ( .A(y[6675]), .B(x[6675]), .Z(n22946) );
  AND U12415 ( .A(n22949), .B(n22946), .Z(n59400) );
  NANDN U12416 ( .A(x[6673]), .B(y[6673]), .Z(n22951) );
  NANDN U12417 ( .A(x[6674]), .B(y[6674]), .Z(n22948) );
  AND U12418 ( .A(n22951), .B(n22948), .Z(n59399) );
  NANDN U12419 ( .A(x[6671]), .B(y[6671]), .Z(n22955) );
  NANDN U12420 ( .A(x[6672]), .B(y[6672]), .Z(n22952) );
  AND U12421 ( .A(n22955), .B(n22952), .Z(n59397) );
  NANDN U12422 ( .A(y[6670]), .B(x[6670]), .Z(n9196) );
  NANDN U12423 ( .A(y[6671]), .B(x[6671]), .Z(n22954) );
  AND U12424 ( .A(n9196), .B(n22954), .Z(n59396) );
  ANDN U12425 ( .B(y[6669]), .A(x[6669]), .Z(n50995) );
  XNOR U12426 ( .A(x[6670]), .B(y[6670]), .Z(n22957) );
  NANDN U12427 ( .A(y[6668]), .B(x[6668]), .Z(n9197) );
  NANDN U12428 ( .A(y[6669]), .B(x[6669]), .Z(n22956) );
  NAND U12429 ( .A(n9197), .B(n22956), .Z(n59394) );
  ANDN U12430 ( .B(y[6665]), .A(x[6665]), .Z(n59391) );
  XNOR U12431 ( .A(x[6666]), .B(y[6666]), .Z(n22959) );
  NANDN U12432 ( .A(y[6664]), .B(x[6664]), .Z(n9198) );
  NANDN U12433 ( .A(y[6665]), .B(x[6665]), .Z(n22958) );
  AND U12434 ( .A(n9198), .B(n22958), .Z(n50999) );
  XNOR U12435 ( .A(x[6664]), .B(y[6664]), .Z(n46755) );
  ANDN U12436 ( .B(y[6663]), .A(x[6663]), .Z(n46751) );
  ANDN U12437 ( .B(n46755), .A(n46751), .Z(n19496) );
  XNOR U12438 ( .A(x[6662]), .B(y[6662]), .Z(n22961) );
  NANDN U12439 ( .A(y[6660]), .B(x[6660]), .Z(n9199) );
  NANDN U12440 ( .A(y[6661]), .B(x[6661]), .Z(n22960) );
  AND U12441 ( .A(n9199), .B(n22960), .Z(n59387) );
  XNOR U12442 ( .A(x[6660]), .B(y[6660]), .Z(n46744) );
  NANDN U12443 ( .A(x[6659]), .B(y[6659]), .Z(n51002) );
  AND U12444 ( .A(n46744), .B(n51002), .Z(n19489) );
  XNOR U12445 ( .A(x[6658]), .B(y[6658]), .Z(n22963) );
  NANDN U12446 ( .A(y[6656]), .B(x[6656]), .Z(n9200) );
  NANDN U12447 ( .A(y[6657]), .B(x[6657]), .Z(n22962) );
  AND U12448 ( .A(n9200), .B(n22962), .Z(n59381) );
  NANDN U12449 ( .A(x[6655]), .B(y[6655]), .Z(n59379) );
  XNOR U12450 ( .A(x[6656]), .B(y[6656]), .Z(n46734) );
  AND U12451 ( .A(n59379), .B(n46734), .Z(n19482) );
  NANDN U12452 ( .A(y[6654]), .B(x[6654]), .Z(n22965) );
  NANDN U12453 ( .A(y[6655]), .B(x[6655]), .Z(n46733) );
  NAND U12454 ( .A(n22965), .B(n46733), .Z(n59378) );
  NANDN U12455 ( .A(x[6653]), .B(y[6653]), .Z(n22967) );
  NANDN U12456 ( .A(x[6654]), .B(y[6654]), .Z(n22964) );
  AND U12457 ( .A(n22967), .B(n22964), .Z(n59377) );
  NANDN U12458 ( .A(y[6652]), .B(x[6652]), .Z(n22969) );
  NANDN U12459 ( .A(y[6653]), .B(x[6653]), .Z(n22966) );
  AND U12460 ( .A(n22969), .B(n22966), .Z(n59376) );
  NANDN U12461 ( .A(x[6651]), .B(y[6651]), .Z(n22971) );
  NANDN U12462 ( .A(x[6652]), .B(y[6652]), .Z(n22968) );
  AND U12463 ( .A(n22971), .B(n22968), .Z(n59375) );
  NANDN U12464 ( .A(y[6650]), .B(x[6650]), .Z(n9201) );
  NANDN U12465 ( .A(y[6651]), .B(x[6651]), .Z(n22970) );
  AND U12466 ( .A(n9201), .B(n22970), .Z(n59374) );
  XNOR U12467 ( .A(y[6650]), .B(x[6650]), .Z(n22974) );
  ANDN U12468 ( .B(y[6649]), .A(x[6649]), .Z(n22975) );
  ANDN U12469 ( .B(n22974), .A(n22975), .Z(n59373) );
  XNOR U12470 ( .A(x[6648]), .B(y[6648]), .Z(n46716) );
  NANDN U12471 ( .A(y[6646]), .B(x[6646]), .Z(n9202) );
  NANDN U12472 ( .A(y[6647]), .B(x[6647]), .Z(n46715) );
  AND U12473 ( .A(n9202), .B(n46715), .Z(n59372) );
  XNOR U12474 ( .A(x[6646]), .B(y[6646]), .Z(n22977) );
  ANDN U12475 ( .B(y[6645]), .A(x[6645]), .Z(n59370) );
  ANDN U12476 ( .B(n22977), .A(n59370), .Z(n19469) );
  XNOR U12477 ( .A(x[6644]), .B(y[6644]), .Z(n46706) );
  NANDN U12478 ( .A(y[6642]), .B(x[6642]), .Z(n9203) );
  NANDN U12479 ( .A(y[6643]), .B(x[6643]), .Z(n46705) );
  AND U12480 ( .A(n9203), .B(n46705), .Z(n59367) );
  XNOR U12481 ( .A(x[6642]), .B(y[6642]), .Z(n22979) );
  ANDN U12482 ( .B(y[6641]), .A(x[6641]), .Z(n59365) );
  ANDN U12483 ( .B(n22979), .A(n59365), .Z(n19462) );
  XNOR U12484 ( .A(x[6640]), .B(y[6640]), .Z(n46696) );
  NANDN U12485 ( .A(y[6638]), .B(x[6638]), .Z(n9204) );
  NANDN U12486 ( .A(y[6639]), .B(x[6639]), .Z(n46695) );
  AND U12487 ( .A(n9204), .B(n46695), .Z(n59363) );
  ANDN U12488 ( .B(y[6637]), .A(x[6637]), .Z(n59361) );
  XNOR U12489 ( .A(x[6638]), .B(y[6638]), .Z(n22981) );
  NANDN U12490 ( .A(y[6636]), .B(x[6636]), .Z(n9205) );
  NANDN U12491 ( .A(y[6637]), .B(x[6637]), .Z(n22980) );
  AND U12492 ( .A(n9205), .B(n22980), .Z(n59360) );
  XNOR U12493 ( .A(x[6636]), .B(y[6636]), .Z(n22983) );
  NANDN U12494 ( .A(y[6634]), .B(x[6634]), .Z(n9206) );
  NANDN U12495 ( .A(y[6635]), .B(x[6635]), .Z(n22982) );
  AND U12496 ( .A(n9206), .B(n22982), .Z(n59357) );
  XNOR U12497 ( .A(y[6634]), .B(x[6634]), .Z(n22985) );
  NANDN U12498 ( .A(x[6633]), .B(y[6633]), .Z(n22986) );
  AND U12499 ( .A(n22985), .B(n22986), .Z(n59356) );
  NANDN U12500 ( .A(y[6632]), .B(x[6632]), .Z(n22988) );
  NANDN U12501 ( .A(y[6633]), .B(x[6633]), .Z(n22984) );
  NAND U12502 ( .A(n22988), .B(n22984), .Z(n59355) );
  NANDN U12503 ( .A(x[6631]), .B(y[6631]), .Z(n22990) );
  NANDN U12504 ( .A(x[6632]), .B(y[6632]), .Z(n22987) );
  AND U12505 ( .A(n22990), .B(n22987), .Z(n59353) );
  XNOR U12506 ( .A(x[6630]), .B(y[6630]), .Z(n22992) );
  NANDN U12507 ( .A(x[6627]), .B(y[6627]), .Z(n46667) );
  NANDN U12508 ( .A(x[6628]), .B(y[6628]), .Z(n22993) );
  AND U12509 ( .A(n46667), .B(n22993), .Z(n59350) );
  NANDN U12510 ( .A(y[6626]), .B(x[6626]), .Z(n9207) );
  NANDN U12511 ( .A(y[6627]), .B(x[6627]), .Z(n22995) );
  AND U12512 ( .A(n9207), .B(n22995), .Z(n59349) );
  XNOR U12513 ( .A(x[6626]), .B(y[6626]), .Z(n22997) );
  ANDN U12514 ( .B(y[6625]), .A(x[6625]), .Z(n22998) );
  NANDN U12515 ( .A(x[6623]), .B(y[6623]), .Z(n23002) );
  NANDN U12516 ( .A(x[6624]), .B(y[6624]), .Z(n22999) );
  AND U12517 ( .A(n23002), .B(n22999), .Z(n59345) );
  NANDN U12518 ( .A(y[6622]), .B(x[6622]), .Z(n23004) );
  NANDN U12519 ( .A(y[6623]), .B(x[6623]), .Z(n23001) );
  AND U12520 ( .A(n23004), .B(n23001), .Z(n59344) );
  NANDN U12521 ( .A(x[6621]), .B(y[6621]), .Z(n23006) );
  NANDN U12522 ( .A(x[6622]), .B(y[6622]), .Z(n23003) );
  NAND U12523 ( .A(n23006), .B(n23003), .Z(n51014) );
  NANDN U12524 ( .A(y[6620]), .B(x[6620]), .Z(n9208) );
  NANDN U12525 ( .A(y[6621]), .B(x[6621]), .Z(n23005) );
  AND U12526 ( .A(n9208), .B(n23005), .Z(n59343) );
  XNOR U12527 ( .A(x[6620]), .B(y[6620]), .Z(n23008) );
  NANDN U12528 ( .A(y[6618]), .B(x[6618]), .Z(n9209) );
  NANDN U12529 ( .A(y[6619]), .B(x[6619]), .Z(n23007) );
  AND U12530 ( .A(n9209), .B(n23007), .Z(n59340) );
  ANDN U12531 ( .B(y[6617]), .A(x[6617]), .Z(n59337) );
  XNOR U12532 ( .A(x[6618]), .B(y[6618]), .Z(n23011) );
  NANDN U12533 ( .A(y[6616]), .B(x[6616]), .Z(n9210) );
  NANDN U12534 ( .A(y[6617]), .B(x[6617]), .Z(n23010) );
  AND U12535 ( .A(n9210), .B(n23010), .Z(n59336) );
  ANDN U12536 ( .B(y[6613]), .A(x[6613]), .Z(n51016) );
  XNOR U12537 ( .A(x[6614]), .B(y[6614]), .Z(n23013) );
  NANDN U12538 ( .A(y[6612]), .B(x[6612]), .Z(n9211) );
  NANDN U12539 ( .A(y[6613]), .B(x[6613]), .Z(n23012) );
  AND U12540 ( .A(n9211), .B(n23012), .Z(n59333) );
  XNOR U12541 ( .A(x[6612]), .B(y[6612]), .Z(n46634) );
  NANDN U12542 ( .A(x[6611]), .B(y[6611]), .Z(n59331) );
  NAND U12543 ( .A(n46634), .B(n59331), .Z(n19419) );
  NANDN U12544 ( .A(y[6610]), .B(x[6610]), .Z(n9212) );
  NANDN U12545 ( .A(y[6611]), .B(x[6611]), .Z(n46633) );
  AND U12546 ( .A(n9212), .B(n46633), .Z(n59330) );
  NANDN U12547 ( .A(x[6609]), .B(y[6609]), .Z(n23016) );
  XNOR U12548 ( .A(x[6610]), .B(y[6610]), .Z(n23015) );
  NAND U12549 ( .A(n23016), .B(n23015), .Z(n19416) );
  NANDN U12550 ( .A(y[6608]), .B(x[6608]), .Z(n9213) );
  NANDN U12551 ( .A(y[6609]), .B(x[6609]), .Z(n23014) );
  AND U12552 ( .A(n9213), .B(n23014), .Z(n59329) );
  ANDN U12553 ( .B(y[6607]), .A(x[6607]), .Z(n23017) );
  XOR U12554 ( .A(x[6608]), .B(y[6608]), .Z(n46624) );
  NOR U12555 ( .A(n23017), .B(n46624), .Z(n19413) );
  XNOR U12556 ( .A(x[6606]), .B(y[6606]), .Z(n23019) );
  NANDN U12557 ( .A(y[6604]), .B(x[6604]), .Z(n9214) );
  NANDN U12558 ( .A(y[6605]), .B(x[6605]), .Z(n23018) );
  AND U12559 ( .A(n9214), .B(n23018), .Z(n59322) );
  XNOR U12560 ( .A(x[6604]), .B(y[6604]), .Z(n23021) );
  NANDN U12561 ( .A(y[6602]), .B(x[6602]), .Z(n9215) );
  NANDN U12562 ( .A(y[6603]), .B(x[6603]), .Z(n23020) );
  NAND U12563 ( .A(n9215), .B(n23020), .Z(n59319) );
  NANDN U12564 ( .A(y[6600]), .B(x[6600]), .Z(n9216) );
  NANDN U12565 ( .A(y[6601]), .B(x[6601]), .Z(n23022) );
  AND U12566 ( .A(n9216), .B(n23022), .Z(n59316) );
  XNOR U12567 ( .A(x[6600]), .B(y[6600]), .Z(n23025) );
  NANDN U12568 ( .A(y[6598]), .B(x[6598]), .Z(n9217) );
  NANDN U12569 ( .A(y[6599]), .B(x[6599]), .Z(n23024) );
  NAND U12570 ( .A(n9217), .B(n23024), .Z(n59315) );
  XNOR U12571 ( .A(x[6598]), .B(y[6598]), .Z(n23027) );
  NANDN U12572 ( .A(x[6597]), .B(y[6597]), .Z(n59313) );
  AND U12573 ( .A(n23027), .B(n59313), .Z(n19397) );
  NANDN U12574 ( .A(y[6596]), .B(x[6596]), .Z(n9218) );
  NANDN U12575 ( .A(y[6597]), .B(x[6597]), .Z(n23026) );
  NAND U12576 ( .A(n9218), .B(n23026), .Z(n59312) );
  XNOR U12577 ( .A(x[6596]), .B(y[6596]), .Z(n23029) );
  NANDN U12578 ( .A(y[6594]), .B(x[6594]), .Z(n9219) );
  NANDN U12579 ( .A(y[6595]), .B(x[6595]), .Z(n23028) );
  AND U12580 ( .A(n9219), .B(n23028), .Z(n59309) );
  NANDN U12581 ( .A(x[6593]), .B(y[6593]), .Z(n59307) );
  XNOR U12582 ( .A(x[6594]), .B(y[6594]), .Z(n23031) );
  NAND U12583 ( .A(n59307), .B(n23031), .Z(n19391) );
  NANDN U12584 ( .A(y[6592]), .B(x[6592]), .Z(n9220) );
  NANDN U12585 ( .A(y[6593]), .B(x[6593]), .Z(n23030) );
  AND U12586 ( .A(n9220), .B(n23030), .Z(n59305) );
  XNOR U12587 ( .A(x[6592]), .B(y[6592]), .Z(n23033) );
  NANDN U12588 ( .A(x[6591]), .B(y[6591]), .Z(n51022) );
  NAND U12589 ( .A(n23033), .B(n51022), .Z(n19388) );
  XNOR U12590 ( .A(x[6590]), .B(y[6590]), .Z(n23035) );
  NANDN U12591 ( .A(y[6588]), .B(x[6588]), .Z(n9221) );
  NANDN U12592 ( .A(y[6589]), .B(x[6589]), .Z(n23034) );
  NAND U12593 ( .A(n9221), .B(n23034), .Z(n59301) );
  XNOR U12594 ( .A(x[6586]), .B(y[6586]), .Z(n23039) );
  NANDN U12595 ( .A(y[6584]), .B(x[6584]), .Z(n9222) );
  NANDN U12596 ( .A(y[6585]), .B(x[6585]), .Z(n23038) );
  NAND U12597 ( .A(n9222), .B(n23038), .Z(n59296) );
  NANDN U12598 ( .A(x[6583]), .B(y[6583]), .Z(n51025) );
  XOR U12599 ( .A(x[6584]), .B(y[6584]), .Z(n46575) );
  ANDN U12600 ( .B(n51025), .A(n46575), .Z(n19374) );
  ANDN U12601 ( .B(x[6583]), .A(y[6583]), .Z(n46574) );
  NANDN U12602 ( .A(y[6582]), .B(x[6582]), .Z(n9223) );
  NANDN U12603 ( .A(n46574), .B(n9223), .Z(n59293) );
  XNOR U12604 ( .A(x[6582]), .B(y[6582]), .Z(n23041) );
  NANDN U12605 ( .A(y[6580]), .B(x[6580]), .Z(n9224) );
  NANDN U12606 ( .A(y[6581]), .B(x[6581]), .Z(n23040) );
  AND U12607 ( .A(n9224), .B(n23040), .Z(n59290) );
  XNOR U12608 ( .A(x[6580]), .B(y[6580]), .Z(n23043) );
  NANDN U12609 ( .A(x[6579]), .B(y[6579]), .Z(n59288) );
  AND U12610 ( .A(n23043), .B(n59288), .Z(n19368) );
  XNOR U12611 ( .A(x[6578]), .B(y[6578]), .Z(n23045) );
  NANDN U12612 ( .A(y[6576]), .B(x[6576]), .Z(n9225) );
  NANDN U12613 ( .A(y[6577]), .B(x[6577]), .Z(n23044) );
  AND U12614 ( .A(n9225), .B(n23044), .Z(n59284) );
  ANDN U12615 ( .B(y[6575]), .A(x[6575]), .Z(n46552) );
  XOR U12616 ( .A(x[6576]), .B(y[6576]), .Z(n9226) );
  NOR U12617 ( .A(n46552), .B(n9226), .Z(n19361) );
  XNOR U12618 ( .A(x[6574]), .B(y[6574]), .Z(n46549) );
  NANDN U12619 ( .A(y[6572]), .B(x[6572]), .Z(n9227) );
  NANDN U12620 ( .A(y[6573]), .B(x[6573]), .Z(n46548) );
  AND U12621 ( .A(n9227), .B(n46548), .Z(n59280) );
  XNOR U12622 ( .A(x[6572]), .B(y[6572]), .Z(n23047) );
  NANDN U12623 ( .A(y[6570]), .B(x[6570]), .Z(n9228) );
  NANDN U12624 ( .A(y[6571]), .B(x[6571]), .Z(n23046) );
  NAND U12625 ( .A(n9228), .B(n23046), .Z(n59276) );
  NANDN U12626 ( .A(y[6568]), .B(x[6568]), .Z(n9229) );
  NANDN U12627 ( .A(y[6569]), .B(x[6569]), .Z(n23048) );
  AND U12628 ( .A(n9229), .B(n23048), .Z(n59273) );
  NANDN U12629 ( .A(x[6567]), .B(y[6567]), .Z(n23052) );
  IV U12630 ( .A(n23052), .Z(n51029) );
  XNOR U12631 ( .A(x[6568]), .B(y[6568]), .Z(n23051) );
  NANDN U12632 ( .A(y[6566]), .B(x[6566]), .Z(n9230) );
  NANDN U12633 ( .A(y[6567]), .B(x[6567]), .Z(n23050) );
  NAND U12634 ( .A(n9230), .B(n23050), .Z(n59272) );
  XNOR U12635 ( .A(x[6566]), .B(y[6566]), .Z(n23054) );
  ANDN U12636 ( .B(y[6565]), .A(x[6565]), .Z(n23055) );
  NANDN U12637 ( .A(x[6563]), .B(y[6563]), .Z(n46524) );
  NANDN U12638 ( .A(x[6564]), .B(y[6564]), .Z(n23056) );
  AND U12639 ( .A(n46524), .B(n23056), .Z(n59269) );
  NANDN U12640 ( .A(y[6562]), .B(x[6562]), .Z(n23059) );
  NANDN U12641 ( .A(y[6563]), .B(x[6563]), .Z(n23058) );
  AND U12642 ( .A(n23059), .B(n23058), .Z(n59268) );
  NANDN U12643 ( .A(x[6561]), .B(y[6561]), .Z(n46520) );
  NANDN U12644 ( .A(x[6562]), .B(y[6562]), .Z(n46525) );
  AND U12645 ( .A(n46520), .B(n46525), .Z(n59267) );
  NANDN U12646 ( .A(y[6560]), .B(x[6560]), .Z(n9231) );
  NANDN U12647 ( .A(y[6561]), .B(x[6561]), .Z(n23060) );
  NAND U12648 ( .A(n9231), .B(n23060), .Z(n59266) );
  XNOR U12649 ( .A(x[6560]), .B(y[6560]), .Z(n23062) );
  NANDN U12650 ( .A(x[6559]), .B(y[6559]), .Z(n59264) );
  AND U12651 ( .A(n23062), .B(n59264), .Z(n19338) );
  NANDN U12652 ( .A(y[6558]), .B(x[6558]), .Z(n9232) );
  NANDN U12653 ( .A(y[6559]), .B(x[6559]), .Z(n23061) );
  NAND U12654 ( .A(n9232), .B(n23061), .Z(n59262) );
  XNOR U12655 ( .A(x[6558]), .B(y[6558]), .Z(n23064) );
  NANDN U12656 ( .A(y[6556]), .B(x[6556]), .Z(n9233) );
  NANDN U12657 ( .A(y[6557]), .B(x[6557]), .Z(n23063) );
  NAND U12658 ( .A(n9233), .B(n23063), .Z(n59259) );
  NANDN U12659 ( .A(x[6555]), .B(y[6555]), .Z(n51032) );
  XOR U12660 ( .A(x[6556]), .B(y[6556]), .Z(n46508) );
  ANDN U12661 ( .B(n51032), .A(n46508), .Z(n19332) );
  ANDN U12662 ( .B(x[6555]), .A(y[6555]), .Z(n46510) );
  NANDN U12663 ( .A(y[6554]), .B(x[6554]), .Z(n9234) );
  NANDN U12664 ( .A(n46510), .B(n9234), .Z(n59258) );
  XNOR U12665 ( .A(x[6554]), .B(y[6554]), .Z(n23066) );
  NANDN U12666 ( .A(y[6552]), .B(x[6552]), .Z(n9235) );
  NANDN U12667 ( .A(y[6553]), .B(x[6553]), .Z(n23065) );
  AND U12668 ( .A(n9235), .B(n23065), .Z(n59255) );
  XNOR U12669 ( .A(x[6552]), .B(y[6552]), .Z(n23068) );
  NANDN U12670 ( .A(x[6551]), .B(y[6551]), .Z(n59253) );
  AND U12671 ( .A(n23068), .B(n59253), .Z(n19326) );
  XNOR U12672 ( .A(x[6550]), .B(y[6550]), .Z(n23070) );
  NANDN U12673 ( .A(y[6548]), .B(x[6548]), .Z(n9236) );
  NANDN U12674 ( .A(y[6549]), .B(x[6549]), .Z(n23069) );
  AND U12675 ( .A(n9236), .B(n23069), .Z(n59249) );
  XNOR U12676 ( .A(y[6548]), .B(x[6548]), .Z(n23072) );
  NANDN U12677 ( .A(x[6547]), .B(y[6547]), .Z(n46488) );
  NAND U12678 ( .A(n23072), .B(n46488), .Z(n59248) );
  NANDN U12679 ( .A(y[6546]), .B(x[6546]), .Z(n9237) );
  NANDN U12680 ( .A(y[6547]), .B(x[6547]), .Z(n23071) );
  AND U12681 ( .A(n9237), .B(n23071), .Z(n59246) );
  XNOR U12682 ( .A(x[6546]), .B(y[6546]), .Z(n23074) );
  NANDN U12683 ( .A(x[6545]), .B(y[6545]), .Z(n59245) );
  NAND U12684 ( .A(n23074), .B(n59245), .Z(n19317) );
  NANDN U12685 ( .A(x[6543]), .B(y[6543]), .Z(n46479) );
  IV U12686 ( .A(n46479), .Z(n59243) );
  XNOR U12687 ( .A(x[6544]), .B(y[6544]), .Z(n23076) );
  NANDN U12688 ( .A(y[6542]), .B(x[6542]), .Z(n9238) );
  NANDN U12689 ( .A(y[6543]), .B(x[6543]), .Z(n23075) );
  NAND U12690 ( .A(n9238), .B(n23075), .Z(n59242) );
  XNOR U12691 ( .A(x[6542]), .B(y[6542]), .Z(n23078) );
  NANDN U12692 ( .A(x[6541]), .B(y[6541]), .Z(n51036) );
  AND U12693 ( .A(n23078), .B(n51036), .Z(n19310) );
  NANDN U12694 ( .A(y[6540]), .B(x[6540]), .Z(n9239) );
  NANDN U12695 ( .A(y[6541]), .B(x[6541]), .Z(n23077) );
  NAND U12696 ( .A(n9239), .B(n23077), .Z(n59241) );
  XNOR U12697 ( .A(x[6540]), .B(y[6540]), .Z(n23080) );
  NANDN U12698 ( .A(y[6538]), .B(x[6538]), .Z(n9240) );
  NANDN U12699 ( .A(y[6539]), .B(x[6539]), .Z(n23079) );
  AND U12700 ( .A(n9240), .B(n23079), .Z(n59238) );
  XNOR U12701 ( .A(x[6538]), .B(y[6538]), .Z(n23082) );
  NANDN U12702 ( .A(x[6537]), .B(y[6537]), .Z(n59236) );
  NAND U12703 ( .A(n23082), .B(n59236), .Z(n19304) );
  NANDN U12704 ( .A(y[6536]), .B(x[6536]), .Z(n9241) );
  NANDN U12705 ( .A(y[6537]), .B(x[6537]), .Z(n23081) );
  AND U12706 ( .A(n9241), .B(n23081), .Z(n51038) );
  XNOR U12707 ( .A(x[6536]), .B(y[6536]), .Z(n23084) );
  NANDN U12708 ( .A(x[6535]), .B(y[6535]), .Z(n59234) );
  NAND U12709 ( .A(n23084), .B(n59234), .Z(n19301) );
  NANDN U12710 ( .A(y[6534]), .B(x[6534]), .Z(n9242) );
  NANDN U12711 ( .A(y[6535]), .B(x[6535]), .Z(n23083) );
  AND U12712 ( .A(n9242), .B(n23083), .Z(n59232) );
  XNOR U12713 ( .A(x[6534]), .B(y[6534]), .Z(n23086) );
  NANDN U12714 ( .A(y[6532]), .B(x[6532]), .Z(n9243) );
  NANDN U12715 ( .A(y[6533]), .B(x[6533]), .Z(n23085) );
  NAND U12716 ( .A(n9243), .B(n23085), .Z(n59231) );
  XNOR U12717 ( .A(y[6532]), .B(x[6532]), .Z(n23087) );
  NANDN U12718 ( .A(x[6531]), .B(y[6531]), .Z(n23089) );
  AND U12719 ( .A(n23087), .B(n23089), .Z(n59230) );
  NANDN U12720 ( .A(y[6530]), .B(x[6530]), .Z(n23091) );
  NANDN U12721 ( .A(y[6531]), .B(x[6531]), .Z(n23088) );
  NAND U12722 ( .A(n23091), .B(n23088), .Z(n59229) );
  NANDN U12723 ( .A(x[6529]), .B(y[6529]), .Z(n46449) );
  NANDN U12724 ( .A(x[6530]), .B(y[6530]), .Z(n23090) );
  AND U12725 ( .A(n46449), .B(n23090), .Z(n59228) );
  NANDN U12726 ( .A(y[6528]), .B(x[6528]), .Z(n9244) );
  NANDN U12727 ( .A(y[6529]), .B(x[6529]), .Z(n23092) );
  AND U12728 ( .A(n9244), .B(n23092), .Z(n59227) );
  XNOR U12729 ( .A(x[6528]), .B(y[6528]), .Z(n23094) );
  NANDN U12730 ( .A(x[6527]), .B(y[6527]), .Z(n51041) );
  NAND U12731 ( .A(n23094), .B(n51041), .Z(n19291) );
  NANDN U12732 ( .A(y[6526]), .B(x[6526]), .Z(n9245) );
  NANDN U12733 ( .A(y[6527]), .B(x[6527]), .Z(n23093) );
  AND U12734 ( .A(n9245), .B(n23093), .Z(n59226) );
  NANDN U12735 ( .A(x[6525]), .B(y[6525]), .Z(n59224) );
  XNOR U12736 ( .A(x[6526]), .B(y[6526]), .Z(n23096) );
  NAND U12737 ( .A(n59224), .B(n23096), .Z(n19288) );
  NANDN U12738 ( .A(y[6524]), .B(x[6524]), .Z(n9246) );
  NANDN U12739 ( .A(y[6525]), .B(x[6525]), .Z(n23095) );
  AND U12740 ( .A(n9246), .B(n23095), .Z(n59223) );
  XNOR U12741 ( .A(x[6524]), .B(y[6524]), .Z(n23098) );
  NANDN U12742 ( .A(y[6522]), .B(x[6522]), .Z(n9247) );
  NANDN U12743 ( .A(y[6523]), .B(x[6523]), .Z(n23097) );
  NAND U12744 ( .A(n9247), .B(n23097), .Z(n59219) );
  NANDN U12745 ( .A(y[6520]), .B(x[6520]), .Z(n9248) );
  NANDN U12746 ( .A(y[6521]), .B(x[6521]), .Z(n23099) );
  AND U12747 ( .A(n9248), .B(n23099), .Z(n59216) );
  XNOR U12748 ( .A(x[6520]), .B(y[6520]), .Z(n23102) );
  NANDN U12749 ( .A(y[6518]), .B(x[6518]), .Z(n9249) );
  NANDN U12750 ( .A(y[6519]), .B(x[6519]), .Z(n23101) );
  NAND U12751 ( .A(n9249), .B(n23101), .Z(n59215) );
  NANDN U12752 ( .A(x[6517]), .B(y[6517]), .Z(n59213) );
  XNOR U12753 ( .A(x[6518]), .B(y[6518]), .Z(n23104) );
  NANDN U12754 ( .A(y[6516]), .B(x[6516]), .Z(n9250) );
  NANDN U12755 ( .A(y[6517]), .B(x[6517]), .Z(n23103) );
  AND U12756 ( .A(n9250), .B(n23103), .Z(n59212) );
  XNOR U12757 ( .A(x[6516]), .B(y[6516]), .Z(n23106) );
  XNOR U12758 ( .A(x[6514]), .B(y[6514]), .Z(n23108) );
  NANDN U12759 ( .A(x[6513]), .B(y[6513]), .Z(n59209) );
  AND U12760 ( .A(n23108), .B(n59209), .Z(n19269) );
  XNOR U12761 ( .A(x[6512]), .B(y[6512]), .Z(n23110) );
  NANDN U12762 ( .A(y[6510]), .B(x[6510]), .Z(n9251) );
  NANDN U12763 ( .A(y[6511]), .B(x[6511]), .Z(n23109) );
  AND U12764 ( .A(n9251), .B(n23109), .Z(n59203) );
  XNOR U12765 ( .A(x[6510]), .B(y[6510]), .Z(n23112) );
  ANDN U12766 ( .B(y[6509]), .A(x[6509]), .Z(n46407) );
  ANDN U12767 ( .B(n23112), .A(n46407), .Z(n19262) );
  XNOR U12768 ( .A(x[6508]), .B(y[6508]), .Z(n23114) );
  NANDN U12769 ( .A(y[6506]), .B(x[6506]), .Z(n9252) );
  NANDN U12770 ( .A(y[6507]), .B(x[6507]), .Z(n23113) );
  AND U12771 ( .A(n9252), .B(n23113), .Z(n59197) );
  NANDN U12772 ( .A(x[6505]), .B(y[6505]), .Z(n59196) );
  XNOR U12773 ( .A(x[6506]), .B(y[6506]), .Z(n23116) );
  NANDN U12774 ( .A(y[6504]), .B(x[6504]), .Z(n9253) );
  NANDN U12775 ( .A(y[6505]), .B(x[6505]), .Z(n23115) );
  NAND U12776 ( .A(n9253), .B(n23115), .Z(n59194) );
  NANDN U12777 ( .A(y[6502]), .B(x[6502]), .Z(n9254) );
  ANDN U12778 ( .B(x[6503]), .A(y[6503]), .Z(n46398) );
  ANDN U12779 ( .B(n9254), .A(n46398), .Z(n59193) );
  XNOR U12780 ( .A(x[6502]), .B(y[6502]), .Z(n23118) );
  NANDN U12781 ( .A(y[6500]), .B(x[6500]), .Z(n9255) );
  NANDN U12782 ( .A(y[6501]), .B(x[6501]), .Z(n23117) );
  NAND U12783 ( .A(n9255), .B(n23117), .Z(n59190) );
  NANDN U12784 ( .A(x[6499]), .B(y[6499]), .Z(n59187) );
  XNOR U12785 ( .A(x[6500]), .B(y[6500]), .Z(n23120) );
  NANDN U12786 ( .A(y[6498]), .B(x[6498]), .Z(n9256) );
  NANDN U12787 ( .A(y[6499]), .B(x[6499]), .Z(n23119) );
  AND U12788 ( .A(n9256), .B(n23119), .Z(n59186) );
  NANDN U12789 ( .A(y[6496]), .B(x[6496]), .Z(n9257) );
  NANDN U12790 ( .A(y[6497]), .B(x[6497]), .Z(n23121) );
  AND U12791 ( .A(n9257), .B(n23121), .Z(n59183) );
  XNOR U12792 ( .A(x[6496]), .B(y[6496]), .Z(n23124) );
  NANDN U12793 ( .A(x[6495]), .B(y[6495]), .Z(n51050) );
  NANDN U12794 ( .A(y[6494]), .B(x[6494]), .Z(n9258) );
  NANDN U12795 ( .A(y[6495]), .B(x[6495]), .Z(n23123) );
  AND U12796 ( .A(n9258), .B(n23123), .Z(n59182) );
  XNOR U12797 ( .A(x[6494]), .B(y[6494]), .Z(n23126) );
  NANDN U12798 ( .A(x[6493]), .B(y[6493]), .Z(n59180) );
  NAND U12799 ( .A(n23126), .B(n59180), .Z(n19255) );
  XNOR U12800 ( .A(x[6492]), .B(y[6492]), .Z(n23128) );
  NANDN U12801 ( .A(y[6490]), .B(x[6490]), .Z(n9259) );
  NANDN U12802 ( .A(y[6491]), .B(x[6491]), .Z(n23127) );
  NAND U12803 ( .A(n9259), .B(n23127), .Z(n59176) );
  NANDN U12804 ( .A(y[6488]), .B(x[6488]), .Z(n9260) );
  NANDN U12805 ( .A(y[6489]), .B(x[6489]), .Z(n23129) );
  AND U12806 ( .A(n9260), .B(n23129), .Z(n59172) );
  XNOR U12807 ( .A(x[6488]), .B(y[6488]), .Z(n23132) );
  NANDN U12808 ( .A(y[6486]), .B(x[6486]), .Z(n9261) );
  NANDN U12809 ( .A(y[6487]), .B(x[6487]), .Z(n23131) );
  NAND U12810 ( .A(n9261), .B(n23131), .Z(n59168) );
  XNOR U12811 ( .A(x[6486]), .B(y[6486]), .Z(n23134) );
  NANDN U12812 ( .A(x[6485]), .B(y[6485]), .Z(n59164) );
  AND U12813 ( .A(n23134), .B(n59164), .Z(n19242) );
  NANDN U12814 ( .A(y[6484]), .B(x[6484]), .Z(n9262) );
  NANDN U12815 ( .A(y[6485]), .B(x[6485]), .Z(n23133) );
  NAND U12816 ( .A(n9262), .B(n23133), .Z(n59161) );
  XNOR U12817 ( .A(x[6484]), .B(y[6484]), .Z(n23136) );
  NANDN U12818 ( .A(y[6482]), .B(x[6482]), .Z(n9263) );
  NANDN U12819 ( .A(y[6483]), .B(x[6483]), .Z(n23135) );
  AND U12820 ( .A(n9263), .B(n23135), .Z(n59156) );
  XNOR U12821 ( .A(x[6482]), .B(y[6482]), .Z(n23138) );
  NANDN U12822 ( .A(x[6481]), .B(y[6481]), .Z(n59154) );
  NAND U12823 ( .A(n23138), .B(n59154), .Z(n19236) );
  NANDN U12824 ( .A(y[6480]), .B(x[6480]), .Z(n9264) );
  NANDN U12825 ( .A(y[6481]), .B(x[6481]), .Z(n23137) );
  AND U12826 ( .A(n9264), .B(n23137), .Z(n59150) );
  XOR U12827 ( .A(x[6480]), .B(y[6480]), .Z(n46347) );
  NANDN U12828 ( .A(x[6479]), .B(y[6479]), .Z(n23139) );
  IV U12829 ( .A(n23139), .Z(n51054) );
  OR U12830 ( .A(n46347), .B(n51054), .Z(n19233) );
  NANDN U12831 ( .A(y[6478]), .B(x[6478]), .Z(n9265) );
  ANDN U12832 ( .B(x[6479]), .A(y[6479]), .Z(n46346) );
  ANDN U12833 ( .B(n9265), .A(n46346), .Z(n59145) );
  XNOR U12834 ( .A(x[6478]), .B(y[6478]), .Z(n23141) );
  XNOR U12835 ( .A(x[6476]), .B(y[6476]), .Z(n23143) );
  NANDN U12836 ( .A(y[6474]), .B(x[6474]), .Z(n9266) );
  NANDN U12837 ( .A(y[6475]), .B(x[6475]), .Z(n23142) );
  NAND U12838 ( .A(n9266), .B(n23142), .Z(n59134) );
  XNOR U12839 ( .A(x[6474]), .B(y[6474]), .Z(n23145) );
  NANDN U12840 ( .A(x[6473]), .B(y[6473]), .Z(n59133) );
  NANDN U12841 ( .A(y[6472]), .B(x[6472]), .Z(n9267) );
  NANDN U12842 ( .A(y[6473]), .B(x[6473]), .Z(n23144) );
  AND U12843 ( .A(n9267), .B(n23144), .Z(n59131) );
  ANDN U12844 ( .B(y[6471]), .A(x[6471]), .Z(n46324) );
  XOR U12845 ( .A(x[6472]), .B(y[6472]), .Z(n9268) );
  NOR U12846 ( .A(n46324), .B(n9268), .Z(n19220) );
  XNOR U12847 ( .A(x[6470]), .B(y[6470]), .Z(n23147) );
  XNOR U12848 ( .A(x[6468]), .B(y[6468]), .Z(n23149) );
  NANDN U12849 ( .A(y[6466]), .B(x[6466]), .Z(n9269) );
  NANDN U12850 ( .A(y[6467]), .B(x[6467]), .Z(n23148) );
  NAND U12851 ( .A(n9269), .B(n23148), .Z(n59124) );
  XNOR U12852 ( .A(x[6466]), .B(y[6466]), .Z(n23151) );
  NANDN U12853 ( .A(x[6465]), .B(y[6465]), .Z(n59123) );
  NANDN U12854 ( .A(y[6464]), .B(x[6464]), .Z(n9270) );
  NANDN U12855 ( .A(y[6465]), .B(x[6465]), .Z(n23150) );
  AND U12856 ( .A(n9270), .B(n23150), .Z(n59121) );
  XNOR U12857 ( .A(x[6464]), .B(y[6464]), .Z(n23153) );
  ANDN U12858 ( .B(y[6463]), .A(x[6463]), .Z(n23154) );
  ANDN U12859 ( .B(n23153), .A(n23154), .Z(n19206) );
  XNOR U12860 ( .A(x[6462]), .B(y[6462]), .Z(n23156) );
  XNOR U12861 ( .A(x[6460]), .B(y[6460]), .Z(n23158) );
  NANDN U12862 ( .A(y[6458]), .B(x[6458]), .Z(n9271) );
  NANDN U12863 ( .A(y[6459]), .B(x[6459]), .Z(n23157) );
  NAND U12864 ( .A(n9271), .B(n23157), .Z(n59113) );
  NANDN U12865 ( .A(x[6457]), .B(y[6457]), .Z(n59112) );
  XNOR U12866 ( .A(x[6458]), .B(y[6458]), .Z(n23160) );
  NANDN U12867 ( .A(y[6456]), .B(x[6456]), .Z(n23162) );
  NANDN U12868 ( .A(y[6457]), .B(x[6457]), .Z(n23159) );
  AND U12869 ( .A(n23162), .B(n23159), .Z(n59110) );
  NANDN U12870 ( .A(x[6455]), .B(y[6455]), .Z(n23164) );
  NANDN U12871 ( .A(x[6456]), .B(y[6456]), .Z(n23161) );
  NAND U12872 ( .A(n23164), .B(n23161), .Z(n59109) );
  NANDN U12873 ( .A(y[6454]), .B(x[6454]), .Z(n23166) );
  NANDN U12874 ( .A(y[6455]), .B(x[6455]), .Z(n23163) );
  AND U12875 ( .A(n23166), .B(n23163), .Z(n59108) );
  NANDN U12876 ( .A(x[6453]), .B(y[6453]), .Z(n46287) );
  NANDN U12877 ( .A(x[6454]), .B(y[6454]), .Z(n23165) );
  NAND U12878 ( .A(n46287), .B(n23165), .Z(n59107) );
  NANDN U12879 ( .A(y[6452]), .B(x[6452]), .Z(n9272) );
  NANDN U12880 ( .A(y[6453]), .B(x[6453]), .Z(n23167) );
  AND U12881 ( .A(n9272), .B(n23167), .Z(n59106) );
  NANDN U12882 ( .A(y[6450]), .B(x[6450]), .Z(n9273) );
  NANDN U12883 ( .A(y[6451]), .B(x[6451]), .Z(n46285) );
  NAND U12884 ( .A(n9273), .B(n46285), .Z(n59102) );
  XNOR U12885 ( .A(x[6450]), .B(y[6450]), .Z(n23169) );
  ANDN U12886 ( .B(y[6449]), .A(x[6449]), .Z(n46276) );
  NANDN U12887 ( .A(x[6447]), .B(y[6447]), .Z(n59097) );
  XNOR U12888 ( .A(x[6448]), .B(y[6448]), .Z(n23171) );
  AND U12889 ( .A(n59097), .B(n23171), .Z(n19181) );
  NANDN U12890 ( .A(y[6446]), .B(x[6446]), .Z(n9274) );
  NANDN U12891 ( .A(y[6447]), .B(x[6447]), .Z(n23170) );
  NAND U12892 ( .A(n9274), .B(n23170), .Z(n59096) );
  XNOR U12893 ( .A(y[6446]), .B(x[6446]), .Z(n23174) );
  NANDN U12894 ( .A(x[6445]), .B(y[6445]), .Z(n23175) );
  AND U12895 ( .A(n23174), .B(n23175), .Z(n59095) );
  NANDN U12896 ( .A(y[6444]), .B(x[6444]), .Z(n23177) );
  NANDN U12897 ( .A(y[6445]), .B(x[6445]), .Z(n23173) );
  NAND U12898 ( .A(n23177), .B(n23173), .Z(n59094) );
  NANDN U12899 ( .A(x[6443]), .B(y[6443]), .Z(n46264) );
  NANDN U12900 ( .A(x[6444]), .B(y[6444]), .Z(n23176) );
  AND U12901 ( .A(n46264), .B(n23176), .Z(n59093) );
  NANDN U12902 ( .A(y[6442]), .B(x[6442]), .Z(n9275) );
  NANDN U12903 ( .A(y[6443]), .B(x[6443]), .Z(n23178) );
  NAND U12904 ( .A(n9275), .B(n23178), .Z(n59092) );
  NANDN U12905 ( .A(y[6440]), .B(x[6440]), .Z(n9276) );
  NANDN U12906 ( .A(y[6441]), .B(x[6441]), .Z(n23179) );
  AND U12907 ( .A(n9276), .B(n23179), .Z(n59089) );
  XNOR U12908 ( .A(x[6440]), .B(y[6440]), .Z(n23182) );
  NANDN U12909 ( .A(y[6439]), .B(x[6439]), .Z(n23181) );
  ANDN U12910 ( .B(x[6438]), .A(y[6438]), .Z(n46254) );
  ANDN U12911 ( .B(n23181), .A(n46254), .Z(n59086) );
  NANDN U12912 ( .A(y[6437]), .B(x[6437]), .Z(n46250) );
  NANDN U12913 ( .A(y[6436]), .B(x[6436]), .Z(n9277) );
  AND U12914 ( .A(n46250), .B(n9277), .Z(n59085) );
  NANDN U12915 ( .A(x[6435]), .B(y[6435]), .Z(n23186) );
  NANDN U12916 ( .A(x[6436]), .B(y[6436]), .Z(n46248) );
  NAND U12917 ( .A(n23186), .B(n46248), .Z(n59082) );
  NANDN U12918 ( .A(y[6434]), .B(x[6434]), .Z(n23188) );
  NANDN U12919 ( .A(y[6435]), .B(x[6435]), .Z(n23185) );
  AND U12920 ( .A(n23188), .B(n23185), .Z(n51063) );
  XNOR U12921 ( .A(y[6430]), .B(x[6430]), .Z(n23194) );
  NANDN U12922 ( .A(x[6429]), .B(y[6429]), .Z(n23195) );
  AND U12923 ( .A(n23194), .B(n23195), .Z(n59079) );
  XNOR U12924 ( .A(x[6428]), .B(y[6428]), .Z(n23197) );
  NANDN U12925 ( .A(y[6426]), .B(x[6426]), .Z(n9278) );
  NANDN U12926 ( .A(y[6427]), .B(x[6427]), .Z(n23196) );
  NAND U12927 ( .A(n9278), .B(n23196), .Z(n59075) );
  XNOR U12928 ( .A(x[6426]), .B(y[6426]), .Z(n23199) );
  NANDN U12929 ( .A(y[6424]), .B(x[6424]), .Z(n9279) );
  NANDN U12930 ( .A(y[6425]), .B(x[6425]), .Z(n23198) );
  NAND U12931 ( .A(n9279), .B(n23198), .Z(n59074) );
  NANDN U12932 ( .A(x[6423]), .B(y[6423]), .Z(n59071) );
  XNOR U12933 ( .A(x[6424]), .B(y[6424]), .Z(n23201) );
  NANDN U12934 ( .A(y[6422]), .B(x[6422]), .Z(n9280) );
  NANDN U12935 ( .A(y[6423]), .B(x[6423]), .Z(n23200) );
  AND U12936 ( .A(n9280), .B(n23200), .Z(n59070) );
  XNOR U12937 ( .A(x[6422]), .B(y[6422]), .Z(n23203) );
  ANDN U12938 ( .B(y[6421]), .A(x[6421]), .Z(n23204) );
  ANDN U12939 ( .B(n23203), .A(n23204), .Z(n19145) );
  ANDN U12940 ( .B(x[6419]), .A(y[6419]), .Z(n46210) );
  NANDN U12941 ( .A(y[6418]), .B(x[6418]), .Z(n9281) );
  NANDN U12942 ( .A(n46210), .B(n9281), .Z(n59065) );
  ANDN U12943 ( .B(y[6417]), .A(x[6417]), .Z(n51070) );
  XNOR U12944 ( .A(x[6418]), .B(y[6418]), .Z(n23206) );
  NANDN U12945 ( .A(y[6416]), .B(x[6416]), .Z(n9282) );
  NANDN U12946 ( .A(y[6417]), .B(x[6417]), .Z(n23205) );
  NAND U12947 ( .A(n9282), .B(n23205), .Z(n59064) );
  XNOR U12948 ( .A(x[6416]), .B(y[6416]), .Z(n46200) );
  ANDN U12949 ( .B(y[6415]), .A(x[6415]), .Z(n46196) );
  NANDN U12950 ( .A(x[6413]), .B(y[6413]), .Z(n59057) );
  XNOR U12951 ( .A(x[6414]), .B(y[6414]), .Z(n23208) );
  AND U12952 ( .A(n59057), .B(n23208), .Z(n19131) );
  NANDN U12953 ( .A(y[6412]), .B(x[6412]), .Z(n9283) );
  NANDN U12954 ( .A(y[6413]), .B(x[6413]), .Z(n23207) );
  NAND U12955 ( .A(n9283), .B(n23207), .Z(n59056) );
  XNOR U12956 ( .A(x[6412]), .B(y[6412]), .Z(n23210) );
  NANDN U12957 ( .A(y[6410]), .B(x[6410]), .Z(n9284) );
  NANDN U12958 ( .A(y[6411]), .B(x[6411]), .Z(n23209) );
  NAND U12959 ( .A(n9284), .B(n23209), .Z(n59053) );
  ANDN U12960 ( .B(y[6409]), .A(x[6409]), .Z(n51072) );
  XNOR U12961 ( .A(x[6410]), .B(y[6410]), .Z(n23212) );
  NANDN U12962 ( .A(y[6408]), .B(x[6408]), .Z(n9285) );
  NANDN U12963 ( .A(y[6409]), .B(x[6409]), .Z(n23211) );
  NAND U12964 ( .A(n9285), .B(n23211), .Z(n59052) );
  XNOR U12965 ( .A(x[6408]), .B(y[6408]), .Z(n46181) );
  NANDN U12966 ( .A(x[6407]), .B(y[6407]), .Z(n59050) );
  NANDN U12967 ( .A(y[6406]), .B(x[6406]), .Z(n9286) );
  NANDN U12968 ( .A(y[6407]), .B(x[6407]), .Z(n46180) );
  AND U12969 ( .A(n9286), .B(n46180), .Z(n59049) );
  XNOR U12970 ( .A(x[6406]), .B(y[6406]), .Z(n23214) );
  ANDN U12971 ( .B(y[6405]), .A(x[6405]), .Z(n59048) );
  ANDN U12972 ( .B(n23214), .A(n59048), .Z(n19119) );
  NANDN U12973 ( .A(y[6404]), .B(x[6404]), .Z(n9287) );
  NANDN U12974 ( .A(y[6405]), .B(x[6405]), .Z(n23213) );
  NAND U12975 ( .A(n9287), .B(n23213), .Z(n59047) );
  XNOR U12976 ( .A(x[6404]), .B(y[6404]), .Z(n46171) );
  NANDN U12977 ( .A(y[6402]), .B(x[6402]), .Z(n9288) );
  NANDN U12978 ( .A(y[6403]), .B(x[6403]), .Z(n46170) );
  NAND U12979 ( .A(n9288), .B(n46170), .Z(n59041) );
  XNOR U12980 ( .A(x[6402]), .B(y[6402]), .Z(n23216) );
  NANDN U12981 ( .A(y[6400]), .B(x[6400]), .Z(n9289) );
  NANDN U12982 ( .A(y[6401]), .B(x[6401]), .Z(n23215) );
  NAND U12983 ( .A(n9289), .B(n23215), .Z(n59040) );
  XNOR U12984 ( .A(x[6400]), .B(y[6400]), .Z(n23218) );
  ANDN U12985 ( .B(y[6399]), .A(x[6399]), .Z(n46159) );
  XNOR U12986 ( .A(x[6398]), .B(y[6398]), .Z(n23220) );
  ANDN U12987 ( .B(y[6397]), .A(x[6397]), .Z(n59035) );
  ANDN U12988 ( .B(n23220), .A(n59035), .Z(n19106) );
  XNOR U12989 ( .A(x[6396]), .B(y[6396]), .Z(n46152) );
  NANDN U12990 ( .A(y[6394]), .B(x[6394]), .Z(n9290) );
  NANDN U12991 ( .A(y[6395]), .B(x[6395]), .Z(n46151) );
  NAND U12992 ( .A(n9290), .B(n46151), .Z(n59034) );
  ANDN U12993 ( .B(y[6393]), .A(x[6393]), .Z(n51080) );
  XNOR U12994 ( .A(x[6394]), .B(y[6394]), .Z(n23222) );
  NANDN U12995 ( .A(y[6392]), .B(x[6392]), .Z(n9291) );
  NANDN U12996 ( .A(y[6393]), .B(x[6393]), .Z(n23221) );
  NAND U12997 ( .A(n9291), .B(n23221), .Z(n59033) );
  XNOR U12998 ( .A(x[6392]), .B(y[6392]), .Z(n46142) );
  ANDN U12999 ( .B(y[6391]), .A(x[6391]), .Z(n46138) );
  XNOR U13000 ( .A(x[6390]), .B(y[6390]), .Z(n23224) );
  ANDN U13001 ( .B(y[6389]), .A(x[6389]), .Z(n59026) );
  ANDN U13002 ( .B(n23224), .A(n59026), .Z(n19092) );
  NANDN U13003 ( .A(y[6388]), .B(x[6388]), .Z(n9292) );
  NANDN U13004 ( .A(y[6389]), .B(x[6389]), .Z(n23223) );
  NAND U13005 ( .A(n9292), .B(n23223), .Z(n59025) );
  XNOR U13006 ( .A(x[6388]), .B(y[6388]), .Z(n46131) );
  NANDN U13007 ( .A(y[6386]), .B(x[6386]), .Z(n9293) );
  NANDN U13008 ( .A(y[6387]), .B(x[6387]), .Z(n46130) );
  NAND U13009 ( .A(n9293), .B(n46130), .Z(n59022) );
  ANDN U13010 ( .B(y[6385]), .A(x[6385]), .Z(n51082) );
  XNOR U13011 ( .A(x[6386]), .B(y[6386]), .Z(n23226) );
  NANDN U13012 ( .A(y[6384]), .B(x[6384]), .Z(n9294) );
  NANDN U13013 ( .A(y[6385]), .B(x[6385]), .Z(n23225) );
  NAND U13014 ( .A(n9294), .B(n23225), .Z(n59021) );
  NANDN U13015 ( .A(x[6383]), .B(y[6383]), .Z(n59019) );
  XNOR U13016 ( .A(x[6384]), .B(y[6384]), .Z(n46121) );
  NANDN U13017 ( .A(y[6382]), .B(x[6382]), .Z(n9295) );
  NANDN U13018 ( .A(y[6383]), .B(x[6383]), .Z(n46120) );
  AND U13019 ( .A(n9295), .B(n46120), .Z(n59018) );
  XNOR U13020 ( .A(x[6382]), .B(y[6382]), .Z(n23228) );
  ANDN U13021 ( .B(y[6381]), .A(x[6381]), .Z(n59014) );
  ANDN U13022 ( .B(n23228), .A(n59014), .Z(n19080) );
  XNOR U13023 ( .A(x[6380]), .B(y[6380]), .Z(n46111) );
  NANDN U13024 ( .A(y[6378]), .B(x[6378]), .Z(n9296) );
  NANDN U13025 ( .A(y[6379]), .B(x[6379]), .Z(n46110) );
  NAND U13026 ( .A(n9296), .B(n46110), .Z(n59011) );
  NANDN U13027 ( .A(x[6377]), .B(y[6377]), .Z(n23231) );
  XNOR U13028 ( .A(x[6378]), .B(y[6378]), .Z(n23230) );
  NANDN U13029 ( .A(y[6376]), .B(x[6376]), .Z(n9297) );
  NANDN U13030 ( .A(y[6377]), .B(x[6377]), .Z(n23229) );
  NAND U13031 ( .A(n9297), .B(n23229), .Z(n59010) );
  XNOR U13032 ( .A(x[6376]), .B(y[6376]), .Z(n23233) );
  ANDN U13033 ( .B(y[6375]), .A(x[6375]), .Z(n23234) );
  NANDN U13034 ( .A(x[6373]), .B(y[6373]), .Z(n23238) );
  NANDN U13035 ( .A(x[6374]), .B(y[6374]), .Z(n23235) );
  NAND U13036 ( .A(n23238), .B(n23235), .Z(n51088) );
  NANDN U13037 ( .A(y[6372]), .B(x[6372]), .Z(n9298) );
  NANDN U13038 ( .A(y[6373]), .B(x[6373]), .Z(n23237) );
  AND U13039 ( .A(n9298), .B(n23237), .Z(n59007) );
  ANDN U13040 ( .B(y[6371]), .A(x[6371]), .Z(n46091) );
  XNOR U13041 ( .A(x[6372]), .B(y[6372]), .Z(n23240) );
  NANDN U13042 ( .A(y[6370]), .B(x[6370]), .Z(n9299) );
  NANDN U13043 ( .A(y[6371]), .B(x[6371]), .Z(n23239) );
  NAND U13044 ( .A(n9299), .B(n23239), .Z(n59004) );
  XNOR U13045 ( .A(x[6370]), .B(y[6370]), .Z(n23242) );
  ANDN U13046 ( .B(y[6369]), .A(x[6369]), .Z(n23243) );
  NANDN U13047 ( .A(y[6369]), .B(x[6369]), .Z(n23241) );
  ANDN U13048 ( .B(x[6368]), .A(y[6368]), .Z(n46084) );
  ANDN U13049 ( .B(n23241), .A(n46084), .Z(n59001) );
  NANDN U13050 ( .A(x[6367]), .B(y[6367]), .Z(n46082) );
  NANDN U13051 ( .A(x[6368]), .B(y[6368]), .Z(n23244) );
  AND U13052 ( .A(n46082), .B(n23244), .Z(n59000) );
  XNOR U13053 ( .A(x[6366]), .B(y[6366]), .Z(n23246) );
  XNOR U13054 ( .A(x[6364]), .B(y[6364]), .Z(n23248) );
  NANDN U13055 ( .A(y[6362]), .B(x[6362]), .Z(n23250) );
  NANDN U13056 ( .A(y[6363]), .B(x[6363]), .Z(n23247) );
  NAND U13057 ( .A(n23250), .B(n23247), .Z(n58995) );
  NANDN U13058 ( .A(x[6362]), .B(y[6362]), .Z(n23249) );
  ANDN U13059 ( .B(y[6361]), .A(x[6361]), .Z(n23252) );
  ANDN U13060 ( .B(n23249), .A(n23252), .Z(n58994) );
  NANDN U13061 ( .A(y[6360]), .B(x[6360]), .Z(n9300) );
  NANDN U13062 ( .A(y[6361]), .B(x[6361]), .Z(n23251) );
  NAND U13063 ( .A(n9300), .B(n23251), .Z(n58993) );
  NANDN U13064 ( .A(y[6358]), .B(x[6358]), .Z(n9301) );
  NANDN U13065 ( .A(y[6359]), .B(x[6359]), .Z(n46064) );
  AND U13066 ( .A(n9301), .B(n46064), .Z(n58992) );
  XNOR U13067 ( .A(x[6358]), .B(y[6358]), .Z(n23254) );
  NANDN U13068 ( .A(y[6356]), .B(x[6356]), .Z(n9302) );
  NANDN U13069 ( .A(y[6357]), .B(x[6357]), .Z(n23253) );
  AND U13070 ( .A(n9302), .B(n23253), .Z(n58988) );
  ANDN U13071 ( .B(y[6355]), .A(x[6355]), .Z(n46051) );
  XNOR U13072 ( .A(x[6356]), .B(y[6356]), .Z(n46055) );
  NANDN U13073 ( .A(y[6354]), .B(x[6354]), .Z(n9303) );
  NANDN U13074 ( .A(y[6355]), .B(x[6355]), .Z(n46054) );
  NAND U13075 ( .A(n9303), .B(n46054), .Z(n58985) );
  XNOR U13076 ( .A(x[6354]), .B(y[6354]), .Z(n23256) );
  ANDN U13077 ( .B(y[6353]), .A(x[6353]), .Z(n58984) );
  NANDN U13078 ( .A(y[6352]), .B(x[6352]), .Z(n9304) );
  NANDN U13079 ( .A(y[6353]), .B(x[6353]), .Z(n23255) );
  AND U13080 ( .A(n9304), .B(n23255), .Z(n58982) );
  NANDN U13081 ( .A(x[6351]), .B(y[6351]), .Z(n51096) );
  XNOR U13082 ( .A(x[6352]), .B(y[6352]), .Z(n46044) );
  AND U13083 ( .A(n51096), .B(n46044), .Z(n19035) );
  NANDN U13084 ( .A(y[6350]), .B(x[6350]), .Z(n9305) );
  NANDN U13085 ( .A(y[6351]), .B(x[6351]), .Z(n46043) );
  NAND U13086 ( .A(n9305), .B(n46043), .Z(n58981) );
  XNOR U13087 ( .A(x[6350]), .B(y[6350]), .Z(n23258) );
  NANDN U13088 ( .A(y[6348]), .B(x[6348]), .Z(n9306) );
  NANDN U13089 ( .A(y[6349]), .B(x[6349]), .Z(n23257) );
  NAND U13090 ( .A(n9306), .B(n23257), .Z(n58978) );
  XNOR U13091 ( .A(x[6348]), .B(y[6348]), .Z(n46034) );
  NANDN U13092 ( .A(y[6346]), .B(x[6346]), .Z(n23260) );
  NANDN U13093 ( .A(y[6347]), .B(x[6347]), .Z(n46033) );
  NAND U13094 ( .A(n23260), .B(n46033), .Z(n58973) );
  NANDN U13095 ( .A(x[6346]), .B(y[6346]), .Z(n23259) );
  ANDN U13096 ( .B(y[6345]), .A(x[6345]), .Z(n46026) );
  ANDN U13097 ( .B(n23259), .A(n46026), .Z(n58972) );
  NANDN U13098 ( .A(y[6342]), .B(x[6342]), .Z(n23266) );
  NANDN U13099 ( .A(y[6343]), .B(x[6343]), .Z(n23263) );
  NAND U13100 ( .A(n23266), .B(n23263), .Z(n58969) );
  NANDN U13101 ( .A(x[6342]), .B(y[6342]), .Z(n23265) );
  ANDN U13102 ( .B(y[6341]), .A(x[6341]), .Z(n46017) );
  ANDN U13103 ( .B(n23265), .A(n46017), .Z(n58968) );
  XNOR U13104 ( .A(x[6340]), .B(y[6340]), .Z(n23269) );
  NANDN U13105 ( .A(x[6339]), .B(y[6339]), .Z(n51098) );
  AND U13106 ( .A(n23269), .B(n51098), .Z(n19019) );
  NANDN U13107 ( .A(x[6337]), .B(y[6337]), .Z(n23273) );
  NANDN U13108 ( .A(x[6338]), .B(y[6338]), .Z(n23270) );
  AND U13109 ( .A(n23273), .B(n23270), .Z(n58965) );
  ANDN U13110 ( .B(x[6336]), .A(y[6336]), .Z(n46005) );
  NANDN U13111 ( .A(y[6337]), .B(x[6337]), .Z(n23272) );
  NANDN U13112 ( .A(n46005), .B(n23272), .Z(n58964) );
  NANDN U13113 ( .A(x[6335]), .B(y[6335]), .Z(n23275) );
  NANDN U13114 ( .A(x[6336]), .B(y[6336]), .Z(n23274) );
  AND U13115 ( .A(n23275), .B(n23274), .Z(n58963) );
  ANDN U13116 ( .B(x[6335]), .A(y[6335]), .Z(n46007) );
  NANDN U13117 ( .A(y[6334]), .B(x[6334]), .Z(n23277) );
  NANDN U13118 ( .A(n46007), .B(n23277), .Z(n58962) );
  NANDN U13119 ( .A(x[6334]), .B(y[6334]), .Z(n23276) );
  ANDN U13120 ( .B(y[6333]), .A(x[6333]), .Z(n45997) );
  ANDN U13121 ( .B(n23276), .A(n45997), .Z(n58961) );
  NANDN U13122 ( .A(x[6331]), .B(y[6331]), .Z(n23281) );
  NANDN U13123 ( .A(x[6332]), .B(y[6332]), .Z(n45999) );
  AND U13124 ( .A(n23281), .B(n45999), .Z(n58959) );
  NANDN U13125 ( .A(y[6330]), .B(x[6330]), .Z(n23283) );
  NANDN U13126 ( .A(y[6331]), .B(x[6331]), .Z(n23280) );
  NAND U13127 ( .A(n23283), .B(n23280), .Z(n58958) );
  NANDN U13128 ( .A(x[6329]), .B(y[6329]), .Z(n23286) );
  NANDN U13129 ( .A(x[6330]), .B(y[6330]), .Z(n23282) );
  AND U13130 ( .A(n23286), .B(n23282), .Z(n58956) );
  NANDN U13131 ( .A(y[6328]), .B(x[6328]), .Z(n23287) );
  NANDN U13132 ( .A(y[6329]), .B(x[6329]), .Z(n23284) );
  NAND U13133 ( .A(n23287), .B(n23284), .Z(n58955) );
  NANDN U13134 ( .A(x[6327]), .B(y[6327]), .Z(n23289) );
  NANDN U13135 ( .A(x[6328]), .B(y[6328]), .Z(n23285) );
  AND U13136 ( .A(n23289), .B(n23285), .Z(n58954) );
  NANDN U13137 ( .A(y[6326]), .B(x[6326]), .Z(n9307) );
  NANDN U13138 ( .A(y[6327]), .B(x[6327]), .Z(n23288) );
  NAND U13139 ( .A(n9307), .B(n23288), .Z(n58953) );
  ANDN U13140 ( .B(y[6325]), .A(x[6325]), .Z(n58951) );
  XNOR U13141 ( .A(x[6326]), .B(y[6326]), .Z(n23291) );
  NANDN U13142 ( .A(y[6324]), .B(x[6324]), .Z(n9308) );
  NANDN U13143 ( .A(y[6325]), .B(x[6325]), .Z(n23290) );
  NAND U13144 ( .A(n9308), .B(n23290), .Z(n58950) );
  XNOR U13145 ( .A(x[6324]), .B(y[6324]), .Z(n45977) );
  NANDN U13146 ( .A(x[6323]), .B(y[6323]), .Z(n58949) );
  NANDN U13147 ( .A(y[6322]), .B(x[6322]), .Z(n9309) );
  NANDN U13148 ( .A(y[6323]), .B(x[6323]), .Z(n45976) );
  AND U13149 ( .A(n9309), .B(n45976), .Z(n58947) );
  XNOR U13150 ( .A(x[6322]), .B(y[6322]), .Z(n23293) );
  ANDN U13151 ( .B(y[6321]), .A(x[6321]), .Z(n51100) );
  ANDN U13152 ( .B(n23293), .A(n51100), .Z(n18998) );
  XNOR U13153 ( .A(x[6320]), .B(y[6320]), .Z(n45967) );
  XNOR U13154 ( .A(x[6318]), .B(y[6318]), .Z(n23295) );
  NANDN U13155 ( .A(y[6316]), .B(x[6316]), .Z(n9310) );
  NANDN U13156 ( .A(y[6317]), .B(x[6317]), .Z(n23294) );
  NAND U13157 ( .A(n9310), .B(n23294), .Z(n58939) );
  XNOR U13158 ( .A(x[6316]), .B(y[6316]), .Z(n45957) );
  NANDN U13159 ( .A(x[6315]), .B(y[6315]), .Z(n58938) );
  NANDN U13160 ( .A(y[6314]), .B(x[6314]), .Z(n9311) );
  NANDN U13161 ( .A(y[6315]), .B(x[6315]), .Z(n45956) );
  AND U13162 ( .A(n9311), .B(n45956), .Z(n58936) );
  ANDN U13163 ( .B(y[6313]), .A(x[6313]), .Z(n51102) );
  NANDN U13164 ( .A(y[6312]), .B(x[6312]), .Z(n9312) );
  NANDN U13165 ( .A(y[6313]), .B(x[6313]), .Z(n23296) );
  AND U13166 ( .A(n9312), .B(n23296), .Z(n58935) );
  ANDN U13167 ( .B(y[6311]), .A(x[6311]), .Z(n45943) );
  XNOR U13168 ( .A(x[6312]), .B(y[6312]), .Z(n45947) );
  XNOR U13169 ( .A(x[6310]), .B(y[6310]), .Z(n23299) );
  NANDN U13170 ( .A(y[6308]), .B(x[6308]), .Z(n9313) );
  NANDN U13171 ( .A(y[6309]), .B(x[6309]), .Z(n23298) );
  NAND U13172 ( .A(n9313), .B(n23298), .Z(n51104) );
  XNOR U13173 ( .A(x[6308]), .B(y[6308]), .Z(n45936) );
  NANDN U13174 ( .A(x[6307]), .B(y[6307]), .Z(n51106) );
  NANDN U13175 ( .A(y[6306]), .B(x[6306]), .Z(n9314) );
  NANDN U13176 ( .A(y[6307]), .B(x[6307]), .Z(n45935) );
  AND U13177 ( .A(n9314), .B(n45935), .Z(n58929) );
  XNOR U13178 ( .A(x[6306]), .B(y[6306]), .Z(n23301) );
  ANDN U13179 ( .B(y[6305]), .A(x[6305]), .Z(n51107) );
  ANDN U13180 ( .B(n23301), .A(n51107), .Z(n18971) );
  XNOR U13181 ( .A(x[6304]), .B(y[6304]), .Z(n45926) );
  XNOR U13182 ( .A(x[6302]), .B(y[6302]), .Z(n23303) );
  NANDN U13183 ( .A(y[6300]), .B(x[6300]), .Z(n9315) );
  NANDN U13184 ( .A(y[6301]), .B(x[6301]), .Z(n23302) );
  NAND U13185 ( .A(n9315), .B(n23302), .Z(n58920) );
  XNOR U13186 ( .A(x[6300]), .B(y[6300]), .Z(n23305) );
  NANDN U13187 ( .A(x[6299]), .B(y[6299]), .Z(n58919) );
  NANDN U13188 ( .A(y[6298]), .B(x[6298]), .Z(n9316) );
  NANDN U13189 ( .A(y[6299]), .B(x[6299]), .Z(n23304) );
  AND U13190 ( .A(n9316), .B(n23304), .Z(n58917) );
  XNOR U13191 ( .A(x[6298]), .B(y[6298]), .Z(n23307) );
  ANDN U13192 ( .B(y[6297]), .A(x[6297]), .Z(n51109) );
  ANDN U13193 ( .B(n23307), .A(n51109), .Z(n18957) );
  XNOR U13194 ( .A(x[6296]), .B(y[6296]), .Z(n45908) );
  XNOR U13195 ( .A(x[6294]), .B(y[6294]), .Z(n23309) );
  NANDN U13196 ( .A(y[6292]), .B(x[6292]), .Z(n9317) );
  NANDN U13197 ( .A(y[6293]), .B(x[6293]), .Z(n23308) );
  NAND U13198 ( .A(n9317), .B(n23308), .Z(n58909) );
  XNOR U13199 ( .A(x[6292]), .B(y[6292]), .Z(n23311) );
  NANDN U13200 ( .A(x[6291]), .B(y[6291]), .Z(n58908) );
  NANDN U13201 ( .A(y[6290]), .B(x[6290]), .Z(n9318) );
  NANDN U13202 ( .A(y[6291]), .B(x[6291]), .Z(n23310) );
  AND U13203 ( .A(n9318), .B(n23310), .Z(n58906) );
  XNOR U13204 ( .A(x[6290]), .B(y[6290]), .Z(n23313) );
  ANDN U13205 ( .B(y[6289]), .A(x[6289]), .Z(n23314) );
  ANDN U13206 ( .B(n23313), .A(n23314), .Z(n18943) );
  XNOR U13207 ( .A(x[6288]), .B(y[6288]), .Z(n23316) );
  XNOR U13208 ( .A(x[6286]), .B(y[6286]), .Z(n23318) );
  NANDN U13209 ( .A(y[6284]), .B(x[6284]), .Z(n9319) );
  NANDN U13210 ( .A(y[6285]), .B(x[6285]), .Z(n23317) );
  NAND U13211 ( .A(n9319), .B(n23317), .Z(n58899) );
  XNOR U13212 ( .A(x[6284]), .B(y[6284]), .Z(n45882) );
  NANDN U13213 ( .A(x[6283]), .B(y[6283]), .Z(n58898) );
  NANDN U13214 ( .A(y[6282]), .B(x[6282]), .Z(n9320) );
  NANDN U13215 ( .A(y[6283]), .B(x[6283]), .Z(n45881) );
  AND U13216 ( .A(n9320), .B(n45881), .Z(n58896) );
  XNOR U13217 ( .A(x[6282]), .B(y[6282]), .Z(n23320) );
  ANDN U13218 ( .B(y[6281]), .A(x[6281]), .Z(n23321) );
  ANDN U13219 ( .B(n23320), .A(n23321), .Z(n18929) );
  NANDN U13220 ( .A(y[6278]), .B(x[6278]), .Z(n9321) );
  ANDN U13221 ( .B(x[6279]), .A(y[6279]), .Z(n45874) );
  ANDN U13222 ( .B(n9321), .A(n45874), .Z(n58891) );
  ANDN U13223 ( .B(y[6277]), .A(x[6277]), .Z(n58889) );
  XNOR U13224 ( .A(x[6278]), .B(y[6278]), .Z(n23323) );
  NANDN U13225 ( .A(y[6276]), .B(x[6276]), .Z(n9322) );
  NANDN U13226 ( .A(y[6277]), .B(x[6277]), .Z(n23322) );
  NAND U13227 ( .A(n9322), .B(n23322), .Z(n58888) );
  XNOR U13228 ( .A(x[6276]), .B(y[6276]), .Z(n45862) );
  NANDN U13229 ( .A(x[6275]), .B(y[6275]), .Z(n58887) );
  NANDN U13230 ( .A(y[6274]), .B(x[6274]), .Z(n9323) );
  NANDN U13231 ( .A(y[6275]), .B(x[6275]), .Z(n45861) );
  AND U13232 ( .A(n9323), .B(n45861), .Z(n58885) );
  XNOR U13233 ( .A(x[6274]), .B(y[6274]), .Z(n23325) );
  ANDN U13234 ( .B(y[6273]), .A(x[6273]), .Z(n51115) );
  ANDN U13235 ( .B(n23325), .A(n51115), .Z(n18915) );
  XNOR U13236 ( .A(x[6272]), .B(y[6272]), .Z(n45852) );
  XNOR U13237 ( .A(x[6270]), .B(y[6270]), .Z(n23327) );
  NANDN U13238 ( .A(y[6268]), .B(x[6268]), .Z(n9324) );
  NANDN U13239 ( .A(y[6269]), .B(x[6269]), .Z(n23326) );
  NAND U13240 ( .A(n9324), .B(n23326), .Z(n58877) );
  XNOR U13241 ( .A(x[6264]), .B(y[6264]), .Z(n23333) );
  XNOR U13242 ( .A(x[6262]), .B(y[6262]), .Z(n23335) );
  NANDN U13243 ( .A(y[6260]), .B(x[6260]), .Z(n9325) );
  NANDN U13244 ( .A(y[6261]), .B(x[6261]), .Z(n23334) );
  NAND U13245 ( .A(n9325), .B(n23334), .Z(n58866) );
  XNOR U13246 ( .A(x[6260]), .B(y[6260]), .Z(n23337) );
  ANDN U13247 ( .B(y[6259]), .A(x[6259]), .Z(n45822) );
  XNOR U13248 ( .A(x[6258]), .B(y[6258]), .Z(n23339) );
  ANDN U13249 ( .B(y[6257]), .A(x[6257]), .Z(n58863) );
  XNOR U13250 ( .A(x[6256]), .B(y[6256]), .Z(n45815) );
  XNOR U13251 ( .A(x[6254]), .B(y[6254]), .Z(n23341) );
  NANDN U13252 ( .A(y[6252]), .B(x[6252]), .Z(n9326) );
  NANDN U13253 ( .A(y[6253]), .B(x[6253]), .Z(n23340) );
  NAND U13254 ( .A(n9326), .B(n23340), .Z(n58856) );
  XNOR U13255 ( .A(x[6252]), .B(y[6252]), .Z(n23343) );
  ANDN U13256 ( .B(y[6251]), .A(x[6251]), .Z(n23344) );
  NANDN U13257 ( .A(y[6248]), .B(x[6248]), .Z(n9327) );
  NANDN U13258 ( .A(y[6249]), .B(x[6249]), .Z(n23345) );
  AND U13259 ( .A(n9327), .B(n23345), .Z(n58851) );
  XNOR U13260 ( .A(x[6248]), .B(y[6248]), .Z(n23348) );
  ANDN U13261 ( .B(y[6247]), .A(x[6247]), .Z(n45795) );
  ANDN U13262 ( .B(n23348), .A(n45795), .Z(n18886) );
  XNOR U13263 ( .A(x[6246]), .B(y[6246]), .Z(n23350) );
  NANDN U13264 ( .A(y[6244]), .B(x[6244]), .Z(n23352) );
  NANDN U13265 ( .A(y[6245]), .B(x[6245]), .Z(n23349) );
  NAND U13266 ( .A(n23352), .B(n23349), .Z(n58847) );
  NANDN U13267 ( .A(x[6243]), .B(y[6243]), .Z(n23354) );
  NANDN U13268 ( .A(x[6244]), .B(y[6244]), .Z(n23351) );
  AND U13269 ( .A(n23354), .B(n23351), .Z(n51126) );
  XNOR U13270 ( .A(x[6240]), .B(y[6240]), .Z(n23360) );
  NANDN U13271 ( .A(y[6238]), .B(x[6238]), .Z(n9328) );
  NANDN U13272 ( .A(y[6239]), .B(x[6239]), .Z(n23359) );
  NAND U13273 ( .A(n9328), .B(n23359), .Z(n58841) );
  ANDN U13274 ( .B(y[6237]), .A(x[6237]), .Z(n51128) );
  XNOR U13275 ( .A(x[6238]), .B(y[6238]), .Z(n23362) );
  NANDN U13276 ( .A(y[6236]), .B(x[6236]), .Z(n9329) );
  NANDN U13277 ( .A(y[6237]), .B(x[6237]), .Z(n23361) );
  NAND U13278 ( .A(n9329), .B(n23361), .Z(n58840) );
  XNOR U13279 ( .A(x[6236]), .B(y[6236]), .Z(n45772) );
  NANDN U13280 ( .A(x[6235]), .B(y[6235]), .Z(n58838) );
  AND U13281 ( .A(n45772), .B(n58838), .Z(n18868) );
  NANDN U13282 ( .A(y[6234]), .B(x[6234]), .Z(n9330) );
  NANDN U13283 ( .A(y[6235]), .B(x[6235]), .Z(n45771) );
  NAND U13284 ( .A(n9330), .B(n45771), .Z(n58837) );
  NANDN U13285 ( .A(y[6232]), .B(x[6232]), .Z(n9331) );
  NANDN U13286 ( .A(y[6233]), .B(x[6233]), .Z(n23363) );
  AND U13287 ( .A(n9331), .B(n23363), .Z(n51130) );
  XNOR U13288 ( .A(x[6232]), .B(y[6232]), .Z(n45762) );
  XNOR U13289 ( .A(x[6230]), .B(y[6230]), .Z(n23366) );
  NANDN U13290 ( .A(y[6228]), .B(x[6228]), .Z(n9332) );
  NANDN U13291 ( .A(y[6229]), .B(x[6229]), .Z(n23365) );
  NAND U13292 ( .A(n9332), .B(n23365), .Z(n58829) );
  XNOR U13293 ( .A(x[6228]), .B(y[6228]), .Z(n45752) );
  NANDN U13294 ( .A(x[6227]), .B(y[6227]), .Z(n58827) );
  AND U13295 ( .A(n45752), .B(n58827), .Z(n18855) );
  NANDN U13296 ( .A(y[6226]), .B(x[6226]), .Z(n9333) );
  NANDN U13297 ( .A(y[6227]), .B(x[6227]), .Z(n45751) );
  NAND U13298 ( .A(n9333), .B(n45751), .Z(n58826) );
  XNOR U13299 ( .A(y[6226]), .B(x[6226]), .Z(n23369) );
  NANDN U13300 ( .A(x[6225]), .B(y[6225]), .Z(n23370) );
  AND U13301 ( .A(n23369), .B(n23370), .Z(n58825) );
  XNOR U13302 ( .A(x[6224]), .B(y[6224]), .Z(n23372) );
  XNOR U13303 ( .A(x[6222]), .B(y[6222]), .Z(n23374) );
  NANDN U13304 ( .A(y[6220]), .B(x[6220]), .Z(n9334) );
  NANDN U13305 ( .A(y[6221]), .B(x[6221]), .Z(n23373) );
  NAND U13306 ( .A(n9334), .B(n23373), .Z(n58820) );
  XNOR U13307 ( .A(x[6220]), .B(y[6220]), .Z(n45733) );
  ANDN U13308 ( .B(y[6219]), .A(x[6219]), .Z(n45729) );
  XNOR U13309 ( .A(x[6218]), .B(y[6218]), .Z(n23376) );
  ANDN U13310 ( .B(y[6217]), .A(x[6217]), .Z(n58816) );
  ANDN U13311 ( .B(n23376), .A(n58816), .Z(n18838) );
  XNOR U13312 ( .A(x[6216]), .B(y[6216]), .Z(n45722) );
  NANDN U13313 ( .A(y[6214]), .B(x[6214]), .Z(n9335) );
  NANDN U13314 ( .A(y[6215]), .B(x[6215]), .Z(n45721) );
  AND U13315 ( .A(n9335), .B(n45721), .Z(n58812) );
  ANDN U13316 ( .B(y[6213]), .A(x[6213]), .Z(n58810) );
  XNOR U13317 ( .A(x[6214]), .B(y[6214]), .Z(n23378) );
  NANDN U13318 ( .A(y[6212]), .B(x[6212]), .Z(n9336) );
  NANDN U13319 ( .A(y[6213]), .B(x[6213]), .Z(n23377) );
  NAND U13320 ( .A(n9336), .B(n23377), .Z(n58809) );
  XNOR U13321 ( .A(x[6212]), .B(y[6212]), .Z(n45712) );
  ANDN U13322 ( .B(y[6211]), .A(x[6211]), .Z(n45708) );
  XNOR U13323 ( .A(x[6210]), .B(y[6210]), .Z(n23380) );
  ANDN U13324 ( .B(y[6209]), .A(x[6209]), .Z(n51139) );
  ANDN U13325 ( .B(n23380), .A(n51139), .Z(n18824) );
  XNOR U13326 ( .A(x[6208]), .B(y[6208]), .Z(n45701) );
  XNOR U13327 ( .A(x[6206]), .B(y[6206]), .Z(n23382) );
  NANDN U13328 ( .A(y[6204]), .B(x[6204]), .Z(n9337) );
  NANDN U13329 ( .A(y[6205]), .B(x[6205]), .Z(n23381) );
  NAND U13330 ( .A(n9337), .B(n23381), .Z(n51142) );
  XNOR U13331 ( .A(x[6204]), .B(y[6204]), .Z(n45691) );
  ANDN U13332 ( .B(y[6203]), .A(x[6203]), .Z(n45687) );
  XNOR U13333 ( .A(x[6202]), .B(y[6202]), .Z(n23385) );
  ANDN U13334 ( .B(y[6201]), .A(x[6201]), .Z(n58798) );
  ANDN U13335 ( .B(n23385), .A(n58798), .Z(n18809) );
  XNOR U13336 ( .A(x[6200]), .B(y[6200]), .Z(n45680) );
  XNOR U13337 ( .A(x[6198]), .B(y[6198]), .Z(n23387) );
  NANDN U13338 ( .A(y[6196]), .B(x[6196]), .Z(n9338) );
  NANDN U13339 ( .A(y[6197]), .B(x[6197]), .Z(n23386) );
  NAND U13340 ( .A(n9338), .B(n23386), .Z(n51146) );
  XNOR U13341 ( .A(x[6196]), .B(y[6196]), .Z(n45670) );
  ANDN U13342 ( .B(y[6195]), .A(x[6195]), .Z(n45666) );
  XNOR U13343 ( .A(x[6194]), .B(y[6194]), .Z(n23390) );
  ANDN U13344 ( .B(y[6193]), .A(x[6193]), .Z(n58789) );
  ANDN U13345 ( .B(n23390), .A(n58789), .Z(n18794) );
  XNOR U13346 ( .A(x[6192]), .B(y[6192]), .Z(n45659) );
  XNOR U13347 ( .A(x[6190]), .B(y[6190]), .Z(n23392) );
  NANDN U13348 ( .A(y[6188]), .B(x[6188]), .Z(n9339) );
  NANDN U13349 ( .A(y[6189]), .B(x[6189]), .Z(n23391) );
  NAND U13350 ( .A(n9339), .B(n23391), .Z(n58783) );
  XNOR U13351 ( .A(x[6188]), .B(y[6188]), .Z(n45649) );
  ANDN U13352 ( .B(y[6187]), .A(x[6187]), .Z(n45645) );
  XNOR U13353 ( .A(x[6186]), .B(y[6186]), .Z(n23394) );
  ANDN U13354 ( .B(y[6185]), .A(x[6185]), .Z(n58779) );
  ANDN U13355 ( .B(n23394), .A(n58779), .Z(n18779) );
  XNOR U13356 ( .A(x[6184]), .B(y[6184]), .Z(n45638) );
  NANDN U13357 ( .A(y[6182]), .B(x[6182]), .Z(n9340) );
  NANDN U13358 ( .A(y[6183]), .B(x[6183]), .Z(n45637) );
  NAND U13359 ( .A(n9340), .B(n45637), .Z(n58776) );
  XNOR U13360 ( .A(x[6182]), .B(y[6182]), .Z(n23396) );
  NANDN U13361 ( .A(y[6180]), .B(x[6180]), .Z(n9341) );
  NANDN U13362 ( .A(y[6181]), .B(x[6181]), .Z(n23395) );
  NAND U13363 ( .A(n9341), .B(n23395), .Z(n58773) );
  XNOR U13364 ( .A(x[6180]), .B(y[6180]), .Z(n45628) );
  ANDN U13365 ( .B(y[6179]), .A(x[6179]), .Z(n45624) );
  NANDN U13366 ( .A(x[6177]), .B(y[6177]), .Z(n58770) );
  XNOR U13367 ( .A(x[6178]), .B(y[6178]), .Z(n23398) );
  NANDN U13368 ( .A(y[6176]), .B(x[6176]), .Z(n9342) );
  NANDN U13369 ( .A(y[6177]), .B(x[6177]), .Z(n23397) );
  NAND U13370 ( .A(n9342), .B(n23397), .Z(n58766) );
  XNOR U13371 ( .A(x[6176]), .B(y[6176]), .Z(n45617) );
  NANDN U13372 ( .A(x[6175]), .B(y[6175]), .Z(n51155) );
  XNOR U13373 ( .A(x[6174]), .B(y[6174]), .Z(n23400) );
  NANDN U13374 ( .A(y[6172]), .B(x[6172]), .Z(n9343) );
  NANDN U13375 ( .A(y[6173]), .B(x[6173]), .Z(n23399) );
  NAND U13376 ( .A(n9343), .B(n23399), .Z(n58760) );
  XNOR U13377 ( .A(x[6172]), .B(y[6172]), .Z(n23402) );
  ANDN U13378 ( .B(y[6171]), .A(x[6171]), .Z(n23403) );
  NANDN U13379 ( .A(x[6169]), .B(y[6169]), .Z(n58757) );
  XNOR U13380 ( .A(x[6170]), .B(y[6170]), .Z(n23405) );
  AND U13381 ( .A(n58757), .B(n23405), .Z(n18751) );
  NANDN U13382 ( .A(y[6166]), .B(x[6166]), .Z(n9344) );
  NANDN U13383 ( .A(y[6167]), .B(x[6167]), .Z(n23408) );
  NAND U13384 ( .A(n9344), .B(n23408), .Z(n51158) );
  XNOR U13385 ( .A(x[6166]), .B(y[6166]), .Z(n23411) );
  NANDN U13386 ( .A(x[6165]), .B(y[6165]), .Z(n58753) );
  AND U13387 ( .A(n23411), .B(n58753), .Z(n18746) );
  NANDN U13388 ( .A(y[6164]), .B(x[6164]), .Z(n23413) );
  NANDN U13389 ( .A(y[6165]), .B(x[6165]), .Z(n23410) );
  NAND U13390 ( .A(n23413), .B(n23410), .Z(n58752) );
  NANDN U13391 ( .A(x[6163]), .B(y[6163]), .Z(n45589) );
  NANDN U13392 ( .A(x[6164]), .B(y[6164]), .Z(n23412) );
  AND U13393 ( .A(n45589), .B(n23412), .Z(n58750) );
  XNOR U13394 ( .A(x[6162]), .B(y[6162]), .Z(n23416) );
  XNOR U13395 ( .A(x[6160]), .B(y[6160]), .Z(n45582) );
  NANDN U13396 ( .A(y[6158]), .B(x[6158]), .Z(n9345) );
  NANDN U13397 ( .A(y[6159]), .B(x[6159]), .Z(n45581) );
  NAND U13398 ( .A(n9345), .B(n45581), .Z(n58745) );
  XNOR U13399 ( .A(x[6158]), .B(y[6158]), .Z(n23418) );
  ANDN U13400 ( .B(y[6157]), .A(x[6157]), .Z(n58743) );
  NANDN U13401 ( .A(x[6155]), .B(y[6155]), .Z(n58742) );
  XNOR U13402 ( .A(x[6156]), .B(y[6156]), .Z(n45572) );
  AND U13403 ( .A(n58742), .B(n45572), .Z(n18729) );
  XNOR U13404 ( .A(x[6154]), .B(y[6154]), .Z(n23420) );
  NANDN U13405 ( .A(y[6152]), .B(x[6152]), .Z(n9346) );
  NANDN U13406 ( .A(y[6153]), .B(x[6153]), .Z(n23419) );
  NAND U13407 ( .A(n9346), .B(n23419), .Z(n58739) );
  XNOR U13408 ( .A(x[6152]), .B(y[6152]), .Z(n45562) );
  NANDN U13409 ( .A(y[6150]), .B(x[6150]), .Z(n9347) );
  NANDN U13410 ( .A(y[6151]), .B(x[6151]), .Z(n45561) );
  NAND U13411 ( .A(n9347), .B(n45561), .Z(n58735) );
  XNOR U13412 ( .A(x[6150]), .B(y[6150]), .Z(n23422) );
  ANDN U13413 ( .B(y[6149]), .A(x[6149]), .Z(n58733) );
  NANDN U13414 ( .A(x[6147]), .B(y[6147]), .Z(n58732) );
  XNOR U13415 ( .A(x[6148]), .B(y[6148]), .Z(n23424) );
  AND U13416 ( .A(n58732), .B(n23424), .Z(n18715) );
  XNOR U13417 ( .A(x[6144]), .B(y[6144]), .Z(n23430) );
  NANDN U13418 ( .A(y[6142]), .B(x[6142]), .Z(n9348) );
  NANDN U13419 ( .A(y[6143]), .B(x[6143]), .Z(n23429) );
  NAND U13420 ( .A(n9348), .B(n23429), .Z(n58727) );
  XNOR U13421 ( .A(x[6142]), .B(y[6142]), .Z(n23432) );
  ANDN U13422 ( .B(y[6141]), .A(x[6141]), .Z(n58724) );
  NANDN U13423 ( .A(y[6140]), .B(x[6140]), .Z(n9349) );
  NANDN U13424 ( .A(y[6141]), .B(x[6141]), .Z(n23431) );
  AND U13425 ( .A(n9349), .B(n23431), .Z(n58722) );
  XNOR U13426 ( .A(y[6140]), .B(x[6140]), .Z(n23434) );
  NANDN U13427 ( .A(x[6139]), .B(y[6139]), .Z(n23435) );
  AND U13428 ( .A(n23434), .B(n23435), .Z(n58721) );
  NANDN U13429 ( .A(y[6138]), .B(x[6138]), .Z(n9350) );
  NANDN U13430 ( .A(y[6139]), .B(x[6139]), .Z(n23433) );
  AND U13431 ( .A(n9350), .B(n23433), .Z(n58720) );
  ANDN U13432 ( .B(y[6137]), .A(x[6137]), .Z(n45529) );
  XNOR U13433 ( .A(x[6138]), .B(y[6138]), .Z(n23437) );
  NANDN U13434 ( .A(y[6136]), .B(x[6136]), .Z(n9351) );
  NANDN U13435 ( .A(y[6137]), .B(x[6137]), .Z(n23436) );
  NAND U13436 ( .A(n9351), .B(n23436), .Z(n58717) );
  XNOR U13437 ( .A(x[6136]), .B(y[6136]), .Z(n23439) );
  ANDN U13438 ( .B(y[6135]), .A(x[6135]), .Z(n45524) );
  NANDN U13439 ( .A(x[6133]), .B(y[6133]), .Z(n58714) );
  XNOR U13440 ( .A(x[6134]), .B(y[6134]), .Z(n23441) );
  AND U13441 ( .A(n58714), .B(n23441), .Z(n18694) );
  XNOR U13442 ( .A(x[6132]), .B(y[6132]), .Z(n23443) );
  NANDN U13443 ( .A(y[6130]), .B(x[6130]), .Z(n9352) );
  NANDN U13444 ( .A(y[6131]), .B(x[6131]), .Z(n23442) );
  NAND U13445 ( .A(n9352), .B(n23442), .Z(n58711) );
  XNOR U13446 ( .A(x[6130]), .B(y[6130]), .Z(n23445) );
  NANDN U13447 ( .A(y[6128]), .B(x[6128]), .Z(n9353) );
  NANDN U13448 ( .A(y[6129]), .B(x[6129]), .Z(n23444) );
  NAND U13449 ( .A(n9353), .B(n23444), .Z(n58707) );
  XNOR U13450 ( .A(x[6128]), .B(y[6128]), .Z(n23447) );
  ANDN U13451 ( .B(y[6127]), .A(x[6127]), .Z(n45507) );
  NANDN U13452 ( .A(x[6125]), .B(y[6125]), .Z(n58704) );
  XNOR U13453 ( .A(x[6126]), .B(y[6126]), .Z(n23449) );
  AND U13454 ( .A(n58704), .B(n23449), .Z(n18680) );
  NANDN U13455 ( .A(x[6123]), .B(y[6123]), .Z(n45497) );
  XOR U13456 ( .A(y[6124]), .B(x[6124]), .Z(n45500) );
  ANDN U13457 ( .B(n45497), .A(n45500), .Z(n58701) );
  XNOR U13458 ( .A(x[6122]), .B(y[6122]), .Z(n23451) );
  NANDN U13459 ( .A(y[6120]), .B(x[6120]), .Z(n9354) );
  NANDN U13460 ( .A(y[6121]), .B(x[6121]), .Z(n23450) );
  NAND U13461 ( .A(n9354), .B(n23450), .Z(n58697) );
  XNOR U13462 ( .A(x[6120]), .B(y[6120]), .Z(n23453) );
  NANDN U13463 ( .A(x[6119]), .B(y[6119]), .Z(n58696) );
  NANDN U13464 ( .A(y[6118]), .B(x[6118]), .Z(n9355) );
  NANDN U13465 ( .A(y[6119]), .B(x[6119]), .Z(n23452) );
  AND U13466 ( .A(n9355), .B(n23452), .Z(n58694) );
  NANDN U13467 ( .A(x[6117]), .B(y[6117]), .Z(n51171) );
  XNOR U13468 ( .A(x[6118]), .B(y[6118]), .Z(n23455) );
  AND U13469 ( .A(n51171), .B(n23455), .Z(n18667) );
  NANDN U13470 ( .A(y[6116]), .B(x[6116]), .Z(n9356) );
  NANDN U13471 ( .A(y[6117]), .B(x[6117]), .Z(n23454) );
  NAND U13472 ( .A(n9356), .B(n23454), .Z(n58693) );
  XNOR U13473 ( .A(x[6116]), .B(y[6116]), .Z(n23457) );
  XNOR U13474 ( .A(x[6114]), .B(y[6114]), .Z(n23459) );
  NANDN U13475 ( .A(y[6112]), .B(x[6112]), .Z(n9357) );
  NANDN U13476 ( .A(y[6113]), .B(x[6113]), .Z(n23458) );
  NAND U13477 ( .A(n9357), .B(n23458), .Z(n58686) );
  XNOR U13478 ( .A(x[6112]), .B(y[6112]), .Z(n23461) );
  NANDN U13479 ( .A(x[6111]), .B(y[6111]), .Z(n58685) );
  NANDN U13480 ( .A(y[6110]), .B(x[6110]), .Z(n9358) );
  NANDN U13481 ( .A(y[6111]), .B(x[6111]), .Z(n23460) );
  AND U13482 ( .A(n9358), .B(n23460), .Z(n58683) );
  XNOR U13483 ( .A(x[6110]), .B(y[6110]), .Z(n23463) );
  ANDN U13484 ( .B(y[6109]), .A(x[6109]), .Z(n45466) );
  ANDN U13485 ( .B(n23463), .A(n45466), .Z(n18654) );
  XNOR U13486 ( .A(x[6108]), .B(y[6108]), .Z(n23465) );
  NANDN U13487 ( .A(y[6106]), .B(x[6106]), .Z(n9359) );
  NANDN U13488 ( .A(y[6107]), .B(x[6107]), .Z(n23464) );
  NAND U13489 ( .A(n9359), .B(n23464), .Z(n51175) );
  XNOR U13490 ( .A(x[6106]), .B(y[6106]), .Z(n23467) );
  NANDN U13491 ( .A(y[6104]), .B(x[6104]), .Z(n9360) );
  NANDN U13492 ( .A(y[6105]), .B(x[6105]), .Z(n23466) );
  NAND U13493 ( .A(n9360), .B(n23466), .Z(n58677) );
  XNOR U13494 ( .A(x[6104]), .B(y[6104]), .Z(n23469) );
  NANDN U13495 ( .A(x[6103]), .B(y[6103]), .Z(n58674) );
  NANDN U13496 ( .A(y[6102]), .B(x[6102]), .Z(n9361) );
  NANDN U13497 ( .A(y[6103]), .B(x[6103]), .Z(n23468) );
  AND U13498 ( .A(n9361), .B(n23468), .Z(n58672) );
  NANDN U13499 ( .A(x[6101]), .B(y[6101]), .Z(n51176) );
  XNOR U13500 ( .A(x[6102]), .B(y[6102]), .Z(n23471) );
  AND U13501 ( .A(n51176), .B(n23471), .Z(n18641) );
  NANDN U13502 ( .A(y[6100]), .B(x[6100]), .Z(n9362) );
  NANDN U13503 ( .A(y[6101]), .B(x[6101]), .Z(n23470) );
  NAND U13504 ( .A(n9362), .B(n23470), .Z(n58671) );
  XNOR U13505 ( .A(x[6100]), .B(y[6100]), .Z(n23473) );
  NANDN U13506 ( .A(y[6098]), .B(x[6098]), .Z(n9363) );
  NANDN U13507 ( .A(y[6099]), .B(x[6099]), .Z(n23472) );
  NAND U13508 ( .A(n9363), .B(n23472), .Z(n58668) );
  XNOR U13509 ( .A(x[6098]), .B(y[6098]), .Z(n23475) );
  NANDN U13510 ( .A(y[6096]), .B(x[6096]), .Z(n9364) );
  NANDN U13511 ( .A(y[6097]), .B(x[6097]), .Z(n23474) );
  NAND U13512 ( .A(n9364), .B(n23474), .Z(n51178) );
  XNOR U13513 ( .A(x[6096]), .B(y[6096]), .Z(n45439) );
  NANDN U13514 ( .A(x[6095]), .B(y[6095]), .Z(n51179) );
  NANDN U13515 ( .A(y[6094]), .B(x[6094]), .Z(n9365) );
  ANDN U13516 ( .B(x[6095]), .A(y[6095]), .Z(n45438) );
  ANDN U13517 ( .B(n9365), .A(n45438), .Z(n58665) );
  NANDN U13518 ( .A(x[6093]), .B(y[6093]), .Z(n51181) );
  XNOR U13519 ( .A(x[6094]), .B(y[6094]), .Z(n23477) );
  AND U13520 ( .A(n51181), .B(n23477), .Z(n18629) );
  NANDN U13521 ( .A(y[6092]), .B(x[6092]), .Z(n9366) );
  NANDN U13522 ( .A(y[6093]), .B(x[6093]), .Z(n23476) );
  NAND U13523 ( .A(n9366), .B(n23476), .Z(n58664) );
  XNOR U13524 ( .A(x[6092]), .B(y[6092]), .Z(n23479) );
  NANDN U13525 ( .A(y[6090]), .B(x[6090]), .Z(n9367) );
  NANDN U13526 ( .A(y[6091]), .B(x[6091]), .Z(n23478) );
  NAND U13527 ( .A(n9367), .B(n23478), .Z(n58660) );
  XNOR U13528 ( .A(x[6090]), .B(y[6090]), .Z(n23481) );
  NANDN U13529 ( .A(y[6088]), .B(x[6088]), .Z(n9368) );
  NANDN U13530 ( .A(y[6089]), .B(x[6089]), .Z(n23480) );
  NAND U13531 ( .A(n9368), .B(n23480), .Z(n58657) );
  XNOR U13532 ( .A(x[6088]), .B(y[6088]), .Z(n23483) );
  NANDN U13533 ( .A(x[6087]), .B(y[6087]), .Z(n58656) );
  NANDN U13534 ( .A(y[6086]), .B(x[6086]), .Z(n9369) );
  NANDN U13535 ( .A(y[6087]), .B(x[6087]), .Z(n23482) );
  AND U13536 ( .A(n9369), .B(n23482), .Z(n58654) );
  NANDN U13537 ( .A(x[6085]), .B(y[6085]), .Z(n51183) );
  XNOR U13538 ( .A(x[6086]), .B(y[6086]), .Z(n23485) );
  AND U13539 ( .A(n51183), .B(n23485), .Z(n18617) );
  NANDN U13540 ( .A(y[6084]), .B(x[6084]), .Z(n9370) );
  NANDN U13541 ( .A(y[6085]), .B(x[6085]), .Z(n23484) );
  NAND U13542 ( .A(n9370), .B(n23484), .Z(n58653) );
  XNOR U13543 ( .A(x[6084]), .B(y[6084]), .Z(n23487) );
  NANDN U13544 ( .A(y[6082]), .B(x[6082]), .Z(n9371) );
  NANDN U13545 ( .A(y[6083]), .B(x[6083]), .Z(n23486) );
  NAND U13546 ( .A(n9371), .B(n23486), .Z(n58650) );
  XNOR U13547 ( .A(x[6082]), .B(y[6082]), .Z(n23489) );
  NANDN U13548 ( .A(y[6080]), .B(x[6080]), .Z(n9372) );
  NANDN U13549 ( .A(y[6081]), .B(x[6081]), .Z(n23488) );
  NAND U13550 ( .A(n9372), .B(n23488), .Z(n58647) );
  XNOR U13551 ( .A(x[6080]), .B(y[6080]), .Z(n23491) );
  NANDN U13552 ( .A(x[6079]), .B(y[6079]), .Z(n58644) );
  AND U13553 ( .A(n23491), .B(n58644), .Z(n18608) );
  NANDN U13554 ( .A(y[6076]), .B(x[6076]), .Z(n9373) );
  NANDN U13555 ( .A(y[6077]), .B(x[6077]), .Z(n23492) );
  AND U13556 ( .A(n9373), .B(n23492), .Z(n58640) );
  XNOR U13557 ( .A(x[6076]), .B(y[6076]), .Z(n23495) );
  XNOR U13558 ( .A(x[6074]), .B(y[6074]), .Z(n23498) );
  NANDN U13559 ( .A(y[6072]), .B(x[6072]), .Z(n9374) );
  NANDN U13560 ( .A(y[6073]), .B(x[6073]), .Z(n23497) );
  NAND U13561 ( .A(n9374), .B(n23497), .Z(n58634) );
  XNOR U13562 ( .A(x[6072]), .B(y[6072]), .Z(n23500) );
  NANDN U13563 ( .A(x[6071]), .B(y[6071]), .Z(n58633) );
  NANDN U13564 ( .A(y[6070]), .B(x[6070]), .Z(n9375) );
  NANDN U13565 ( .A(y[6071]), .B(x[6071]), .Z(n23499) );
  AND U13566 ( .A(n9375), .B(n23499), .Z(n58631) );
  XNOR U13567 ( .A(x[6070]), .B(y[6070]), .Z(n23502) );
  ANDN U13568 ( .B(y[6069]), .A(x[6069]), .Z(n23503) );
  ANDN U13569 ( .B(n23502), .A(n23503), .Z(n18591) );
  NANDN U13570 ( .A(x[6067]), .B(y[6067]), .Z(n23507) );
  NANDN U13571 ( .A(x[6068]), .B(y[6068]), .Z(n23504) );
  AND U13572 ( .A(n23507), .B(n23504), .Z(n58629) );
  NANDN U13573 ( .A(y[6066]), .B(x[6066]), .Z(n23509) );
  NANDN U13574 ( .A(y[6067]), .B(x[6067]), .Z(n23506) );
  NAND U13575 ( .A(n23509), .B(n23506), .Z(n58628) );
  NANDN U13576 ( .A(x[6065]), .B(y[6065]), .Z(n45375) );
  NANDN U13577 ( .A(x[6066]), .B(y[6066]), .Z(n23508) );
  AND U13578 ( .A(n45375), .B(n23508), .Z(n58627) );
  NANDN U13579 ( .A(y[6064]), .B(x[6064]), .Z(n9376) );
  NANDN U13580 ( .A(y[6065]), .B(x[6065]), .Z(n23510) );
  NAND U13581 ( .A(n9376), .B(n23510), .Z(n58625) );
  XNOR U13582 ( .A(x[6064]), .B(y[6064]), .Z(n23512) );
  NANDN U13583 ( .A(x[6063]), .B(y[6063]), .Z(n51189) );
  AND U13584 ( .A(n23512), .B(n51189), .Z(n18584) );
  NANDN U13585 ( .A(x[6061]), .B(y[6061]), .Z(n23516) );
  NANDN U13586 ( .A(x[6062]), .B(y[6062]), .Z(n23513) );
  AND U13587 ( .A(n23516), .B(n23513), .Z(n58623) );
  NANDN U13588 ( .A(y[6060]), .B(x[6060]), .Z(n23518) );
  NANDN U13589 ( .A(y[6061]), .B(x[6061]), .Z(n23515) );
  NAND U13590 ( .A(n23518), .B(n23515), .Z(n58622) );
  NANDN U13591 ( .A(x[6059]), .B(y[6059]), .Z(n45363) );
  NANDN U13592 ( .A(x[6060]), .B(y[6060]), .Z(n23517) );
  AND U13593 ( .A(n45363), .B(n23517), .Z(n58621) );
  NANDN U13594 ( .A(y[6058]), .B(x[6058]), .Z(n9377) );
  NANDN U13595 ( .A(y[6059]), .B(x[6059]), .Z(n23519) );
  NAND U13596 ( .A(n9377), .B(n23519), .Z(n58620) );
  XNOR U13597 ( .A(x[6058]), .B(y[6058]), .Z(n23521) );
  NANDN U13598 ( .A(x[6057]), .B(y[6057]), .Z(n51191) );
  AND U13599 ( .A(n23521), .B(n51191), .Z(n18577) );
  NANDN U13600 ( .A(y[6056]), .B(x[6056]), .Z(n9378) );
  NANDN U13601 ( .A(y[6057]), .B(x[6057]), .Z(n23520) );
  NAND U13602 ( .A(n9378), .B(n23520), .Z(n58619) );
  XNOR U13603 ( .A(x[6056]), .B(y[6056]), .Z(n23523) );
  NANDN U13604 ( .A(x[6055]), .B(y[6055]), .Z(n58617) );
  NANDN U13605 ( .A(y[6054]), .B(x[6054]), .Z(n23525) );
  NANDN U13606 ( .A(y[6055]), .B(x[6055]), .Z(n23522) );
  NAND U13607 ( .A(n23525), .B(n23522), .Z(n58616) );
  NANDN U13608 ( .A(y[6052]), .B(x[6052]), .Z(n23529) );
  NANDN U13609 ( .A(y[6053]), .B(x[6053]), .Z(n23526) );
  AND U13610 ( .A(n23529), .B(n23526), .Z(n58614) );
  NANDN U13611 ( .A(x[6051]), .B(y[6051]), .Z(n23531) );
  NANDN U13612 ( .A(x[6052]), .B(y[6052]), .Z(n23528) );
  NAND U13613 ( .A(n23531), .B(n23528), .Z(n58613) );
  NANDN U13614 ( .A(y[6050]), .B(x[6050]), .Z(n23533) );
  NANDN U13615 ( .A(y[6051]), .B(x[6051]), .Z(n23530) );
  AND U13616 ( .A(n23533), .B(n23530), .Z(n58612) );
  NANDN U13617 ( .A(x[6049]), .B(y[6049]), .Z(n45341) );
  NANDN U13618 ( .A(x[6050]), .B(y[6050]), .Z(n23532) );
  NAND U13619 ( .A(n45341), .B(n23532), .Z(n58610) );
  NANDN U13620 ( .A(y[6048]), .B(x[6048]), .Z(n9379) );
  NANDN U13621 ( .A(y[6049]), .B(x[6049]), .Z(n23534) );
  AND U13622 ( .A(n9379), .B(n23534), .Z(n58609) );
  NANDN U13623 ( .A(y[6046]), .B(x[6046]), .Z(n9380) );
  NANDN U13624 ( .A(y[6047]), .B(x[6047]), .Z(n23535) );
  AND U13625 ( .A(n9380), .B(n23535), .Z(n58606) );
  NANDN U13626 ( .A(x[6045]), .B(y[6045]), .Z(n51193) );
  XNOR U13627 ( .A(x[6046]), .B(y[6046]), .Z(n23538) );
  AND U13628 ( .A(n51193), .B(n23538), .Z(n18562) );
  NANDN U13629 ( .A(y[6044]), .B(x[6044]), .Z(n9381) );
  NANDN U13630 ( .A(y[6045]), .B(x[6045]), .Z(n23537) );
  NAND U13631 ( .A(n9381), .B(n23537), .Z(n58605) );
  XNOR U13632 ( .A(x[6044]), .B(y[6044]), .Z(n23540) );
  NANDN U13633 ( .A(y[6042]), .B(x[6042]), .Z(n9382) );
  NANDN U13634 ( .A(y[6043]), .B(x[6043]), .Z(n23539) );
  NAND U13635 ( .A(n9382), .B(n23539), .Z(n58602) );
  XNOR U13636 ( .A(x[6042]), .B(y[6042]), .Z(n23542) );
  NANDN U13637 ( .A(y[6040]), .B(x[6040]), .Z(n9383) );
  NANDN U13638 ( .A(y[6041]), .B(x[6041]), .Z(n23541) );
  NAND U13639 ( .A(n9383), .B(n23541), .Z(n58599) );
  XNOR U13640 ( .A(x[6040]), .B(y[6040]), .Z(n45322) );
  NANDN U13641 ( .A(x[6039]), .B(y[6039]), .Z(n58598) );
  NANDN U13642 ( .A(y[6038]), .B(x[6038]), .Z(n9384) );
  NANDN U13643 ( .A(y[6039]), .B(x[6039]), .Z(n45323) );
  AND U13644 ( .A(n9384), .B(n45323), .Z(n58596) );
  XNOR U13645 ( .A(y[6038]), .B(x[6038]), .Z(n45316) );
  NANDN U13646 ( .A(x[6037]), .B(y[6037]), .Z(n45312) );
  NAND U13647 ( .A(n45316), .B(n45312), .Z(n58595) );
  NANDN U13648 ( .A(y[6036]), .B(x[6036]), .Z(n9385) );
  NANDN U13649 ( .A(y[6037]), .B(x[6037]), .Z(n45315) );
  AND U13650 ( .A(n9385), .B(n45315), .Z(n58594) );
  ANDN U13651 ( .B(y[6035]), .A(x[6035]), .Z(n23546) );
  XNOR U13652 ( .A(x[6036]), .B(y[6036]), .Z(n23545) );
  NANDN U13653 ( .A(y[6034]), .B(x[6034]), .Z(n9386) );
  NANDN U13654 ( .A(y[6035]), .B(x[6035]), .Z(n23544) );
  NAND U13655 ( .A(n9386), .B(n23544), .Z(n58591) );
  XNOR U13656 ( .A(x[6034]), .B(y[6034]), .Z(n23548) );
  NANDN U13657 ( .A(x[6033]), .B(y[6033]), .Z(n58590) );
  NANDN U13658 ( .A(y[6032]), .B(x[6032]), .Z(n9387) );
  NANDN U13659 ( .A(y[6033]), .B(x[6033]), .Z(n23547) );
  AND U13660 ( .A(n9387), .B(n23547), .Z(n58588) );
  XNOR U13661 ( .A(x[6032]), .B(y[6032]), .Z(n45302) );
  XNOR U13662 ( .A(x[6030]), .B(y[6030]), .Z(n23550) );
  NANDN U13663 ( .A(x[6029]), .B(y[6029]), .Z(n58585) );
  AND U13664 ( .A(n23550), .B(n58585), .Z(n18538) );
  XNOR U13665 ( .A(x[6028]), .B(y[6028]), .Z(n23552) );
  XNOR U13666 ( .A(x[6026]), .B(y[6026]), .Z(n23554) );
  NANDN U13667 ( .A(y[6024]), .B(x[6024]), .Z(n9388) );
  NANDN U13668 ( .A(y[6025]), .B(x[6025]), .Z(n23553) );
  NAND U13669 ( .A(n9388), .B(n23553), .Z(n58575) );
  XNOR U13670 ( .A(x[6024]), .B(y[6024]), .Z(n23556) );
  NANDN U13671 ( .A(x[6023]), .B(y[6023]), .Z(n51198) );
  AND U13672 ( .A(n23556), .B(n51198), .Z(n18527) );
  XNOR U13673 ( .A(y[6022]), .B(x[6022]), .Z(n23559) );
  NANDN U13674 ( .A(x[6021]), .B(y[6021]), .Z(n45277) );
  AND U13675 ( .A(n23559), .B(n45277), .Z(n58573) );
  XNOR U13676 ( .A(x[6020]), .B(y[6020]), .Z(n45275) );
  XNOR U13677 ( .A(x[6018]), .B(y[6018]), .Z(n23561) );
  NANDN U13678 ( .A(y[6016]), .B(x[6016]), .Z(n9389) );
  NANDN U13679 ( .A(y[6017]), .B(x[6017]), .Z(n23560) );
  NAND U13680 ( .A(n9389), .B(n23560), .Z(n58568) );
  XNOR U13681 ( .A(x[6016]), .B(y[6016]), .Z(n23563) );
  ANDN U13682 ( .B(y[6015]), .A(x[6015]), .Z(n45262) );
  XNOR U13683 ( .A(x[6014]), .B(y[6014]), .Z(n23565) );
  ANDN U13684 ( .B(y[6013]), .A(x[6013]), .Z(n45257) );
  ANDN U13685 ( .B(n23565), .A(n45257), .Z(n18509) );
  XNOR U13686 ( .A(x[6012]), .B(y[6012]), .Z(n23567) );
  XNOR U13687 ( .A(x[6010]), .B(y[6010]), .Z(n23569) );
  NANDN U13688 ( .A(y[6008]), .B(x[6008]), .Z(n9390) );
  NANDN U13689 ( .A(y[6009]), .B(x[6009]), .Z(n23568) );
  NAND U13690 ( .A(n9390), .B(n23568), .Z(n58558) );
  XNOR U13691 ( .A(x[6008]), .B(y[6008]), .Z(n23571) );
  ANDN U13692 ( .B(y[6007]), .A(x[6007]), .Z(n45244) );
  XNOR U13693 ( .A(x[6006]), .B(y[6006]), .Z(n23573) );
  ANDN U13694 ( .B(y[6005]), .A(x[6005]), .Z(n45239) );
  ANDN U13695 ( .B(n23573), .A(n45239), .Z(n18494) );
  XNOR U13696 ( .A(x[6004]), .B(y[6004]), .Z(n23575) );
  XNOR U13697 ( .A(x[6002]), .B(y[6002]), .Z(n23577) );
  NANDN U13698 ( .A(y[6000]), .B(x[6000]), .Z(n9391) );
  NANDN U13699 ( .A(y[6001]), .B(x[6001]), .Z(n23576) );
  NAND U13700 ( .A(n9391), .B(n23576), .Z(n58547) );
  XNOR U13701 ( .A(x[6000]), .B(y[6000]), .Z(n23579) );
  ANDN U13702 ( .B(y[5999]), .A(x[5999]), .Z(n45226) );
  XNOR U13703 ( .A(x[5998]), .B(y[5998]), .Z(n23581) );
  NANDN U13704 ( .A(y[5996]), .B(x[5996]), .Z(n9392) );
  NANDN U13705 ( .A(y[5997]), .B(x[5997]), .Z(n23580) );
  AND U13706 ( .A(n9392), .B(n23580), .Z(n51208) );
  NANDN U13707 ( .A(x[5995]), .B(y[5995]), .Z(n58540) );
  XNOR U13708 ( .A(x[5996]), .B(y[5996]), .Z(n23583) );
  XNOR U13709 ( .A(x[5994]), .B(y[5994]), .Z(n23585) );
  NANDN U13710 ( .A(y[5992]), .B(x[5992]), .Z(n9393) );
  NANDN U13711 ( .A(y[5993]), .B(x[5993]), .Z(n23584) );
  NAND U13712 ( .A(n9393), .B(n23584), .Z(n58537) );
  XNOR U13713 ( .A(x[5992]), .B(y[5992]), .Z(n23587) );
  ANDN U13714 ( .B(y[5991]), .A(x[5991]), .Z(n23588) );
  XNOR U13715 ( .A(x[5990]), .B(y[5990]), .Z(n23590) );
  ANDN U13716 ( .B(y[5989]), .A(x[5989]), .Z(n45204) );
  ANDN U13717 ( .B(n23590), .A(n45204), .Z(n18465) );
  XNOR U13718 ( .A(x[5988]), .B(y[5988]), .Z(n23592) );
  XNOR U13719 ( .A(x[5986]), .B(y[5986]), .Z(n23594) );
  NANDN U13720 ( .A(y[5984]), .B(x[5984]), .Z(n9394) );
  NANDN U13721 ( .A(y[5985]), .B(x[5985]), .Z(n23593) );
  NAND U13722 ( .A(n9394), .B(n23593), .Z(n58528) );
  XNOR U13723 ( .A(x[5984]), .B(y[5984]), .Z(n23596) );
  ANDN U13724 ( .B(y[5983]), .A(x[5983]), .Z(n58525) );
  ANDN U13725 ( .B(y[5981]), .A(x[5981]), .Z(n45187) );
  NANDN U13726 ( .A(y[5980]), .B(x[5980]), .Z(n9395) );
  NANDN U13727 ( .A(y[5981]), .B(x[5981]), .Z(n23597) );
  AND U13728 ( .A(n9395), .B(n23597), .Z(n51214) );
  XNOR U13729 ( .A(x[5980]), .B(y[5980]), .Z(n23600) );
  XNOR U13730 ( .A(x[5978]), .B(y[5978]), .Z(n23602) );
  NANDN U13731 ( .A(y[5976]), .B(x[5976]), .Z(n9396) );
  NANDN U13732 ( .A(y[5977]), .B(x[5977]), .Z(n23601) );
  NAND U13733 ( .A(n9396), .B(n23601), .Z(n58516) );
  XNOR U13734 ( .A(x[5976]), .B(y[5976]), .Z(n23604) );
  ANDN U13735 ( .B(y[5975]), .A(x[5975]), .Z(n23605) );
  NANDN U13736 ( .A(x[5973]), .B(y[5973]), .Z(n58511) );
  XNOR U13737 ( .A(x[5974]), .B(y[5974]), .Z(n23607) );
  AND U13738 ( .A(n58511), .B(n23607), .Z(n18436) );
  NANDN U13739 ( .A(y[5972]), .B(x[5972]), .Z(n9397) );
  NANDN U13740 ( .A(y[5973]), .B(x[5973]), .Z(n23606) );
  NAND U13741 ( .A(n9397), .B(n23606), .Z(n58510) );
  XNOR U13742 ( .A(x[5972]), .B(y[5972]), .Z(n23609) );
  XNOR U13743 ( .A(x[5970]), .B(y[5970]), .Z(n23611) );
  ANDN U13744 ( .B(x[5968]), .A(y[5968]), .Z(n45160) );
  NANDN U13745 ( .A(y[5969]), .B(x[5969]), .Z(n23610) );
  NANDN U13746 ( .A(n45160), .B(n23610), .Z(n58503) );
  NANDN U13747 ( .A(x[5967]), .B(y[5967]), .Z(n23613) );
  NANDN U13748 ( .A(x[5968]), .B(y[5968]), .Z(n23612) );
  AND U13749 ( .A(n23613), .B(n23612), .Z(n58502) );
  NANDN U13750 ( .A(y[5966]), .B(x[5966]), .Z(n23615) );
  NANDN U13751 ( .A(y[5967]), .B(x[5967]), .Z(n45161) );
  NAND U13752 ( .A(n23615), .B(n45161), .Z(n58501) );
  NANDN U13753 ( .A(x[5965]), .B(y[5965]), .Z(n45152) );
  NANDN U13754 ( .A(x[5966]), .B(y[5966]), .Z(n23614) );
  AND U13755 ( .A(n45152), .B(n23614), .Z(n58500) );
  NANDN U13756 ( .A(y[5964]), .B(x[5964]), .Z(n9398) );
  NANDN U13757 ( .A(y[5965]), .B(x[5965]), .Z(n23616) );
  NAND U13758 ( .A(n9398), .B(n23616), .Z(n58499) );
  XNOR U13759 ( .A(x[5964]), .B(y[5964]), .Z(n23618) );
  NANDN U13760 ( .A(y[5962]), .B(x[5962]), .Z(n9399) );
  NANDN U13761 ( .A(y[5963]), .B(x[5963]), .Z(n23617) );
  NAND U13762 ( .A(n9399), .B(n23617), .Z(n58498) );
  XNOR U13763 ( .A(x[5962]), .B(y[5962]), .Z(n23620) );
  ANDN U13764 ( .B(y[5961]), .A(x[5961]), .Z(n23621) );
  NANDN U13765 ( .A(x[5959]), .B(y[5959]), .Z(n45140) );
  NANDN U13766 ( .A(x[5960]), .B(y[5960]), .Z(n23622) );
  AND U13767 ( .A(n45140), .B(n23622), .Z(n58495) );
  XNOR U13768 ( .A(x[5958]), .B(y[5958]), .Z(n23626) );
  XNOR U13769 ( .A(x[5956]), .B(y[5956]), .Z(n45133) );
  ANDN U13770 ( .B(x[5955]), .A(y[5955]), .Z(n45132) );
  NANDN U13771 ( .A(y[5954]), .B(x[5954]), .Z(n23628) );
  NANDN U13772 ( .A(n45132), .B(n23628), .Z(n58489) );
  NANDN U13773 ( .A(x[5953]), .B(y[5953]), .Z(n45124) );
  NANDN U13774 ( .A(x[5954]), .B(y[5954]), .Z(n23627) );
  AND U13775 ( .A(n45124), .B(n23627), .Z(n58488) );
  NANDN U13776 ( .A(y[5952]), .B(x[5952]), .Z(n9400) );
  NANDN U13777 ( .A(y[5953]), .B(x[5953]), .Z(n23629) );
  NAND U13778 ( .A(n9400), .B(n23629), .Z(n58487) );
  NANDN U13779 ( .A(y[5950]), .B(x[5950]), .Z(n9401) );
  NANDN U13780 ( .A(y[5951]), .B(x[5951]), .Z(n45120) );
  AND U13781 ( .A(n9401), .B(n45120), .Z(n58486) );
  XNOR U13782 ( .A(x[5950]), .B(y[5950]), .Z(n23631) );
  NANDN U13783 ( .A(y[5948]), .B(x[5948]), .Z(n9402) );
  NANDN U13784 ( .A(y[5949]), .B(x[5949]), .Z(n23630) );
  AND U13785 ( .A(n9402), .B(n23630), .Z(n58483) );
  ANDN U13786 ( .B(y[5947]), .A(x[5947]), .Z(n45108) );
  XNOR U13787 ( .A(x[5948]), .B(y[5948]), .Z(n23633) );
  NANDN U13788 ( .A(y[5946]), .B(x[5946]), .Z(n9403) );
  NANDN U13789 ( .A(y[5947]), .B(x[5947]), .Z(n23632) );
  NAND U13790 ( .A(n9403), .B(n23632), .Z(n58480) );
  XNOR U13791 ( .A(x[5946]), .B(y[5946]), .Z(n23635) );
  NANDN U13792 ( .A(x[5945]), .B(y[5945]), .Z(n58477) );
  AND U13793 ( .A(n23635), .B(n58477), .Z(n18395) );
  NANDN U13794 ( .A(y[5942]), .B(x[5942]), .Z(n9404) );
  NANDN U13795 ( .A(y[5943]), .B(x[5943]), .Z(n23636) );
  AND U13796 ( .A(n9404), .B(n23636), .Z(n58473) );
  XNOR U13797 ( .A(x[5942]), .B(y[5942]), .Z(n23639) );
  XNOR U13798 ( .A(x[5940]), .B(y[5940]), .Z(n23641) );
  NANDN U13799 ( .A(y[5938]), .B(x[5938]), .Z(n9405) );
  NANDN U13800 ( .A(y[5939]), .B(x[5939]), .Z(n23640) );
  NAND U13801 ( .A(n9405), .B(n23640), .Z(n58467) );
  XNOR U13802 ( .A(x[5938]), .B(y[5938]), .Z(n23643) );
  NANDN U13803 ( .A(x[5937]), .B(y[5937]), .Z(n58466) );
  AND U13804 ( .A(n23643), .B(n58466), .Z(n18381) );
  XNOR U13805 ( .A(x[5934]), .B(y[5934]), .Z(n23647) );
  XNOR U13806 ( .A(x[5932]), .B(y[5932]), .Z(n45074) );
  ANDN U13807 ( .B(x[5931]), .A(y[5931]), .Z(n45073) );
  NANDN U13808 ( .A(y[5930]), .B(x[5930]), .Z(n9406) );
  NANDN U13809 ( .A(n45073), .B(n9406), .Z(n58458) );
  XNOR U13810 ( .A(x[5930]), .B(y[5930]), .Z(n23649) );
  ANDN U13811 ( .B(y[5929]), .A(x[5929]), .Z(n45066) );
  NANDN U13812 ( .A(y[5928]), .B(x[5928]), .Z(n9407) );
  NANDN U13813 ( .A(y[5929]), .B(x[5929]), .Z(n23648) );
  AND U13814 ( .A(n9407), .B(n23648), .Z(n58457) );
  XNOR U13815 ( .A(x[5928]), .B(y[5928]), .Z(n23651) );
  NANDN U13816 ( .A(x[5927]), .B(y[5927]), .Z(n58455) );
  AND U13817 ( .A(n23651), .B(n58455), .Z(n18364) );
  NANDN U13818 ( .A(x[5925]), .B(y[5925]), .Z(n58452) );
  XNOR U13819 ( .A(x[5926]), .B(y[5926]), .Z(n23653) );
  AND U13820 ( .A(n58452), .B(n23653), .Z(n18360) );
  NANDN U13821 ( .A(y[5924]), .B(x[5924]), .Z(n9408) );
  NANDN U13822 ( .A(y[5925]), .B(x[5925]), .Z(n23652) );
  NAND U13823 ( .A(n9408), .B(n23652), .Z(n58451) );
  XNOR U13824 ( .A(x[5924]), .B(y[5924]), .Z(n23654) );
  NANDN U13825 ( .A(y[5922]), .B(x[5922]), .Z(n23657) );
  NANDN U13826 ( .A(y[5923]), .B(x[5923]), .Z(n23655) );
  AND U13827 ( .A(n23657), .B(n23655), .Z(n58447) );
  NANDN U13828 ( .A(x[5921]), .B(y[5921]), .Z(n45049) );
  NANDN U13829 ( .A(x[5922]), .B(y[5922]), .Z(n23656) );
  AND U13830 ( .A(n45049), .B(n23656), .Z(n51233) );
  XNOR U13831 ( .A(x[5918]), .B(y[5918]), .Z(n23662) );
  NANDN U13832 ( .A(y[5916]), .B(x[5916]), .Z(n9409) );
  NANDN U13833 ( .A(y[5917]), .B(x[5917]), .Z(n23661) );
  NAND U13834 ( .A(n9409), .B(n23661), .Z(n58442) );
  XNOR U13835 ( .A(x[5916]), .B(y[5916]), .Z(n23664) );
  NANDN U13836 ( .A(y[5914]), .B(x[5914]), .Z(n9410) );
  NANDN U13837 ( .A(y[5915]), .B(x[5915]), .Z(n23663) );
  NAND U13838 ( .A(n9410), .B(n23663), .Z(n58441) );
  XNOR U13839 ( .A(x[5914]), .B(y[5914]), .Z(n23666) );
  ANDN U13840 ( .B(y[5913]), .A(x[5913]), .Z(n45030) );
  NANDN U13841 ( .A(x[5911]), .B(y[5911]), .Z(n58434) );
  XNOR U13842 ( .A(x[5912]), .B(y[5912]), .Z(n23668) );
  AND U13843 ( .A(n58434), .B(n23668), .Z(n18338) );
  NANDN U13844 ( .A(y[5910]), .B(x[5910]), .Z(n9411) );
  NANDN U13845 ( .A(y[5911]), .B(x[5911]), .Z(n23667) );
  NAND U13846 ( .A(n9411), .B(n23667), .Z(n58433) );
  XNOR U13847 ( .A(x[5910]), .B(y[5910]), .Z(n23670) );
  NANDN U13848 ( .A(y[5908]), .B(x[5908]), .Z(n9412) );
  NANDN U13849 ( .A(y[5909]), .B(x[5909]), .Z(n23669) );
  NAND U13850 ( .A(n9412), .B(n23669), .Z(n58430) );
  XNOR U13851 ( .A(x[5908]), .B(y[5908]), .Z(n23672) );
  NANDN U13852 ( .A(y[5906]), .B(x[5906]), .Z(n9413) );
  NANDN U13853 ( .A(y[5907]), .B(x[5907]), .Z(n23671) );
  NAND U13854 ( .A(n9413), .B(n23671), .Z(n58429) );
  XNOR U13855 ( .A(x[5906]), .B(y[5906]), .Z(n23674) );
  ANDN U13856 ( .B(y[5905]), .A(x[5905]), .Z(n45013) );
  NANDN U13857 ( .A(x[5903]), .B(y[5903]), .Z(n58424) );
  XNOR U13858 ( .A(x[5904]), .B(y[5904]), .Z(n23676) );
  AND U13859 ( .A(n58424), .B(n23676), .Z(n18325) );
  NANDN U13860 ( .A(y[5902]), .B(x[5902]), .Z(n9414) );
  NANDN U13861 ( .A(y[5903]), .B(x[5903]), .Z(n23675) );
  NAND U13862 ( .A(n9414), .B(n23675), .Z(n58423) );
  XNOR U13863 ( .A(x[5902]), .B(y[5902]), .Z(n23678) );
  NANDN U13864 ( .A(y[5900]), .B(x[5900]), .Z(n9415) );
  NANDN U13865 ( .A(y[5901]), .B(x[5901]), .Z(n23677) );
  NAND U13866 ( .A(n9415), .B(n23677), .Z(n58417) );
  XNOR U13867 ( .A(x[5900]), .B(y[5900]), .Z(n23680) );
  NANDN U13868 ( .A(y[5898]), .B(x[5898]), .Z(n9416) );
  NANDN U13869 ( .A(y[5899]), .B(x[5899]), .Z(n23679) );
  NAND U13870 ( .A(n9416), .B(n23679), .Z(n58416) );
  XNOR U13871 ( .A(x[5898]), .B(y[5898]), .Z(n23682) );
  ANDN U13872 ( .B(y[5897]), .A(x[5897]), .Z(n44996) );
  NANDN U13873 ( .A(x[5895]), .B(y[5895]), .Z(n58411) );
  XNOR U13874 ( .A(x[5896]), .B(y[5896]), .Z(n23684) );
  AND U13875 ( .A(n58411), .B(n23684), .Z(n18312) );
  NANDN U13876 ( .A(y[5894]), .B(x[5894]), .Z(n9417) );
  NANDN U13877 ( .A(y[5895]), .B(x[5895]), .Z(n23683) );
  NAND U13878 ( .A(n9417), .B(n23683), .Z(n58410) );
  XNOR U13879 ( .A(x[5894]), .B(y[5894]), .Z(n23686) );
  NANDN U13880 ( .A(y[5892]), .B(x[5892]), .Z(n9418) );
  NANDN U13881 ( .A(y[5893]), .B(x[5893]), .Z(n23685) );
  NAND U13882 ( .A(n9418), .B(n23685), .Z(n58407) );
  XNOR U13883 ( .A(x[5892]), .B(y[5892]), .Z(n23688) );
  NANDN U13884 ( .A(y[5890]), .B(x[5890]), .Z(n9419) );
  NANDN U13885 ( .A(y[5891]), .B(x[5891]), .Z(n23687) );
  NAND U13886 ( .A(n9419), .B(n23687), .Z(n58406) );
  XNOR U13887 ( .A(x[5890]), .B(y[5890]), .Z(n23690) );
  ANDN U13888 ( .B(y[5889]), .A(x[5889]), .Z(n44979) );
  NANDN U13889 ( .A(x[5887]), .B(y[5887]), .Z(n58400) );
  XNOR U13890 ( .A(x[5888]), .B(y[5888]), .Z(n23692) );
  AND U13891 ( .A(n58400), .B(n23692), .Z(n18299) );
  NANDN U13892 ( .A(y[5886]), .B(x[5886]), .Z(n9420) );
  NANDN U13893 ( .A(y[5887]), .B(x[5887]), .Z(n23691) );
  NAND U13894 ( .A(n9420), .B(n23691), .Z(n58399) );
  XNOR U13895 ( .A(x[5886]), .B(y[5886]), .Z(n23694) );
  NANDN U13896 ( .A(y[5884]), .B(x[5884]), .Z(n9421) );
  NANDN U13897 ( .A(y[5885]), .B(x[5885]), .Z(n23693) );
  NAND U13898 ( .A(n9421), .B(n23693), .Z(n58396) );
  XNOR U13899 ( .A(x[5884]), .B(y[5884]), .Z(n23696) );
  NANDN U13900 ( .A(y[5882]), .B(x[5882]), .Z(n9422) );
  NANDN U13901 ( .A(y[5883]), .B(x[5883]), .Z(n23695) );
  NAND U13902 ( .A(n9422), .B(n23695), .Z(n58395) );
  XNOR U13903 ( .A(x[5882]), .B(y[5882]), .Z(n23698) );
  ANDN U13904 ( .B(y[5881]), .A(x[5881]), .Z(n44962) );
  XNOR U13905 ( .A(x[5880]), .B(y[5880]), .Z(n23700) );
  ANDN U13906 ( .B(y[5879]), .A(x[5879]), .Z(n58390) );
  ANDN U13907 ( .B(n23700), .A(n58390), .Z(n18286) );
  NANDN U13908 ( .A(y[5878]), .B(x[5878]), .Z(n9423) );
  NANDN U13909 ( .A(y[5879]), .B(x[5879]), .Z(n23699) );
  NAND U13910 ( .A(n9423), .B(n23699), .Z(n58389) );
  XNOR U13911 ( .A(x[5878]), .B(y[5878]), .Z(n44955) );
  NANDN U13912 ( .A(y[5876]), .B(x[5876]), .Z(n9424) );
  NANDN U13913 ( .A(y[5877]), .B(x[5877]), .Z(n44954) );
  NAND U13914 ( .A(n9424), .B(n44954), .Z(n58385) );
  NANDN U13915 ( .A(x[5875]), .B(y[5875]), .Z(n51245) );
  XNOR U13916 ( .A(x[5876]), .B(y[5876]), .Z(n23702) );
  NANDN U13917 ( .A(y[5874]), .B(x[5874]), .Z(n9425) );
  NANDN U13918 ( .A(y[5875]), .B(x[5875]), .Z(n23701) );
  NAND U13919 ( .A(n9425), .B(n23701), .Z(n58384) );
  XNOR U13920 ( .A(x[5874]), .B(y[5874]), .Z(n23704) );
  ANDN U13921 ( .B(y[5873]), .A(x[5873]), .Z(n23705) );
  NANDN U13922 ( .A(x[5871]), .B(y[5871]), .Z(n44940) );
  NANDN U13923 ( .A(x[5872]), .B(y[5872]), .Z(n23706) );
  NAND U13924 ( .A(n44940), .B(n23706), .Z(n51248) );
  NANDN U13925 ( .A(y[5870]), .B(x[5870]), .Z(n9426) );
  NANDN U13926 ( .A(y[5871]), .B(x[5871]), .Z(n23708) );
  AND U13927 ( .A(n9426), .B(n23708), .Z(n58381) );
  ANDN U13928 ( .B(y[5869]), .A(x[5869]), .Z(n44934) );
  XNOR U13929 ( .A(x[5870]), .B(y[5870]), .Z(n23710) );
  NANDN U13930 ( .A(y[5868]), .B(x[5868]), .Z(n9427) );
  NANDN U13931 ( .A(y[5869]), .B(x[5869]), .Z(n23709) );
  NAND U13932 ( .A(n9427), .B(n23709), .Z(n58379) );
  XNOR U13933 ( .A(x[5868]), .B(y[5868]), .Z(n23712) );
  ANDN U13934 ( .B(y[5867]), .A(x[5867]), .Z(n23713) );
  NANDN U13935 ( .A(x[5865]), .B(y[5865]), .Z(n44925) );
  NANDN U13936 ( .A(x[5866]), .B(y[5866]), .Z(n23714) );
  AND U13937 ( .A(n44925), .B(n23714), .Z(n58376) );
  XNOR U13938 ( .A(x[5864]), .B(y[5864]), .Z(n23718) );
  XNOR U13939 ( .A(x[5862]), .B(y[5862]), .Z(n23720) );
  NANDN U13940 ( .A(y[5860]), .B(x[5860]), .Z(n23723) );
  NANDN U13941 ( .A(y[5861]), .B(x[5861]), .Z(n23719) );
  NAND U13942 ( .A(n23723), .B(n23719), .Z(n58370) );
  NANDN U13943 ( .A(x[5859]), .B(y[5859]), .Z(n23724) );
  NANDN U13944 ( .A(x[5860]), .B(y[5860]), .Z(n23721) );
  AND U13945 ( .A(n23724), .B(n23721), .Z(n58369) );
  NANDN U13946 ( .A(y[5858]), .B(x[5858]), .Z(n23726) );
  NANDN U13947 ( .A(y[5859]), .B(x[5859]), .Z(n23722) );
  NAND U13948 ( .A(n23726), .B(n23722), .Z(n58368) );
  NANDN U13949 ( .A(x[5857]), .B(y[5857]), .Z(n44909) );
  NANDN U13950 ( .A(x[5858]), .B(y[5858]), .Z(n23725) );
  AND U13951 ( .A(n44909), .B(n23725), .Z(n58367) );
  NANDN U13952 ( .A(y[5856]), .B(x[5856]), .Z(n9428) );
  NANDN U13953 ( .A(y[5857]), .B(x[5857]), .Z(n23727) );
  NAND U13954 ( .A(n9428), .B(n23727), .Z(n58365) );
  XNOR U13955 ( .A(x[5856]), .B(y[5856]), .Z(n23729) );
  NANDN U13956 ( .A(y[5854]), .B(x[5854]), .Z(n9429) );
  NANDN U13957 ( .A(y[5855]), .B(x[5855]), .Z(n23728) );
  NAND U13958 ( .A(n9429), .B(n23728), .Z(n58362) );
  XNOR U13959 ( .A(x[5854]), .B(y[5854]), .Z(n23731) );
  ANDN U13960 ( .B(y[5853]), .A(x[5853]), .Z(n44899) );
  NANDN U13961 ( .A(x[5851]), .B(y[5851]), .Z(n58359) );
  XOR U13962 ( .A(x[5852]), .B(y[5852]), .Z(n44896) );
  ANDN U13963 ( .B(n58359), .A(n44896), .Z(n18245) );
  XNOR U13964 ( .A(x[5850]), .B(y[5850]), .Z(n23733) );
  XNOR U13965 ( .A(x[5848]), .B(y[5848]), .Z(n23735) );
  NANDN U13966 ( .A(y[5846]), .B(x[5846]), .Z(n9430) );
  NANDN U13967 ( .A(y[5847]), .B(x[5847]), .Z(n23734) );
  NAND U13968 ( .A(n9430), .B(n23734), .Z(n58353) );
  XNOR U13969 ( .A(x[5846]), .B(y[5846]), .Z(n23737) );
  ANDN U13970 ( .B(y[5845]), .A(x[5845]), .Z(n44880) );
  NANDN U13971 ( .A(x[5843]), .B(y[5843]), .Z(n58349) );
  XNOR U13972 ( .A(x[5844]), .B(y[5844]), .Z(n23739) );
  AND U13973 ( .A(n58349), .B(n23739), .Z(n18230) );
  XNOR U13974 ( .A(x[5842]), .B(y[5842]), .Z(n23741) );
  NANDN U13975 ( .A(y[5840]), .B(x[5840]), .Z(n9431) );
  NANDN U13976 ( .A(y[5841]), .B(x[5841]), .Z(n23740) );
  NAND U13977 ( .A(n9431), .B(n23740), .Z(n58346) );
  XNOR U13978 ( .A(x[5840]), .B(y[5840]), .Z(n23743) );
  NANDN U13979 ( .A(y[5838]), .B(x[5838]), .Z(n9432) );
  NANDN U13980 ( .A(y[5839]), .B(x[5839]), .Z(n23742) );
  NAND U13981 ( .A(n9432), .B(n23742), .Z(n58343) );
  XNOR U13982 ( .A(x[5838]), .B(y[5838]), .Z(n23745) );
  ANDN U13983 ( .B(y[5837]), .A(x[5837]), .Z(n44863) );
  NANDN U13984 ( .A(x[5835]), .B(y[5835]), .Z(n58340) );
  NANDN U13985 ( .A(y[5834]), .B(x[5834]), .Z(n9433) );
  NANDN U13986 ( .A(y[5835]), .B(x[5835]), .Z(n23746) );
  AND U13987 ( .A(n9433), .B(n23746), .Z(n58338) );
  XNOR U13988 ( .A(y[5834]), .B(x[5834]), .Z(n23750) );
  NANDN U13989 ( .A(x[5833]), .B(y[5833]), .Z(n44854) );
  AND U13990 ( .A(n23750), .B(n44854), .Z(n58337) );
  NANDN U13991 ( .A(y[5832]), .B(x[5832]), .Z(n9434) );
  NANDN U13992 ( .A(y[5833]), .B(x[5833]), .Z(n23749) );
  AND U13993 ( .A(n9434), .B(n23749), .Z(n58336) );
  ANDN U13994 ( .B(y[5831]), .A(x[5831]), .Z(n23753) );
  XNOR U13995 ( .A(x[5832]), .B(y[5832]), .Z(n23752) );
  NANDN U13996 ( .A(y[5830]), .B(x[5830]), .Z(n9435) );
  NANDN U13997 ( .A(y[5831]), .B(x[5831]), .Z(n23751) );
  NAND U13998 ( .A(n9435), .B(n23751), .Z(n58332) );
  XNOR U13999 ( .A(x[5830]), .B(y[5830]), .Z(n23755) );
  ANDN U14000 ( .B(y[5829]), .A(x[5829]), .Z(n44845) );
  NANDN U14001 ( .A(x[5827]), .B(y[5827]), .Z(n58329) );
  NANDN U14002 ( .A(y[5826]), .B(x[5826]), .Z(n9436) );
  ANDN U14003 ( .B(x[5827]), .A(y[5827]), .Z(n44842) );
  ANDN U14004 ( .B(n9436), .A(n44842), .Z(n58327) );
  NANDN U14005 ( .A(x[5825]), .B(y[5825]), .Z(n51262) );
  XNOR U14006 ( .A(x[5826]), .B(y[5826]), .Z(n23757) );
  NANDN U14007 ( .A(x[5823]), .B(y[5823]), .Z(n23761) );
  NANDN U14008 ( .A(x[5824]), .B(y[5824]), .Z(n23758) );
  AND U14009 ( .A(n23761), .B(n23758), .Z(n58325) );
  NANDN U14010 ( .A(y[5822]), .B(x[5822]), .Z(n9437) );
  NANDN U14011 ( .A(y[5823]), .B(x[5823]), .Z(n23760) );
  NAND U14012 ( .A(n9437), .B(n23760), .Z(n58324) );
  XNOR U14013 ( .A(x[5822]), .B(y[5822]), .Z(n23763) );
  ANDN U14014 ( .B(y[5821]), .A(x[5821]), .Z(n44826) );
  NANDN U14015 ( .A(y[5820]), .B(x[5820]), .Z(n9438) );
  NANDN U14016 ( .A(y[5821]), .B(x[5821]), .Z(n23762) );
  AND U14017 ( .A(n9438), .B(n23762), .Z(n58321) );
  NANDN U14018 ( .A(x[5819]), .B(y[5819]), .Z(n51265) );
  XNOR U14019 ( .A(x[5820]), .B(y[5820]), .Z(n23765) );
  AND U14020 ( .A(n51265), .B(n23765), .Z(n18208) );
  XNOR U14021 ( .A(y[5818]), .B(x[5818]), .Z(n23768) );
  NANDN U14022 ( .A(x[5817]), .B(y[5817]), .Z(n44817) );
  AND U14023 ( .A(n23768), .B(n44817), .Z(n58318) );
  NANDN U14024 ( .A(y[5816]), .B(x[5816]), .Z(n9439) );
  NANDN U14025 ( .A(y[5817]), .B(x[5817]), .Z(n23767) );
  NAND U14026 ( .A(n9439), .B(n23767), .Z(n58316) );
  XNOR U14027 ( .A(x[5816]), .B(y[5816]), .Z(n23770) );
  NANDN U14028 ( .A(x[5815]), .B(y[5815]), .Z(n51266) );
  AND U14029 ( .A(n23770), .B(n51266), .Z(n18202) );
  NANDN U14030 ( .A(y[5814]), .B(x[5814]), .Z(n23771) );
  NANDN U14031 ( .A(y[5815]), .B(x[5815]), .Z(n23769) );
  NAND U14032 ( .A(n23771), .B(n23769), .Z(n58312) );
  NANDN U14033 ( .A(x[5813]), .B(y[5813]), .Z(n44808) );
  NANDN U14034 ( .A(x[5814]), .B(y[5814]), .Z(n44812) );
  AND U14035 ( .A(n44808), .B(n44812), .Z(n58310) );
  XNOR U14036 ( .A(x[5812]), .B(y[5812]), .Z(n23774) );
  XNOR U14037 ( .A(x[5810]), .B(y[5810]), .Z(n23776) );
  NANDN U14038 ( .A(y[5808]), .B(x[5808]), .Z(n9440) );
  NANDN U14039 ( .A(y[5809]), .B(x[5809]), .Z(n23775) );
  NAND U14040 ( .A(n9440), .B(n23775), .Z(n58296) );
  XNOR U14041 ( .A(x[5808]), .B(y[5808]), .Z(n23778) );
  NANDN U14042 ( .A(x[5807]), .B(y[5807]), .Z(n58292) );
  NANDN U14043 ( .A(y[5806]), .B(x[5806]), .Z(n9441) );
  NANDN U14044 ( .A(y[5807]), .B(x[5807]), .Z(n23777) );
  AND U14045 ( .A(n9441), .B(n23777), .Z(n58290) );
  XNOR U14046 ( .A(x[5806]), .B(y[5806]), .Z(n23780) );
  ANDN U14047 ( .B(y[5805]), .A(x[5805]), .Z(n44790) );
  ANDN U14048 ( .B(n23780), .A(n44790), .Z(n18186) );
  XNOR U14049 ( .A(x[5804]), .B(y[5804]), .Z(n23782) );
  XNOR U14050 ( .A(x[5802]), .B(y[5802]), .Z(n23784) );
  NANDN U14051 ( .A(y[5800]), .B(x[5800]), .Z(n9442) );
  NANDN U14052 ( .A(y[5801]), .B(x[5801]), .Z(n23783) );
  NAND U14053 ( .A(n9442), .B(n23783), .Z(n58277) );
  XOR U14054 ( .A(x[5800]), .B(y[5800]), .Z(n44780) );
  NANDN U14055 ( .A(x[5799]), .B(y[5799]), .Z(n58276) );
  NANDN U14056 ( .A(y[5798]), .B(x[5798]), .Z(n9443) );
  ANDN U14057 ( .B(x[5799]), .A(y[5799]), .Z(n44779) );
  ANDN U14058 ( .B(n9443), .A(n44779), .Z(n58274) );
  XNOR U14059 ( .A(x[5798]), .B(y[5798]), .Z(n23786) );
  ANDN U14060 ( .B(y[5797]), .A(x[5797]), .Z(n44771) );
  ANDN U14061 ( .B(n23786), .A(n44771), .Z(n18172) );
  XNOR U14062 ( .A(x[5796]), .B(y[5796]), .Z(n23788) );
  XNOR U14063 ( .A(x[5794]), .B(y[5794]), .Z(n23790) );
  NANDN U14064 ( .A(y[5792]), .B(x[5792]), .Z(n9444) );
  NANDN U14065 ( .A(y[5793]), .B(x[5793]), .Z(n23789) );
  NAND U14066 ( .A(n9444), .B(n23789), .Z(n51270) );
  XNOR U14067 ( .A(x[5792]), .B(y[5792]), .Z(n44761) );
  NANDN U14068 ( .A(x[5791]), .B(y[5791]), .Z(n51271) );
  NANDN U14069 ( .A(y[5790]), .B(x[5790]), .Z(n9445) );
  ANDN U14070 ( .B(x[5791]), .A(y[5791]), .Z(n44760) );
  ANDN U14071 ( .B(n9445), .A(n44760), .Z(n58263) );
  XNOR U14072 ( .A(x[5790]), .B(y[5790]), .Z(n44754) );
  ANDN U14073 ( .B(y[5789]), .A(x[5789]), .Z(n44750) );
  ANDN U14074 ( .B(n44754), .A(n44750), .Z(n18158) );
  XNOR U14075 ( .A(x[5788]), .B(y[5788]), .Z(n23792) );
  NANDN U14076 ( .A(y[5786]), .B(x[5786]), .Z(n9446) );
  NANDN U14077 ( .A(y[5787]), .B(x[5787]), .Z(n23791) );
  NAND U14078 ( .A(n9446), .B(n23791), .Z(n58259) );
  XNOR U14079 ( .A(x[5786]), .B(y[5786]), .Z(n23794) );
  NANDN U14080 ( .A(y[5784]), .B(x[5784]), .Z(n9447) );
  NANDN U14081 ( .A(y[5785]), .B(x[5785]), .Z(n23793) );
  NAND U14082 ( .A(n9447), .B(n23793), .Z(n58256) );
  XNOR U14083 ( .A(x[5784]), .B(y[5784]), .Z(n23796) );
  NANDN U14084 ( .A(x[5783]), .B(y[5783]), .Z(n58255) );
  NANDN U14085 ( .A(y[5782]), .B(x[5782]), .Z(n9448) );
  NANDN U14086 ( .A(y[5783]), .B(x[5783]), .Z(n23795) );
  AND U14087 ( .A(n9448), .B(n23795), .Z(n58253) );
  NANDN U14088 ( .A(x[5781]), .B(y[5781]), .Z(n51276) );
  XNOR U14089 ( .A(x[5782]), .B(y[5782]), .Z(n23798) );
  AND U14090 ( .A(n51276), .B(n23798), .Z(n18145) );
  XNOR U14091 ( .A(x[5780]), .B(y[5780]), .Z(n23800) );
  NANDN U14092 ( .A(y[5778]), .B(x[5778]), .Z(n23802) );
  NANDN U14093 ( .A(y[5779]), .B(x[5779]), .Z(n23799) );
  NAND U14094 ( .A(n23802), .B(n23799), .Z(n58248) );
  NANDN U14095 ( .A(x[5777]), .B(y[5777]), .Z(n23804) );
  NANDN U14096 ( .A(x[5778]), .B(y[5778]), .Z(n23801) );
  AND U14097 ( .A(n23804), .B(n23801), .Z(n58247) );
  NANDN U14098 ( .A(y[5776]), .B(x[5776]), .Z(n23806) );
  NANDN U14099 ( .A(y[5777]), .B(x[5777]), .Z(n23803) );
  NAND U14100 ( .A(n23806), .B(n23803), .Z(n58246) );
  NANDN U14101 ( .A(x[5775]), .B(y[5775]), .Z(n23808) );
  NANDN U14102 ( .A(x[5776]), .B(y[5776]), .Z(n23805) );
  AND U14103 ( .A(n23808), .B(n23805), .Z(n58245) );
  XNOR U14104 ( .A(x[5774]), .B(y[5774]), .Z(n23810) );
  NANDN U14105 ( .A(y[5772]), .B(x[5772]), .Z(n44715) );
  NANDN U14106 ( .A(y[5773]), .B(x[5773]), .Z(n23809) );
  AND U14107 ( .A(n44715), .B(n23809), .Z(n51277) );
  NANDN U14108 ( .A(x[5769]), .B(y[5769]), .Z(n23814) );
  NANDN U14109 ( .A(x[5770]), .B(y[5770]), .Z(n23813) );
  NAND U14110 ( .A(n23814), .B(n23813), .Z(n58240) );
  NANDN U14111 ( .A(y[5769]), .B(x[5769]), .Z(n44709) );
  ANDN U14112 ( .B(x[5768]), .A(y[5768]), .Z(n44703) );
  ANDN U14113 ( .B(n44709), .A(n44703), .Z(n58239) );
  NANDN U14114 ( .A(x[5763]), .B(y[5763]), .Z(n23825) );
  NANDN U14115 ( .A(x[5764]), .B(y[5764]), .Z(n23821) );
  NAND U14116 ( .A(n23825), .B(n23821), .Z(n58232) );
  NANDN U14117 ( .A(y[5762]), .B(x[5762]), .Z(n23826) );
  NANDN U14118 ( .A(y[5763]), .B(x[5763]), .Z(n23823) );
  AND U14119 ( .A(n23826), .B(n23823), .Z(n51280) );
  XNOR U14120 ( .A(x[5758]), .B(y[5758]), .Z(n23831) );
  NANDN U14121 ( .A(y[5756]), .B(x[5756]), .Z(n9449) );
  NANDN U14122 ( .A(y[5757]), .B(x[5757]), .Z(n23830) );
  AND U14123 ( .A(n9449), .B(n23830), .Z(n58227) );
  XNOR U14124 ( .A(x[5756]), .B(y[5756]), .Z(n23833) );
  NANDN U14125 ( .A(x[5755]), .B(y[5755]), .Z(n58225) );
  XNOR U14126 ( .A(x[5754]), .B(y[5754]), .Z(n23835) );
  NANDN U14127 ( .A(y[5752]), .B(x[5752]), .Z(n9450) );
  NANDN U14128 ( .A(y[5753]), .B(x[5753]), .Z(n23834) );
  NAND U14129 ( .A(n9450), .B(n23834), .Z(n58220) );
  XNOR U14130 ( .A(x[5752]), .B(y[5752]), .Z(n23837) );
  NANDN U14131 ( .A(x[5751]), .B(y[5751]), .Z(n51284) );
  NANDN U14132 ( .A(y[5750]), .B(x[5750]), .Z(n9451) );
  NANDN U14133 ( .A(y[5751]), .B(x[5751]), .Z(n23836) );
  AND U14134 ( .A(n9451), .B(n23836), .Z(n58219) );
  XNOR U14135 ( .A(x[5750]), .B(y[5750]), .Z(n23839) );
  ANDN U14136 ( .B(y[5749]), .A(x[5749]), .Z(n44659) );
  ANDN U14137 ( .B(n23839), .A(n44659), .Z(n18100) );
  NANDN U14138 ( .A(x[5747]), .B(y[5747]), .Z(n44654) );
  NANDN U14139 ( .A(x[5748]), .B(y[5748]), .Z(n44661) );
  AND U14140 ( .A(n44654), .B(n44661), .Z(n58216) );
  XNOR U14141 ( .A(x[5746]), .B(y[5746]), .Z(n23843) );
  NANDN U14142 ( .A(y[5744]), .B(x[5744]), .Z(n9452) );
  NANDN U14143 ( .A(y[5745]), .B(x[5745]), .Z(n23842) );
  NAND U14144 ( .A(n9452), .B(n23842), .Z(n58214) );
  XNOR U14145 ( .A(x[5744]), .B(y[5744]), .Z(n23845) );
  NANDN U14146 ( .A(x[5743]), .B(y[5743]), .Z(n58211) );
  NANDN U14147 ( .A(y[5742]), .B(x[5742]), .Z(n9453) );
  NANDN U14148 ( .A(y[5743]), .B(x[5743]), .Z(n23844) );
  AND U14149 ( .A(n9453), .B(n23844), .Z(n58210) );
  NANDN U14150 ( .A(x[5741]), .B(y[5741]), .Z(n58209) );
  XNOR U14151 ( .A(x[5742]), .B(y[5742]), .Z(n23847) );
  AND U14152 ( .A(n58209), .B(n23847), .Z(n18088) );
  NANDN U14153 ( .A(y[5740]), .B(x[5740]), .Z(n9454) );
  NANDN U14154 ( .A(y[5741]), .B(x[5741]), .Z(n23846) );
  NAND U14155 ( .A(n9454), .B(n23846), .Z(n58208) );
  XNOR U14156 ( .A(x[5740]), .B(y[5740]), .Z(n23849) );
  NANDN U14157 ( .A(y[5738]), .B(x[5738]), .Z(n9455) );
  NANDN U14158 ( .A(y[5739]), .B(x[5739]), .Z(n23848) );
  NAND U14159 ( .A(n9455), .B(n23848), .Z(n58205) );
  XNOR U14160 ( .A(x[5738]), .B(y[5738]), .Z(n23851) );
  NANDN U14161 ( .A(y[5736]), .B(x[5736]), .Z(n9456) );
  NANDN U14162 ( .A(y[5737]), .B(x[5737]), .Z(n23850) );
  NAND U14163 ( .A(n9456), .B(n23850), .Z(n58204) );
  XNOR U14164 ( .A(x[5736]), .B(y[5736]), .Z(n44631) );
  ANDN U14165 ( .B(y[5735]), .A(x[5735]), .Z(n58202) );
  NANDN U14166 ( .A(y[5734]), .B(x[5734]), .Z(n9457) );
  ANDN U14167 ( .B(x[5735]), .A(y[5735]), .Z(n44630) );
  ANDN U14168 ( .B(n9457), .A(n44630), .Z(n58201) );
  XNOR U14169 ( .A(x[5734]), .B(y[5734]), .Z(n44625) );
  ANDN U14170 ( .B(y[5733]), .A(x[5733]), .Z(n44620) );
  ANDN U14171 ( .B(n44625), .A(n44620), .Z(n18076) );
  ANDN U14172 ( .B(x[5731]), .A(y[5731]), .Z(n44617) );
  NANDN U14173 ( .A(y[5730]), .B(x[5730]), .Z(n9458) );
  NANDN U14174 ( .A(n44617), .B(n9458), .Z(n51293) );
  XNOR U14175 ( .A(x[5730]), .B(y[5730]), .Z(n23853) );
  NANDN U14176 ( .A(x[5729]), .B(y[5729]), .Z(n58195) );
  NANDN U14177 ( .A(y[5728]), .B(x[5728]), .Z(n9459) );
  NANDN U14178 ( .A(y[5729]), .B(x[5729]), .Z(n23852) );
  AND U14179 ( .A(n9459), .B(n23852), .Z(n58194) );
  XNOR U14180 ( .A(x[5728]), .B(y[5728]), .Z(n23855) );
  ANDN U14181 ( .B(y[5727]), .A(x[5727]), .Z(n44604) );
  ANDN U14182 ( .B(n23855), .A(n44604), .Z(n18067) );
  XNOR U14183 ( .A(x[5726]), .B(y[5726]), .Z(n23857) );
  XNOR U14184 ( .A(x[5724]), .B(y[5724]), .Z(n23859) );
  NANDN U14185 ( .A(y[5722]), .B(x[5722]), .Z(n9460) );
  NANDN U14186 ( .A(y[5723]), .B(x[5723]), .Z(n23858) );
  NAND U14187 ( .A(n9460), .B(n23858), .Z(n58187) );
  XNOR U14188 ( .A(x[5722]), .B(y[5722]), .Z(n23861) );
  NANDN U14189 ( .A(x[5721]), .B(y[5721]), .Z(n58185) );
  NANDN U14190 ( .A(y[5720]), .B(x[5720]), .Z(n9461) );
  NANDN U14191 ( .A(y[5721]), .B(x[5721]), .Z(n23860) );
  AND U14192 ( .A(n9461), .B(n23860), .Z(n58184) );
  XNOR U14193 ( .A(x[5720]), .B(y[5720]), .Z(n23863) );
  NANDN U14194 ( .A(x[5719]), .B(y[5719]), .Z(n58182) );
  AND U14195 ( .A(n23863), .B(n58182), .Z(n18053) );
  NANDN U14196 ( .A(x[5717]), .B(y[5717]), .Z(n58181) );
  XNOR U14197 ( .A(x[5718]), .B(y[5718]), .Z(n23865) );
  AND U14198 ( .A(n58181), .B(n23865), .Z(n18049) );
  NANDN U14199 ( .A(y[5714]), .B(x[5714]), .Z(n9462) );
  NANDN U14200 ( .A(y[5715]), .B(x[5715]), .Z(n23866) );
  NAND U14201 ( .A(n9462), .B(n23866), .Z(n51299) );
  XNOR U14202 ( .A(x[5714]), .B(y[5714]), .Z(n23869) );
  ANDN U14203 ( .B(y[5713]), .A(x[5713]), .Z(n44573) );
  NANDN U14204 ( .A(x[5711]), .B(y[5711]), .Z(n23870) );
  IV U14205 ( .A(n23870), .Z(n58174) );
  XOR U14206 ( .A(x[5712]), .B(y[5712]), .Z(n44570) );
  NOR U14207 ( .A(n58174), .B(n44570), .Z(n18039) );
  XNOR U14208 ( .A(x[5710]), .B(y[5710]), .Z(n23872) );
  XNOR U14209 ( .A(x[5708]), .B(y[5708]), .Z(n44561) );
  ANDN U14210 ( .B(x[5707]), .A(y[5707]), .Z(n44560) );
  NANDN U14211 ( .A(y[5706]), .B(x[5706]), .Z(n23874) );
  NANDN U14212 ( .A(n44560), .B(n23874), .Z(n58169) );
  NANDN U14213 ( .A(x[5705]), .B(y[5705]), .Z(n23876) );
  NANDN U14214 ( .A(x[5706]), .B(y[5706]), .Z(n23873) );
  AND U14215 ( .A(n23876), .B(n23873), .Z(n58168) );
  NANDN U14216 ( .A(y[5704]), .B(x[5704]), .Z(n23878) );
  NANDN U14217 ( .A(y[5705]), .B(x[5705]), .Z(n23875) );
  NAND U14218 ( .A(n23878), .B(n23875), .Z(n58167) );
  NANDN U14219 ( .A(x[5703]), .B(y[5703]), .Z(n44549) );
  NANDN U14220 ( .A(x[5704]), .B(y[5704]), .Z(n23877) );
  AND U14221 ( .A(n44549), .B(n23877), .Z(n58166) );
  XNOR U14222 ( .A(x[5702]), .B(y[5702]), .Z(n23881) );
  NANDN U14223 ( .A(y[5700]), .B(x[5700]), .Z(n9463) );
  NANDN U14224 ( .A(y[5701]), .B(x[5701]), .Z(n23880) );
  NAND U14225 ( .A(n9463), .B(n23880), .Z(n58162) );
  XNOR U14226 ( .A(y[5700]), .B(x[5700]), .Z(n23883) );
  NANDN U14227 ( .A(x[5699]), .B(y[5699]), .Z(n23884) );
  AND U14228 ( .A(n23883), .B(n23884), .Z(n58161) );
  NANDN U14229 ( .A(y[5698]), .B(x[5698]), .Z(n9464) );
  NANDN U14230 ( .A(y[5699]), .B(x[5699]), .Z(n23882) );
  NAND U14231 ( .A(n9464), .B(n23882), .Z(n58159) );
  NANDN U14232 ( .A(y[5696]), .B(x[5696]), .Z(n9465) );
  NANDN U14233 ( .A(y[5697]), .B(x[5697]), .Z(n23885) );
  AND U14234 ( .A(n9465), .B(n23885), .Z(n58158) );
  XNOR U14235 ( .A(x[5696]), .B(y[5696]), .Z(n23888) );
  XNOR U14236 ( .A(x[5694]), .B(y[5694]), .Z(n23891) );
  NANDN U14237 ( .A(y[5692]), .B(x[5692]), .Z(n23893) );
  NANDN U14238 ( .A(y[5693]), .B(x[5693]), .Z(n23890) );
  NAND U14239 ( .A(n23893), .B(n23890), .Z(n58155) );
  NANDN U14240 ( .A(x[5691]), .B(y[5691]), .Z(n44523) );
  NANDN U14241 ( .A(x[5692]), .B(y[5692]), .Z(n23892) );
  AND U14242 ( .A(n44523), .B(n23892), .Z(n58154) );
  NANDN U14243 ( .A(y[5690]), .B(x[5690]), .Z(n9466) );
  NANDN U14244 ( .A(y[5691]), .B(x[5691]), .Z(n23894) );
  NAND U14245 ( .A(n9466), .B(n23894), .Z(n58153) );
  NANDN U14246 ( .A(y[5688]), .B(x[5688]), .Z(n9467) );
  NANDN U14247 ( .A(y[5689]), .B(x[5689]), .Z(n23895) );
  AND U14248 ( .A(n9467), .B(n23895), .Z(n58150) );
  XNOR U14249 ( .A(x[5688]), .B(y[5688]), .Z(n23898) );
  XNOR U14250 ( .A(x[5686]), .B(y[5686]), .Z(n23901) );
  NANDN U14251 ( .A(y[5684]), .B(x[5684]), .Z(n9468) );
  NANDN U14252 ( .A(y[5685]), .B(x[5685]), .Z(n23900) );
  NAND U14253 ( .A(n9468), .B(n23900), .Z(n58144) );
  XNOR U14254 ( .A(x[5684]), .B(y[5684]), .Z(n44508) );
  ANDN U14255 ( .B(y[5683]), .A(x[5683]), .Z(n23902) );
  NANDN U14256 ( .A(y[5682]), .B(x[5682]), .Z(n9469) );
  ANDN U14257 ( .B(x[5683]), .A(y[5683]), .Z(n44507) );
  ANDN U14258 ( .B(n9469), .A(n44507), .Z(n58143) );
  XNOR U14259 ( .A(x[5682]), .B(y[5682]), .Z(n23904) );
  ANDN U14260 ( .B(y[5681]), .A(x[5681]), .Z(n44499) );
  ANDN U14261 ( .B(n23904), .A(n44499), .Z(n17993) );
  XNOR U14262 ( .A(x[5680]), .B(y[5680]), .Z(n23906) );
  XNOR U14263 ( .A(x[5678]), .B(y[5678]), .Z(n23908) );
  NANDN U14264 ( .A(y[5676]), .B(x[5676]), .Z(n9470) );
  NANDN U14265 ( .A(y[5677]), .B(x[5677]), .Z(n23907) );
  NAND U14266 ( .A(n9470), .B(n23907), .Z(n58131) );
  XNOR U14267 ( .A(x[5676]), .B(y[5676]), .Z(n23910) );
  NANDN U14268 ( .A(x[5675]), .B(y[5675]), .Z(n58129) );
  NANDN U14269 ( .A(y[5674]), .B(x[5674]), .Z(n9471) );
  NANDN U14270 ( .A(y[5675]), .B(x[5675]), .Z(n23909) );
  AND U14271 ( .A(n9471), .B(n23909), .Z(n58128) );
  NANDN U14272 ( .A(x[5671]), .B(y[5671]), .Z(n44479) );
  NANDN U14273 ( .A(x[5672]), .B(y[5672]), .Z(n23913) );
  NAND U14274 ( .A(n44479), .B(n23913), .Z(n51314) );
  NANDN U14275 ( .A(y[5670]), .B(x[5670]), .Z(n9472) );
  NANDN U14276 ( .A(y[5671]), .B(x[5671]), .Z(n23915) );
  AND U14277 ( .A(n9472), .B(n23915), .Z(n58126) );
  ANDN U14278 ( .B(y[5669]), .A(x[5669]), .Z(n44473) );
  XNOR U14279 ( .A(x[5670]), .B(y[5670]), .Z(n23917) );
  NANDN U14280 ( .A(y[5668]), .B(x[5668]), .Z(n9473) );
  NANDN U14281 ( .A(y[5669]), .B(x[5669]), .Z(n23916) );
  AND U14282 ( .A(n9473), .B(n23916), .Z(n58125) );
  NANDN U14283 ( .A(x[5667]), .B(y[5667]), .Z(n58123) );
  XNOR U14284 ( .A(x[5668]), .B(y[5668]), .Z(n23919) );
  AND U14285 ( .A(n58123), .B(n23919), .Z(n17971) );
  NANDN U14286 ( .A(y[5666]), .B(x[5666]), .Z(n23921) );
  NANDN U14287 ( .A(y[5667]), .B(x[5667]), .Z(n23918) );
  NAND U14288 ( .A(n23921), .B(n23918), .Z(n58122) );
  NANDN U14289 ( .A(x[5665]), .B(y[5665]), .Z(n44464) );
  NANDN U14290 ( .A(x[5666]), .B(y[5666]), .Z(n23920) );
  AND U14291 ( .A(n44464), .B(n23920), .Z(n58121) );
  XNOR U14292 ( .A(x[5664]), .B(y[5664]), .Z(n23924) );
  NANDN U14293 ( .A(y[5662]), .B(x[5662]), .Z(n9474) );
  NANDN U14294 ( .A(y[5663]), .B(x[5663]), .Z(n23923) );
  NAND U14295 ( .A(n9474), .B(n23923), .Z(n58118) );
  XNOR U14296 ( .A(x[5662]), .B(y[5662]), .Z(n23926) );
  NANDN U14297 ( .A(y[5660]), .B(x[5660]), .Z(n9475) );
  NANDN U14298 ( .A(y[5661]), .B(x[5661]), .Z(n23925) );
  NAND U14299 ( .A(n9475), .B(n23925), .Z(n58115) );
  XNOR U14300 ( .A(x[5660]), .B(y[5660]), .Z(n23928) );
  ANDN U14301 ( .B(y[5659]), .A(x[5659]), .Z(n23929) );
  XNOR U14302 ( .A(x[5658]), .B(y[5658]), .Z(n23931) );
  NANDN U14303 ( .A(x[5657]), .B(y[5657]), .Z(n58112) );
  AND U14304 ( .A(n23931), .B(n58112), .Z(n17955) );
  XNOR U14305 ( .A(x[5654]), .B(y[5654]), .Z(n23933) );
  NANDN U14306 ( .A(y[5652]), .B(x[5652]), .Z(n9476) );
  NANDN U14307 ( .A(y[5653]), .B(x[5653]), .Z(n23932) );
  NAND U14308 ( .A(n9476), .B(n23932), .Z(n58104) );
  XNOR U14309 ( .A(y[5652]), .B(x[5652]), .Z(n23935) );
  NANDN U14310 ( .A(x[5651]), .B(y[5651]), .Z(n23936) );
  AND U14311 ( .A(n23935), .B(n23936), .Z(n58103) );
  NANDN U14312 ( .A(y[5650]), .B(x[5650]), .Z(n9477) );
  NANDN U14313 ( .A(y[5651]), .B(x[5651]), .Z(n23934) );
  NAND U14314 ( .A(n9477), .B(n23934), .Z(n58102) );
  NANDN U14315 ( .A(y[5648]), .B(x[5648]), .Z(n9478) );
  NANDN U14316 ( .A(y[5649]), .B(x[5649]), .Z(n23937) );
  AND U14317 ( .A(n9478), .B(n23937), .Z(n58101) );
  XNOR U14318 ( .A(x[5648]), .B(y[5648]), .Z(n23940) );
  XNOR U14319 ( .A(x[5646]), .B(y[5646]), .Z(n23943) );
  NANDN U14320 ( .A(y[5644]), .B(x[5644]), .Z(n9479) );
  NANDN U14321 ( .A(y[5645]), .B(x[5645]), .Z(n23942) );
  NAND U14322 ( .A(n9479), .B(n23942), .Z(n58095) );
  XNOR U14323 ( .A(x[5644]), .B(y[5644]), .Z(n23945) );
  NANDN U14324 ( .A(x[5643]), .B(y[5643]), .Z(n58094) );
  NANDN U14325 ( .A(y[5642]), .B(x[5642]), .Z(n9480) );
  NANDN U14326 ( .A(y[5643]), .B(x[5643]), .Z(n23944) );
  AND U14327 ( .A(n9480), .B(n23944), .Z(n58092) );
  XNOR U14328 ( .A(x[5642]), .B(y[5642]), .Z(n23947) );
  ANDN U14329 ( .B(y[5641]), .A(x[5641]), .Z(n44412) );
  ANDN U14330 ( .B(n23947), .A(n44412), .Z(n17929) );
  XNOR U14331 ( .A(x[5640]), .B(y[5640]), .Z(n23949) );
  XNOR U14332 ( .A(x[5638]), .B(y[5638]), .Z(n23951) );
  NANDN U14333 ( .A(y[5636]), .B(x[5636]), .Z(n9481) );
  NANDN U14334 ( .A(y[5637]), .B(x[5637]), .Z(n23950) );
  NAND U14335 ( .A(n9481), .B(n23950), .Z(n58083) );
  XNOR U14336 ( .A(x[5636]), .B(y[5636]), .Z(n23953) );
  NANDN U14337 ( .A(x[5635]), .B(y[5635]), .Z(n58082) );
  NANDN U14338 ( .A(y[5634]), .B(x[5634]), .Z(n9482) );
  NANDN U14339 ( .A(y[5635]), .B(x[5635]), .Z(n23952) );
  AND U14340 ( .A(n9482), .B(n23952), .Z(n58080) );
  XNOR U14341 ( .A(x[5634]), .B(y[5634]), .Z(n23955) );
  ANDN U14342 ( .B(y[5633]), .A(x[5633]), .Z(n44395) );
  ANDN U14343 ( .B(n23955), .A(n44395), .Z(n17915) );
  XNOR U14344 ( .A(x[5632]), .B(y[5632]), .Z(n44393) );
  ANDN U14345 ( .B(x[5631]), .A(y[5631]), .Z(n44392) );
  NANDN U14346 ( .A(y[5630]), .B(x[5630]), .Z(n9483) );
  NANDN U14347 ( .A(n44392), .B(n9483), .Z(n58076) );
  XNOR U14348 ( .A(x[5630]), .B(y[5630]), .Z(n23957) );
  NANDN U14349 ( .A(y[5628]), .B(x[5628]), .Z(n9484) );
  NANDN U14350 ( .A(y[5629]), .B(x[5629]), .Z(n23956) );
  NAND U14351 ( .A(n9484), .B(n23956), .Z(n58071) );
  XNOR U14352 ( .A(x[5628]), .B(y[5628]), .Z(n23959) );
  NANDN U14353 ( .A(x[5627]), .B(y[5627]), .Z(n58070) );
  NANDN U14354 ( .A(y[5626]), .B(x[5626]), .Z(n9485) );
  NANDN U14355 ( .A(y[5627]), .B(x[5627]), .Z(n23958) );
  AND U14356 ( .A(n9485), .B(n23958), .Z(n58068) );
  XNOR U14357 ( .A(x[5626]), .B(y[5626]), .Z(n23961) );
  NANDN U14358 ( .A(x[5625]), .B(y[5625]), .Z(n51328) );
  AND U14359 ( .A(n23961), .B(n51328), .Z(n17902) );
  XNOR U14360 ( .A(x[5624]), .B(y[5624]), .Z(n23963) );
  NANDN U14361 ( .A(x[5621]), .B(y[5621]), .Z(n44368) );
  NANDN U14362 ( .A(x[5622]), .B(y[5622]), .Z(n23964) );
  AND U14363 ( .A(n44368), .B(n23964), .Z(n58063) );
  NANDN U14364 ( .A(y[5620]), .B(x[5620]), .Z(n9486) );
  NANDN U14365 ( .A(y[5621]), .B(x[5621]), .Z(n23966) );
  NAND U14366 ( .A(n9486), .B(n23966), .Z(n58062) );
  NANDN U14367 ( .A(x[5619]), .B(y[5619]), .Z(n51330) );
  XNOR U14368 ( .A(x[5620]), .B(y[5620]), .Z(n23968) );
  NANDN U14369 ( .A(y[5618]), .B(x[5618]), .Z(n9487) );
  NANDN U14370 ( .A(y[5619]), .B(x[5619]), .Z(n23967) );
  AND U14371 ( .A(n9487), .B(n23967), .Z(n58061) );
  XNOR U14372 ( .A(y[5618]), .B(x[5618]), .Z(n23971) );
  NANDN U14373 ( .A(x[5617]), .B(y[5617]), .Z(n44358) );
  NAND U14374 ( .A(n23971), .B(n44358), .Z(n58060) );
  NANDN U14375 ( .A(y[5616]), .B(x[5616]), .Z(n9488) );
  NANDN U14376 ( .A(y[5617]), .B(x[5617]), .Z(n23970) );
  AND U14377 ( .A(n9488), .B(n23970), .Z(n51332) );
  XNOR U14378 ( .A(x[5612]), .B(y[5612]), .Z(n44346) );
  ANDN U14379 ( .B(y[5611]), .A(x[5611]), .Z(n23976) );
  ANDN U14380 ( .B(n44346), .A(n23976), .Z(n17881) );
  NANDN U14381 ( .A(x[5609]), .B(y[5609]), .Z(n44337) );
  NANDN U14382 ( .A(x[5610]), .B(y[5610]), .Z(n23977) );
  AND U14383 ( .A(n44337), .B(n23977), .Z(n58052) );
  NANDN U14384 ( .A(y[5608]), .B(x[5608]), .Z(n9489) );
  NANDN U14385 ( .A(y[5609]), .B(x[5609]), .Z(n23979) );
  NAND U14386 ( .A(n9489), .B(n23979), .Z(n58051) );
  XNOR U14387 ( .A(x[5608]), .B(y[5608]), .Z(n23980) );
  NANDN U14388 ( .A(x[5607]), .B(y[5607]), .Z(n51336) );
  AND U14389 ( .A(n23980), .B(n51336), .Z(n17876) );
  NANDN U14390 ( .A(y[5606]), .B(x[5606]), .Z(n23983) );
  NANDN U14391 ( .A(y[5607]), .B(x[5607]), .Z(n23981) );
  NAND U14392 ( .A(n23983), .B(n23981), .Z(n58050) );
  NANDN U14393 ( .A(x[5605]), .B(y[5605]), .Z(n44328) );
  NANDN U14394 ( .A(x[5606]), .B(y[5606]), .Z(n23982) );
  AND U14395 ( .A(n44328), .B(n23982), .Z(n58049) );
  XNOR U14396 ( .A(x[5604]), .B(y[5604]), .Z(n23986) );
  XNOR U14397 ( .A(x[5602]), .B(y[5602]), .Z(n23988) );
  NANDN U14398 ( .A(y[5600]), .B(x[5600]), .Z(n23990) );
  NANDN U14399 ( .A(y[5601]), .B(x[5601]), .Z(n23987) );
  NAND U14400 ( .A(n23990), .B(n23987), .Z(n58042) );
  NANDN U14401 ( .A(x[5599]), .B(y[5599]), .Z(n23992) );
  NANDN U14402 ( .A(x[5600]), .B(y[5600]), .Z(n23989) );
  AND U14403 ( .A(n23992), .B(n23989), .Z(n58041) );
  NANDN U14404 ( .A(y[5598]), .B(x[5598]), .Z(n9490) );
  NANDN U14405 ( .A(y[5599]), .B(x[5599]), .Z(n23991) );
  NAND U14406 ( .A(n9490), .B(n23991), .Z(n58040) );
  XNOR U14407 ( .A(x[5598]), .B(y[5598]), .Z(n23994) );
  NANDN U14408 ( .A(x[5597]), .B(y[5597]), .Z(n58039) );
  AND U14409 ( .A(n23994), .B(n58039), .Z(n17861) );
  XNOR U14410 ( .A(y[5596]), .B(x[5596]), .Z(n23996) );
  NANDN U14411 ( .A(x[5595]), .B(y[5595]), .Z(n23997) );
  AND U14412 ( .A(n23996), .B(n23997), .Z(n58036) );
  NANDN U14413 ( .A(y[5594]), .B(x[5594]), .Z(n9491) );
  NANDN U14414 ( .A(y[5595]), .B(x[5595]), .Z(n23995) );
  NAND U14415 ( .A(n9491), .B(n23995), .Z(n58035) );
  XNOR U14416 ( .A(y[5594]), .B(x[5594]), .Z(n24000) );
  NANDN U14417 ( .A(x[5593]), .B(y[5593]), .Z(n24001) );
  AND U14418 ( .A(n24000), .B(n24001), .Z(n58034) );
  NANDN U14419 ( .A(y[5592]), .B(x[5592]), .Z(n24003) );
  NANDN U14420 ( .A(y[5593]), .B(x[5593]), .Z(n23999) );
  NAND U14421 ( .A(n24003), .B(n23999), .Z(n58033) );
  NANDN U14422 ( .A(x[5591]), .B(y[5591]), .Z(n44299) );
  NANDN U14423 ( .A(x[5592]), .B(y[5592]), .Z(n24002) );
  AND U14424 ( .A(n44299), .B(n24002), .Z(n58032) );
  NANDN U14425 ( .A(y[5590]), .B(x[5590]), .Z(n9492) );
  NANDN U14426 ( .A(y[5591]), .B(x[5591]), .Z(n24004) );
  NAND U14427 ( .A(n9492), .B(n24004), .Z(n58031) );
  XNOR U14428 ( .A(x[5590]), .B(y[5590]), .Z(n24006) );
  NANDN U14429 ( .A(x[5587]), .B(y[5587]), .Z(n24010) );
  NANDN U14430 ( .A(x[5588]), .B(y[5588]), .Z(n24007) );
  AND U14431 ( .A(n24010), .B(n24007), .Z(n58028) );
  XNOR U14432 ( .A(x[5586]), .B(y[5586]), .Z(n24012) );
  NANDN U14433 ( .A(x[5585]), .B(y[5585]), .Z(n58026) );
  AND U14434 ( .A(n24012), .B(n58026), .Z(n17845) );
  NANDN U14435 ( .A(y[5584]), .B(x[5584]), .Z(n9493) );
  NANDN U14436 ( .A(y[5585]), .B(x[5585]), .Z(n24011) );
  AND U14437 ( .A(n9493), .B(n24011), .Z(n58024) );
  NANDN U14438 ( .A(x[5583]), .B(y[5583]), .Z(n51343) );
  XNOR U14439 ( .A(x[5584]), .B(y[5584]), .Z(n24014) );
  AND U14440 ( .A(n51343), .B(n24014), .Z(n17842) );
  XNOR U14441 ( .A(y[5582]), .B(x[5582]), .Z(n24016) );
  NANDN U14442 ( .A(x[5581]), .B(y[5581]), .Z(n44276) );
  AND U14443 ( .A(n24016), .B(n44276), .Z(n58022) );
  NANDN U14444 ( .A(y[5580]), .B(x[5580]), .Z(n9494) );
  NANDN U14445 ( .A(y[5581]), .B(x[5581]), .Z(n24015) );
  NAND U14446 ( .A(n9494), .B(n24015), .Z(n58021) );
  NANDN U14447 ( .A(x[5579]), .B(y[5579]), .Z(n58020) );
  XNOR U14448 ( .A(x[5580]), .B(y[5580]), .Z(n44274) );
  ANDN U14449 ( .B(x[5578]), .A(y[5578]), .Z(n44269) );
  ANDN U14450 ( .B(x[5579]), .A(y[5579]), .Z(n44273) );
  NOR U14451 ( .A(n44269), .B(n44273), .Z(n58018) );
  NANDN U14452 ( .A(x[5577]), .B(y[5577]), .Z(n44262) );
  NANDN U14453 ( .A(x[5578]), .B(y[5578]), .Z(n24017) );
  NAND U14454 ( .A(n44262), .B(n24017), .Z(n58017) );
  NANDN U14455 ( .A(y[5577]), .B(x[5577]), .Z(n44265) );
  NANDN U14456 ( .A(y[5576]), .B(x[5576]), .Z(n9495) );
  AND U14457 ( .A(n44265), .B(n9495), .Z(n58016) );
  NANDN U14458 ( .A(x[5575]), .B(y[5575]), .Z(n44256) );
  NANDN U14459 ( .A(x[5576]), .B(y[5576]), .Z(n44263) );
  NAND U14460 ( .A(n44256), .B(n44263), .Z(n58015) );
  NANDN U14461 ( .A(y[5574]), .B(x[5574]), .Z(n9496) );
  NANDN U14462 ( .A(y[5575]), .B(x[5575]), .Z(n24018) );
  AND U14463 ( .A(n9496), .B(n24018), .Z(n58013) );
  ANDN U14464 ( .B(y[5573]), .A(x[5573]), .Z(n44251) );
  XNOR U14465 ( .A(y[5574]), .B(x[5574]), .Z(n24020) );
  NANDN U14466 ( .A(n44251), .B(n24020), .Z(n58012) );
  XNOR U14467 ( .A(y[5572]), .B(x[5572]), .Z(n24022) );
  NANDN U14468 ( .A(x[5571]), .B(y[5571]), .Z(n24023) );
  AND U14469 ( .A(n24022), .B(n24023), .Z(n58010) );
  NANDN U14470 ( .A(y[5570]), .B(x[5570]), .Z(n24025) );
  NANDN U14471 ( .A(y[5571]), .B(x[5571]), .Z(n24021) );
  NAND U14472 ( .A(n24025), .B(n24021), .Z(n58009) );
  NANDN U14473 ( .A(x[5569]), .B(y[5569]), .Z(n24027) );
  NANDN U14474 ( .A(x[5570]), .B(y[5570]), .Z(n24024) );
  AND U14475 ( .A(n24027), .B(n24024), .Z(n58008) );
  NANDN U14476 ( .A(y[5568]), .B(x[5568]), .Z(n24029) );
  NANDN U14477 ( .A(y[5569]), .B(x[5569]), .Z(n24026) );
  NAND U14478 ( .A(n24029), .B(n24026), .Z(n58007) );
  NANDN U14479 ( .A(x[5567]), .B(y[5567]), .Z(n44237) );
  NANDN U14480 ( .A(x[5568]), .B(y[5568]), .Z(n24028) );
  AND U14481 ( .A(n44237), .B(n24028), .Z(n58006) );
  XNOR U14482 ( .A(x[5566]), .B(y[5566]), .Z(n24032) );
  XNOR U14483 ( .A(x[5564]), .B(y[5564]), .Z(n44230) );
  NANDN U14484 ( .A(y[5562]), .B(x[5562]), .Z(n9497) );
  NANDN U14485 ( .A(y[5563]), .B(x[5563]), .Z(n44229) );
  NAND U14486 ( .A(n9497), .B(n44229), .Z(n57999) );
  XNOR U14487 ( .A(x[5562]), .B(y[5562]), .Z(n24034) );
  ANDN U14488 ( .B(y[5561]), .A(x[5561]), .Z(n57997) );
  NANDN U14489 ( .A(y[5560]), .B(x[5560]), .Z(n9498) );
  NANDN U14490 ( .A(y[5561]), .B(x[5561]), .Z(n24033) );
  AND U14491 ( .A(n9498), .B(n24033), .Z(n57995) );
  XNOR U14492 ( .A(x[5560]), .B(y[5560]), .Z(n44220) );
  ANDN U14493 ( .B(y[5559]), .A(x[5559]), .Z(n44216) );
  ANDN U14494 ( .B(n44220), .A(n44216), .Z(n17809) );
  XNOR U14495 ( .A(x[5558]), .B(y[5558]), .Z(n24036) );
  XNOR U14496 ( .A(x[5556]), .B(y[5556]), .Z(n44209) );
  NANDN U14497 ( .A(y[5554]), .B(x[5554]), .Z(n9499) );
  NANDN U14498 ( .A(y[5555]), .B(x[5555]), .Z(n44208) );
  NAND U14499 ( .A(n9499), .B(n44208), .Z(n57987) );
  XNOR U14500 ( .A(x[5554]), .B(y[5554]), .Z(n24038) );
  ANDN U14501 ( .B(y[5553]), .A(x[5553]), .Z(n57986) );
  NANDN U14502 ( .A(y[5552]), .B(x[5552]), .Z(n9500) );
  NANDN U14503 ( .A(y[5553]), .B(x[5553]), .Z(n24037) );
  AND U14504 ( .A(n9500), .B(n24037), .Z(n57984) );
  XNOR U14505 ( .A(x[5552]), .B(y[5552]), .Z(n44199) );
  ANDN U14506 ( .B(y[5551]), .A(x[5551]), .Z(n44195) );
  ANDN U14507 ( .B(n44199), .A(n44195), .Z(n17795) );
  XNOR U14508 ( .A(x[5550]), .B(y[5550]), .Z(n24040) );
  NANDN U14509 ( .A(y[5548]), .B(x[5548]), .Z(n9501) );
  NANDN U14510 ( .A(y[5549]), .B(x[5549]), .Z(n24039) );
  AND U14511 ( .A(n9501), .B(n24039), .Z(n57979) );
  ANDN U14512 ( .B(y[5547]), .A(x[5547]), .Z(n44184) );
  XNOR U14513 ( .A(x[5548]), .B(y[5548]), .Z(n44188) );
  NANDN U14514 ( .A(y[5546]), .B(x[5546]), .Z(n9502) );
  NANDN U14515 ( .A(y[5547]), .B(x[5547]), .Z(n44187) );
  NAND U14516 ( .A(n9502), .B(n44187), .Z(n51348) );
  XNOR U14517 ( .A(x[5546]), .B(y[5546]), .Z(n24042) );
  NANDN U14518 ( .A(x[5545]), .B(y[5545]), .Z(n51350) );
  NANDN U14519 ( .A(y[5544]), .B(x[5544]), .Z(n24044) );
  NANDN U14520 ( .A(y[5545]), .B(x[5545]), .Z(n24041) );
  AND U14521 ( .A(n24044), .B(n24041), .Z(n57976) );
  NANDN U14522 ( .A(x[5543]), .B(y[5543]), .Z(n24046) );
  NANDN U14523 ( .A(x[5544]), .B(y[5544]), .Z(n24043) );
  NAND U14524 ( .A(n24046), .B(n24043), .Z(n57975) );
  NANDN U14525 ( .A(y[5542]), .B(x[5542]), .Z(n9503) );
  NANDN U14526 ( .A(y[5543]), .B(x[5543]), .Z(n24045) );
  AND U14527 ( .A(n9503), .B(n24045), .Z(n57974) );
  XNOR U14528 ( .A(x[5542]), .B(y[5542]), .Z(n24048) );
  NANDN U14529 ( .A(y[5540]), .B(x[5540]), .Z(n9504) );
  NANDN U14530 ( .A(y[5541]), .B(x[5541]), .Z(n24047) );
  NAND U14531 ( .A(n9504), .B(n24047), .Z(n57971) );
  XNOR U14532 ( .A(y[5540]), .B(x[5540]), .Z(n24050) );
  NANDN U14533 ( .A(x[5539]), .B(y[5539]), .Z(n24051) );
  AND U14534 ( .A(n24050), .B(n24051), .Z(n57969) );
  NANDN U14535 ( .A(y[5538]), .B(x[5538]), .Z(n24053) );
  NANDN U14536 ( .A(y[5539]), .B(x[5539]), .Z(n24049) );
  NAND U14537 ( .A(n24053), .B(n24049), .Z(n57968) );
  NANDN U14538 ( .A(x[5538]), .B(y[5538]), .Z(n24052) );
  ANDN U14539 ( .B(y[5537]), .A(x[5537]), .Z(n24055) );
  ANDN U14540 ( .B(n24052), .A(n24055), .Z(n57967) );
  XNOR U14541 ( .A(x[5536]), .B(y[5536]), .Z(n44160) );
  XNOR U14542 ( .A(x[5534]), .B(y[5534]), .Z(n24057) );
  NANDN U14543 ( .A(y[5532]), .B(x[5532]), .Z(n9505) );
  NANDN U14544 ( .A(y[5533]), .B(x[5533]), .Z(n24056) );
  NAND U14545 ( .A(n9505), .B(n24056), .Z(n57960) );
  XNOR U14546 ( .A(x[5532]), .B(y[5532]), .Z(n24059) );
  NANDN U14547 ( .A(x[5531]), .B(y[5531]), .Z(n57959) );
  NANDN U14548 ( .A(y[5530]), .B(x[5530]), .Z(n9506) );
  NANDN U14549 ( .A(y[5531]), .B(x[5531]), .Z(n24058) );
  AND U14550 ( .A(n9506), .B(n24058), .Z(n57957) );
  XNOR U14551 ( .A(x[5530]), .B(y[5530]), .Z(n24061) );
  NANDN U14552 ( .A(x[5529]), .B(y[5529]), .Z(n51351) );
  AND U14553 ( .A(n24061), .B(n51351), .Z(n17762) );
  NANDN U14554 ( .A(y[5528]), .B(x[5528]), .Z(n24063) );
  NANDN U14555 ( .A(y[5529]), .B(x[5529]), .Z(n24060) );
  AND U14556 ( .A(n24063), .B(n24060), .Z(n57955) );
  NANDN U14557 ( .A(x[5527]), .B(y[5527]), .Z(n44140) );
  NANDN U14558 ( .A(x[5528]), .B(y[5528]), .Z(n24062) );
  NAND U14559 ( .A(n44140), .B(n24062), .Z(n57954) );
  NANDN U14560 ( .A(y[5526]), .B(x[5526]), .Z(n9507) );
  NANDN U14561 ( .A(y[5527]), .B(x[5527]), .Z(n24064) );
  AND U14562 ( .A(n9507), .B(n24064), .Z(n51353) );
  ANDN U14563 ( .B(y[5525]), .A(x[5525]), .Z(n57953) );
  XNOR U14564 ( .A(x[5526]), .B(y[5526]), .Z(n24066) );
  NANDN U14565 ( .A(y[5524]), .B(x[5524]), .Z(n9508) );
  NANDN U14566 ( .A(y[5525]), .B(x[5525]), .Z(n24065) );
  NAND U14567 ( .A(n9508), .B(n24065), .Z(n57951) );
  XNOR U14568 ( .A(x[5524]), .B(y[5524]), .Z(n44133) );
  ANDN U14569 ( .B(y[5523]), .A(x[5523]), .Z(n44129) );
  NANDN U14570 ( .A(x[5521]), .B(y[5521]), .Z(n57948) );
  XNOR U14571 ( .A(x[5522]), .B(y[5522]), .Z(n24068) );
  AND U14572 ( .A(n57948), .B(n24068), .Z(n17750) );
  NANDN U14573 ( .A(y[5520]), .B(x[5520]), .Z(n24069) );
  NANDN U14574 ( .A(y[5521]), .B(x[5521]), .Z(n24067) );
  NAND U14575 ( .A(n24069), .B(n24067), .Z(n57947) );
  NANDN U14576 ( .A(y[5516]), .B(x[5516]), .Z(n24074) );
  NANDN U14577 ( .A(y[5517]), .B(x[5517]), .Z(n24073) );
  NAND U14578 ( .A(n24074), .B(n24073), .Z(n57938) );
  NANDN U14579 ( .A(x[5515]), .B(y[5515]), .Z(n44112) );
  NANDN U14580 ( .A(x[5516]), .B(y[5516]), .Z(n44118) );
  AND U14581 ( .A(n44112), .B(n44118), .Z(n51356) );
  NANDN U14582 ( .A(y[5512]), .B(x[5512]), .Z(n9509) );
  NANDN U14583 ( .A(y[5513]), .B(x[5513]), .Z(n24076) );
  AND U14584 ( .A(n9509), .B(n24076), .Z(n57936) );
  XNOR U14585 ( .A(x[5512]), .B(y[5512]), .Z(n24079) );
  NANDN U14586 ( .A(y[5510]), .B(x[5510]), .Z(n9510) );
  NANDN U14587 ( .A(y[5511]), .B(x[5511]), .Z(n24078) );
  NAND U14588 ( .A(n9510), .B(n24078), .Z(n57935) );
  XNOR U14589 ( .A(y[5510]), .B(x[5510]), .Z(n24082) );
  ANDN U14590 ( .B(y[5509]), .A(x[5509]), .Z(n24083) );
  ANDN U14591 ( .B(n24082), .A(n24083), .Z(n57934) );
  NANDN U14592 ( .A(y[5508]), .B(x[5508]), .Z(n9511) );
  NANDN U14593 ( .A(y[5509]), .B(x[5509]), .Z(n24081) );
  NAND U14594 ( .A(n9511), .B(n24081), .Z(n57933) );
  NANDN U14595 ( .A(y[5506]), .B(x[5506]), .Z(n9512) );
  NANDN U14596 ( .A(y[5507]), .B(x[5507]), .Z(n44095) );
  AND U14597 ( .A(n9512), .B(n44095), .Z(n57929) );
  XNOR U14598 ( .A(x[5506]), .B(y[5506]), .Z(n24085) );
  NANDN U14599 ( .A(y[5504]), .B(x[5504]), .Z(n9513) );
  NANDN U14600 ( .A(y[5505]), .B(x[5505]), .Z(n24084) );
  AND U14601 ( .A(n9513), .B(n24084), .Z(n51361) );
  NANDN U14602 ( .A(x[5503]), .B(y[5503]), .Z(n57926) );
  XNOR U14603 ( .A(x[5504]), .B(y[5504]), .Z(n44086) );
  NANDN U14604 ( .A(y[5502]), .B(x[5502]), .Z(n9514) );
  NANDN U14605 ( .A(y[5503]), .B(x[5503]), .Z(n44085) );
  NAND U14606 ( .A(n9514), .B(n44085), .Z(n57924) );
  XNOR U14607 ( .A(y[5502]), .B(x[5502]), .Z(n24087) );
  NANDN U14608 ( .A(x[5501]), .B(y[5501]), .Z(n24088) );
  AND U14609 ( .A(n24087), .B(n24088), .Z(n51362) );
  NANDN U14610 ( .A(x[5499]), .B(y[5499]), .Z(n57923) );
  XNOR U14611 ( .A(x[5500]), .B(y[5500]), .Z(n24090) );
  AND U14612 ( .A(n57923), .B(n24090), .Z(n17718) );
  NANDN U14613 ( .A(y[5498]), .B(x[5498]), .Z(n9515) );
  NANDN U14614 ( .A(y[5499]), .B(x[5499]), .Z(n24089) );
  NAND U14615 ( .A(n9515), .B(n24089), .Z(n57922) );
  XNOR U14616 ( .A(x[5498]), .B(y[5498]), .Z(n24092) );
  NANDN U14617 ( .A(y[5496]), .B(x[5496]), .Z(n24094) );
  NANDN U14618 ( .A(y[5497]), .B(x[5497]), .Z(n24091) );
  NAND U14619 ( .A(n24094), .B(n24091), .Z(n57917) );
  NANDN U14620 ( .A(x[5495]), .B(y[5495]), .Z(n44065) );
  NANDN U14621 ( .A(x[5496]), .B(y[5496]), .Z(n24093) );
  AND U14622 ( .A(n44065), .B(n24093), .Z(n57916) );
  NANDN U14623 ( .A(y[5494]), .B(x[5494]), .Z(n9516) );
  NANDN U14624 ( .A(y[5495]), .B(x[5495]), .Z(n24095) );
  NAND U14625 ( .A(n9516), .B(n24095), .Z(n57915) );
  XNOR U14626 ( .A(x[5494]), .B(y[5494]), .Z(n24097) );
  ANDN U14627 ( .B(y[5493]), .A(x[5493]), .Z(n57913) );
  ANDN U14628 ( .B(n24097), .A(n57913), .Z(n17710) );
  XNOR U14629 ( .A(x[5492]), .B(y[5492]), .Z(n44058) );
  NANDN U14630 ( .A(y[5490]), .B(x[5490]), .Z(n9517) );
  NANDN U14631 ( .A(y[5491]), .B(x[5491]), .Z(n44057) );
  AND U14632 ( .A(n9517), .B(n44057), .Z(n51365) );
  NANDN U14633 ( .A(x[5489]), .B(y[5489]), .Z(n57909) );
  XNOR U14634 ( .A(x[5490]), .B(y[5490]), .Z(n24099) );
  NANDN U14635 ( .A(y[5488]), .B(x[5488]), .Z(n24100) );
  NANDN U14636 ( .A(y[5489]), .B(x[5489]), .Z(n24098) );
  NAND U14637 ( .A(n24100), .B(n24098), .Z(n57907) );
  NANDN U14638 ( .A(x[5487]), .B(y[5487]), .Z(n44044) );
  NANDN U14639 ( .A(x[5488]), .B(y[5488]), .Z(n44050) );
  AND U14640 ( .A(n44044), .B(n44050), .Z(n57906) );
  NANDN U14641 ( .A(y[5486]), .B(x[5486]), .Z(n9518) );
  NANDN U14642 ( .A(y[5487]), .B(x[5487]), .Z(n24101) );
  NAND U14643 ( .A(n9518), .B(n24101), .Z(n57904) );
  XNOR U14644 ( .A(x[5486]), .B(y[5486]), .Z(n24103) );
  NANDN U14645 ( .A(x[5485]), .B(y[5485]), .Z(n57902) );
  AND U14646 ( .A(n24103), .B(n57902), .Z(n17698) );
  NANDN U14647 ( .A(x[5483]), .B(y[5483]), .Z(n24107) );
  NANDN U14648 ( .A(x[5484]), .B(y[5484]), .Z(n24104) );
  AND U14649 ( .A(n24107), .B(n24104), .Z(n57900) );
  NANDN U14650 ( .A(y[5482]), .B(x[5482]), .Z(n24109) );
  NANDN U14651 ( .A(y[5483]), .B(x[5483]), .Z(n24105) );
  NAND U14652 ( .A(n24109), .B(n24105), .Z(n57899) );
  NANDN U14653 ( .A(x[5481]), .B(y[5481]), .Z(n24111) );
  NANDN U14654 ( .A(x[5482]), .B(y[5482]), .Z(n24108) );
  AND U14655 ( .A(n24111), .B(n24108), .Z(n51366) );
  XNOR U14656 ( .A(x[5478]), .B(y[5478]), .Z(n24117) );
  NANDN U14657 ( .A(y[5476]), .B(x[5476]), .Z(n24118) );
  NANDN U14658 ( .A(y[5477]), .B(x[5477]), .Z(n24116) );
  NAND U14659 ( .A(n24118), .B(n24116), .Z(n57894) );
  NANDN U14660 ( .A(x[5475]), .B(y[5475]), .Z(n24120) );
  NANDN U14661 ( .A(x[5476]), .B(y[5476]), .Z(n44024) );
  AND U14662 ( .A(n24120), .B(n44024), .Z(n51368) );
  NANDN U14663 ( .A(x[5474]), .B(y[5474]), .Z(n24121) );
  ANDN U14664 ( .B(y[5473]), .A(x[5473]), .Z(n24124) );
  ANDN U14665 ( .B(n24121), .A(n24124), .Z(n57891) );
  XNOR U14666 ( .A(x[5472]), .B(y[5472]), .Z(n44012) );
  XNOR U14667 ( .A(x[5470]), .B(y[5470]), .Z(n24126) );
  NANDN U14668 ( .A(y[5468]), .B(x[5468]), .Z(n9519) );
  NANDN U14669 ( .A(y[5469]), .B(x[5469]), .Z(n24125) );
  NAND U14670 ( .A(n9519), .B(n24125), .Z(n57886) );
  XNOR U14671 ( .A(x[5468]), .B(y[5468]), .Z(n44002) );
  ANDN U14672 ( .B(y[5467]), .A(x[5467]), .Z(n43997) );
  XNOR U14673 ( .A(y[5466]), .B(x[5466]), .Z(n24129) );
  NANDN U14674 ( .A(x[5465]), .B(y[5465]), .Z(n24130) );
  AND U14675 ( .A(n24129), .B(n24130), .Z(n57883) );
  XNOR U14676 ( .A(x[5464]), .B(y[5464]), .Z(n24132) );
  XNOR U14677 ( .A(y[5462]), .B(x[5462]), .Z(n24135) );
  ANDN U14678 ( .B(y[5461]), .A(x[5461]), .Z(n24136) );
  ANDN U14679 ( .B(n24135), .A(n24136), .Z(n57879) );
  NANDN U14680 ( .A(y[5460]), .B(x[5460]), .Z(n9520) );
  NANDN U14681 ( .A(y[5461]), .B(x[5461]), .Z(n24134) );
  NAND U14682 ( .A(n9520), .B(n24134), .Z(n57878) );
  XNOR U14683 ( .A(x[5460]), .B(y[5460]), .Z(n43982) );
  NANDN U14684 ( .A(x[5459]), .B(y[5459]), .Z(n57877) );
  NANDN U14685 ( .A(y[5458]), .B(x[5458]), .Z(n9521) );
  NANDN U14686 ( .A(y[5459]), .B(x[5459]), .Z(n43981) );
  AND U14687 ( .A(n9521), .B(n43981), .Z(n57875) );
  XNOR U14688 ( .A(x[5458]), .B(y[5458]), .Z(n24138) );
  ANDN U14689 ( .B(y[5457]), .A(x[5457]), .Z(n51375) );
  ANDN U14690 ( .B(n24138), .A(n51375), .Z(n17657) );
  NANDN U14691 ( .A(y[5456]), .B(x[5456]), .Z(n9522) );
  NANDN U14692 ( .A(y[5457]), .B(x[5457]), .Z(n24137) );
  NAND U14693 ( .A(n9522), .B(n24137), .Z(n57874) );
  XNOR U14694 ( .A(x[5456]), .B(y[5456]), .Z(n43972) );
  NANDN U14695 ( .A(y[5454]), .B(x[5454]), .Z(n9523) );
  NANDN U14696 ( .A(y[5455]), .B(x[5455]), .Z(n43971) );
  NAND U14697 ( .A(n9523), .B(n43971), .Z(n57871) );
  XNOR U14698 ( .A(x[5454]), .B(y[5454]), .Z(n24140) );
  NANDN U14699 ( .A(y[5452]), .B(x[5452]), .Z(n9524) );
  NANDN U14700 ( .A(y[5453]), .B(x[5453]), .Z(n24139) );
  NAND U14701 ( .A(n9524), .B(n24139), .Z(n57868) );
  NANDN U14702 ( .A(x[5451]), .B(y[5451]), .Z(n57865) );
  XNOR U14703 ( .A(x[5452]), .B(y[5452]), .Z(n24142) );
  NANDN U14704 ( .A(y[5450]), .B(x[5450]), .Z(n9525) );
  NANDN U14705 ( .A(y[5451]), .B(x[5451]), .Z(n24141) );
  AND U14706 ( .A(n9525), .B(n24141), .Z(n57864) );
  XNOR U14707 ( .A(x[5450]), .B(y[5450]), .Z(n24144) );
  ANDN U14708 ( .B(y[5449]), .A(x[5449]), .Z(n51377) );
  ANDN U14709 ( .B(n24144), .A(n51377), .Z(n17645) );
  NANDN U14710 ( .A(y[5448]), .B(x[5448]), .Z(n9526) );
  NANDN U14711 ( .A(y[5449]), .B(x[5449]), .Z(n24143) );
  NAND U14712 ( .A(n9526), .B(n24143), .Z(n57862) );
  XNOR U14713 ( .A(x[5448]), .B(y[5448]), .Z(n43954) );
  NANDN U14714 ( .A(y[5446]), .B(x[5446]), .Z(n9527) );
  NANDN U14715 ( .A(y[5447]), .B(x[5447]), .Z(n43953) );
  NAND U14716 ( .A(n9527), .B(n43953), .Z(n57859) );
  ANDN U14717 ( .B(y[5445]), .A(x[5445]), .Z(n57857) );
  XNOR U14718 ( .A(x[5446]), .B(y[5446]), .Z(n24146) );
  NANDN U14719 ( .A(y[5444]), .B(x[5444]), .Z(n9528) );
  NANDN U14720 ( .A(y[5445]), .B(x[5445]), .Z(n24145) );
  NAND U14721 ( .A(n9528), .B(n24145), .Z(n57856) );
  XNOR U14722 ( .A(x[5444]), .B(y[5444]), .Z(n43944) );
  NANDN U14723 ( .A(x[5443]), .B(y[5443]), .Z(n57855) );
  NANDN U14724 ( .A(y[5442]), .B(x[5442]), .Z(n9529) );
  NANDN U14725 ( .A(y[5443]), .B(x[5443]), .Z(n43943) );
  AND U14726 ( .A(n9529), .B(n43943), .Z(n57853) );
  XNOR U14727 ( .A(x[5442]), .B(y[5442]), .Z(n24148) );
  ANDN U14728 ( .B(y[5441]), .A(x[5441]), .Z(n51379) );
  ANDN U14729 ( .B(n24148), .A(n51379), .Z(n17633) );
  NANDN U14730 ( .A(y[5440]), .B(x[5440]), .Z(n9530) );
  NANDN U14731 ( .A(y[5441]), .B(x[5441]), .Z(n24147) );
  NAND U14732 ( .A(n9530), .B(n24147), .Z(n57852) );
  XNOR U14733 ( .A(x[5440]), .B(y[5440]), .Z(n43934) );
  NANDN U14734 ( .A(y[5438]), .B(x[5438]), .Z(n9531) );
  NANDN U14735 ( .A(y[5439]), .B(x[5439]), .Z(n43933) );
  NAND U14736 ( .A(n9531), .B(n43933), .Z(n57848) );
  ANDN U14737 ( .B(y[5437]), .A(x[5437]), .Z(n57846) );
  XNOR U14738 ( .A(x[5438]), .B(y[5438]), .Z(n24150) );
  NANDN U14739 ( .A(y[5436]), .B(x[5436]), .Z(n9532) );
  NANDN U14740 ( .A(y[5437]), .B(x[5437]), .Z(n24149) );
  NAND U14741 ( .A(n9532), .B(n24149), .Z(n57845) );
  XNOR U14742 ( .A(x[5436]), .B(y[5436]), .Z(n43924) );
  NANDN U14743 ( .A(x[5435]), .B(y[5435]), .Z(n57844) );
  NANDN U14744 ( .A(y[5434]), .B(x[5434]), .Z(n9533) );
  NANDN U14745 ( .A(y[5435]), .B(x[5435]), .Z(n43923) );
  AND U14746 ( .A(n9533), .B(n43923), .Z(n57842) );
  XNOR U14747 ( .A(x[5434]), .B(y[5434]), .Z(n24152) );
  ANDN U14748 ( .B(y[5433]), .A(x[5433]), .Z(n51381) );
  ANDN U14749 ( .B(n24152), .A(n51381), .Z(n17621) );
  NANDN U14750 ( .A(y[5432]), .B(x[5432]), .Z(n9534) );
  NANDN U14751 ( .A(y[5433]), .B(x[5433]), .Z(n24151) );
  NAND U14752 ( .A(n9534), .B(n24151), .Z(n57841) );
  XNOR U14753 ( .A(x[5432]), .B(y[5432]), .Z(n43914) );
  NANDN U14754 ( .A(y[5430]), .B(x[5430]), .Z(n9535) );
  NANDN U14755 ( .A(y[5431]), .B(x[5431]), .Z(n43913) );
  NAND U14756 ( .A(n9535), .B(n43913), .Z(n57838) );
  XNOR U14757 ( .A(x[5430]), .B(y[5430]), .Z(n24154) );
  NANDN U14758 ( .A(y[5428]), .B(x[5428]), .Z(n9536) );
  NANDN U14759 ( .A(y[5429]), .B(x[5429]), .Z(n24153) );
  NAND U14760 ( .A(n9536), .B(n24153), .Z(n57835) );
  XNOR U14761 ( .A(x[5428]), .B(y[5428]), .Z(n24156) );
  ANDN U14762 ( .B(y[5427]), .A(x[5427]), .Z(n43902) );
  NANDN U14763 ( .A(y[5426]), .B(x[5426]), .Z(n9537) );
  NANDN U14764 ( .A(y[5427]), .B(x[5427]), .Z(n24155) );
  AND U14765 ( .A(n9537), .B(n24155), .Z(n57832) );
  NANDN U14766 ( .A(x[5425]), .B(y[5425]), .Z(n51383) );
  XNOR U14767 ( .A(x[5426]), .B(y[5426]), .Z(n24158) );
  AND U14768 ( .A(n51383), .B(n24158), .Z(n17609) );
  NANDN U14769 ( .A(y[5424]), .B(x[5424]), .Z(n9538) );
  NANDN U14770 ( .A(y[5425]), .B(x[5425]), .Z(n24157) );
  NAND U14771 ( .A(n9538), .B(n24157), .Z(n57829) );
  ANDN U14772 ( .B(x[5423]), .A(y[5423]), .Z(n43897) );
  NANDN U14773 ( .A(y[5422]), .B(x[5422]), .Z(n9539) );
  NANDN U14774 ( .A(n43897), .B(n9539), .Z(n51385) );
  ANDN U14775 ( .B(y[5421]), .A(x[5421]), .Z(n57825) );
  XNOR U14776 ( .A(x[5422]), .B(y[5422]), .Z(n24160) );
  NANDN U14777 ( .A(y[5420]), .B(x[5420]), .Z(n9540) );
  NANDN U14778 ( .A(y[5421]), .B(x[5421]), .Z(n24159) );
  NAND U14779 ( .A(n9540), .B(n24159), .Z(n57824) );
  XNOR U14780 ( .A(x[5420]), .B(y[5420]), .Z(n43885) );
  NANDN U14781 ( .A(x[5419]), .B(y[5419]), .Z(n57823) );
  NANDN U14782 ( .A(y[5418]), .B(x[5418]), .Z(n9541) );
  NANDN U14783 ( .A(y[5419]), .B(x[5419]), .Z(n43884) );
  AND U14784 ( .A(n9541), .B(n43884), .Z(n57821) );
  XNOR U14785 ( .A(x[5418]), .B(y[5418]), .Z(n24162) );
  ANDN U14786 ( .B(y[5417]), .A(x[5417]), .Z(n51386) );
  ANDN U14787 ( .B(n24162), .A(n51386), .Z(n17597) );
  NANDN U14788 ( .A(y[5416]), .B(x[5416]), .Z(n9542) );
  NANDN U14789 ( .A(y[5417]), .B(x[5417]), .Z(n24161) );
  NAND U14790 ( .A(n9542), .B(n24161), .Z(n57820) );
  XNOR U14791 ( .A(x[5416]), .B(y[5416]), .Z(n43875) );
  NANDN U14792 ( .A(y[5414]), .B(x[5414]), .Z(n9543) );
  NANDN U14793 ( .A(y[5415]), .B(x[5415]), .Z(n43874) );
  NAND U14794 ( .A(n9543), .B(n43874), .Z(n51388) );
  ANDN U14795 ( .B(y[5413]), .A(x[5413]), .Z(n57813) );
  XNOR U14796 ( .A(x[5414]), .B(y[5414]), .Z(n24164) );
  NANDN U14797 ( .A(y[5412]), .B(x[5412]), .Z(n9544) );
  NANDN U14798 ( .A(y[5413]), .B(x[5413]), .Z(n24163) );
  NAND U14799 ( .A(n9544), .B(n24163), .Z(n57812) );
  XNOR U14800 ( .A(x[5412]), .B(y[5412]), .Z(n43865) );
  NANDN U14801 ( .A(x[5411]), .B(y[5411]), .Z(n57810) );
  AND U14802 ( .A(n43865), .B(n57810), .Z(n17588) );
  NANDN U14803 ( .A(y[5408]), .B(x[5408]), .Z(n9545) );
  NANDN U14804 ( .A(y[5409]), .B(x[5409]), .Z(n24165) );
  AND U14805 ( .A(n9545), .B(n24165), .Z(n57808) );
  XNOR U14806 ( .A(x[5408]), .B(y[5408]), .Z(n43855) );
  XNOR U14807 ( .A(x[5406]), .B(y[5406]), .Z(n24168) );
  NANDN U14808 ( .A(y[5404]), .B(x[5404]), .Z(n9546) );
  NANDN U14809 ( .A(y[5405]), .B(x[5405]), .Z(n24167) );
  NAND U14810 ( .A(n9546), .B(n24167), .Z(n57801) );
  XNOR U14811 ( .A(x[5404]), .B(y[5404]), .Z(n43844) );
  NANDN U14812 ( .A(x[5403]), .B(y[5403]), .Z(n57799) );
  AND U14813 ( .A(n43844), .B(n57799), .Z(n17574) );
  NANDN U14814 ( .A(x[5401]), .B(y[5401]), .Z(n24172) );
  NANDN U14815 ( .A(x[5402]), .B(y[5402]), .Z(n24169) );
  AND U14816 ( .A(n24172), .B(n24169), .Z(n57797) );
  XNOR U14817 ( .A(x[5400]), .B(y[5400]), .Z(n24174) );
  XNOR U14818 ( .A(x[5398]), .B(y[5398]), .Z(n24176) );
  NANDN U14819 ( .A(y[5396]), .B(x[5396]), .Z(n9547) );
  NANDN U14820 ( .A(y[5397]), .B(x[5397]), .Z(n24175) );
  NAND U14821 ( .A(n9547), .B(n24175), .Z(n57790) );
  XNOR U14822 ( .A(x[5396]), .B(y[5396]), .Z(n24178) );
  NANDN U14823 ( .A(x[5395]), .B(y[5395]), .Z(n57789) );
  NANDN U14824 ( .A(y[5394]), .B(x[5394]), .Z(n9548) );
  NANDN U14825 ( .A(y[5395]), .B(x[5395]), .Z(n24177) );
  AND U14826 ( .A(n9548), .B(n24177), .Z(n57787) );
  ANDN U14827 ( .B(y[5393]), .A(x[5393]), .Z(n51391) );
  NANDN U14828 ( .A(y[5392]), .B(x[5392]), .Z(n9549) );
  NANDN U14829 ( .A(y[5393]), .B(x[5393]), .Z(n24179) );
  AND U14830 ( .A(n9549), .B(n24179), .Z(n57785) );
  XNOR U14831 ( .A(x[5392]), .B(y[5392]), .Z(n43818) );
  XNOR U14832 ( .A(x[5390]), .B(y[5390]), .Z(n24182) );
  NANDN U14833 ( .A(y[5388]), .B(x[5388]), .Z(n9550) );
  NANDN U14834 ( .A(y[5389]), .B(x[5389]), .Z(n24181) );
  NAND U14835 ( .A(n9550), .B(n24181), .Z(n57779) );
  XNOR U14836 ( .A(x[5388]), .B(y[5388]), .Z(n43807) );
  NANDN U14837 ( .A(x[5387]), .B(y[5387]), .Z(n57778) );
  NANDN U14838 ( .A(y[5386]), .B(x[5386]), .Z(n9551) );
  NANDN U14839 ( .A(y[5387]), .B(x[5387]), .Z(n43806) );
  AND U14840 ( .A(n9551), .B(n43806), .Z(n57776) );
  XNOR U14841 ( .A(y[5386]), .B(x[5386]), .Z(n24184) );
  ANDN U14842 ( .B(y[5385]), .A(x[5385]), .Z(n24185) );
  ANDN U14843 ( .B(n24184), .A(n24185), .Z(n57775) );
  XNOR U14844 ( .A(x[5384]), .B(y[5384]), .Z(n43796) );
  NANDN U14845 ( .A(y[5382]), .B(x[5382]), .Z(n9552) );
  NANDN U14846 ( .A(y[5383]), .B(x[5383]), .Z(n43795) );
  NAND U14847 ( .A(n9552), .B(n43795), .Z(n57772) );
  NANDN U14848 ( .A(x[5381]), .B(y[5381]), .Z(n57770) );
  XNOR U14849 ( .A(x[5382]), .B(y[5382]), .Z(n24187) );
  NANDN U14850 ( .A(y[5380]), .B(x[5380]), .Z(n9553) );
  NANDN U14851 ( .A(y[5381]), .B(x[5381]), .Z(n24186) );
  NAND U14852 ( .A(n9553), .B(n24186), .Z(n57766) );
  NANDN U14853 ( .A(x[5379]), .B(y[5379]), .Z(n51395) );
  XNOR U14854 ( .A(x[5380]), .B(y[5380]), .Z(n43786) );
  NANDN U14855 ( .A(y[5378]), .B(x[5378]), .Z(n24189) );
  NANDN U14856 ( .A(y[5379]), .B(x[5379]), .Z(n43785) );
  AND U14857 ( .A(n24189), .B(n43785), .Z(n57765) );
  NANDN U14858 ( .A(x[5377]), .B(y[5377]), .Z(n24191) );
  NANDN U14859 ( .A(x[5378]), .B(y[5378]), .Z(n24188) );
  NAND U14860 ( .A(n24191), .B(n24188), .Z(n57764) );
  NANDN U14861 ( .A(y[5376]), .B(x[5376]), .Z(n9554) );
  NANDN U14862 ( .A(y[5377]), .B(x[5377]), .Z(n24190) );
  AND U14863 ( .A(n9554), .B(n24190), .Z(n51397) );
  NANDN U14864 ( .A(x[5375]), .B(y[5375]), .Z(n57763) );
  XNOR U14865 ( .A(x[5376]), .B(y[5376]), .Z(n24193) );
  NANDN U14866 ( .A(y[5374]), .B(x[5374]), .Z(n9555) );
  NANDN U14867 ( .A(y[5375]), .B(x[5375]), .Z(n24192) );
  NAND U14868 ( .A(n9555), .B(n24192), .Z(n57761) );
  XNOR U14869 ( .A(x[5374]), .B(y[5374]), .Z(n24195) );
  ANDN U14870 ( .B(y[5373]), .A(x[5373]), .Z(n51398) );
  NANDN U14871 ( .A(x[5371]), .B(y[5371]), .Z(n57758) );
  XNOR U14872 ( .A(x[5372]), .B(y[5372]), .Z(n43768) );
  AND U14873 ( .A(n57758), .B(n43768), .Z(n17524) );
  NANDN U14874 ( .A(y[5370]), .B(x[5370]), .Z(n9556) );
  NANDN U14875 ( .A(y[5371]), .B(x[5371]), .Z(n43767) );
  NAND U14876 ( .A(n9556), .B(n43767), .Z(n57756) );
  XNOR U14877 ( .A(y[5370]), .B(x[5370]), .Z(n24197) );
  NANDN U14878 ( .A(x[5369]), .B(y[5369]), .Z(n24198) );
  AND U14879 ( .A(n24197), .B(n24198), .Z(n57755) );
  NANDN U14880 ( .A(y[5368]), .B(x[5368]), .Z(n9557) );
  NANDN U14881 ( .A(y[5369]), .B(x[5369]), .Z(n24196) );
  NAND U14882 ( .A(n9557), .B(n24196), .Z(n57754) );
  XNOR U14883 ( .A(y[5368]), .B(x[5368]), .Z(n24201) );
  NANDN U14884 ( .A(x[5367]), .B(y[5367]), .Z(n24202) );
  AND U14885 ( .A(n24201), .B(n24202), .Z(n51400) );
  XNOR U14886 ( .A(y[5366]), .B(x[5366]), .Z(n24205) );
  ANDN U14887 ( .B(y[5365]), .A(x[5365]), .Z(n24206) );
  ANDN U14888 ( .B(n24205), .A(n24206), .Z(n57753) );
  XNOR U14889 ( .A(x[5364]), .B(y[5364]), .Z(n43749) );
  XNOR U14890 ( .A(x[5362]), .B(y[5362]), .Z(n24208) );
  NANDN U14891 ( .A(y[5360]), .B(x[5360]), .Z(n9558) );
  NANDN U14892 ( .A(y[5361]), .B(x[5361]), .Z(n24207) );
  NAND U14893 ( .A(n9558), .B(n24207), .Z(n57747) );
  XNOR U14894 ( .A(x[5360]), .B(y[5360]), .Z(n43739) );
  ANDN U14895 ( .B(y[5359]), .A(x[5359]), .Z(n43735) );
  XNOR U14896 ( .A(x[5358]), .B(y[5358]), .Z(n24211) );
  ANDN U14897 ( .B(y[5357]), .A(x[5357]), .Z(n57743) );
  ANDN U14898 ( .B(n24211), .A(n57743), .Z(n17502) );
  NANDN U14899 ( .A(y[5354]), .B(x[5354]), .Z(n24216) );
  NANDN U14900 ( .A(y[5355]), .B(x[5355]), .Z(n24213) );
  NAND U14901 ( .A(n24216), .B(n24213), .Z(n51407) );
  NANDN U14902 ( .A(x[5354]), .B(y[5354]), .Z(n24215) );
  ANDN U14903 ( .B(y[5353]), .A(x[5353]), .Z(n24218) );
  ANDN U14904 ( .B(n24215), .A(n24218), .Z(n57741) );
  XNOR U14905 ( .A(x[5352]), .B(y[5352]), .Z(n43719) );
  NANDN U14906 ( .A(x[5351]), .B(y[5351]), .Z(n57738) );
  AND U14907 ( .A(n43719), .B(n57738), .Z(n17494) );
  XNOR U14908 ( .A(x[5350]), .B(y[5350]), .Z(n24220) );
  NANDN U14909 ( .A(y[5348]), .B(x[5348]), .Z(n9559) );
  NANDN U14910 ( .A(y[5349]), .B(x[5349]), .Z(n24219) );
  NAND U14911 ( .A(n9559), .B(n24219), .Z(n51409) );
  XNOR U14912 ( .A(y[5348]), .B(x[5348]), .Z(n24223) );
  NANDN U14913 ( .A(x[5347]), .B(y[5347]), .Z(n24224) );
  AND U14914 ( .A(n24223), .B(n24224), .Z(n57733) );
  NANDN U14915 ( .A(y[5342]), .B(x[5342]), .Z(n9560) );
  NANDN U14916 ( .A(y[5343]), .B(x[5343]), .Z(n24230) );
  NAND U14917 ( .A(n9560), .B(n24230), .Z(n51411) );
  XNOR U14918 ( .A(y[5342]), .B(x[5342]), .Z(n24235) );
  ANDN U14919 ( .B(y[5341]), .A(x[5341]), .Z(n24236) );
  ANDN U14920 ( .B(n24235), .A(n24236), .Z(n57729) );
  XNOR U14921 ( .A(x[5340]), .B(y[5340]), .Z(n43693) );
  NANDN U14922 ( .A(x[5339]), .B(y[5339]), .Z(n57725) );
  AND U14923 ( .A(n43693), .B(n57725), .Z(n17476) );
  NANDN U14924 ( .A(y[5336]), .B(x[5336]), .Z(n9561) );
  NANDN U14925 ( .A(y[5337]), .B(x[5337]), .Z(n24239) );
  AND U14926 ( .A(n9561), .B(n24239), .Z(n57721) );
  XNOR U14927 ( .A(x[5336]), .B(y[5336]), .Z(n24242) );
  ANDN U14928 ( .B(y[5335]), .A(x[5335]), .Z(n24243) );
  ANDN U14929 ( .B(n24242), .A(n24243), .Z(n17471) );
  XNOR U14930 ( .A(x[5334]), .B(y[5334]), .Z(n24245) );
  NANDN U14931 ( .A(x[5333]), .B(y[5333]), .Z(n57719) );
  AND U14932 ( .A(n24245), .B(n57719), .Z(n17467) );
  NANDN U14933 ( .A(y[5332]), .B(x[5332]), .Z(n24247) );
  NANDN U14934 ( .A(y[5333]), .B(x[5333]), .Z(n24244) );
  AND U14935 ( .A(n24247), .B(n24244), .Z(n57717) );
  ANDN U14936 ( .B(y[5329]), .A(x[5329]), .Z(n57713) );
  XNOR U14937 ( .A(x[5330]), .B(y[5330]), .Z(n24250) );
  NANDN U14938 ( .A(y[5328]), .B(x[5328]), .Z(n9562) );
  NANDN U14939 ( .A(y[5329]), .B(x[5329]), .Z(n24249) );
  NAND U14940 ( .A(n9562), .B(n24249), .Z(n57712) );
  XNOR U14941 ( .A(x[5328]), .B(y[5328]), .Z(n43666) );
  NANDN U14942 ( .A(y[5326]), .B(x[5326]), .Z(n9563) );
  NANDN U14943 ( .A(y[5327]), .B(x[5327]), .Z(n43665) );
  NAND U14944 ( .A(n9563), .B(n43665), .Z(n57707) );
  XNOR U14945 ( .A(x[5326]), .B(y[5326]), .Z(n24252) );
  ANDN U14946 ( .B(y[5325]), .A(x[5325]), .Z(n57706) );
  NANDN U14947 ( .A(y[5324]), .B(x[5324]), .Z(n9564) );
  NANDN U14948 ( .A(y[5325]), .B(x[5325]), .Z(n24251) );
  AND U14949 ( .A(n9564), .B(n24251), .Z(n57704) );
  NANDN U14950 ( .A(x[5323]), .B(y[5323]), .Z(n51416) );
  NANDN U14951 ( .A(y[5322]), .B(x[5322]), .Z(n9565) );
  NANDN U14952 ( .A(y[5323]), .B(x[5323]), .Z(n43655) );
  AND U14953 ( .A(n9565), .B(n43655), .Z(n57703) );
  XNOR U14954 ( .A(x[5322]), .B(y[5322]), .Z(n24254) );
  ANDN U14955 ( .B(y[5321]), .A(x[5321]), .Z(n24255) );
  NANDN U14956 ( .A(x[5319]), .B(y[5319]), .Z(n43643) );
  NANDN U14957 ( .A(x[5320]), .B(y[5320]), .Z(n43649) );
  AND U14958 ( .A(n43643), .B(n43649), .Z(n57700) );
  NANDN U14959 ( .A(y[5318]), .B(x[5318]), .Z(n9566) );
  NANDN U14960 ( .A(y[5319]), .B(x[5319]), .Z(n24257) );
  NAND U14961 ( .A(n9566), .B(n24257), .Z(n57699) );
  XNOR U14962 ( .A(x[5318]), .B(y[5318]), .Z(n24259) );
  ANDN U14963 ( .B(y[5317]), .A(x[5317]), .Z(n24260) );
  XNOR U14964 ( .A(x[5316]), .B(y[5316]), .Z(n24262) );
  ANDN U14965 ( .B(y[5315]), .A(x[5315]), .Z(n24263) );
  NANDN U14966 ( .A(x[5313]), .B(y[5313]), .Z(n24267) );
  NANDN U14967 ( .A(x[5314]), .B(y[5314]), .Z(n24264) );
  AND U14968 ( .A(n24267), .B(n24264), .Z(n57694) );
  NANDN U14969 ( .A(y[5312]), .B(x[5312]), .Z(n9567) );
  NANDN U14970 ( .A(y[5313]), .B(x[5313]), .Z(n24266) );
  NAND U14971 ( .A(n9567), .B(n24266), .Z(n57693) );
  NANDN U14972 ( .A(x[5311]), .B(y[5311]), .Z(n51421) );
  XOR U14973 ( .A(x[5312]), .B(y[5312]), .Z(n43630) );
  ANDN U14974 ( .B(x[5311]), .A(y[5311]), .Z(n43628) );
  NANDN U14975 ( .A(y[5310]), .B(x[5310]), .Z(n24269) );
  NANDN U14976 ( .A(n43628), .B(n24269), .Z(n57692) );
  NANDN U14977 ( .A(x[5309]), .B(y[5309]), .Z(n24271) );
  NANDN U14978 ( .A(x[5310]), .B(y[5310]), .Z(n24268) );
  AND U14979 ( .A(n24271), .B(n24268), .Z(n57691) );
  XNOR U14980 ( .A(x[5308]), .B(y[5308]), .Z(n24273) );
  XNOR U14981 ( .A(x[5306]), .B(y[5306]), .Z(n24275) );
  NANDN U14982 ( .A(y[5304]), .B(x[5304]), .Z(n9568) );
  NANDN U14983 ( .A(y[5305]), .B(x[5305]), .Z(n24274) );
  NAND U14984 ( .A(n9568), .B(n24274), .Z(n57687) );
  XNOR U14985 ( .A(x[5304]), .B(y[5304]), .Z(n43610) );
  ANDN U14986 ( .B(y[5303]), .A(x[5303]), .Z(n24276) );
  ANDN U14987 ( .B(y[5301]), .A(x[5301]), .Z(n24280) );
  NANDN U14988 ( .A(x[5302]), .B(y[5302]), .Z(n24277) );
  NANDN U14989 ( .A(n24280), .B(n24277), .Z(n57683) );
  NANDN U14990 ( .A(y[5300]), .B(x[5300]), .Z(n9569) );
  NANDN U14991 ( .A(y[5301]), .B(x[5301]), .Z(n24279) );
  AND U14992 ( .A(n9569), .B(n24279), .Z(n57682) );
  XNOR U14993 ( .A(x[5300]), .B(y[5300]), .Z(n43600) );
  NANDN U14994 ( .A(y[5298]), .B(x[5298]), .Z(n24283) );
  NANDN U14995 ( .A(y[5299]), .B(x[5299]), .Z(n43599) );
  NAND U14996 ( .A(n24283), .B(n43599), .Z(n57681) );
  NANDN U14997 ( .A(x[5297]), .B(y[5297]), .Z(n24285) );
  NANDN U14998 ( .A(x[5298]), .B(y[5298]), .Z(n24282) );
  AND U14999 ( .A(n24285), .B(n24282), .Z(n57680) );
  NANDN U15000 ( .A(y[5296]), .B(x[5296]), .Z(n24287) );
  NANDN U15001 ( .A(y[5297]), .B(x[5297]), .Z(n24284) );
  NAND U15002 ( .A(n24287), .B(n24284), .Z(n57679) );
  NANDN U15003 ( .A(x[5295]), .B(y[5295]), .Z(n24289) );
  NANDN U15004 ( .A(x[5296]), .B(y[5296]), .Z(n24286) );
  AND U15005 ( .A(n24289), .B(n24286), .Z(n57678) );
  NANDN U15006 ( .A(x[5293]), .B(y[5293]), .Z(n24293) );
  NANDN U15007 ( .A(x[5294]), .B(y[5294]), .Z(n24290) );
  AND U15008 ( .A(n24293), .B(n24290), .Z(n57676) );
  NANDN U15009 ( .A(y[5292]), .B(x[5292]), .Z(n9570) );
  NANDN U15010 ( .A(y[5293]), .B(x[5293]), .Z(n24292) );
  NAND U15011 ( .A(n9570), .B(n24292), .Z(n57675) );
  NANDN U15012 ( .A(x[5291]), .B(y[5291]), .Z(n57673) );
  NANDN U15013 ( .A(x[5290]), .B(y[5290]), .Z(n24296) );
  ANDN U15014 ( .B(y[5289]), .A(x[5289]), .Z(n43576) );
  ANDN U15015 ( .B(n24296), .A(n43576), .Z(n57671) );
  NANDN U15016 ( .A(y[5286]), .B(x[5286]), .Z(n24303) );
  NANDN U15017 ( .A(y[5287]), .B(x[5287]), .Z(n24300) );
  NAND U15018 ( .A(n24303), .B(n24300), .Z(n51430) );
  NANDN U15019 ( .A(x[5286]), .B(y[5286]), .Z(n24302) );
  ANDN U15020 ( .B(y[5285]), .A(x[5285]), .Z(n24305) );
  ANDN U15021 ( .B(n24302), .A(n24305), .Z(n57666) );
  XNOR U15022 ( .A(x[5284]), .B(y[5284]), .Z(n43564) );
  NANDN U15023 ( .A(x[5283]), .B(y[5283]), .Z(n57664) );
  NANDN U15024 ( .A(y[5280]), .B(x[5280]), .Z(n24311) );
  NANDN U15025 ( .A(y[5281]), .B(x[5281]), .Z(n24308) );
  NAND U15026 ( .A(n24311), .B(n24308), .Z(n51432) );
  NANDN U15027 ( .A(x[5279]), .B(y[5279]), .Z(n43552) );
  NANDN U15028 ( .A(x[5280]), .B(y[5280]), .Z(n24310) );
  AND U15029 ( .A(n43552), .B(n24310), .Z(n57661) );
  NANDN U15030 ( .A(x[5277]), .B(y[5277]), .Z(n57658) );
  XNOR U15031 ( .A(x[5278]), .B(y[5278]), .Z(n24314) );
  AND U15032 ( .A(n57658), .B(n24314), .Z(n17424) );
  NANDN U15033 ( .A(y[5274]), .B(x[5274]), .Z(n24320) );
  NANDN U15034 ( .A(y[5275]), .B(x[5275]), .Z(n24317) );
  NAND U15035 ( .A(n24320), .B(n24317), .Z(n51434) );
  NANDN U15036 ( .A(x[5273]), .B(y[5273]), .Z(n24322) );
  NANDN U15037 ( .A(x[5274]), .B(y[5274]), .Z(n24319) );
  AND U15038 ( .A(n24322), .B(n24319), .Z(n57653) );
  NANDN U15039 ( .A(x[5271]), .B(y[5271]), .Z(n57650) );
  XOR U15040 ( .A(x[5272]), .B(y[5272]), .Z(n43539) );
  ANDN U15041 ( .B(n57650), .A(n43539), .Z(n17416) );
  NANDN U15042 ( .A(y[5268]), .B(x[5268]), .Z(n24327) );
  NANDN U15043 ( .A(y[5269]), .B(x[5269]), .Z(n24323) );
  NAND U15044 ( .A(n24327), .B(n24323), .Z(n51436) );
  NANDN U15045 ( .A(x[5267]), .B(y[5267]), .Z(n24329) );
  NANDN U15046 ( .A(x[5268]), .B(y[5268]), .Z(n24326) );
  AND U15047 ( .A(n24329), .B(n24326), .Z(n57648) );
  NANDN U15048 ( .A(y[5264]), .B(x[5264]), .Z(n9571) );
  NANDN U15049 ( .A(y[5265]), .B(x[5265]), .Z(n24330) );
  AND U15050 ( .A(n9571), .B(n24330), .Z(n57641) );
  XNOR U15051 ( .A(x[5264]), .B(y[5264]), .Z(n43518) );
  NANDN U15052 ( .A(y[5262]), .B(x[5262]), .Z(n9572) );
  NANDN U15053 ( .A(y[5263]), .B(x[5263]), .Z(n43517) );
  AND U15054 ( .A(n9572), .B(n43517), .Z(n57640) );
  ANDN U15055 ( .B(y[5261]), .A(x[5261]), .Z(n57638) );
  XNOR U15056 ( .A(x[5262]), .B(y[5262]), .Z(n24334) );
  NANDN U15057 ( .A(y[5260]), .B(x[5260]), .Z(n9573) );
  NANDN U15058 ( .A(y[5261]), .B(x[5261]), .Z(n24333) );
  NAND U15059 ( .A(n9573), .B(n24333), .Z(n57637) );
  XNOR U15060 ( .A(x[5260]), .B(y[5260]), .Z(n43507) );
  ANDN U15061 ( .B(y[5259]), .A(x[5259]), .Z(n24335) );
  ANDN U15062 ( .B(y[5257]), .A(x[5257]), .Z(n24339) );
  NANDN U15063 ( .A(x[5258]), .B(y[5258]), .Z(n24336) );
  NANDN U15064 ( .A(n24339), .B(n24336), .Z(n57633) );
  NANDN U15065 ( .A(y[5256]), .B(x[5256]), .Z(n9574) );
  NANDN U15066 ( .A(y[5257]), .B(x[5257]), .Z(n24338) );
  AND U15067 ( .A(n9574), .B(n24338), .Z(n57632) );
  ANDN U15068 ( .B(y[5255]), .A(x[5255]), .Z(n43493) );
  XNOR U15069 ( .A(x[5256]), .B(y[5256]), .Z(n43497) );
  NANDN U15070 ( .A(y[5254]), .B(x[5254]), .Z(n9575) );
  NANDN U15071 ( .A(y[5255]), .B(x[5255]), .Z(n43496) );
  NAND U15072 ( .A(n9575), .B(n43496), .Z(n57628) );
  XNOR U15073 ( .A(x[5254]), .B(y[5254]), .Z(n24341) );
  ANDN U15074 ( .B(y[5253]), .A(x[5253]), .Z(n24342) );
  NANDN U15075 ( .A(y[5250]), .B(x[5250]), .Z(n24346) );
  NANDN U15076 ( .A(y[5251]), .B(x[5251]), .Z(n24343) );
  AND U15077 ( .A(n24346), .B(n24343), .Z(n57623) );
  NANDN U15078 ( .A(x[5249]), .B(y[5249]), .Z(n43481) );
  NANDN U15079 ( .A(x[5250]), .B(y[5250]), .Z(n24345) );
  NAND U15080 ( .A(n43481), .B(n24345), .Z(n57622) );
  NANDN U15081 ( .A(y[5248]), .B(x[5248]), .Z(n9576) );
  NANDN U15082 ( .A(y[5249]), .B(x[5249]), .Z(n24347) );
  AND U15083 ( .A(n9576), .B(n24347), .Z(n57621) );
  ANDN U15084 ( .B(y[5247]), .A(x[5247]), .Z(n43475) );
  XNOR U15085 ( .A(x[5248]), .B(y[5248]), .Z(n24349) );
  NANDN U15086 ( .A(y[5246]), .B(x[5246]), .Z(n9577) );
  NANDN U15087 ( .A(y[5247]), .B(x[5247]), .Z(n24348) );
  NAND U15088 ( .A(n9577), .B(n24348), .Z(n57619) );
  XNOR U15089 ( .A(x[5246]), .B(y[5246]), .Z(n24351) );
  NANDN U15090 ( .A(x[5245]), .B(y[5245]), .Z(n57618) );
  NANDN U15091 ( .A(y[5244]), .B(x[5244]), .Z(n24353) );
  NANDN U15092 ( .A(y[5245]), .B(x[5245]), .Z(n24350) );
  AND U15093 ( .A(n24353), .B(n24350), .Z(n57616) );
  NANDN U15094 ( .A(x[5243]), .B(y[5243]), .Z(n24355) );
  NANDN U15095 ( .A(x[5244]), .B(y[5244]), .Z(n24352) );
  AND U15096 ( .A(n24355), .B(n24352), .Z(n57615) );
  XNOR U15097 ( .A(x[5242]), .B(y[5242]), .Z(n24357) );
  NANDN U15098 ( .A(y[5240]), .B(x[5240]), .Z(n9578) );
  NANDN U15099 ( .A(y[5241]), .B(x[5241]), .Z(n24356) );
  NAND U15100 ( .A(n9578), .B(n24356), .Z(n57610) );
  XNOR U15101 ( .A(x[5240]), .B(y[5240]), .Z(n43460) );
  NANDN U15102 ( .A(y[5238]), .B(x[5238]), .Z(n9579) );
  NANDN U15103 ( .A(y[5239]), .B(x[5239]), .Z(n43459) );
  NAND U15104 ( .A(n9579), .B(n43459), .Z(n57607) );
  XNOR U15105 ( .A(x[5238]), .B(y[5238]), .Z(n24359) );
  ANDN U15106 ( .B(y[5237]), .A(x[5237]), .Z(n57606) );
  NANDN U15107 ( .A(y[5236]), .B(x[5236]), .Z(n9580) );
  NANDN U15108 ( .A(y[5237]), .B(x[5237]), .Z(n24358) );
  AND U15109 ( .A(n9580), .B(n24358), .Z(n57604) );
  NANDN U15110 ( .A(x[5235]), .B(y[5235]), .Z(n57603) );
  XNOR U15111 ( .A(x[5236]), .B(y[5236]), .Z(n43450) );
  AND U15112 ( .A(n57603), .B(n43450), .Z(n17363) );
  NANDN U15113 ( .A(x[5234]), .B(y[5234]), .Z(n24360) );
  ANDN U15114 ( .B(y[5233]), .A(x[5233]), .Z(n24363) );
  ANDN U15115 ( .B(n24360), .A(n24363), .Z(n57600) );
  NANDN U15116 ( .A(y[5232]), .B(x[5232]), .Z(n9581) );
  NANDN U15117 ( .A(y[5233]), .B(x[5233]), .Z(n24362) );
  AND U15118 ( .A(n9581), .B(n24362), .Z(n57599) );
  XNOR U15119 ( .A(x[5232]), .B(y[5232]), .Z(n43440) );
  NANDN U15120 ( .A(y[5230]), .B(x[5230]), .Z(n9582) );
  NANDN U15121 ( .A(y[5231]), .B(x[5231]), .Z(n43439) );
  AND U15122 ( .A(n9582), .B(n43439), .Z(n57596) );
  NANDN U15123 ( .A(x[5229]), .B(y[5229]), .Z(n51441) );
  XNOR U15124 ( .A(x[5230]), .B(y[5230]), .Z(n24365) );
  NAND U15125 ( .A(n51441), .B(n24365), .Z(n17355) );
  NANDN U15126 ( .A(y[5228]), .B(x[5228]), .Z(n24367) );
  NANDN U15127 ( .A(y[5229]), .B(x[5229]), .Z(n24364) );
  AND U15128 ( .A(n24367), .B(n24364), .Z(n57593) );
  NANDN U15129 ( .A(x[5227]), .B(y[5227]), .Z(n24369) );
  NANDN U15130 ( .A(x[5228]), .B(y[5228]), .Z(n24366) );
  NAND U15131 ( .A(n24369), .B(n24366), .Z(n57592) );
  NANDN U15132 ( .A(y[5226]), .B(x[5226]), .Z(n9583) );
  NANDN U15133 ( .A(y[5227]), .B(x[5227]), .Z(n24368) );
  AND U15134 ( .A(n9583), .B(n24368), .Z(n51443) );
  NANDN U15135 ( .A(y[5224]), .B(x[5224]), .Z(n9584) );
  NANDN U15136 ( .A(y[5225]), .B(x[5225]), .Z(n24370) );
  AND U15137 ( .A(n9584), .B(n24370), .Z(n57589) );
  NANDN U15138 ( .A(y[5222]), .B(x[5222]), .Z(n9585) );
  NANDN U15139 ( .A(y[5223]), .B(x[5223]), .Z(n43421) );
  AND U15140 ( .A(n9585), .B(n43421), .Z(n57588) );
  ANDN U15141 ( .B(y[5221]), .A(x[5221]), .Z(n24374) );
  XNOR U15142 ( .A(y[5222]), .B(x[5222]), .Z(n24373) );
  NANDN U15143 ( .A(n24374), .B(n24373), .Z(n57587) );
  NANDN U15144 ( .A(y[5220]), .B(x[5220]), .Z(n9586) );
  NANDN U15145 ( .A(y[5221]), .B(x[5221]), .Z(n24372) );
  AND U15146 ( .A(n9586), .B(n24372), .Z(n51446) );
  XNOR U15147 ( .A(x[5220]), .B(y[5220]), .Z(n43411) );
  NANDN U15148 ( .A(y[5218]), .B(x[5218]), .Z(n9587) );
  NANDN U15149 ( .A(y[5219]), .B(x[5219]), .Z(n43410) );
  NAND U15150 ( .A(n9587), .B(n43410), .Z(n57582) );
  XNOR U15151 ( .A(y[5218]), .B(x[5218]), .Z(n24376) );
  NANDN U15152 ( .A(x[5217]), .B(y[5217]), .Z(n24377) );
  AND U15153 ( .A(n24376), .B(n24377), .Z(n51447) );
  NANDN U15154 ( .A(x[5215]), .B(y[5215]), .Z(n57581) );
  XNOR U15155 ( .A(x[5216]), .B(y[5216]), .Z(n24379) );
  AND U15156 ( .A(n57581), .B(n24379), .Z(n17336) );
  NANDN U15157 ( .A(y[5214]), .B(x[5214]), .Z(n9588) );
  NANDN U15158 ( .A(y[5215]), .B(x[5215]), .Z(n24378) );
  NAND U15159 ( .A(n9588), .B(n24378), .Z(n57580) );
  XNOR U15160 ( .A(x[5214]), .B(y[5214]), .Z(n24381) );
  XNOR U15161 ( .A(x[5212]), .B(y[5212]), .Z(n43392) );
  NANDN U15162 ( .A(y[5210]), .B(x[5210]), .Z(n9589) );
  NANDN U15163 ( .A(y[5211]), .B(x[5211]), .Z(n43391) );
  NAND U15164 ( .A(n9589), .B(n43391), .Z(n57576) );
  XNOR U15165 ( .A(x[5210]), .B(y[5210]), .Z(n24383) );
  ANDN U15166 ( .B(y[5209]), .A(x[5209]), .Z(n57572) );
  XNOR U15167 ( .A(x[5208]), .B(y[5208]), .Z(n43382) );
  NANDN U15168 ( .A(x[5207]), .B(y[5207]), .Z(n57570) );
  AND U15169 ( .A(n43382), .B(n57570), .Z(n17322) );
  NANDN U15170 ( .A(y[5204]), .B(x[5204]), .Z(n24389) );
  NANDN U15171 ( .A(y[5205]), .B(x[5205]), .Z(n24386) );
  NAND U15172 ( .A(n24389), .B(n24386), .Z(n51454) );
  NANDN U15173 ( .A(x[5203]), .B(y[5203]), .Z(n24391) );
  NANDN U15174 ( .A(x[5204]), .B(y[5204]), .Z(n24388) );
  AND U15175 ( .A(n24391), .B(n24388), .Z(n57568) );
  XNOR U15176 ( .A(x[5202]), .B(y[5202]), .Z(n24393) );
  ANDN U15177 ( .B(y[5201]), .A(x[5201]), .Z(n51456) );
  NANDN U15178 ( .A(y[5200]), .B(x[5200]), .Z(n9590) );
  NANDN U15179 ( .A(y[5201]), .B(x[5201]), .Z(n24392) );
  AND U15180 ( .A(n9590), .B(n24392), .Z(n57566) );
  XNOR U15181 ( .A(x[5200]), .B(y[5200]), .Z(n43364) );
  XNOR U15182 ( .A(x[5198]), .B(y[5198]), .Z(n24395) );
  NANDN U15183 ( .A(y[5196]), .B(x[5196]), .Z(n9591) );
  NANDN U15184 ( .A(y[5197]), .B(x[5197]), .Z(n24394) );
  NAND U15185 ( .A(n9591), .B(n24394), .Z(n57560) );
  XNOR U15186 ( .A(x[5196]), .B(y[5196]), .Z(n43353) );
  ANDN U15187 ( .B(y[5195]), .A(x[5195]), .Z(n43349) );
  XNOR U15188 ( .A(x[5194]), .B(y[5194]), .Z(n24397) );
  NANDN U15189 ( .A(x[5193]), .B(y[5193]), .Z(n57557) );
  AND U15190 ( .A(n24397), .B(n57557), .Z(n17300) );
  XNOR U15191 ( .A(x[5192]), .B(y[5192]), .Z(n24399) );
  NANDN U15192 ( .A(x[5190]), .B(y[5190]), .Z(n24400) );
  ANDN U15193 ( .B(y[5189]), .A(x[5189]), .Z(n24403) );
  ANDN U15194 ( .B(n24400), .A(n24403), .Z(n57552) );
  NANDN U15195 ( .A(y[5188]), .B(x[5188]), .Z(n9592) );
  NANDN U15196 ( .A(y[5189]), .B(x[5189]), .Z(n24402) );
  NAND U15197 ( .A(n9592), .B(n24402), .Z(n51462) );
  XNOR U15198 ( .A(x[5188]), .B(y[5188]), .Z(n43334) );
  ANDN U15199 ( .B(y[5187]), .A(x[5187]), .Z(n24404) );
  NANDN U15200 ( .A(x[5185]), .B(y[5185]), .Z(n24408) );
  NANDN U15201 ( .A(x[5186]), .B(y[5186]), .Z(n24405) );
  NAND U15202 ( .A(n24408), .B(n24405), .Z(n57549) );
  NANDN U15203 ( .A(y[5184]), .B(x[5184]), .Z(n9593) );
  NANDN U15204 ( .A(y[5185]), .B(x[5185]), .Z(n24407) );
  AND U15205 ( .A(n9593), .B(n24407), .Z(n57548) );
  ANDN U15206 ( .B(y[5183]), .A(x[5183]), .Z(n24409) );
  ANDN U15207 ( .B(x[5183]), .A(y[5183]), .Z(n43324) );
  NANDN U15208 ( .A(y[5182]), .B(x[5182]), .Z(n9594) );
  NANDN U15209 ( .A(n43324), .B(n9594), .Z(n57545) );
  XNOR U15210 ( .A(x[5182]), .B(y[5182]), .Z(n24411) );
  ANDN U15211 ( .B(y[5181]), .A(x[5181]), .Z(n57543) );
  NANDN U15212 ( .A(y[5180]), .B(x[5180]), .Z(n9595) );
  NANDN U15213 ( .A(y[5181]), .B(x[5181]), .Z(n24410) );
  AND U15214 ( .A(n9595), .B(n24410), .Z(n51465) );
  XNOR U15215 ( .A(x[5180]), .B(y[5180]), .Z(n43314) );
  NANDN U15216 ( .A(x[5179]), .B(y[5179]), .Z(n57539) );
  AND U15217 ( .A(n43314), .B(n57539), .Z(n17280) );
  NANDN U15218 ( .A(y[5178]), .B(x[5178]), .Z(n24413) );
  NANDN U15219 ( .A(y[5179]), .B(x[5179]), .Z(n43313) );
  AND U15220 ( .A(n24413), .B(n43313), .Z(n57538) );
  ANDN U15221 ( .B(y[5177]), .A(x[5177]), .Z(n24415) );
  NANDN U15222 ( .A(x[5178]), .B(y[5178]), .Z(n24412) );
  NANDN U15223 ( .A(n24415), .B(n24412), .Z(n57537) );
  NANDN U15224 ( .A(y[5176]), .B(x[5176]), .Z(n9596) );
  NANDN U15225 ( .A(y[5177]), .B(x[5177]), .Z(n24414) );
  AND U15226 ( .A(n9596), .B(n24414), .Z(n57536) );
  ANDN U15227 ( .B(y[5175]), .A(x[5175]), .Z(n43300) );
  XNOR U15228 ( .A(x[5176]), .B(y[5176]), .Z(n43304) );
  NANDN U15229 ( .A(y[5174]), .B(x[5174]), .Z(n9597) );
  NANDN U15230 ( .A(y[5175]), .B(x[5175]), .Z(n43303) );
  NAND U15231 ( .A(n9597), .B(n43303), .Z(n57533) );
  XNOR U15232 ( .A(x[5174]), .B(y[5174]), .Z(n24417) );
  ANDN U15233 ( .B(y[5173]), .A(x[5173]), .Z(n57532) );
  NANDN U15234 ( .A(y[5172]), .B(x[5172]), .Z(n9598) );
  NANDN U15235 ( .A(y[5173]), .B(x[5173]), .Z(n24416) );
  AND U15236 ( .A(n9598), .B(n24416), .Z(n57530) );
  XNOR U15237 ( .A(x[5172]), .B(y[5172]), .Z(n43293) );
  NANDN U15238 ( .A(x[5171]), .B(y[5171]), .Z(n51466) );
  AND U15239 ( .A(n43293), .B(n51466), .Z(n17269) );
  XNOR U15240 ( .A(x[5170]), .B(y[5170]), .Z(n24419) );
  NANDN U15241 ( .A(x[5167]), .B(y[5167]), .Z(n43281) );
  NANDN U15242 ( .A(x[5168]), .B(y[5168]), .Z(n24420) );
  AND U15243 ( .A(n43281), .B(n24420), .Z(n57525) );
  NANDN U15244 ( .A(y[5166]), .B(x[5166]), .Z(n9599) );
  NANDN U15245 ( .A(y[5167]), .B(x[5167]), .Z(n24422) );
  NAND U15246 ( .A(n9599), .B(n24422), .Z(n57524) );
  XNOR U15247 ( .A(x[5166]), .B(y[5166]), .Z(n24424) );
  ANDN U15248 ( .B(y[5165]), .A(x[5165]), .Z(n24425) );
  NANDN U15249 ( .A(x[5163]), .B(y[5163]), .Z(n57520) );
  XNOR U15250 ( .A(x[5164]), .B(y[5164]), .Z(n24427) );
  AND U15251 ( .A(n57520), .B(n24427), .Z(n17256) );
  NANDN U15252 ( .A(y[5162]), .B(x[5162]), .Z(n24429) );
  NANDN U15253 ( .A(y[5163]), .B(x[5163]), .Z(n24426) );
  NAND U15254 ( .A(n24429), .B(n24426), .Z(n57519) );
  NANDN U15255 ( .A(x[5161]), .B(y[5161]), .Z(n43268) );
  NANDN U15256 ( .A(x[5162]), .B(y[5162]), .Z(n24428) );
  AND U15257 ( .A(n43268), .B(n24428), .Z(n57518) );
  NANDN U15258 ( .A(y[5160]), .B(x[5160]), .Z(n24431) );
  NANDN U15259 ( .A(y[5161]), .B(x[5161]), .Z(n24430) );
  NAND U15260 ( .A(n24431), .B(n24430), .Z(n57517) );
  NANDN U15261 ( .A(x[5159]), .B(y[5159]), .Z(n43262) );
  NANDN U15262 ( .A(x[5160]), .B(y[5160]), .Z(n43269) );
  AND U15263 ( .A(n43262), .B(n43269), .Z(n57516) );
  NANDN U15264 ( .A(y[5158]), .B(x[5158]), .Z(n9600) );
  NANDN U15265 ( .A(y[5159]), .B(x[5159]), .Z(n24432) );
  NAND U15266 ( .A(n9600), .B(n24432), .Z(n57515) );
  XNOR U15267 ( .A(x[5158]), .B(y[5158]), .Z(n24434) );
  NANDN U15268 ( .A(x[5157]), .B(y[5157]), .Z(n57513) );
  AND U15269 ( .A(n24434), .B(n57513), .Z(n17249) );
  XNOR U15270 ( .A(x[5156]), .B(y[5156]), .Z(n24436) );
  NANDN U15271 ( .A(y[5152]), .B(x[5152]), .Z(n9601) );
  NANDN U15272 ( .A(y[5153]), .B(x[5153]), .Z(n24439) );
  NAND U15273 ( .A(n9601), .B(n24439), .Z(n51471) );
  XNOR U15274 ( .A(y[5152]), .B(x[5152]), .Z(n43247) );
  NANDN U15275 ( .A(x[5151]), .B(y[5151]), .Z(n57505) );
  NANDN U15276 ( .A(y[5150]), .B(x[5150]), .Z(n24441) );
  ANDN U15277 ( .B(x[5151]), .A(y[5151]), .Z(n43249) );
  ANDN U15278 ( .B(n24441), .A(n43249), .Z(n57504) );
  ANDN U15279 ( .B(y[5149]), .A(x[5149]), .Z(n24443) );
  NANDN U15280 ( .A(x[5150]), .B(y[5150]), .Z(n43243) );
  NANDN U15281 ( .A(n24443), .B(n43243), .Z(n51472) );
  NANDN U15282 ( .A(y[5148]), .B(x[5148]), .Z(n9602) );
  NANDN U15283 ( .A(y[5149]), .B(x[5149]), .Z(n24442) );
  AND U15284 ( .A(n9602), .B(n24442), .Z(n57503) );
  ANDN U15285 ( .B(y[5147]), .A(x[5147]), .Z(n43232) );
  XNOR U15286 ( .A(x[5148]), .B(y[5148]), .Z(n43236) );
  NANDN U15287 ( .A(y[5146]), .B(x[5146]), .Z(n9603) );
  NANDN U15288 ( .A(y[5147]), .B(x[5147]), .Z(n43235) );
  NAND U15289 ( .A(n9603), .B(n43235), .Z(n57502) );
  NANDN U15290 ( .A(x[5145]), .B(y[5145]), .Z(n57500) );
  NANDN U15291 ( .A(x[5143]), .B(y[5143]), .Z(n24449) );
  NANDN U15292 ( .A(x[5144]), .B(y[5144]), .Z(n24446) );
  AND U15293 ( .A(n24449), .B(n24446), .Z(n57498) );
  NANDN U15294 ( .A(y[5140]), .B(x[5140]), .Z(n24455) );
  NANDN U15295 ( .A(y[5141]), .B(x[5141]), .Z(n24451) );
  NAND U15296 ( .A(n24455), .B(n24451), .Z(n51476) );
  NANDN U15297 ( .A(x[5139]), .B(y[5139]), .Z(n24457) );
  NANDN U15298 ( .A(x[5140]), .B(y[5140]), .Z(n24454) );
  AND U15299 ( .A(n24457), .B(n24454), .Z(n57494) );
  NANDN U15300 ( .A(y[5136]), .B(x[5136]), .Z(n9604) );
  NANDN U15301 ( .A(y[5137]), .B(x[5137]), .Z(n24458) );
  AND U15302 ( .A(n9604), .B(n24458), .Z(n57490) );
  XNOR U15303 ( .A(x[5136]), .B(y[5136]), .Z(n43209) );
  XNOR U15304 ( .A(x[5134]), .B(y[5134]), .Z(n24462) );
  NANDN U15305 ( .A(y[5132]), .B(x[5132]), .Z(n9605) );
  NANDN U15306 ( .A(y[5133]), .B(x[5133]), .Z(n24461) );
  NAND U15307 ( .A(n9605), .B(n24461), .Z(n57486) );
  XNOR U15308 ( .A(x[5132]), .B(y[5132]), .Z(n43198) );
  ANDN U15309 ( .B(y[5131]), .A(x[5131]), .Z(n43194) );
  XNOR U15310 ( .A(x[5130]), .B(y[5130]), .Z(n24464) );
  ANDN U15311 ( .B(y[5129]), .A(x[5129]), .Z(n57481) );
  ANDN U15312 ( .B(n24464), .A(n57481), .Z(n17206) );
  XNOR U15313 ( .A(x[5128]), .B(y[5128]), .Z(n43187) );
  NANDN U15314 ( .A(y[5126]), .B(x[5126]), .Z(n9606) );
  NANDN U15315 ( .A(y[5127]), .B(x[5127]), .Z(n43186) );
  AND U15316 ( .A(n9606), .B(n43186), .Z(n57478) );
  NANDN U15317 ( .A(y[5124]), .B(x[5124]), .Z(n9607) );
  NANDN U15318 ( .A(y[5125]), .B(x[5125]), .Z(n24465) );
  AND U15319 ( .A(n9607), .B(n24465), .Z(n57476) );
  XNOR U15320 ( .A(y[5124]), .B(x[5124]), .Z(n24470) );
  NANDN U15321 ( .A(x[5123]), .B(y[5123]), .Z(n24471) );
  NAND U15322 ( .A(n24470), .B(n24471), .Z(n57475) );
  NANDN U15323 ( .A(y[5122]), .B(x[5122]), .Z(n9608) );
  NANDN U15324 ( .A(y[5123]), .B(x[5123]), .Z(n24469) );
  AND U15325 ( .A(n9608), .B(n24469), .Z(n57474) );
  XNOR U15326 ( .A(y[5122]), .B(x[5122]), .Z(n24474) );
  NANDN U15327 ( .A(x[5121]), .B(y[5121]), .Z(n24475) );
  NAND U15328 ( .A(n24474), .B(n24475), .Z(n57473) );
  NANDN U15329 ( .A(y[5120]), .B(x[5120]), .Z(n24477) );
  NANDN U15330 ( .A(y[5121]), .B(x[5121]), .Z(n24473) );
  AND U15331 ( .A(n24477), .B(n24473), .Z(n57472) );
  NANDN U15332 ( .A(y[5118]), .B(x[5118]), .Z(n9609) );
  NANDN U15333 ( .A(y[5119]), .B(x[5119]), .Z(n24478) );
  AND U15334 ( .A(n9609), .B(n24478), .Z(n57470) );
  NANDN U15335 ( .A(x[5117]), .B(y[5117]), .Z(n57469) );
  XNOR U15336 ( .A(x[5118]), .B(y[5118]), .Z(n24481) );
  AND U15337 ( .A(n57469), .B(n24481), .Z(n17191) );
  XNOR U15338 ( .A(x[5116]), .B(y[5116]), .Z(n24483) );
  NANDN U15339 ( .A(y[5114]), .B(x[5114]), .Z(n9610) );
  NANDN U15340 ( .A(y[5115]), .B(x[5115]), .Z(n24482) );
  NAND U15341 ( .A(n9610), .B(n24482), .Z(n57464) );
  ANDN U15342 ( .B(y[5113]), .A(x[5113]), .Z(n57462) );
  XNOR U15343 ( .A(x[5114]), .B(y[5114]), .Z(n24485) );
  NANDN U15344 ( .A(y[5112]), .B(x[5112]), .Z(n9611) );
  NANDN U15345 ( .A(y[5113]), .B(x[5113]), .Z(n24484) );
  NAND U15346 ( .A(n9611), .B(n24484), .Z(n57461) );
  XNOR U15347 ( .A(x[5112]), .B(y[5112]), .Z(n43152) );
  ANDN U15348 ( .B(y[5111]), .A(x[5111]), .Z(n43148) );
  NANDN U15349 ( .A(y[5110]), .B(x[5110]), .Z(n9612) );
  NANDN U15350 ( .A(y[5111]), .B(x[5111]), .Z(n43151) );
  AND U15351 ( .A(n9612), .B(n43151), .Z(n57458) );
  XNOR U15352 ( .A(x[5110]), .B(y[5110]), .Z(n24487) );
  NANDN U15353 ( .A(x[5109]), .B(y[5109]), .Z(n51484) );
  AND U15354 ( .A(n24487), .B(n51484), .Z(n17178) );
  XNOR U15355 ( .A(x[5108]), .B(y[5108]), .Z(n24489) );
  XNOR U15356 ( .A(x[5106]), .B(y[5106]), .Z(n24491) );
  NANDN U15357 ( .A(y[5104]), .B(x[5104]), .Z(n9613) );
  NANDN U15358 ( .A(y[5105]), .B(x[5105]), .Z(n24490) );
  NAND U15359 ( .A(n9613), .B(n24490), .Z(n57452) );
  XNOR U15360 ( .A(y[5104]), .B(x[5104]), .Z(n24494) );
  NANDN U15361 ( .A(x[5103]), .B(y[5103]), .Z(n24495) );
  AND U15362 ( .A(n24494), .B(n24495), .Z(n57451) );
  NANDN U15363 ( .A(y[5102]), .B(x[5102]), .Z(n24497) );
  NANDN U15364 ( .A(y[5103]), .B(x[5103]), .Z(n24493) );
  NAND U15365 ( .A(n24497), .B(n24493), .Z(n57450) );
  NANDN U15366 ( .A(x[5101]), .B(y[5101]), .Z(n43127) );
  XNOR U15367 ( .A(x[5102]), .B(y[5102]), .Z(n9614) );
  AND U15368 ( .A(n43127), .B(n9614), .Z(n57449) );
  NANDN U15369 ( .A(y[5100]), .B(x[5100]), .Z(n24499) );
  NANDN U15370 ( .A(y[5101]), .B(x[5101]), .Z(n24498) );
  NAND U15371 ( .A(n24499), .B(n24498), .Z(n57448) );
  NANDN U15372 ( .A(x[5099]), .B(y[5099]), .Z(n43120) );
  NANDN U15373 ( .A(x[5100]), .B(y[5100]), .Z(n43128) );
  AND U15374 ( .A(n43120), .B(n43128), .Z(n57447) );
  NANDN U15375 ( .A(y[5098]), .B(x[5098]), .Z(n24501) );
  NANDN U15376 ( .A(y[5099]), .B(x[5099]), .Z(n24500) );
  NAND U15377 ( .A(n24501), .B(n24500), .Z(n57446) );
  NANDN U15378 ( .A(x[5098]), .B(y[5098]), .Z(n43121) );
  ANDN U15379 ( .B(y[5097]), .A(x[5097]), .Z(n24503) );
  ANDN U15380 ( .B(n43121), .A(n24503), .Z(n57445) );
  NANDN U15381 ( .A(y[5096]), .B(x[5096]), .Z(n9615) );
  NANDN U15382 ( .A(y[5097]), .B(x[5097]), .Z(n24502) );
  NAND U15383 ( .A(n9615), .B(n24502), .Z(n57444) );
  XNOR U15384 ( .A(x[5096]), .B(y[5096]), .Z(n43113) );
  ANDN U15385 ( .B(y[5095]), .A(x[5095]), .Z(n43109) );
  XNOR U15386 ( .A(x[5094]), .B(y[5094]), .Z(n24505) );
  NANDN U15387 ( .A(y[5092]), .B(x[5092]), .Z(n24507) );
  NANDN U15388 ( .A(y[5093]), .B(x[5093]), .Z(n24504) );
  NAND U15389 ( .A(n24507), .B(n24504), .Z(n57440) );
  NANDN U15390 ( .A(x[5091]), .B(y[5091]), .Z(n24509) );
  NANDN U15391 ( .A(x[5092]), .B(y[5092]), .Z(n24506) );
  AND U15392 ( .A(n24509), .B(n24506), .Z(n57439) );
  NANDN U15393 ( .A(y[5090]), .B(x[5090]), .Z(n24511) );
  NANDN U15394 ( .A(y[5091]), .B(x[5091]), .Z(n24508) );
  NAND U15395 ( .A(n24511), .B(n24508), .Z(n57438) );
  NANDN U15396 ( .A(x[5089]), .B(y[5089]), .Z(n24513) );
  NANDN U15397 ( .A(x[5090]), .B(y[5090]), .Z(n24510) );
  AND U15398 ( .A(n24513), .B(n24510), .Z(n57437) );
  NANDN U15399 ( .A(y[5088]), .B(x[5088]), .Z(n9616) );
  NANDN U15400 ( .A(y[5089]), .B(x[5089]), .Z(n24512) );
  NAND U15401 ( .A(n9616), .B(n24512), .Z(n57434) );
  XNOR U15402 ( .A(x[5088]), .B(y[5088]), .Z(n24515) );
  NANDN U15403 ( .A(y[5086]), .B(x[5086]), .Z(n9617) );
  NANDN U15404 ( .A(y[5087]), .B(x[5087]), .Z(n24514) );
  NAND U15405 ( .A(n9617), .B(n24514), .Z(n57431) );
  XNOR U15406 ( .A(x[5086]), .B(y[5086]), .Z(n24517) );
  ANDN U15407 ( .B(y[5085]), .A(x[5085]), .Z(n57429) );
  NANDN U15408 ( .A(y[5084]), .B(x[5084]), .Z(n9618) );
  NANDN U15409 ( .A(y[5085]), .B(x[5085]), .Z(n24516) );
  AND U15410 ( .A(n9618), .B(n24516), .Z(n51490) );
  XNOR U15411 ( .A(x[5084]), .B(y[5084]), .Z(n43086) );
  NANDN U15412 ( .A(x[5083]), .B(y[5083]), .Z(n57427) );
  AND U15413 ( .A(n43086), .B(n57427), .Z(n17142) );
  NANDN U15414 ( .A(y[5082]), .B(x[5082]), .Z(n9619) );
  NANDN U15415 ( .A(y[5083]), .B(x[5083]), .Z(n43085) );
  AND U15416 ( .A(n9619), .B(n43085), .Z(n57426) );
  XNOR U15417 ( .A(x[5082]), .B(y[5082]), .Z(n24519) );
  ANDN U15418 ( .B(y[5081]), .A(x[5081]), .Z(n51492) );
  ANDN U15419 ( .B(n24519), .A(n51492), .Z(n17139) );
  XNOR U15420 ( .A(x[5080]), .B(y[5080]), .Z(n43076) );
  NANDN U15421 ( .A(y[5078]), .B(x[5078]), .Z(n24521) );
  NANDN U15422 ( .A(y[5079]), .B(x[5079]), .Z(n43075) );
  NAND U15423 ( .A(n24521), .B(n43075), .Z(n57422) );
  NANDN U15424 ( .A(x[5078]), .B(y[5078]), .Z(n24520) );
  ANDN U15425 ( .B(y[5077]), .A(x[5077]), .Z(n24523) );
  ANDN U15426 ( .B(n24520), .A(n24523), .Z(n57420) );
  NANDN U15427 ( .A(y[5076]), .B(x[5076]), .Z(n9620) );
  NANDN U15428 ( .A(y[5077]), .B(x[5077]), .Z(n24522) );
  NAND U15429 ( .A(n9620), .B(n24522), .Z(n57419) );
  NANDN U15430 ( .A(x[5075]), .B(y[5075]), .Z(n51494) );
  XNOR U15431 ( .A(x[5076]), .B(y[5076]), .Z(n43066) );
  AND U15432 ( .A(n51494), .B(n43066), .Z(n17130) );
  NANDN U15433 ( .A(y[5074]), .B(x[5074]), .Z(n24525) );
  NANDN U15434 ( .A(y[5075]), .B(x[5075]), .Z(n43065) );
  NAND U15435 ( .A(n24525), .B(n43065), .Z(n57418) );
  NANDN U15436 ( .A(x[5073]), .B(y[5073]), .Z(n24527) );
  NANDN U15437 ( .A(x[5074]), .B(y[5074]), .Z(n24524) );
  AND U15438 ( .A(n24527), .B(n24524), .Z(n57417) );
  NANDN U15439 ( .A(y[5072]), .B(x[5072]), .Z(n9621) );
  NANDN U15440 ( .A(y[5073]), .B(x[5073]), .Z(n24526) );
  NAND U15441 ( .A(n9621), .B(n24526), .Z(n57416) );
  XNOR U15442 ( .A(x[5072]), .B(y[5072]), .Z(n24529) );
  NANDN U15443 ( .A(x[5071]), .B(y[5071]), .Z(n57415) );
  AND U15444 ( .A(n24529), .B(n57415), .Z(n17125) );
  NANDN U15445 ( .A(x[5070]), .B(y[5070]), .Z(n24530) );
  ANDN U15446 ( .B(y[5069]), .A(x[5069]), .Z(n24533) );
  ANDN U15447 ( .B(n24530), .A(n24533), .Z(n57412) );
  XNOR U15448 ( .A(x[5068]), .B(y[5068]), .Z(n43048) );
  NANDN U15449 ( .A(y[5066]), .B(x[5066]), .Z(n9622) );
  NANDN U15450 ( .A(y[5067]), .B(x[5067]), .Z(n43047) );
  NAND U15451 ( .A(n9622), .B(n43047), .Z(n57407) );
  XNOR U15452 ( .A(x[5066]), .B(y[5066]), .Z(n24535) );
  NANDN U15453 ( .A(y[5064]), .B(x[5064]), .Z(n9623) );
  NANDN U15454 ( .A(y[5065]), .B(x[5065]), .Z(n24534) );
  NAND U15455 ( .A(n9623), .B(n24534), .Z(n57404) );
  XNOR U15456 ( .A(x[5064]), .B(y[5064]), .Z(n43038) );
  NANDN U15457 ( .A(x[5063]), .B(y[5063]), .Z(n57403) );
  NANDN U15458 ( .A(y[5062]), .B(x[5062]), .Z(n9624) );
  NANDN U15459 ( .A(y[5063]), .B(x[5063]), .Z(n43037) );
  AND U15460 ( .A(n9624), .B(n43037), .Z(n57401) );
  XNOR U15461 ( .A(x[5062]), .B(y[5062]), .Z(n24537) );
  ANDN U15462 ( .B(y[5061]), .A(x[5061]), .Z(n51496) );
  ANDN U15463 ( .B(n24537), .A(n51496), .Z(n17110) );
  XNOR U15464 ( .A(x[5060]), .B(y[5060]), .Z(n43028) );
  NANDN U15465 ( .A(y[5058]), .B(x[5058]), .Z(n24539) );
  NANDN U15466 ( .A(y[5059]), .B(x[5059]), .Z(n43027) );
  NAND U15467 ( .A(n24539), .B(n43027), .Z(n57397) );
  NANDN U15468 ( .A(x[5057]), .B(y[5057]), .Z(n24541) );
  NANDN U15469 ( .A(x[5058]), .B(y[5058]), .Z(n24538) );
  AND U15470 ( .A(n24541), .B(n24538), .Z(n57396) );
  NANDN U15471 ( .A(y[5056]), .B(x[5056]), .Z(n24543) );
  NANDN U15472 ( .A(y[5057]), .B(x[5057]), .Z(n24540) );
  NAND U15473 ( .A(n24543), .B(n24540), .Z(n57395) );
  NANDN U15474 ( .A(x[5055]), .B(y[5055]), .Z(n24545) );
  NANDN U15475 ( .A(x[5056]), .B(y[5056]), .Z(n24542) );
  AND U15476 ( .A(n24545), .B(n24542), .Z(n57394) );
  XNOR U15477 ( .A(x[5054]), .B(y[5054]), .Z(n24547) );
  NANDN U15478 ( .A(y[5052]), .B(x[5052]), .Z(n9625) );
  NANDN U15479 ( .A(y[5053]), .B(x[5053]), .Z(n24546) );
  NAND U15480 ( .A(n9625), .B(n24546), .Z(n57389) );
  XNOR U15481 ( .A(x[5052]), .B(y[5052]), .Z(n43010) );
  NANDN U15482 ( .A(y[5050]), .B(x[5050]), .Z(n9626) );
  NANDN U15483 ( .A(y[5051]), .B(x[5051]), .Z(n43009) );
  NAND U15484 ( .A(n9626), .B(n43009), .Z(n57386) );
  NANDN U15485 ( .A(x[5047]), .B(y[5047]), .Z(n24553) );
  NANDN U15486 ( .A(x[5048]), .B(y[5048]), .Z(n24550) );
  AND U15487 ( .A(n24553), .B(n24550), .Z(n57384) );
  XNOR U15488 ( .A(x[5046]), .B(y[5046]), .Z(n24555) );
  NANDN U15489 ( .A(y[5044]), .B(x[5044]), .Z(n24557) );
  NANDN U15490 ( .A(y[5045]), .B(x[5045]), .Z(n24554) );
  NAND U15491 ( .A(n24557), .B(n24554), .Z(n57380) );
  NANDN U15492 ( .A(x[5043]), .B(y[5043]), .Z(n42990) );
  NANDN U15493 ( .A(x[5044]), .B(y[5044]), .Z(n24556) );
  AND U15494 ( .A(n42990), .B(n24556), .Z(n51499) );
  NANDN U15495 ( .A(x[5041]), .B(y[5041]), .Z(n57377) );
  XNOR U15496 ( .A(x[5042]), .B(y[5042]), .Z(n24560) );
  AND U15497 ( .A(n57377), .B(n24560), .Z(n17080) );
  NANDN U15498 ( .A(y[5040]), .B(x[5040]), .Z(n24562) );
  NANDN U15499 ( .A(y[5041]), .B(x[5041]), .Z(n24559) );
  NAND U15500 ( .A(n24562), .B(n24559), .Z(n57376) );
  NANDN U15501 ( .A(x[5039]), .B(y[5039]), .Z(n24564) );
  NANDN U15502 ( .A(x[5040]), .B(y[5040]), .Z(n24561) );
  AND U15503 ( .A(n24564), .B(n24561), .Z(n57375) );
  NANDN U15504 ( .A(y[5038]), .B(x[5038]), .Z(n9627) );
  NANDN U15505 ( .A(y[5039]), .B(x[5039]), .Z(n24563) );
  NAND U15506 ( .A(n9627), .B(n24563), .Z(n57374) );
  XNOR U15507 ( .A(x[5038]), .B(y[5038]), .Z(n24566) );
  NANDN U15508 ( .A(x[5037]), .B(y[5037]), .Z(n51501) );
  AND U15509 ( .A(n24566), .B(n51501), .Z(n17075) );
  NANDN U15510 ( .A(y[5036]), .B(x[5036]), .Z(n24567) );
  NANDN U15511 ( .A(y[5037]), .B(x[5037]), .Z(n24565) );
  NAND U15512 ( .A(n24567), .B(n24565), .Z(n57373) );
  NANDN U15513 ( .A(x[5035]), .B(y[5035]), .Z(n24569) );
  ANDN U15514 ( .B(y[5036]), .A(x[5036]), .Z(n42977) );
  ANDN U15515 ( .B(n24569), .A(n42977), .Z(n57372) );
  NANDN U15516 ( .A(x[5033]), .B(y[5033]), .Z(n24573) );
  NANDN U15517 ( .A(x[5034]), .B(y[5034]), .Z(n24570) );
  AND U15518 ( .A(n24573), .B(n24570), .Z(n57370) );
  NANDN U15519 ( .A(y[5032]), .B(x[5032]), .Z(n24575) );
  NANDN U15520 ( .A(y[5033]), .B(x[5033]), .Z(n24572) );
  NAND U15521 ( .A(n24575), .B(n24572), .Z(n57369) );
  NANDN U15522 ( .A(x[5031]), .B(y[5031]), .Z(n24577) );
  NANDN U15523 ( .A(x[5032]), .B(y[5032]), .Z(n24574) );
  AND U15524 ( .A(n24577), .B(n24574), .Z(n57368) );
  NANDN U15525 ( .A(y[5030]), .B(x[5030]), .Z(n9628) );
  NANDN U15526 ( .A(y[5031]), .B(x[5031]), .Z(n24576) );
  NAND U15527 ( .A(n9628), .B(n24576), .Z(n57367) );
  XNOR U15528 ( .A(x[5030]), .B(y[5030]), .Z(n24579) );
  ANDN U15529 ( .B(y[5029]), .A(x[5029]), .Z(n57365) );
  ANDN U15530 ( .B(n24579), .A(n57365), .Z(n17066) );
  NANDN U15531 ( .A(y[5028]), .B(x[5028]), .Z(n9629) );
  NANDN U15532 ( .A(y[5029]), .B(x[5029]), .Z(n24578) );
  NAND U15533 ( .A(n9629), .B(n24578), .Z(n57364) );
  XNOR U15534 ( .A(x[5028]), .B(y[5028]), .Z(n42958) );
  NANDN U15535 ( .A(y[5026]), .B(x[5026]), .Z(n9630) );
  NANDN U15536 ( .A(y[5027]), .B(x[5027]), .Z(n42957) );
  NAND U15537 ( .A(n9630), .B(n42957), .Z(n57359) );
  XNOR U15538 ( .A(y[5026]), .B(x[5026]), .Z(n24581) );
  ANDN U15539 ( .B(y[5025]), .A(x[5025]), .Z(n42951) );
  ANDN U15540 ( .B(n24581), .A(n42951), .Z(n57358) );
  XNOR U15541 ( .A(x[5024]), .B(y[5024]), .Z(n24583) );
  NANDN U15542 ( .A(x[5023]), .B(y[5023]), .Z(n57356) );
  AND U15543 ( .A(n24583), .B(n57356), .Z(n17057) );
  XNOR U15544 ( .A(x[5022]), .B(y[5022]), .Z(n24585) );
  NANDN U15545 ( .A(y[5018]), .B(x[5018]), .Z(n9631) );
  NANDN U15546 ( .A(y[5019]), .B(x[5019]), .Z(n24588) );
  NAND U15547 ( .A(n9631), .B(n24588), .Z(n51505) );
  XNOR U15548 ( .A(x[5018]), .B(y[5018]), .Z(n24590) );
  ANDN U15549 ( .B(y[5017]), .A(x[5017]), .Z(n57349) );
  NANDN U15550 ( .A(x[5015]), .B(y[5015]), .Z(n57346) );
  XNOR U15551 ( .A(x[5016]), .B(y[5016]), .Z(n42929) );
  AND U15552 ( .A(n57346), .B(n42929), .Z(n17044) );
  NANDN U15553 ( .A(x[5013]), .B(y[5013]), .Z(n24594) );
  NANDN U15554 ( .A(x[5014]), .B(y[5014]), .Z(n24591) );
  AND U15555 ( .A(n24594), .B(n24591), .Z(n57343) );
  NANDN U15556 ( .A(y[5012]), .B(x[5012]), .Z(n9632) );
  NANDN U15557 ( .A(y[5013]), .B(x[5013]), .Z(n24593) );
  NAND U15558 ( .A(n9632), .B(n24593), .Z(n57342) );
  XNOR U15559 ( .A(x[5012]), .B(y[5012]), .Z(n24596) );
  ANDN U15560 ( .B(y[5011]), .A(x[5011]), .Z(n24597) );
  NANDN U15561 ( .A(x[5007]), .B(y[5007]), .Z(n57336) );
  XNOR U15562 ( .A(x[5008]), .B(y[5008]), .Z(n42911) );
  AND U15563 ( .A(n57336), .B(n42911), .Z(n17031) );
  NANDN U15564 ( .A(x[5006]), .B(y[5006]), .Z(n24600) );
  ANDN U15565 ( .B(y[5005]), .A(x[5005]), .Z(n24603) );
  ANDN U15566 ( .B(n24600), .A(n24603), .Z(n57333) );
  NANDN U15567 ( .A(y[5004]), .B(x[5004]), .Z(n9633) );
  NANDN U15568 ( .A(y[5005]), .B(x[5005]), .Z(n24602) );
  NAND U15569 ( .A(n9633), .B(n24602), .Z(n51508) );
  XNOR U15570 ( .A(x[5004]), .B(y[5004]), .Z(n42901) );
  ANDN U15571 ( .B(y[5003]), .A(x[5003]), .Z(n42897) );
  NANDN U15572 ( .A(x[5001]), .B(y[5001]), .Z(n57329) );
  XNOR U15573 ( .A(x[5002]), .B(y[5002]), .Z(n24605) );
  AND U15574 ( .A(n57329), .B(n24605), .Z(n17022) );
  NANDN U15575 ( .A(x[4999]), .B(y[4999]), .Z(n42889) );
  NANDN U15576 ( .A(x[5000]), .B(y[5000]), .Z(n24606) );
  AND U15577 ( .A(n42889), .B(n24606), .Z(n57326) );
  XNOR U15578 ( .A(x[4998]), .B(y[4998]), .Z(n24610) );
  NANDN U15579 ( .A(y[4996]), .B(x[4996]), .Z(n9634) );
  NANDN U15580 ( .A(y[4997]), .B(x[4997]), .Z(n24609) );
  NAND U15581 ( .A(n9634), .B(n24609), .Z(n57322) );
  XNOR U15582 ( .A(y[4996]), .B(x[4996]), .Z(n42881) );
  ANDN U15583 ( .B(y[4995]), .A(x[4995]), .Z(n42876) );
  NANDN U15584 ( .A(y[4994]), .B(x[4994]), .Z(n24611) );
  ANDN U15585 ( .B(x[4995]), .A(y[4995]), .Z(n42882) );
  ANDN U15586 ( .B(n24611), .A(n42882), .Z(n57319) );
  ANDN U15587 ( .B(y[4993]), .A(x[4993]), .Z(n24613) );
  NANDN U15588 ( .A(x[4994]), .B(y[4994]), .Z(n42877) );
  NANDN U15589 ( .A(n24613), .B(n42877), .Z(n57318) );
  NANDN U15590 ( .A(y[4992]), .B(x[4992]), .Z(n9635) );
  NANDN U15591 ( .A(y[4993]), .B(x[4993]), .Z(n24612) );
  AND U15592 ( .A(n9635), .B(n24612), .Z(n57317) );
  ANDN U15593 ( .B(y[4991]), .A(x[4991]), .Z(n42865) );
  XNOR U15594 ( .A(x[4992]), .B(y[4992]), .Z(n42869) );
  NANDN U15595 ( .A(y[4990]), .B(x[4990]), .Z(n9636) );
  NANDN U15596 ( .A(y[4991]), .B(x[4991]), .Z(n42868) );
  NAND U15597 ( .A(n9636), .B(n42868), .Z(n57313) );
  XNOR U15598 ( .A(x[4990]), .B(y[4990]), .Z(n24615) );
  ANDN U15599 ( .B(y[4989]), .A(x[4989]), .Z(n57311) );
  NANDN U15600 ( .A(x[4987]), .B(y[4987]), .Z(n57310) );
  XNOR U15601 ( .A(x[4988]), .B(y[4988]), .Z(n42858) );
  AND U15602 ( .A(n57310), .B(n42858), .Z(n17001) );
  XNOR U15603 ( .A(x[4986]), .B(y[4986]), .Z(n24617) );
  XNOR U15604 ( .A(x[4984]), .B(y[4984]), .Z(n42848) );
  NANDN U15605 ( .A(y[4982]), .B(x[4982]), .Z(n9637) );
  NANDN U15606 ( .A(y[4983]), .B(x[4983]), .Z(n42847) );
  NAND U15607 ( .A(n9637), .B(n42847), .Z(n57302) );
  XNOR U15608 ( .A(x[4982]), .B(y[4982]), .Z(n24619) );
  ANDN U15609 ( .B(y[4981]), .A(x[4981]), .Z(n57299) );
  NANDN U15610 ( .A(y[4980]), .B(x[4980]), .Z(n9638) );
  NANDN U15611 ( .A(y[4981]), .B(x[4981]), .Z(n24618) );
  AND U15612 ( .A(n9638), .B(n24618), .Z(n57298) );
  NANDN U15613 ( .A(x[4979]), .B(y[4979]), .Z(n51511) );
  XNOR U15614 ( .A(x[4980]), .B(y[4980]), .Z(n42838) );
  NAND U15615 ( .A(n51511), .B(n42838), .Z(n16987) );
  NANDN U15616 ( .A(y[4978]), .B(x[4978]), .Z(n9639) );
  NANDN U15617 ( .A(y[4979]), .B(x[4979]), .Z(n42837) );
  AND U15618 ( .A(n9639), .B(n42837), .Z(n57295) );
  NANDN U15619 ( .A(y[4974]), .B(x[4974]), .Z(n9640) );
  NANDN U15620 ( .A(y[4975]), .B(x[4975]), .Z(n24625) );
  AND U15621 ( .A(n9640), .B(n24625), .Z(n57293) );
  XNOR U15622 ( .A(y[4974]), .B(x[4974]), .Z(n24629) );
  NANDN U15623 ( .A(x[4973]), .B(y[4973]), .Z(n24630) );
  NAND U15624 ( .A(n24629), .B(n24630), .Z(n57292) );
  NANDN U15625 ( .A(y[4972]), .B(x[4972]), .Z(n24632) );
  NANDN U15626 ( .A(y[4973]), .B(x[4973]), .Z(n24628) );
  AND U15627 ( .A(n24632), .B(n24628), .Z(n57291) );
  NANDN U15628 ( .A(x[4971]), .B(y[4971]), .Z(n24634) );
  NANDN U15629 ( .A(x[4972]), .B(y[4972]), .Z(n24631) );
  NAND U15630 ( .A(n24634), .B(n24631), .Z(n57290) );
  NANDN U15631 ( .A(y[4970]), .B(x[4970]), .Z(n9641) );
  NANDN U15632 ( .A(y[4971]), .B(x[4971]), .Z(n24633) );
  AND U15633 ( .A(n9641), .B(n24633), .Z(n57289) );
  NANDN U15634 ( .A(y[4968]), .B(x[4968]), .Z(n24638) );
  NANDN U15635 ( .A(y[4969]), .B(x[4969]), .Z(n24635) );
  AND U15636 ( .A(n24638), .B(n24635), .Z(n57286) );
  NANDN U15637 ( .A(x[4967]), .B(y[4967]), .Z(n42809) );
  NANDN U15638 ( .A(x[4968]), .B(y[4968]), .Z(n24637) );
  AND U15639 ( .A(n42809), .B(n24637), .Z(n57285) );
  NANDN U15640 ( .A(y[4966]), .B(x[4966]), .Z(n9642) );
  NANDN U15641 ( .A(y[4967]), .B(x[4967]), .Z(n24639) );
  AND U15642 ( .A(n9642), .B(n24639), .Z(n57284) );
  ANDN U15643 ( .B(y[4965]), .A(x[4965]), .Z(n57280) );
  XNOR U15644 ( .A(x[4966]), .B(y[4966]), .Z(n24641) );
  NANDN U15645 ( .A(y[4964]), .B(x[4964]), .Z(n9643) );
  NANDN U15646 ( .A(y[4965]), .B(x[4965]), .Z(n24640) );
  NAND U15647 ( .A(n9643), .B(n24640), .Z(n57279) );
  XNOR U15648 ( .A(x[4964]), .B(y[4964]), .Z(n42802) );
  ANDN U15649 ( .B(y[4963]), .A(x[4963]), .Z(n42798) );
  NANDN U15650 ( .A(y[4962]), .B(x[4962]), .Z(n9644) );
  NANDN U15651 ( .A(y[4963]), .B(x[4963]), .Z(n42801) );
  AND U15652 ( .A(n9644), .B(n42801), .Z(n57276) );
  NANDN U15653 ( .A(x[4961]), .B(y[4961]), .Z(n51516) );
  XNOR U15654 ( .A(x[4962]), .B(y[4962]), .Z(n24643) );
  AND U15655 ( .A(n51516), .B(n24643), .Z(n16965) );
  XNOR U15656 ( .A(x[4960]), .B(y[4960]), .Z(n24645) );
  NANDN U15657 ( .A(y[4958]), .B(x[4958]), .Z(n9645) );
  NANDN U15658 ( .A(y[4959]), .B(x[4959]), .Z(n24644) );
  NAND U15659 ( .A(n9645), .B(n24644), .Z(n57274) );
  XNOR U15660 ( .A(x[4958]), .B(y[4958]), .Z(n24647) );
  NANDN U15661 ( .A(y[4956]), .B(x[4956]), .Z(n9646) );
  NANDN U15662 ( .A(y[4957]), .B(x[4957]), .Z(n24646) );
  NAND U15663 ( .A(n9646), .B(n24646), .Z(n57271) );
  XNOR U15664 ( .A(x[4956]), .B(y[4956]), .Z(n42783) );
  ANDN U15665 ( .B(y[4955]), .A(x[4955]), .Z(n42779) );
  NANDN U15666 ( .A(x[4953]), .B(y[4953]), .Z(n57266) );
  NANDN U15667 ( .A(y[4952]), .B(x[4952]), .Z(n24651) );
  NANDN U15668 ( .A(y[4953]), .B(x[4953]), .Z(n24648) );
  AND U15669 ( .A(n24651), .B(n24648), .Z(n57264) );
  NANDN U15670 ( .A(x[4951]), .B(y[4951]), .Z(n24653) );
  NANDN U15671 ( .A(x[4952]), .B(y[4952]), .Z(n24650) );
  NAND U15672 ( .A(n24653), .B(n24650), .Z(n57263) );
  NANDN U15673 ( .A(y[4950]), .B(x[4950]), .Z(n9647) );
  NANDN U15674 ( .A(y[4951]), .B(x[4951]), .Z(n24652) );
  AND U15675 ( .A(n9647), .B(n24652), .Z(n57262) );
  ANDN U15676 ( .B(y[4949]), .A(x[4949]), .Z(n57261) );
  XNOR U15677 ( .A(x[4950]), .B(y[4950]), .Z(n24655) );
  NANDN U15678 ( .A(y[4948]), .B(x[4948]), .Z(n9648) );
  NANDN U15679 ( .A(y[4949]), .B(x[4949]), .Z(n24654) );
  NAND U15680 ( .A(n9648), .B(n24654), .Z(n57260) );
  XNOR U15681 ( .A(x[4948]), .B(y[4948]), .Z(n42764) );
  NANDN U15682 ( .A(x[4947]), .B(y[4947]), .Z(n57259) );
  NANDN U15683 ( .A(y[4946]), .B(x[4946]), .Z(n9649) );
  NANDN U15684 ( .A(y[4947]), .B(x[4947]), .Z(n42763) );
  AND U15685 ( .A(n9649), .B(n42763), .Z(n57257) );
  ANDN U15686 ( .B(y[4945]), .A(x[4945]), .Z(n51521) );
  XNOR U15687 ( .A(x[4946]), .B(y[4946]), .Z(n24657) );
  NANDN U15688 ( .A(n51521), .B(n24657), .Z(n16957) );
  NANDN U15689 ( .A(y[4944]), .B(x[4944]), .Z(n9650) );
  NANDN U15690 ( .A(y[4945]), .B(x[4945]), .Z(n24656) );
  AND U15691 ( .A(n9650), .B(n24656), .Z(n57256) );
  XNOR U15692 ( .A(x[4944]), .B(y[4944]), .Z(n42754) );
  NANDN U15693 ( .A(x[4943]), .B(y[4943]), .Z(n57254) );
  XNOR U15694 ( .A(x[4942]), .B(y[4942]), .Z(n24659) );
  NANDN U15695 ( .A(y[4940]), .B(x[4940]), .Z(n9651) );
  NANDN U15696 ( .A(y[4941]), .B(x[4941]), .Z(n24658) );
  NAND U15697 ( .A(n9651), .B(n24658), .Z(n57249) );
  XOR U15698 ( .A(x[4940]), .B(y[4940]), .Z(n42745) );
  NANDN U15699 ( .A(x[4939]), .B(y[4939]), .Z(n57248) );
  NANDN U15700 ( .A(y[4938]), .B(x[4938]), .Z(n24661) );
  ANDN U15701 ( .B(x[4939]), .A(y[4939]), .Z(n42744) );
  ANDN U15702 ( .B(n24661), .A(n42744), .Z(n57246) );
  NANDN U15703 ( .A(x[4937]), .B(y[4937]), .Z(n42737) );
  NANDN U15704 ( .A(x[4938]), .B(y[4938]), .Z(n24660) );
  NAND U15705 ( .A(n42737), .B(n24660), .Z(n57245) );
  NANDN U15706 ( .A(y[4936]), .B(x[4936]), .Z(n9652) );
  NANDN U15707 ( .A(y[4937]), .B(x[4937]), .Z(n24662) );
  AND U15708 ( .A(n9652), .B(n24662), .Z(n57244) );
  ANDN U15709 ( .B(y[4935]), .A(x[4935]), .Z(n24665) );
  XNOR U15710 ( .A(x[4936]), .B(y[4936]), .Z(n24664) );
  NANDN U15711 ( .A(y[4934]), .B(x[4934]), .Z(n9653) );
  NANDN U15712 ( .A(y[4935]), .B(x[4935]), .Z(n24663) );
  NAND U15713 ( .A(n9653), .B(n24663), .Z(n57242) );
  XNOR U15714 ( .A(x[4934]), .B(y[4934]), .Z(n24667) );
  NANDN U15715 ( .A(x[4933]), .B(y[4933]), .Z(n57240) );
  AND U15716 ( .A(n24667), .B(n57240), .Z(n16939) );
  NANDN U15717 ( .A(x[4932]), .B(y[4932]), .Z(n24668) );
  ANDN U15718 ( .B(y[4931]), .A(x[4931]), .Z(n42724) );
  ANDN U15719 ( .B(n24668), .A(n42724), .Z(n57238) );
  XNOR U15720 ( .A(x[4930]), .B(y[4930]), .Z(n24672) );
  NANDN U15721 ( .A(y[4928]), .B(x[4928]), .Z(n9654) );
  NANDN U15722 ( .A(y[4929]), .B(x[4929]), .Z(n24671) );
  NAND U15723 ( .A(n9654), .B(n24671), .Z(n57234) );
  XNOR U15724 ( .A(x[4928]), .B(y[4928]), .Z(n24674) );
  NANDN U15725 ( .A(y[4926]), .B(x[4926]), .Z(n9655) );
  NANDN U15726 ( .A(y[4927]), .B(x[4927]), .Z(n24673) );
  NAND U15727 ( .A(n9655), .B(n24673), .Z(n57231) );
  XNOR U15728 ( .A(x[4926]), .B(y[4926]), .Z(n24676) );
  ANDN U15729 ( .B(y[4925]), .A(x[4925]), .Z(n42710) );
  XNOR U15730 ( .A(x[4924]), .B(y[4924]), .Z(n42708) );
  NANDN U15731 ( .A(x[4923]), .B(y[4923]), .Z(n57228) );
  AND U15732 ( .A(n42708), .B(n57228), .Z(n16923) );
  NANDN U15733 ( .A(y[4920]), .B(x[4920]), .Z(n24682) );
  NANDN U15734 ( .A(y[4921]), .B(x[4921]), .Z(n24679) );
  NAND U15735 ( .A(n24682), .B(n24679), .Z(n57224) );
  NANDN U15736 ( .A(x[4919]), .B(y[4919]), .Z(n42696) );
  NANDN U15737 ( .A(x[4920]), .B(y[4920]), .Z(n24681) );
  AND U15738 ( .A(n42696), .B(n24681), .Z(n51528) );
  XNOR U15739 ( .A(x[4918]), .B(y[4918]), .Z(n24685) );
  NANDN U15740 ( .A(x[4917]), .B(y[4917]), .Z(n57223) );
  AND U15741 ( .A(n24685), .B(n57223), .Z(n16915) );
  NANDN U15742 ( .A(x[4915]), .B(y[4915]), .Z(n57220) );
  XNOR U15743 ( .A(x[4916]), .B(y[4916]), .Z(n24687) );
  AND U15744 ( .A(n57220), .B(n24687), .Z(n16911) );
  NANDN U15745 ( .A(y[4914]), .B(x[4914]), .Z(n9656) );
  NANDN U15746 ( .A(y[4915]), .B(x[4915]), .Z(n24686) );
  NAND U15747 ( .A(n9656), .B(n24686), .Z(n57219) );
  XNOR U15748 ( .A(x[4914]), .B(y[4914]), .Z(n24689) );
  ANDN U15749 ( .B(x[4912]), .A(y[4912]), .Z(n42680) );
  NANDN U15750 ( .A(y[4913]), .B(x[4913]), .Z(n24688) );
  NANDN U15751 ( .A(n42680), .B(n24688), .Z(n57216) );
  NANDN U15752 ( .A(x[4909]), .B(y[4909]), .Z(n24695) );
  NANDN U15753 ( .A(x[4910]), .B(y[4910]), .Z(n24692) );
  NAND U15754 ( .A(n24695), .B(n24692), .Z(n57212) );
  NANDN U15755 ( .A(y[4908]), .B(x[4908]), .Z(n24697) );
  NANDN U15756 ( .A(y[4909]), .B(x[4909]), .Z(n24694) );
  AND U15757 ( .A(n24697), .B(n24694), .Z(n51531) );
  ANDN U15758 ( .B(y[4905]), .A(x[4905]), .Z(n24702) );
  XNOR U15759 ( .A(x[4906]), .B(y[4906]), .Z(n24701) );
  NANDN U15760 ( .A(y[4905]), .B(x[4905]), .Z(n24700) );
  ANDN U15761 ( .B(x[4904]), .A(y[4904]), .Z(n42662) );
  ANDN U15762 ( .B(n24700), .A(n42662), .Z(n57210) );
  NANDN U15763 ( .A(x[4903]), .B(y[4903]), .Z(n24704) );
  NANDN U15764 ( .A(x[4904]), .B(y[4904]), .Z(n24703) );
  NAND U15765 ( .A(n24704), .B(n24703), .Z(n57209) );
  NANDN U15766 ( .A(y[4902]), .B(x[4902]), .Z(n24706) );
  NANDN U15767 ( .A(y[4903]), .B(x[4903]), .Z(n42663) );
  AND U15768 ( .A(n24706), .B(n42663), .Z(n57208) );
  NANDN U15769 ( .A(x[4901]), .B(y[4901]), .Z(n24708) );
  NANDN U15770 ( .A(x[4902]), .B(y[4902]), .Z(n24705) );
  NAND U15771 ( .A(n24708), .B(n24705), .Z(n57207) );
  NANDN U15772 ( .A(y[4901]), .B(x[4901]), .Z(n24707) );
  ANDN U15773 ( .B(x[4900]), .A(y[4900]), .Z(n42652) );
  ANDN U15774 ( .B(n24707), .A(n42652), .Z(n57206) );
  NANDN U15775 ( .A(y[4898]), .B(x[4898]), .Z(n24712) );
  NANDN U15776 ( .A(y[4899]), .B(x[4899]), .Z(n42653) );
  AND U15777 ( .A(n24712), .B(n42653), .Z(n57204) );
  NANDN U15778 ( .A(x[4897]), .B(y[4897]), .Z(n24714) );
  NANDN U15779 ( .A(x[4898]), .B(y[4898]), .Z(n24711) );
  NAND U15780 ( .A(n24714), .B(n24711), .Z(n57202) );
  NANDN U15781 ( .A(y[4897]), .B(x[4897]), .Z(n24713) );
  ANDN U15782 ( .B(x[4896]), .A(y[4896]), .Z(n42642) );
  ANDN U15783 ( .B(n24713), .A(n42642), .Z(n57201) );
  NANDN U15784 ( .A(x[4893]), .B(y[4893]), .Z(n24720) );
  NANDN U15785 ( .A(x[4894]), .B(y[4894]), .Z(n24717) );
  NAND U15786 ( .A(n24720), .B(n24717), .Z(n57198) );
  NANDN U15787 ( .A(x[4891]), .B(y[4891]), .Z(n24722) );
  NANDN U15788 ( .A(x[4892]), .B(y[4892]), .Z(n24721) );
  AND U15789 ( .A(n24722), .B(n24721), .Z(n57196) );
  NANDN U15790 ( .A(y[4890]), .B(x[4890]), .Z(n24724) );
  NANDN U15791 ( .A(y[4891]), .B(x[4891]), .Z(n42633) );
  NAND U15792 ( .A(n24724), .B(n42633), .Z(n57195) );
  NANDN U15793 ( .A(x[4889]), .B(y[4889]), .Z(n24726) );
  NANDN U15794 ( .A(x[4890]), .B(y[4890]), .Z(n24723) );
  AND U15795 ( .A(n24726), .B(n24723), .Z(n57194) );
  NANDN U15796 ( .A(y[4888]), .B(x[4888]), .Z(n24728) );
  NANDN U15797 ( .A(y[4889]), .B(x[4889]), .Z(n24725) );
  NAND U15798 ( .A(n24728), .B(n24725), .Z(n57193) );
  NANDN U15799 ( .A(x[4887]), .B(y[4887]), .Z(n42621) );
  NANDN U15800 ( .A(x[4888]), .B(y[4888]), .Z(n24727) );
  AND U15801 ( .A(n42621), .B(n24727), .Z(n57192) );
  XNOR U15802 ( .A(x[4886]), .B(y[4886]), .Z(n24731) );
  NANDN U15803 ( .A(x[4883]), .B(y[4883]), .Z(n24735) );
  NANDN U15804 ( .A(x[4884]), .B(y[4884]), .Z(n24732) );
  AND U15805 ( .A(n24735), .B(n24732), .Z(n57187) );
  XNOR U15806 ( .A(y[4882]), .B(x[4882]), .Z(n24738) );
  NANDN U15807 ( .A(x[4881]), .B(y[4881]), .Z(n42606) );
  AND U15808 ( .A(n24738), .B(n42606), .Z(n57184) );
  NANDN U15809 ( .A(y[4880]), .B(x[4880]), .Z(n9657) );
  NANDN U15810 ( .A(y[4881]), .B(x[4881]), .Z(n24737) );
  AND U15811 ( .A(n9657), .B(n24737), .Z(n51535) );
  XNOR U15812 ( .A(y[4880]), .B(x[4880]), .Z(n24740) );
  NANDN U15813 ( .A(x[4879]), .B(y[4879]), .Z(n24741) );
  NAND U15814 ( .A(n24740), .B(n24741), .Z(n51536) );
  NANDN U15815 ( .A(y[4878]), .B(x[4878]), .Z(n9658) );
  NANDN U15816 ( .A(y[4879]), .B(x[4879]), .Z(n24739) );
  AND U15817 ( .A(n9658), .B(n24739), .Z(n57182) );
  NANDN U15818 ( .A(x[4873]), .B(y[4873]), .Z(n57175) );
  XNOR U15819 ( .A(x[4874]), .B(y[4874]), .Z(n24749) );
  AND U15820 ( .A(n57175), .B(n24749), .Z(n16859) );
  NANDN U15821 ( .A(y[4872]), .B(x[4872]), .Z(n9659) );
  NANDN U15822 ( .A(y[4873]), .B(x[4873]), .Z(n24748) );
  NAND U15823 ( .A(n9659), .B(n24748), .Z(n57174) );
  XNOR U15824 ( .A(x[4872]), .B(y[4872]), .Z(n24751) );
  XNOR U15825 ( .A(x[4870]), .B(y[4870]), .Z(n24753) );
  NANDN U15826 ( .A(y[4868]), .B(x[4868]), .Z(n9660) );
  NANDN U15827 ( .A(y[4869]), .B(x[4869]), .Z(n24752) );
  NAND U15828 ( .A(n9660), .B(n24752), .Z(n57167) );
  XNOR U15829 ( .A(x[4868]), .B(y[4868]), .Z(n42579) );
  ANDN U15830 ( .B(y[4867]), .A(x[4867]), .Z(n24754) );
  NANDN U15831 ( .A(y[4866]), .B(x[4866]), .Z(n9661) );
  ANDN U15832 ( .B(x[4867]), .A(y[4867]), .Z(n42578) );
  ANDN U15833 ( .B(n9661), .A(n42578), .Z(n57164) );
  XNOR U15834 ( .A(x[4866]), .B(y[4866]), .Z(n24756) );
  ANDN U15835 ( .B(y[4865]), .A(x[4865]), .Z(n42570) );
  ANDN U15836 ( .B(n24756), .A(n42570), .Z(n16846) );
  XNOR U15837 ( .A(x[4864]), .B(y[4864]), .Z(n24758) );
  NANDN U15838 ( .A(y[4862]), .B(x[4862]), .Z(n9662) );
  NANDN U15839 ( .A(y[4863]), .B(x[4863]), .Z(n24757) );
  NAND U15840 ( .A(n9662), .B(n24757), .Z(n57159) );
  XNOR U15841 ( .A(x[4862]), .B(y[4862]), .Z(n24760) );
  NANDN U15842 ( .A(y[4860]), .B(x[4860]), .Z(n9663) );
  NANDN U15843 ( .A(y[4861]), .B(x[4861]), .Z(n24759) );
  NAND U15844 ( .A(n9663), .B(n24759), .Z(n57158) );
  XNOR U15845 ( .A(x[4860]), .B(y[4860]), .Z(n24762) );
  ANDN U15846 ( .B(y[4859]), .A(x[4859]), .Z(n42557) );
  NANDN U15847 ( .A(x[4857]), .B(y[4857]), .Z(n57152) );
  XNOR U15848 ( .A(x[4858]), .B(y[4858]), .Z(n24764) );
  AND U15849 ( .A(n57152), .B(n24764), .Z(n16832) );
  NANDN U15850 ( .A(y[4856]), .B(x[4856]), .Z(n9664) );
  NANDN U15851 ( .A(y[4857]), .B(x[4857]), .Z(n24763) );
  NAND U15852 ( .A(n9664), .B(n24763), .Z(n57151) );
  XNOR U15853 ( .A(x[4856]), .B(y[4856]), .Z(n24766) );
  XNOR U15854 ( .A(x[4854]), .B(y[4854]), .Z(n24768) );
  NANDN U15855 ( .A(y[4852]), .B(x[4852]), .Z(n24770) );
  NANDN U15856 ( .A(y[4853]), .B(x[4853]), .Z(n24767) );
  NAND U15857 ( .A(n24770), .B(n24767), .Z(n57147) );
  NANDN U15858 ( .A(x[4851]), .B(y[4851]), .Z(n42541) );
  NANDN U15859 ( .A(x[4852]), .B(y[4852]), .Z(n24769) );
  AND U15860 ( .A(n42541), .B(n24769), .Z(n57146) );
  NANDN U15861 ( .A(y[4850]), .B(x[4850]), .Z(n9665) );
  NANDN U15862 ( .A(y[4851]), .B(x[4851]), .Z(n24771) );
  NAND U15863 ( .A(n9665), .B(n24771), .Z(n57145) );
  XNOR U15864 ( .A(x[4850]), .B(y[4850]), .Z(n24773) );
  NANDN U15865 ( .A(x[4849]), .B(y[4849]), .Z(n57143) );
  AND U15866 ( .A(n24773), .B(n57143), .Z(n16820) );
  NANDN U15867 ( .A(x[4847]), .B(y[4847]), .Z(n42531) );
  NANDN U15868 ( .A(x[4848]), .B(y[4848]), .Z(n24774) );
  AND U15869 ( .A(n42531), .B(n24774), .Z(n57138) );
  NANDN U15870 ( .A(y[4846]), .B(x[4846]), .Z(n9666) );
  NANDN U15871 ( .A(y[4847]), .B(x[4847]), .Z(n24776) );
  NAND U15872 ( .A(n9666), .B(n24776), .Z(n57137) );
  XNOR U15873 ( .A(x[4846]), .B(y[4846]), .Z(n24778) );
  ANDN U15874 ( .B(y[4845]), .A(x[4845]), .Z(n42526) );
  NANDN U15875 ( .A(x[4843]), .B(y[4843]), .Z(n57132) );
  XNOR U15876 ( .A(x[4844]), .B(y[4844]), .Z(n24780) );
  AND U15877 ( .A(n57132), .B(n24780), .Z(n16811) );
  NANDN U15878 ( .A(y[4842]), .B(x[4842]), .Z(n9667) );
  NANDN U15879 ( .A(y[4843]), .B(x[4843]), .Z(n24779) );
  NAND U15880 ( .A(n9667), .B(n24779), .Z(n57131) );
  XNOR U15881 ( .A(x[4842]), .B(y[4842]), .Z(n24782) );
  ANDN U15882 ( .B(x[4839]), .A(y[4839]), .Z(n42515) );
  NANDN U15883 ( .A(y[4838]), .B(x[4838]), .Z(n9668) );
  NANDN U15884 ( .A(n42515), .B(n9668), .Z(n51545) );
  XNOR U15885 ( .A(y[4838]), .B(x[4838]), .Z(n24785) );
  NANDN U15886 ( .A(x[4837]), .B(y[4837]), .Z(n42507) );
  AND U15887 ( .A(n24785), .B(n42507), .Z(n57126) );
  NANDN U15888 ( .A(y[4836]), .B(x[4836]), .Z(n9669) );
  NANDN U15889 ( .A(y[4837]), .B(x[4837]), .Z(n24784) );
  NAND U15890 ( .A(n9669), .B(n24784), .Z(n57124) );
  XNOR U15891 ( .A(x[4836]), .B(y[4836]), .Z(n24787) );
  NANDN U15892 ( .A(x[4835]), .B(y[4835]), .Z(n57123) );
  AND U15893 ( .A(n24787), .B(n57123), .Z(n16799) );
  XNOR U15894 ( .A(y[4834]), .B(x[4834]), .Z(n24790) );
  NANDN U15895 ( .A(x[4833]), .B(y[4833]), .Z(n42497) );
  AND U15896 ( .A(n24790), .B(n42497), .Z(n57120) );
  NANDN U15897 ( .A(y[4832]), .B(x[4832]), .Z(n9670) );
  NANDN U15898 ( .A(y[4833]), .B(x[4833]), .Z(n24789) );
  NAND U15899 ( .A(n9670), .B(n24789), .Z(n57119) );
  XNOR U15900 ( .A(y[4832]), .B(x[4832]), .Z(n24792) );
  NANDN U15901 ( .A(x[4831]), .B(y[4831]), .Z(n24793) );
  AND U15902 ( .A(n24792), .B(n24793), .Z(n57118) );
  NANDN U15903 ( .A(y[4830]), .B(x[4830]), .Z(n9671) );
  NANDN U15904 ( .A(y[4831]), .B(x[4831]), .Z(n24791) );
  NAND U15905 ( .A(n9671), .B(n24791), .Z(n57117) );
  XNOR U15906 ( .A(y[4830]), .B(x[4830]), .Z(n24796) );
  NANDN U15907 ( .A(x[4829]), .B(y[4829]), .Z(n42488) );
  AND U15908 ( .A(n24796), .B(n42488), .Z(n57116) );
  XNOR U15909 ( .A(x[4828]), .B(y[4828]), .Z(n24798) );
  NANDN U15910 ( .A(y[4826]), .B(x[4826]), .Z(n9672) );
  NANDN U15911 ( .A(y[4827]), .B(x[4827]), .Z(n24797) );
  NAND U15912 ( .A(n9672), .B(n24797), .Z(n57114) );
  XNOR U15913 ( .A(y[4826]), .B(x[4826]), .Z(n24801) );
  NANDN U15914 ( .A(x[4825]), .B(y[4825]), .Z(n24802) );
  AND U15915 ( .A(n24801), .B(n24802), .Z(n57113) );
  NANDN U15916 ( .A(y[4822]), .B(x[4822]), .Z(n9673) );
  NANDN U15917 ( .A(y[4823]), .B(x[4823]), .Z(n24805) );
  NAND U15918 ( .A(n9673), .B(n24805), .Z(n57108) );
  XNOR U15919 ( .A(x[4822]), .B(y[4822]), .Z(n24807) );
  ANDN U15920 ( .B(x[4820]), .A(y[4820]), .Z(n42468) );
  NANDN U15921 ( .A(y[4821]), .B(x[4821]), .Z(n24806) );
  NANDN U15922 ( .A(n42468), .B(n24806), .Z(n57107) );
  NANDN U15923 ( .A(x[4819]), .B(y[4819]), .Z(n24809) );
  NANDN U15924 ( .A(x[4820]), .B(y[4820]), .Z(n24808) );
  AND U15925 ( .A(n24809), .B(n24808), .Z(n57106) );
  NANDN U15926 ( .A(y[4818]), .B(x[4818]), .Z(n24811) );
  NANDN U15927 ( .A(y[4819]), .B(x[4819]), .Z(n42469) );
  NAND U15928 ( .A(n24811), .B(n42469), .Z(n57105) );
  NANDN U15929 ( .A(x[4817]), .B(y[4817]), .Z(n24813) );
  XNOR U15930 ( .A(x[4818]), .B(y[4818]), .Z(n9674) );
  AND U15931 ( .A(n24813), .B(n9674), .Z(n57104) );
  ANDN U15932 ( .B(x[4816]), .A(y[4816]), .Z(n42458) );
  NANDN U15933 ( .A(y[4817]), .B(x[4817]), .Z(n24812) );
  NANDN U15934 ( .A(n42458), .B(n24812), .Z(n57103) );
  NANDN U15935 ( .A(x[4813]), .B(y[4813]), .Z(n24819) );
  NANDN U15936 ( .A(x[4814]), .B(y[4814]), .Z(n24816) );
  NAND U15937 ( .A(n24819), .B(n24816), .Z(n57100) );
  NANDN U15938 ( .A(y[4812]), .B(x[4812]), .Z(n24822) );
  NANDN U15939 ( .A(y[4813]), .B(x[4813]), .Z(n24818) );
  AND U15940 ( .A(n24822), .B(n24818), .Z(n51550) );
  XNOR U15941 ( .A(x[4810]), .B(y[4810]), .Z(n42444) );
  NANDN U15942 ( .A(x[4809]), .B(y[4809]), .Z(n51554) );
  NAND U15943 ( .A(n42444), .B(n51554), .Z(n16766) );
  XNOR U15944 ( .A(x[4808]), .B(y[4808]), .Z(n24823) );
  NANDN U15945 ( .A(x[4807]), .B(y[4807]), .Z(n24825) );
  AND U15946 ( .A(n24823), .B(n24825), .Z(n16762) );
  ANDN U15947 ( .B(y[4805]), .A(x[4805]), .Z(n24828) );
  NANDN U15948 ( .A(y[4804]), .B(x[4804]), .Z(n57092) );
  NANDN U15949 ( .A(x[4803]), .B(y[4803]), .Z(n24832) );
  NANDN U15950 ( .A(x[4804]), .B(y[4804]), .Z(n24829) );
  NAND U15951 ( .A(n24832), .B(n24829), .Z(n57091) );
  NANDN U15952 ( .A(y[4802]), .B(x[4802]), .Z(n24833) );
  NANDN U15953 ( .A(y[4803]), .B(x[4803]), .Z(n24830) );
  AND U15954 ( .A(n24833), .B(n24830), .Z(n57090) );
  NANDN U15955 ( .A(x[4801]), .B(y[4801]), .Z(n24835) );
  NANDN U15956 ( .A(x[4802]), .B(y[4802]), .Z(n24831) );
  NAND U15957 ( .A(n24835), .B(n24831), .Z(n57089) );
  NANDN U15958 ( .A(y[4800]), .B(x[4800]), .Z(n42422) );
  NANDN U15959 ( .A(y[4801]), .B(x[4801]), .Z(n24834) );
  AND U15960 ( .A(n42422), .B(n24834), .Z(n57088) );
  NANDN U15961 ( .A(x[4799]), .B(y[4799]), .Z(n24837) );
  NANDN U15962 ( .A(x[4800]), .B(y[4800]), .Z(n24836) );
  NAND U15963 ( .A(n24837), .B(n24836), .Z(n57087) );
  NANDN U15964 ( .A(y[4798]), .B(x[4798]), .Z(n42416) );
  NANDN U15965 ( .A(y[4799]), .B(x[4799]), .Z(n42423) );
  AND U15966 ( .A(n42416), .B(n42423), .Z(n57086) );
  NANDN U15967 ( .A(x[4797]), .B(y[4797]), .Z(n24839) );
  NANDN U15968 ( .A(x[4798]), .B(y[4798]), .Z(n24838) );
  NAND U15969 ( .A(n24839), .B(n24838), .Z(n57085) );
  NANDN U15970 ( .A(y[4796]), .B(x[4796]), .Z(n42411) );
  NANDN U15971 ( .A(y[4797]), .B(x[4797]), .Z(n42417) );
  AND U15972 ( .A(n42411), .B(n42417), .Z(n57084) );
  NANDN U15973 ( .A(x[4793]), .B(y[4793]), .Z(n24842) );
  NANDN U15974 ( .A(x[4794]), .B(y[4794]), .Z(n24841) );
  NAND U15975 ( .A(n24842), .B(n24841), .Z(n57079) );
  NANDN U15976 ( .A(y[4792]), .B(x[4792]), .Z(n9675) );
  NANDN U15977 ( .A(y[4793]), .B(x[4793]), .Z(n42406) );
  AND U15978 ( .A(n9675), .B(n42406), .Z(n51558) );
  XNOR U15979 ( .A(y[4792]), .B(x[4792]), .Z(n42401) );
  NANDN U15980 ( .A(x[4791]), .B(y[4791]), .Z(n24844) );
  AND U15981 ( .A(n42401), .B(n24844), .Z(n57078) );
  NANDN U15982 ( .A(y[4790]), .B(x[4790]), .Z(n9676) );
  NANDN U15983 ( .A(y[4791]), .B(x[4791]), .Z(n42400) );
  NAND U15984 ( .A(n9676), .B(n42400), .Z(n57077) );
  XNOR U15985 ( .A(y[4790]), .B(x[4790]), .Z(n42395) );
  NANDN U15986 ( .A(x[4789]), .B(y[4789]), .Z(n24846) );
  AND U15987 ( .A(n42395), .B(n24846), .Z(n57076) );
  NANDN U15988 ( .A(y[4788]), .B(x[4788]), .Z(n9677) );
  NANDN U15989 ( .A(y[4789]), .B(x[4789]), .Z(n42394) );
  NAND U15990 ( .A(n9677), .B(n42394), .Z(n57075) );
  XNOR U15991 ( .A(y[4788]), .B(x[4788]), .Z(n42389) );
  NANDN U15992 ( .A(x[4787]), .B(y[4787]), .Z(n24848) );
  AND U15993 ( .A(n42389), .B(n24848), .Z(n57074) );
  NANDN U15994 ( .A(y[4786]), .B(x[4786]), .Z(n9678) );
  NANDN U15995 ( .A(y[4787]), .B(x[4787]), .Z(n42388) );
  NAND U15996 ( .A(n9678), .B(n42388), .Z(n57073) );
  XNOR U15997 ( .A(y[4784]), .B(x[4784]), .Z(n42377) );
  NANDN U15998 ( .A(x[4783]), .B(y[4783]), .Z(n24852) );
  NAND U15999 ( .A(n42377), .B(n24852), .Z(n57070) );
  NANDN U16000 ( .A(y[4782]), .B(x[4782]), .Z(n9679) );
  NANDN U16001 ( .A(y[4783]), .B(x[4783]), .Z(n42376) );
  AND U16002 ( .A(n9679), .B(n42376), .Z(n51559) );
  XNOR U16003 ( .A(y[4782]), .B(x[4782]), .Z(n42371) );
  NANDN U16004 ( .A(x[4781]), .B(y[4781]), .Z(n42367) );
  AND U16005 ( .A(n42371), .B(n42367), .Z(n57069) );
  NANDN U16006 ( .A(y[4780]), .B(x[4780]), .Z(n9680) );
  NANDN U16007 ( .A(y[4781]), .B(x[4781]), .Z(n42370) );
  NAND U16008 ( .A(n9680), .B(n42370), .Z(n57067) );
  XNOR U16009 ( .A(y[4780]), .B(x[4780]), .Z(n24855) );
  NANDN U16010 ( .A(x[4779]), .B(y[4779]), .Z(n24856) );
  AND U16011 ( .A(n24855), .B(n24856), .Z(n57066) );
  NANDN U16012 ( .A(y[4778]), .B(x[4778]), .Z(n9681) );
  NANDN U16013 ( .A(y[4779]), .B(x[4779]), .Z(n24854) );
  NAND U16014 ( .A(n9681), .B(n24854), .Z(n57065) );
  NANDN U16015 ( .A(x[4777]), .B(y[4777]), .Z(n57063) );
  XNOR U16016 ( .A(x[4778]), .B(y[4778]), .Z(n24858) );
  NANDN U16017 ( .A(y[4776]), .B(x[4776]), .Z(n9682) );
  NANDN U16018 ( .A(y[4777]), .B(x[4777]), .Z(n24857) );
  AND U16019 ( .A(n9682), .B(n24857), .Z(n51560) );
  NANDN U16020 ( .A(x[4775]), .B(y[4775]), .Z(n57062) );
  XNOR U16021 ( .A(x[4776]), .B(y[4776]), .Z(n42355) );
  NANDN U16022 ( .A(y[4774]), .B(x[4774]), .Z(n9683) );
  NANDN U16023 ( .A(y[4775]), .B(x[4775]), .Z(n42354) );
  NAND U16024 ( .A(n9683), .B(n42354), .Z(n57060) );
  XNOR U16025 ( .A(y[4774]), .B(x[4774]), .Z(n42349) );
  NANDN U16026 ( .A(x[4773]), .B(y[4773]), .Z(n24860) );
  AND U16027 ( .A(n42349), .B(n24860), .Z(n57059) );
  NANDN U16028 ( .A(y[4772]), .B(x[4772]), .Z(n9684) );
  NANDN U16029 ( .A(y[4773]), .B(x[4773]), .Z(n42348) );
  NAND U16030 ( .A(n9684), .B(n42348), .Z(n57058) );
  XNOR U16031 ( .A(y[4772]), .B(x[4772]), .Z(n24863) );
  NANDN U16032 ( .A(x[4771]), .B(y[4771]), .Z(n24864) );
  AND U16033 ( .A(n24863), .B(n24864), .Z(n57057) );
  XNOR U16034 ( .A(x[4770]), .B(y[4770]), .Z(n24866) );
  NANDN U16035 ( .A(y[4768]), .B(x[4768]), .Z(n9685) );
  NANDN U16036 ( .A(y[4769]), .B(x[4769]), .Z(n24865) );
  NAND U16037 ( .A(n9685), .B(n24865), .Z(n57051) );
  XNOR U16038 ( .A(y[4768]), .B(x[4768]), .Z(n42335) );
  NANDN U16039 ( .A(x[4767]), .B(y[4767]), .Z(n42332) );
  AND U16040 ( .A(n42335), .B(n42332), .Z(n51561) );
  NANDN U16041 ( .A(x[4765]), .B(y[4765]), .Z(n57048) );
  XNOR U16042 ( .A(x[4766]), .B(y[4766]), .Z(n42328) );
  NANDN U16043 ( .A(y[4764]), .B(x[4764]), .Z(n9686) );
  NANDN U16044 ( .A(y[4765]), .B(x[4765]), .Z(n42327) );
  AND U16045 ( .A(n9686), .B(n42327), .Z(n51564) );
  XNOR U16046 ( .A(y[4760]), .B(x[4760]), .Z(n42310) );
  NANDN U16047 ( .A(x[4759]), .B(y[4759]), .Z(n24873) );
  NAND U16048 ( .A(n42310), .B(n24873), .Z(n57045) );
  NANDN U16049 ( .A(y[4758]), .B(x[4758]), .Z(n9687) );
  NANDN U16050 ( .A(y[4759]), .B(x[4759]), .Z(n42309) );
  AND U16051 ( .A(n9687), .B(n42309), .Z(n57044) );
  XNOR U16052 ( .A(y[4758]), .B(x[4758]), .Z(n42304) );
  NANDN U16053 ( .A(x[4757]), .B(y[4757]), .Z(n24875) );
  NAND U16054 ( .A(n42304), .B(n24875), .Z(n57043) );
  NANDN U16055 ( .A(y[4756]), .B(x[4756]), .Z(n9688) );
  NANDN U16056 ( .A(y[4757]), .B(x[4757]), .Z(n42303) );
  AND U16057 ( .A(n9688), .B(n42303), .Z(n57042) );
  XNOR U16058 ( .A(y[4756]), .B(x[4756]), .Z(n42298) );
  NANDN U16059 ( .A(x[4755]), .B(y[4755]), .Z(n24877) );
  NAND U16060 ( .A(n42298), .B(n24877), .Z(n57040) );
  NANDN U16061 ( .A(y[4752]), .B(x[4752]), .Z(n9689) );
  NANDN U16062 ( .A(y[4753]), .B(x[4753]), .Z(n42291) );
  NAND U16063 ( .A(n9689), .B(n42291), .Z(n57037) );
  XNOR U16064 ( .A(y[4752]), .B(x[4752]), .Z(n42286) );
  NANDN U16065 ( .A(x[4751]), .B(y[4751]), .Z(n24881) );
  AND U16066 ( .A(n42286), .B(n24881), .Z(n51567) );
  XNOR U16067 ( .A(x[4748]), .B(y[4748]), .Z(n24886) );
  NANDN U16068 ( .A(y[4746]), .B(x[4746]), .Z(n24887) );
  NANDN U16069 ( .A(y[4747]), .B(x[4747]), .Z(n24885) );
  NAND U16070 ( .A(n24887), .B(n24885), .Z(n57033) );
  NANDN U16071 ( .A(x[4745]), .B(y[4745]), .Z(n42268) );
  NANDN U16072 ( .A(x[4746]), .B(y[4746]), .Z(n42274) );
  AND U16073 ( .A(n42268), .B(n42274), .Z(n57032) );
  NANDN U16074 ( .A(y[4744]), .B(x[4744]), .Z(n9690) );
  NANDN U16075 ( .A(y[4745]), .B(x[4745]), .Z(n24888) );
  NAND U16076 ( .A(n9690), .B(n24888), .Z(n57031) );
  XNOR U16077 ( .A(x[4744]), .B(y[4744]), .Z(n42266) );
  NANDN U16078 ( .A(x[4743]), .B(y[4743]), .Z(n57028) );
  AND U16079 ( .A(n42266), .B(n57028), .Z(n16680) );
  XNOR U16080 ( .A(y[4742]), .B(x[4742]), .Z(n42259) );
  NANDN U16081 ( .A(x[4741]), .B(y[4741]), .Z(n42253) );
  AND U16082 ( .A(n42259), .B(n42253), .Z(n57026) );
  ANDN U16083 ( .B(x[4741]), .A(y[4741]), .Z(n42258) );
  NANDN U16084 ( .A(y[4740]), .B(x[4740]), .Z(n9691) );
  NANDN U16085 ( .A(n42258), .B(n9691), .Z(n57025) );
  XNOR U16086 ( .A(y[4740]), .B(x[4740]), .Z(n24890) );
  NANDN U16087 ( .A(x[4739]), .B(y[4739]), .Z(n42247) );
  AND U16088 ( .A(n24890), .B(n42247), .Z(n57024) );
  NANDN U16089 ( .A(y[4738]), .B(x[4738]), .Z(n9692) );
  NANDN U16090 ( .A(y[4739]), .B(x[4739]), .Z(n24889) );
  NAND U16091 ( .A(n9692), .B(n24889), .Z(n57023) );
  XNOR U16092 ( .A(y[4738]), .B(x[4738]), .Z(n42245) );
  NANDN U16093 ( .A(x[4737]), .B(y[4737]), .Z(n42239) );
  AND U16094 ( .A(n42245), .B(n42239), .Z(n57022) );
  XNOR U16095 ( .A(y[4736]), .B(x[4736]), .Z(n42237) );
  NANDN U16096 ( .A(x[4735]), .B(y[4735]), .Z(n42231) );
  AND U16097 ( .A(n42237), .B(n42231), .Z(n57020) );
  ANDN U16098 ( .B(x[4735]), .A(y[4735]), .Z(n42236) );
  NANDN U16099 ( .A(y[4734]), .B(x[4734]), .Z(n9693) );
  NANDN U16100 ( .A(n42236), .B(n9693), .Z(n57019) );
  XNOR U16101 ( .A(y[4734]), .B(x[4734]), .Z(n42229) );
  NANDN U16102 ( .A(x[4733]), .B(y[4733]), .Z(n42224) );
  AND U16103 ( .A(n42229), .B(n42224), .Z(n57018) );
  ANDN U16104 ( .B(x[4733]), .A(y[4733]), .Z(n42228) );
  NANDN U16105 ( .A(y[4732]), .B(x[4732]), .Z(n9694) );
  NANDN U16106 ( .A(n42228), .B(n9694), .Z(n57017) );
  NANDN U16107 ( .A(y[4730]), .B(x[4730]), .Z(n9695) );
  NANDN U16108 ( .A(y[4731]), .B(x[4731]), .Z(n24891) );
  AND U16109 ( .A(n9695), .B(n24891), .Z(n51570) );
  XOR U16110 ( .A(x[4730]), .B(y[4730]), .Z(n42219) );
  NANDN U16111 ( .A(y[4728]), .B(x[4728]), .Z(n9696) );
  ANDN U16112 ( .B(x[4729]), .A(y[4729]), .Z(n42217) );
  ANDN U16113 ( .B(n9696), .A(n42217), .Z(n57012) );
  ANDN U16114 ( .B(y[4727]), .A(x[4727]), .Z(n24896) );
  XNOR U16115 ( .A(x[4728]), .B(y[4728]), .Z(n24895) );
  NANDN U16116 ( .A(y[4726]), .B(x[4726]), .Z(n9697) );
  NANDN U16117 ( .A(y[4727]), .B(x[4727]), .Z(n24894) );
  NAND U16118 ( .A(n9697), .B(n24894), .Z(n57009) );
  XNOR U16119 ( .A(x[4726]), .B(y[4726]), .Z(n24898) );
  ANDN U16120 ( .B(y[4725]), .A(x[4725]), .Z(n24899) );
  XNOR U16121 ( .A(x[4724]), .B(y[4724]), .Z(n24901) );
  NANDN U16122 ( .A(x[4723]), .B(y[4723]), .Z(n57005) );
  AND U16123 ( .A(n24901), .B(n57005), .Z(n16652) );
  NANDN U16124 ( .A(x[4721]), .B(y[4721]), .Z(n42196) );
  NANDN U16125 ( .A(x[4722]), .B(y[4722]), .Z(n42202) );
  AND U16126 ( .A(n42196), .B(n42202), .Z(n57003) );
  NANDN U16127 ( .A(y[4720]), .B(x[4720]), .Z(n24904) );
  NANDN U16128 ( .A(y[4721]), .B(x[4721]), .Z(n24903) );
  NAND U16129 ( .A(n24904), .B(n24903), .Z(n57002) );
  NANDN U16130 ( .A(x[4719]), .B(y[4719]), .Z(n24906) );
  XNOR U16131 ( .A(y[4720]), .B(x[4720]), .Z(n9698) );
  AND U16132 ( .A(n24906), .B(n9698), .Z(n57001) );
  NANDN U16133 ( .A(y[4718]), .B(x[4718]), .Z(n24908) );
  NANDN U16134 ( .A(y[4719]), .B(x[4719]), .Z(n24905) );
  NAND U16135 ( .A(n24908), .B(n24905), .Z(n57000) );
  NANDN U16136 ( .A(x[4717]), .B(y[4717]), .Z(n42186) );
  NANDN U16137 ( .A(x[4718]), .B(y[4718]), .Z(n24907) );
  AND U16138 ( .A(n42186), .B(n24907), .Z(n56999) );
  XNOR U16139 ( .A(y[4716]), .B(x[4716]), .Z(n42183) );
  NANDN U16140 ( .A(x[4715]), .B(y[4715]), .Z(n42177) );
  AND U16141 ( .A(n42183), .B(n42177), .Z(n56997) );
  ANDN U16142 ( .B(x[4715]), .A(y[4715]), .Z(n42182) );
  NANDN U16143 ( .A(y[4714]), .B(x[4714]), .Z(n9699) );
  NANDN U16144 ( .A(n42182), .B(n9699), .Z(n56996) );
  XNOR U16145 ( .A(y[4714]), .B(x[4714]), .Z(n24911) );
  NANDN U16146 ( .A(x[4713]), .B(y[4713]), .Z(n24912) );
  AND U16147 ( .A(n24911), .B(n24912), .Z(n56995) );
  NANDN U16148 ( .A(y[4712]), .B(x[4712]), .Z(n9700) );
  NANDN U16149 ( .A(y[4713]), .B(x[4713]), .Z(n24910) );
  NAND U16150 ( .A(n9700), .B(n24910), .Z(n56994) );
  XNOR U16151 ( .A(y[4712]), .B(x[4712]), .Z(n42170) );
  NANDN U16152 ( .A(x[4711]), .B(y[4711]), .Z(n24914) );
  AND U16153 ( .A(n42170), .B(n24914), .Z(n56993) );
  ANDN U16154 ( .B(x[4711]), .A(y[4711]), .Z(n42172) );
  NANDN U16155 ( .A(y[4710]), .B(x[4710]), .Z(n9701) );
  NANDN U16156 ( .A(n42172), .B(n9701), .Z(n56991) );
  NANDN U16157 ( .A(y[4706]), .B(x[4706]), .Z(n24918) );
  NANDN U16158 ( .A(y[4707]), .B(x[4707]), .Z(n24915) );
  AND U16159 ( .A(n24918), .B(n24915), .Z(n56986) );
  NANDN U16160 ( .A(x[4705]), .B(y[4705]), .Z(n24920) );
  NANDN U16161 ( .A(x[4706]), .B(y[4706]), .Z(n24917) );
  NAND U16162 ( .A(n24920), .B(n24917), .Z(n56985) );
  NANDN U16163 ( .A(y[4704]), .B(x[4704]), .Z(n9702) );
  NANDN U16164 ( .A(y[4705]), .B(x[4705]), .Z(n24919) );
  AND U16165 ( .A(n9702), .B(n24919), .Z(n56984) );
  XNOR U16166 ( .A(y[4704]), .B(x[4704]), .Z(n42150) );
  NANDN U16167 ( .A(x[4703]), .B(y[4703]), .Z(n24922) );
  NAND U16168 ( .A(n42150), .B(n24922), .Z(n56983) );
  NANDN U16169 ( .A(y[4702]), .B(x[4702]), .Z(n9703) );
  NANDN U16170 ( .A(y[4703]), .B(x[4703]), .Z(n42149) );
  AND U16171 ( .A(n9703), .B(n42149), .Z(n56982) );
  NANDN U16172 ( .A(y[4700]), .B(x[4700]), .Z(n9704) );
  NANDN U16173 ( .A(y[4701]), .B(x[4701]), .Z(n42143) );
  AND U16174 ( .A(n9704), .B(n42143), .Z(n56980) );
  ANDN U16175 ( .B(y[4699]), .A(x[4699]), .Z(n42135) );
  XNOR U16176 ( .A(y[4700]), .B(x[4700]), .Z(n42138) );
  NANDN U16177 ( .A(n42135), .B(n42138), .Z(n56979) );
  NANDN U16178 ( .A(y[4698]), .B(x[4698]), .Z(n9705) );
  NANDN U16179 ( .A(y[4699]), .B(x[4699]), .Z(n42137) );
  AND U16180 ( .A(n9705), .B(n42137), .Z(n56978) );
  XNOR U16181 ( .A(y[4698]), .B(x[4698]), .Z(n24927) );
  NANDN U16182 ( .A(x[4697]), .B(y[4697]), .Z(n24928) );
  NAND U16183 ( .A(n24927), .B(n24928), .Z(n56977) );
  NANDN U16184 ( .A(y[4696]), .B(x[4696]), .Z(n9706) );
  NANDN U16185 ( .A(y[4697]), .B(x[4697]), .Z(n24926) );
  AND U16186 ( .A(n9706), .B(n24926), .Z(n56976) );
  NANDN U16187 ( .A(y[4694]), .B(x[4694]), .Z(n9707) );
  NANDN U16188 ( .A(y[4695]), .B(x[4695]), .Z(n24929) );
  AND U16189 ( .A(n9707), .B(n24929), .Z(n56972) );
  ANDN U16190 ( .B(y[4693]), .A(x[4693]), .Z(n42120) );
  XNOR U16191 ( .A(y[4694]), .B(x[4694]), .Z(n24932) );
  NANDN U16192 ( .A(n42120), .B(n24932), .Z(n56970) );
  NANDN U16193 ( .A(y[4692]), .B(x[4692]), .Z(n9708) );
  NANDN U16194 ( .A(y[4693]), .B(x[4693]), .Z(n24931) );
  AND U16195 ( .A(n9708), .B(n24931), .Z(n56969) );
  ANDN U16196 ( .B(y[4691]), .A(x[4691]), .Z(n42114) );
  XNOR U16197 ( .A(x[4692]), .B(y[4692]), .Z(n24934) );
  NANDN U16198 ( .A(y[4690]), .B(x[4690]), .Z(n9709) );
  NANDN U16199 ( .A(y[4691]), .B(x[4691]), .Z(n24933) );
  NAND U16200 ( .A(n9709), .B(n24933), .Z(n56966) );
  XNOR U16201 ( .A(x[4690]), .B(y[4690]), .Z(n42112) );
  NANDN U16202 ( .A(x[4689]), .B(y[4689]), .Z(n56965) );
  NANDN U16203 ( .A(y[4688]), .B(x[4688]), .Z(n9710) );
  ANDN U16204 ( .B(x[4689]), .A(y[4689]), .Z(n42111) );
  ANDN U16205 ( .B(n9710), .A(n42111), .Z(n56963) );
  XNOR U16206 ( .A(x[4688]), .B(y[4688]), .Z(n24936) );
  ANDN U16207 ( .B(y[4687]), .A(x[4687]), .Z(n42102) );
  ANDN U16208 ( .B(n24936), .A(n42102), .Z(n16608) );
  XNOR U16209 ( .A(y[4686]), .B(x[4686]), .Z(n24938) );
  NANDN U16210 ( .A(x[4685]), .B(y[4685]), .Z(n24939) );
  AND U16211 ( .A(n24938), .B(n24939), .Z(n56961) );
  NANDN U16212 ( .A(y[4684]), .B(x[4684]), .Z(n9711) );
  NANDN U16213 ( .A(y[4685]), .B(x[4685]), .Z(n24937) );
  NAND U16214 ( .A(n9711), .B(n24937), .Z(n56960) );
  XNOR U16215 ( .A(y[4684]), .B(x[4684]), .Z(n42095) );
  NANDN U16216 ( .A(x[4683]), .B(y[4683]), .Z(n24941) );
  AND U16217 ( .A(n42095), .B(n24941), .Z(n56959) );
  ANDN U16218 ( .B(x[4683]), .A(y[4683]), .Z(n42097) );
  NANDN U16219 ( .A(y[4682]), .B(x[4682]), .Z(n9712) );
  NANDN U16220 ( .A(n42097), .B(n9712), .Z(n56958) );
  NANDN U16221 ( .A(y[4680]), .B(x[4680]), .Z(n9713) );
  NANDN U16222 ( .A(y[4681]), .B(x[4681]), .Z(n42090) );
  AND U16223 ( .A(n9713), .B(n42090), .Z(n56956) );
  XNOR U16224 ( .A(x[4680]), .B(y[4680]), .Z(n24943) );
  NANDN U16225 ( .A(y[4678]), .B(x[4678]), .Z(n9714) );
  NANDN U16226 ( .A(y[4679]), .B(x[4679]), .Z(n24942) );
  NAND U16227 ( .A(n9714), .B(n24942), .Z(n56952) );
  XNOR U16228 ( .A(y[4678]), .B(x[4678]), .Z(n42079) );
  NANDN U16229 ( .A(x[4677]), .B(y[4677]), .Z(n24945) );
  AND U16230 ( .A(n42079), .B(n24945), .Z(n56951) );
  XNOR U16231 ( .A(x[4676]), .B(y[4676]), .Z(n42073) );
  NANDN U16232 ( .A(x[4675]), .B(y[4675]), .Z(n51579) );
  AND U16233 ( .A(n42073), .B(n51579), .Z(n16591) );
  XNOR U16234 ( .A(y[4674]), .B(x[4674]), .Z(n42067) );
  NANDN U16235 ( .A(x[4673]), .B(y[4673]), .Z(n24947) );
  AND U16236 ( .A(n42067), .B(n24947), .Z(n56948) );
  NANDN U16237 ( .A(y[4672]), .B(x[4672]), .Z(n9715) );
  NANDN U16238 ( .A(y[4673]), .B(x[4673]), .Z(n42066) );
  NAND U16239 ( .A(n9715), .B(n42066), .Z(n56947) );
  XNOR U16240 ( .A(y[4672]), .B(x[4672]), .Z(n42061) );
  NANDN U16241 ( .A(x[4671]), .B(y[4671]), .Z(n24949) );
  AND U16242 ( .A(n42061), .B(n24949), .Z(n56946) );
  NANDN U16243 ( .A(y[4670]), .B(x[4670]), .Z(n9716) );
  NANDN U16244 ( .A(y[4671]), .B(x[4671]), .Z(n42060) );
  NAND U16245 ( .A(n9716), .B(n42060), .Z(n56945) );
  XNOR U16246 ( .A(y[4670]), .B(x[4670]), .Z(n42055) );
  NANDN U16247 ( .A(x[4669]), .B(y[4669]), .Z(n24951) );
  AND U16248 ( .A(n42055), .B(n24951), .Z(n56944) );
  XNOR U16249 ( .A(y[4668]), .B(x[4668]), .Z(n42049) );
  NANDN U16250 ( .A(x[4667]), .B(y[4667]), .Z(n42044) );
  AND U16251 ( .A(n42049), .B(n42044), .Z(n56942) );
  NANDN U16252 ( .A(y[4666]), .B(x[4666]), .Z(n24953) );
  NANDN U16253 ( .A(y[4667]), .B(x[4667]), .Z(n42048) );
  NAND U16254 ( .A(n24953), .B(n42048), .Z(n56941) );
  NANDN U16255 ( .A(x[4666]), .B(y[4666]), .Z(n42045) );
  ANDN U16256 ( .B(y[4665]), .A(x[4665]), .Z(n42039) );
  ANDN U16257 ( .B(n42045), .A(n42039), .Z(n56940) );
  NANDN U16258 ( .A(y[4664]), .B(x[4664]), .Z(n24955) );
  NANDN U16259 ( .A(y[4665]), .B(x[4665]), .Z(n24954) );
  NAND U16260 ( .A(n24955), .B(n24954), .Z(n56939) );
  ANDN U16261 ( .B(y[4663]), .A(x[4663]), .Z(n42034) );
  ANDN U16262 ( .B(y[4664]), .A(x[4664]), .Z(n42040) );
  NOR U16263 ( .A(n42034), .B(n42040), .Z(n56938) );
  XNOR U16264 ( .A(x[4662]), .B(y[4662]), .Z(n24958) );
  NANDN U16265 ( .A(y[4660]), .B(x[4660]), .Z(n9717) );
  NANDN U16266 ( .A(y[4661]), .B(x[4661]), .Z(n24957) );
  NAND U16267 ( .A(n9717), .B(n24957), .Z(n56934) );
  XNOR U16268 ( .A(y[4660]), .B(x[4660]), .Z(n24960) );
  NANDN U16269 ( .A(x[4659]), .B(y[4659]), .Z(n42022) );
  AND U16270 ( .A(n24960), .B(n42022), .Z(n56933) );
  NANDN U16271 ( .A(y[4658]), .B(x[4658]), .Z(n9718) );
  NANDN U16272 ( .A(y[4659]), .B(x[4659]), .Z(n24959) );
  NAND U16273 ( .A(n9718), .B(n24959), .Z(n56932) );
  XNOR U16274 ( .A(y[4658]), .B(x[4658]), .Z(n42020) );
  NANDN U16275 ( .A(x[4657]), .B(y[4657]), .Z(n42014) );
  AND U16276 ( .A(n42020), .B(n42014), .Z(n56931) );
  XNOR U16277 ( .A(y[4656]), .B(x[4656]), .Z(n42012) );
  NANDN U16278 ( .A(x[4655]), .B(y[4655]), .Z(n42006) );
  AND U16279 ( .A(n42012), .B(n42006), .Z(n56929) );
  ANDN U16280 ( .B(x[4655]), .A(y[4655]), .Z(n42011) );
  NANDN U16281 ( .A(y[4654]), .B(x[4654]), .Z(n9719) );
  NANDN U16282 ( .A(n42011), .B(n9719), .Z(n56928) );
  XNOR U16283 ( .A(y[4654]), .B(x[4654]), .Z(n42004) );
  NANDN U16284 ( .A(x[4653]), .B(y[4653]), .Z(n41999) );
  AND U16285 ( .A(n42004), .B(n41999), .Z(n56927) );
  ANDN U16286 ( .B(x[4653]), .A(y[4653]), .Z(n42003) );
  NANDN U16287 ( .A(y[4652]), .B(x[4652]), .Z(n9720) );
  NANDN U16288 ( .A(n42003), .B(n9720), .Z(n56926) );
  XNOR U16289 ( .A(x[4652]), .B(y[4652]), .Z(n24962) );
  NANDN U16290 ( .A(x[4651]), .B(y[4651]), .Z(n56924) );
  AND U16291 ( .A(n24962), .B(n56924), .Z(n16561) );
  ANDN U16292 ( .B(x[4649]), .A(y[4649]), .Z(n56920) );
  NANDN U16293 ( .A(y[4648]), .B(x[4648]), .Z(n9721) );
  NANDN U16294 ( .A(n56920), .B(n9721), .Z(n16556) );
  XNOR U16295 ( .A(x[4648]), .B(y[4648]), .Z(n24965) );
  NANDN U16296 ( .A(x[4647]), .B(y[4647]), .Z(n56918) );
  AND U16297 ( .A(n24965), .B(n56918), .Z(n16554) );
  ANDN U16298 ( .B(x[4647]), .A(y[4647]), .Z(n24964) );
  XNOR U16299 ( .A(y[4646]), .B(x[4646]), .Z(n24967) );
  NANDN U16300 ( .A(x[4645]), .B(y[4645]), .Z(n51584) );
  NANDN U16301 ( .A(y[4644]), .B(x[4644]), .Z(n9722) );
  NANDN U16302 ( .A(y[4645]), .B(x[4645]), .Z(n24966) );
  AND U16303 ( .A(n9722), .B(n24966), .Z(n56916) );
  XNOR U16304 ( .A(x[4644]), .B(y[4644]), .Z(n41979) );
  ANDN U16305 ( .B(y[4643]), .A(x[4643]), .Z(n56914) );
  ANDN U16306 ( .B(n41979), .A(n56914), .Z(n16547) );
  XNOR U16307 ( .A(y[4642]), .B(x[4642]), .Z(n41973) );
  NANDN U16308 ( .A(x[4641]), .B(y[4641]), .Z(n24969) );
  AND U16309 ( .A(n41973), .B(n24969), .Z(n56913) );
  NANDN U16310 ( .A(y[4640]), .B(x[4640]), .Z(n9723) );
  NANDN U16311 ( .A(y[4641]), .B(x[4641]), .Z(n41972) );
  AND U16312 ( .A(n9723), .B(n41972), .Z(n56912) );
  NANDN U16313 ( .A(x[4638]), .B(y[4638]), .Z(n56908) );
  NANDN U16314 ( .A(y[4637]), .B(x[4637]), .Z(n41963) );
  NANDN U16315 ( .A(y[4636]), .B(x[4636]), .Z(n56905) );
  NANDN U16316 ( .A(x[4635]), .B(y[4635]), .Z(n41955) );
  NANDN U16317 ( .A(x[4636]), .B(y[4636]), .Z(n24972) );
  NAND U16318 ( .A(n41955), .B(n24972), .Z(n56904) );
  NANDN U16319 ( .A(y[4634]), .B(x[4634]), .Z(n9724) );
  NANDN U16320 ( .A(y[4635]), .B(x[4635]), .Z(n24973) );
  AND U16321 ( .A(n9724), .B(n24973), .Z(n56903) );
  XNOR U16322 ( .A(y[4634]), .B(x[4634]), .Z(n41951) );
  NANDN U16323 ( .A(x[4633]), .B(y[4633]), .Z(n41946) );
  NAND U16324 ( .A(n41951), .B(n41946), .Z(n56902) );
  NANDN U16325 ( .A(y[4632]), .B(x[4632]), .Z(n9725) );
  NANDN U16326 ( .A(y[4633]), .B(x[4633]), .Z(n41950) );
  AND U16327 ( .A(n9725), .B(n41950), .Z(n56901) );
  XNOR U16328 ( .A(y[4632]), .B(x[4632]), .Z(n41944) );
  NANDN U16329 ( .A(x[4631]), .B(y[4631]), .Z(n41938) );
  NAND U16330 ( .A(n41944), .B(n41938), .Z(n56900) );
  ANDN U16331 ( .B(x[4629]), .A(y[4629]), .Z(n41935) );
  NANDN U16332 ( .A(y[4628]), .B(x[4628]), .Z(n9726) );
  NANDN U16333 ( .A(n41935), .B(n9726), .Z(n51589) );
  XNOR U16334 ( .A(y[4628]), .B(x[4628]), .Z(n41928) );
  NANDN U16335 ( .A(x[4627]), .B(y[4627]), .Z(n41922) );
  AND U16336 ( .A(n41928), .B(n41922), .Z(n56898) );
  NANDN U16337 ( .A(y[4622]), .B(x[4622]), .Z(n9727) );
  NANDN U16338 ( .A(y[4623]), .B(x[4623]), .Z(n24975) );
  NAND U16339 ( .A(n9727), .B(n24975), .Z(n51591) );
  XNOR U16340 ( .A(y[4622]), .B(x[4622]), .Z(n41905) );
  NANDN U16341 ( .A(x[4621]), .B(y[4621]), .Z(n41901) );
  AND U16342 ( .A(n41905), .B(n41901), .Z(n56892) );
  XNOR U16343 ( .A(x[4620]), .B(y[4620]), .Z(n41899) );
  NANDN U16344 ( .A(x[4619]), .B(y[4619]), .Z(n56889) );
  AND U16345 ( .A(n41899), .B(n56889), .Z(n16514) );
  XNOR U16346 ( .A(x[4618]), .B(y[4618]), .Z(n24977) );
  NANDN U16347 ( .A(y[4616]), .B(x[4616]), .Z(n9728) );
  NANDN U16348 ( .A(y[4617]), .B(x[4617]), .Z(n24976) );
  NAND U16349 ( .A(n9728), .B(n24976), .Z(n56886) );
  XNOR U16350 ( .A(y[4616]), .B(x[4616]), .Z(n41888) );
  NANDN U16351 ( .A(x[4615]), .B(y[4615]), .Z(n24979) );
  AND U16352 ( .A(n41888), .B(n24979), .Z(n56885) );
  NANDN U16353 ( .A(x[4614]), .B(y[4614]), .Z(n24980) );
  ANDN U16354 ( .B(y[4613]), .A(x[4613]), .Z(n41880) );
  ANDN U16355 ( .B(n24980), .A(n41880), .Z(n56882) );
  XNOR U16356 ( .A(x[4612]), .B(y[4612]), .Z(n24982) );
  NANDN U16357 ( .A(y[4610]), .B(x[4610]), .Z(n9729) );
  NANDN U16358 ( .A(y[4611]), .B(x[4611]), .Z(n24981) );
  NAND U16359 ( .A(n9729), .B(n24981), .Z(n56880) );
  XNOR U16360 ( .A(y[4610]), .B(x[4610]), .Z(n24985) );
  NANDN U16361 ( .A(x[4609]), .B(y[4609]), .Z(n24986) );
  AND U16362 ( .A(n24985), .B(n24986), .Z(n56879) );
  NANDN U16363 ( .A(y[4608]), .B(x[4608]), .Z(n9730) );
  NANDN U16364 ( .A(y[4609]), .B(x[4609]), .Z(n24984) );
  NAND U16365 ( .A(n9730), .B(n24984), .Z(n56878) );
  XNOR U16366 ( .A(x[4608]), .B(y[4608]), .Z(n41867) );
  NANDN U16367 ( .A(x[4607]), .B(y[4607]), .Z(n56877) );
  AND U16368 ( .A(n41867), .B(n56877), .Z(n16497) );
  NANDN U16369 ( .A(y[4604]), .B(x[4604]), .Z(n9731) );
  NANDN U16370 ( .A(y[4605]), .B(x[4605]), .Z(n41860) );
  NAND U16371 ( .A(n9731), .B(n41860), .Z(n51597) );
  XNOR U16372 ( .A(y[4604]), .B(x[4604]), .Z(n41855) );
  NANDN U16373 ( .A(x[4603]), .B(y[4603]), .Z(n24990) );
  AND U16374 ( .A(n41855), .B(n24990), .Z(n56873) );
  NANDN U16375 ( .A(y[4598]), .B(x[4598]), .Z(n9732) );
  NANDN U16376 ( .A(y[4599]), .B(x[4599]), .Z(n24992) );
  NAND U16377 ( .A(n9732), .B(n24992), .Z(n51599) );
  XNOR U16378 ( .A(y[4598]), .B(x[4598]), .Z(n24995) );
  NANDN U16379 ( .A(x[4597]), .B(y[4597]), .Z(n24996) );
  AND U16380 ( .A(n24995), .B(n24996), .Z(n56867) );
  XNOR U16381 ( .A(y[4594]), .B(x[4594]), .Z(n41827) );
  NANDN U16382 ( .A(x[4593]), .B(y[4593]), .Z(n25002) );
  AND U16383 ( .A(n41827), .B(n25002), .Z(n56864) );
  NANDN U16384 ( .A(y[4592]), .B(x[4592]), .Z(n9733) );
  NANDN U16385 ( .A(y[4593]), .B(x[4593]), .Z(n41826) );
  NAND U16386 ( .A(n9733), .B(n41826), .Z(n56863) );
  XNOR U16387 ( .A(y[4592]), .B(x[4592]), .Z(n41821) );
  ANDN U16388 ( .B(y[4591]), .A(x[4591]), .Z(n41817) );
  ANDN U16389 ( .B(n41821), .A(n41817), .Z(n56862) );
  NANDN U16390 ( .A(y[4590]), .B(x[4590]), .Z(n25004) );
  NANDN U16391 ( .A(y[4591]), .B(x[4591]), .Z(n41820) );
  NAND U16392 ( .A(n25004), .B(n41820), .Z(n56861) );
  NANDN U16393 ( .A(x[4590]), .B(y[4590]), .Z(n41819) );
  ANDN U16394 ( .B(y[4589]), .A(x[4589]), .Z(n41812) );
  ANDN U16395 ( .B(n41819), .A(n41812), .Z(n56860) );
  NANDN U16396 ( .A(y[4588]), .B(x[4588]), .Z(n9734) );
  NANDN U16397 ( .A(y[4589]), .B(x[4589]), .Z(n25005) );
  NAND U16398 ( .A(n9734), .B(n25005), .Z(n56858) );
  ANDN U16399 ( .B(y[4587]), .A(x[4587]), .Z(n56856) );
  XNOR U16400 ( .A(x[4588]), .B(y[4588]), .Z(n25007) );
  NANDN U16401 ( .A(y[4586]), .B(x[4586]), .Z(n9735) );
  NANDN U16402 ( .A(y[4587]), .B(x[4587]), .Z(n25006) );
  NAND U16403 ( .A(n9735), .B(n25006), .Z(n56855) );
  NANDN U16404 ( .A(x[4585]), .B(y[4585]), .Z(n56854) );
  NANDN U16405 ( .A(y[4584]), .B(x[4584]), .Z(n9736) );
  NANDN U16406 ( .A(y[4585]), .B(x[4585]), .Z(n25008) );
  AND U16407 ( .A(n9736), .B(n25008), .Z(n56852) );
  XNOR U16408 ( .A(y[4584]), .B(x[4584]), .Z(n41800) );
  NANDN U16409 ( .A(x[4583]), .B(y[4583]), .Z(n41794) );
  NAND U16410 ( .A(n41800), .B(n41794), .Z(n56851) );
  NANDN U16411 ( .A(y[4582]), .B(x[4582]), .Z(n9737) );
  ANDN U16412 ( .B(x[4583]), .A(y[4583]), .Z(n41799) );
  ANDN U16413 ( .B(n9737), .A(n41799), .Z(n56850) );
  XNOR U16414 ( .A(y[4582]), .B(x[4582]), .Z(n41792) );
  NANDN U16415 ( .A(x[4581]), .B(y[4581]), .Z(n41786) );
  NAND U16416 ( .A(n41792), .B(n41786), .Z(n56849) );
  NANDN U16417 ( .A(y[4580]), .B(x[4580]), .Z(n9738) );
  ANDN U16418 ( .B(x[4581]), .A(y[4581]), .Z(n41791) );
  ANDN U16419 ( .B(n9738), .A(n41791), .Z(n56848) );
  NANDN U16420 ( .A(y[4578]), .B(x[4578]), .Z(n9739) );
  ANDN U16421 ( .B(x[4579]), .A(y[4579]), .Z(n41783) );
  ANDN U16422 ( .B(n9739), .A(n41783), .Z(n56846) );
  XNOR U16423 ( .A(y[4578]), .B(x[4578]), .Z(n41775) );
  NANDN U16424 ( .A(x[4577]), .B(y[4577]), .Z(n41770) );
  NAND U16425 ( .A(n41775), .B(n41770), .Z(n56845) );
  NANDN U16426 ( .A(y[4576]), .B(x[4576]), .Z(n9740) );
  NANDN U16427 ( .A(y[4577]), .B(x[4577]), .Z(n41774) );
  AND U16428 ( .A(n9740), .B(n41774), .Z(n56844) );
  XNOR U16429 ( .A(y[4576]), .B(x[4576]), .Z(n41768) );
  NANDN U16430 ( .A(x[4575]), .B(y[4575]), .Z(n41763) );
  NAND U16431 ( .A(n41768), .B(n41763), .Z(n56843) );
  NANDN U16432 ( .A(y[4574]), .B(x[4574]), .Z(n9741) );
  ANDN U16433 ( .B(x[4575]), .A(y[4575]), .Z(n41767) );
  ANDN U16434 ( .B(n9741), .A(n41767), .Z(n56842) );
  NANDN U16435 ( .A(x[4573]), .B(y[4573]), .Z(n56838) );
  XNOR U16436 ( .A(x[4574]), .B(y[4574]), .Z(n41760) );
  NAND U16437 ( .A(n56838), .B(n41760), .Z(n16454) );
  NANDN U16438 ( .A(x[4571]), .B(y[4571]), .Z(n25011) );
  NANDN U16439 ( .A(x[4572]), .B(y[4572]), .Z(n25010) );
  AND U16440 ( .A(n25011), .B(n25010), .Z(n56836) );
  XNOR U16441 ( .A(x[4570]), .B(y[4570]), .Z(n41748) );
  NANDN U16442 ( .A(y[4568]), .B(x[4568]), .Z(n9742) );
  NANDN U16443 ( .A(y[4569]), .B(x[4569]), .Z(n41749) );
  NAND U16444 ( .A(n9742), .B(n41749), .Z(n56832) );
  XNOR U16445 ( .A(x[4568]), .B(y[4568]), .Z(n25013) );
  NANDN U16446 ( .A(y[4566]), .B(x[4566]), .Z(n9743) );
  NANDN U16447 ( .A(y[4567]), .B(x[4567]), .Z(n25012) );
  NAND U16448 ( .A(n9743), .B(n25012), .Z(n56829) );
  XNOR U16449 ( .A(x[4566]), .B(y[4566]), .Z(n25015) );
  NANDN U16450 ( .A(x[4565]), .B(y[4565]), .Z(n56828) );
  NANDN U16451 ( .A(y[4564]), .B(x[4564]), .Z(n9744) );
  NANDN U16452 ( .A(y[4565]), .B(x[4565]), .Z(n25014) );
  AND U16453 ( .A(n9744), .B(n25014), .Z(n56826) );
  XNOR U16454 ( .A(x[4564]), .B(y[4564]), .Z(n25017) );
  ANDN U16455 ( .B(y[4563]), .A(x[4563]), .Z(n51601) );
  ANDN U16456 ( .B(n25017), .A(n51601), .Z(n16439) );
  XNOR U16457 ( .A(y[4562]), .B(x[4562]), .Z(n25019) );
  ANDN U16458 ( .B(y[4561]), .A(x[4561]), .Z(n41727) );
  ANDN U16459 ( .B(n25019), .A(n41727), .Z(n56824) );
  NANDN U16460 ( .A(y[4560]), .B(x[4560]), .Z(n9745) );
  NANDN U16461 ( .A(y[4561]), .B(x[4561]), .Z(n25018) );
  NAND U16462 ( .A(n9745), .B(n25018), .Z(n56823) );
  XNOR U16463 ( .A(y[4560]), .B(x[4560]), .Z(n41723) );
  NANDN U16464 ( .A(x[4559]), .B(y[4559]), .Z(n25020) );
  AND U16465 ( .A(n41723), .B(n25020), .Z(n56822) );
  NANDN U16466 ( .A(y[4558]), .B(x[4558]), .Z(n9746) );
  NANDN U16467 ( .A(y[4559]), .B(x[4559]), .Z(n41722) );
  NAND U16468 ( .A(n9746), .B(n41722), .Z(n56820) );
  XNOR U16469 ( .A(y[4558]), .B(x[4558]), .Z(n25023) );
  NANDN U16470 ( .A(x[4557]), .B(y[4557]), .Z(n25024) );
  AND U16471 ( .A(n25023), .B(n25024), .Z(n56819) );
  NANDN U16472 ( .A(x[4555]), .B(y[4555]), .Z(n41709) );
  XOR U16473 ( .A(y[4556]), .B(x[4556]), .Z(n41714) );
  ANDN U16474 ( .B(n41709), .A(n41714), .Z(n56817) );
  ANDN U16475 ( .B(x[4555]), .A(y[4555]), .Z(n41712) );
  NANDN U16476 ( .A(y[4554]), .B(x[4554]), .Z(n9747) );
  NANDN U16477 ( .A(n41712), .B(n9747), .Z(n56816) );
  XNOR U16478 ( .A(y[4554]), .B(x[4554]), .Z(n41705) );
  NANDN U16479 ( .A(x[4553]), .B(y[4553]), .Z(n25026) );
  AND U16480 ( .A(n41705), .B(n25026), .Z(n56815) );
  ANDN U16481 ( .B(x[4553]), .A(y[4553]), .Z(n41707) );
  NANDN U16482 ( .A(y[4552]), .B(x[4552]), .Z(n9748) );
  NANDN U16483 ( .A(n41707), .B(n9748), .Z(n56814) );
  XNOR U16484 ( .A(x[4552]), .B(y[4552]), .Z(n41699) );
  XNOR U16485 ( .A(x[4550]), .B(y[4550]), .Z(n25028) );
  NANDN U16486 ( .A(x[4549]), .B(y[4549]), .Z(n56811) );
  AND U16487 ( .A(n25028), .B(n56811), .Z(n16420) );
  XNOR U16488 ( .A(x[4548]), .B(y[4548]), .Z(n25030) );
  NANDN U16489 ( .A(y[4546]), .B(x[4546]), .Z(n9749) );
  NANDN U16490 ( .A(y[4547]), .B(x[4547]), .Z(n25029) );
  NAND U16491 ( .A(n9749), .B(n25029), .Z(n56807) );
  XNOR U16492 ( .A(y[4546]), .B(x[4546]), .Z(n41685) );
  NANDN U16493 ( .A(x[4545]), .B(y[4545]), .Z(n25032) );
  AND U16494 ( .A(n41685), .B(n25032), .Z(n56806) );
  NANDN U16495 ( .A(y[4544]), .B(x[4544]), .Z(n9750) );
  NANDN U16496 ( .A(y[4545]), .B(x[4545]), .Z(n41684) );
  NAND U16497 ( .A(n9750), .B(n41684), .Z(n56804) );
  XNOR U16498 ( .A(y[4544]), .B(x[4544]), .Z(n41679) );
  NANDN U16499 ( .A(x[4543]), .B(y[4543]), .Z(n25034) );
  AND U16500 ( .A(n41679), .B(n25034), .Z(n56802) );
  NANDN U16501 ( .A(x[4541]), .B(y[4541]), .Z(n25036) );
  NANDN U16502 ( .A(x[4542]), .B(y[4542]), .Z(n25035) );
  AND U16503 ( .A(n25036), .B(n25035), .Z(n56798) );
  NANDN U16504 ( .A(y[4540]), .B(x[4540]), .Z(n9751) );
  NANDN U16505 ( .A(y[4541]), .B(x[4541]), .Z(n41673) );
  NAND U16506 ( .A(n9751), .B(n41673), .Z(n56796) );
  XNOR U16507 ( .A(y[4540]), .B(x[4540]), .Z(n41667) );
  NANDN U16508 ( .A(x[4539]), .B(y[4539]), .Z(n25038) );
  AND U16509 ( .A(n41667), .B(n25038), .Z(n56794) );
  NANDN U16510 ( .A(y[4538]), .B(x[4538]), .Z(n9752) );
  NANDN U16511 ( .A(y[4539]), .B(x[4539]), .Z(n41666) );
  NAND U16512 ( .A(n9752), .B(n41666), .Z(n56791) );
  XNOR U16513 ( .A(x[4538]), .B(y[4538]), .Z(n25040) );
  NANDN U16514 ( .A(x[4537]), .B(y[4537]), .Z(n56788) );
  AND U16515 ( .A(n25040), .B(n56788), .Z(n16405) );
  XNOR U16516 ( .A(y[4536]), .B(x[4536]), .Z(n25042) );
  NANDN U16517 ( .A(x[4535]), .B(y[4535]), .Z(n41654) );
  AND U16518 ( .A(n25042), .B(n41654), .Z(n56784) );
  NANDN U16519 ( .A(y[4534]), .B(x[4534]), .Z(n25043) );
  NANDN U16520 ( .A(y[4535]), .B(x[4535]), .Z(n25041) );
  NAND U16521 ( .A(n25043), .B(n25041), .Z(n56782) );
  NANDN U16522 ( .A(x[4533]), .B(y[4533]), .Z(n41648) );
  NANDN U16523 ( .A(x[4534]), .B(y[4534]), .Z(n41655) );
  AND U16524 ( .A(n41648), .B(n41655), .Z(n56780) );
  NANDN U16525 ( .A(y[4532]), .B(x[4532]), .Z(n9753) );
  NANDN U16526 ( .A(y[4533]), .B(x[4533]), .Z(n25044) );
  NAND U16527 ( .A(n9753), .B(n25044), .Z(n56777) );
  NANDN U16528 ( .A(y[4530]), .B(x[4530]), .Z(n9754) );
  ANDN U16529 ( .B(x[4531]), .A(y[4531]), .Z(n41645) );
  ANDN U16530 ( .B(n9754), .A(n41645), .Z(n56772) );
  XNOR U16531 ( .A(x[4530]), .B(y[4530]), .Z(n41639) );
  NANDN U16532 ( .A(y[4528]), .B(x[4528]), .Z(n9755) );
  NANDN U16533 ( .A(y[4529]), .B(x[4529]), .Z(n41640) );
  AND U16534 ( .A(n9755), .B(n41640), .Z(n56766) );
  XNOR U16535 ( .A(y[4528]), .B(x[4528]), .Z(n41633) );
  NANDN U16536 ( .A(x[4527]), .B(y[4527]), .Z(n25047) );
  NAND U16537 ( .A(n41633), .B(n25047), .Z(n56764) );
  NANDN U16538 ( .A(y[4526]), .B(x[4526]), .Z(n9756) );
  NANDN U16539 ( .A(y[4527]), .B(x[4527]), .Z(n41634) );
  AND U16540 ( .A(n9756), .B(n41634), .Z(n56763) );
  ANDN U16541 ( .B(y[4525]), .A(x[4525]), .Z(n41623) );
  XNOR U16542 ( .A(y[4526]), .B(x[4526]), .Z(n41627) );
  NANDN U16543 ( .A(n41623), .B(n41627), .Z(n56762) );
  NANDN U16544 ( .A(y[4524]), .B(x[4524]), .Z(n41619) );
  NANDN U16545 ( .A(y[4525]), .B(x[4525]), .Z(n41628) );
  AND U16546 ( .A(n41619), .B(n41628), .Z(n56761) );
  NANDN U16547 ( .A(x[4523]), .B(y[4523]), .Z(n25049) );
  ANDN U16548 ( .B(y[4524]), .A(x[4524]), .Z(n41625) );
  ANDN U16549 ( .B(n25049), .A(n41625), .Z(n56760) );
  NANDN U16550 ( .A(y[4522]), .B(x[4522]), .Z(n41612) );
  NANDN U16551 ( .A(y[4523]), .B(x[4523]), .Z(n41621) );
  NAND U16552 ( .A(n41612), .B(n41621), .Z(n56759) );
  NANDN U16553 ( .A(x[4521]), .B(y[4521]), .Z(n25051) );
  NANDN U16554 ( .A(x[4522]), .B(y[4522]), .Z(n25050) );
  AND U16555 ( .A(n25051), .B(n25050), .Z(n51605) );
  XNOR U16556 ( .A(y[4520]), .B(x[4520]), .Z(n41607) );
  ANDN U16557 ( .B(y[4519]), .A(x[4519]), .Z(n41604) );
  ANDN U16558 ( .B(n41607), .A(n41604), .Z(n56758) );
  XNOR U16559 ( .A(x[4518]), .B(y[4518]), .Z(n25054) );
  NANDN U16560 ( .A(y[4516]), .B(x[4516]), .Z(n9757) );
  NANDN U16561 ( .A(y[4517]), .B(x[4517]), .Z(n25053) );
  NAND U16562 ( .A(n9757), .B(n25053), .Z(n56754) );
  XNOR U16563 ( .A(y[4516]), .B(x[4516]), .Z(n25057) );
  NANDN U16564 ( .A(x[4515]), .B(y[4515]), .Z(n25058) );
  AND U16565 ( .A(n25057), .B(n25058), .Z(n51607) );
  NANDN U16566 ( .A(y[4512]), .B(x[4512]), .Z(n9758) );
  NANDN U16567 ( .A(y[4513]), .B(x[4513]), .Z(n41591) );
  NAND U16568 ( .A(n9758), .B(n41591), .Z(n56750) );
  NANDN U16569 ( .A(y[4510]), .B(x[4510]), .Z(n9759) );
  NANDN U16570 ( .A(y[4511]), .B(x[4511]), .Z(n41585) );
  AND U16571 ( .A(n9759), .B(n41585), .Z(n56749) );
  XNOR U16572 ( .A(y[4510]), .B(x[4510]), .Z(n25063) );
  NANDN U16573 ( .A(x[4509]), .B(y[4509]), .Z(n41576) );
  NAND U16574 ( .A(n25063), .B(n41576), .Z(n56748) );
  NANDN U16575 ( .A(y[4508]), .B(x[4508]), .Z(n25064) );
  NANDN U16576 ( .A(y[4509]), .B(x[4509]), .Z(n25062) );
  AND U16577 ( .A(n25064), .B(n25062), .Z(n56747) );
  NANDN U16578 ( .A(x[4507]), .B(y[4507]), .Z(n41570) );
  NANDN U16579 ( .A(x[4508]), .B(y[4508]), .Z(n41577) );
  NAND U16580 ( .A(n41570), .B(n41577), .Z(n56746) );
  NANDN U16581 ( .A(y[4506]), .B(x[4506]), .Z(n25066) );
  NANDN U16582 ( .A(y[4507]), .B(x[4507]), .Z(n25065) );
  AND U16583 ( .A(n25066), .B(n25065), .Z(n56745) );
  NANDN U16584 ( .A(y[4504]), .B(x[4504]), .Z(n25070) );
  NANDN U16585 ( .A(y[4505]), .B(x[4505]), .Z(n25067) );
  AND U16586 ( .A(n25070), .B(n25067), .Z(n56743) );
  NANDN U16587 ( .A(x[4503]), .B(y[4503]), .Z(n41560) );
  NANDN U16588 ( .A(x[4504]), .B(y[4504]), .Z(n25069) );
  NAND U16589 ( .A(n41560), .B(n25069), .Z(n56742) );
  NANDN U16590 ( .A(y[4502]), .B(x[4502]), .Z(n9760) );
  NANDN U16591 ( .A(y[4503]), .B(x[4503]), .Z(n25071) );
  AND U16592 ( .A(n9760), .B(n25071), .Z(n56741) );
  XNOR U16593 ( .A(y[4502]), .B(x[4502]), .Z(n41557) );
  NANDN U16594 ( .A(x[4501]), .B(y[4501]), .Z(n41551) );
  NAND U16595 ( .A(n41557), .B(n41551), .Z(n56740) );
  NANDN U16596 ( .A(y[4500]), .B(x[4500]), .Z(n9761) );
  ANDN U16597 ( .B(x[4501]), .A(y[4501]), .Z(n41556) );
  ANDN U16598 ( .B(n9761), .A(n41556), .Z(n56739) );
  NANDN U16599 ( .A(y[4498]), .B(x[4498]), .Z(n9762) );
  ANDN U16600 ( .B(x[4499]), .A(y[4499]), .Z(n41548) );
  ANDN U16601 ( .B(n9762), .A(n41548), .Z(n56736) );
  XNOR U16602 ( .A(y[4498]), .B(x[4498]), .Z(n41540) );
  NANDN U16603 ( .A(x[4497]), .B(y[4497]), .Z(n41535) );
  NAND U16604 ( .A(n41540), .B(n41535), .Z(n51610) );
  NANDN U16605 ( .A(y[4496]), .B(x[4496]), .Z(n9763) );
  NANDN U16606 ( .A(y[4497]), .B(x[4497]), .Z(n41539) );
  AND U16607 ( .A(n9763), .B(n41539), .Z(n56735) );
  ANDN U16608 ( .B(x[4490]), .A(y[4490]), .Z(n25081) );
  NANDN U16609 ( .A(x[4489]), .B(y[4489]), .Z(n56728) );
  NANDN U16610 ( .A(y[4488]), .B(x[4488]), .Z(n56727) );
  NANDN U16611 ( .A(y[4489]), .B(x[4489]), .Z(n25082) );
  AND U16612 ( .A(n56727), .B(n25082), .Z(n16343) );
  XNOR U16613 ( .A(x[4486]), .B(y[4486]), .Z(n25086) );
  NANDN U16614 ( .A(x[4485]), .B(y[4485]), .Z(n56723) );
  AND U16615 ( .A(n25086), .B(n56723), .Z(n16338) );
  XNOR U16616 ( .A(y[4484]), .B(x[4484]), .Z(n25088) );
  ANDN U16617 ( .B(y[4483]), .A(x[4483]), .Z(n41504) );
  ANDN U16618 ( .B(n25088), .A(n41504), .Z(n56720) );
  NANDN U16619 ( .A(y[4482]), .B(x[4482]), .Z(n9764) );
  NANDN U16620 ( .A(y[4483]), .B(x[4483]), .Z(n25087) );
  NAND U16621 ( .A(n9764), .B(n25087), .Z(n56719) );
  XNOR U16622 ( .A(y[4482]), .B(x[4482]), .Z(n25090) );
  NANDN U16623 ( .A(x[4481]), .B(y[4481]), .Z(n25091) );
  AND U16624 ( .A(n25090), .B(n25091), .Z(n56718) );
  NANDN U16625 ( .A(y[4480]), .B(x[4480]), .Z(n25093) );
  NANDN U16626 ( .A(y[4481]), .B(x[4481]), .Z(n25089) );
  NAND U16627 ( .A(n25093), .B(n25089), .Z(n56717) );
  NANDN U16628 ( .A(x[4479]), .B(y[4479]), .Z(n41494) );
  NANDN U16629 ( .A(x[4480]), .B(y[4480]), .Z(n25092) );
  AND U16630 ( .A(n41494), .B(n25092), .Z(n56716) );
  NANDN U16631 ( .A(y[4478]), .B(x[4478]), .Z(n9765) );
  NANDN U16632 ( .A(y[4479]), .B(x[4479]), .Z(n25094) );
  NAND U16633 ( .A(n9765), .B(n25094), .Z(n56715) );
  XNOR U16634 ( .A(x[4478]), .B(y[4478]), .Z(n41491) );
  NANDN U16635 ( .A(x[4477]), .B(y[4477]), .Z(n51612) );
  NANDN U16636 ( .A(y[4476]), .B(x[4476]), .Z(n9766) );
  NANDN U16637 ( .A(y[4477]), .B(x[4477]), .Z(n41492) );
  NAND U16638 ( .A(n9766), .B(n41492), .Z(n56714) );
  ANDN U16639 ( .B(y[4473]), .A(x[4473]), .Z(n41475) );
  XNOR U16640 ( .A(y[4474]), .B(x[4474]), .Z(n41479) );
  NANDN U16641 ( .A(n41475), .B(n41479), .Z(n51615) );
  NANDN U16642 ( .A(y[4472]), .B(x[4472]), .Z(n9767) );
  NANDN U16643 ( .A(y[4473]), .B(x[4473]), .Z(n41480) );
  AND U16644 ( .A(n9767), .B(n41480), .Z(n56712) );
  NANDN U16645 ( .A(y[4470]), .B(x[4470]), .Z(n9768) );
  NANDN U16646 ( .A(y[4471]), .B(x[4471]), .Z(n41473) );
  AND U16647 ( .A(n9768), .B(n41473), .Z(n56709) );
  XNOR U16648 ( .A(y[4470]), .B(x[4470]), .Z(n41465) );
  NANDN U16649 ( .A(x[4469]), .B(y[4469]), .Z(n25100) );
  NAND U16650 ( .A(n41465), .B(n25100), .Z(n56707) );
  NANDN U16651 ( .A(y[4466]), .B(x[4466]), .Z(n9769) );
  NANDN U16652 ( .A(y[4467]), .B(x[4467]), .Z(n41458) );
  NAND U16653 ( .A(n9769), .B(n41458), .Z(n56704) );
  XNOR U16654 ( .A(y[4466]), .B(x[4466]), .Z(n25105) );
  ANDN U16655 ( .B(y[4465]), .A(x[4465]), .Z(n41452) );
  ANDN U16656 ( .B(n25105), .A(n41452), .Z(n56703) );
  XNOR U16657 ( .A(y[4464]), .B(x[4464]), .Z(n25107) );
  ANDN U16658 ( .B(y[4463]), .A(x[4463]), .Z(n41446) );
  ANDN U16659 ( .B(n25107), .A(n41446), .Z(n56702) );
  XNOR U16660 ( .A(x[4462]), .B(y[4462]), .Z(n41442) );
  XNOR U16661 ( .A(x[4460]), .B(y[4460]), .Z(n25109) );
  NANDN U16662 ( .A(y[4458]), .B(x[4458]), .Z(n9770) );
  NANDN U16663 ( .A(y[4459]), .B(x[4459]), .Z(n25108) );
  NAND U16664 ( .A(n9770), .B(n25108), .Z(n56695) );
  XNOR U16665 ( .A(y[4458]), .B(x[4458]), .Z(n25112) );
  NANDN U16666 ( .A(x[4457]), .B(y[4457]), .Z(n41429) );
  AND U16667 ( .A(n25112), .B(n41429), .Z(n56694) );
  NANDN U16668 ( .A(y[4454]), .B(x[4454]), .Z(n25115) );
  NANDN U16669 ( .A(y[4455]), .B(x[4455]), .Z(n41425) );
  NAND U16670 ( .A(n25115), .B(n41425), .Z(n56691) );
  NANDN U16671 ( .A(x[4453]), .B(y[4453]), .Z(n41418) );
  NANDN U16672 ( .A(x[4454]), .B(y[4454]), .Z(n25114) );
  AND U16673 ( .A(n41418), .B(n25114), .Z(n51620) );
  XNOR U16674 ( .A(x[4450]), .B(y[4450]), .Z(n25117) );
  NANDN U16675 ( .A(y[4448]), .B(x[4448]), .Z(n9771) );
  NANDN U16676 ( .A(y[4449]), .B(x[4449]), .Z(n25118) );
  NAND U16677 ( .A(n9771), .B(n25118), .Z(n51623) );
  NANDN U16678 ( .A(y[4446]), .B(x[4446]), .Z(n9772) );
  ANDN U16679 ( .B(x[4447]), .A(y[4447]), .Z(n41402) );
  ANDN U16680 ( .B(n9772), .A(n41402), .Z(n56686) );
  XNOR U16681 ( .A(y[4446]), .B(x[4446]), .Z(n25119) );
  NANDN U16682 ( .A(x[4445]), .B(y[4445]), .Z(n41391) );
  NAND U16683 ( .A(n25119), .B(n41391), .Z(n56685) );
  NANDN U16684 ( .A(y[4444]), .B(x[4444]), .Z(n9773) );
  NANDN U16685 ( .A(y[4445]), .B(x[4445]), .Z(n25120) );
  AND U16686 ( .A(n9773), .B(n25120), .Z(n56684) );
  XNOR U16687 ( .A(y[4444]), .B(x[4444]), .Z(n41389) );
  NANDN U16688 ( .A(x[4443]), .B(y[4443]), .Z(n41383) );
  NAND U16689 ( .A(n41389), .B(n41383), .Z(n56683) );
  NANDN U16690 ( .A(y[4442]), .B(x[4442]), .Z(n9774) );
  ANDN U16691 ( .B(x[4443]), .A(y[4443]), .Z(n41388) );
  ANDN U16692 ( .B(n9774), .A(n41388), .Z(n56682) );
  XNOR U16693 ( .A(y[4442]), .B(x[4442]), .Z(n41380) );
  NANDN U16694 ( .A(x[4441]), .B(y[4441]), .Z(n41375) );
  NAND U16695 ( .A(n41380), .B(n41375), .Z(n56681) );
  ANDN U16696 ( .B(x[4439]), .A(y[4439]), .Z(n41372) );
  NANDN U16697 ( .A(y[4438]), .B(x[4438]), .Z(n9775) );
  NANDN U16698 ( .A(n41372), .B(n9775), .Z(n56678) );
  XNOR U16699 ( .A(y[4438]), .B(x[4438]), .Z(n41365) );
  NANDN U16700 ( .A(x[4437]), .B(y[4437]), .Z(n41359) );
  AND U16701 ( .A(n41365), .B(n41359), .Z(n51625) );
  XNOR U16702 ( .A(y[4436]), .B(x[4436]), .Z(n41357) );
  NANDN U16703 ( .A(x[4435]), .B(y[4435]), .Z(n41351) );
  AND U16704 ( .A(n41357), .B(n41351), .Z(n56676) );
  XNOR U16705 ( .A(y[4434]), .B(x[4434]), .Z(n41348) );
  NANDN U16706 ( .A(x[4433]), .B(y[4433]), .Z(n25121) );
  AND U16707 ( .A(n41348), .B(n25121), .Z(n56674) );
  NANDN U16708 ( .A(y[4432]), .B(x[4432]), .Z(n41342) );
  NANDN U16709 ( .A(y[4433]), .B(x[4433]), .Z(n41349) );
  NAND U16710 ( .A(n41342), .B(n41349), .Z(n56673) );
  NANDN U16711 ( .A(x[4431]), .B(y[4431]), .Z(n25123) );
  NANDN U16712 ( .A(x[4432]), .B(y[4432]), .Z(n25122) );
  AND U16713 ( .A(n25123), .B(n25122), .Z(n56672) );
  NANDN U16714 ( .A(y[4430]), .B(x[4430]), .Z(n9776) );
  NANDN U16715 ( .A(y[4431]), .B(x[4431]), .Z(n41343) );
  NAND U16716 ( .A(n9776), .B(n41343), .Z(n56670) );
  NANDN U16717 ( .A(y[4428]), .B(x[4428]), .Z(n9777) );
  NANDN U16718 ( .A(y[4429]), .B(x[4429]), .Z(n41337) );
  AND U16719 ( .A(n9777), .B(n41337), .Z(n56667) );
  XNOR U16720 ( .A(x[4428]), .B(y[4428]), .Z(n25125) );
  NANDN U16721 ( .A(y[4426]), .B(x[4426]), .Z(n9778) );
  NANDN U16722 ( .A(y[4427]), .B(x[4427]), .Z(n25124) );
  AND U16723 ( .A(n9778), .B(n25124), .Z(n51626) );
  XNOR U16724 ( .A(y[4424]), .B(x[4424]), .Z(n25133) );
  NANDN U16725 ( .A(x[4423]), .B(y[4423]), .Z(n41320) );
  NAND U16726 ( .A(n25133), .B(n41320), .Z(n56663) );
  NANDN U16727 ( .A(y[4422]), .B(x[4422]), .Z(n9779) );
  NANDN U16728 ( .A(y[4423]), .B(x[4423]), .Z(n25132) );
  AND U16729 ( .A(n9779), .B(n25132), .Z(n51628) );
  NANDN U16730 ( .A(x[4417]), .B(y[4417]), .Z(n25140) );
  NANDN U16731 ( .A(x[4418]), .B(y[4418]), .Z(n41309) );
  NAND U16732 ( .A(n25140), .B(n41309), .Z(n56658) );
  NANDN U16733 ( .A(y[4416]), .B(x[4416]), .Z(n25142) );
  NANDN U16734 ( .A(y[4417]), .B(x[4417]), .Z(n25139) );
  AND U16735 ( .A(n25142), .B(n25139), .Z(n51630) );
  NANDN U16736 ( .A(y[4412]), .B(x[4412]), .Z(n9780) );
  NANDN U16737 ( .A(y[4413]), .B(x[4413]), .Z(n41294) );
  AND U16738 ( .A(n9780), .B(n41294), .Z(n56654) );
  ANDN U16739 ( .B(y[4411]), .A(x[4411]), .Z(n25144) );
  NANDN U16740 ( .A(x[4409]), .B(y[4409]), .Z(n25146) );
  NANDN U16741 ( .A(x[4410]), .B(y[4410]), .Z(n25145) );
  NAND U16742 ( .A(n25146), .B(n25145), .Z(n51633) );
  NANDN U16743 ( .A(y[4408]), .B(x[4408]), .Z(n9781) );
  NANDN U16744 ( .A(y[4409]), .B(x[4409]), .Z(n41284) );
  AND U16745 ( .A(n9781), .B(n41284), .Z(n56649) );
  ANDN U16746 ( .B(y[4407]), .A(x[4407]), .Z(n51634) );
  XNOR U16747 ( .A(x[4408]), .B(y[4408]), .Z(n41277) );
  NANDN U16748 ( .A(n51634), .B(n41277), .Z(n16254) );
  XNOR U16749 ( .A(x[4406]), .B(y[4406]), .Z(n25148) );
  NANDN U16750 ( .A(y[4404]), .B(x[4404]), .Z(n9782) );
  NANDN U16751 ( .A(y[4405]), .B(x[4405]), .Z(n25147) );
  AND U16752 ( .A(n9782), .B(n25147), .Z(n51636) );
  XNOR U16753 ( .A(y[4404]), .B(x[4404]), .Z(n25152) );
  NANDN U16754 ( .A(x[4403]), .B(y[4403]), .Z(n25153) );
  AND U16755 ( .A(n25152), .B(n25153), .Z(n56645) );
  NANDN U16756 ( .A(y[4402]), .B(x[4402]), .Z(n9783) );
  NANDN U16757 ( .A(y[4403]), .B(x[4403]), .Z(n25151) );
  NAND U16758 ( .A(n9783), .B(n25151), .Z(n56644) );
  XNOR U16759 ( .A(y[4402]), .B(x[4402]), .Z(n41263) );
  NANDN U16760 ( .A(x[4401]), .B(y[4401]), .Z(n25155) );
  AND U16761 ( .A(n41263), .B(n25155), .Z(n56643) );
  NANDN U16762 ( .A(y[4400]), .B(x[4400]), .Z(n9784) );
  NANDN U16763 ( .A(y[4401]), .B(x[4401]), .Z(n41262) );
  NAND U16764 ( .A(n9784), .B(n41262), .Z(n56642) );
  XOR U16765 ( .A(y[4400]), .B(x[4400]), .Z(n41259) );
  ANDN U16766 ( .B(y[4399]), .A(x[4399]), .Z(n41253) );
  NOR U16767 ( .A(n41259), .B(n41253), .Z(n56641) );
  XNOR U16768 ( .A(y[4398]), .B(x[4398]), .Z(n25158) );
  NANDN U16769 ( .A(x[4397]), .B(y[4397]), .Z(n41246) );
  AND U16770 ( .A(n25158), .B(n41246), .Z(n56639) );
  NANDN U16771 ( .A(y[4396]), .B(x[4396]), .Z(n9785) );
  NANDN U16772 ( .A(y[4397]), .B(x[4397]), .Z(n25157) );
  NAND U16773 ( .A(n9785), .B(n25157), .Z(n56637) );
  XNOR U16774 ( .A(y[4396]), .B(x[4396]), .Z(n25160) );
  NANDN U16775 ( .A(x[4395]), .B(y[4395]), .Z(n41242) );
  AND U16776 ( .A(n25160), .B(n41242), .Z(n56636) );
  XNOR U16777 ( .A(x[4394]), .B(y[4394]), .Z(n25162) );
  NANDN U16778 ( .A(x[4393]), .B(y[4393]), .Z(n56633) );
  AND U16779 ( .A(n25162), .B(n56633), .Z(n16235) );
  NANDN U16780 ( .A(x[4392]), .B(y[4392]), .Z(n41236) );
  ANDN U16781 ( .B(y[4391]), .A(x[4391]), .Z(n41233) );
  ANDN U16782 ( .B(n41236), .A(n41233), .Z(n56631) );
  NANDN U16783 ( .A(y[4390]), .B(x[4390]), .Z(n9786) );
  NANDN U16784 ( .A(y[4391]), .B(x[4391]), .Z(n25164) );
  NAND U16785 ( .A(n9786), .B(n25164), .Z(n56630) );
  NANDN U16786 ( .A(x[4389]), .B(y[4389]), .Z(n25165) );
  NANDN U16787 ( .A(x[4390]), .B(y[4390]), .Z(n9787) );
  AND U16788 ( .A(n25165), .B(n9787), .Z(n51637) );
  NANDN U16789 ( .A(y[4386]), .B(x[4386]), .Z(n9788) );
  NANDN U16790 ( .A(y[4387]), .B(x[4387]), .Z(n41222) );
  NAND U16791 ( .A(n9788), .B(n41222), .Z(n56628) );
  NANDN U16792 ( .A(y[4384]), .B(x[4384]), .Z(n9789) );
  NANDN U16793 ( .A(y[4385]), .B(x[4385]), .Z(n41216) );
  AND U16794 ( .A(n9789), .B(n41216), .Z(n56625) );
  ANDN U16795 ( .B(y[4383]), .A(x[4383]), .Z(n41204) );
  XNOR U16796 ( .A(y[4384]), .B(x[4384]), .Z(n25170) );
  NANDN U16797 ( .A(n41204), .B(n25170), .Z(n56624) );
  NANDN U16798 ( .A(y[4382]), .B(x[4382]), .Z(n9790) );
  NANDN U16799 ( .A(y[4383]), .B(x[4383]), .Z(n25169) );
  AND U16800 ( .A(n9790), .B(n25169), .Z(n51639) );
  NANDN U16801 ( .A(x[4377]), .B(y[4377]), .Z(n25175) );
  NANDN U16802 ( .A(x[4378]), .B(y[4378]), .Z(n41192) );
  NAND U16803 ( .A(n25175), .B(n41192), .Z(n56620) );
  NANDN U16804 ( .A(y[4376]), .B(x[4376]), .Z(n25177) );
  NANDN U16805 ( .A(y[4377]), .B(x[4377]), .Z(n25174) );
  AND U16806 ( .A(n25177), .B(n25174), .Z(n51641) );
  NANDN U16807 ( .A(y[4372]), .B(x[4372]), .Z(n25180) );
  ANDN U16808 ( .B(x[4373]), .A(y[4373]), .Z(n41178) );
  ANDN U16809 ( .B(n25180), .A(n41178), .Z(n56615) );
  NANDN U16810 ( .A(x[4371]), .B(y[4371]), .Z(n25182) );
  NANDN U16811 ( .A(x[4372]), .B(y[4372]), .Z(n25179) );
  NAND U16812 ( .A(n25182), .B(n25179), .Z(n56614) );
  NANDN U16813 ( .A(y[4371]), .B(x[4371]), .Z(n25181) );
  ANDN U16814 ( .B(x[4370]), .A(y[4370]), .Z(n41168) );
  ANDN U16815 ( .B(n25181), .A(n41168), .Z(n56613) );
  ANDN U16816 ( .B(x[4368]), .A(y[4368]), .Z(n41162) );
  ANDN U16817 ( .B(x[4369]), .A(y[4369]), .Z(n41169) );
  NOR U16818 ( .A(n41162), .B(n41169), .Z(n56612) );
  NANDN U16819 ( .A(y[4366]), .B(x[4366]), .Z(n9791) );
  ANDN U16820 ( .B(x[4367]), .A(y[4367]), .Z(n41163) );
  ANDN U16821 ( .B(n9791), .A(n41163), .Z(n56610) );
  XNOR U16822 ( .A(x[4366]), .B(y[4366]), .Z(n25187) );
  ANDN U16823 ( .B(y[4365]), .A(x[4365]), .Z(n25188) );
  ANDN U16824 ( .B(n25187), .A(n25188), .Z(n16202) );
  XNOR U16825 ( .A(x[4364]), .B(y[4364]), .Z(n25190) );
  NANDN U16826 ( .A(y[4362]), .B(x[4362]), .Z(n9792) );
  NANDN U16827 ( .A(y[4363]), .B(x[4363]), .Z(n25189) );
  NAND U16828 ( .A(n9792), .B(n25189), .Z(n56605) );
  XNOR U16829 ( .A(y[4362]), .B(x[4362]), .Z(n41147) );
  NANDN U16830 ( .A(x[4361]), .B(y[4361]), .Z(n25192) );
  AND U16831 ( .A(n41147), .B(n25192), .Z(n56604) );
  NANDN U16832 ( .A(y[4360]), .B(x[4360]), .Z(n9793) );
  NANDN U16833 ( .A(y[4361]), .B(x[4361]), .Z(n41146) );
  NAND U16834 ( .A(n9793), .B(n41146), .Z(n56602) );
  XNOR U16835 ( .A(x[4360]), .B(y[4360]), .Z(n25194) );
  NANDN U16836 ( .A(x[4359]), .B(y[4359]), .Z(n56600) );
  AND U16837 ( .A(n25194), .B(n56600), .Z(n16193) );
  NANDN U16838 ( .A(y[4356]), .B(x[4356]), .Z(n41129) );
  NANDN U16839 ( .A(y[4357]), .B(x[4357]), .Z(n25195) );
  NAND U16840 ( .A(n41129), .B(n25195), .Z(n56598) );
  NANDN U16841 ( .A(x[4355]), .B(y[4355]), .Z(n25197) );
  NANDN U16842 ( .A(x[4356]), .B(y[4356]), .Z(n41135) );
  AND U16843 ( .A(n25197), .B(n41135), .Z(n51649) );
  ANDN U16844 ( .B(x[4351]), .A(y[4351]), .Z(n41120) );
  NANDN U16845 ( .A(y[4350]), .B(x[4350]), .Z(n25199) );
  NANDN U16846 ( .A(n41120), .B(n25199), .Z(n56591) );
  NANDN U16847 ( .A(x[4350]), .B(y[4350]), .Z(n41118) );
  NANDN U16848 ( .A(x[4349]), .B(y[4349]), .Z(n25201) );
  AND U16849 ( .A(n41118), .B(n25201), .Z(n51651) );
  NANDN U16850 ( .A(y[4346]), .B(x[4346]), .Z(n41103) );
  NANDN U16851 ( .A(y[4347]), .B(x[4347]), .Z(n41110) );
  NAND U16852 ( .A(n41103), .B(n41110), .Z(n56589) );
  NANDN U16853 ( .A(x[4345]), .B(y[4345]), .Z(n25205) );
  NANDN U16854 ( .A(x[4346]), .B(y[4346]), .Z(n25204) );
  AND U16855 ( .A(n25205), .B(n25204), .Z(n51653) );
  NANDN U16856 ( .A(y[4340]), .B(x[4340]), .Z(n41085) );
  NANDN U16857 ( .A(y[4341]), .B(x[4341]), .Z(n41092) );
  NAND U16858 ( .A(n41085), .B(n41092), .Z(n56584) );
  NANDN U16859 ( .A(x[4339]), .B(y[4339]), .Z(n25211) );
  XNOR U16860 ( .A(x[4340]), .B(y[4340]), .Z(n9794) );
  AND U16861 ( .A(n25211), .B(n9794), .Z(n51655) );
  NANDN U16862 ( .A(y[4336]), .B(x[4336]), .Z(n9795) );
  NANDN U16863 ( .A(y[4337]), .B(x[4337]), .Z(n41080) );
  NAND U16864 ( .A(n9795), .B(n41080), .Z(n56580) );
  NANDN U16865 ( .A(x[4335]), .B(y[4335]), .Z(n51657) );
  XNOR U16866 ( .A(x[4336]), .B(y[4336]), .Z(n41074) );
  NANDN U16867 ( .A(y[4334]), .B(x[4334]), .Z(n25214) );
  NANDN U16868 ( .A(y[4335]), .B(x[4335]), .Z(n41073) );
  NAND U16869 ( .A(n25214), .B(n41073), .Z(n51658) );
  NANDN U16870 ( .A(x[4333]), .B(y[4333]), .Z(n41065) );
  NANDN U16871 ( .A(x[4334]), .B(y[4334]), .Z(n41071) );
  AND U16872 ( .A(n41065), .B(n41071), .Z(n56578) );
  NANDN U16873 ( .A(y[4332]), .B(x[4332]), .Z(n25216) );
  NANDN U16874 ( .A(y[4333]), .B(x[4333]), .Z(n25215) );
  NAND U16875 ( .A(n25216), .B(n25215), .Z(n56577) );
  NANDN U16876 ( .A(x[4331]), .B(y[4331]), .Z(n41059) );
  NANDN U16877 ( .A(x[4332]), .B(y[4332]), .Z(n41066) );
  AND U16878 ( .A(n41059), .B(n41066), .Z(n56576) );
  NANDN U16879 ( .A(y[4330]), .B(x[4330]), .Z(n25218) );
  NANDN U16880 ( .A(y[4331]), .B(x[4331]), .Z(n25217) );
  NAND U16881 ( .A(n25218), .B(n25217), .Z(n56575) );
  NANDN U16882 ( .A(x[4329]), .B(y[4329]), .Z(n25220) );
  NANDN U16883 ( .A(x[4330]), .B(y[4330]), .Z(n41060) );
  AND U16884 ( .A(n25220), .B(n41060), .Z(n56574) );
  NANDN U16885 ( .A(y[4328]), .B(x[4328]), .Z(n25222) );
  NANDN U16886 ( .A(y[4329]), .B(x[4329]), .Z(n25219) );
  NAND U16887 ( .A(n25222), .B(n25219), .Z(n56573) );
  NANDN U16888 ( .A(x[4327]), .B(y[4327]), .Z(n41049) );
  NANDN U16889 ( .A(x[4328]), .B(y[4328]), .Z(n25221) );
  AND U16890 ( .A(n41049), .B(n25221), .Z(n56572) );
  XNOR U16891 ( .A(y[4326]), .B(x[4326]), .Z(n41046) );
  NANDN U16892 ( .A(x[4325]), .B(y[4325]), .Z(n41040) );
  AND U16893 ( .A(n41046), .B(n41040), .Z(n56569) );
  ANDN U16894 ( .B(x[4325]), .A(y[4325]), .Z(n41045) );
  NANDN U16895 ( .A(y[4324]), .B(x[4324]), .Z(n9796) );
  NANDN U16896 ( .A(n41045), .B(n9796), .Z(n56568) );
  XNOR U16897 ( .A(y[4324]), .B(x[4324]), .Z(n41037) );
  NANDN U16898 ( .A(x[4323]), .B(y[4323]), .Z(n41033) );
  AND U16899 ( .A(n41037), .B(n41033), .Z(n56567) );
  NANDN U16900 ( .A(y[4322]), .B(x[4322]), .Z(n9797) );
  NANDN U16901 ( .A(y[4323]), .B(x[4323]), .Z(n41036) );
  NAND U16902 ( .A(n9797), .B(n41036), .Z(n56566) );
  NANDN U16903 ( .A(x[4321]), .B(y[4321]), .Z(n56564) );
  XNOR U16904 ( .A(x[4322]), .B(y[4322]), .Z(n41030) );
  AND U16905 ( .A(n56564), .B(n41030), .Z(n16147) );
  NANDN U16906 ( .A(y[4320]), .B(x[4320]), .Z(n25224) );
  NANDN U16907 ( .A(y[4321]), .B(x[4321]), .Z(n41031) );
  NAND U16908 ( .A(n25224), .B(n41031), .Z(n56563) );
  NANDN U16909 ( .A(x[4319]), .B(y[4319]), .Z(n41020) );
  NANDN U16910 ( .A(x[4320]), .B(y[4320]), .Z(n41026) );
  AND U16911 ( .A(n41020), .B(n41026), .Z(n56562) );
  NANDN U16912 ( .A(y[4318]), .B(x[4318]), .Z(n41016) );
  NANDN U16913 ( .A(y[4319]), .B(x[4319]), .Z(n25225) );
  NAND U16914 ( .A(n41016), .B(n25225), .Z(n56561) );
  NANDN U16915 ( .A(x[4317]), .B(y[4317]), .Z(n41015) );
  XNOR U16916 ( .A(y[4318]), .B(x[4318]), .Z(n9798) );
  AND U16917 ( .A(n41015), .B(n9798), .Z(n56560) );
  NANDN U16918 ( .A(y[4316]), .B(x[4316]), .Z(n25226) );
  NANDN U16919 ( .A(y[4317]), .B(x[4317]), .Z(n41017) );
  NAND U16920 ( .A(n25226), .B(n41017), .Z(n56559) );
  NANDN U16921 ( .A(x[4315]), .B(y[4315]), .Z(n41006) );
  XNOR U16922 ( .A(y[4316]), .B(x[4316]), .Z(n9799) );
  AND U16923 ( .A(n41006), .B(n9799), .Z(n56558) );
  NANDN U16924 ( .A(y[4314]), .B(x[4314]), .Z(n25228) );
  NANDN U16925 ( .A(y[4315]), .B(x[4315]), .Z(n25227) );
  NAND U16926 ( .A(n25228), .B(n25227), .Z(n56557) );
  NANDN U16927 ( .A(x[4313]), .B(y[4313]), .Z(n41000) );
  NANDN U16928 ( .A(x[4314]), .B(y[4314]), .Z(n41007) );
  AND U16929 ( .A(n41000), .B(n41007), .Z(n56556) );
  NANDN U16930 ( .A(y[4312]), .B(x[4312]), .Z(n25230) );
  NANDN U16931 ( .A(y[4313]), .B(x[4313]), .Z(n25229) );
  NAND U16932 ( .A(n25230), .B(n25229), .Z(n56555) );
  NANDN U16933 ( .A(x[4311]), .B(y[4311]), .Z(n40994) );
  NANDN U16934 ( .A(x[4312]), .B(y[4312]), .Z(n41001) );
  AND U16935 ( .A(n40994), .B(n41001), .Z(n56554) );
  NANDN U16936 ( .A(y[4308]), .B(x[4308]), .Z(n40984) );
  NANDN U16937 ( .A(y[4309]), .B(x[4309]), .Z(n25233) );
  NAND U16938 ( .A(n40984), .B(n25233), .Z(n51660) );
  NANDN U16939 ( .A(x[4307]), .B(y[4307]), .Z(n25234) );
  NANDN U16940 ( .A(x[4308]), .B(y[4308]), .Z(n40989) );
  AND U16941 ( .A(n25234), .B(n40989), .Z(n56551) );
  NANDN U16942 ( .A(y[4306]), .B(x[4306]), .Z(n25236) );
  NANDN U16943 ( .A(y[4307]), .B(x[4307]), .Z(n40985) );
  NAND U16944 ( .A(n25236), .B(n40985), .Z(n56550) );
  NANDN U16945 ( .A(x[4305]), .B(y[4305]), .Z(n40977) );
  NANDN U16946 ( .A(x[4306]), .B(y[4306]), .Z(n25235) );
  AND U16947 ( .A(n40977), .B(n25235), .Z(n56549) );
  NANDN U16948 ( .A(y[4304]), .B(x[4304]), .Z(n9800) );
  NANDN U16949 ( .A(y[4305]), .B(x[4305]), .Z(n25237) );
  NAND U16950 ( .A(n9800), .B(n25237), .Z(n56548) );
  XNOR U16951 ( .A(x[4304]), .B(y[4304]), .Z(n40975) );
  ANDN U16952 ( .B(x[4303]), .A(y[4303]), .Z(n40974) );
  NANDN U16953 ( .A(y[4302]), .B(x[4302]), .Z(n9801) );
  NANDN U16954 ( .A(n40974), .B(n9801), .Z(n56547) );
  XNOR U16955 ( .A(x[4302]), .B(y[4302]), .Z(n25239) );
  NANDN U16956 ( .A(x[4301]), .B(y[4301]), .Z(n56545) );
  NANDN U16957 ( .A(y[4300]), .B(x[4300]), .Z(n9802) );
  NANDN U16958 ( .A(y[4301]), .B(x[4301]), .Z(n25238) );
  AND U16959 ( .A(n9802), .B(n25238), .Z(n56544) );
  NANDN U16960 ( .A(x[4299]), .B(y[4299]), .Z(n25241) );
  XOR U16961 ( .A(y[4300]), .B(x[4300]), .Z(n40964) );
  ANDN U16962 ( .B(n25241), .A(n40964), .Z(n56543) );
  NANDN U16963 ( .A(x[4297]), .B(y[4297]), .Z(n25243) );
  XOR U16964 ( .A(y[4298]), .B(x[4298]), .Z(n40958) );
  ANDN U16965 ( .B(n25243), .A(n40958), .Z(n56541) );
  ANDN U16966 ( .B(x[4297]), .A(y[4297]), .Z(n40959) );
  NANDN U16967 ( .A(y[4296]), .B(x[4296]), .Z(n25245) );
  NANDN U16968 ( .A(n40959), .B(n25245), .Z(n51663) );
  NANDN U16969 ( .A(x[4296]), .B(y[4296]), .Z(n25244) );
  ANDN U16970 ( .B(y[4295]), .A(x[4295]), .Z(n25247) );
  ANDN U16971 ( .B(n25244), .A(n25247), .Z(n56540) );
  NANDN U16972 ( .A(y[4292]), .B(x[4292]), .Z(n40941) );
  NANDN U16973 ( .A(y[4293]), .B(x[4293]), .Z(n40947) );
  NAND U16974 ( .A(n40941), .B(n40947), .Z(n56535) );
  NANDN U16975 ( .A(y[4290]), .B(x[4290]), .Z(n25251) );
  NANDN U16976 ( .A(y[4291]), .B(x[4291]), .Z(n40942) );
  AND U16977 ( .A(n25251), .B(n40942), .Z(n56534) );
  ANDN U16978 ( .B(y[4289]), .A(x[4289]), .Z(n40932) );
  NANDN U16979 ( .A(x[4290]), .B(y[4290]), .Z(n40938) );
  NANDN U16980 ( .A(n40932), .B(n40938), .Z(n56533) );
  NANDN U16981 ( .A(y[4288]), .B(x[4288]), .Z(n25253) );
  NANDN U16982 ( .A(y[4289]), .B(x[4289]), .Z(n25252) );
  AND U16983 ( .A(n25253), .B(n25252), .Z(n56532) );
  ANDN U16984 ( .B(y[4288]), .A(x[4288]), .Z(n40933) );
  NANDN U16985 ( .A(x[4287]), .B(y[4287]), .Z(n40926) );
  NANDN U16986 ( .A(n40933), .B(n40926), .Z(n56531) );
  NANDN U16987 ( .A(y[4286]), .B(x[4286]), .Z(n25255) );
  NANDN U16988 ( .A(y[4287]), .B(x[4287]), .Z(n25254) );
  AND U16989 ( .A(n25255), .B(n25254), .Z(n56530) );
  NANDN U16990 ( .A(x[4283]), .B(y[4283]), .Z(n25259) );
  NANDN U16991 ( .A(x[4284]), .B(y[4284]), .Z(n40921) );
  NAND U16992 ( .A(n25259), .B(n40921), .Z(n51667) );
  NANDN U16993 ( .A(y[4282]), .B(x[4282]), .Z(n25261) );
  NANDN U16994 ( .A(y[4283]), .B(x[4283]), .Z(n25258) );
  AND U16995 ( .A(n25261), .B(n25258), .Z(n56529) );
  XNOR U16996 ( .A(y[4280]), .B(x[4280]), .Z(n40907) );
  NANDN U16997 ( .A(x[4279]), .B(y[4279]), .Z(n25263) );
  NAND U16998 ( .A(n40907), .B(n25263), .Z(n56524) );
  NANDN U16999 ( .A(x[4277]), .B(y[4277]), .Z(n25265) );
  XNOR U17000 ( .A(y[4278]), .B(x[4278]), .Z(n9803) );
  AND U17001 ( .A(n25265), .B(n9803), .Z(n56522) );
  NANDN U17002 ( .A(y[4276]), .B(x[4276]), .Z(n40894) );
  NANDN U17003 ( .A(y[4277]), .B(x[4277]), .Z(n40901) );
  NAND U17004 ( .A(n40894), .B(n40901), .Z(n56521) );
  NANDN U17005 ( .A(x[4275]), .B(y[4275]), .Z(n25267) );
  NANDN U17006 ( .A(x[4276]), .B(y[4276]), .Z(n25266) );
  AND U17007 ( .A(n25267), .B(n25266), .Z(n56520) );
  NANDN U17008 ( .A(y[4274]), .B(x[4274]), .Z(n9804) );
  NANDN U17009 ( .A(y[4275]), .B(x[4275]), .Z(n40895) );
  NAND U17010 ( .A(n9804), .B(n40895), .Z(n56519) );
  ANDN U17011 ( .B(y[4273]), .A(x[4273]), .Z(n25268) );
  NANDN U17012 ( .A(y[4272]), .B(x[4272]), .Z(n25270) );
  NANDN U17013 ( .A(y[4273]), .B(x[4273]), .Z(n40889) );
  AND U17014 ( .A(n25270), .B(n40889), .Z(n56516) );
  NANDN U17015 ( .A(x[4271]), .B(y[4271]), .Z(n25272) );
  NANDN U17016 ( .A(x[4272]), .B(y[4272]), .Z(n25269) );
  NAND U17017 ( .A(n25272), .B(n25269), .Z(n56515) );
  NANDN U17018 ( .A(y[4270]), .B(x[4270]), .Z(n9805) );
  NANDN U17019 ( .A(y[4271]), .B(x[4271]), .Z(n25271) );
  AND U17020 ( .A(n9805), .B(n25271), .Z(n56514) );
  XNOR U17021 ( .A(x[4270]), .B(y[4270]), .Z(n25274) );
  NANDN U17022 ( .A(y[4268]), .B(x[4268]), .Z(n25277) );
  NANDN U17023 ( .A(y[4269]), .B(x[4269]), .Z(n25273) );
  NAND U17024 ( .A(n25277), .B(n25273), .Z(n56513) );
  NANDN U17025 ( .A(x[4267]), .B(y[4267]), .Z(n40872) );
  NANDN U17026 ( .A(x[4268]), .B(y[4268]), .Z(n25276) );
  AND U17027 ( .A(n40872), .B(n25276), .Z(n56512) );
  NANDN U17028 ( .A(y[4266]), .B(x[4266]), .Z(n25279) );
  NANDN U17029 ( .A(y[4267]), .B(x[4267]), .Z(n25278) );
  NAND U17030 ( .A(n25279), .B(n25278), .Z(n56510) );
  XNOR U17031 ( .A(y[4266]), .B(x[4266]), .Z(n9806) );
  ANDN U17032 ( .B(y[4265]), .A(x[4265]), .Z(n40866) );
  ANDN U17033 ( .B(n9806), .A(n40866), .Z(n56509) );
  NANDN U17034 ( .A(y[4264]), .B(x[4264]), .Z(n9807) );
  NANDN U17035 ( .A(y[4265]), .B(x[4265]), .Z(n25280) );
  AND U17036 ( .A(n9807), .B(n25280), .Z(n56508) );
  NANDN U17037 ( .A(x[4259]), .B(y[4259]), .Z(n40849) );
  ANDN U17038 ( .B(y[4260]), .A(x[4260]), .Z(n40858) );
  ANDN U17039 ( .B(n40849), .A(n40858), .Z(n56505) );
  NANDN U17040 ( .A(x[4255]), .B(y[4255]), .Z(n40835) );
  NANDN U17041 ( .A(x[4256]), .B(y[4256]), .Z(n40843) );
  AND U17042 ( .A(n40835), .B(n40843), .Z(n56500) );
  NANDN U17043 ( .A(y[4254]), .B(x[4254]), .Z(n25289) );
  NANDN U17044 ( .A(y[4255]), .B(x[4255]), .Z(n25288) );
  NAND U17045 ( .A(n25289), .B(n25288), .Z(n56499) );
  NANDN U17046 ( .A(x[4253]), .B(y[4253]), .Z(n40829) );
  NANDN U17047 ( .A(x[4254]), .B(y[4254]), .Z(n40836) );
  AND U17048 ( .A(n40829), .B(n40836), .Z(n51672) );
  NANDN U17049 ( .A(y[4250]), .B(x[4250]), .Z(n25293) );
  NANDN U17050 ( .A(y[4251]), .B(x[4251]), .Z(n40826) );
  NAND U17051 ( .A(n25293), .B(n40826), .Z(n56495) );
  NANDN U17052 ( .A(x[4249]), .B(y[4249]), .Z(n40818) );
  NANDN U17053 ( .A(x[4250]), .B(y[4250]), .Z(n25292) );
  AND U17054 ( .A(n40818), .B(n25292), .Z(n56494) );
  XNOR U17055 ( .A(x[4248]), .B(y[4248]), .Z(n40816) );
  NANDN U17056 ( .A(x[4247]), .B(y[4247]), .Z(n51674) );
  AND U17057 ( .A(n40816), .B(n51674), .Z(n16060) );
  XNOR U17058 ( .A(y[4246]), .B(x[4246]), .Z(n40809) );
  NANDN U17059 ( .A(x[4245]), .B(y[4245]), .Z(n25295) );
  AND U17060 ( .A(n40809), .B(n25295), .Z(n56491) );
  ANDN U17061 ( .B(x[4245]), .A(y[4245]), .Z(n40808) );
  NANDN U17062 ( .A(y[4244]), .B(x[4244]), .Z(n25298) );
  NANDN U17063 ( .A(n40808), .B(n25298), .Z(n56490) );
  NANDN U17064 ( .A(x[4243]), .B(y[4243]), .Z(n25299) );
  NANDN U17065 ( .A(x[4244]), .B(y[4244]), .Z(n25296) );
  AND U17066 ( .A(n25299), .B(n25296), .Z(n56489) );
  NANDN U17067 ( .A(y[4242]), .B(x[4242]), .Z(n40797) );
  NANDN U17068 ( .A(y[4243]), .B(x[4243]), .Z(n25297) );
  NAND U17069 ( .A(n40797), .B(n25297), .Z(n56488) );
  NANDN U17070 ( .A(x[4241]), .B(y[4241]), .Z(n40794) );
  NANDN U17071 ( .A(x[4242]), .B(y[4242]), .Z(n25300) );
  AND U17072 ( .A(n40794), .B(n25300), .Z(n56487) );
  NANDN U17073 ( .A(x[4239]), .B(y[4239]), .Z(n25303) );
  NANDN U17074 ( .A(x[4240]), .B(y[4240]), .Z(n40796) );
  AND U17075 ( .A(n25303), .B(n40796), .Z(n56485) );
  NANDN U17076 ( .A(y[4238]), .B(x[4238]), .Z(n9808) );
  NANDN U17077 ( .A(y[4239]), .B(x[4239]), .Z(n25302) );
  NAND U17078 ( .A(n9808), .B(n25302), .Z(n56484) );
  XNOR U17079 ( .A(y[4238]), .B(x[4238]), .Z(n40786) );
  NANDN U17080 ( .A(x[4237]), .B(y[4237]), .Z(n25305) );
  AND U17081 ( .A(n40786), .B(n25305), .Z(n56482) );
  ANDN U17082 ( .B(x[4237]), .A(y[4237]), .Z(n40788) );
  NANDN U17083 ( .A(y[4236]), .B(x[4236]), .Z(n9809) );
  NANDN U17084 ( .A(n40788), .B(n9809), .Z(n56480) );
  NANDN U17085 ( .A(x[4235]), .B(y[4235]), .Z(n51676) );
  XNOR U17086 ( .A(x[4236]), .B(y[4236]), .Z(n40780) );
  AND U17087 ( .A(n51676), .B(n40780), .Z(n16046) );
  NANDN U17088 ( .A(y[4234]), .B(x[4234]), .Z(n25307) );
  NANDN U17089 ( .A(y[4235]), .B(x[4235]), .Z(n40781) );
  NAND U17090 ( .A(n25307), .B(n40781), .Z(n56476) );
  NANDN U17091 ( .A(x[4233]), .B(y[4233]), .Z(n25309) );
  NANDN U17092 ( .A(x[4234]), .B(y[4234]), .Z(n25306) );
  AND U17093 ( .A(n25309), .B(n25306), .Z(n56474) );
  NANDN U17094 ( .A(y[4232]), .B(x[4232]), .Z(n9810) );
  NANDN U17095 ( .A(y[4233]), .B(x[4233]), .Z(n25308) );
  NAND U17096 ( .A(n9810), .B(n25308), .Z(n56472) );
  NANDN U17097 ( .A(x[4231]), .B(y[4231]), .Z(n56470) );
  XNOR U17098 ( .A(x[4232]), .B(y[4232]), .Z(n25311) );
  NANDN U17099 ( .A(y[4230]), .B(x[4230]), .Z(n40765) );
  NANDN U17100 ( .A(y[4231]), .B(x[4231]), .Z(n25310) );
  AND U17101 ( .A(n40765), .B(n25310), .Z(n56466) );
  NANDN U17102 ( .A(x[4229]), .B(y[4229]), .Z(n40762) );
  XNOR U17103 ( .A(x[4230]), .B(y[4230]), .Z(n9811) );
  NAND U17104 ( .A(n40762), .B(n9811), .Z(n56464) );
  NANDN U17105 ( .A(y[4228]), .B(x[4228]), .Z(n25313) );
  NANDN U17106 ( .A(y[4229]), .B(x[4229]), .Z(n40766) );
  AND U17107 ( .A(n25313), .B(n40766), .Z(n56462) );
  NANDN U17108 ( .A(x[4227]), .B(y[4227]), .Z(n40756) );
  NANDN U17109 ( .A(x[4228]), .B(y[4228]), .Z(n40763) );
  NAND U17110 ( .A(n40756), .B(n40763), .Z(n56460) );
  NANDN U17111 ( .A(y[4226]), .B(x[4226]), .Z(n25315) );
  NANDN U17112 ( .A(y[4227]), .B(x[4227]), .Z(n25314) );
  AND U17113 ( .A(n25315), .B(n25314), .Z(n56458) );
  NANDN U17114 ( .A(x[4225]), .B(y[4225]), .Z(n40750) );
  NANDN U17115 ( .A(x[4226]), .B(y[4226]), .Z(n40757) );
  NAND U17116 ( .A(n40750), .B(n40757), .Z(n56456) );
  NANDN U17117 ( .A(y[4224]), .B(x[4224]), .Z(n25317) );
  NANDN U17118 ( .A(y[4225]), .B(x[4225]), .Z(n25316) );
  AND U17119 ( .A(n25317), .B(n25316), .Z(n56453) );
  NANDN U17120 ( .A(x[4223]), .B(y[4223]), .Z(n25319) );
  NANDN U17121 ( .A(x[4224]), .B(y[4224]), .Z(n40751) );
  AND U17122 ( .A(n25319), .B(n40751), .Z(n56452) );
  ANDN U17123 ( .B(x[4222]), .A(y[4222]), .Z(n40741) );
  NANDN U17124 ( .A(y[4223]), .B(x[4223]), .Z(n25318) );
  NANDN U17125 ( .A(n40741), .B(n25318), .Z(n56450) );
  NANDN U17126 ( .A(x[4221]), .B(y[4221]), .Z(n40738) );
  NANDN U17127 ( .A(x[4222]), .B(y[4222]), .Z(n25320) );
  AND U17128 ( .A(n40738), .B(n25320), .Z(n56448) );
  ANDN U17129 ( .B(x[4221]), .A(y[4221]), .Z(n40744) );
  NANDN U17130 ( .A(y[4220]), .B(x[4220]), .Z(n9812) );
  NANDN U17131 ( .A(n40744), .B(n9812), .Z(n56446) );
  XNOR U17132 ( .A(y[4220]), .B(x[4220]), .Z(n40734) );
  NANDN U17133 ( .A(x[4219]), .B(y[4219]), .Z(n25321) );
  AND U17134 ( .A(n40734), .B(n25321), .Z(n56444) );
  NANDN U17135 ( .A(x[4217]), .B(y[4217]), .Z(n25323) );
  NANDN U17136 ( .A(x[4218]), .B(y[4218]), .Z(n25322) );
  AND U17137 ( .A(n25323), .B(n25322), .Z(n56442) );
  NANDN U17138 ( .A(y[4216]), .B(x[4216]), .Z(n40722) );
  NANDN U17139 ( .A(y[4217]), .B(x[4217]), .Z(n40729) );
  NAND U17140 ( .A(n40722), .B(n40729), .Z(n56441) );
  NANDN U17141 ( .A(x[4216]), .B(y[4216]), .Z(n25324) );
  ANDN U17142 ( .B(y[4215]), .A(x[4215]), .Z(n40720) );
  ANDN U17143 ( .B(n25324), .A(n40720), .Z(n56440) );
  NANDN U17144 ( .A(y[4214]), .B(x[4214]), .Z(n9813) );
  NANDN U17145 ( .A(y[4215]), .B(x[4215]), .Z(n40723) );
  NAND U17146 ( .A(n9813), .B(n40723), .Z(n56439) );
  NANDN U17147 ( .A(x[4213]), .B(y[4213]), .Z(n51679) );
  XNOR U17148 ( .A(x[4214]), .B(y[4214]), .Z(n25326) );
  AND U17149 ( .A(n51679), .B(n25326), .Z(n16022) );
  NANDN U17150 ( .A(y[4212]), .B(x[4212]), .Z(n25328) );
  NANDN U17151 ( .A(y[4213]), .B(x[4213]), .Z(n25325) );
  NAND U17152 ( .A(n25328), .B(n25325), .Z(n56438) );
  NANDN U17153 ( .A(x[4211]), .B(y[4211]), .Z(n25330) );
  NANDN U17154 ( .A(x[4212]), .B(y[4212]), .Z(n25327) );
  AND U17155 ( .A(n25330), .B(n25327), .Z(n56437) );
  NANDN U17156 ( .A(y[4210]), .B(x[4210]), .Z(n40706) );
  NANDN U17157 ( .A(y[4211]), .B(x[4211]), .Z(n25329) );
  AND U17158 ( .A(n40706), .B(n25329), .Z(n56436) );
  NANDN U17159 ( .A(y[4208]), .B(x[4208]), .Z(n40700) );
  NANDN U17160 ( .A(y[4209]), .B(x[4209]), .Z(n40707) );
  AND U17161 ( .A(n40700), .B(n40707), .Z(n56434) );
  NANDN U17162 ( .A(x[4207]), .B(y[4207]), .Z(n25334) );
  NANDN U17163 ( .A(x[4208]), .B(y[4208]), .Z(n25333) );
  NAND U17164 ( .A(n25334), .B(n25333), .Z(n56433) );
  NANDN U17165 ( .A(y[4206]), .B(x[4206]), .Z(n40694) );
  NANDN U17166 ( .A(y[4207]), .B(x[4207]), .Z(n40701) );
  AND U17167 ( .A(n40694), .B(n40701), .Z(n56432) );
  NANDN U17168 ( .A(x[4205]), .B(y[4205]), .Z(n25336) );
  NANDN U17169 ( .A(x[4206]), .B(y[4206]), .Z(n25335) );
  NAND U17170 ( .A(n25336), .B(n25335), .Z(n56431) );
  NANDN U17171 ( .A(y[4204]), .B(x[4204]), .Z(n9814) );
  NANDN U17172 ( .A(y[4205]), .B(x[4205]), .Z(n40695) );
  AND U17173 ( .A(n9814), .B(n40695), .Z(n56430) );
  XNOR U17174 ( .A(x[4204]), .B(y[4204]), .Z(n40689) );
  NANDN U17175 ( .A(y[4202]), .B(x[4202]), .Z(n9815) );
  NANDN U17176 ( .A(y[4203]), .B(x[4203]), .Z(n40688) );
  NAND U17177 ( .A(n9815), .B(n40688), .Z(n56424) );
  NANDN U17178 ( .A(x[4201]), .B(y[4201]), .Z(n25337) );
  XNOR U17179 ( .A(x[4202]), .B(y[4202]), .Z(n40683) );
  NANDN U17180 ( .A(y[4200]), .B(x[4200]), .Z(n25338) );
  NANDN U17181 ( .A(y[4201]), .B(x[4201]), .Z(n40682) );
  AND U17182 ( .A(n25338), .B(n40682), .Z(n56423) );
  NANDN U17183 ( .A(x[4199]), .B(y[4199]), .Z(n40674) );
  NANDN U17184 ( .A(x[4200]), .B(y[4200]), .Z(n40681) );
  NAND U17185 ( .A(n40674), .B(n40681), .Z(n56422) );
  NANDN U17186 ( .A(y[4198]), .B(x[4198]), .Z(n9816) );
  NANDN U17187 ( .A(y[4199]), .B(x[4199]), .Z(n25339) );
  AND U17188 ( .A(n9816), .B(n25339), .Z(n56421) );
  ANDN U17189 ( .B(y[4197]), .A(x[4197]), .Z(n40667) );
  XNOR U17190 ( .A(y[4198]), .B(x[4198]), .Z(n25341) );
  NANDN U17191 ( .A(n40667), .B(n25341), .Z(n56420) );
  NANDN U17192 ( .A(y[4196]), .B(x[4196]), .Z(n25342) );
  NANDN U17193 ( .A(y[4197]), .B(x[4197]), .Z(n25340) );
  AND U17194 ( .A(n25342), .B(n25340), .Z(n56419) );
  NANDN U17195 ( .A(x[4195]), .B(y[4195]), .Z(n40661) );
  NANDN U17196 ( .A(x[4196]), .B(y[4196]), .Z(n40669) );
  NAND U17197 ( .A(n40661), .B(n40669), .Z(n56418) );
  NANDN U17198 ( .A(y[4192]), .B(x[4192]), .Z(n9817) );
  NANDN U17199 ( .A(y[4193]), .B(x[4193]), .Z(n40657) );
  NAND U17200 ( .A(n9817), .B(n40657), .Z(n56415) );
  XNOR U17201 ( .A(y[4192]), .B(x[4192]), .Z(n25345) );
  NANDN U17202 ( .A(x[4191]), .B(y[4191]), .Z(n40648) );
  AND U17203 ( .A(n25345), .B(n40648), .Z(n51682) );
  NANDN U17204 ( .A(x[4189]), .B(y[4189]), .Z(n40640) );
  NANDN U17205 ( .A(x[4190]), .B(y[4190]), .Z(n40649) );
  AND U17206 ( .A(n40640), .B(n40649), .Z(n56413) );
  NANDN U17207 ( .A(x[4187]), .B(y[4187]), .Z(n40633) );
  NANDN U17208 ( .A(x[4188]), .B(y[4188]), .Z(n40642) );
  AND U17209 ( .A(n40633), .B(n40642), .Z(n56410) );
  NANDN U17210 ( .A(y[4186]), .B(x[4186]), .Z(n25348) );
  NANDN U17211 ( .A(y[4187]), .B(x[4187]), .Z(n25347) );
  NAND U17212 ( .A(n25348), .B(n25347), .Z(n56409) );
  NANDN U17213 ( .A(x[4185]), .B(y[4185]), .Z(n40627) );
  NANDN U17214 ( .A(x[4186]), .B(y[4186]), .Z(n40634) );
  AND U17215 ( .A(n40627), .B(n40634), .Z(n56408) );
  NANDN U17216 ( .A(y[4184]), .B(x[4184]), .Z(n25350) );
  NANDN U17217 ( .A(y[4185]), .B(x[4185]), .Z(n25349) );
  NAND U17218 ( .A(n25350), .B(n25349), .Z(n56407) );
  NANDN U17219 ( .A(x[4183]), .B(y[4183]), .Z(n40621) );
  NANDN U17220 ( .A(x[4184]), .B(y[4184]), .Z(n40628) );
  AND U17221 ( .A(n40621), .B(n40628), .Z(n56406) );
  NANDN U17222 ( .A(y[4182]), .B(x[4182]), .Z(n25352) );
  NANDN U17223 ( .A(y[4183]), .B(x[4183]), .Z(n25351) );
  NAND U17224 ( .A(n25352), .B(n25351), .Z(n56405) );
  NANDN U17225 ( .A(x[4179]), .B(y[4179]), .Z(n25354) );
  XNOR U17226 ( .A(x[4180]), .B(y[4180]), .Z(n9818) );
  NAND U17227 ( .A(n25354), .B(n9818), .Z(n56402) );
  NANDN U17228 ( .A(y[4178]), .B(x[4178]), .Z(n40606) );
  NANDN U17229 ( .A(y[4179]), .B(x[4179]), .Z(n40613) );
  AND U17230 ( .A(n40606), .B(n40613), .Z(n51683) );
  NANDN U17231 ( .A(y[4176]), .B(x[4176]), .Z(n40600) );
  NANDN U17232 ( .A(y[4177]), .B(x[4177]), .Z(n40607) );
  AND U17233 ( .A(n40600), .B(n40607), .Z(n56400) );
  NANDN U17234 ( .A(y[4174]), .B(x[4174]), .Z(n40592) );
  NANDN U17235 ( .A(y[4175]), .B(x[4175]), .Z(n40601) );
  AND U17236 ( .A(n40592), .B(n40601), .Z(n56398) );
  ANDN U17237 ( .B(y[4174]), .A(x[4174]), .Z(n40598) );
  NANDN U17238 ( .A(x[4173]), .B(y[4173]), .Z(n25358) );
  NANDN U17239 ( .A(n40598), .B(n25358), .Z(n56397) );
  NANDN U17240 ( .A(y[4172]), .B(x[4172]), .Z(n40585) );
  NANDN U17241 ( .A(y[4173]), .B(x[4173]), .Z(n40594) );
  AND U17242 ( .A(n40585), .B(n40594), .Z(n56396) );
  NANDN U17243 ( .A(x[4171]), .B(y[4171]), .Z(n25360) );
  NANDN U17244 ( .A(x[4172]), .B(y[4172]), .Z(n25359) );
  NAND U17245 ( .A(n25360), .B(n25359), .Z(n56394) );
  NANDN U17246 ( .A(y[4170]), .B(x[4170]), .Z(n40579) );
  NANDN U17247 ( .A(y[4171]), .B(x[4171]), .Z(n40586) );
  AND U17248 ( .A(n40579), .B(n40586), .Z(n56393) );
  NANDN U17249 ( .A(x[4169]), .B(y[4169]), .Z(n25362) );
  NANDN U17250 ( .A(x[4170]), .B(y[4170]), .Z(n25361) );
  AND U17251 ( .A(n25362), .B(n25361), .Z(n56392) );
  NANDN U17252 ( .A(x[4168]), .B(y[4168]), .Z(n25363) );
  ANDN U17253 ( .B(y[4167]), .A(x[4167]), .Z(n40571) );
  ANDN U17254 ( .B(n25363), .A(n40571), .Z(n56391) );
  XNOR U17255 ( .A(y[4166]), .B(x[4166]), .Z(n25365) );
  NANDN U17256 ( .A(x[4165]), .B(y[4165]), .Z(n25367) );
  AND U17257 ( .A(n25365), .B(n25367), .Z(n56390) );
  NANDN U17258 ( .A(y[4164]), .B(x[4164]), .Z(n25368) );
  NANDN U17259 ( .A(y[4165]), .B(x[4165]), .Z(n25364) );
  NAND U17260 ( .A(n25368), .B(n25364), .Z(n51686) );
  NANDN U17261 ( .A(x[4163]), .B(y[4163]), .Z(n25370) );
  NANDN U17262 ( .A(x[4164]), .B(y[4164]), .Z(n25366) );
  AND U17263 ( .A(n25370), .B(n25366), .Z(n51687) );
  NANDN U17264 ( .A(y[4160]), .B(x[4160]), .Z(n40551) );
  NANDN U17265 ( .A(y[4161]), .B(x[4161]), .Z(n40558) );
  NAND U17266 ( .A(n40551), .B(n40558), .Z(n56388) );
  NANDN U17267 ( .A(y[4158]), .B(x[4158]), .Z(n9819) );
  NANDN U17268 ( .A(y[4159]), .B(x[4159]), .Z(n40552) );
  AND U17269 ( .A(n9819), .B(n40552), .Z(n56385) );
  XNOR U17270 ( .A(y[4158]), .B(x[4158]), .Z(n40546) );
  NANDN U17271 ( .A(x[4157]), .B(y[4157]), .Z(n25376) );
  NAND U17272 ( .A(n40546), .B(n25376), .Z(n56384) );
  NANDN U17273 ( .A(y[4156]), .B(x[4156]), .Z(n9820) );
  NANDN U17274 ( .A(y[4157]), .B(x[4157]), .Z(n40545) );
  AND U17275 ( .A(n9820), .B(n40545), .Z(n51690) );
  NANDN U17276 ( .A(y[4154]), .B(x[4154]), .Z(n9821) );
  NANDN U17277 ( .A(y[4155]), .B(x[4155]), .Z(n40539) );
  AND U17278 ( .A(n9821), .B(n40539), .Z(n56383) );
  XNOR U17279 ( .A(x[4154]), .B(y[4154]), .Z(n40534) );
  NANDN U17280 ( .A(y[4152]), .B(x[4152]), .Z(n9822) );
  NANDN U17281 ( .A(y[4153]), .B(x[4153]), .Z(n40533) );
  NAND U17282 ( .A(n9822), .B(n40533), .Z(n56382) );
  XNOR U17283 ( .A(x[4152]), .B(y[4152]), .Z(n25380) );
  ANDN U17284 ( .B(y[4151]), .A(x[4151]), .Z(n40525) );
  NANDN U17285 ( .A(x[4149]), .B(y[4149]), .Z(n40520) );
  NANDN U17286 ( .A(x[4150]), .B(y[4150]), .Z(n40527) );
  AND U17287 ( .A(n40520), .B(n40527), .Z(n56379) );
  XNOR U17288 ( .A(x[4148]), .B(y[4148]), .Z(n25384) );
  NANDN U17289 ( .A(y[4146]), .B(x[4146]), .Z(n25385) );
  NANDN U17290 ( .A(y[4147]), .B(x[4147]), .Z(n25383) );
  AND U17291 ( .A(n25385), .B(n25383), .Z(n56375) );
  NANDN U17292 ( .A(x[4143]), .B(y[4143]), .Z(n40503) );
  NANDN U17293 ( .A(x[4144]), .B(y[4144]), .Z(n40510) );
  NAND U17294 ( .A(n40503), .B(n40510), .Z(n51698) );
  NANDN U17295 ( .A(y[4142]), .B(x[4142]), .Z(n40500) );
  NANDN U17296 ( .A(y[4143]), .B(x[4143]), .Z(n25388) );
  AND U17297 ( .A(n40500), .B(n25388), .Z(n56373) );
  NANDN U17298 ( .A(x[4137]), .B(y[4137]), .Z(n25393) );
  NANDN U17299 ( .A(x[4138]), .B(y[4138]), .Z(n25392) );
  NAND U17300 ( .A(n25393), .B(n25392), .Z(n51700) );
  NANDN U17301 ( .A(y[4136]), .B(x[4136]), .Z(n25395) );
  NANDN U17302 ( .A(y[4137]), .B(x[4137]), .Z(n40489) );
  AND U17303 ( .A(n25395), .B(n40489), .Z(n56368) );
  NANDN U17304 ( .A(x[4131]), .B(y[4131]), .Z(n40468) );
  NANDN U17305 ( .A(x[4132]), .B(y[4132]), .Z(n25398) );
  NAND U17306 ( .A(n40468), .B(n25398), .Z(n51702) );
  NANDN U17307 ( .A(y[4130]), .B(x[4130]), .Z(n40463) );
  NANDN U17308 ( .A(y[4131]), .B(x[4131]), .Z(n40472) );
  AND U17309 ( .A(n40463), .B(n40472), .Z(n56363) );
  XNOR U17310 ( .A(x[4128]), .B(y[4128]), .Z(n40458) );
  NANDN U17311 ( .A(x[4127]), .B(y[4127]), .Z(n56358) );
  NAND U17312 ( .A(n40458), .B(n56358), .Z(n15923) );
  NANDN U17313 ( .A(x[4125]), .B(y[4125]), .Z(n40450) );
  NANDN U17314 ( .A(x[4126]), .B(y[4126]), .Z(n25400) );
  AND U17315 ( .A(n40450), .B(n25400), .Z(n56357) );
  NANDN U17316 ( .A(x[4123]), .B(y[4123]), .Z(n40444) );
  NANDN U17317 ( .A(x[4124]), .B(y[4124]), .Z(n40451) );
  AND U17318 ( .A(n40444), .B(n40451), .Z(n56355) );
  NANDN U17319 ( .A(y[4122]), .B(x[4122]), .Z(n25405) );
  NANDN U17320 ( .A(y[4123]), .B(x[4123]), .Z(n25404) );
  NAND U17321 ( .A(n25405), .B(n25404), .Z(n56354) );
  NANDN U17322 ( .A(x[4121]), .B(y[4121]), .Z(n40438) );
  NANDN U17323 ( .A(x[4122]), .B(y[4122]), .Z(n40445) );
  AND U17324 ( .A(n40438), .B(n40445), .Z(n56353) );
  ANDN U17325 ( .B(x[4118]), .A(y[4118]), .Z(n40428) );
  NANDN U17326 ( .A(y[4119]), .B(x[4119]), .Z(n25408) );
  NANDN U17327 ( .A(n40428), .B(n25408), .Z(n51705) );
  NANDN U17328 ( .A(y[4116]), .B(x[4116]), .Z(n25409) );
  ANDN U17329 ( .B(x[4117]), .A(y[4117]), .Z(n40430) );
  ANDN U17330 ( .B(n25409), .A(n40430), .Z(n56350) );
  NANDN U17331 ( .A(x[4115]), .B(y[4115]), .Z(n40417) );
  NANDN U17332 ( .A(x[4116]), .B(y[4116]), .Z(n40426) );
  NAND U17333 ( .A(n40417), .B(n40426), .Z(n56349) );
  NANDN U17334 ( .A(y[4114]), .B(x[4114]), .Z(n25411) );
  NANDN U17335 ( .A(y[4115]), .B(x[4115]), .Z(n25410) );
  AND U17336 ( .A(n25411), .B(n25410), .Z(n56348) );
  NANDN U17337 ( .A(x[4113]), .B(y[4113]), .Z(n40411) );
  NANDN U17338 ( .A(x[4114]), .B(y[4114]), .Z(n40418) );
  NAND U17339 ( .A(n40411), .B(n40418), .Z(n56347) );
  NANDN U17340 ( .A(y[4112]), .B(x[4112]), .Z(n25413) );
  NANDN U17341 ( .A(y[4113]), .B(x[4113]), .Z(n25412) );
  AND U17342 ( .A(n25413), .B(n25412), .Z(n56345) );
  NANDN U17343 ( .A(y[4110]), .B(x[4110]), .Z(n25415) );
  NANDN U17344 ( .A(y[4111]), .B(x[4111]), .Z(n25414) );
  AND U17345 ( .A(n25415), .B(n25414), .Z(n56343) );
  NANDN U17346 ( .A(x[4109]), .B(y[4109]), .Z(n40399) );
  NANDN U17347 ( .A(x[4110]), .B(y[4110]), .Z(n40406) );
  NAND U17348 ( .A(n40399), .B(n40406), .Z(n56342) );
  NANDN U17349 ( .A(y[4108]), .B(x[4108]), .Z(n25417) );
  NANDN U17350 ( .A(y[4109]), .B(x[4109]), .Z(n25416) );
  AND U17351 ( .A(n25417), .B(n25416), .Z(n56341) );
  NANDN U17352 ( .A(x[4105]), .B(y[4105]), .Z(n40387) );
  NANDN U17353 ( .A(x[4106]), .B(y[4106]), .Z(n40394) );
  NAND U17354 ( .A(n40387), .B(n40394), .Z(n51707) );
  NANDN U17355 ( .A(y[4104]), .B(x[4104]), .Z(n25421) );
  NANDN U17356 ( .A(y[4105]), .B(x[4105]), .Z(n25420) );
  AND U17357 ( .A(n25421), .B(n25420), .Z(n56339) );
  NANDN U17358 ( .A(x[4099]), .B(y[4099]), .Z(n25425) );
  NANDN U17359 ( .A(x[4100]), .B(y[4100]), .Z(n40376) );
  NAND U17360 ( .A(n25425), .B(n40376), .Z(n51709) );
  NANDN U17361 ( .A(y[4098]), .B(x[4098]), .Z(n40366) );
  NANDN U17362 ( .A(y[4099]), .B(x[4099]), .Z(n40373) );
  AND U17363 ( .A(n40366), .B(n40373), .Z(n56333) );
  XNOR U17364 ( .A(x[4096]), .B(y[4096]), .Z(n40360) );
  NANDN U17365 ( .A(x[4095]), .B(y[4095]), .Z(n56329) );
  NAND U17366 ( .A(n40360), .B(n56329), .Z(n15888) );
  NANDN U17367 ( .A(x[4093]), .B(y[4093]), .Z(n25431) );
  NANDN U17368 ( .A(x[4094]), .B(y[4094]), .Z(n25428) );
  AND U17369 ( .A(n25431), .B(n25428), .Z(n56328) );
  XNOR U17370 ( .A(x[4092]), .B(y[4092]), .Z(n25433) );
  NANDN U17371 ( .A(y[4090]), .B(x[4090]), .Z(n40345) );
  NANDN U17372 ( .A(y[4091]), .B(x[4091]), .Z(n25432) );
  NAND U17373 ( .A(n40345), .B(n25432), .Z(n56326) );
  ANDN U17374 ( .B(y[4087]), .A(x[4087]), .Z(n40336) );
  XNOR U17375 ( .A(y[4088]), .B(x[4088]), .Z(n40340) );
  NANDN U17376 ( .A(n40336), .B(n40340), .Z(n51714) );
  NANDN U17377 ( .A(y[4086]), .B(x[4086]), .Z(n25437) );
  NANDN U17378 ( .A(y[4087]), .B(x[4087]), .Z(n40339) );
  AND U17379 ( .A(n25437), .B(n40339), .Z(n56323) );
  NANDN U17380 ( .A(x[4081]), .B(y[4081]), .Z(n56320) );
  XNOR U17381 ( .A(x[4082]), .B(y[4082]), .Z(n25442) );
  AND U17382 ( .A(n56320), .B(n25442), .Z(n15867) );
  NANDN U17383 ( .A(y[4078]), .B(x[4078]), .Z(n25446) );
  ANDN U17384 ( .B(x[4079]), .A(y[4079]), .Z(n40318) );
  ANDN U17385 ( .B(n25446), .A(n40318), .Z(n56317) );
  NANDN U17386 ( .A(y[4076]), .B(x[4076]), .Z(n25449) );
  NANDN U17387 ( .A(y[4077]), .B(x[4077]), .Z(n25445) );
  AND U17388 ( .A(n25449), .B(n25445), .Z(n56314) );
  NANDN U17389 ( .A(x[4075]), .B(y[4075]), .Z(n40305) );
  NANDN U17390 ( .A(x[4076]), .B(y[4076]), .Z(n25448) );
  NAND U17391 ( .A(n40305), .B(n25448), .Z(n56313) );
  NANDN U17392 ( .A(y[4074]), .B(x[4074]), .Z(n40302) );
  NANDN U17393 ( .A(y[4075]), .B(x[4075]), .Z(n25450) );
  AND U17394 ( .A(n40302), .B(n25450), .Z(n56312) );
  NANDN U17395 ( .A(x[4073]), .B(y[4073]), .Z(n25451) );
  NANDN U17396 ( .A(x[4074]), .B(y[4074]), .Z(n40306) );
  NAND U17397 ( .A(n25451), .B(n40306), .Z(n56311) );
  NANDN U17398 ( .A(y[4072]), .B(x[4072]), .Z(n40296) );
  NANDN U17399 ( .A(y[4073]), .B(x[4073]), .Z(n40303) );
  AND U17400 ( .A(n40296), .B(n40303), .Z(n56310) );
  NANDN U17401 ( .A(x[4071]), .B(y[4071]), .Z(n25453) );
  NANDN U17402 ( .A(x[4072]), .B(y[4072]), .Z(n25452) );
  NAND U17403 ( .A(n25453), .B(n25452), .Z(n56309) );
  NANDN U17404 ( .A(y[4068]), .B(x[4068]), .Z(n9823) );
  NANDN U17405 ( .A(y[4069]), .B(x[4069]), .Z(n40291) );
  NAND U17406 ( .A(n9823), .B(n40291), .Z(n51720) );
  XNOR U17407 ( .A(y[4068]), .B(x[4068]), .Z(n40284) );
  NANDN U17408 ( .A(x[4067]), .B(y[4067]), .Z(n25457) );
  AND U17409 ( .A(n40284), .B(n25457), .Z(n56307) );
  NANDN U17410 ( .A(x[4063]), .B(y[4063]), .Z(n25463) );
  NANDN U17411 ( .A(x[4064]), .B(y[4064]), .Z(n25462) );
  AND U17412 ( .A(n25463), .B(n25462), .Z(n56303) );
  ANDN U17413 ( .B(x[4063]), .A(y[4063]), .Z(n40274) );
  NANDN U17414 ( .A(y[4062]), .B(x[4062]), .Z(n40267) );
  NANDN U17415 ( .A(n40274), .B(n40267), .Z(n56301) );
  NANDN U17416 ( .A(x[4061]), .B(y[4061]), .Z(n25465) );
  NANDN U17417 ( .A(x[4062]), .B(y[4062]), .Z(n25464) );
  AND U17418 ( .A(n25465), .B(n25464), .Z(n56300) );
  NANDN U17419 ( .A(y[4060]), .B(x[4060]), .Z(n9824) );
  NANDN U17420 ( .A(y[4061]), .B(x[4061]), .Z(n40268) );
  NAND U17421 ( .A(n9824), .B(n40268), .Z(n56299) );
  XNOR U17422 ( .A(y[4060]), .B(x[4060]), .Z(n40262) );
  NANDN U17423 ( .A(x[4059]), .B(y[4059]), .Z(n40258) );
  AND U17424 ( .A(n40262), .B(n40258), .Z(n56298) );
  NANDN U17425 ( .A(y[4058]), .B(x[4058]), .Z(n40253) );
  NANDN U17426 ( .A(y[4059]), .B(x[4059]), .Z(n40261) );
  NAND U17427 ( .A(n40253), .B(n40261), .Z(n56297) );
  NANDN U17428 ( .A(x[4055]), .B(y[4055]), .Z(n40244) );
  NANDN U17429 ( .A(x[4056]), .B(y[4056]), .Z(n25468) );
  NAND U17430 ( .A(n40244), .B(n25468), .Z(n51723) );
  NANDN U17431 ( .A(y[4054]), .B(x[4054]), .Z(n25469) );
  NANDN U17432 ( .A(y[4055]), .B(x[4055]), .Z(n40248) );
  AND U17433 ( .A(n25469), .B(n40248), .Z(n56295) );
  NANDN U17434 ( .A(y[4050]), .B(x[4050]), .Z(n25473) );
  NANDN U17435 ( .A(y[4051]), .B(x[4051]), .Z(n25472) );
  AND U17436 ( .A(n25473), .B(n25472), .Z(n56292) );
  NANDN U17437 ( .A(x[4049]), .B(y[4049]), .Z(n25475) );
  NANDN U17438 ( .A(x[4050]), .B(y[4050]), .Z(n40233) );
  NAND U17439 ( .A(n25475), .B(n40233), .Z(n56291) );
  NANDN U17440 ( .A(y[4048]), .B(x[4048]), .Z(n25477) );
  NANDN U17441 ( .A(y[4049]), .B(x[4049]), .Z(n25474) );
  AND U17442 ( .A(n25477), .B(n25474), .Z(n56289) );
  NANDN U17443 ( .A(x[4047]), .B(y[4047]), .Z(n40222) );
  XNOR U17444 ( .A(y[4048]), .B(x[4048]), .Z(n9825) );
  NAND U17445 ( .A(n40222), .B(n9825), .Z(n56288) );
  NANDN U17446 ( .A(y[4046]), .B(x[4046]), .Z(n9826) );
  NANDN U17447 ( .A(y[4047]), .B(x[4047]), .Z(n25478) );
  AND U17448 ( .A(n9826), .B(n25478), .Z(n56287) );
  XNOR U17449 ( .A(y[4046]), .B(x[4046]), .Z(n40218) );
  NANDN U17450 ( .A(x[4045]), .B(y[4045]), .Z(n25479) );
  NAND U17451 ( .A(n40218), .B(n25479), .Z(n56286) );
  NANDN U17452 ( .A(y[4042]), .B(x[4042]), .Z(n40206) );
  NANDN U17453 ( .A(y[4043]), .B(x[4043]), .Z(n40213) );
  NAND U17454 ( .A(n40206), .B(n40213), .Z(n51726) );
  NANDN U17455 ( .A(x[4041]), .B(y[4041]), .Z(n25483) );
  NANDN U17456 ( .A(x[4042]), .B(y[4042]), .Z(n25482) );
  AND U17457 ( .A(n25483), .B(n25482), .Z(n56284) );
  NANDN U17458 ( .A(x[4039]), .B(y[4039]), .Z(n25487) );
  NANDN U17459 ( .A(x[4040]), .B(y[4040]), .Z(n25484) );
  AND U17460 ( .A(n25487), .B(n25484), .Z(n56283) );
  ANDN U17461 ( .B(x[4037]), .A(y[4037]), .Z(n40196) );
  NANDN U17462 ( .A(y[4036]), .B(x[4036]), .Z(n40189) );
  NANDN U17463 ( .A(n40196), .B(n40189), .Z(n51730) );
  NANDN U17464 ( .A(x[4035]), .B(y[4035]), .Z(n25491) );
  NANDN U17465 ( .A(x[4036]), .B(y[4036]), .Z(n25490) );
  AND U17466 ( .A(n25491), .B(n25490), .Z(n56281) );
  XNOR U17467 ( .A(x[4034]), .B(y[4034]), .Z(n40184) );
  NANDN U17468 ( .A(x[4033]), .B(y[4033]), .Z(n56278) );
  AND U17469 ( .A(n40184), .B(n56278), .Z(n15815) );
  XNOR U17470 ( .A(x[4032]), .B(y[4032]), .Z(n40178) );
  NANDN U17471 ( .A(y[4030]), .B(x[4030]), .Z(n25493) );
  NANDN U17472 ( .A(y[4031]), .B(x[4031]), .Z(n40177) );
  NAND U17473 ( .A(n25493), .B(n40177), .Z(n51732) );
  NANDN U17474 ( .A(x[4029]), .B(y[4029]), .Z(n25495) );
  NANDN U17475 ( .A(x[4030]), .B(y[4030]), .Z(n25492) );
  AND U17476 ( .A(n25495), .B(n25492), .Z(n56275) );
  NANDN U17477 ( .A(y[4028]), .B(x[4028]), .Z(n9827) );
  NANDN U17478 ( .A(y[4029]), .B(x[4029]), .Z(n25494) );
  NAND U17479 ( .A(n9827), .B(n25494), .Z(n56274) );
  XNOR U17480 ( .A(x[4028]), .B(y[4028]), .Z(n25497) );
  NANDN U17481 ( .A(x[4027]), .B(y[4027]), .Z(n56273) );
  NANDN U17482 ( .A(y[4026]), .B(x[4026]), .Z(n40163) );
  NANDN U17483 ( .A(y[4027]), .B(x[4027]), .Z(n25496) );
  AND U17484 ( .A(n40163), .B(n25496), .Z(n56270) );
  NANDN U17485 ( .A(x[4025]), .B(y[4025]), .Z(n25499) );
  NANDN U17486 ( .A(x[4026]), .B(y[4026]), .Z(n25498) );
  AND U17487 ( .A(n25499), .B(n25498), .Z(n51733) );
  NANDN U17488 ( .A(y[4024]), .B(x[4024]), .Z(n40157) );
  NANDN U17489 ( .A(y[4025]), .B(x[4025]), .Z(n40164) );
  NAND U17490 ( .A(n40157), .B(n40164), .Z(n51734) );
  NANDN U17491 ( .A(x[4023]), .B(y[4023]), .Z(n25501) );
  NANDN U17492 ( .A(x[4024]), .B(y[4024]), .Z(n25500) );
  AND U17493 ( .A(n25501), .B(n25500), .Z(n56267) );
  NANDN U17494 ( .A(y[4020]), .B(x[4020]), .Z(n40145) );
  NANDN U17495 ( .A(y[4021]), .B(x[4021]), .Z(n40152) );
  NAND U17496 ( .A(n40145), .B(n40152), .Z(n51736) );
  NANDN U17497 ( .A(y[4018]), .B(x[4018]), .Z(n40139) );
  NANDN U17498 ( .A(y[4019]), .B(x[4019]), .Z(n40146) );
  AND U17499 ( .A(n40139), .B(n40146), .Z(n56264) );
  NANDN U17500 ( .A(x[4017]), .B(y[4017]), .Z(n25507) );
  NANDN U17501 ( .A(x[4018]), .B(y[4018]), .Z(n25506) );
  NAND U17502 ( .A(n25507), .B(n25506), .Z(n56263) );
  NANDN U17503 ( .A(y[4016]), .B(x[4016]), .Z(n40133) );
  NANDN U17504 ( .A(y[4017]), .B(x[4017]), .Z(n40140) );
  AND U17505 ( .A(n40133), .B(n40140), .Z(n56262) );
  NANDN U17506 ( .A(x[4015]), .B(y[4015]), .Z(n25509) );
  NANDN U17507 ( .A(x[4016]), .B(y[4016]), .Z(n25508) );
  AND U17508 ( .A(n25509), .B(n25508), .Z(n51737) );
  NANDN U17509 ( .A(y[4014]), .B(x[4014]), .Z(n9828) );
  NANDN U17510 ( .A(y[4015]), .B(x[4015]), .Z(n40134) );
  NAND U17511 ( .A(n9828), .B(n40134), .Z(n51738) );
  XNOR U17512 ( .A(y[4014]), .B(x[4014]), .Z(n40128) );
  NANDN U17513 ( .A(x[4013]), .B(y[4013]), .Z(n40123) );
  AND U17514 ( .A(n40128), .B(n40123), .Z(n56259) );
  XNOR U17515 ( .A(y[4012]), .B(x[4012]), .Z(n9829) );
  ANDN U17516 ( .B(y[4011]), .A(x[4011]), .Z(n40118) );
  ANDN U17517 ( .B(n9829), .A(n40118), .Z(n56257) );
  NANDN U17518 ( .A(y[4010]), .B(x[4010]), .Z(n25513) );
  NANDN U17519 ( .A(y[4011]), .B(x[4011]), .Z(n25512) );
  NAND U17520 ( .A(n25513), .B(n25512), .Z(n56256) );
  NANDN U17521 ( .A(x[4009]), .B(y[4009]), .Z(n40112) );
  ANDN U17522 ( .B(y[4010]), .A(x[4010]), .Z(n40119) );
  ANDN U17523 ( .B(n40112), .A(n40119), .Z(n56255) );
  NANDN U17524 ( .A(y[4004]), .B(x[4004]), .Z(n25521) );
  NANDN U17525 ( .A(y[4005]), .B(x[4005]), .Z(n25518) );
  NAND U17526 ( .A(n25521), .B(n25518), .Z(n51740) );
  NANDN U17527 ( .A(x[4003]), .B(y[4003]), .Z(n40096) );
  NANDN U17528 ( .A(x[4004]), .B(y[4004]), .Z(n25520) );
  AND U17529 ( .A(n40096), .B(n25520), .Z(n56251) );
  XNOR U17530 ( .A(x[4002]), .B(y[4002]), .Z(n25524) );
  NANDN U17531 ( .A(x[4001]), .B(y[4001]), .Z(n56245) );
  AND U17532 ( .A(n25524), .B(n56245), .Z(n15777) );
  XNOR U17533 ( .A(x[3998]), .B(y[3998]), .Z(n25526) );
  NANDN U17534 ( .A(y[3996]), .B(x[3996]), .Z(n25528) );
  NANDN U17535 ( .A(y[3997]), .B(x[3997]), .Z(n25525) );
  NAND U17536 ( .A(n25528), .B(n25525), .Z(n56240) );
  NANDN U17537 ( .A(x[3995]), .B(y[3995]), .Z(n25530) );
  NANDN U17538 ( .A(x[3996]), .B(y[3996]), .Z(n25527) );
  AND U17539 ( .A(n25530), .B(n25527), .Z(n56239) );
  NANDN U17540 ( .A(y[3994]), .B(x[3994]), .Z(n9830) );
  NANDN U17541 ( .A(y[3995]), .B(x[3995]), .Z(n25529) );
  NAND U17542 ( .A(n9830), .B(n25529), .Z(n56238) );
  NANDN U17543 ( .A(x[3993]), .B(y[3993]), .Z(n51743) );
  XNOR U17544 ( .A(x[3994]), .B(y[3994]), .Z(n40075) );
  AND U17545 ( .A(n51743), .B(n40075), .Z(n15764) );
  NANDN U17546 ( .A(y[3992]), .B(x[3992]), .Z(n9831) );
  NANDN U17547 ( .A(y[3993]), .B(x[3993]), .Z(n40074) );
  NAND U17548 ( .A(n9831), .B(n40074), .Z(n56237) );
  XNOR U17549 ( .A(x[3992]), .B(y[3992]), .Z(n25532) );
  NANDN U17550 ( .A(y[3990]), .B(x[3990]), .Z(n25533) );
  NANDN U17551 ( .A(y[3991]), .B(x[3991]), .Z(n25531) );
  NAND U17552 ( .A(n25533), .B(n25531), .Z(n56234) );
  NANDN U17553 ( .A(x[3989]), .B(y[3989]), .Z(n25535) );
  NANDN U17554 ( .A(x[3990]), .B(y[3990]), .Z(n40067) );
  AND U17555 ( .A(n25535), .B(n40067), .Z(n56233) );
  NANDN U17556 ( .A(y[3988]), .B(x[3988]), .Z(n9832) );
  NANDN U17557 ( .A(y[3989]), .B(x[3989]), .Z(n25534) );
  NAND U17558 ( .A(n9832), .B(n25534), .Z(n56232) );
  XNOR U17559 ( .A(x[3988]), .B(y[3988]), .Z(n25537) );
  NANDN U17560 ( .A(x[3985]), .B(y[3985]), .Z(n40054) );
  ANDN U17561 ( .B(y[3986]), .A(x[3986]), .Z(n40060) );
  ANDN U17562 ( .B(n40054), .A(n40060), .Z(n56229) );
  XNOR U17563 ( .A(x[3984]), .B(y[3984]), .Z(n25541) );
  NANDN U17564 ( .A(y[3982]), .B(x[3982]), .Z(n40046) );
  NANDN U17565 ( .A(y[3983]), .B(x[3983]), .Z(n25540) );
  NAND U17566 ( .A(n40046), .B(n25540), .Z(n56225) );
  NANDN U17567 ( .A(x[3981]), .B(y[3981]), .Z(n25543) );
  NANDN U17568 ( .A(x[3982]), .B(y[3982]), .Z(n25542) );
  AND U17569 ( .A(n25543), .B(n25542), .Z(n51747) );
  NANDN U17570 ( .A(y[3978]), .B(x[3978]), .Z(n40034) );
  NANDN U17571 ( .A(y[3979]), .B(x[3979]), .Z(n40041) );
  NAND U17572 ( .A(n40034), .B(n40041), .Z(n56223) );
  NANDN U17573 ( .A(y[3976]), .B(x[3976]), .Z(n40028) );
  NANDN U17574 ( .A(y[3977]), .B(x[3977]), .Z(n40035) );
  AND U17575 ( .A(n40028), .B(n40035), .Z(n56220) );
  ANDN U17576 ( .B(y[3975]), .A(x[3975]), .Z(n40026) );
  XNOR U17577 ( .A(x[3976]), .B(y[3976]), .Z(n9833) );
  NANDN U17578 ( .A(n40026), .B(n9833), .Z(n56219) );
  NANDN U17579 ( .A(y[3974]), .B(x[3974]), .Z(n9834) );
  NANDN U17580 ( .A(y[3975]), .B(x[3975]), .Z(n40029) );
  AND U17581 ( .A(n9834), .B(n40029), .Z(n51750) );
  XNOR U17582 ( .A(y[3970]), .B(x[3970]), .Z(n40012) );
  NANDN U17583 ( .A(x[3969]), .B(y[3969]), .Z(n40007) );
  AND U17584 ( .A(n40012), .B(n40007), .Z(n56215) );
  NANDN U17585 ( .A(x[3967]), .B(y[3967]), .Z(n25557) );
  NANDN U17586 ( .A(x[3968]), .B(y[3968]), .Z(n40008) );
  AND U17587 ( .A(n25557), .B(n40008), .Z(n56213) );
  NANDN U17588 ( .A(y[3966]), .B(x[3966]), .Z(n25559) );
  NANDN U17589 ( .A(y[3967]), .B(x[3967]), .Z(n40006) );
  NAND U17590 ( .A(n25559), .B(n40006), .Z(n56212) );
  NANDN U17591 ( .A(x[3965]), .B(y[3965]), .Z(n39997) );
  NANDN U17592 ( .A(x[3966]), .B(y[3966]), .Z(n25558) );
  AND U17593 ( .A(n39997), .B(n25558), .Z(n56211) );
  NANDN U17594 ( .A(y[3964]), .B(x[3964]), .Z(n9835) );
  NANDN U17595 ( .A(y[3965]), .B(x[3965]), .Z(n25560) );
  NAND U17596 ( .A(n9835), .B(n25560), .Z(n56210) );
  NANDN U17597 ( .A(x[3963]), .B(y[3963]), .Z(n56206) );
  XNOR U17598 ( .A(x[3964]), .B(y[3964]), .Z(n25562) );
  AND U17599 ( .A(n56206), .B(n25562), .Z(n15726) );
  NANDN U17600 ( .A(y[3962]), .B(x[3962]), .Z(n25563) );
  NANDN U17601 ( .A(y[3963]), .B(x[3963]), .Z(n25561) );
  NAND U17602 ( .A(n25563), .B(n25561), .Z(n56205) );
  NANDN U17603 ( .A(x[3961]), .B(y[3961]), .Z(n25565) );
  NANDN U17604 ( .A(x[3962]), .B(y[3962]), .Z(n39992) );
  AND U17605 ( .A(n25565), .B(n39992), .Z(n56204) );
  NANDN U17606 ( .A(y[3960]), .B(x[3960]), .Z(n25567) );
  NANDN U17607 ( .A(y[3961]), .B(x[3961]), .Z(n25564) );
  NAND U17608 ( .A(n25567), .B(n25564), .Z(n56203) );
  NANDN U17609 ( .A(x[3959]), .B(y[3959]), .Z(n39982) );
  NANDN U17610 ( .A(x[3960]), .B(y[3960]), .Z(n25566) );
  AND U17611 ( .A(n39982), .B(n25566), .Z(n56202) );
  NANDN U17612 ( .A(y[3958]), .B(x[3958]), .Z(n9836) );
  NANDN U17613 ( .A(y[3959]), .B(x[3959]), .Z(n25568) );
  NAND U17614 ( .A(n9836), .B(n25568), .Z(n56201) );
  NANDN U17615 ( .A(x[3957]), .B(y[3957]), .Z(n56199) );
  XNOR U17616 ( .A(x[3958]), .B(y[3958]), .Z(n39980) );
  AND U17617 ( .A(n56199), .B(n39980), .Z(n15719) );
  ANDN U17618 ( .B(x[3957]), .A(y[3957]), .Z(n39979) );
  NANDN U17619 ( .A(y[3956]), .B(x[3956]), .Z(n39973) );
  NANDN U17620 ( .A(n39979), .B(n39973), .Z(n56198) );
  NANDN U17621 ( .A(x[3955]), .B(y[3955]), .Z(n25570) );
  NANDN U17622 ( .A(x[3956]), .B(y[3956]), .Z(n25569) );
  AND U17623 ( .A(n25570), .B(n25569), .Z(n56197) );
  NANDN U17624 ( .A(y[3954]), .B(x[3954]), .Z(n39968) );
  NANDN U17625 ( .A(y[3955]), .B(x[3955]), .Z(n39974) );
  NAND U17626 ( .A(n39968), .B(n39974), .Z(n56196) );
  NANDN U17627 ( .A(y[3952]), .B(x[3952]), .Z(n9837) );
  NANDN U17628 ( .A(y[3953]), .B(x[3953]), .Z(n51752) );
  AND U17629 ( .A(n9837), .B(n51752), .Z(n56195) );
  IV U17630 ( .A(x[3952]), .Z(n9838) );
  XOR U17631 ( .A(n9838), .B(y[3952]), .Z(n15711) );
  ANDN U17632 ( .B(y[3951]), .A(x[3951]), .Z(n25574) );
  NANDN U17633 ( .A(x[3949]), .B(y[3949]), .Z(n25578) );
  NANDN U17634 ( .A(x[3950]), .B(y[3950]), .Z(n25575) );
  NAND U17635 ( .A(n25578), .B(n25575), .Z(n51756) );
  NANDN U17636 ( .A(y[3948]), .B(x[3948]), .Z(n25580) );
  NANDN U17637 ( .A(y[3949]), .B(x[3949]), .Z(n25577) );
  AND U17638 ( .A(n25580), .B(n25577), .Z(n56192) );
  ANDN U17639 ( .B(y[3945]), .A(x[3945]), .Z(n39947) );
  XNOR U17640 ( .A(x[3946]), .B(y[3946]), .Z(n9839) );
  NANDN U17641 ( .A(n39947), .B(n9839), .Z(n51758) );
  NANDN U17642 ( .A(y[3944]), .B(x[3944]), .Z(n9840) );
  NANDN U17643 ( .A(y[3945]), .B(x[3945]), .Z(n25583) );
  AND U17644 ( .A(n9840), .B(n25583), .Z(n56190) );
  XNOR U17645 ( .A(y[3944]), .B(x[3944]), .Z(n25585) );
  NANDN U17646 ( .A(x[3943]), .B(y[3943]), .Z(n25586) );
  NAND U17647 ( .A(n25585), .B(n25586), .Z(n56189) );
  NANDN U17648 ( .A(y[3942]), .B(x[3942]), .Z(n25588) );
  NANDN U17649 ( .A(y[3943]), .B(x[3943]), .Z(n25584) );
  AND U17650 ( .A(n25588), .B(n25584), .Z(n56188) );
  NANDN U17651 ( .A(x[3941]), .B(y[3941]), .Z(n39937) );
  NANDN U17652 ( .A(x[3942]), .B(y[3942]), .Z(n25587) );
  NAND U17653 ( .A(n39937), .B(n25587), .Z(n56187) );
  NANDN U17654 ( .A(y[3938]), .B(x[3938]), .Z(n25592) );
  NANDN U17655 ( .A(y[3939]), .B(x[3939]), .Z(n25591) );
  NAND U17656 ( .A(n25592), .B(n25591), .Z(n56184) );
  NANDN U17657 ( .A(x[3937]), .B(y[3937]), .Z(n25594) );
  NANDN U17658 ( .A(x[3938]), .B(y[3938]), .Z(n39932) );
  AND U17659 ( .A(n25594), .B(n39932), .Z(n51759) );
  XNOR U17660 ( .A(x[3934]), .B(y[3934]), .Z(n39918) );
  NANDN U17661 ( .A(y[3932]), .B(x[3932]), .Z(n9841) );
  NANDN U17662 ( .A(y[3933]), .B(x[3933]), .Z(n39917) );
  NAND U17663 ( .A(n9841), .B(n39917), .Z(n56177) );
  NANDN U17664 ( .A(x[3931]), .B(y[3931]), .Z(n51761) );
  XNOR U17665 ( .A(x[3932]), .B(y[3932]), .Z(n39913) );
  ANDN U17666 ( .B(x[3931]), .A(y[3931]), .Z(n39912) );
  NANDN U17667 ( .A(y[3930]), .B(x[3930]), .Z(n25600) );
  NANDN U17668 ( .A(n39912), .B(n25600), .Z(n56176) );
  NANDN U17669 ( .A(x[3929]), .B(y[3929]), .Z(n25601) );
  NANDN U17670 ( .A(x[3930]), .B(y[3930]), .Z(n25598) );
  AND U17671 ( .A(n25601), .B(n25598), .Z(n56175) );
  NANDN U17672 ( .A(y[3926]), .B(x[3926]), .Z(n25605) );
  NANDN U17673 ( .A(y[3927]), .B(x[3927]), .Z(n25604) );
  NAND U17674 ( .A(n25605), .B(n25604), .Z(n56171) );
  NANDN U17675 ( .A(x[3925]), .B(y[3925]), .Z(n39893) );
  NANDN U17676 ( .A(x[3926]), .B(y[3926]), .Z(n39900) );
  AND U17677 ( .A(n39893), .B(n39900), .Z(n51763) );
  NANDN U17678 ( .A(y[3920]), .B(x[3920]), .Z(n39878) );
  NANDN U17679 ( .A(y[3921]), .B(x[3921]), .Z(n25610) );
  NAND U17680 ( .A(n39878), .B(n25610), .Z(n56166) );
  NANDN U17681 ( .A(x[3919]), .B(y[3919]), .Z(n25611) );
  NANDN U17682 ( .A(x[3920]), .B(y[3920]), .Z(n39882) );
  AND U17683 ( .A(n25611), .B(n39882), .Z(n56165) );
  NANDN U17684 ( .A(y[3918]), .B(x[3918]), .Z(n39872) );
  NANDN U17685 ( .A(y[3919]), .B(x[3919]), .Z(n39879) );
  NAND U17686 ( .A(n39872), .B(n39879), .Z(n56164) );
  NANDN U17687 ( .A(x[3917]), .B(y[3917]), .Z(n25613) );
  NANDN U17688 ( .A(x[3918]), .B(y[3918]), .Z(n25612) );
  AND U17689 ( .A(n25613), .B(n25612), .Z(n56163) );
  NANDN U17690 ( .A(y[3916]), .B(x[3916]), .Z(n39866) );
  NANDN U17691 ( .A(y[3917]), .B(x[3917]), .Z(n39873) );
  NAND U17692 ( .A(n39866), .B(n39873), .Z(n56162) );
  NANDN U17693 ( .A(x[3913]), .B(y[3913]), .Z(n25619) );
  NANDN U17694 ( .A(x[3914]), .B(y[3914]), .Z(n25616) );
  NAND U17695 ( .A(n25619), .B(n25616), .Z(n56159) );
  NANDN U17696 ( .A(y[3912]), .B(x[3912]), .Z(n39858) );
  NANDN U17697 ( .A(y[3913]), .B(x[3913]), .Z(n25618) );
  AND U17698 ( .A(n39858), .B(n25618), .Z(n51766) );
  NANDN U17699 ( .A(y[3910]), .B(x[3910]), .Z(n39849) );
  ANDN U17700 ( .B(x[3911]), .A(y[3911]), .Z(n39856) );
  ANDN U17701 ( .B(n39849), .A(n39856), .Z(n56156) );
  NANDN U17702 ( .A(x[3907]), .B(y[3907]), .Z(n25625) );
  XNOR U17703 ( .A(x[3908]), .B(y[3908]), .Z(n9842) );
  NAND U17704 ( .A(n25625), .B(n9842), .Z(n51769) );
  NANDN U17705 ( .A(y[3906]), .B(x[3906]), .Z(n39837) );
  NANDN U17706 ( .A(y[3907]), .B(x[3907]), .Z(n39844) );
  AND U17707 ( .A(n39837), .B(n39844), .Z(n56154) );
  NANDN U17708 ( .A(x[3905]), .B(y[3905]), .Z(n25627) );
  NANDN U17709 ( .A(x[3906]), .B(y[3906]), .Z(n25626) );
  NAND U17710 ( .A(n25627), .B(n25626), .Z(n56153) );
  NANDN U17711 ( .A(y[3904]), .B(x[3904]), .Z(n9843) );
  NANDN U17712 ( .A(y[3905]), .B(x[3905]), .Z(n39838) );
  AND U17713 ( .A(n9843), .B(n39838), .Z(n56152) );
  XNOR U17714 ( .A(y[3904]), .B(x[3904]), .Z(n39832) );
  NANDN U17715 ( .A(x[3903]), .B(y[3903]), .Z(n25629) );
  NAND U17716 ( .A(n39832), .B(n25629), .Z(n56151) );
  NANDN U17717 ( .A(y[3902]), .B(x[3902]), .Z(n9844) );
  NANDN U17718 ( .A(y[3903]), .B(x[3903]), .Z(n39831) );
  AND U17719 ( .A(n9844), .B(n39831), .Z(n56150) );
  XNOR U17720 ( .A(y[3902]), .B(x[3902]), .Z(n39826) );
  NANDN U17721 ( .A(x[3901]), .B(y[3901]), .Z(n39821) );
  NAND U17722 ( .A(n39826), .B(n39821), .Z(n56149) );
  NANDN U17723 ( .A(y[3900]), .B(x[3900]), .Z(n39818) );
  NANDN U17724 ( .A(y[3901]), .B(x[3901]), .Z(n39825) );
  AND U17725 ( .A(n39818), .B(n39825), .Z(n56148) );
  NANDN U17726 ( .A(x[3897]), .B(y[3897]), .Z(n39810) );
  XNOR U17727 ( .A(x[3898]), .B(y[3898]), .Z(n9845) );
  NAND U17728 ( .A(n39810), .B(n9845), .Z(n51771) );
  NANDN U17729 ( .A(y[3896]), .B(x[3896]), .Z(n25635) );
  NANDN U17730 ( .A(y[3897]), .B(x[3897]), .Z(n25634) );
  AND U17731 ( .A(n25635), .B(n25634), .Z(n56145) );
  ANDN U17732 ( .B(y[3893]), .A(x[3893]), .Z(n39798) );
  NANDN U17733 ( .A(x[3894]), .B(y[3894]), .Z(n39805) );
  NANDN U17734 ( .A(n39798), .B(n39805), .Z(n56142) );
  NANDN U17735 ( .A(x[3891]), .B(y[3891]), .Z(n25641) );
  ANDN U17736 ( .B(y[3892]), .A(x[3892]), .Z(n39799) );
  ANDN U17737 ( .B(n25641), .A(n39799), .Z(n56141) );
  NANDN U17738 ( .A(y[3890]), .B(x[3890]), .Z(n25643) );
  NANDN U17739 ( .A(y[3891]), .B(x[3891]), .Z(n25640) );
  NAND U17740 ( .A(n25643), .B(n25640), .Z(n56140) );
  NANDN U17741 ( .A(x[3889]), .B(y[3889]), .Z(n39788) );
  NANDN U17742 ( .A(x[3890]), .B(y[3890]), .Z(n25642) );
  AND U17743 ( .A(n39788), .B(n25642), .Z(n56139) );
  NANDN U17744 ( .A(y[3888]), .B(x[3888]), .Z(n9846) );
  NANDN U17745 ( .A(y[3889]), .B(x[3889]), .Z(n25644) );
  NAND U17746 ( .A(n9846), .B(n25644), .Z(n56138) );
  XNOR U17747 ( .A(x[3888]), .B(y[3888]), .Z(n39785) );
  NANDN U17748 ( .A(x[3887]), .B(y[3887]), .Z(n56136) );
  AND U17749 ( .A(n39785), .B(n56136), .Z(n15640) );
  NANDN U17750 ( .A(x[3885]), .B(y[3885]), .Z(n25648) );
  NANDN U17751 ( .A(x[3886]), .B(y[3886]), .Z(n25645) );
  AND U17752 ( .A(n25648), .B(n25645), .Z(n56134) );
  NANDN U17753 ( .A(y[3884]), .B(x[3884]), .Z(n25650) );
  NANDN U17754 ( .A(y[3885]), .B(x[3885]), .Z(n25646) );
  NAND U17755 ( .A(n25650), .B(n25646), .Z(n56132) );
  NANDN U17756 ( .A(x[3883]), .B(y[3883]), .Z(n25652) );
  NANDN U17757 ( .A(x[3884]), .B(y[3884]), .Z(n25649) );
  AND U17758 ( .A(n25652), .B(n25649), .Z(n56131) );
  NANDN U17759 ( .A(y[3882]), .B(x[3882]), .Z(n9847) );
  NANDN U17760 ( .A(y[3883]), .B(x[3883]), .Z(n25651) );
  NAND U17761 ( .A(n9847), .B(n25651), .Z(n56130) );
  NANDN U17762 ( .A(y[3880]), .B(x[3880]), .Z(n9848) );
  NANDN U17763 ( .A(y[3881]), .B(x[3881]), .Z(n39772) );
  AND U17764 ( .A(n9848), .B(n39772), .Z(n51773) );
  XNOR U17765 ( .A(x[3880]), .B(y[3880]), .Z(n39765) );
  NANDN U17766 ( .A(y[3878]), .B(x[3878]), .Z(n9849) );
  NANDN U17767 ( .A(y[3879]), .B(x[3879]), .Z(n39766) );
  AND U17768 ( .A(n9849), .B(n39766), .Z(n56125) );
  ANDN U17769 ( .B(y[3877]), .A(x[3877]), .Z(n25655) );
  XNOR U17770 ( .A(x[3878]), .B(y[3878]), .Z(n25654) );
  NANDN U17771 ( .A(y[3876]), .B(x[3876]), .Z(n25657) );
  NANDN U17772 ( .A(y[3877]), .B(x[3877]), .Z(n25653) );
  NAND U17773 ( .A(n25657), .B(n25653), .Z(n56124) );
  NANDN U17774 ( .A(x[3875]), .B(y[3875]), .Z(n25659) );
  NANDN U17775 ( .A(x[3876]), .B(y[3876]), .Z(n25656) );
  AND U17776 ( .A(n25659), .B(n25656), .Z(n56123) );
  NANDN U17777 ( .A(y[3874]), .B(x[3874]), .Z(n9850) );
  NANDN U17778 ( .A(y[3875]), .B(x[3875]), .Z(n25658) );
  NAND U17779 ( .A(n9850), .B(n25658), .Z(n56122) );
  XNOR U17780 ( .A(x[3874]), .B(y[3874]), .Z(n39751) );
  NANDN U17781 ( .A(y[3870]), .B(x[3870]), .Z(n25662) );
  NANDN U17782 ( .A(y[3871]), .B(x[3871]), .Z(n39746) );
  NAND U17783 ( .A(n25662), .B(n39746), .Z(n51777) );
  NANDN U17784 ( .A(x[3869]), .B(y[3869]), .Z(n39736) );
  NANDN U17785 ( .A(x[3870]), .B(y[3870]), .Z(n25661) );
  AND U17786 ( .A(n39736), .B(n25661), .Z(n56116) );
  NANDN U17787 ( .A(x[3867]), .B(y[3867]), .Z(n39730) );
  ANDN U17788 ( .B(y[3868]), .A(x[3868]), .Z(n39738) );
  ANDN U17789 ( .B(n39730), .A(n39738), .Z(n56114) );
  NANDN U17790 ( .A(y[3866]), .B(x[3866]), .Z(n25666) );
  NANDN U17791 ( .A(y[3867]), .B(x[3867]), .Z(n25665) );
  NAND U17792 ( .A(n25666), .B(n25665), .Z(n56113) );
  NANDN U17793 ( .A(y[3864]), .B(x[3864]), .Z(n25670) );
  NANDN U17794 ( .A(y[3865]), .B(x[3865]), .Z(n25667) );
  AND U17795 ( .A(n25670), .B(n25667), .Z(n56112) );
  NANDN U17796 ( .A(x[3863]), .B(y[3863]), .Z(n39720) );
  NANDN U17797 ( .A(x[3864]), .B(y[3864]), .Z(n25669) );
  NAND U17798 ( .A(n39720), .B(n25669), .Z(n56111) );
  NANDN U17799 ( .A(y[3862]), .B(x[3862]), .Z(n9851) );
  NANDN U17800 ( .A(y[3863]), .B(x[3863]), .Z(n25671) );
  AND U17801 ( .A(n9851), .B(n25671), .Z(n56110) );
  XNOR U17802 ( .A(y[3862]), .B(x[3862]), .Z(n39716) );
  NANDN U17803 ( .A(x[3861]), .B(y[3861]), .Z(n25672) );
  NAND U17804 ( .A(n39716), .B(n25672), .Z(n56109) );
  NANDN U17805 ( .A(y[3860]), .B(x[3860]), .Z(n39710) );
  NANDN U17806 ( .A(y[3861]), .B(x[3861]), .Z(n39717) );
  AND U17807 ( .A(n39710), .B(n39717), .Z(n56108) );
  NANDN U17808 ( .A(x[3857]), .B(y[3857]), .Z(n25676) );
  NANDN U17809 ( .A(x[3858]), .B(y[3858]), .Z(n25675) );
  NAND U17810 ( .A(n25676), .B(n25675), .Z(n51780) );
  NANDN U17811 ( .A(y[3856]), .B(x[3856]), .Z(n39698) );
  NANDN U17812 ( .A(y[3857]), .B(x[3857]), .Z(n39705) );
  AND U17813 ( .A(n39698), .B(n39705), .Z(n56105) );
  ANDN U17814 ( .B(y[3853]), .A(x[3853]), .Z(n25680) );
  XNOR U17815 ( .A(x[3854]), .B(y[3854]), .Z(n25679) );
  NANDN U17816 ( .A(y[3852]), .B(x[3852]), .Z(n25682) );
  NANDN U17817 ( .A(y[3853]), .B(x[3853]), .Z(n25678) );
  AND U17818 ( .A(n25682), .B(n25678), .Z(n56100) );
  NANDN U17819 ( .A(x[3851]), .B(y[3851]), .Z(n25685) );
  NANDN U17820 ( .A(x[3852]), .B(y[3852]), .Z(n25681) );
  NAND U17821 ( .A(n25685), .B(n25681), .Z(n51781) );
  NANDN U17822 ( .A(y[3850]), .B(x[3850]), .Z(n39683) );
  NANDN U17823 ( .A(y[3851]), .B(x[3851]), .Z(n25683) );
  AND U17824 ( .A(n39683), .B(n25683), .Z(n56099) );
  NANDN U17825 ( .A(y[3848]), .B(x[3848]), .Z(n25686) );
  ANDN U17826 ( .B(x[3849]), .A(y[3849]), .Z(n39685) );
  ANDN U17827 ( .B(n25686), .A(n39685), .Z(n56097) );
  NANDN U17828 ( .A(x[3845]), .B(y[3845]), .Z(n25690) );
  NANDN U17829 ( .A(x[3846]), .B(y[3846]), .Z(n39674) );
  NAND U17830 ( .A(n25690), .B(n39674), .Z(n51783) );
  NANDN U17831 ( .A(y[3844]), .B(x[3844]), .Z(n25692) );
  NANDN U17832 ( .A(y[3845]), .B(x[3845]), .Z(n25689) );
  AND U17833 ( .A(n25692), .B(n25689), .Z(n56093) );
  NANDN U17834 ( .A(y[3842]), .B(x[3842]), .Z(n9852) );
  NANDN U17835 ( .A(y[3843]), .B(x[3843]), .Z(n25693) );
  AND U17836 ( .A(n9852), .B(n25693), .Z(n51784) );
  XNOR U17837 ( .A(x[3842]), .B(y[3842]), .Z(n39660) );
  NANDN U17838 ( .A(y[3840]), .B(x[3840]), .Z(n9853) );
  NANDN U17839 ( .A(y[3841]), .B(x[3841]), .Z(n39659) );
  NAND U17840 ( .A(n9853), .B(n39659), .Z(n56089) );
  NANDN U17841 ( .A(x[3839]), .B(y[3839]), .Z(n56088) );
  XNOR U17842 ( .A(x[3840]), .B(y[3840]), .Z(n39654) );
  NANDN U17843 ( .A(y[3838]), .B(x[3838]), .Z(n39648) );
  NANDN U17844 ( .A(y[3839]), .B(x[3839]), .Z(n39655) );
  AND U17845 ( .A(n39648), .B(n39655), .Z(n56086) );
  NANDN U17846 ( .A(x[3837]), .B(y[3837]), .Z(n25695) );
  NANDN U17847 ( .A(x[3838]), .B(y[3838]), .Z(n25694) );
  NAND U17848 ( .A(n25695), .B(n25694), .Z(n56085) );
  NANDN U17849 ( .A(y[3836]), .B(x[3836]), .Z(n9854) );
  NANDN U17850 ( .A(y[3837]), .B(x[3837]), .Z(n39649) );
  AND U17851 ( .A(n9854), .B(n39649), .Z(n56084) );
  NANDN U17852 ( .A(x[3835]), .B(y[3835]), .Z(n56080) );
  XNOR U17853 ( .A(x[3836]), .B(y[3836]), .Z(n39642) );
  NANDN U17854 ( .A(y[3834]), .B(x[3834]), .Z(n9855) );
  NANDN U17855 ( .A(y[3835]), .B(x[3835]), .Z(n39643) );
  NAND U17856 ( .A(n9855), .B(n39643), .Z(n56079) );
  NANDN U17857 ( .A(x[3833]), .B(y[3833]), .Z(n51786) );
  XNOR U17858 ( .A(x[3834]), .B(y[3834]), .Z(n25697) );
  XNOR U17859 ( .A(x[3832]), .B(y[3832]), .Z(n25699) );
  NANDN U17860 ( .A(x[3831]), .B(y[3831]), .Z(n51787) );
  AND U17861 ( .A(n25699), .B(n51787), .Z(n15572) );
  NANDN U17862 ( .A(x[3829]), .B(y[3829]), .Z(n25701) );
  NANDN U17863 ( .A(x[3830]), .B(y[3830]), .Z(n25700) );
  NAND U17864 ( .A(n25701), .B(n25700), .Z(n56076) );
  NANDN U17865 ( .A(y[3828]), .B(x[3828]), .Z(n9856) );
  NANDN U17866 ( .A(y[3829]), .B(x[3829]), .Z(n39628) );
  AND U17867 ( .A(n9856), .B(n39628), .Z(n51789) );
  XNOR U17868 ( .A(y[3826]), .B(x[3826]), .Z(n39616) );
  NANDN U17869 ( .A(x[3825]), .B(y[3825]), .Z(n25705) );
  NAND U17870 ( .A(n39616), .B(n25705), .Z(n56072) );
  NANDN U17871 ( .A(y[3824]), .B(x[3824]), .Z(n9857) );
  NANDN U17872 ( .A(y[3825]), .B(x[3825]), .Z(n39615) );
  AND U17873 ( .A(n9857), .B(n39615), .Z(n56071) );
  XNOR U17874 ( .A(y[3820]), .B(x[3820]), .Z(n25712) );
  NANDN U17875 ( .A(x[3819]), .B(y[3819]), .Z(n39596) );
  NAND U17876 ( .A(n25712), .B(n39596), .Z(n56068) );
  NANDN U17877 ( .A(y[3818]), .B(x[3818]), .Z(n9858) );
  NANDN U17878 ( .A(y[3819]), .B(x[3819]), .Z(n25711) );
  AND U17879 ( .A(n9858), .B(n25711), .Z(n51793) );
  NANDN U17880 ( .A(y[3817]), .B(x[3817]), .Z(n25713) );
  ANDN U17881 ( .B(x[3816]), .A(y[3816]), .Z(n39586) );
  ANDN U17882 ( .B(n25713), .A(n39586), .Z(n56066) );
  NANDN U17883 ( .A(x[3815]), .B(y[3815]), .Z(n39582) );
  NANDN U17884 ( .A(x[3816]), .B(y[3816]), .Z(n39591) );
  NAND U17885 ( .A(n39582), .B(n39591), .Z(n56065) );
  NANDN U17886 ( .A(y[3812]), .B(x[3812]), .Z(n25717) );
  NANDN U17887 ( .A(y[3813]), .B(x[3813]), .Z(n25716) );
  NAND U17888 ( .A(n25717), .B(n25716), .Z(n56060) );
  NANDN U17889 ( .A(x[3811]), .B(y[3811]), .Z(n39569) );
  NANDN U17890 ( .A(x[3812]), .B(y[3812]), .Z(n39576) );
  AND U17891 ( .A(n39569), .B(n39576), .Z(n56059) );
  NANDN U17892 ( .A(y[3806]), .B(x[3806]), .Z(n39553) );
  NANDN U17893 ( .A(y[3807]), .B(x[3807]), .Z(n25722) );
  NAND U17894 ( .A(n39553), .B(n25722), .Z(n56056) );
  NANDN U17895 ( .A(x[3805]), .B(y[3805]), .Z(n39550) );
  NANDN U17896 ( .A(x[3806]), .B(y[3806]), .Z(n39558) );
  AND U17897 ( .A(n39550), .B(n39558), .Z(n51796) );
  NANDN U17898 ( .A(x[3803]), .B(y[3803]), .Z(n25725) );
  NANDN U17899 ( .A(x[3804]), .B(y[3804]), .Z(n39552) );
  AND U17900 ( .A(n25725), .B(n39552), .Z(n56054) );
  ANDN U17901 ( .B(x[3802]), .A(y[3802]), .Z(n39543) );
  NANDN U17902 ( .A(y[3803]), .B(x[3803]), .Z(n25724) );
  NANDN U17903 ( .A(n39543), .B(n25724), .Z(n56053) );
  NANDN U17904 ( .A(x[3802]), .B(y[3802]), .Z(n56049) );
  ANDN U17905 ( .B(x[3801]), .A(y[3801]), .Z(n56050) );
  NANDN U17906 ( .A(y[3800]), .B(x[3800]), .Z(n25728) );
  NANDN U17907 ( .A(n56050), .B(n25728), .Z(n56048) );
  NANDN U17908 ( .A(y[3798]), .B(x[3798]), .Z(n9859) );
  NANDN U17909 ( .A(y[3799]), .B(x[3799]), .Z(n25729) );
  AND U17910 ( .A(n9859), .B(n25729), .Z(n56046) );
  NANDN U17911 ( .A(x[3797]), .B(y[3797]), .Z(n51798) );
  XNOR U17912 ( .A(x[3798]), .B(y[3798]), .Z(n25731) );
  AND U17913 ( .A(n51798), .B(n25731), .Z(n15532) );
  NANDN U17914 ( .A(x[3795]), .B(y[3795]), .Z(n39527) );
  XNOR U17915 ( .A(x[3796]), .B(y[3796]), .Z(n9860) );
  AND U17916 ( .A(n39527), .B(n9860), .Z(n56044) );
  NANDN U17917 ( .A(y[3794]), .B(x[3794]), .Z(n25734) );
  NANDN U17918 ( .A(y[3795]), .B(x[3795]), .Z(n25733) );
  AND U17919 ( .A(n25734), .B(n25733), .Z(n56043) );
  NANDN U17920 ( .A(y[3792]), .B(x[3792]), .Z(n25738) );
  NANDN U17921 ( .A(y[3793]), .B(x[3793]), .Z(n25735) );
  AND U17922 ( .A(n25738), .B(n25735), .Z(n56041) );
  NANDN U17923 ( .A(x[3791]), .B(y[3791]), .Z(n39517) );
  NANDN U17924 ( .A(x[3792]), .B(y[3792]), .Z(n25737) );
  NAND U17925 ( .A(n39517), .B(n25737), .Z(n56040) );
  NANDN U17926 ( .A(y[3790]), .B(x[3790]), .Z(n9861) );
  NANDN U17927 ( .A(y[3791]), .B(x[3791]), .Z(n25739) );
  AND U17928 ( .A(n9861), .B(n25739), .Z(n56039) );
  XNOR U17929 ( .A(y[3790]), .B(x[3790]), .Z(n39514) );
  NANDN U17930 ( .A(x[3789]), .B(y[3789]), .Z(n25740) );
  NAND U17931 ( .A(n39514), .B(n25740), .Z(n56038) );
  NANDN U17932 ( .A(y[3788]), .B(x[3788]), .Z(n25743) );
  ANDN U17933 ( .B(x[3789]), .A(y[3789]), .Z(n39513) );
  ANDN U17934 ( .B(n25743), .A(n39513), .Z(n56037) );
  NANDN U17935 ( .A(x[3787]), .B(y[3787]), .Z(n25744) );
  NANDN U17936 ( .A(x[3788]), .B(y[3788]), .Z(n25741) );
  NAND U17937 ( .A(n25744), .B(n25741), .Z(n56036) );
  NANDN U17938 ( .A(x[3785]), .B(y[3785]), .Z(n39500) );
  NANDN U17939 ( .A(x[3786]), .B(y[3786]), .Z(n25745) );
  AND U17940 ( .A(n39500), .B(n25745), .Z(n56033) );
  NANDN U17941 ( .A(y[3784]), .B(x[3784]), .Z(n39497) );
  NANDN U17942 ( .A(y[3785]), .B(x[3785]), .Z(n25747) );
  NAND U17943 ( .A(n39497), .B(n25747), .Z(n56032) );
  NANDN U17944 ( .A(x[3783]), .B(y[3783]), .Z(n25748) );
  NANDN U17945 ( .A(x[3784]), .B(y[3784]), .Z(n39501) );
  AND U17946 ( .A(n25748), .B(n39501), .Z(n56031) );
  NANDN U17947 ( .A(y[3782]), .B(x[3782]), .Z(n39491) );
  NANDN U17948 ( .A(y[3783]), .B(x[3783]), .Z(n39498) );
  NAND U17949 ( .A(n39491), .B(n39498), .Z(n56030) );
  NANDN U17950 ( .A(x[3781]), .B(y[3781]), .Z(n25750) );
  NANDN U17951 ( .A(x[3782]), .B(y[3782]), .Z(n25749) );
  AND U17952 ( .A(n25750), .B(n25749), .Z(n56029) );
  XNOR U17953 ( .A(x[3780]), .B(y[3780]), .Z(n39485) );
  XNOR U17954 ( .A(x[3778]), .B(y[3778]), .Z(n25752) );
  NANDN U17955 ( .A(y[3776]), .B(x[3776]), .Z(n9862) );
  NANDN U17956 ( .A(y[3777]), .B(x[3777]), .Z(n25751) );
  NAND U17957 ( .A(n9862), .B(n25751), .Z(n56022) );
  XNOR U17958 ( .A(x[3776]), .B(y[3776]), .Z(n25754) );
  NANDN U17959 ( .A(x[3775]), .B(y[3775]), .Z(n56021) );
  AND U17960 ( .A(n25754), .B(n56021), .Z(n15505) );
  XNOR U17961 ( .A(x[3772]), .B(y[3772]), .Z(n39465) );
  NANDN U17962 ( .A(y[3770]), .B(x[3770]), .Z(n25757) );
  NANDN U17963 ( .A(y[3771]), .B(x[3771]), .Z(n39464) );
  AND U17964 ( .A(n25757), .B(n39464), .Z(n51801) );
  NANDN U17965 ( .A(x[3767]), .B(y[3767]), .Z(n25763) );
  NANDN U17966 ( .A(x[3768]), .B(y[3768]), .Z(n25760) );
  NAND U17967 ( .A(n25763), .B(n25760), .Z(n56014) );
  NANDN U17968 ( .A(y[3766]), .B(x[3766]), .Z(n39452) );
  NANDN U17969 ( .A(y[3767]), .B(x[3767]), .Z(n25762) );
  AND U17970 ( .A(n39452), .B(n25762), .Z(n51803) );
  NANDN U17971 ( .A(y[3764]), .B(x[3764]), .Z(n39443) );
  ANDN U17972 ( .B(x[3765]), .A(y[3765]), .Z(n39450) );
  ANDN U17973 ( .B(n39443), .A(n39450), .Z(n56012) );
  NANDN U17974 ( .A(y[3762]), .B(x[3762]), .Z(n39437) );
  NANDN U17975 ( .A(y[3763]), .B(x[3763]), .Z(n39444) );
  AND U17976 ( .A(n39437), .B(n39444), .Z(n56010) );
  NANDN U17977 ( .A(x[3761]), .B(y[3761]), .Z(n39433) );
  NANDN U17978 ( .A(x[3762]), .B(y[3762]), .Z(n25768) );
  NAND U17979 ( .A(n39433), .B(n25768), .Z(n56008) );
  NANDN U17980 ( .A(y[3760]), .B(x[3760]), .Z(n25769) );
  NANDN U17981 ( .A(y[3761]), .B(x[3761]), .Z(n39438) );
  AND U17982 ( .A(n25769), .B(n39438), .Z(n56007) );
  ANDN U17983 ( .B(y[3759]), .A(x[3759]), .Z(n39428) );
  NANDN U17984 ( .A(x[3760]), .B(y[3760]), .Z(n39434) );
  NANDN U17985 ( .A(n39428), .B(n39434), .Z(n56006) );
  NANDN U17986 ( .A(y[3758]), .B(x[3758]), .Z(n25771) );
  NANDN U17987 ( .A(y[3759]), .B(x[3759]), .Z(n25770) );
  AND U17988 ( .A(n25771), .B(n25770), .Z(n56005) );
  ANDN U17989 ( .B(y[3757]), .A(x[3757]), .Z(n39422) );
  ANDN U17990 ( .B(y[3758]), .A(x[3758]), .Z(n39429) );
  OR U17991 ( .A(n39422), .B(n39429), .Z(n56004) );
  XNOR U17992 ( .A(y[3756]), .B(x[3756]), .Z(n25774) );
  ANDN U17993 ( .B(y[3755]), .A(x[3755]), .Z(n39416) );
  ANDN U17994 ( .B(n25774), .A(n39416), .Z(n56002) );
  NANDN U17995 ( .A(y[3754]), .B(x[3754]), .Z(n9863) );
  NANDN U17996 ( .A(y[3755]), .B(x[3755]), .Z(n25773) );
  NAND U17997 ( .A(n9863), .B(n25773), .Z(n56001) );
  XNOR U17998 ( .A(y[3754]), .B(x[3754]), .Z(n25776) );
  NANDN U17999 ( .A(x[3753]), .B(y[3753]), .Z(n25777) );
  AND U18000 ( .A(n25776), .B(n25777), .Z(n51804) );
  NANDN U18001 ( .A(x[3751]), .B(y[3751]), .Z(n39406) );
  NANDN U18002 ( .A(x[3752]), .B(y[3752]), .Z(n25778) );
  AND U18003 ( .A(n39406), .B(n25778), .Z(n55999) );
  XNOR U18004 ( .A(y[3750]), .B(x[3750]), .Z(n39403) );
  NANDN U18005 ( .A(x[3749]), .B(y[3749]), .Z(n25781) );
  AND U18006 ( .A(n39403), .B(n25781), .Z(n55997) );
  ANDN U18007 ( .B(x[3749]), .A(y[3749]), .Z(n39402) );
  NANDN U18008 ( .A(y[3748]), .B(x[3748]), .Z(n25784) );
  NANDN U18009 ( .A(n39402), .B(n25784), .Z(n51805) );
  NANDN U18010 ( .A(x[3747]), .B(y[3747]), .Z(n25785) );
  NANDN U18011 ( .A(x[3748]), .B(y[3748]), .Z(n25782) );
  AND U18012 ( .A(n25785), .B(n25782), .Z(n51806) );
  NANDN U18013 ( .A(y[3744]), .B(x[3744]), .Z(n39386) );
  NANDN U18014 ( .A(y[3745]), .B(x[3745]), .Z(n39393) );
  NAND U18015 ( .A(n39386), .B(n39393), .Z(n55994) );
  NANDN U18016 ( .A(y[3742]), .B(x[3742]), .Z(n39380) );
  NANDN U18017 ( .A(y[3743]), .B(x[3743]), .Z(n39387) );
  AND U18018 ( .A(n39380), .B(n39387), .Z(n55993) );
  NANDN U18019 ( .A(x[3741]), .B(y[3741]), .Z(n25791) );
  NANDN U18020 ( .A(x[3742]), .B(y[3742]), .Z(n25790) );
  NAND U18021 ( .A(n25791), .B(n25790), .Z(n55992) );
  NANDN U18022 ( .A(y[3740]), .B(x[3740]), .Z(n25793) );
  NANDN U18023 ( .A(y[3741]), .B(x[3741]), .Z(n39381) );
  AND U18024 ( .A(n25793), .B(n39381), .Z(n51809) );
  NANDN U18025 ( .A(y[3736]), .B(x[3736]), .Z(n39363) );
  ANDN U18026 ( .B(x[3737]), .A(y[3737]), .Z(n39370) );
  ANDN U18027 ( .B(n39363), .A(n39370), .Z(n55988) );
  NANDN U18028 ( .A(x[3735]), .B(y[3735]), .Z(n25799) );
  NANDN U18029 ( .A(x[3736]), .B(y[3736]), .Z(n25798) );
  NAND U18030 ( .A(n25799), .B(n25798), .Z(n55987) );
  NANDN U18031 ( .A(y[3734]), .B(x[3734]), .Z(n39357) );
  NANDN U18032 ( .A(y[3735]), .B(x[3735]), .Z(n39364) );
  AND U18033 ( .A(n39357), .B(n39364), .Z(n51811) );
  NANDN U18034 ( .A(x[3729]), .B(y[3729]), .Z(n55983) );
  XNOR U18035 ( .A(x[3730]), .B(y[3730]), .Z(n39346) );
  AND U18036 ( .A(n55983), .B(n39346), .Z(n15451) );
  NANDN U18037 ( .A(y[3728]), .B(x[3728]), .Z(n25804) );
  NANDN U18038 ( .A(y[3729]), .B(x[3729]), .Z(n39345) );
  NAND U18039 ( .A(n25804), .B(n39345), .Z(n55982) );
  NANDN U18040 ( .A(x[3727]), .B(y[3727]), .Z(n39338) );
  NANDN U18041 ( .A(x[3728]), .B(y[3728]), .Z(n25803) );
  AND U18042 ( .A(n39338), .B(n25803), .Z(n55981) );
  NANDN U18043 ( .A(y[3726]), .B(x[3726]), .Z(n25806) );
  NANDN U18044 ( .A(y[3727]), .B(x[3727]), .Z(n25805) );
  NAND U18045 ( .A(n25806), .B(n25805), .Z(n55980) );
  NANDN U18046 ( .A(x[3725]), .B(y[3725]), .Z(n39333) );
  NANDN U18047 ( .A(x[3726]), .B(y[3726]), .Z(n39339) );
  AND U18048 ( .A(n39333), .B(n39339), .Z(n55979) );
  NANDN U18049 ( .A(y[3724]), .B(x[3724]), .Z(n9864) );
  NANDN U18050 ( .A(y[3725]), .B(x[3725]), .Z(n25807) );
  NAND U18051 ( .A(n9864), .B(n25807), .Z(n55978) );
  NANDN U18052 ( .A(y[3722]), .B(x[3722]), .Z(n9865) );
  ANDN U18053 ( .B(x[3723]), .A(y[3723]), .Z(n39331) );
  ANDN U18054 ( .B(n9865), .A(n39331), .Z(n55973) );
  XNOR U18055 ( .A(x[3722]), .B(y[3722]), .Z(n25809) );
  NANDN U18056 ( .A(y[3720]), .B(x[3720]), .Z(n25812) );
  NANDN U18057 ( .A(y[3721]), .B(x[3721]), .Z(n25808) );
  AND U18058 ( .A(n25812), .B(n25808), .Z(n55970) );
  NANDN U18059 ( .A(x[3719]), .B(y[3719]), .Z(n39316) );
  NANDN U18060 ( .A(x[3720]), .B(y[3720]), .Z(n25811) );
  AND U18061 ( .A(n39316), .B(n25811), .Z(n51815) );
  NANDN U18062 ( .A(y[3718]), .B(x[3718]), .Z(n25814) );
  NANDN U18063 ( .A(y[3719]), .B(x[3719]), .Z(n25813) );
  NAND U18064 ( .A(n25814), .B(n25813), .Z(n51816) );
  NANDN U18065 ( .A(x[3717]), .B(y[3717]), .Z(n39310) );
  NANDN U18066 ( .A(x[3718]), .B(y[3718]), .Z(n39317) );
  AND U18067 ( .A(n39310), .B(n39317), .Z(n55969) );
  NANDN U18068 ( .A(y[3714]), .B(x[3714]), .Z(n25818) );
  NANDN U18069 ( .A(y[3715]), .B(x[3715]), .Z(n25817) );
  NAND U18070 ( .A(n25818), .B(n25817), .Z(n55967) );
  NANDN U18071 ( .A(x[3713]), .B(y[3713]), .Z(n39298) );
  NANDN U18072 ( .A(x[3714]), .B(y[3714]), .Z(n39305) );
  AND U18073 ( .A(n39298), .B(n39305), .Z(n55966) );
  NANDN U18074 ( .A(y[3712]), .B(x[3712]), .Z(n39295) );
  NANDN U18075 ( .A(y[3713]), .B(x[3713]), .Z(n25819) );
  NAND U18076 ( .A(n39295), .B(n25819), .Z(n55965) );
  NANDN U18077 ( .A(x[3711]), .B(y[3711]), .Z(n25820) );
  NANDN U18078 ( .A(x[3712]), .B(y[3712]), .Z(n39299) );
  AND U18079 ( .A(n25820), .B(n39299), .Z(n55964) );
  NANDN U18080 ( .A(x[3709]), .B(y[3709]), .Z(n25822) );
  NANDN U18081 ( .A(x[3710]), .B(y[3710]), .Z(n25821) );
  AND U18082 ( .A(n25822), .B(n25821), .Z(n55961) );
  NANDN U18083 ( .A(y[3708]), .B(x[3708]), .Z(n39283) );
  NANDN U18084 ( .A(y[3709]), .B(x[3709]), .Z(n39290) );
  NAND U18085 ( .A(n39283), .B(n39290), .Z(n55960) );
  NANDN U18086 ( .A(x[3708]), .B(y[3708]), .Z(n25823) );
  ANDN U18087 ( .B(y[3707]), .A(x[3707]), .Z(n39279) );
  ANDN U18088 ( .B(n25823), .A(n39279), .Z(n55959) );
  NANDN U18089 ( .A(y[3706]), .B(x[3706]), .Z(n9866) );
  NANDN U18090 ( .A(y[3707]), .B(x[3707]), .Z(n39284) );
  NAND U18091 ( .A(n9866), .B(n39284), .Z(n55958) );
  NANDN U18092 ( .A(x[3705]), .B(y[3705]), .Z(n55957) );
  XNOR U18093 ( .A(x[3706]), .B(y[3706]), .Z(n25825) );
  AND U18094 ( .A(n55957), .B(n25825), .Z(n15424) );
  NANDN U18095 ( .A(y[3702]), .B(x[3702]), .Z(n25831) );
  NANDN U18096 ( .A(y[3703]), .B(x[3703]), .Z(n25828) );
  NAND U18097 ( .A(n25831), .B(n25828), .Z(n51819) );
  NANDN U18098 ( .A(x[3701]), .B(y[3701]), .Z(n39266) );
  NANDN U18099 ( .A(x[3702]), .B(y[3702]), .Z(n25830) );
  AND U18100 ( .A(n39266), .B(n25830), .Z(n55954) );
  NANDN U18101 ( .A(x[3699]), .B(y[3699]), .Z(n39260) );
  ANDN U18102 ( .B(y[3700]), .A(x[3700]), .Z(n39268) );
  ANDN U18103 ( .B(n39260), .A(n39268), .Z(n55952) );
  NANDN U18104 ( .A(y[3698]), .B(x[3698]), .Z(n25835) );
  NANDN U18105 ( .A(y[3699]), .B(x[3699]), .Z(n25834) );
  NAND U18106 ( .A(n25835), .B(n25834), .Z(n55951) );
  NANDN U18107 ( .A(x[3697]), .B(y[3697]), .Z(n25837) );
  NANDN U18108 ( .A(x[3698]), .B(y[3698]), .Z(n39261) );
  AND U18109 ( .A(n25837), .B(n39261), .Z(n51820) );
  XNOR U18110 ( .A(x[3694]), .B(y[3694]), .Z(n39248) );
  ANDN U18111 ( .B(x[3693]), .A(y[3693]), .Z(n39247) );
  NANDN U18112 ( .A(y[3692]), .B(x[3692]), .Z(n25843) );
  NANDN U18113 ( .A(n39247), .B(n25843), .Z(n55945) );
  NANDN U18114 ( .A(x[3691]), .B(y[3691]), .Z(n25844) );
  NANDN U18115 ( .A(x[3692]), .B(y[3692]), .Z(n25841) );
  AND U18116 ( .A(n25844), .B(n25841), .Z(n51822) );
  NANDN U18117 ( .A(y[3686]), .B(x[3686]), .Z(n25850) );
  NANDN U18118 ( .A(y[3687]), .B(x[3687]), .Z(n25849) );
  NAND U18119 ( .A(n25850), .B(n25849), .Z(n55941) );
  NANDN U18120 ( .A(x[3685]), .B(y[3685]), .Z(n39222) );
  NANDN U18121 ( .A(x[3686]), .B(y[3686]), .Z(n39229) );
  AND U18122 ( .A(n39222), .B(n39229), .Z(n55940) );
  NANDN U18123 ( .A(y[3684]), .B(x[3684]), .Z(n25852) );
  NANDN U18124 ( .A(y[3685]), .B(x[3685]), .Z(n25851) );
  NAND U18125 ( .A(n25852), .B(n25851), .Z(n55939) );
  NANDN U18126 ( .A(x[3683]), .B(y[3683]), .Z(n39216) );
  NANDN U18127 ( .A(x[3684]), .B(y[3684]), .Z(n39223) );
  AND U18128 ( .A(n39216), .B(n39223), .Z(n55938) );
  NANDN U18129 ( .A(x[3677]), .B(y[3677]), .Z(n39201) );
  NANDN U18130 ( .A(x[3678]), .B(y[3678]), .Z(n25859) );
  NAND U18131 ( .A(n39201), .B(n25859), .Z(n51826) );
  NANDN U18132 ( .A(y[3676]), .B(x[3676]), .Z(n25863) );
  NANDN U18133 ( .A(y[3677]), .B(x[3677]), .Z(n25861) );
  AND U18134 ( .A(n25863), .B(n25861), .Z(n55933) );
  NANDN U18135 ( .A(x[3673]), .B(y[3673]), .Z(n25868) );
  NANDN U18136 ( .A(x[3674]), .B(y[3674]), .Z(n25865) );
  NAND U18137 ( .A(n25868), .B(n25865), .Z(n51828) );
  NANDN U18138 ( .A(y[3670]), .B(x[3670]), .Z(n9867) );
  NANDN U18139 ( .A(y[3671]), .B(x[3671]), .Z(n25871) );
  NAND U18140 ( .A(n9867), .B(n25871), .Z(n51830) );
  XNOR U18141 ( .A(y[3670]), .B(x[3670]), .Z(n39183) );
  NANDN U18142 ( .A(x[3669]), .B(y[3669]), .Z(n25872) );
  AND U18143 ( .A(n39183), .B(n25872), .Z(n55927) );
  NANDN U18144 ( .A(y[3664]), .B(x[3664]), .Z(n25878) );
  NANDN U18145 ( .A(y[3665]), .B(x[3665]), .Z(n39172) );
  NAND U18146 ( .A(n25878), .B(n39172), .Z(n51832) );
  NANDN U18147 ( .A(x[3664]), .B(y[3664]), .Z(n25877) );
  ANDN U18148 ( .B(y[3663]), .A(x[3663]), .Z(n39165) );
  ANDN U18149 ( .B(n25877), .A(n39165), .Z(n55922) );
  NANDN U18150 ( .A(x[3661]), .B(y[3661]), .Z(n55920) );
  XNOR U18151 ( .A(x[3662]), .B(y[3662]), .Z(n25881) );
  AND U18152 ( .A(n55920), .B(n25881), .Z(n15376) );
  NANDN U18153 ( .A(y[3658]), .B(x[3658]), .Z(n25887) );
  NANDN U18154 ( .A(y[3659]), .B(x[3659]), .Z(n25884) );
  NAND U18155 ( .A(n25887), .B(n25884), .Z(n51834) );
  NANDN U18156 ( .A(x[3657]), .B(y[3657]), .Z(n25889) );
  NANDN U18157 ( .A(x[3658]), .B(y[3658]), .Z(n25886) );
  AND U18158 ( .A(n25889), .B(n25886), .Z(n55917) );
  XNOR U18159 ( .A(x[3656]), .B(y[3656]), .Z(n25891) );
  NANDN U18160 ( .A(x[3655]), .B(y[3655]), .Z(n55914) );
  AND U18161 ( .A(n25891), .B(n55914), .Z(n15368) );
  NANDN U18162 ( .A(x[3654]), .B(y[3654]), .Z(n25892) );
  ANDN U18163 ( .B(y[3653]), .A(x[3653]), .Z(n39143) );
  ANDN U18164 ( .B(n25892), .A(n39143), .Z(n55912) );
  NANDN U18165 ( .A(y[3652]), .B(x[3652]), .Z(n9868) );
  NANDN U18166 ( .A(y[3653]), .B(x[3653]), .Z(n25894) );
  NAND U18167 ( .A(n9868), .B(n25894), .Z(n51835) );
  XNOR U18168 ( .A(y[3652]), .B(x[3652]), .Z(n25896) );
  ANDN U18169 ( .B(y[3651]), .A(x[3651]), .Z(n39136) );
  ANDN U18170 ( .B(n25896), .A(n39136), .Z(n55910) );
  XNOR U18171 ( .A(y[3650]), .B(x[3650]), .Z(n25897) );
  NANDN U18172 ( .A(x[3649]), .B(y[3649]), .Z(n25898) );
  AND U18173 ( .A(n25897), .B(n25898), .Z(n55908) );
  NANDN U18174 ( .A(y[3648]), .B(x[3648]), .Z(n25899) );
  NANDN U18175 ( .A(y[3649]), .B(x[3649]), .Z(n55907) );
  NAND U18176 ( .A(n25899), .B(n55907), .Z(n55905) );
  NANDN U18177 ( .A(x[3647]), .B(y[3647]), .Z(n55904) );
  NANDN U18178 ( .A(y[3646]), .B(x[3646]), .Z(n9869) );
  NANDN U18179 ( .A(y[3647]), .B(x[3647]), .Z(n25900) );
  NAND U18180 ( .A(n9869), .B(n25900), .Z(n55903) );
  XNOR U18181 ( .A(x[3646]), .B(y[3646]), .Z(n39124) );
  NANDN U18182 ( .A(x[3645]), .B(y[3645]), .Z(n51837) );
  NANDN U18183 ( .A(y[3644]), .B(x[3644]), .Z(n9870) );
  NANDN U18184 ( .A(y[3645]), .B(x[3645]), .Z(n39125) );
  AND U18185 ( .A(n9870), .B(n39125), .Z(n55902) );
  XNOR U18186 ( .A(y[3644]), .B(x[3644]), .Z(n39118) );
  NANDN U18187 ( .A(x[3643]), .B(y[3643]), .Z(n25902) );
  NAND U18188 ( .A(n39118), .B(n25902), .Z(n55899) );
  NANDN U18189 ( .A(y[3642]), .B(x[3642]), .Z(n39112) );
  NANDN U18190 ( .A(y[3643]), .B(x[3643]), .Z(n39119) );
  AND U18191 ( .A(n39112), .B(n39119), .Z(n51838) );
  ANDN U18192 ( .B(y[3640]), .A(x[3640]), .Z(n39110) );
  NANDN U18193 ( .A(x[3639]), .B(y[3639]), .Z(n25904) );
  NANDN U18194 ( .A(n39110), .B(n25904), .Z(n55897) );
  NANDN U18195 ( .A(y[3638]), .B(x[3638]), .Z(n39097) );
  NANDN U18196 ( .A(y[3639]), .B(x[3639]), .Z(n39106) );
  AND U18197 ( .A(n39097), .B(n39106), .Z(n51840) );
  NANDN U18198 ( .A(x[3633]), .B(y[3633]), .Z(n25910) );
  NANDN U18199 ( .A(x[3634]), .B(y[3634]), .Z(n25909) );
  NAND U18200 ( .A(n25910), .B(n25909), .Z(n55892) );
  NANDN U18201 ( .A(y[3632]), .B(x[3632]), .Z(n39079) );
  NANDN U18202 ( .A(y[3633]), .B(x[3633]), .Z(n39086) );
  AND U18203 ( .A(n39079), .B(n39086), .Z(n51842) );
  NANDN U18204 ( .A(x[3627]), .B(y[3627]), .Z(n39064) );
  NANDN U18205 ( .A(x[3628]), .B(y[3628]), .Z(n39071) );
  NAND U18206 ( .A(n39064), .B(n39071), .Z(n55887) );
  NANDN U18207 ( .A(y[3626]), .B(x[3626]), .Z(n25915) );
  NANDN U18208 ( .A(y[3627]), .B(x[3627]), .Z(n25914) );
  AND U18209 ( .A(n25915), .B(n25914), .Z(n51846) );
  NANDN U18210 ( .A(x[3623]), .B(y[3623]), .Z(n39051) );
  NANDN U18211 ( .A(x[3624]), .B(y[3624]), .Z(n39059) );
  NAND U18212 ( .A(n39051), .B(n39059), .Z(n55885) );
  NANDN U18213 ( .A(y[3622]), .B(x[3622]), .Z(n25919) );
  NANDN U18214 ( .A(y[3623]), .B(x[3623]), .Z(n25918) );
  AND U18215 ( .A(n25919), .B(n25918), .Z(n51848) );
  NANDN U18216 ( .A(x[3617]), .B(y[3617]), .Z(n25923) );
  NANDN U18217 ( .A(x[3618]), .B(y[3618]), .Z(n39040) );
  NAND U18218 ( .A(n25923), .B(n39040), .Z(n55880) );
  NANDN U18219 ( .A(y[3616]), .B(x[3616]), .Z(n25925) );
  NANDN U18220 ( .A(y[3617]), .B(x[3617]), .Z(n39036) );
  AND U18221 ( .A(n25925), .B(n39036), .Z(n51850) );
  XNOR U18222 ( .A(x[3614]), .B(y[3614]), .Z(n25928) );
  NANDN U18223 ( .A(x[3613]), .B(y[3613]), .Z(n51852) );
  NAND U18224 ( .A(n25928), .B(n51852), .Z(n15318) );
  NANDN U18225 ( .A(x[3611]), .B(y[3611]), .Z(n39017) );
  NANDN U18226 ( .A(x[3612]), .B(y[3612]), .Z(n39023) );
  AND U18227 ( .A(n39017), .B(n39023), .Z(n55876) );
  NANDN U18228 ( .A(x[3609]), .B(y[3609]), .Z(n39011) );
  NANDN U18229 ( .A(x[3610]), .B(y[3610]), .Z(n39018) );
  AND U18230 ( .A(n39011), .B(n39018), .Z(n55873) );
  NANDN U18231 ( .A(y[3608]), .B(x[3608]), .Z(n25933) );
  NANDN U18232 ( .A(y[3609]), .B(x[3609]), .Z(n25932) );
  NAND U18233 ( .A(n25933), .B(n25932), .Z(n55872) );
  NANDN U18234 ( .A(x[3607]), .B(y[3607]), .Z(n39005) );
  NANDN U18235 ( .A(x[3608]), .B(y[3608]), .Z(n39012) );
  AND U18236 ( .A(n39005), .B(n39012), .Z(n55871) );
  NANDN U18237 ( .A(y[3606]), .B(x[3606]), .Z(n25935) );
  NANDN U18238 ( .A(y[3607]), .B(x[3607]), .Z(n25934) );
  NAND U18239 ( .A(n25935), .B(n25934), .Z(n55870) );
  NANDN U18240 ( .A(x[3605]), .B(y[3605]), .Z(n38999) );
  NANDN U18241 ( .A(x[3606]), .B(y[3606]), .Z(n39006) );
  AND U18242 ( .A(n38999), .B(n39006), .Z(n55869) );
  NANDN U18243 ( .A(y[3604]), .B(x[3604]), .Z(n38996) );
  NANDN U18244 ( .A(y[3605]), .B(x[3605]), .Z(n25936) );
  NAND U18245 ( .A(n38996), .B(n25936), .Z(n55868) );
  NANDN U18246 ( .A(y[3602]), .B(x[3602]), .Z(n38990) );
  NANDN U18247 ( .A(y[3603]), .B(x[3603]), .Z(n38997) );
  AND U18248 ( .A(n38990), .B(n38997), .Z(n55867) );
  NANDN U18249 ( .A(x[3601]), .B(y[3601]), .Z(n25939) );
  NANDN U18250 ( .A(x[3602]), .B(y[3602]), .Z(n25938) );
  NAND U18251 ( .A(n25939), .B(n25938), .Z(n55866) );
  NANDN U18252 ( .A(y[3600]), .B(x[3600]), .Z(n38984) );
  NANDN U18253 ( .A(y[3601]), .B(x[3601]), .Z(n38991) );
  AND U18254 ( .A(n38984), .B(n38991), .Z(n55865) );
  NANDN U18255 ( .A(x[3599]), .B(y[3599]), .Z(n25941) );
  NANDN U18256 ( .A(x[3600]), .B(y[3600]), .Z(n25940) );
  NAND U18257 ( .A(n25941), .B(n25940), .Z(n55864) );
  ANDN U18258 ( .B(y[3595]), .A(x[3595]), .Z(n25945) );
  NANDN U18259 ( .A(x[3596]), .B(y[3596]), .Z(n38974) );
  NANDN U18260 ( .A(n25945), .B(n38974), .Z(n55860) );
  NANDN U18261 ( .A(y[3594]), .B(x[3594]), .Z(n9871) );
  NANDN U18262 ( .A(y[3595]), .B(x[3595]), .Z(n25944) );
  AND U18263 ( .A(n9871), .B(n25944), .Z(n51857) );
  XNOR U18264 ( .A(y[3594]), .B(x[3594]), .Z(n38966) );
  NANDN U18265 ( .A(x[3593]), .B(y[3593]), .Z(n25947) );
  NAND U18266 ( .A(n38966), .B(n25947), .Z(n55859) );
  NANDN U18267 ( .A(y[3592]), .B(x[3592]), .Z(n38959) );
  NANDN U18268 ( .A(y[3593]), .B(x[3593]), .Z(n38965) );
  AND U18269 ( .A(n38959), .B(n38965), .Z(n55858) );
  NANDN U18270 ( .A(x[3591]), .B(y[3591]), .Z(n38955) );
  NANDN U18271 ( .A(x[3592]), .B(y[3592]), .Z(n25948) );
  NAND U18272 ( .A(n38955), .B(n25948), .Z(n55857) );
  NANDN U18273 ( .A(x[3590]), .B(y[3590]), .Z(n38956) );
  ANDN U18274 ( .B(y[3589]), .A(x[3589]), .Z(n38950) );
  ANDN U18275 ( .B(n38956), .A(n38950), .Z(n55855) );
  NANDN U18276 ( .A(y[3588]), .B(x[3588]), .Z(n9872) );
  NANDN U18277 ( .A(y[3589]), .B(x[3589]), .Z(n25950) );
  NAND U18278 ( .A(n9872), .B(n25950), .Z(n55854) );
  XNOR U18279 ( .A(y[3588]), .B(x[3588]), .Z(n38946) );
  NANDN U18280 ( .A(x[3587]), .B(y[3587]), .Z(n25951) );
  AND U18281 ( .A(n38946), .B(n25951), .Z(n55853) );
  NANDN U18282 ( .A(y[3586]), .B(x[3586]), .Z(n9873) );
  NANDN U18283 ( .A(y[3587]), .B(x[3587]), .Z(n38948) );
  NAND U18284 ( .A(n9873), .B(n38948), .Z(n55852) );
  XNOR U18285 ( .A(y[3586]), .B(x[3586]), .Z(n38940) );
  NANDN U18286 ( .A(x[3585]), .B(y[3585]), .Z(n25953) );
  AND U18287 ( .A(n38940), .B(n25953), .Z(n55851) );
  XNOR U18288 ( .A(x[3584]), .B(y[3584]), .Z(n38934) );
  NANDN U18289 ( .A(y[3582]), .B(x[3582]), .Z(n25955) );
  NANDN U18290 ( .A(y[3583]), .B(x[3583]), .Z(n38933) );
  AND U18291 ( .A(n25955), .B(n38933), .Z(n55847) );
  NANDN U18292 ( .A(x[3581]), .B(y[3581]), .Z(n38926) );
  NANDN U18293 ( .A(x[3582]), .B(y[3582]), .Z(n25954) );
  NAND U18294 ( .A(n38926), .B(n25954), .Z(n55846) );
  NANDN U18295 ( .A(y[3581]), .B(x[3581]), .Z(n25956) );
  ANDN U18296 ( .B(x[3580]), .A(y[3580]), .Z(n38922) );
  ANDN U18297 ( .B(n25956), .A(n38922), .Z(n55845) );
  NANDN U18298 ( .A(x[3579]), .B(y[3579]), .Z(n38918) );
  NANDN U18299 ( .A(x[3580]), .B(y[3580]), .Z(n38927) );
  NAND U18300 ( .A(n38918), .B(n38927), .Z(n51858) );
  NANDN U18301 ( .A(y[3578]), .B(x[3578]), .Z(n25957) );
  ANDN U18302 ( .B(x[3579]), .A(y[3579]), .Z(n38924) );
  ANDN U18303 ( .B(n25957), .A(n38924), .Z(n55843) );
  NANDN U18304 ( .A(y[3574]), .B(x[3574]), .Z(n25961) );
  NANDN U18305 ( .A(y[3575]), .B(x[3575]), .Z(n25960) );
  AND U18306 ( .A(n25961), .B(n25960), .Z(n55840) );
  NANDN U18307 ( .A(x[3573]), .B(y[3573]), .Z(n38901) );
  NANDN U18308 ( .A(x[3574]), .B(y[3574]), .Z(n38906) );
  NAND U18309 ( .A(n38901), .B(n38906), .Z(n55839) );
  NANDN U18310 ( .A(y[3572]), .B(x[3572]), .Z(n9874) );
  NANDN U18311 ( .A(y[3573]), .B(x[3573]), .Z(n25962) );
  AND U18312 ( .A(n9874), .B(n25962), .Z(n55838) );
  ANDN U18313 ( .B(y[3571]), .A(x[3571]), .Z(n25965) );
  XNOR U18314 ( .A(x[3572]), .B(y[3572]), .Z(n25964) );
  NANDN U18315 ( .A(y[3570]), .B(x[3570]), .Z(n25967) );
  NANDN U18316 ( .A(y[3571]), .B(x[3571]), .Z(n25963) );
  NAND U18317 ( .A(n25967), .B(n25963), .Z(n55835) );
  NANDN U18318 ( .A(x[3569]), .B(y[3569]), .Z(n38891) );
  NANDN U18319 ( .A(x[3570]), .B(y[3570]), .Z(n25966) );
  AND U18320 ( .A(n38891), .B(n25966), .Z(n55834) );
  NANDN U18321 ( .A(y[3568]), .B(x[3568]), .Z(n9875) );
  NANDN U18322 ( .A(y[3569]), .B(x[3569]), .Z(n25968) );
  NAND U18323 ( .A(n9875), .B(n25968), .Z(n55833) );
  XNOR U18324 ( .A(x[3568]), .B(y[3568]), .Z(n38889) );
  NANDN U18325 ( .A(x[3567]), .B(y[3567]), .Z(n55831) );
  AND U18326 ( .A(n38889), .B(n55831), .Z(n15267) );
  NANDN U18327 ( .A(y[3564]), .B(x[3564]), .Z(n25974) );
  NANDN U18328 ( .A(y[3565]), .B(x[3565]), .Z(n25970) );
  NAND U18329 ( .A(n25974), .B(n25970), .Z(n55829) );
  NANDN U18330 ( .A(x[3563]), .B(y[3563]), .Z(n38875) );
  NANDN U18331 ( .A(x[3564]), .B(y[3564]), .Z(n25973) );
  AND U18332 ( .A(n38875), .B(n25973), .Z(n55827) );
  NANDN U18333 ( .A(y[3562]), .B(x[3562]), .Z(n25976) );
  NANDN U18334 ( .A(y[3563]), .B(x[3563]), .Z(n25975) );
  NAND U18335 ( .A(n25976), .B(n25975), .Z(n55826) );
  NANDN U18336 ( .A(x[3561]), .B(y[3561]), .Z(n38869) );
  NANDN U18337 ( .A(x[3562]), .B(y[3562]), .Z(n38876) );
  AND U18338 ( .A(n38869), .B(n38876), .Z(n55825) );
  NANDN U18339 ( .A(y[3560]), .B(x[3560]), .Z(n25978) );
  NANDN U18340 ( .A(y[3561]), .B(x[3561]), .Z(n25977) );
  NAND U18341 ( .A(n25978), .B(n25977), .Z(n55824) );
  NANDN U18342 ( .A(y[3558]), .B(x[3558]), .Z(n25980) );
  NANDN U18343 ( .A(y[3559]), .B(x[3559]), .Z(n25979) );
  AND U18344 ( .A(n25980), .B(n25979), .Z(n55823) );
  NANDN U18345 ( .A(x[3557]), .B(y[3557]), .Z(n38857) );
  NANDN U18346 ( .A(x[3558]), .B(y[3558]), .Z(n38864) );
  NAND U18347 ( .A(n38857), .B(n38864), .Z(n55822) );
  NANDN U18348 ( .A(y[3556]), .B(x[3556]), .Z(n38853) );
  NANDN U18349 ( .A(y[3557]), .B(x[3557]), .Z(n25981) );
  AND U18350 ( .A(n38853), .B(n25981), .Z(n55821) );
  NANDN U18351 ( .A(x[3555]), .B(y[3555]), .Z(n38850) );
  NANDN U18352 ( .A(x[3556]), .B(y[3556]), .Z(n38858) );
  NAND U18353 ( .A(n38850), .B(n38858), .Z(n55820) );
  NANDN U18354 ( .A(y[3553]), .B(x[3553]), .Z(n25983) );
  ANDN U18355 ( .B(x[3552]), .A(y[3552]), .Z(n38842) );
  ANDN U18356 ( .B(n25983), .A(n38842), .Z(n55819) );
  NANDN U18357 ( .A(x[3551]), .B(y[3551]), .Z(n25986) );
  NANDN U18358 ( .A(x[3552]), .B(y[3552]), .Z(n25985) );
  NAND U18359 ( .A(n25986), .B(n25985), .Z(n55818) );
  NANDN U18360 ( .A(y[3550]), .B(x[3550]), .Z(n9876) );
  ANDN U18361 ( .B(x[3551]), .A(y[3551]), .Z(n38843) );
  ANDN U18362 ( .B(n9876), .A(n38843), .Z(n55817) );
  NANDN U18363 ( .A(x[3549]), .B(y[3549]), .Z(n55814) );
  NANDN U18364 ( .A(y[3548]), .B(x[3548]), .Z(n25987) );
  ANDN U18365 ( .B(x[3549]), .A(y[3549]), .Z(n38837) );
  ANDN U18366 ( .B(n25987), .A(n38837), .Z(n55812) );
  NANDN U18367 ( .A(x[3547]), .B(y[3547]), .Z(n25989) );
  NANDN U18368 ( .A(x[3548]), .B(y[3548]), .Z(n38832) );
  NAND U18369 ( .A(n25989), .B(n38832), .Z(n55811) );
  NANDN U18370 ( .A(y[3546]), .B(x[3546]), .Z(n38827) );
  NANDN U18371 ( .A(y[3547]), .B(x[3547]), .Z(n25988) );
  AND U18372 ( .A(n38827), .B(n25988), .Z(n55810) );
  NANDN U18373 ( .A(x[3545]), .B(y[3545]), .Z(n25991) );
  NANDN U18374 ( .A(x[3546]), .B(y[3546]), .Z(n25990) );
  NAND U18375 ( .A(n25991), .B(n25990), .Z(n55809) );
  NANDN U18376 ( .A(y[3544]), .B(x[3544]), .Z(n38818) );
  ANDN U18377 ( .B(x[3545]), .A(y[3545]), .Z(n38825) );
  ANDN U18378 ( .B(n38818), .A(n38825), .Z(n55808) );
  NANDN U18379 ( .A(y[3540]), .B(x[3540]), .Z(n25995) );
  NANDN U18380 ( .A(y[3541]), .B(x[3541]), .Z(n38812) );
  AND U18381 ( .A(n25995), .B(n38812), .Z(n55806) );
  ANDN U18382 ( .B(y[3539]), .A(x[3539]), .Z(n38805) );
  NANDN U18383 ( .A(x[3540]), .B(y[3540]), .Z(n25994) );
  NANDN U18384 ( .A(n38805), .B(n25994), .Z(n55805) );
  NANDN U18385 ( .A(y[3538]), .B(x[3538]), .Z(n25997) );
  NANDN U18386 ( .A(y[3539]), .B(x[3539]), .Z(n25996) );
  AND U18387 ( .A(n25997), .B(n25996), .Z(n55804) );
  ANDN U18388 ( .B(y[3537]), .A(x[3537]), .Z(n38800) );
  ANDN U18389 ( .B(y[3538]), .A(x[3538]), .Z(n38806) );
  OR U18390 ( .A(n38800), .B(n38806), .Z(n55803) );
  NANDN U18391 ( .A(y[3536]), .B(x[3536]), .Z(n9877) );
  NANDN U18392 ( .A(y[3537]), .B(x[3537]), .Z(n25998) );
  AND U18393 ( .A(n9877), .B(n25998), .Z(n55802) );
  NANDN U18394 ( .A(x[3533]), .B(y[3533]), .Z(n38790) );
  NANDN U18395 ( .A(x[3534]), .B(y[3534]), .Z(n26002) );
  NAND U18396 ( .A(n38790), .B(n26002), .Z(n51868) );
  NANDN U18397 ( .A(y[3532]), .B(x[3532]), .Z(n9878) );
  NANDN U18398 ( .A(y[3533]), .B(x[3533]), .Z(n26004) );
  AND U18399 ( .A(n9878), .B(n26004), .Z(n55798) );
  XNOR U18400 ( .A(x[3532]), .B(y[3532]), .Z(n38787) );
  NANDN U18401 ( .A(y[3530]), .B(x[3530]), .Z(n38781) );
  NANDN U18402 ( .A(y[3531]), .B(x[3531]), .Z(n38788) );
  NAND U18403 ( .A(n38781), .B(n38788), .Z(n51871) );
  NANDN U18404 ( .A(x[3529]), .B(y[3529]), .Z(n26007) );
  NANDN U18405 ( .A(x[3530]), .B(y[3530]), .Z(n26006) );
  AND U18406 ( .A(n26007), .B(n26006), .Z(n51872) );
  NANDN U18407 ( .A(x[3528]), .B(y[3528]), .Z(n26008) );
  ANDN U18408 ( .B(y[3527]), .A(x[3527]), .Z(n38773) );
  ANDN U18409 ( .B(n26008), .A(n38773), .Z(n55797) );
  NANDN U18410 ( .A(y[3526]), .B(x[3526]), .Z(n9879) );
  NANDN U18411 ( .A(y[3527]), .B(x[3527]), .Z(n38776) );
  NAND U18412 ( .A(n9879), .B(n38776), .Z(n55796) );
  XNOR U18413 ( .A(x[3526]), .B(y[3526]), .Z(n26010) );
  NANDN U18414 ( .A(y[3524]), .B(x[3524]), .Z(n26012) );
  NANDN U18415 ( .A(y[3525]), .B(x[3525]), .Z(n26009) );
  NAND U18416 ( .A(n26012), .B(n26009), .Z(n55793) );
  NANDN U18417 ( .A(x[3523]), .B(y[3523]), .Z(n26014) );
  NANDN U18418 ( .A(x[3524]), .B(y[3524]), .Z(n26011) );
  AND U18419 ( .A(n26014), .B(n26011), .Z(n55792) );
  NANDN U18420 ( .A(y[3522]), .B(x[3522]), .Z(n38759) );
  NANDN U18421 ( .A(y[3523]), .B(x[3523]), .Z(n26013) );
  NAND U18422 ( .A(n38759), .B(n26013), .Z(n55790) );
  NANDN U18423 ( .A(x[3521]), .B(y[3521]), .Z(n38756) );
  NANDN U18424 ( .A(x[3522]), .B(y[3522]), .Z(n26015) );
  AND U18425 ( .A(n38756), .B(n26015), .Z(n55789) );
  NANDN U18426 ( .A(y[3520]), .B(x[3520]), .Z(n38751) );
  NANDN U18427 ( .A(y[3521]), .B(x[3521]), .Z(n38760) );
  NAND U18428 ( .A(n38751), .B(n38760), .Z(n55788) );
  NANDN U18429 ( .A(x[3519]), .B(y[3519]), .Z(n26016) );
  NANDN U18430 ( .A(x[3520]), .B(y[3520]), .Z(n38757) );
  NAND U18431 ( .A(n26016), .B(n38757), .Z(n55787) );
  NANDN U18432 ( .A(y[3518]), .B(x[3518]), .Z(n9880) );
  NANDN U18433 ( .A(y[3519]), .B(x[3519]), .Z(n38752) );
  AND U18434 ( .A(n9880), .B(n38752), .Z(n55786) );
  XNOR U18435 ( .A(y[3518]), .B(x[3518]), .Z(n38746) );
  NANDN U18436 ( .A(x[3517]), .B(y[3517]), .Z(n38742) );
  NAND U18437 ( .A(n38746), .B(n38742), .Z(n55785) );
  NANDN U18438 ( .A(y[3516]), .B(x[3516]), .Z(n9881) );
  NANDN U18439 ( .A(y[3517]), .B(x[3517]), .Z(n38745) );
  AND U18440 ( .A(n9881), .B(n38745), .Z(n55784) );
  XNOR U18441 ( .A(y[3516]), .B(x[3516]), .Z(n26019) );
  NANDN U18442 ( .A(x[3515]), .B(y[3515]), .Z(n38736) );
  NAND U18443 ( .A(n26019), .B(n38736), .Z(n55783) );
  NANDN U18444 ( .A(y[3514]), .B(x[3514]), .Z(n26020) );
  NANDN U18445 ( .A(y[3515]), .B(x[3515]), .Z(n26018) );
  NAND U18446 ( .A(n26020), .B(n26018), .Z(n51874) );
  NANDN U18447 ( .A(x[3513]), .B(y[3513]), .Z(n38730) );
  NANDN U18448 ( .A(x[3514]), .B(y[3514]), .Z(n38737) );
  AND U18449 ( .A(n38730), .B(n38737), .Z(n51875) );
  NANDN U18450 ( .A(y[3510]), .B(x[3510]), .Z(n26024) );
  NANDN U18451 ( .A(y[3511]), .B(x[3511]), .Z(n26023) );
  NAND U18452 ( .A(n26024), .B(n26023), .Z(n55781) );
  NANDN U18453 ( .A(x[3509]), .B(y[3509]), .Z(n26026) );
  NANDN U18454 ( .A(x[3510]), .B(y[3510]), .Z(n38725) );
  NAND U18455 ( .A(n26026), .B(n38725), .Z(n55780) );
  NANDN U18456 ( .A(y[3508]), .B(x[3508]), .Z(n26028) );
  NANDN U18457 ( .A(y[3509]), .B(x[3509]), .Z(n26025) );
  AND U18458 ( .A(n26028), .B(n26025), .Z(n55779) );
  NANDN U18459 ( .A(x[3507]), .B(y[3507]), .Z(n38714) );
  NANDN U18460 ( .A(x[3508]), .B(y[3508]), .Z(n26027) );
  NAND U18461 ( .A(n38714), .B(n26027), .Z(n55777) );
  NANDN U18462 ( .A(y[3506]), .B(x[3506]), .Z(n9882) );
  NANDN U18463 ( .A(y[3507]), .B(x[3507]), .Z(n26029) );
  AND U18464 ( .A(n9882), .B(n26029), .Z(n55776) );
  NANDN U18465 ( .A(y[3504]), .B(x[3504]), .Z(n38705) );
  NANDN U18466 ( .A(y[3505]), .B(x[3505]), .Z(n38712) );
  AND U18467 ( .A(n38705), .B(n38712), .Z(n55773) );
  NANDN U18468 ( .A(x[3503]), .B(y[3503]), .Z(n26031) );
  NANDN U18469 ( .A(x[3504]), .B(y[3504]), .Z(n26030) );
  NAND U18470 ( .A(n26031), .B(n26030), .Z(n55772) );
  NANDN U18471 ( .A(y[3502]), .B(x[3502]), .Z(n38699) );
  NANDN U18472 ( .A(y[3503]), .B(x[3503]), .Z(n38706) );
  AND U18473 ( .A(n38699), .B(n38706), .Z(n55771) );
  NANDN U18474 ( .A(x[3501]), .B(y[3501]), .Z(n26033) );
  NANDN U18475 ( .A(x[3502]), .B(y[3502]), .Z(n26032) );
  NAND U18476 ( .A(n26033), .B(n26032), .Z(n55770) );
  NANDN U18477 ( .A(y[3500]), .B(x[3500]), .Z(n26035) );
  NANDN U18478 ( .A(y[3501]), .B(x[3501]), .Z(n38700) );
  AND U18479 ( .A(n26035), .B(n38700), .Z(n55769) );
  NANDN U18480 ( .A(y[3498]), .B(x[3498]), .Z(n26038) );
  NANDN U18481 ( .A(y[3499]), .B(x[3499]), .Z(n26036) );
  AND U18482 ( .A(n26038), .B(n26036), .Z(n55767) );
  NANDN U18483 ( .A(x[3498]), .B(y[3498]), .Z(n55766) );
  NANDN U18484 ( .A(y[3496]), .B(x[3496]), .Z(n9883) );
  NANDN U18485 ( .A(y[3497]), .B(x[3497]), .Z(n51878) );
  AND U18486 ( .A(n9883), .B(n51878), .Z(n55765) );
  NANDN U18487 ( .A(x[3495]), .B(y[3495]), .Z(n55764) );
  NANDN U18488 ( .A(y[3494]), .B(x[3494]), .Z(n26043) );
  NANDN U18489 ( .A(y[3495]), .B(x[3495]), .Z(n26040) );
  AND U18490 ( .A(n26043), .B(n26040), .Z(n55763) );
  NANDN U18491 ( .A(x[3493]), .B(y[3493]), .Z(n26045) );
  NANDN U18492 ( .A(x[3494]), .B(y[3494]), .Z(n26042) );
  NAND U18493 ( .A(n26045), .B(n26042), .Z(n55762) );
  NANDN U18494 ( .A(x[3491]), .B(y[3491]), .Z(n26047) );
  NANDN U18495 ( .A(x[3492]), .B(y[3492]), .Z(n26046) );
  NAND U18496 ( .A(n26047), .B(n26046), .Z(n51880) );
  NANDN U18497 ( .A(y[3490]), .B(x[3490]), .Z(n38671) );
  NANDN U18498 ( .A(y[3491]), .B(x[3491]), .Z(n38678) );
  NAND U18499 ( .A(n38671), .B(n38678), .Z(n55759) );
  NANDN U18500 ( .A(x[3489]), .B(y[3489]), .Z(n26049) );
  NANDN U18501 ( .A(x[3490]), .B(y[3490]), .Z(n26048) );
  AND U18502 ( .A(n26049), .B(n26048), .Z(n55758) );
  NANDN U18503 ( .A(y[3488]), .B(x[3488]), .Z(n26051) );
  NANDN U18504 ( .A(y[3489]), .B(x[3489]), .Z(n38672) );
  NAND U18505 ( .A(n26051), .B(n38672), .Z(n55757) );
  NANDN U18506 ( .A(x[3487]), .B(y[3487]), .Z(n38664) );
  XNOR U18507 ( .A(x[3488]), .B(y[3488]), .Z(n9884) );
  AND U18508 ( .A(n38664), .B(n9884), .Z(n55756) );
  NANDN U18509 ( .A(y[3486]), .B(x[3486]), .Z(n9885) );
  NANDN U18510 ( .A(y[3487]), .B(x[3487]), .Z(n26052) );
  NAND U18511 ( .A(n9885), .B(n26052), .Z(n55755) );
  XNOR U18512 ( .A(y[3486]), .B(x[3486]), .Z(n38660) );
  NANDN U18513 ( .A(x[3485]), .B(y[3485]), .Z(n38656) );
  NAND U18514 ( .A(n38660), .B(n38656), .Z(n55754) );
  NANDN U18515 ( .A(y[3484]), .B(x[3484]), .Z(n9886) );
  NANDN U18516 ( .A(y[3485]), .B(x[3485]), .Z(n38659) );
  AND U18517 ( .A(n9886), .B(n38659), .Z(n55753) );
  XNOR U18518 ( .A(y[3484]), .B(x[3484]), .Z(n26054) );
  NANDN U18519 ( .A(x[3483]), .B(y[3483]), .Z(n38650) );
  NAND U18520 ( .A(n26054), .B(n38650), .Z(n55752) );
  NANDN U18521 ( .A(y[3482]), .B(x[3482]), .Z(n26055) );
  NANDN U18522 ( .A(y[3483]), .B(x[3483]), .Z(n26053) );
  AND U18523 ( .A(n26055), .B(n26053), .Z(n55751) );
  NANDN U18524 ( .A(x[3481]), .B(y[3481]), .Z(n26057) );
  NANDN U18525 ( .A(x[3482]), .B(y[3482]), .Z(n38651) );
  NAND U18526 ( .A(n26057), .B(n38651), .Z(n55750) );
  NANDN U18527 ( .A(y[3480]), .B(x[3480]), .Z(n26059) );
  NANDN U18528 ( .A(y[3481]), .B(x[3481]), .Z(n26056) );
  NAND U18529 ( .A(n26059), .B(n26056), .Z(n55749) );
  NANDN U18530 ( .A(x[3479]), .B(y[3479]), .Z(n38640) );
  NANDN U18531 ( .A(x[3480]), .B(y[3480]), .Z(n26058) );
  AND U18532 ( .A(n38640), .B(n26058), .Z(n55748) );
  NANDN U18533 ( .A(y[3478]), .B(x[3478]), .Z(n9887) );
  NANDN U18534 ( .A(y[3479]), .B(x[3479]), .Z(n26060) );
  NAND U18535 ( .A(n9887), .B(n26060), .Z(n55747) );
  NANDN U18536 ( .A(x[3477]), .B(y[3477]), .Z(n51881) );
  XNOR U18537 ( .A(x[3478]), .B(y[3478]), .Z(n38637) );
  AND U18538 ( .A(n51881), .B(n38637), .Z(n15166) );
  NANDN U18539 ( .A(y[3476]), .B(x[3476]), .Z(n26063) );
  NANDN U18540 ( .A(y[3477]), .B(x[3477]), .Z(n38636) );
  AND U18541 ( .A(n26063), .B(n38636), .Z(n55746) );
  NANDN U18542 ( .A(x[3475]), .B(y[3475]), .Z(n26064) );
  NANDN U18543 ( .A(x[3476]), .B(y[3476]), .Z(n26061) );
  NAND U18544 ( .A(n26064), .B(n26061), .Z(n55745) );
  NANDN U18545 ( .A(y[3474]), .B(x[3474]), .Z(n26066) );
  NANDN U18546 ( .A(y[3475]), .B(x[3475]), .Z(n26062) );
  AND U18547 ( .A(n26066), .B(n26062), .Z(n55744) );
  NANDN U18548 ( .A(x[3473]), .B(y[3473]), .Z(n38624) );
  NANDN U18549 ( .A(x[3474]), .B(y[3474]), .Z(n26065) );
  NAND U18550 ( .A(n38624), .B(n26065), .Z(n55742) );
  NANDN U18551 ( .A(y[3472]), .B(x[3472]), .Z(n38621) );
  NANDN U18552 ( .A(y[3473]), .B(x[3473]), .Z(n26067) );
  AND U18553 ( .A(n38621), .B(n26067), .Z(n55740) );
  NANDN U18554 ( .A(x[3471]), .B(y[3471]), .Z(n26068) );
  NANDN U18555 ( .A(x[3472]), .B(y[3472]), .Z(n38625) );
  NAND U18556 ( .A(n26068), .B(n38625), .Z(n55738) );
  NANDN U18557 ( .A(y[3470]), .B(x[3470]), .Z(n38615) );
  NANDN U18558 ( .A(y[3471]), .B(x[3471]), .Z(n38622) );
  NAND U18559 ( .A(n38615), .B(n38622), .Z(n55736) );
  NANDN U18560 ( .A(x[3469]), .B(y[3469]), .Z(n26070) );
  NANDN U18561 ( .A(x[3470]), .B(y[3470]), .Z(n26069) );
  AND U18562 ( .A(n26070), .B(n26069), .Z(n55734) );
  NANDN U18563 ( .A(y[3468]), .B(x[3468]), .Z(n38609) );
  NANDN U18564 ( .A(y[3469]), .B(x[3469]), .Z(n38616) );
  NAND U18565 ( .A(n38609), .B(n38616), .Z(n55732) );
  NANDN U18566 ( .A(x[3467]), .B(y[3467]), .Z(n26072) );
  NANDN U18567 ( .A(x[3468]), .B(y[3468]), .Z(n26071) );
  AND U18568 ( .A(n26072), .B(n26071), .Z(n55730) );
  NANDN U18569 ( .A(y[3466]), .B(x[3466]), .Z(n38603) );
  NANDN U18570 ( .A(y[3467]), .B(x[3467]), .Z(n38610) );
  NAND U18571 ( .A(n38603), .B(n38610), .Z(n55728) );
  NANDN U18572 ( .A(x[3465]), .B(y[3465]), .Z(n26074) );
  NANDN U18573 ( .A(x[3466]), .B(y[3466]), .Z(n26073) );
  NAND U18574 ( .A(n26074), .B(n26073), .Z(n55726) );
  NANDN U18575 ( .A(y[3464]), .B(x[3464]), .Z(n38597) );
  NANDN U18576 ( .A(y[3465]), .B(x[3465]), .Z(n38604) );
  AND U18577 ( .A(n38597), .B(n38604), .Z(n55724) );
  NANDN U18578 ( .A(x[3463]), .B(y[3463]), .Z(n26076) );
  NANDN U18579 ( .A(x[3464]), .B(y[3464]), .Z(n26075) );
  NAND U18580 ( .A(n26076), .B(n26075), .Z(n55722) );
  NANDN U18581 ( .A(y[3462]), .B(x[3462]), .Z(n9888) );
  NANDN U18582 ( .A(y[3463]), .B(x[3463]), .Z(n38598) );
  AND U18583 ( .A(n9888), .B(n38598), .Z(n55720) );
  NANDN U18584 ( .A(y[3460]), .B(x[3460]), .Z(n26078) );
  NANDN U18585 ( .A(y[3461]), .B(x[3461]), .Z(n38590) );
  NAND U18586 ( .A(n26078), .B(n38590), .Z(n55714) );
  NANDN U18587 ( .A(x[3459]), .B(y[3459]), .Z(n26080) );
  NANDN U18588 ( .A(x[3460]), .B(y[3460]), .Z(n26077) );
  AND U18589 ( .A(n26080), .B(n26077), .Z(n55712) );
  NANDN U18590 ( .A(y[3458]), .B(x[3458]), .Z(n26082) );
  NANDN U18591 ( .A(y[3459]), .B(x[3459]), .Z(n26079) );
  NAND U18592 ( .A(n26082), .B(n26079), .Z(n55710) );
  NANDN U18593 ( .A(x[3457]), .B(y[3457]), .Z(n26084) );
  NANDN U18594 ( .A(x[3458]), .B(y[3458]), .Z(n26081) );
  AND U18595 ( .A(n26084), .B(n26081), .Z(n55708) );
  NANDN U18596 ( .A(y[3456]), .B(x[3456]), .Z(n26086) );
  NANDN U18597 ( .A(y[3457]), .B(x[3457]), .Z(n26083) );
  NAND U18598 ( .A(n26086), .B(n26083), .Z(n55706) );
  NANDN U18599 ( .A(x[3455]), .B(y[3455]), .Z(n26089) );
  NANDN U18600 ( .A(x[3456]), .B(y[3456]), .Z(n26085) );
  NAND U18601 ( .A(n26089), .B(n26085), .Z(n55704) );
  NANDN U18602 ( .A(y[3454]), .B(x[3454]), .Z(n26090) );
  NANDN U18603 ( .A(y[3455]), .B(x[3455]), .Z(n26087) );
  AND U18604 ( .A(n26090), .B(n26087), .Z(n55702) );
  NANDN U18605 ( .A(x[3453]), .B(y[3453]), .Z(n26092) );
  NANDN U18606 ( .A(x[3454]), .B(y[3454]), .Z(n26088) );
  NAND U18607 ( .A(n26092), .B(n26088), .Z(n55700) );
  NANDN U18608 ( .A(y[3452]), .B(x[3452]), .Z(n26094) );
  NANDN U18609 ( .A(y[3453]), .B(x[3453]), .Z(n26091) );
  AND U18610 ( .A(n26094), .B(n26091), .Z(n55698) );
  NANDN U18611 ( .A(x[3451]), .B(y[3451]), .Z(n38567) );
  NANDN U18612 ( .A(x[3452]), .B(y[3452]), .Z(n26093) );
  NAND U18613 ( .A(n38567), .B(n26093), .Z(n55696) );
  NANDN U18614 ( .A(y[3450]), .B(x[3450]), .Z(n9889) );
  NANDN U18615 ( .A(y[3451]), .B(x[3451]), .Z(n26095) );
  NAND U18616 ( .A(n9889), .B(n26095), .Z(n55694) );
  XNOR U18617 ( .A(y[3450]), .B(x[3450]), .Z(n26097) );
  NANDN U18618 ( .A(x[3449]), .B(y[3449]), .Z(n38561) );
  AND U18619 ( .A(n26097), .B(n38561), .Z(n55692) );
  NANDN U18620 ( .A(y[3448]), .B(x[3448]), .Z(n26098) );
  NANDN U18621 ( .A(y[3449]), .B(x[3449]), .Z(n26096) );
  NAND U18622 ( .A(n26098), .B(n26096), .Z(n55690) );
  NANDN U18623 ( .A(x[3447]), .B(y[3447]), .Z(n38555) );
  NANDN U18624 ( .A(x[3448]), .B(y[3448]), .Z(n38562) );
  AND U18625 ( .A(n38555), .B(n38562), .Z(n55688) );
  NANDN U18626 ( .A(y[3446]), .B(x[3446]), .Z(n26100) );
  NANDN U18627 ( .A(y[3447]), .B(x[3447]), .Z(n26099) );
  NAND U18628 ( .A(n26100), .B(n26099), .Z(n55686) );
  NANDN U18629 ( .A(x[3445]), .B(y[3445]), .Z(n26102) );
  NANDN U18630 ( .A(x[3446]), .B(y[3446]), .Z(n38556) );
  NAND U18631 ( .A(n26102), .B(n38556), .Z(n55684) );
  NANDN U18632 ( .A(y[3444]), .B(x[3444]), .Z(n26104) );
  NANDN U18633 ( .A(y[3445]), .B(x[3445]), .Z(n26101) );
  AND U18634 ( .A(n26104), .B(n26101), .Z(n55682) );
  NANDN U18635 ( .A(x[3443]), .B(y[3443]), .Z(n38547) );
  NANDN U18636 ( .A(x[3444]), .B(y[3444]), .Z(n26103) );
  NAND U18637 ( .A(n38547), .B(n26103), .Z(n55680) );
  NANDN U18638 ( .A(y[3442]), .B(x[3442]), .Z(n26106) );
  NANDN U18639 ( .A(y[3443]), .B(x[3443]), .Z(n26105) );
  AND U18640 ( .A(n26106), .B(n26105), .Z(n55678) );
  ANDN U18641 ( .B(y[3442]), .A(x[3442]), .Z(n38545) );
  NANDN U18642 ( .A(x[3441]), .B(y[3441]), .Z(n38538) );
  NANDN U18643 ( .A(n38545), .B(n38538), .Z(n55676) );
  NANDN U18644 ( .A(y[3440]), .B(x[3440]), .Z(n26108) );
  NANDN U18645 ( .A(y[3441]), .B(x[3441]), .Z(n26107) );
  NAND U18646 ( .A(n26108), .B(n26107), .Z(n55674) );
  NANDN U18647 ( .A(x[3439]), .B(y[3439]), .Z(n26110) );
  NANDN U18648 ( .A(x[3440]), .B(y[3440]), .Z(n38539) );
  AND U18649 ( .A(n26110), .B(n38539), .Z(n55672) );
  NANDN U18650 ( .A(y[3438]), .B(x[3438]), .Z(n38531) );
  NANDN U18651 ( .A(y[3439]), .B(x[3439]), .Z(n26109) );
  NAND U18652 ( .A(n38531), .B(n26109), .Z(n55670) );
  NANDN U18653 ( .A(x[3437]), .B(y[3437]), .Z(n38526) );
  XNOR U18654 ( .A(y[3438]), .B(x[3438]), .Z(n9890) );
  AND U18655 ( .A(n38526), .B(n9890), .Z(n55668) );
  NANDN U18656 ( .A(y[3436]), .B(x[3436]), .Z(n9891) );
  NANDN U18657 ( .A(y[3437]), .B(x[3437]), .Z(n38532) );
  NAND U18658 ( .A(n9891), .B(n38532), .Z(n55666) );
  XNOR U18659 ( .A(y[3436]), .B(x[3436]), .Z(n26113) );
  NANDN U18660 ( .A(x[3435]), .B(y[3435]), .Z(n38520) );
  NAND U18661 ( .A(n26113), .B(n38520), .Z(n55664) );
  NANDN U18662 ( .A(y[3434]), .B(x[3434]), .Z(n26114) );
  NANDN U18663 ( .A(y[3435]), .B(x[3435]), .Z(n26112) );
  AND U18664 ( .A(n26114), .B(n26112), .Z(n55662) );
  NANDN U18665 ( .A(x[3433]), .B(y[3433]), .Z(n38515) );
  NANDN U18666 ( .A(x[3434]), .B(y[3434]), .Z(n38521) );
  NAND U18667 ( .A(n38515), .B(n38521), .Z(n55661) );
  NANDN U18668 ( .A(y[3432]), .B(x[3432]), .Z(n9892) );
  NANDN U18669 ( .A(y[3433]), .B(x[3433]), .Z(n26115) );
  AND U18670 ( .A(n9892), .B(n26115), .Z(n55660) );
  XNOR U18671 ( .A(x[3432]), .B(y[3432]), .Z(n38513) );
  NANDN U18672 ( .A(y[3428]), .B(x[3428]), .Z(n26121) );
  NANDN U18673 ( .A(y[3429]), .B(x[3429]), .Z(n26117) );
  NAND U18674 ( .A(n26121), .B(n26117), .Z(n55655) );
  NANDN U18675 ( .A(x[3427]), .B(y[3427]), .Z(n38499) );
  NANDN U18676 ( .A(x[3428]), .B(y[3428]), .Z(n26120) );
  NAND U18677 ( .A(n38499), .B(n26120), .Z(n55654) );
  NANDN U18678 ( .A(y[3426]), .B(x[3426]), .Z(n38495) );
  NANDN U18679 ( .A(y[3427]), .B(x[3427]), .Z(n26122) );
  AND U18680 ( .A(n38495), .B(n26122), .Z(n55653) );
  NANDN U18681 ( .A(x[3425]), .B(y[3425]), .Z(n38492) );
  NANDN U18682 ( .A(x[3426]), .B(y[3426]), .Z(n38500) );
  NAND U18683 ( .A(n38492), .B(n38500), .Z(n55652) );
  NANDN U18684 ( .A(y[3424]), .B(x[3424]), .Z(n9893) );
  NANDN U18685 ( .A(y[3425]), .B(x[3425]), .Z(n38496) );
  AND U18686 ( .A(n9893), .B(n38496), .Z(n55651) );
  NANDN U18687 ( .A(y[3422]), .B(x[3422]), .Z(n38483) );
  NANDN U18688 ( .A(y[3423]), .B(x[3423]), .Z(n38490) );
  NAND U18689 ( .A(n38483), .B(n38490), .Z(n55648) );
  NANDN U18690 ( .A(x[3421]), .B(y[3421]), .Z(n26124) );
  NANDN U18691 ( .A(x[3422]), .B(y[3422]), .Z(n26123) );
  AND U18692 ( .A(n26124), .B(n26123), .Z(n55647) );
  NANDN U18693 ( .A(y[3420]), .B(x[3420]), .Z(n38477) );
  NANDN U18694 ( .A(y[3421]), .B(x[3421]), .Z(n38484) );
  NAND U18695 ( .A(n38477), .B(n38484), .Z(n55646) );
  NANDN U18696 ( .A(x[3420]), .B(y[3420]), .Z(n26125) );
  ANDN U18697 ( .B(y[3419]), .A(x[3419]), .Z(n38475) );
  ANDN U18698 ( .B(n26125), .A(n38475), .Z(n55644) );
  NANDN U18699 ( .A(y[3418]), .B(x[3418]), .Z(n9894) );
  NANDN U18700 ( .A(y[3419]), .B(x[3419]), .Z(n38478) );
  NAND U18701 ( .A(n9894), .B(n38478), .Z(n55643) );
  NANDN U18702 ( .A(x[3417]), .B(y[3417]), .Z(n55641) );
  NANDN U18703 ( .A(y[3416]), .B(x[3416]), .Z(n26129) );
  NANDN U18704 ( .A(y[3417]), .B(x[3417]), .Z(n26126) );
  AND U18705 ( .A(n26129), .B(n26126), .Z(n55640) );
  NANDN U18706 ( .A(x[3415]), .B(y[3415]), .Z(n26131) );
  NANDN U18707 ( .A(x[3416]), .B(y[3416]), .Z(n26128) );
  NAND U18708 ( .A(n26131), .B(n26128), .Z(n55639) );
  NANDN U18709 ( .A(y[3414]), .B(x[3414]), .Z(n38461) );
  NANDN U18710 ( .A(y[3415]), .B(x[3415]), .Z(n26130) );
  AND U18711 ( .A(n38461), .B(n26130), .Z(n55638) );
  NANDN U18712 ( .A(x[3413]), .B(y[3413]), .Z(n26133) );
  NANDN U18713 ( .A(x[3414]), .B(y[3414]), .Z(n26132) );
  NAND U18714 ( .A(n26133), .B(n26132), .Z(n55637) );
  NANDN U18715 ( .A(y[3412]), .B(x[3412]), .Z(n38455) );
  NANDN U18716 ( .A(y[3413]), .B(x[3413]), .Z(n38462) );
  NAND U18717 ( .A(n38455), .B(n38462), .Z(n55636) );
  NANDN U18718 ( .A(x[3411]), .B(y[3411]), .Z(n26135) );
  NANDN U18719 ( .A(x[3412]), .B(y[3412]), .Z(n26134) );
  AND U18720 ( .A(n26135), .B(n26134), .Z(n55635) );
  NANDN U18721 ( .A(y[3410]), .B(x[3410]), .Z(n38449) );
  NANDN U18722 ( .A(y[3411]), .B(x[3411]), .Z(n38456) );
  NAND U18723 ( .A(n38449), .B(n38456), .Z(n55634) );
  NANDN U18724 ( .A(x[3409]), .B(y[3409]), .Z(n26137) );
  NANDN U18725 ( .A(x[3410]), .B(y[3410]), .Z(n26136) );
  AND U18726 ( .A(n26137), .B(n26136), .Z(n55633) );
  NANDN U18727 ( .A(y[3408]), .B(x[3408]), .Z(n9895) );
  NANDN U18728 ( .A(y[3409]), .B(x[3409]), .Z(n38450) );
  NAND U18729 ( .A(n9895), .B(n38450), .Z(n55632) );
  NANDN U18730 ( .A(x[3407]), .B(y[3407]), .Z(n51883) );
  XNOR U18731 ( .A(x[3408]), .B(y[3408]), .Z(n38444) );
  NANDN U18732 ( .A(y[3406]), .B(x[3406]), .Z(n38437) );
  NANDN U18733 ( .A(y[3407]), .B(x[3407]), .Z(n38443) );
  NAND U18734 ( .A(n38437), .B(n38443), .Z(n51884) );
  NANDN U18735 ( .A(x[3405]), .B(y[3405]), .Z(n26139) );
  NANDN U18736 ( .A(x[3406]), .B(y[3406]), .Z(n26138) );
  AND U18737 ( .A(n26139), .B(n26138), .Z(n55628) );
  NANDN U18738 ( .A(y[3402]), .B(x[3402]), .Z(n38425) );
  NANDN U18739 ( .A(y[3403]), .B(x[3403]), .Z(n38432) );
  NAND U18740 ( .A(n38425), .B(n38432), .Z(n55626) );
  NANDN U18741 ( .A(x[3401]), .B(y[3401]), .Z(n26143) );
  NANDN U18742 ( .A(x[3402]), .B(y[3402]), .Z(n26142) );
  AND U18743 ( .A(n26143), .B(n26142), .Z(n55625) );
  NANDN U18744 ( .A(y[3400]), .B(x[3400]), .Z(n9896) );
  NANDN U18745 ( .A(y[3401]), .B(x[3401]), .Z(n38426) );
  NAND U18746 ( .A(n9896), .B(n38426), .Z(n55624) );
  XNOR U18747 ( .A(y[3400]), .B(x[3400]), .Z(n38420) );
  NANDN U18748 ( .A(x[3399]), .B(y[3399]), .Z(n26145) );
  AND U18749 ( .A(n38420), .B(n26145), .Z(n55623) );
  NANDN U18750 ( .A(y[3398]), .B(x[3398]), .Z(n9897) );
  NANDN U18751 ( .A(y[3399]), .B(x[3399]), .Z(n38419) );
  NAND U18752 ( .A(n9897), .B(n38419), .Z(n55622) );
  XNOR U18753 ( .A(x[3398]), .B(y[3398]), .Z(n38414) );
  NANDN U18754 ( .A(x[3395]), .B(y[3395]), .Z(n55618) );
  XNOR U18755 ( .A(x[3396]), .B(y[3396]), .Z(n26147) );
  AND U18756 ( .A(n55618), .B(n26147), .Z(n15076) );
  NANDN U18757 ( .A(y[3394]), .B(x[3394]), .Z(n26148) );
  NANDN U18758 ( .A(y[3395]), .B(x[3395]), .Z(n26146) );
  AND U18759 ( .A(n26148), .B(n26146), .Z(n51886) );
  NANDN U18760 ( .A(x[3393]), .B(y[3393]), .Z(n26150) );
  NANDN U18761 ( .A(x[3394]), .B(y[3394]), .Z(n38407) );
  NAND U18762 ( .A(n26150), .B(n38407), .Z(n51887) );
  NANDN U18763 ( .A(y[3392]), .B(x[3392]), .Z(n26152) );
  NANDN U18764 ( .A(y[3393]), .B(x[3393]), .Z(n26149) );
  AND U18765 ( .A(n26152), .B(n26149), .Z(n55615) );
  XNOR U18766 ( .A(x[3390]), .B(y[3390]), .Z(n26154) );
  NANDN U18767 ( .A(y[3386]), .B(x[3386]), .Z(n38386) );
  NANDN U18768 ( .A(y[3387]), .B(x[3387]), .Z(n26159) );
  NAND U18769 ( .A(n38386), .B(n26159), .Z(n55608) );
  NANDN U18770 ( .A(x[3385]), .B(y[3385]), .Z(n26162) );
  NANDN U18771 ( .A(x[3386]), .B(y[3386]), .Z(n26161) );
  NAND U18772 ( .A(n26162), .B(n26161), .Z(n51890) );
  NANDN U18773 ( .A(y[3384]), .B(x[3384]), .Z(n38380) );
  NANDN U18774 ( .A(y[3385]), .B(x[3385]), .Z(n38387) );
  AND U18775 ( .A(n38380), .B(n38387), .Z(n55607) );
  XNOR U18776 ( .A(x[3382]), .B(y[3382]), .Z(n38373) );
  NANDN U18777 ( .A(y[3378]), .B(x[3378]), .Z(n38360) );
  NANDN U18778 ( .A(y[3379]), .B(x[3379]), .Z(n38367) );
  NAND U18779 ( .A(n38360), .B(n38367), .Z(n55599) );
  NANDN U18780 ( .A(x[3377]), .B(y[3377]), .Z(n38356) );
  NANDN U18781 ( .A(x[3378]), .B(y[3378]), .Z(n26166) );
  NAND U18782 ( .A(n38356), .B(n26166), .Z(n55598) );
  NANDN U18783 ( .A(y[3376]), .B(x[3376]), .Z(n38355) );
  NANDN U18784 ( .A(y[3377]), .B(x[3377]), .Z(n38361) );
  AND U18785 ( .A(n38355), .B(n38361), .Z(n51892) );
  NANDN U18786 ( .A(y[3374]), .B(x[3374]), .Z(n38346) );
  ANDN U18787 ( .B(x[3375]), .A(y[3375]), .Z(n38353) );
  ANDN U18788 ( .B(n38346), .A(n38353), .Z(n55597) );
  NANDN U18789 ( .A(x[3373]), .B(y[3373]), .Z(n26169) );
  NANDN U18790 ( .A(x[3374]), .B(y[3374]), .Z(n26168) );
  NAND U18791 ( .A(n26169), .B(n26168), .Z(n55596) );
  NANDN U18792 ( .A(y[3372]), .B(x[3372]), .Z(n38340) );
  NANDN U18793 ( .A(y[3373]), .B(x[3373]), .Z(n38347) );
  NAND U18794 ( .A(n38340), .B(n38347), .Z(n55595) );
  NANDN U18795 ( .A(x[3371]), .B(y[3371]), .Z(n26171) );
  NANDN U18796 ( .A(x[3372]), .B(y[3372]), .Z(n26170) );
  AND U18797 ( .A(n26171), .B(n26170), .Z(n51894) );
  NANDN U18798 ( .A(y[3368]), .B(x[3368]), .Z(n9898) );
  NANDN U18799 ( .A(y[3369]), .B(x[3369]), .Z(n38335) );
  NAND U18800 ( .A(n9898), .B(n38335), .Z(n55593) );
  XNOR U18801 ( .A(y[3368]), .B(x[3368]), .Z(n38329) );
  NANDN U18802 ( .A(x[3367]), .B(y[3367]), .Z(n26175) );
  NAND U18803 ( .A(n38329), .B(n26175), .Z(n55592) );
  NANDN U18804 ( .A(y[3366]), .B(x[3366]), .Z(n38322) );
  NANDN U18805 ( .A(y[3367]), .B(x[3367]), .Z(n38328) );
  AND U18806 ( .A(n38322), .B(n38328), .Z(n51896) );
  NANDN U18807 ( .A(x[3363]), .B(y[3363]), .Z(n26179) );
  NANDN U18808 ( .A(x[3364]), .B(y[3364]), .Z(n26178) );
  NAND U18809 ( .A(n26179), .B(n26178), .Z(n55589) );
  NANDN U18810 ( .A(y[3362]), .B(x[3362]), .Z(n38310) );
  NANDN U18811 ( .A(y[3363]), .B(x[3363]), .Z(n38317) );
  NAND U18812 ( .A(n38310), .B(n38317), .Z(n55588) );
  NANDN U18813 ( .A(x[3361]), .B(y[3361]), .Z(n26181) );
  NANDN U18814 ( .A(x[3362]), .B(y[3362]), .Z(n26180) );
  AND U18815 ( .A(n26181), .B(n26180), .Z(n55587) );
  NANDN U18816 ( .A(y[3360]), .B(x[3360]), .Z(n38304) );
  NANDN U18817 ( .A(y[3361]), .B(x[3361]), .Z(n38311) );
  NAND U18818 ( .A(n38304), .B(n38311), .Z(n55586) );
  NANDN U18819 ( .A(x[3359]), .B(y[3359]), .Z(n26183) );
  NANDN U18820 ( .A(x[3360]), .B(y[3360]), .Z(n26182) );
  AND U18821 ( .A(n26183), .B(n26182), .Z(n55585) );
  NANDN U18822 ( .A(y[3358]), .B(x[3358]), .Z(n38298) );
  NANDN U18823 ( .A(y[3359]), .B(x[3359]), .Z(n38305) );
  NAND U18824 ( .A(n38298), .B(n38305), .Z(n55584) );
  NANDN U18825 ( .A(x[3357]), .B(y[3357]), .Z(n26185) );
  NANDN U18826 ( .A(x[3358]), .B(y[3358]), .Z(n26184) );
  NAND U18827 ( .A(n26185), .B(n26184), .Z(n55583) );
  NANDN U18828 ( .A(y[3356]), .B(x[3356]), .Z(n26187) );
  NANDN U18829 ( .A(y[3357]), .B(x[3357]), .Z(n38299) );
  AND U18830 ( .A(n26187), .B(n38299), .Z(n51898) );
  NANDN U18831 ( .A(y[3352]), .B(x[3352]), .Z(n26191) );
  NANDN U18832 ( .A(y[3353]), .B(x[3353]), .Z(n26189) );
  NAND U18833 ( .A(n26191), .B(n26189), .Z(n51902) );
  NANDN U18834 ( .A(x[3351]), .B(y[3351]), .Z(n26193) );
  NANDN U18835 ( .A(x[3352]), .B(y[3352]), .Z(n38287) );
  AND U18836 ( .A(n26193), .B(n38287), .Z(n51903) );
  NANDN U18837 ( .A(y[3348]), .B(x[3348]), .Z(n26197) );
  NANDN U18838 ( .A(y[3349]), .B(x[3349]), .Z(n26196) );
  NAND U18839 ( .A(n26197), .B(n26196), .Z(n55578) );
  NANDN U18840 ( .A(x[3347]), .B(y[3347]), .Z(n26199) );
  NANDN U18841 ( .A(x[3348]), .B(y[3348]), .Z(n38279) );
  NAND U18842 ( .A(n26199), .B(n38279), .Z(n55577) );
  NANDN U18843 ( .A(y[3346]), .B(x[3346]), .Z(n9899) );
  NANDN U18844 ( .A(y[3347]), .B(x[3347]), .Z(n26198) );
  AND U18845 ( .A(n9899), .B(n26198), .Z(n55576) );
  XNOR U18846 ( .A(y[3346]), .B(x[3346]), .Z(n38270) );
  NANDN U18847 ( .A(x[3345]), .B(y[3345]), .Z(n26201) );
  NAND U18848 ( .A(n38270), .B(n26201), .Z(n55575) );
  NANDN U18849 ( .A(y[3344]), .B(x[3344]), .Z(n55573) );
  ANDN U18850 ( .B(x[3345]), .A(y[3345]), .Z(n55574) );
  ANDN U18851 ( .B(n55573), .A(n55574), .Z(n15018) );
  NANDN U18852 ( .A(y[3342]), .B(x[3342]), .Z(n26203) );
  NANDN U18853 ( .A(y[3343]), .B(x[3343]), .Z(n38265) );
  NAND U18854 ( .A(n26203), .B(n38265), .Z(n51907) );
  NANDN U18855 ( .A(x[3341]), .B(y[3341]), .Z(n26206) );
  NANDN U18856 ( .A(x[3342]), .B(y[3342]), .Z(n26202) );
  AND U18857 ( .A(n26206), .B(n26202), .Z(n55570) );
  NANDN U18858 ( .A(y[3338]), .B(x[3338]), .Z(n38250) );
  NANDN U18859 ( .A(y[3339]), .B(x[3339]), .Z(n26208) );
  NAND U18860 ( .A(n38250), .B(n26208), .Z(n55568) );
  NANDN U18861 ( .A(x[3337]), .B(y[3337]), .Z(n26211) );
  NANDN U18862 ( .A(x[3338]), .B(y[3338]), .Z(n26210) );
  NAND U18863 ( .A(n26211), .B(n26210), .Z(n51909) );
  NANDN U18864 ( .A(y[3336]), .B(x[3336]), .Z(n38244) );
  NANDN U18865 ( .A(y[3337]), .B(x[3337]), .Z(n38251) );
  AND U18866 ( .A(n38244), .B(n38251), .Z(n55567) );
  NANDN U18867 ( .A(x[3333]), .B(y[3333]), .Z(n26215) );
  XNOR U18868 ( .A(x[3334]), .B(y[3334]), .Z(n9900) );
  NAND U18869 ( .A(n26215), .B(n9900), .Z(n51911) );
  NANDN U18870 ( .A(y[3332]), .B(x[3332]), .Z(n9901) );
  NANDN U18871 ( .A(y[3333]), .B(x[3333]), .Z(n38239) );
  NAND U18872 ( .A(n9901), .B(n38239), .Z(n55565) );
  XNOR U18873 ( .A(y[3332]), .B(x[3332]), .Z(n38233) );
  NANDN U18874 ( .A(x[3331]), .B(y[3331]), .Z(n26217) );
  AND U18875 ( .A(n38233), .B(n26217), .Z(n55563) );
  NANDN U18876 ( .A(y[3330]), .B(x[3330]), .Z(n38226) );
  NANDN U18877 ( .A(y[3331]), .B(x[3331]), .Z(n38232) );
  NAND U18878 ( .A(n38226), .B(n38232), .Z(n55562) );
  NANDN U18879 ( .A(x[3329]), .B(y[3329]), .Z(n26219) );
  NANDN U18880 ( .A(x[3330]), .B(y[3330]), .Z(n26218) );
  AND U18881 ( .A(n26219), .B(n26218), .Z(n55561) );
  NANDN U18882 ( .A(y[3328]), .B(x[3328]), .Z(n9902) );
  NANDN U18883 ( .A(y[3329]), .B(x[3329]), .Z(n38227) );
  NAND U18884 ( .A(n9902), .B(n38227), .Z(n55560) );
  XNOR U18885 ( .A(y[3328]), .B(x[3328]), .Z(n38221) );
  NANDN U18886 ( .A(x[3327]), .B(y[3327]), .Z(n38216) );
  NAND U18887 ( .A(n38221), .B(n38216), .Z(n51912) );
  NANDN U18888 ( .A(y[3326]), .B(x[3326]), .Z(n38215) );
  NANDN U18889 ( .A(y[3327]), .B(x[3327]), .Z(n38220) );
  AND U18890 ( .A(n38215), .B(n38220), .Z(n55559) );
  NANDN U18891 ( .A(y[3324]), .B(x[3324]), .Z(n38206) );
  ANDN U18892 ( .B(x[3325]), .A(y[3325]), .Z(n38213) );
  ANDN U18893 ( .B(n38206), .A(n38213), .Z(n55557) );
  NANDN U18894 ( .A(x[3323]), .B(y[3323]), .Z(n26223) );
  NANDN U18895 ( .A(x[3324]), .B(y[3324]), .Z(n26222) );
  NAND U18896 ( .A(n26223), .B(n26222), .Z(n55556) );
  NANDN U18897 ( .A(y[3322]), .B(x[3322]), .Z(n38200) );
  NANDN U18898 ( .A(y[3323]), .B(x[3323]), .Z(n38207) );
  NAND U18899 ( .A(n38200), .B(n38207), .Z(n51913) );
  NANDN U18900 ( .A(x[3321]), .B(y[3321]), .Z(n26225) );
  NANDN U18901 ( .A(x[3322]), .B(y[3322]), .Z(n26224) );
  AND U18902 ( .A(n26225), .B(n26224), .Z(n55555) );
  NANDN U18903 ( .A(y[3318]), .B(x[3318]), .Z(n38188) );
  NANDN U18904 ( .A(y[3319]), .B(x[3319]), .Z(n38195) );
  NAND U18905 ( .A(n38188), .B(n38195), .Z(n55552) );
  NANDN U18906 ( .A(x[3317]), .B(y[3317]), .Z(n26229) );
  NANDN U18907 ( .A(x[3318]), .B(y[3318]), .Z(n26228) );
  NAND U18908 ( .A(n26229), .B(n26228), .Z(n51915) );
  NANDN U18909 ( .A(y[3316]), .B(x[3316]), .Z(n38182) );
  NANDN U18910 ( .A(y[3317]), .B(x[3317]), .Z(n38189) );
  AND U18911 ( .A(n38182), .B(n38189), .Z(n55551) );
  NANDN U18912 ( .A(x[3313]), .B(y[3313]), .Z(n26233) );
  NANDN U18913 ( .A(x[3314]), .B(y[3314]), .Z(n26232) );
  NAND U18914 ( .A(n26233), .B(n26232), .Z(n55549) );
  NANDN U18915 ( .A(y[3312]), .B(x[3312]), .Z(n38170) );
  NANDN U18916 ( .A(y[3313]), .B(x[3313]), .Z(n38177) );
  NAND U18917 ( .A(n38170), .B(n38177), .Z(n51917) );
  NANDN U18918 ( .A(x[3311]), .B(y[3311]), .Z(n26235) );
  NANDN U18919 ( .A(x[3312]), .B(y[3312]), .Z(n26234) );
  AND U18920 ( .A(n26235), .B(n26234), .Z(n55548) );
  NANDN U18921 ( .A(y[3308]), .B(x[3308]), .Z(n38158) );
  NANDN U18922 ( .A(y[3309]), .B(x[3309]), .Z(n38165) );
  NAND U18923 ( .A(n38158), .B(n38165), .Z(n55546) );
  NANDN U18924 ( .A(x[3307]), .B(y[3307]), .Z(n26239) );
  NANDN U18925 ( .A(x[3308]), .B(y[3308]), .Z(n26238) );
  NAND U18926 ( .A(n26239), .B(n26238), .Z(n51919) );
  NANDN U18927 ( .A(y[3306]), .B(x[3306]), .Z(n38152) );
  NANDN U18928 ( .A(y[3307]), .B(x[3307]), .Z(n38159) );
  AND U18929 ( .A(n38152), .B(n38159), .Z(n55543) );
  NANDN U18930 ( .A(y[3302]), .B(x[3302]), .Z(n38140) );
  NANDN U18931 ( .A(y[3303]), .B(x[3303]), .Z(n38146) );
  NAND U18932 ( .A(n38140), .B(n38146), .Z(n55539) );
  NANDN U18933 ( .A(x[3301]), .B(y[3301]), .Z(n26243) );
  NANDN U18934 ( .A(x[3302]), .B(y[3302]), .Z(n26242) );
  AND U18935 ( .A(n26243), .B(n26242), .Z(n51921) );
  NANDN U18936 ( .A(y[3300]), .B(x[3300]), .Z(n9903) );
  NANDN U18937 ( .A(y[3301]), .B(x[3301]), .Z(n38141) );
  NAND U18938 ( .A(n9903), .B(n38141), .Z(n55538) );
  XNOR U18939 ( .A(y[3300]), .B(x[3300]), .Z(n38135) );
  NANDN U18940 ( .A(x[3299]), .B(y[3299]), .Z(n26245) );
  AND U18941 ( .A(n38135), .B(n26245), .Z(n55537) );
  NANDN U18942 ( .A(y[3298]), .B(x[3298]), .Z(n38128) );
  NANDN U18943 ( .A(y[3299]), .B(x[3299]), .Z(n38134) );
  NAND U18944 ( .A(n38128), .B(n38134), .Z(n55536) );
  NANDN U18945 ( .A(x[3297]), .B(y[3297]), .Z(n26247) );
  NANDN U18946 ( .A(x[3298]), .B(y[3298]), .Z(n26246) );
  NAND U18947 ( .A(n26247), .B(n26246), .Z(n55535) );
  NANDN U18948 ( .A(y[3296]), .B(x[3296]), .Z(n38122) );
  NANDN U18949 ( .A(y[3297]), .B(x[3297]), .Z(n38129) );
  AND U18950 ( .A(n38122), .B(n38129), .Z(n51922) );
  NANDN U18951 ( .A(x[3295]), .B(y[3295]), .Z(n26249) );
  NANDN U18952 ( .A(x[3296]), .B(y[3296]), .Z(n26248) );
  NAND U18953 ( .A(n26249), .B(n26248), .Z(n55534) );
  NANDN U18954 ( .A(y[3294]), .B(x[3294]), .Z(n38116) );
  NANDN U18955 ( .A(y[3295]), .B(x[3295]), .Z(n38123) );
  AND U18956 ( .A(n38116), .B(n38123), .Z(n55532) );
  NANDN U18957 ( .A(x[3293]), .B(y[3293]), .Z(n26251) );
  NANDN U18958 ( .A(x[3294]), .B(y[3294]), .Z(n26250) );
  NAND U18959 ( .A(n26251), .B(n26250), .Z(n55531) );
  NANDN U18960 ( .A(y[3292]), .B(x[3292]), .Z(n38110) );
  NANDN U18961 ( .A(y[3293]), .B(x[3293]), .Z(n38117) );
  NAND U18962 ( .A(n38110), .B(n38117), .Z(n55530) );
  NANDN U18963 ( .A(x[3291]), .B(y[3291]), .Z(n26253) );
  NANDN U18964 ( .A(x[3292]), .B(y[3292]), .Z(n26252) );
  AND U18965 ( .A(n26253), .B(n26252), .Z(n51923) );
  NANDN U18966 ( .A(y[3290]), .B(x[3290]), .Z(n38104) );
  NANDN U18967 ( .A(y[3291]), .B(x[3291]), .Z(n38111) );
  NAND U18968 ( .A(n38104), .B(n38111), .Z(n55529) );
  NANDN U18969 ( .A(x[3289]), .B(y[3289]), .Z(n26255) );
  NANDN U18970 ( .A(x[3290]), .B(y[3290]), .Z(n26254) );
  AND U18971 ( .A(n26255), .B(n26254), .Z(n55528) );
  NANDN U18972 ( .A(y[3288]), .B(x[3288]), .Z(n9904) );
  NANDN U18973 ( .A(y[3289]), .B(x[3289]), .Z(n38105) );
  NAND U18974 ( .A(n9904), .B(n38105), .Z(n55527) );
  XNOR U18975 ( .A(y[3288]), .B(x[3288]), .Z(n38099) );
  NANDN U18976 ( .A(x[3287]), .B(y[3287]), .Z(n26257) );
  NAND U18977 ( .A(n38099), .B(n26257), .Z(n55526) );
  NANDN U18978 ( .A(y[3286]), .B(x[3286]), .Z(n38092) );
  NANDN U18979 ( .A(y[3287]), .B(x[3287]), .Z(n38098) );
  AND U18980 ( .A(n38092), .B(n38098), .Z(n51924) );
  NANDN U18981 ( .A(x[3285]), .B(y[3285]), .Z(n26259) );
  NANDN U18982 ( .A(x[3286]), .B(y[3286]), .Z(n26258) );
  NAND U18983 ( .A(n26259), .B(n26258), .Z(n55525) );
  NANDN U18984 ( .A(y[3284]), .B(x[3284]), .Z(n9905) );
  NANDN U18985 ( .A(y[3285]), .B(x[3285]), .Z(n38093) );
  AND U18986 ( .A(n9905), .B(n38093), .Z(n55524) );
  XNOR U18987 ( .A(y[3284]), .B(x[3284]), .Z(n38087) );
  NANDN U18988 ( .A(x[3283]), .B(y[3283]), .Z(n26261) );
  NAND U18989 ( .A(n38087), .B(n26261), .Z(n55523) );
  NANDN U18990 ( .A(y[3282]), .B(x[3282]), .Z(n9906) );
  NANDN U18991 ( .A(y[3283]), .B(x[3283]), .Z(n38086) );
  NAND U18992 ( .A(n9906), .B(n38086), .Z(n55522) );
  XNOR U18993 ( .A(y[3282]), .B(x[3282]), .Z(n38081) );
  NANDN U18994 ( .A(x[3281]), .B(y[3281]), .Z(n26263) );
  AND U18995 ( .A(n38081), .B(n26263), .Z(n51925) );
  NANDN U18996 ( .A(y[3280]), .B(x[3280]), .Z(n38074) );
  NANDN U18997 ( .A(y[3281]), .B(x[3281]), .Z(n38080) );
  NAND U18998 ( .A(n38074), .B(n38080), .Z(n55520) );
  NANDN U18999 ( .A(x[3279]), .B(y[3279]), .Z(n26265) );
  NANDN U19000 ( .A(x[3280]), .B(y[3280]), .Z(n26264) );
  AND U19001 ( .A(n26265), .B(n26264), .Z(n55519) );
  NANDN U19002 ( .A(y[3278]), .B(x[3278]), .Z(n38068) );
  NANDN U19003 ( .A(y[3279]), .B(x[3279]), .Z(n38075) );
  NAND U19004 ( .A(n38068), .B(n38075), .Z(n55518) );
  NANDN U19005 ( .A(x[3277]), .B(y[3277]), .Z(n26267) );
  NANDN U19006 ( .A(x[3278]), .B(y[3278]), .Z(n26266) );
  NAND U19007 ( .A(n26267), .B(n26266), .Z(n55517) );
  NANDN U19008 ( .A(y[3276]), .B(x[3276]), .Z(n38062) );
  NANDN U19009 ( .A(y[3277]), .B(x[3277]), .Z(n38069) );
  AND U19010 ( .A(n38062), .B(n38069), .Z(n51926) );
  NANDN U19011 ( .A(x[3275]), .B(y[3275]), .Z(n26269) );
  NANDN U19012 ( .A(x[3276]), .B(y[3276]), .Z(n26268) );
  NAND U19013 ( .A(n26269), .B(n26268), .Z(n55516) );
  NANDN U19014 ( .A(y[3274]), .B(x[3274]), .Z(n38056) );
  NANDN U19015 ( .A(y[3275]), .B(x[3275]), .Z(n38063) );
  AND U19016 ( .A(n38056), .B(n38063), .Z(n55515) );
  NANDN U19017 ( .A(x[3273]), .B(y[3273]), .Z(n38052) );
  NANDN U19018 ( .A(x[3274]), .B(y[3274]), .Z(n26270) );
  NAND U19019 ( .A(n38052), .B(n26270), .Z(n55514) );
  NANDN U19020 ( .A(y[3272]), .B(x[3272]), .Z(n26271) );
  NANDN U19021 ( .A(y[3273]), .B(x[3273]), .Z(n38057) );
  NAND U19022 ( .A(n26271), .B(n38057), .Z(n55513) );
  NANDN U19023 ( .A(x[3271]), .B(y[3271]), .Z(n26273) );
  NANDN U19024 ( .A(x[3272]), .B(y[3272]), .Z(n38053) );
  AND U19025 ( .A(n26273), .B(n38053), .Z(n51927) );
  NANDN U19026 ( .A(y[3270]), .B(x[3270]), .Z(n26275) );
  NANDN U19027 ( .A(y[3271]), .B(x[3271]), .Z(n26272) );
  NAND U19028 ( .A(n26275), .B(n26272), .Z(n55512) );
  NANDN U19029 ( .A(x[3269]), .B(y[3269]), .Z(n26277) );
  NANDN U19030 ( .A(x[3270]), .B(y[3270]), .Z(n26274) );
  AND U19031 ( .A(n26277), .B(n26274), .Z(n55511) );
  NANDN U19032 ( .A(y[3268]), .B(x[3268]), .Z(n9907) );
  NANDN U19033 ( .A(y[3269]), .B(x[3269]), .Z(n26276) );
  NAND U19034 ( .A(n9907), .B(n26276), .Z(n55510) );
  NANDN U19035 ( .A(y[3266]), .B(x[3266]), .Z(n38036) );
  NANDN U19036 ( .A(y[3267]), .B(x[3267]), .Z(n26278) );
  AND U19037 ( .A(n38036), .B(n26278), .Z(n55509) );
  NANDN U19038 ( .A(x[3265]), .B(y[3265]), .Z(n26281) );
  NANDN U19039 ( .A(x[3266]), .B(y[3266]), .Z(n26280) );
  NAND U19040 ( .A(n26281), .B(n26280), .Z(n55507) );
  NANDN U19041 ( .A(y[3264]), .B(x[3264]), .Z(n38030) );
  NANDN U19042 ( .A(y[3265]), .B(x[3265]), .Z(n38037) );
  NAND U19043 ( .A(n38030), .B(n38037), .Z(n51930) );
  NANDN U19044 ( .A(x[3263]), .B(y[3263]), .Z(n26283) );
  NANDN U19045 ( .A(x[3264]), .B(y[3264]), .Z(n26282) );
  AND U19046 ( .A(n26283), .B(n26282), .Z(n55506) );
  NANDN U19047 ( .A(y[3260]), .B(x[3260]), .Z(n38018) );
  NANDN U19048 ( .A(y[3261]), .B(x[3261]), .Z(n38025) );
  NAND U19049 ( .A(n38018), .B(n38025), .Z(n55503) );
  NANDN U19050 ( .A(x[3259]), .B(y[3259]), .Z(n26287) );
  NANDN U19051 ( .A(x[3260]), .B(y[3260]), .Z(n26286) );
  NAND U19052 ( .A(n26287), .B(n26286), .Z(n55502) );
  NANDN U19053 ( .A(y[3258]), .B(x[3258]), .Z(n38012) );
  NANDN U19054 ( .A(y[3259]), .B(x[3259]), .Z(n38019) );
  AND U19055 ( .A(n38012), .B(n38019), .Z(n55501) );
  NANDN U19056 ( .A(x[3255]), .B(y[3255]), .Z(n26291) );
  NANDN U19057 ( .A(x[3256]), .B(y[3256]), .Z(n26290) );
  NAND U19058 ( .A(n26291), .B(n26290), .Z(n55499) );
  NANDN U19059 ( .A(y[3254]), .B(x[3254]), .Z(n9908) );
  NANDN U19060 ( .A(y[3255]), .B(x[3255]), .Z(n38007) );
  NAND U19061 ( .A(n9908), .B(n38007), .Z(n51932) );
  XNOR U19062 ( .A(y[3254]), .B(x[3254]), .Z(n38001) );
  NANDN U19063 ( .A(x[3253]), .B(y[3253]), .Z(n37997) );
  AND U19064 ( .A(n38001), .B(n37997), .Z(n55497) );
  NANDN U19065 ( .A(y[3250]), .B(x[3250]), .Z(n26295) );
  NANDN U19066 ( .A(y[3251]), .B(x[3251]), .Z(n26294) );
  NAND U19067 ( .A(n26295), .B(n26294), .Z(n55495) );
  NANDN U19068 ( .A(x[3249]), .B(y[3249]), .Z(n37985) );
  NANDN U19069 ( .A(x[3250]), .B(y[3250]), .Z(n37992) );
  NAND U19070 ( .A(n37985), .B(n37992), .Z(n51934) );
  NANDN U19071 ( .A(y[3248]), .B(x[3248]), .Z(n26297) );
  NANDN U19072 ( .A(y[3249]), .B(x[3249]), .Z(n26296) );
  AND U19073 ( .A(n26297), .B(n26296), .Z(n55494) );
  NANDN U19074 ( .A(x[3245]), .B(y[3245]), .Z(n37977) );
  NANDN U19075 ( .A(x[3246]), .B(y[3246]), .Z(n26300) );
  NAND U19076 ( .A(n37977), .B(n26300), .Z(n55492) );
  NANDN U19077 ( .A(y[3244]), .B(x[3244]), .Z(n26303) );
  NANDN U19078 ( .A(y[3245]), .B(x[3245]), .Z(n26302) );
  NAND U19079 ( .A(n26303), .B(n26302), .Z(n51936) );
  NANDN U19080 ( .A(x[3243]), .B(y[3243]), .Z(n37968) );
  ANDN U19081 ( .B(y[3244]), .A(x[3244]), .Z(n37975) );
  ANDN U19082 ( .B(n37968), .A(n37975), .Z(n55491) );
  NANDN U19083 ( .A(y[3240]), .B(x[3240]), .Z(n37959) );
  NANDN U19084 ( .A(y[3241]), .B(x[3241]), .Z(n26306) );
  NAND U19085 ( .A(n37959), .B(n26306), .Z(n51938) );
  NANDN U19086 ( .A(x[3239]), .B(y[3239]), .Z(n26307) );
  NANDN U19087 ( .A(x[3240]), .B(y[3240]), .Z(n37963) );
  NAND U19088 ( .A(n26307), .B(n37963), .Z(n55487) );
  NANDN U19089 ( .A(y[3238]), .B(x[3238]), .Z(n37953) );
  NANDN U19090 ( .A(y[3239]), .B(x[3239]), .Z(n37960) );
  AND U19091 ( .A(n37953), .B(n37960), .Z(n55486) );
  NANDN U19092 ( .A(x[3237]), .B(y[3237]), .Z(n26309) );
  NANDN U19093 ( .A(x[3238]), .B(y[3238]), .Z(n26308) );
  NAND U19094 ( .A(n26309), .B(n26308), .Z(n55485) );
  NANDN U19095 ( .A(y[3236]), .B(x[3236]), .Z(n37947) );
  NANDN U19096 ( .A(y[3237]), .B(x[3237]), .Z(n37954) );
  AND U19097 ( .A(n37947), .B(n37954), .Z(n55484) );
  NANDN U19098 ( .A(x[3235]), .B(y[3235]), .Z(n26311) );
  NANDN U19099 ( .A(x[3236]), .B(y[3236]), .Z(n26310) );
  NAND U19100 ( .A(n26311), .B(n26310), .Z(n55483) );
  NANDN U19101 ( .A(y[3234]), .B(x[3234]), .Z(n37941) );
  NANDN U19102 ( .A(y[3235]), .B(x[3235]), .Z(n37948) );
  NAND U19103 ( .A(n37941), .B(n37948), .Z(n51939) );
  NANDN U19104 ( .A(x[3234]), .B(y[3234]), .Z(n26312) );
  ANDN U19105 ( .B(y[3233]), .A(x[3233]), .Z(n37939) );
  ANDN U19106 ( .B(n26312), .A(n37939), .Z(n55482) );
  NANDN U19107 ( .A(x[3231]), .B(y[3231]), .Z(n55479) );
  XNOR U19108 ( .A(x[3232]), .B(y[3232]), .Z(n26314) );
  AND U19109 ( .A(n55479), .B(n26314), .Z(n14897) );
  NANDN U19110 ( .A(y[3230]), .B(x[3230]), .Z(n26316) );
  NANDN U19111 ( .A(y[3231]), .B(x[3231]), .Z(n26313) );
  AND U19112 ( .A(n26316), .B(n26313), .Z(n55478) );
  NANDN U19113 ( .A(x[3229]), .B(y[3229]), .Z(n26318) );
  NANDN U19114 ( .A(x[3230]), .B(y[3230]), .Z(n26315) );
  NAND U19115 ( .A(n26318), .B(n26315), .Z(n55476) );
  NANDN U19116 ( .A(y[3228]), .B(x[3228]), .Z(n9909) );
  NANDN U19117 ( .A(y[3229]), .B(x[3229]), .Z(n26317) );
  AND U19118 ( .A(n9909), .B(n26317), .Z(n51940) );
  NANDN U19119 ( .A(x[3227]), .B(y[3227]), .Z(n55472) );
  NANDN U19120 ( .A(y[3226]), .B(x[3226]), .Z(n37919) );
  NANDN U19121 ( .A(y[3227]), .B(x[3227]), .Z(n37925) );
  AND U19122 ( .A(n37919), .B(n37925), .Z(n55471) );
  NANDN U19123 ( .A(x[3225]), .B(y[3225]), .Z(n26320) );
  NANDN U19124 ( .A(x[3226]), .B(y[3226]), .Z(n26319) );
  NAND U19125 ( .A(n26320), .B(n26319), .Z(n55470) );
  NANDN U19126 ( .A(y[3224]), .B(x[3224]), .Z(n37913) );
  NANDN U19127 ( .A(y[3225]), .B(x[3225]), .Z(n37920) );
  AND U19128 ( .A(n37913), .B(n37920), .Z(n55469) );
  NANDN U19129 ( .A(x[3223]), .B(y[3223]), .Z(n26322) );
  NANDN U19130 ( .A(x[3224]), .B(y[3224]), .Z(n26321) );
  NAND U19131 ( .A(n26322), .B(n26321), .Z(n55468) );
  NANDN U19132 ( .A(y[3222]), .B(x[3222]), .Z(n37907) );
  NANDN U19133 ( .A(y[3223]), .B(x[3223]), .Z(n37914) );
  AND U19134 ( .A(n37907), .B(n37914), .Z(n51941) );
  XNOR U19135 ( .A(y[3220]), .B(x[3220]), .Z(n37902) );
  NANDN U19136 ( .A(x[3219]), .B(y[3219]), .Z(n26326) );
  NAND U19137 ( .A(n37902), .B(n26326), .Z(n55466) );
  NANDN U19138 ( .A(y[3218]), .B(x[3218]), .Z(n37895) );
  NANDN U19139 ( .A(y[3219]), .B(x[3219]), .Z(n37901) );
  NAND U19140 ( .A(n37895), .B(n37901), .Z(n55465) );
  NANDN U19141 ( .A(x[3217]), .B(y[3217]), .Z(n26328) );
  NANDN U19142 ( .A(x[3218]), .B(y[3218]), .Z(n26327) );
  AND U19143 ( .A(n26328), .B(n26327), .Z(n51943) );
  NANDN U19144 ( .A(y[3214]), .B(x[3214]), .Z(n9910) );
  NANDN U19145 ( .A(y[3215]), .B(x[3215]), .Z(n37889) );
  NAND U19146 ( .A(n9910), .B(n37889), .Z(n55462) );
  XNOR U19147 ( .A(y[3214]), .B(x[3214]), .Z(n37884) );
  NANDN U19148 ( .A(x[3213]), .B(y[3213]), .Z(n26332) );
  NAND U19149 ( .A(n37884), .B(n26332), .Z(n55461) );
  NANDN U19150 ( .A(y[3212]), .B(x[3212]), .Z(n9911) );
  NANDN U19151 ( .A(y[3213]), .B(x[3213]), .Z(n37883) );
  AND U19152 ( .A(n9911), .B(n37883), .Z(n51945) );
  NANDN U19153 ( .A(x[3209]), .B(y[3209]), .Z(n26336) );
  NANDN U19154 ( .A(x[3210]), .B(y[3210]), .Z(n26335) );
  NAND U19155 ( .A(n26336), .B(n26335), .Z(n55459) );
  NANDN U19156 ( .A(y[3208]), .B(x[3208]), .Z(n37865) );
  NANDN U19157 ( .A(y[3209]), .B(x[3209]), .Z(n37872) );
  AND U19158 ( .A(n37865), .B(n37872), .Z(n51947) );
  NANDN U19159 ( .A(x[3207]), .B(y[3207]), .Z(n26338) );
  NANDN U19160 ( .A(x[3208]), .B(y[3208]), .Z(n26337) );
  NAND U19161 ( .A(n26338), .B(n26337), .Z(n55458) );
  NANDN U19162 ( .A(y[3206]), .B(x[3206]), .Z(n37859) );
  NANDN U19163 ( .A(y[3207]), .B(x[3207]), .Z(n37866) );
  AND U19164 ( .A(n37859), .B(n37866), .Z(n55457) );
  NANDN U19165 ( .A(x[3205]), .B(y[3205]), .Z(n26340) );
  NANDN U19166 ( .A(x[3206]), .B(y[3206]), .Z(n26339) );
  NAND U19167 ( .A(n26340), .B(n26339), .Z(n55456) );
  NANDN U19168 ( .A(y[3204]), .B(x[3204]), .Z(n37853) );
  NANDN U19169 ( .A(y[3205]), .B(x[3205]), .Z(n37860) );
  AND U19170 ( .A(n37853), .B(n37860), .Z(n55455) );
  NANDN U19171 ( .A(x[3203]), .B(y[3203]), .Z(n26342) );
  NANDN U19172 ( .A(x[3204]), .B(y[3204]), .Z(n26341) );
  NAND U19173 ( .A(n26342), .B(n26341), .Z(n55454) );
  NANDN U19174 ( .A(y[3202]), .B(x[3202]), .Z(n37847) );
  NANDN U19175 ( .A(y[3203]), .B(x[3203]), .Z(n37854) );
  AND U19176 ( .A(n37847), .B(n37854), .Z(n51948) );
  XNOR U19177 ( .A(x[3200]), .B(y[3200]), .Z(n37842) );
  NANDN U19178 ( .A(y[3196]), .B(x[3196]), .Z(n26349) );
  NANDN U19179 ( .A(y[3197]), .B(x[3197]), .Z(n26348) );
  NAND U19180 ( .A(n26349), .B(n26348), .Z(n51953) );
  NANDN U19181 ( .A(x[3195]), .B(y[3195]), .Z(n37828) );
  NANDN U19182 ( .A(x[3196]), .B(y[3196]), .Z(n37835) );
  NAND U19183 ( .A(n37828), .B(n37835), .Z(n55450) );
  NANDN U19184 ( .A(y[3194]), .B(x[3194]), .Z(n37824) );
  NANDN U19185 ( .A(y[3195]), .B(x[3195]), .Z(n26350) );
  AND U19186 ( .A(n37824), .B(n26350), .Z(n55449) );
  NANDN U19187 ( .A(x[3193]), .B(y[3193]), .Z(n26352) );
  NANDN U19188 ( .A(x[3194]), .B(y[3194]), .Z(n37829) );
  NAND U19189 ( .A(n26352), .B(n37829), .Z(n55448) );
  NANDN U19190 ( .A(y[3192]), .B(x[3192]), .Z(n51955) );
  NANDN U19191 ( .A(y[3193]), .B(x[3193]), .Z(n51954) );
  AND U19192 ( .A(n51955), .B(n51954), .Z(n14852) );
  ANDN U19193 ( .B(y[3189]), .A(x[3189]), .Z(n26356) );
  XNOR U19194 ( .A(x[3190]), .B(y[3190]), .Z(n26354) );
  NANDN U19195 ( .A(y[3186]), .B(x[3186]), .Z(n26360) );
  NANDN U19196 ( .A(y[3187]), .B(x[3187]), .Z(n26359) );
  NAND U19197 ( .A(n26360), .B(n26359), .Z(n51960) );
  NANDN U19198 ( .A(y[3184]), .B(x[3184]), .Z(n37797) );
  NANDN U19199 ( .A(y[3185]), .B(x[3185]), .Z(n26361) );
  AND U19200 ( .A(n37797), .B(n26361), .Z(n55442) );
  NANDN U19201 ( .A(x[3183]), .B(y[3183]), .Z(n26362) );
  NANDN U19202 ( .A(x[3184]), .B(y[3184]), .Z(n37802) );
  NAND U19203 ( .A(n26362), .B(n37802), .Z(n55441) );
  NANDN U19204 ( .A(y[3182]), .B(x[3182]), .Z(n26364) );
  NANDN U19205 ( .A(y[3183]), .B(x[3183]), .Z(n37798) );
  NAND U19206 ( .A(n26364), .B(n37798), .Z(n55440) );
  NANDN U19207 ( .A(x[3181]), .B(y[3181]), .Z(n26366) );
  NANDN U19208 ( .A(x[3182]), .B(y[3182]), .Z(n26363) );
  AND U19209 ( .A(n26366), .B(n26363), .Z(n55439) );
  NANDN U19210 ( .A(y[3180]), .B(x[3180]), .Z(n26369) );
  NANDN U19211 ( .A(y[3181]), .B(x[3181]), .Z(n26365) );
  NAND U19212 ( .A(n26369), .B(n26365), .Z(n55438) );
  NANDN U19213 ( .A(x[3180]), .B(y[3180]), .Z(n26367) );
  ANDN U19214 ( .B(y[3179]), .A(x[3179]), .Z(n37786) );
  ANDN U19215 ( .B(n26367), .A(n37786), .Z(n55437) );
  NANDN U19216 ( .A(y[3178]), .B(x[3178]), .Z(n9912) );
  NANDN U19217 ( .A(y[3179]), .B(x[3179]), .Z(n26368) );
  NAND U19218 ( .A(n9912), .B(n26368), .Z(n55436) );
  XNOR U19219 ( .A(y[3178]), .B(x[3178]), .Z(n26371) );
  NANDN U19220 ( .A(x[3177]), .B(y[3177]), .Z(n26372) );
  NAND U19221 ( .A(n26371), .B(n26372), .Z(n55434) );
  NANDN U19222 ( .A(y[3176]), .B(x[3176]), .Z(n9913) );
  NANDN U19223 ( .A(y[3177]), .B(x[3177]), .Z(n26370) );
  AND U19224 ( .A(n9913), .B(n26370), .Z(n55433) );
  XNOR U19225 ( .A(y[3176]), .B(x[3176]), .Z(n26375) );
  NANDN U19226 ( .A(x[3175]), .B(y[3175]), .Z(n37775) );
  NAND U19227 ( .A(n26375), .B(n37775), .Z(n55432) );
  NANDN U19228 ( .A(y[3174]), .B(x[3174]), .Z(n26376) );
  NANDN U19229 ( .A(y[3175]), .B(x[3175]), .Z(n26374) );
  AND U19230 ( .A(n26376), .B(n26374), .Z(n55431) );
  NANDN U19231 ( .A(x[3173]), .B(y[3173]), .Z(n37769) );
  NANDN U19232 ( .A(x[3174]), .B(y[3174]), .Z(n37776) );
  NAND U19233 ( .A(n37769), .B(n37776), .Z(n55430) );
  NANDN U19234 ( .A(y[3172]), .B(x[3172]), .Z(n26378) );
  NANDN U19235 ( .A(y[3173]), .B(x[3173]), .Z(n26377) );
  NAND U19236 ( .A(n26378), .B(n26377), .Z(n55429) );
  NANDN U19237 ( .A(x[3171]), .B(y[3171]), .Z(n37763) );
  NANDN U19238 ( .A(x[3172]), .B(y[3172]), .Z(n37770) );
  AND U19239 ( .A(n37763), .B(n37770), .Z(n55428) );
  NANDN U19240 ( .A(y[3170]), .B(x[3170]), .Z(n37760) );
  NANDN U19241 ( .A(y[3171]), .B(x[3171]), .Z(n26379) );
  NAND U19242 ( .A(n37760), .B(n26379), .Z(n55427) );
  NANDN U19243 ( .A(x[3169]), .B(y[3169]), .Z(n26380) );
  NANDN U19244 ( .A(x[3170]), .B(y[3170]), .Z(n37764) );
  AND U19245 ( .A(n26380), .B(n37764), .Z(n55426) );
  NANDN U19246 ( .A(y[3168]), .B(x[3168]), .Z(n37754) );
  NANDN U19247 ( .A(y[3169]), .B(x[3169]), .Z(n37761) );
  NAND U19248 ( .A(n37754), .B(n37761), .Z(n55425) );
  NANDN U19249 ( .A(x[3167]), .B(y[3167]), .Z(n26382) );
  NANDN U19250 ( .A(x[3168]), .B(y[3168]), .Z(n26381) );
  NAND U19251 ( .A(n26382), .B(n26381), .Z(n55424) );
  NANDN U19252 ( .A(y[3166]), .B(x[3166]), .Z(n37748) );
  NANDN U19253 ( .A(y[3167]), .B(x[3167]), .Z(n37755) );
  AND U19254 ( .A(n37748), .B(n37755), .Z(n55423) );
  ANDN U19255 ( .B(y[3165]), .A(x[3165]), .Z(n37746) );
  NANDN U19256 ( .A(x[3166]), .B(y[3166]), .Z(n26383) );
  NANDN U19257 ( .A(n37746), .B(n26383), .Z(n55422) );
  NANDN U19258 ( .A(y[3164]), .B(x[3164]), .Z(n9914) );
  NANDN U19259 ( .A(y[3165]), .B(x[3165]), .Z(n37749) );
  AND U19260 ( .A(n9914), .B(n37749), .Z(n55421) );
  XNOR U19261 ( .A(x[3164]), .B(y[3164]), .Z(n26385) );
  NANDN U19262 ( .A(y[3162]), .B(x[3162]), .Z(n9915) );
  NANDN U19263 ( .A(y[3163]), .B(x[3163]), .Z(n26384) );
  AND U19264 ( .A(n9915), .B(n26384), .Z(n55418) );
  XNOR U19265 ( .A(x[3162]), .B(y[3162]), .Z(n26387) );
  ANDN U19266 ( .B(y[3161]), .A(x[3161]), .Z(n26388) );
  ANDN U19267 ( .B(n26387), .A(n26388), .Z(n14816) );
  NANDN U19268 ( .A(x[3159]), .B(y[3159]), .Z(n26390) );
  NANDN U19269 ( .A(x[3160]), .B(y[3160]), .Z(n26389) );
  AND U19270 ( .A(n26390), .B(n26389), .Z(n55414) );
  NANDN U19271 ( .A(y[3158]), .B(x[3158]), .Z(n9916) );
  NANDN U19272 ( .A(y[3159]), .B(x[3159]), .Z(n37733) );
  NAND U19273 ( .A(n9916), .B(n37733), .Z(n55413) );
  NANDN U19274 ( .A(x[3157]), .B(y[3157]), .Z(n51962) );
  NANDN U19275 ( .A(x[3155]), .B(y[3155]), .Z(n26392) );
  NANDN U19276 ( .A(x[3156]), .B(y[3156]), .Z(n26391) );
  AND U19277 ( .A(n26392), .B(n26391), .Z(n55411) );
  NANDN U19278 ( .A(y[3154]), .B(x[3154]), .Z(n37714) );
  NANDN U19279 ( .A(y[3155]), .B(x[3155]), .Z(n37721) );
  NAND U19280 ( .A(n37714), .B(n37721), .Z(n55410) );
  NANDN U19281 ( .A(x[3153]), .B(y[3153]), .Z(n37710) );
  NANDN U19282 ( .A(x[3154]), .B(y[3154]), .Z(n26393) );
  NAND U19283 ( .A(n37710), .B(n26393), .Z(n55409) );
  NANDN U19284 ( .A(y[3152]), .B(x[3152]), .Z(n37709) );
  NANDN U19285 ( .A(y[3153]), .B(x[3153]), .Z(n37715) );
  AND U19286 ( .A(n37709), .B(n37715), .Z(n55408) );
  NANDN U19287 ( .A(x[3151]), .B(y[3151]), .Z(n26394) );
  NANDN U19288 ( .A(x[3152]), .B(y[3152]), .Z(n37711) );
  NAND U19289 ( .A(n26394), .B(n37711), .Z(n55407) );
  NANDN U19290 ( .A(y[3150]), .B(x[3150]), .Z(n37700) );
  ANDN U19291 ( .B(x[3151]), .A(y[3151]), .Z(n37707) );
  ANDN U19292 ( .B(n37700), .A(n37707), .Z(n55406) );
  NANDN U19293 ( .A(x[3149]), .B(y[3149]), .Z(n26396) );
  NANDN U19294 ( .A(x[3150]), .B(y[3150]), .Z(n26395) );
  NAND U19295 ( .A(n26396), .B(n26395), .Z(n55405) );
  NANDN U19296 ( .A(y[3148]), .B(x[3148]), .Z(n9917) );
  NANDN U19297 ( .A(y[3149]), .B(x[3149]), .Z(n37701) );
  NAND U19298 ( .A(n9917), .B(n37701), .Z(n55404) );
  XNOR U19299 ( .A(y[3148]), .B(x[3148]), .Z(n37695) );
  NANDN U19300 ( .A(x[3147]), .B(y[3147]), .Z(n26398) );
  AND U19301 ( .A(n37695), .B(n26398), .Z(n55403) );
  NANDN U19302 ( .A(y[3146]), .B(x[3146]), .Z(n37688) );
  NANDN U19303 ( .A(y[3147]), .B(x[3147]), .Z(n37694) );
  NAND U19304 ( .A(n37688), .B(n37694), .Z(n55402) );
  NANDN U19305 ( .A(x[3145]), .B(y[3145]), .Z(n26400) );
  NANDN U19306 ( .A(x[3146]), .B(y[3146]), .Z(n26399) );
  AND U19307 ( .A(n26400), .B(n26399), .Z(n55401) );
  NANDN U19308 ( .A(y[3144]), .B(x[3144]), .Z(n37682) );
  NANDN U19309 ( .A(y[3145]), .B(x[3145]), .Z(n37689) );
  NAND U19310 ( .A(n37682), .B(n37689), .Z(n55400) );
  NANDN U19311 ( .A(x[3143]), .B(y[3143]), .Z(n26402) );
  NANDN U19312 ( .A(x[3144]), .B(y[3144]), .Z(n26401) );
  NAND U19313 ( .A(n26402), .B(n26401), .Z(n55399) );
  NANDN U19314 ( .A(y[3142]), .B(x[3142]), .Z(n9918) );
  NANDN U19315 ( .A(y[3143]), .B(x[3143]), .Z(n37683) );
  AND U19316 ( .A(n9918), .B(n37683), .Z(n55397) );
  XNOR U19317 ( .A(y[3142]), .B(x[3142]), .Z(n26405) );
  NANDN U19318 ( .A(x[3141]), .B(y[3141]), .Z(n26406) );
  NAND U19319 ( .A(n26405), .B(n26406), .Z(n55396) );
  NANDN U19320 ( .A(y[3140]), .B(x[3140]), .Z(n9919) );
  NANDN U19321 ( .A(y[3141]), .B(x[3141]), .Z(n26404) );
  AND U19322 ( .A(n9919), .B(n26404), .Z(n55395) );
  NANDN U19323 ( .A(y[3138]), .B(x[3138]), .Z(n37668) );
  NANDN U19324 ( .A(y[3139]), .B(x[3139]), .Z(n26407) );
  NAND U19325 ( .A(n37668), .B(n26407), .Z(n55392) );
  NANDN U19326 ( .A(x[3137]), .B(y[3137]), .Z(n26410) );
  NANDN U19327 ( .A(x[3138]), .B(y[3138]), .Z(n26409) );
  AND U19328 ( .A(n26410), .B(n26409), .Z(n55391) );
  NANDN U19329 ( .A(y[3136]), .B(x[3136]), .Z(n9920) );
  NANDN U19330 ( .A(y[3137]), .B(x[3137]), .Z(n37669) );
  NAND U19331 ( .A(n9920), .B(n37669), .Z(n55390) );
  XNOR U19332 ( .A(y[3136]), .B(x[3136]), .Z(n37663) );
  NANDN U19333 ( .A(x[3135]), .B(y[3135]), .Z(n26412) );
  AND U19334 ( .A(n37663), .B(n26412), .Z(n55389) );
  NANDN U19335 ( .A(y[3132]), .B(x[3132]), .Z(n37650) );
  NANDN U19336 ( .A(y[3133]), .B(x[3133]), .Z(n37657) );
  NAND U19337 ( .A(n37650), .B(n37657), .Z(n51965) );
  NANDN U19338 ( .A(y[3130]), .B(x[3130]), .Z(n37644) );
  NANDN U19339 ( .A(y[3131]), .B(x[3131]), .Z(n37651) );
  AND U19340 ( .A(n37644), .B(n37651), .Z(n55386) );
  NANDN U19341 ( .A(x[3129]), .B(y[3129]), .Z(n37641) );
  NANDN U19342 ( .A(x[3130]), .B(y[3130]), .Z(n26417) );
  NAND U19343 ( .A(n37641), .B(n26417), .Z(n55385) );
  NANDN U19344 ( .A(y[3128]), .B(x[3128]), .Z(n26418) );
  NANDN U19345 ( .A(y[3129]), .B(x[3129]), .Z(n37645) );
  NAND U19346 ( .A(n26418), .B(n37645), .Z(n55383) );
  NANDN U19347 ( .A(x[3127]), .B(y[3127]), .Z(n37635) );
  NANDN U19348 ( .A(x[3128]), .B(y[3128]), .Z(n37642) );
  AND U19349 ( .A(n37635), .B(n37642), .Z(n51966) );
  NANDN U19350 ( .A(x[3125]), .B(y[3125]), .Z(n37629) );
  NANDN U19351 ( .A(x[3126]), .B(y[3126]), .Z(n37636) );
  AND U19352 ( .A(n37629), .B(n37636), .Z(n55379) );
  NANDN U19353 ( .A(y[3124]), .B(x[3124]), .Z(n26422) );
  NANDN U19354 ( .A(y[3125]), .B(x[3125]), .Z(n26421) );
  NAND U19355 ( .A(n26422), .B(n26421), .Z(n55378) );
  NANDN U19356 ( .A(x[3123]), .B(y[3123]), .Z(n26424) );
  NANDN U19357 ( .A(x[3124]), .B(y[3124]), .Z(n37630) );
  NAND U19358 ( .A(n26424), .B(n37630), .Z(n55377) );
  NANDN U19359 ( .A(y[3122]), .B(x[3122]), .Z(n26427) );
  NANDN U19360 ( .A(y[3123]), .B(x[3123]), .Z(n26423) );
  AND U19361 ( .A(n26427), .B(n26423), .Z(n55376) );
  NANDN U19362 ( .A(x[3121]), .B(y[3121]), .Z(n26428) );
  NANDN U19363 ( .A(x[3122]), .B(y[3122]), .Z(n26425) );
  NAND U19364 ( .A(n26428), .B(n26425), .Z(n55375) );
  NANDN U19365 ( .A(y[3121]), .B(x[3121]), .Z(n26426) );
  ANDN U19366 ( .B(x[3120]), .A(y[3120]), .Z(n26430) );
  ANDN U19367 ( .B(n26426), .A(n26430), .Z(n55374) );
  NANDN U19368 ( .A(x[3119]), .B(y[3119]), .Z(n9921) );
  NANDN U19369 ( .A(x[3120]), .B(y[3120]), .Z(n26429) );
  NAND U19370 ( .A(n9921), .B(n26429), .Z(n55373) );
  NANDN U19371 ( .A(y[3117]), .B(x[3117]), .Z(n37609) );
  NANDN U19372 ( .A(y[3116]), .B(x[3116]), .Z(n9922) );
  AND U19373 ( .A(n37609), .B(n9922), .Z(n55370) );
  NANDN U19374 ( .A(x[3115]), .B(y[3115]), .Z(n26432) );
  ANDN U19375 ( .B(y[3116]), .A(x[3116]), .Z(n37610) );
  ANDN U19376 ( .B(n26432), .A(n37610), .Z(n55369) );
  NANDN U19377 ( .A(y[3114]), .B(x[3114]), .Z(n26434) );
  NANDN U19378 ( .A(y[3115]), .B(x[3115]), .Z(n37607) );
  NAND U19379 ( .A(n26434), .B(n37607), .Z(n55368) );
  NANDN U19380 ( .A(x[3113]), .B(y[3113]), .Z(n26436) );
  NANDN U19381 ( .A(x[3114]), .B(y[3114]), .Z(n26433) );
  AND U19382 ( .A(n26436), .B(n26433), .Z(n55367) );
  NANDN U19383 ( .A(y[3112]), .B(x[3112]), .Z(n26438) );
  NANDN U19384 ( .A(y[3113]), .B(x[3113]), .Z(n26435) );
  NAND U19385 ( .A(n26438), .B(n26435), .Z(n55366) );
  NANDN U19386 ( .A(x[3111]), .B(y[3111]), .Z(n37595) );
  NANDN U19387 ( .A(x[3112]), .B(y[3112]), .Z(n26437) );
  NAND U19388 ( .A(n37595), .B(n26437), .Z(n55365) );
  NANDN U19389 ( .A(y[3110]), .B(x[3110]), .Z(n26440) );
  NANDN U19390 ( .A(y[3111]), .B(x[3111]), .Z(n26439) );
  AND U19391 ( .A(n26440), .B(n26439), .Z(n55364) );
  ANDN U19392 ( .B(y[3110]), .A(x[3110]), .Z(n37597) );
  NANDN U19393 ( .A(x[3109]), .B(y[3109]), .Z(n37589) );
  NANDN U19394 ( .A(n37597), .B(n37589), .Z(n55363) );
  NANDN U19395 ( .A(y[3108]), .B(x[3108]), .Z(n26442) );
  NANDN U19396 ( .A(y[3109]), .B(x[3109]), .Z(n26441) );
  AND U19397 ( .A(n26442), .B(n26441), .Z(n55362) );
  NANDN U19398 ( .A(x[3107]), .B(y[3107]), .Z(n37583) );
  NANDN U19399 ( .A(x[3108]), .B(y[3108]), .Z(n37590) );
  NAND U19400 ( .A(n37583), .B(n37590), .Z(n55360) );
  NANDN U19401 ( .A(y[3106]), .B(x[3106]), .Z(n26444) );
  NANDN U19402 ( .A(y[3107]), .B(x[3107]), .Z(n26443) );
  NAND U19403 ( .A(n26444), .B(n26443), .Z(n55358) );
  NANDN U19404 ( .A(x[3105]), .B(y[3105]), .Z(n26446) );
  NANDN U19405 ( .A(x[3106]), .B(y[3106]), .Z(n37584) );
  AND U19406 ( .A(n26446), .B(n37584), .Z(n55356) );
  NANDN U19407 ( .A(y[3104]), .B(x[3104]), .Z(n26448) );
  NANDN U19408 ( .A(y[3105]), .B(x[3105]), .Z(n26445) );
  NAND U19409 ( .A(n26448), .B(n26445), .Z(n55354) );
  NANDN U19410 ( .A(x[3103]), .B(y[3103]), .Z(n37573) );
  NANDN U19411 ( .A(x[3104]), .B(y[3104]), .Z(n26447) );
  AND U19412 ( .A(n37573), .B(n26447), .Z(n55352) );
  NANDN U19413 ( .A(y[3102]), .B(x[3102]), .Z(n9923) );
  NANDN U19414 ( .A(y[3103]), .B(x[3103]), .Z(n26449) );
  NAND U19415 ( .A(n9923), .B(n26449), .Z(n55350) );
  XNOR U19416 ( .A(y[3102]), .B(x[3102]), .Z(n37570) );
  NANDN U19417 ( .A(x[3101]), .B(y[3101]), .Z(n26450) );
  NAND U19418 ( .A(n37570), .B(n26450), .Z(n55348) );
  NANDN U19419 ( .A(y[3100]), .B(x[3100]), .Z(n26453) );
  ANDN U19420 ( .B(x[3101]), .A(y[3101]), .Z(n37569) );
  ANDN U19421 ( .B(n26453), .A(n37569), .Z(n55346) );
  NANDN U19422 ( .A(x[3099]), .B(y[3099]), .Z(n26454) );
  NANDN U19423 ( .A(x[3100]), .B(y[3100]), .Z(n26451) );
  NAND U19424 ( .A(n26454), .B(n26451), .Z(n55344) );
  NANDN U19425 ( .A(y[3098]), .B(x[3098]), .Z(n26456) );
  NANDN U19426 ( .A(y[3099]), .B(x[3099]), .Z(n26452) );
  AND U19427 ( .A(n26456), .B(n26452), .Z(n55342) );
  NANDN U19428 ( .A(x[3097]), .B(y[3097]), .Z(n37556) );
  NANDN U19429 ( .A(x[3098]), .B(y[3098]), .Z(n26455) );
  NAND U19430 ( .A(n37556), .B(n26455), .Z(n55340) );
  NANDN U19431 ( .A(y[3096]), .B(x[3096]), .Z(n37553) );
  NANDN U19432 ( .A(y[3097]), .B(x[3097]), .Z(n26457) );
  NAND U19433 ( .A(n37553), .B(n26457), .Z(n55338) );
  NANDN U19434 ( .A(x[3095]), .B(y[3095]), .Z(n26458) );
  NANDN U19435 ( .A(x[3096]), .B(y[3096]), .Z(n37557) );
  AND U19436 ( .A(n26458), .B(n37557), .Z(n55336) );
  NANDN U19437 ( .A(y[3094]), .B(x[3094]), .Z(n37547) );
  NANDN U19438 ( .A(y[3095]), .B(x[3095]), .Z(n37554) );
  NAND U19439 ( .A(n37547), .B(n37554), .Z(n55334) );
  NANDN U19440 ( .A(x[3093]), .B(y[3093]), .Z(n26460) );
  NANDN U19441 ( .A(x[3094]), .B(y[3094]), .Z(n26459) );
  AND U19442 ( .A(n26460), .B(n26459), .Z(n55332) );
  NANDN U19443 ( .A(y[3092]), .B(x[3092]), .Z(n37541) );
  NANDN U19444 ( .A(y[3093]), .B(x[3093]), .Z(n37548) );
  NAND U19445 ( .A(n37541), .B(n37548), .Z(n55330) );
  NANDN U19446 ( .A(x[3091]), .B(y[3091]), .Z(n26462) );
  NANDN U19447 ( .A(x[3092]), .B(y[3092]), .Z(n26461) );
  NAND U19448 ( .A(n26462), .B(n26461), .Z(n55328) );
  NANDN U19449 ( .A(y[3090]), .B(x[3090]), .Z(n37535) );
  NANDN U19450 ( .A(y[3091]), .B(x[3091]), .Z(n37542) );
  AND U19451 ( .A(n37535), .B(n37542), .Z(n55326) );
  NANDN U19452 ( .A(x[3089]), .B(y[3089]), .Z(n26464) );
  NANDN U19453 ( .A(x[3090]), .B(y[3090]), .Z(n26463) );
  NAND U19454 ( .A(n26464), .B(n26463), .Z(n55324) );
  NANDN U19455 ( .A(y[3088]), .B(x[3088]), .Z(n9924) );
  NANDN U19456 ( .A(y[3089]), .B(x[3089]), .Z(n37536) );
  AND U19457 ( .A(n9924), .B(n37536), .Z(n55322) );
  XNOR U19458 ( .A(x[3088]), .B(y[3088]), .Z(n37529) );
  NANDN U19459 ( .A(y[3086]), .B(x[3086]), .Z(n37522) );
  NANDN U19460 ( .A(y[3087]), .B(x[3087]), .Z(n37528) );
  AND U19461 ( .A(n37522), .B(n37528), .Z(n55318) );
  NANDN U19462 ( .A(x[3085]), .B(y[3085]), .Z(n26466) );
  NANDN U19463 ( .A(x[3086]), .B(y[3086]), .Z(n26465) );
  NAND U19464 ( .A(n26466), .B(n26465), .Z(n55317) );
  NANDN U19465 ( .A(y[3084]), .B(x[3084]), .Z(n37516) );
  NANDN U19466 ( .A(y[3085]), .B(x[3085]), .Z(n37523) );
  AND U19467 ( .A(n37516), .B(n37523), .Z(n55316) );
  NANDN U19468 ( .A(x[3083]), .B(y[3083]), .Z(n26468) );
  NANDN U19469 ( .A(x[3084]), .B(y[3084]), .Z(n26467) );
  NAND U19470 ( .A(n26468), .B(n26467), .Z(n55315) );
  NANDN U19471 ( .A(y[3082]), .B(x[3082]), .Z(n37510) );
  NANDN U19472 ( .A(y[3083]), .B(x[3083]), .Z(n37517) );
  AND U19473 ( .A(n37510), .B(n37517), .Z(n55314) );
  NANDN U19474 ( .A(x[3081]), .B(y[3081]), .Z(n26470) );
  NANDN U19475 ( .A(x[3082]), .B(y[3082]), .Z(n26469) );
  NAND U19476 ( .A(n26470), .B(n26469), .Z(n55313) );
  NANDN U19477 ( .A(y[3080]), .B(x[3080]), .Z(n9925) );
  NANDN U19478 ( .A(y[3081]), .B(x[3081]), .Z(n37511) );
  AND U19479 ( .A(n9925), .B(n37511), .Z(n55312) );
  XNOR U19480 ( .A(x[3080]), .B(y[3080]), .Z(n26472) );
  NANDN U19481 ( .A(y[3078]), .B(x[3078]), .Z(n26473) );
  NANDN U19482 ( .A(y[3079]), .B(x[3079]), .Z(n26471) );
  AND U19483 ( .A(n26473), .B(n26471), .Z(n55310) );
  ANDN U19484 ( .B(y[3077]), .A(x[3077]), .Z(n37499) );
  ANDN U19485 ( .B(y[3078]), .A(x[3078]), .Z(n37504) );
  OR U19486 ( .A(n37499), .B(n37504), .Z(n55309) );
  NANDN U19487 ( .A(y[3076]), .B(x[3076]), .Z(n9926) );
  NANDN U19488 ( .A(y[3077]), .B(x[3077]), .Z(n26474) );
  AND U19489 ( .A(n9926), .B(n26474), .Z(n51968) );
  NANDN U19490 ( .A(x[3075]), .B(y[3075]), .Z(n55306) );
  XNOR U19491 ( .A(x[3076]), .B(y[3076]), .Z(n37496) );
  NANDN U19492 ( .A(y[3074]), .B(x[3074]), .Z(n37489) );
  NANDN U19493 ( .A(y[3075]), .B(x[3075]), .Z(n37495) );
  NAND U19494 ( .A(n37489), .B(n37495), .Z(n51969) );
  NANDN U19495 ( .A(x[3073]), .B(y[3073]), .Z(n26476) );
  NANDN U19496 ( .A(x[3074]), .B(y[3074]), .Z(n26475) );
  AND U19497 ( .A(n26476), .B(n26475), .Z(n55305) );
  NANDN U19498 ( .A(x[3069]), .B(y[3069]), .Z(n26480) );
  NANDN U19499 ( .A(x[3070]), .B(y[3070]), .Z(n26479) );
  AND U19500 ( .A(n26480), .B(n26479), .Z(n55302) );
  NANDN U19501 ( .A(y[3068]), .B(x[3068]), .Z(n26482) );
  NANDN U19502 ( .A(y[3069]), .B(x[3069]), .Z(n37478) );
  NAND U19503 ( .A(n26482), .B(n37478), .Z(n55301) );
  NANDN U19504 ( .A(x[3067]), .B(y[3067]), .Z(n26485) );
  XNOR U19505 ( .A(x[3068]), .B(y[3068]), .Z(n9927) );
  NAND U19506 ( .A(n26485), .B(n9927), .Z(n55300) );
  NANDN U19507 ( .A(y[3066]), .B(x[3066]), .Z(n26486) );
  NANDN U19508 ( .A(y[3067]), .B(x[3067]), .Z(n26483) );
  AND U19509 ( .A(n26486), .B(n26483), .Z(n51971) );
  NANDN U19510 ( .A(y[3064]), .B(x[3064]), .Z(n37462) );
  NANDN U19511 ( .A(y[3065]), .B(x[3065]), .Z(n26487) );
  AND U19512 ( .A(n37462), .B(n26487), .Z(n55298) );
  NANDN U19513 ( .A(x[3063]), .B(y[3063]), .Z(n26490) );
  XNOR U19514 ( .A(x[3064]), .B(y[3064]), .Z(n9928) );
  NAND U19515 ( .A(n26490), .B(n9928), .Z(n55296) );
  NANDN U19516 ( .A(y[3062]), .B(x[3062]), .Z(n9929) );
  NANDN U19517 ( .A(y[3063]), .B(x[3063]), .Z(n37463) );
  NAND U19518 ( .A(n9929), .B(n37463), .Z(n51972) );
  XNOR U19519 ( .A(y[3062]), .B(x[3062]), .Z(n37457) );
  NANDN U19520 ( .A(x[3061]), .B(y[3061]), .Z(n26492) );
  AND U19521 ( .A(n37457), .B(n26492), .Z(n55295) );
  NANDN U19522 ( .A(y[3058]), .B(x[3058]), .Z(n37444) );
  NANDN U19523 ( .A(y[3059]), .B(x[3059]), .Z(n37450) );
  NAND U19524 ( .A(n37444), .B(n37450), .Z(n55293) );
  NANDN U19525 ( .A(x[3057]), .B(y[3057]), .Z(n26496) );
  NANDN U19526 ( .A(x[3058]), .B(y[3058]), .Z(n26495) );
  NAND U19527 ( .A(n26496), .B(n26495), .Z(n51974) );
  NANDN U19528 ( .A(y[3056]), .B(x[3056]), .Z(n37438) );
  NANDN U19529 ( .A(y[3057]), .B(x[3057]), .Z(n37445) );
  AND U19530 ( .A(n37438), .B(n37445), .Z(n55292) );
  ANDN U19531 ( .B(y[3053]), .A(x[3053]), .Z(n37431) );
  NANDN U19532 ( .A(x[3054]), .B(y[3054]), .Z(n26499) );
  NANDN U19533 ( .A(n37431), .B(n26499), .Z(n55290) );
  NANDN U19534 ( .A(y[3052]), .B(x[3052]), .Z(n26502) );
  NANDN U19535 ( .A(y[3053]), .B(x[3053]), .Z(n26501) );
  NAND U19536 ( .A(n26502), .B(n26501), .Z(n51976) );
  NANDN U19537 ( .A(x[3051]), .B(y[3051]), .Z(n37425) );
  ANDN U19538 ( .B(y[3052]), .A(x[3052]), .Z(n37432) );
  ANDN U19539 ( .B(n37425), .A(n37432), .Z(n55287) );
  NANDN U19540 ( .A(x[3049]), .B(y[3049]), .Z(n55284) );
  XNOR U19541 ( .A(x[3050]), .B(y[3050]), .Z(n26505) );
  AND U19542 ( .A(n55284), .B(n26505), .Z(n14692) );
  NANDN U19543 ( .A(y[3048]), .B(x[3048]), .Z(n26507) );
  NANDN U19544 ( .A(y[3049]), .B(x[3049]), .Z(n26504) );
  NAND U19545 ( .A(n26507), .B(n26504), .Z(n55283) );
  NANDN U19546 ( .A(x[3047]), .B(y[3047]), .Z(n37417) );
  NANDN U19547 ( .A(x[3048]), .B(y[3048]), .Z(n26506) );
  AND U19548 ( .A(n37417), .B(n26506), .Z(n55282) );
  NANDN U19549 ( .A(y[3046]), .B(x[3046]), .Z(n9930) );
  NANDN U19550 ( .A(y[3047]), .B(x[3047]), .Z(n26508) );
  NAND U19551 ( .A(n9930), .B(n26508), .Z(n55281) );
  NANDN U19552 ( .A(x[3045]), .B(y[3045]), .Z(n55279) );
  NANDN U19553 ( .A(x[3041]), .B(y[3041]), .Z(n26510) );
  ANDN U19554 ( .B(y[3042]), .A(x[3042]), .Z(n37405) );
  ANDN U19555 ( .B(n26510), .A(n37405), .Z(n55274) );
  NANDN U19556 ( .A(y[3040]), .B(x[3040]), .Z(n26511) );
  NANDN U19557 ( .A(y[3041]), .B(x[3041]), .Z(n55272) );
  AND U19558 ( .A(n26511), .B(n55272), .Z(n55271) );
  NANDN U19559 ( .A(y[3038]), .B(x[3038]), .Z(n37391) );
  NANDN U19560 ( .A(y[3039]), .B(x[3039]), .Z(n26512) );
  AND U19561 ( .A(n37391), .B(n26512), .Z(n55267) );
  NANDN U19562 ( .A(x[3037]), .B(y[3037]), .Z(n26513) );
  NANDN U19563 ( .A(x[3038]), .B(y[3038]), .Z(n37396) );
  NAND U19564 ( .A(n26513), .B(n37396), .Z(n55265) );
  NANDN U19565 ( .A(y[3036]), .B(x[3036]), .Z(n37385) );
  NANDN U19566 ( .A(y[3037]), .B(x[3037]), .Z(n37392) );
  NAND U19567 ( .A(n37385), .B(n37392), .Z(n55263) );
  NANDN U19568 ( .A(x[3035]), .B(y[3035]), .Z(n26515) );
  NANDN U19569 ( .A(x[3036]), .B(y[3036]), .Z(n26514) );
  AND U19570 ( .A(n26515), .B(n26514), .Z(n55261) );
  NANDN U19571 ( .A(y[3034]), .B(x[3034]), .Z(n37379) );
  NANDN U19572 ( .A(y[3035]), .B(x[3035]), .Z(n37386) );
  NAND U19573 ( .A(n37379), .B(n37386), .Z(n55259) );
  NANDN U19574 ( .A(x[3033]), .B(y[3033]), .Z(n26517) );
  NANDN U19575 ( .A(x[3034]), .B(y[3034]), .Z(n26516) );
  AND U19576 ( .A(n26517), .B(n26516), .Z(n55257) );
  NANDN U19577 ( .A(y[3032]), .B(x[3032]), .Z(n37373) );
  NANDN U19578 ( .A(y[3033]), .B(x[3033]), .Z(n37380) );
  NAND U19579 ( .A(n37373), .B(n37380), .Z(n55255) );
  NANDN U19580 ( .A(x[3031]), .B(y[3031]), .Z(n37369) );
  NANDN U19581 ( .A(x[3032]), .B(y[3032]), .Z(n26518) );
  NAND U19582 ( .A(n37369), .B(n26518), .Z(n55253) );
  NANDN U19583 ( .A(y[3030]), .B(x[3030]), .Z(n37368) );
  NANDN U19584 ( .A(y[3031]), .B(x[3031]), .Z(n37374) );
  AND U19585 ( .A(n37368), .B(n37374), .Z(n55251) );
  NANDN U19586 ( .A(x[3029]), .B(y[3029]), .Z(n26519) );
  XNOR U19587 ( .A(x[3030]), .B(y[3030]), .Z(n9931) );
  NAND U19588 ( .A(n26519), .B(n9931), .Z(n55249) );
  NANDN U19589 ( .A(y[3028]), .B(x[3028]), .Z(n9932) );
  ANDN U19590 ( .B(x[3029]), .A(y[3029]), .Z(n37366) );
  ANDN U19591 ( .B(n9932), .A(n37366), .Z(n55247) );
  XNOR U19592 ( .A(y[3028]), .B(x[3028]), .Z(n37360) );
  NANDN U19593 ( .A(x[3027]), .B(y[3027]), .Z(n26521) );
  NAND U19594 ( .A(n37360), .B(n26521), .Z(n55245) );
  NANDN U19595 ( .A(y[3026]), .B(x[3026]), .Z(n37353) );
  NANDN U19596 ( .A(y[3027]), .B(x[3027]), .Z(n37359) );
  NAND U19597 ( .A(n37353), .B(n37359), .Z(n55243) );
  NANDN U19598 ( .A(x[3025]), .B(y[3025]), .Z(n26523) );
  NANDN U19599 ( .A(x[3026]), .B(y[3026]), .Z(n26522) );
  AND U19600 ( .A(n26523), .B(n26522), .Z(n55241) );
  NANDN U19601 ( .A(y[3024]), .B(x[3024]), .Z(n37347) );
  NANDN U19602 ( .A(y[3025]), .B(x[3025]), .Z(n37354) );
  NAND U19603 ( .A(n37347), .B(n37354), .Z(n55239) );
  NANDN U19604 ( .A(x[3023]), .B(y[3023]), .Z(n37344) );
  NANDN U19605 ( .A(x[3024]), .B(y[3024]), .Z(n26524) );
  AND U19606 ( .A(n37344), .B(n26524), .Z(n55237) );
  NANDN U19607 ( .A(y[3022]), .B(x[3022]), .Z(n26525) );
  NANDN U19608 ( .A(y[3023]), .B(x[3023]), .Z(n37348) );
  NAND U19609 ( .A(n26525), .B(n37348), .Z(n55235) );
  NANDN U19610 ( .A(x[3021]), .B(y[3021]), .Z(n37338) );
  NANDN U19611 ( .A(x[3022]), .B(y[3022]), .Z(n37345) );
  NAND U19612 ( .A(n37338), .B(n37345), .Z(n55233) );
  NANDN U19613 ( .A(y[3020]), .B(x[3020]), .Z(n26527) );
  NANDN U19614 ( .A(y[3021]), .B(x[3021]), .Z(n26526) );
  AND U19615 ( .A(n26527), .B(n26526), .Z(n55231) );
  NANDN U19616 ( .A(x[3019]), .B(y[3019]), .Z(n37332) );
  NANDN U19617 ( .A(x[3020]), .B(y[3020]), .Z(n37339) );
  NAND U19618 ( .A(n37332), .B(n37339), .Z(n55229) );
  NANDN U19619 ( .A(y[3019]), .B(x[3019]), .Z(n26528) );
  ANDN U19620 ( .B(x[3018]), .A(y[3018]), .Z(n37327) );
  ANDN U19621 ( .B(n26528), .A(n37327), .Z(n55227) );
  ANDN U19622 ( .B(y[3017]), .A(x[3017]), .Z(n37323) );
  NANDN U19623 ( .A(x[3018]), .B(y[3018]), .Z(n37333) );
  NANDN U19624 ( .A(n37323), .B(n37333), .Z(n55226) );
  ANDN U19625 ( .B(x[3017]), .A(y[3017]), .Z(n37328) );
  NANDN U19626 ( .A(y[3016]), .B(x[3016]), .Z(n37320) );
  NANDN U19627 ( .A(n37328), .B(n37320), .Z(n55225) );
  NANDN U19628 ( .A(x[3015]), .B(y[3015]), .Z(n26529) );
  ANDN U19629 ( .B(y[3016]), .A(x[3016]), .Z(n37326) );
  ANDN U19630 ( .B(n26529), .A(n37326), .Z(n55224) );
  NANDN U19631 ( .A(y[3014]), .B(x[3014]), .Z(n9933) );
  NANDN U19632 ( .A(y[3015]), .B(x[3015]), .Z(n37321) );
  NAND U19633 ( .A(n9933), .B(n37321), .Z(n55223) );
  XNOR U19634 ( .A(x[3014]), .B(y[3014]), .Z(n37314) );
  ANDN U19635 ( .B(y[3013]), .A(x[3013]), .Z(n51977) );
  ANDN U19636 ( .B(n37314), .A(n51977), .Z(n14650) );
  NANDN U19637 ( .A(y[3012]), .B(x[3012]), .Z(n37307) );
  NANDN U19638 ( .A(y[3013]), .B(x[3013]), .Z(n37315) );
  AND U19639 ( .A(n37307), .B(n37315), .Z(n55222) );
  ANDN U19640 ( .B(y[3012]), .A(x[3012]), .Z(n37311) );
  NANDN U19641 ( .A(x[3011]), .B(y[3011]), .Z(n26530) );
  NANDN U19642 ( .A(n37311), .B(n26530), .Z(n55221) );
  NANDN U19643 ( .A(y[3010]), .B(x[3010]), .Z(n37300) );
  NANDN U19644 ( .A(y[3011]), .B(x[3011]), .Z(n37309) );
  AND U19645 ( .A(n37300), .B(n37309), .Z(n55220) );
  NANDN U19646 ( .A(x[3009]), .B(y[3009]), .Z(n26532) );
  NANDN U19647 ( .A(x[3010]), .B(y[3010]), .Z(n26531) );
  NAND U19648 ( .A(n26532), .B(n26531), .Z(n55219) );
  NANDN U19649 ( .A(y[3008]), .B(x[3008]), .Z(n9934) );
  NANDN U19650 ( .A(y[3009]), .B(x[3009]), .Z(n37301) );
  AND U19651 ( .A(n9934), .B(n37301), .Z(n55218) );
  XNOR U19652 ( .A(x[3008]), .B(y[3008]), .Z(n37295) );
  NANDN U19653 ( .A(y[3004]), .B(x[3004]), .Z(n37282) );
  NANDN U19654 ( .A(y[3005]), .B(x[3005]), .Z(n37289) );
  NAND U19655 ( .A(n37282), .B(n37289), .Z(n55212) );
  NANDN U19656 ( .A(x[3003]), .B(y[3003]), .Z(n26536) );
  NANDN U19657 ( .A(x[3004]), .B(y[3004]), .Z(n26535) );
  NAND U19658 ( .A(n26536), .B(n26535), .Z(n55211) );
  NANDN U19659 ( .A(y[3002]), .B(x[3002]), .Z(n37276) );
  NANDN U19660 ( .A(y[3003]), .B(x[3003]), .Z(n37283) );
  AND U19661 ( .A(n37276), .B(n37283), .Z(n55209) );
  NANDN U19662 ( .A(x[3001]), .B(y[3001]), .Z(n26538) );
  NANDN U19663 ( .A(x[3002]), .B(y[3002]), .Z(n26537) );
  NAND U19664 ( .A(n26538), .B(n26537), .Z(n55208) );
  NANDN U19665 ( .A(y[3000]), .B(x[3000]), .Z(n37270) );
  NANDN U19666 ( .A(y[3001]), .B(x[3001]), .Z(n37277) );
  AND U19667 ( .A(n37270), .B(n37277), .Z(n55207) );
  NANDN U19668 ( .A(x[2999]), .B(y[2999]), .Z(n26540) );
  NANDN U19669 ( .A(x[3000]), .B(y[3000]), .Z(n26539) );
  NAND U19670 ( .A(n26540), .B(n26539), .Z(n55206) );
  NANDN U19671 ( .A(y[2998]), .B(x[2998]), .Z(n37264) );
  NANDN U19672 ( .A(y[2999]), .B(x[2999]), .Z(n37271) );
  NAND U19673 ( .A(n37264), .B(n37271), .Z(n55205) );
  NANDN U19674 ( .A(x[2997]), .B(y[2997]), .Z(n26542) );
  NANDN U19675 ( .A(x[2998]), .B(y[2998]), .Z(n26541) );
  AND U19676 ( .A(n26542), .B(n26541), .Z(n55204) );
  NANDN U19677 ( .A(y[2996]), .B(x[2996]), .Z(n37258) );
  NANDN U19678 ( .A(y[2997]), .B(x[2997]), .Z(n37265) );
  NAND U19679 ( .A(n37258), .B(n37265), .Z(n55203) );
  NANDN U19680 ( .A(x[2995]), .B(y[2995]), .Z(n26544) );
  XNOR U19681 ( .A(y[2996]), .B(x[2996]), .Z(n9935) );
  AND U19682 ( .A(n26544), .B(n9935), .Z(n55202) );
  NANDN U19683 ( .A(y[2992]), .B(x[2992]), .Z(n37246) );
  NANDN U19684 ( .A(y[2993]), .B(x[2993]), .Z(n37252) );
  NAND U19685 ( .A(n37246), .B(n37252), .Z(n51980) );
  NANDN U19686 ( .A(y[2990]), .B(x[2990]), .Z(n37240) );
  NANDN U19687 ( .A(y[2991]), .B(x[2991]), .Z(n37247) );
  AND U19688 ( .A(n37240), .B(n37247), .Z(n55199) );
  NANDN U19689 ( .A(x[2989]), .B(y[2989]), .Z(n37236) );
  NANDN U19690 ( .A(x[2990]), .B(y[2990]), .Z(n26549) );
  NAND U19691 ( .A(n37236), .B(n26549), .Z(n55198) );
  NANDN U19692 ( .A(y[2988]), .B(x[2988]), .Z(n26550) );
  NANDN U19693 ( .A(y[2989]), .B(x[2989]), .Z(n37241) );
  NAND U19694 ( .A(n26550), .B(n37241), .Z(n55197) );
  NANDN U19695 ( .A(x[2988]), .B(y[2988]), .Z(n37237) );
  ANDN U19696 ( .B(y[2987]), .A(x[2987]), .Z(n37231) );
  ANDN U19697 ( .B(n37237), .A(n37231), .Z(n55196) );
  NANDN U19698 ( .A(y[2986]), .B(x[2986]), .Z(n26552) );
  NANDN U19699 ( .A(y[2987]), .B(x[2987]), .Z(n26551) );
  NAND U19700 ( .A(n26552), .B(n26551), .Z(n55195) );
  NANDN U19701 ( .A(x[2985]), .B(y[2985]), .Z(n26554) );
  ANDN U19702 ( .B(y[2986]), .A(x[2986]), .Z(n37232) );
  ANDN U19703 ( .B(n26554), .A(n37232), .Z(n55193) );
  NANDN U19704 ( .A(y[2984]), .B(x[2984]), .Z(n26556) );
  NANDN U19705 ( .A(y[2985]), .B(x[2985]), .Z(n26553) );
  NAND U19706 ( .A(n26556), .B(n26553), .Z(n55192) );
  NANDN U19707 ( .A(x[2983]), .B(y[2983]), .Z(n26559) );
  NANDN U19708 ( .A(x[2984]), .B(y[2984]), .Z(n26555) );
  NAND U19709 ( .A(n26559), .B(n26555), .Z(n55191) );
  NANDN U19710 ( .A(y[2982]), .B(x[2982]), .Z(n26560) );
  NANDN U19711 ( .A(y[2983]), .B(x[2983]), .Z(n26557) );
  AND U19712 ( .A(n26560), .B(n26557), .Z(n51981) );
  NANDN U19713 ( .A(y[2980]), .B(x[2980]), .Z(n26564) );
  NANDN U19714 ( .A(y[2981]), .B(x[2981]), .Z(n26561) );
  AND U19715 ( .A(n26564), .B(n26561), .Z(n55189) );
  NANDN U19716 ( .A(x[2979]), .B(y[2979]), .Z(n26566) );
  XNOR U19717 ( .A(x[2980]), .B(y[2980]), .Z(n9936) );
  NAND U19718 ( .A(n26566), .B(n9936), .Z(n55188) );
  NANDN U19719 ( .A(y[2978]), .B(x[2978]), .Z(n9937) );
  NANDN U19720 ( .A(y[2979]), .B(x[2979]), .Z(n26565) );
  NAND U19721 ( .A(n9937), .B(n26565), .Z(n55187) );
  XNOR U19722 ( .A(y[2978]), .B(x[2978]), .Z(n26569) );
  NANDN U19723 ( .A(x[2977]), .B(y[2977]), .Z(n26570) );
  AND U19724 ( .A(n26569), .B(n26570), .Z(n55186) );
  NANDN U19725 ( .A(y[2976]), .B(x[2976]), .Z(n37206) );
  NANDN U19726 ( .A(y[2977]), .B(x[2977]), .Z(n26568) );
  NAND U19727 ( .A(n37206), .B(n26568), .Z(n55185) );
  NANDN U19728 ( .A(x[2975]), .B(y[2975]), .Z(n26572) );
  NANDN U19729 ( .A(x[2976]), .B(y[2976]), .Z(n26571) );
  AND U19730 ( .A(n26572), .B(n26571), .Z(n55184) );
  NANDN U19731 ( .A(y[2974]), .B(x[2974]), .Z(n37200) );
  NANDN U19732 ( .A(y[2975]), .B(x[2975]), .Z(n37207) );
  NAND U19733 ( .A(n37200), .B(n37207), .Z(n55183) );
  NANDN U19734 ( .A(x[2973]), .B(y[2973]), .Z(n26574) );
  NANDN U19735 ( .A(x[2974]), .B(y[2974]), .Z(n26573) );
  NAND U19736 ( .A(n26574), .B(n26573), .Z(n55182) );
  NANDN U19737 ( .A(y[2972]), .B(x[2972]), .Z(n37194) );
  NANDN U19738 ( .A(y[2973]), .B(x[2973]), .Z(n37201) );
  AND U19739 ( .A(n37194), .B(n37201), .Z(n55181) );
  NANDN U19740 ( .A(x[2971]), .B(y[2971]), .Z(n26576) );
  NANDN U19741 ( .A(x[2972]), .B(y[2972]), .Z(n26575) );
  NAND U19742 ( .A(n26576), .B(n26575), .Z(n55180) );
  NANDN U19743 ( .A(y[2970]), .B(x[2970]), .Z(n9938) );
  NANDN U19744 ( .A(y[2971]), .B(x[2971]), .Z(n37195) );
  AND U19745 ( .A(n9938), .B(n37195), .Z(n55179) );
  NANDN U19746 ( .A(x[2967]), .B(y[2967]), .Z(n26579) );
  NANDN U19747 ( .A(x[2968]), .B(y[2968]), .Z(n26578) );
  NAND U19748 ( .A(n26579), .B(n26578), .Z(n51983) );
  NANDN U19749 ( .A(y[2966]), .B(x[2966]), .Z(n37176) );
  NANDN U19750 ( .A(y[2967]), .B(x[2967]), .Z(n37183) );
  AND U19751 ( .A(n37176), .B(n37183), .Z(n55174) );
  NANDN U19752 ( .A(y[2962]), .B(x[2962]), .Z(n26582) );
  NANDN U19753 ( .A(y[2963]), .B(x[2963]), .Z(n37170) );
  NAND U19754 ( .A(n26582), .B(n37170), .Z(n51985) );
  NANDN U19755 ( .A(x[2961]), .B(y[2961]), .Z(n37162) );
  NANDN U19756 ( .A(x[2962]), .B(y[2962]), .Z(n37168) );
  AND U19757 ( .A(n37162), .B(n37168), .Z(n51986) );
  NANDN U19758 ( .A(y[2958]), .B(x[2958]), .Z(n26586) );
  NANDN U19759 ( .A(y[2959]), .B(x[2959]), .Z(n26585) );
  NAND U19760 ( .A(n26586), .B(n26585), .Z(n55166) );
  NANDN U19761 ( .A(x[2957]), .B(y[2957]), .Z(n26588) );
  NANDN U19762 ( .A(x[2958]), .B(y[2958]), .Z(n37157) );
  NAND U19763 ( .A(n26588), .B(n37157), .Z(n55165) );
  NANDN U19764 ( .A(y[2956]), .B(x[2956]), .Z(n26591) );
  NANDN U19765 ( .A(y[2957]), .B(x[2957]), .Z(n26587) );
  AND U19766 ( .A(n26591), .B(n26587), .Z(n55164) );
  NANDN U19767 ( .A(x[2955]), .B(y[2955]), .Z(n26592) );
  NANDN U19768 ( .A(x[2956]), .B(y[2956]), .Z(n26589) );
  NAND U19769 ( .A(n26592), .B(n26589), .Z(n55163) );
  NANDN U19770 ( .A(y[2954]), .B(x[2954]), .Z(n26593) );
  NANDN U19771 ( .A(y[2955]), .B(x[2955]), .Z(n26590) );
  AND U19772 ( .A(n26593), .B(n26590), .Z(n55162) );
  NANDN U19773 ( .A(y[2953]), .B(x[2953]), .Z(n26594) );
  NANDN U19774 ( .A(y[2952]), .B(x[2952]), .Z(n26596) );
  NANDN U19775 ( .A(x[2953]), .B(y[2953]), .Z(n9939) );
  NANDN U19776 ( .A(x[2952]), .B(y[2952]), .Z(n9940) );
  AND U19777 ( .A(n9940), .B(n9939), .Z(n37144) );
  NANDN U19778 ( .A(x[2951]), .B(y[2951]), .Z(n26597) );
  NAND U19779 ( .A(n37144), .B(n26597), .Z(n55159) );
  NANDN U19780 ( .A(x[2949]), .B(y[2949]), .Z(n26599) );
  NANDN U19781 ( .A(x[2950]), .B(y[2950]), .Z(n26598) );
  AND U19782 ( .A(n26599), .B(n26598), .Z(n55157) );
  NANDN U19783 ( .A(y[2946]), .B(x[2946]), .Z(n37124) );
  NANDN U19784 ( .A(y[2947]), .B(x[2947]), .Z(n37131) );
  NAND U19785 ( .A(n37124), .B(n37131), .Z(n51989) );
  NANDN U19786 ( .A(y[2944]), .B(x[2944]), .Z(n26605) );
  NANDN U19787 ( .A(y[2945]), .B(x[2945]), .Z(n37125) );
  AND U19788 ( .A(n26605), .B(n37125), .Z(n55154) );
  NANDN U19789 ( .A(x[2943]), .B(y[2943]), .Z(n26607) );
  NANDN U19790 ( .A(x[2944]), .B(y[2944]), .Z(n26604) );
  NAND U19791 ( .A(n26607), .B(n26604), .Z(n55153) );
  NANDN U19792 ( .A(y[2942]), .B(x[2942]), .Z(n37116) );
  NANDN U19793 ( .A(y[2943]), .B(x[2943]), .Z(n26606) );
  NAND U19794 ( .A(n37116), .B(n26606), .Z(n55152) );
  NANDN U19795 ( .A(x[2941]), .B(y[2941]), .Z(n26609) );
  NANDN U19796 ( .A(x[2942]), .B(y[2942]), .Z(n26608) );
  AND U19797 ( .A(n26609), .B(n26608), .Z(n55151) );
  ANDN U19798 ( .B(x[2941]), .A(y[2941]), .Z(n37114) );
  NANDN U19799 ( .A(y[2940]), .B(x[2940]), .Z(n37107) );
  NANDN U19800 ( .A(n37114), .B(n37107), .Z(n55149) );
  NANDN U19801 ( .A(x[2939]), .B(y[2939]), .Z(n26611) );
  NANDN U19802 ( .A(x[2940]), .B(y[2940]), .Z(n26610) );
  AND U19803 ( .A(n26611), .B(n26610), .Z(n55148) );
  NANDN U19804 ( .A(y[2938]), .B(x[2938]), .Z(n9941) );
  NANDN U19805 ( .A(y[2939]), .B(x[2939]), .Z(n37108) );
  NAND U19806 ( .A(n9941), .B(n37108), .Z(n55147) );
  NANDN U19807 ( .A(x[2937]), .B(y[2937]), .Z(n55145) );
  NANDN U19808 ( .A(y[2936]), .B(x[2936]), .Z(n37095) );
  NANDN U19809 ( .A(y[2937]), .B(x[2937]), .Z(n37101) );
  AND U19810 ( .A(n37095), .B(n37101), .Z(n55144) );
  NANDN U19811 ( .A(x[2935]), .B(y[2935]), .Z(n26613) );
  NANDN U19812 ( .A(x[2936]), .B(y[2936]), .Z(n26612) );
  NAND U19813 ( .A(n26613), .B(n26612), .Z(n55143) );
  NANDN U19814 ( .A(y[2934]), .B(x[2934]), .Z(n37089) );
  NANDN U19815 ( .A(y[2935]), .B(x[2935]), .Z(n37096) );
  AND U19816 ( .A(n37089), .B(n37096), .Z(n55142) );
  NANDN U19817 ( .A(x[2933]), .B(y[2933]), .Z(n26615) );
  NANDN U19818 ( .A(x[2934]), .B(y[2934]), .Z(n26614) );
  NAND U19819 ( .A(n26615), .B(n26614), .Z(n55141) );
  NANDN U19820 ( .A(y[2932]), .B(x[2932]), .Z(n37083) );
  NANDN U19821 ( .A(y[2933]), .B(x[2933]), .Z(n37090) );
  NAND U19822 ( .A(n37083), .B(n37090), .Z(n55140) );
  NANDN U19823 ( .A(x[2931]), .B(y[2931]), .Z(n26617) );
  NANDN U19824 ( .A(x[2932]), .B(y[2932]), .Z(n26616) );
  AND U19825 ( .A(n26617), .B(n26616), .Z(n55139) );
  NANDN U19826 ( .A(y[2930]), .B(x[2930]), .Z(n37077) );
  NANDN U19827 ( .A(y[2931]), .B(x[2931]), .Z(n37084) );
  NAND U19828 ( .A(n37077), .B(n37084), .Z(n55138) );
  NANDN U19829 ( .A(x[2929]), .B(y[2929]), .Z(n26619) );
  NANDN U19830 ( .A(x[2930]), .B(y[2930]), .Z(n26618) );
  AND U19831 ( .A(n26619), .B(n26618), .Z(n55137) );
  NANDN U19832 ( .A(y[2928]), .B(x[2928]), .Z(n37071) );
  NANDN U19833 ( .A(y[2929]), .B(x[2929]), .Z(n37078) );
  NAND U19834 ( .A(n37071), .B(n37078), .Z(n55136) );
  NANDN U19835 ( .A(x[2927]), .B(y[2927]), .Z(n26621) );
  NANDN U19836 ( .A(x[2928]), .B(y[2928]), .Z(n26620) );
  NAND U19837 ( .A(n26621), .B(n26620), .Z(n55135) );
  NANDN U19838 ( .A(y[2926]), .B(x[2926]), .Z(n37065) );
  NANDN U19839 ( .A(y[2927]), .B(x[2927]), .Z(n37072) );
  AND U19840 ( .A(n37065), .B(n37072), .Z(n55134) );
  NANDN U19841 ( .A(x[2925]), .B(y[2925]), .Z(n26623) );
  NANDN U19842 ( .A(x[2926]), .B(y[2926]), .Z(n26622) );
  NAND U19843 ( .A(n26623), .B(n26622), .Z(n55133) );
  NANDN U19844 ( .A(y[2924]), .B(x[2924]), .Z(n37059) );
  NANDN U19845 ( .A(y[2925]), .B(x[2925]), .Z(n37066) );
  AND U19846 ( .A(n37059), .B(n37066), .Z(n55132) );
  NANDN U19847 ( .A(x[2923]), .B(y[2923]), .Z(n26625) );
  NANDN U19848 ( .A(x[2924]), .B(y[2924]), .Z(n26624) );
  NAND U19849 ( .A(n26625), .B(n26624), .Z(n55131) );
  NANDN U19850 ( .A(y[2922]), .B(x[2922]), .Z(n37053) );
  NANDN U19851 ( .A(y[2923]), .B(x[2923]), .Z(n37060) );
  NAND U19852 ( .A(n37053), .B(n37060), .Z(n55129) );
  NANDN U19853 ( .A(x[2921]), .B(y[2921]), .Z(n26627) );
  NANDN U19854 ( .A(x[2922]), .B(y[2922]), .Z(n26626) );
  AND U19855 ( .A(n26627), .B(n26626), .Z(n55128) );
  NANDN U19856 ( .A(y[2920]), .B(x[2920]), .Z(n37047) );
  NANDN U19857 ( .A(y[2921]), .B(x[2921]), .Z(n37054) );
  NAND U19858 ( .A(n37047), .B(n37054), .Z(n55127) );
  NANDN U19859 ( .A(x[2919]), .B(y[2919]), .Z(n26629) );
  NANDN U19860 ( .A(x[2920]), .B(y[2920]), .Z(n26628) );
  AND U19861 ( .A(n26629), .B(n26628), .Z(n55126) );
  NANDN U19862 ( .A(y[2918]), .B(x[2918]), .Z(n37041) );
  NANDN U19863 ( .A(y[2919]), .B(x[2919]), .Z(n37048) );
  NAND U19864 ( .A(n37041), .B(n37048), .Z(n55125) );
  NANDN U19865 ( .A(x[2917]), .B(y[2917]), .Z(n26631) );
  NANDN U19866 ( .A(x[2918]), .B(y[2918]), .Z(n26630) );
  NAND U19867 ( .A(n26631), .B(n26630), .Z(n55124) );
  NANDN U19868 ( .A(y[2916]), .B(x[2916]), .Z(n37035) );
  NANDN U19869 ( .A(y[2917]), .B(x[2917]), .Z(n37042) );
  AND U19870 ( .A(n37035), .B(n37042), .Z(n55123) );
  NANDN U19871 ( .A(x[2915]), .B(y[2915]), .Z(n26633) );
  NANDN U19872 ( .A(x[2916]), .B(y[2916]), .Z(n26632) );
  NAND U19873 ( .A(n26633), .B(n26632), .Z(n55122) );
  NANDN U19874 ( .A(y[2914]), .B(x[2914]), .Z(n26635) );
  NANDN U19875 ( .A(y[2915]), .B(x[2915]), .Z(n37036) );
  AND U19876 ( .A(n26635), .B(n37036), .Z(n55121) );
  ANDN U19877 ( .B(y[2913]), .A(x[2913]), .Z(n37028) );
  XNOR U19878 ( .A(y[2914]), .B(x[2914]), .Z(n9942) );
  NANDN U19879 ( .A(n37028), .B(n9942), .Z(n55120) );
  NANDN U19880 ( .A(y[2912]), .B(x[2912]), .Z(n26637) );
  NANDN U19881 ( .A(y[2913]), .B(x[2913]), .Z(n26636) );
  NAND U19882 ( .A(n26637), .B(n26636), .Z(n55119) );
  ANDN U19883 ( .B(y[2911]), .A(x[2911]), .Z(n37022) );
  ANDN U19884 ( .B(y[2912]), .A(x[2912]), .Z(n37029) );
  NOR U19885 ( .A(n37022), .B(n37029), .Z(n55118) );
  NANDN U19886 ( .A(y[2910]), .B(x[2910]), .Z(n9943) );
  NANDN U19887 ( .A(y[2911]), .B(x[2911]), .Z(n26638) );
  NAND U19888 ( .A(n9943), .B(n26638), .Z(n55117) );
  XNOR U19889 ( .A(y[2910]), .B(x[2910]), .Z(n26640) );
  NANDN U19890 ( .A(x[2909]), .B(y[2909]), .Z(n26641) );
  AND U19891 ( .A(n26640), .B(n26641), .Z(n55116) );
  NANDN U19892 ( .A(y[2908]), .B(x[2908]), .Z(n26643) );
  NANDN U19893 ( .A(y[2909]), .B(x[2909]), .Z(n26639) );
  NAND U19894 ( .A(n26643), .B(n26639), .Z(n55115) );
  NANDN U19895 ( .A(x[2907]), .B(y[2907]), .Z(n37012) );
  XNOR U19896 ( .A(x[2908]), .B(y[2908]), .Z(n9944) );
  NAND U19897 ( .A(n37012), .B(n9944), .Z(n55114) );
  NANDN U19898 ( .A(y[2906]), .B(x[2906]), .Z(n9945) );
  NANDN U19899 ( .A(y[2907]), .B(x[2907]), .Z(n26644) );
  AND U19900 ( .A(n9945), .B(n26644), .Z(n51990) );
  XNOR U19901 ( .A(y[2906]), .B(x[2906]), .Z(n37009) );
  NANDN U19902 ( .A(x[2905]), .B(y[2905]), .Z(n26645) );
  NAND U19903 ( .A(n37009), .B(n26645), .Z(n55112) );
  NANDN U19904 ( .A(y[2904]), .B(x[2904]), .Z(n26648) );
  ANDN U19905 ( .B(x[2905]), .A(y[2905]), .Z(n37008) );
  ANDN U19906 ( .B(n26648), .A(n37008), .Z(n55111) );
  NANDN U19907 ( .A(x[2903]), .B(y[2903]), .Z(n26649) );
  NANDN U19908 ( .A(x[2904]), .B(y[2904]), .Z(n26646) );
  NAND U19909 ( .A(n26649), .B(n26646), .Z(n55110) );
  NANDN U19910 ( .A(y[2902]), .B(x[2902]), .Z(n26651) );
  NANDN U19911 ( .A(y[2903]), .B(x[2903]), .Z(n26647) );
  NAND U19912 ( .A(n26651), .B(n26647), .Z(n55109) );
  NANDN U19913 ( .A(x[2901]), .B(y[2901]), .Z(n36995) );
  NANDN U19914 ( .A(x[2902]), .B(y[2902]), .Z(n26650) );
  AND U19915 ( .A(n36995), .B(n26650), .Z(n51991) );
  NANDN U19916 ( .A(y[2900]), .B(x[2900]), .Z(n26653) );
  NANDN U19917 ( .A(y[2901]), .B(x[2901]), .Z(n26652) );
  NAND U19918 ( .A(n26653), .B(n26652), .Z(n55108) );
  NANDN U19919 ( .A(x[2899]), .B(y[2899]), .Z(n36989) );
  NANDN U19920 ( .A(x[2900]), .B(y[2900]), .Z(n36996) );
  AND U19921 ( .A(n36989), .B(n36996), .Z(n55107) );
  NANDN U19922 ( .A(y[2898]), .B(x[2898]), .Z(n26655) );
  NANDN U19923 ( .A(y[2899]), .B(x[2899]), .Z(n26654) );
  NAND U19924 ( .A(n26655), .B(n26654), .Z(n55106) );
  NANDN U19925 ( .A(x[2897]), .B(y[2897]), .Z(n36983) );
  NANDN U19926 ( .A(x[2898]), .B(y[2898]), .Z(n36990) );
  NAND U19927 ( .A(n36983), .B(n36990), .Z(n55105) );
  NANDN U19928 ( .A(y[2896]), .B(x[2896]), .Z(n26657) );
  NANDN U19929 ( .A(y[2897]), .B(x[2897]), .Z(n26656) );
  AND U19930 ( .A(n26657), .B(n26656), .Z(n51992) );
  NANDN U19931 ( .A(x[2895]), .B(y[2895]), .Z(n36977) );
  NANDN U19932 ( .A(x[2896]), .B(y[2896]), .Z(n36984) );
  NAND U19933 ( .A(n36977), .B(n36984), .Z(n55104) );
  NANDN U19934 ( .A(y[2894]), .B(x[2894]), .Z(n26659) );
  NANDN U19935 ( .A(y[2895]), .B(x[2895]), .Z(n26658) );
  AND U19936 ( .A(n26659), .B(n26658), .Z(n55103) );
  NANDN U19937 ( .A(x[2893]), .B(y[2893]), .Z(n36971) );
  NANDN U19938 ( .A(x[2894]), .B(y[2894]), .Z(n36978) );
  NAND U19939 ( .A(n36971), .B(n36978), .Z(n55102) );
  NANDN U19940 ( .A(y[2892]), .B(x[2892]), .Z(n26661) );
  NANDN U19941 ( .A(y[2893]), .B(x[2893]), .Z(n26660) );
  NAND U19942 ( .A(n26661), .B(n26660), .Z(n55101) );
  NANDN U19943 ( .A(x[2891]), .B(y[2891]), .Z(n26663) );
  NANDN U19944 ( .A(x[2892]), .B(y[2892]), .Z(n36972) );
  AND U19945 ( .A(n26663), .B(n36972), .Z(n55098) );
  NANDN U19946 ( .A(x[2889]), .B(y[2889]), .Z(n14514) );
  ANDN U19947 ( .B(x[2889]), .A(y[2889]), .Z(n55095) );
  NANDN U19948 ( .A(y[2888]), .B(x[2888]), .Z(n55094) );
  NANDN U19949 ( .A(n55095), .B(n55094), .Z(n9946) );
  AND U19950 ( .A(n14514), .B(n9946), .Z(n14517) );
  NANDN U19951 ( .A(y[2884]), .B(x[2884]), .Z(n26668) );
  NANDN U19952 ( .A(y[2885]), .B(x[2885]), .Z(n26667) );
  NAND U19953 ( .A(n26668), .B(n26667), .Z(n55092) );
  NANDN U19954 ( .A(x[2883]), .B(y[2883]), .Z(n36948) );
  NANDN U19955 ( .A(x[2884]), .B(y[2884]), .Z(n36955) );
  AND U19956 ( .A(n36948), .B(n36955), .Z(n51996) );
  NANDN U19957 ( .A(y[2882]), .B(x[2882]), .Z(n26670) );
  NANDN U19958 ( .A(y[2883]), .B(x[2883]), .Z(n26669) );
  NAND U19959 ( .A(n26670), .B(n26669), .Z(n55091) );
  NANDN U19960 ( .A(x[2881]), .B(y[2881]), .Z(n36942) );
  NANDN U19961 ( .A(x[2882]), .B(y[2882]), .Z(n36949) );
  AND U19962 ( .A(n36942), .B(n36949), .Z(n55090) );
  NANDN U19963 ( .A(y[2880]), .B(x[2880]), .Z(n26672) );
  NANDN U19964 ( .A(y[2881]), .B(x[2881]), .Z(n26671) );
  NAND U19965 ( .A(n26672), .B(n26671), .Z(n55088) );
  NANDN U19966 ( .A(x[2879]), .B(y[2879]), .Z(n36936) );
  NANDN U19967 ( .A(x[2880]), .B(y[2880]), .Z(n36943) );
  AND U19968 ( .A(n36936), .B(n36943), .Z(n55087) );
  NANDN U19969 ( .A(y[2878]), .B(x[2878]), .Z(n26674) );
  NANDN U19970 ( .A(y[2879]), .B(x[2879]), .Z(n26673) );
  NAND U19971 ( .A(n26674), .B(n26673), .Z(n55086) );
  NANDN U19972 ( .A(x[2877]), .B(y[2877]), .Z(n26676) );
  XNOR U19973 ( .A(x[2878]), .B(y[2878]), .Z(n9947) );
  AND U19974 ( .A(n26676), .B(n9947), .Z(n51997) );
  NANDN U19975 ( .A(y[2874]), .B(x[2874]), .Z(n9948) );
  NANDN U19976 ( .A(y[2875]), .B(x[2875]), .Z(n26679) );
  NAND U19977 ( .A(n9948), .B(n26679), .Z(n55084) );
  XNOR U19978 ( .A(y[2874]), .B(x[2874]), .Z(n26680) );
  NANDN U19979 ( .A(x[2873]), .B(y[2873]), .Z(n26682) );
  NAND U19980 ( .A(n26680), .B(n26682), .Z(n55083) );
  NANDN U19981 ( .A(y[2872]), .B(x[2872]), .Z(n26684) );
  NANDN U19982 ( .A(y[2873]), .B(x[2873]), .Z(n26681) );
  AND U19983 ( .A(n26684), .B(n26681), .Z(n51999) );
  NANDN U19984 ( .A(x[2869]), .B(y[2869]), .Z(n36909) );
  NANDN U19985 ( .A(x[2870]), .B(y[2870]), .Z(n36916) );
  NAND U19986 ( .A(n36909), .B(n36916), .Z(n55080) );
  NANDN U19987 ( .A(y[2868]), .B(x[2868]), .Z(n26688) );
  NANDN U19988 ( .A(y[2869]), .B(x[2869]), .Z(n26687) );
  NAND U19989 ( .A(n26688), .B(n26687), .Z(n55079) );
  NANDN U19990 ( .A(x[2867]), .B(y[2867]), .Z(n36903) );
  NANDN U19991 ( .A(x[2868]), .B(y[2868]), .Z(n36910) );
  AND U19992 ( .A(n36903), .B(n36910), .Z(n52001) );
  NANDN U19993 ( .A(y[2864]), .B(x[2864]), .Z(n26692) );
  NANDN U19994 ( .A(y[2865]), .B(x[2865]), .Z(n26691) );
  NAND U19995 ( .A(n26692), .B(n26691), .Z(n55076) );
  NANDN U19996 ( .A(x[2863]), .B(y[2863]), .Z(n36891) );
  NANDN U19997 ( .A(x[2864]), .B(y[2864]), .Z(n36898) );
  NAND U19998 ( .A(n36891), .B(n36898), .Z(n55075) );
  NANDN U19999 ( .A(y[2862]), .B(x[2862]), .Z(n36888) );
  NANDN U20000 ( .A(y[2863]), .B(x[2863]), .Z(n26693) );
  AND U20001 ( .A(n36888), .B(n26693), .Z(n52003) );
  NANDN U20002 ( .A(x[2859]), .B(y[2859]), .Z(n26696) );
  NANDN U20003 ( .A(x[2860]), .B(y[2860]), .Z(n26695) );
  NAND U20004 ( .A(n26696), .B(n26695), .Z(n55073) );
  NANDN U20005 ( .A(y[2858]), .B(x[2858]), .Z(n36876) );
  NANDN U20006 ( .A(y[2859]), .B(x[2859]), .Z(n36883) );
  NAND U20007 ( .A(n36876), .B(n36883), .Z(n55072) );
  NANDN U20008 ( .A(x[2858]), .B(y[2858]), .Z(n26697) );
  ANDN U20009 ( .B(y[2857]), .A(x[2857]), .Z(n36872) );
  ANDN U20010 ( .B(n26697), .A(n36872), .Z(n55071) );
  NANDN U20011 ( .A(x[2855]), .B(y[2855]), .Z(n26698) );
  ANDN U20012 ( .B(y[2856]), .A(x[2856]), .Z(n36874) );
  ANDN U20013 ( .B(n26698), .A(n36874), .Z(n55068) );
  NANDN U20014 ( .A(y[2852]), .B(x[2852]), .Z(n36855) );
  NANDN U20015 ( .A(y[2853]), .B(x[2853]), .Z(n36862) );
  NAND U20016 ( .A(n36855), .B(n36862), .Z(n55066) );
  NANDN U20017 ( .A(x[2849]), .B(y[2849]), .Z(n36845) );
  NANDN U20018 ( .A(x[2850]), .B(y[2850]), .Z(n26703) );
  NAND U20019 ( .A(n36845), .B(n26703), .Z(n55063) );
  NANDN U20020 ( .A(y[2848]), .B(x[2848]), .Z(n36842) );
  NANDN U20021 ( .A(y[2849]), .B(x[2849]), .Z(n36850) );
  NAND U20022 ( .A(n36842), .B(n36850), .Z(n55062) );
  NANDN U20023 ( .A(x[2847]), .B(y[2847]), .Z(n26704) );
  NANDN U20024 ( .A(x[2848]), .B(y[2848]), .Z(n36846) );
  AND U20025 ( .A(n26704), .B(n36846), .Z(n52007) );
  XNOR U20026 ( .A(x[2846]), .B(y[2846]), .Z(n9949) );
  ANDN U20027 ( .B(y[2845]), .A(x[2845]), .Z(n36834) );
  ANDN U20028 ( .B(n9949), .A(n36834), .Z(n55061) );
  NANDN U20029 ( .A(y[2844]), .B(x[2844]), .Z(n26708) );
  NANDN U20030 ( .A(y[2845]), .B(x[2845]), .Z(n26707) );
  NAND U20031 ( .A(n26708), .B(n26707), .Z(n55060) );
  NANDN U20032 ( .A(y[2842]), .B(x[2842]), .Z(n9950) );
  NANDN U20033 ( .A(y[2843]), .B(x[2843]), .Z(n26709) );
  AND U20034 ( .A(n9950), .B(n26709), .Z(n55057) );
  XNOR U20035 ( .A(y[2842]), .B(x[2842]), .Z(n26711) );
  NANDN U20036 ( .A(x[2841]), .B(y[2841]), .Z(n26712) );
  NAND U20037 ( .A(n26711), .B(n26712), .Z(n55056) );
  NANDN U20038 ( .A(y[2840]), .B(x[2840]), .Z(n26714) );
  NANDN U20039 ( .A(y[2841]), .B(x[2841]), .Z(n26710) );
  AND U20040 ( .A(n26714), .B(n26710), .Z(n52009) );
  XNOR U20041 ( .A(y[2838]), .B(x[2838]), .Z(n26716) );
  NANDN U20042 ( .A(x[2837]), .B(y[2837]), .Z(n26718) );
  NAND U20043 ( .A(n26716), .B(n26718), .Z(n55054) );
  NANDN U20044 ( .A(y[2836]), .B(x[2836]), .Z(n9951) );
  NANDN U20045 ( .A(y[2837]), .B(x[2837]), .Z(n26717) );
  AND U20046 ( .A(n9951), .B(n26717), .Z(n52011) );
  NANDN U20047 ( .A(x[2835]), .B(y[2835]), .Z(n55052) );
  NANDN U20048 ( .A(y[2834]), .B(x[2834]), .Z(n26721) );
  NANDN U20049 ( .A(y[2835]), .B(x[2835]), .Z(n26719) );
  AND U20050 ( .A(n26721), .B(n26719), .Z(n55051) );
  NANDN U20051 ( .A(x[2833]), .B(y[2833]), .Z(n36802) );
  NANDN U20052 ( .A(x[2834]), .B(y[2834]), .Z(n36808) );
  NAND U20053 ( .A(n36802), .B(n36808), .Z(n55050) );
  NANDN U20054 ( .A(y[2832]), .B(x[2832]), .Z(n26723) );
  NANDN U20055 ( .A(y[2833]), .B(x[2833]), .Z(n26722) );
  AND U20056 ( .A(n26723), .B(n26722), .Z(n55049) );
  NANDN U20057 ( .A(x[2831]), .B(y[2831]), .Z(n36796) );
  NANDN U20058 ( .A(x[2832]), .B(y[2832]), .Z(n36803) );
  NAND U20059 ( .A(n36796), .B(n36803), .Z(n55048) );
  NANDN U20060 ( .A(y[2830]), .B(x[2830]), .Z(n26725) );
  NANDN U20061 ( .A(y[2831]), .B(x[2831]), .Z(n26724) );
  NAND U20062 ( .A(n26725), .B(n26724), .Z(n55047) );
  NANDN U20063 ( .A(x[2829]), .B(y[2829]), .Z(n36790) );
  NANDN U20064 ( .A(x[2830]), .B(y[2830]), .Z(n36797) );
  AND U20065 ( .A(n36790), .B(n36797), .Z(n55045) );
  NANDN U20066 ( .A(y[2828]), .B(x[2828]), .Z(n36786) );
  NANDN U20067 ( .A(y[2829]), .B(x[2829]), .Z(n26726) );
  NAND U20068 ( .A(n36786), .B(n26726), .Z(n55044) );
  NANDN U20069 ( .A(x[2827]), .B(y[2827]), .Z(n36783) );
  NANDN U20070 ( .A(x[2828]), .B(y[2828]), .Z(n36791) );
  AND U20071 ( .A(n36783), .B(n36791), .Z(n55043) );
  NANDN U20072 ( .A(y[2826]), .B(x[2826]), .Z(n26727) );
  NANDN U20073 ( .A(y[2827]), .B(x[2827]), .Z(n36787) );
  NAND U20074 ( .A(n26727), .B(n36787), .Z(n55042) );
  NANDN U20075 ( .A(x[2825]), .B(y[2825]), .Z(n26729) );
  NANDN U20076 ( .A(x[2826]), .B(y[2826]), .Z(n36785) );
  NAND U20077 ( .A(n26729), .B(n36785), .Z(n55041) );
  NANDN U20078 ( .A(y[2824]), .B(x[2824]), .Z(n36775) );
  NANDN U20079 ( .A(y[2825]), .B(x[2825]), .Z(n26728) );
  AND U20080 ( .A(n36775), .B(n26728), .Z(n55040) );
  NANDN U20081 ( .A(x[2823]), .B(y[2823]), .Z(n26731) );
  NANDN U20082 ( .A(x[2824]), .B(y[2824]), .Z(n26730) );
  NAND U20083 ( .A(n26731), .B(n26730), .Z(n55039) );
  NANDN U20084 ( .A(y[2822]), .B(x[2822]), .Z(n9952) );
  ANDN U20085 ( .B(x[2823]), .A(y[2823]), .Z(n36777) );
  ANDN U20086 ( .B(n9952), .A(n36777), .Z(n55038) );
  XNOR U20087 ( .A(x[2822]), .B(y[2822]), .Z(n36769) );
  NANDN U20088 ( .A(y[2820]), .B(x[2820]), .Z(n26734) );
  NANDN U20089 ( .A(y[2821]), .B(x[2821]), .Z(n36770) );
  AND U20090 ( .A(n26734), .B(n36770), .Z(n55036) );
  NANDN U20091 ( .A(x[2819]), .B(y[2819]), .Z(n26736) );
  NANDN U20092 ( .A(x[2820]), .B(y[2820]), .Z(n26733) );
  NAND U20093 ( .A(n26736), .B(n26733), .Z(n55035) );
  NANDN U20094 ( .A(y[2818]), .B(x[2818]), .Z(n9953) );
  NANDN U20095 ( .A(y[2819]), .B(x[2819]), .Z(n26735) );
  AND U20096 ( .A(n9953), .B(n26735), .Z(n52013) );
  ANDN U20097 ( .B(y[2817]), .A(x[2817]), .Z(n26739) );
  XNOR U20098 ( .A(x[2818]), .B(y[2818]), .Z(n26738) );
  NANDN U20099 ( .A(y[2816]), .B(x[2816]), .Z(n9954) );
  NANDN U20100 ( .A(y[2817]), .B(x[2817]), .Z(n26737) );
  NAND U20101 ( .A(n9954), .B(n26737), .Z(n55032) );
  NANDN U20102 ( .A(x[2815]), .B(y[2815]), .Z(n55030) );
  XNOR U20103 ( .A(x[2816]), .B(y[2816]), .Z(n36755) );
  NANDN U20104 ( .A(y[2814]), .B(x[2814]), .Z(n36748) );
  NANDN U20105 ( .A(y[2815]), .B(x[2815]), .Z(n36754) );
  NAND U20106 ( .A(n36748), .B(n36754), .Z(n55028) );
  NANDN U20107 ( .A(x[2813]), .B(y[2813]), .Z(n26741) );
  NANDN U20108 ( .A(x[2814]), .B(y[2814]), .Z(n26740) );
  AND U20109 ( .A(n26741), .B(n26740), .Z(n55027) );
  NANDN U20110 ( .A(y[2812]), .B(x[2812]), .Z(n36742) );
  NANDN U20111 ( .A(y[2813]), .B(x[2813]), .Z(n36749) );
  NAND U20112 ( .A(n36742), .B(n36749), .Z(n55026) );
  NANDN U20113 ( .A(x[2811]), .B(y[2811]), .Z(n26743) );
  NANDN U20114 ( .A(x[2812]), .B(y[2812]), .Z(n26742) );
  AND U20115 ( .A(n26743), .B(n26742), .Z(n55025) );
  NANDN U20116 ( .A(y[2810]), .B(x[2810]), .Z(n36736) );
  NANDN U20117 ( .A(y[2811]), .B(x[2811]), .Z(n36743) );
  NAND U20118 ( .A(n36736), .B(n36743), .Z(n55024) );
  NANDN U20119 ( .A(x[2809]), .B(y[2809]), .Z(n26745) );
  NANDN U20120 ( .A(x[2810]), .B(y[2810]), .Z(n26744) );
  NAND U20121 ( .A(n26745), .B(n26744), .Z(n55023) );
  NANDN U20122 ( .A(y[2808]), .B(x[2808]), .Z(n36730) );
  NANDN U20123 ( .A(y[2809]), .B(x[2809]), .Z(n36737) );
  AND U20124 ( .A(n36730), .B(n36737), .Z(n55022) );
  NANDN U20125 ( .A(x[2807]), .B(y[2807]), .Z(n26747) );
  NANDN U20126 ( .A(x[2808]), .B(y[2808]), .Z(n26746) );
  NAND U20127 ( .A(n26747), .B(n26746), .Z(n55021) );
  NANDN U20128 ( .A(y[2806]), .B(x[2806]), .Z(n36724) );
  NANDN U20129 ( .A(y[2807]), .B(x[2807]), .Z(n36731) );
  AND U20130 ( .A(n36724), .B(n36731), .Z(n55020) );
  NANDN U20131 ( .A(x[2805]), .B(y[2805]), .Z(n36721) );
  NANDN U20132 ( .A(x[2806]), .B(y[2806]), .Z(n26748) );
  NAND U20133 ( .A(n36721), .B(n26748), .Z(n55019) );
  NANDN U20134 ( .A(y[2804]), .B(x[2804]), .Z(n26749) );
  NANDN U20135 ( .A(y[2805]), .B(x[2805]), .Z(n36725) );
  NAND U20136 ( .A(n26749), .B(n36725), .Z(n55018) );
  NANDN U20137 ( .A(x[2803]), .B(y[2803]), .Z(n36715) );
  NANDN U20138 ( .A(x[2804]), .B(y[2804]), .Z(n36722) );
  AND U20139 ( .A(n36715), .B(n36722), .Z(n52014) );
  NANDN U20140 ( .A(x[2801]), .B(y[2801]), .Z(n36709) );
  NANDN U20141 ( .A(x[2802]), .B(y[2802]), .Z(n36716) );
  AND U20142 ( .A(n36709), .B(n36716), .Z(n55016) );
  NANDN U20143 ( .A(y[2800]), .B(x[2800]), .Z(n26753) );
  NANDN U20144 ( .A(y[2801]), .B(x[2801]), .Z(n26752) );
  NAND U20145 ( .A(n26753), .B(n26752), .Z(n55015) );
  NANDN U20146 ( .A(x[2799]), .B(y[2799]), .Z(n26755) );
  NANDN U20147 ( .A(x[2800]), .B(y[2800]), .Z(n36710) );
  NAND U20148 ( .A(n26755), .B(n36710), .Z(n55013) );
  NANDN U20149 ( .A(y[2799]), .B(x[2799]), .Z(n26754) );
  ANDN U20150 ( .B(x[2798]), .A(y[2798]), .Z(n36703) );
  ANDN U20151 ( .B(n26754), .A(n36703), .Z(n55012) );
  NANDN U20152 ( .A(x[2797]), .B(y[2797]), .Z(n36701) );
  NANDN U20153 ( .A(x[2798]), .B(y[2798]), .Z(n26756) );
  NAND U20154 ( .A(n36701), .B(n26756), .Z(n55011) );
  NANDN U20155 ( .A(x[2796]), .B(y[2796]), .Z(n36698) );
  NANDN U20156 ( .A(x[2795]), .B(y[2795]), .Z(n26757) );
  NAND U20157 ( .A(n36698), .B(n26757), .Z(n55009) );
  NANDN U20158 ( .A(y[2795]), .B(x[2795]), .Z(n36696) );
  NANDN U20159 ( .A(y[2794]), .B(x[2794]), .Z(n36690) );
  NAND U20160 ( .A(n36696), .B(n36690), .Z(n55008) );
  NANDN U20161 ( .A(x[2794]), .B(y[2794]), .Z(n26758) );
  ANDN U20162 ( .B(y[2793]), .A(x[2793]), .Z(n36688) );
  ANDN U20163 ( .B(n26758), .A(n36688), .Z(n55007) );
  NANDN U20164 ( .A(y[2792]), .B(x[2792]), .Z(n9955) );
  NANDN U20165 ( .A(y[2793]), .B(x[2793]), .Z(n36691) );
  NAND U20166 ( .A(n9955), .B(n36691), .Z(n55006) );
  XNOR U20167 ( .A(y[2792]), .B(x[2792]), .Z(n26760) );
  ANDN U20168 ( .B(y[2791]), .A(x[2791]), .Z(n26761) );
  ANDN U20169 ( .B(n26760), .A(n26761), .Z(n55005) );
  NANDN U20170 ( .A(y[2790]), .B(x[2790]), .Z(n9956) );
  NANDN U20171 ( .A(y[2791]), .B(x[2791]), .Z(n26759) );
  NAND U20172 ( .A(n9956), .B(n26759), .Z(n55004) );
  ANDN U20173 ( .B(y[2789]), .A(x[2789]), .Z(n26762) );
  NANDN U20174 ( .A(x[2787]), .B(y[2787]), .Z(n36668) );
  NANDN U20175 ( .A(x[2788]), .B(y[2788]), .Z(n26763) );
  NAND U20176 ( .A(n36668), .B(n26763), .Z(n52017) );
  NANDN U20177 ( .A(y[2786]), .B(x[2786]), .Z(n36663) );
  NANDN U20178 ( .A(y[2787]), .B(x[2787]), .Z(n36672) );
  NAND U20179 ( .A(n36663), .B(n36672), .Z(n55002) );
  NANDN U20180 ( .A(x[2785]), .B(y[2785]), .Z(n26764) );
  NANDN U20181 ( .A(x[2786]), .B(y[2786]), .Z(n36669) );
  AND U20182 ( .A(n26764), .B(n36669), .Z(n55001) );
  NANDN U20183 ( .A(y[2784]), .B(x[2784]), .Z(n36657) );
  NANDN U20184 ( .A(y[2785]), .B(x[2785]), .Z(n36664) );
  NAND U20185 ( .A(n36657), .B(n36664), .Z(n54999) );
  NANDN U20186 ( .A(x[2783]), .B(y[2783]), .Z(n36653) );
  NANDN U20187 ( .A(x[2784]), .B(y[2784]), .Z(n26765) );
  AND U20188 ( .A(n36653), .B(n26765), .Z(n54998) );
  NANDN U20189 ( .A(y[2782]), .B(x[2782]), .Z(n26766) );
  NANDN U20190 ( .A(y[2783]), .B(x[2783]), .Z(n36658) );
  NAND U20191 ( .A(n26766), .B(n36658), .Z(n54996) );
  ANDN U20192 ( .B(y[2781]), .A(x[2781]), .Z(n36648) );
  NANDN U20193 ( .A(x[2782]), .B(y[2782]), .Z(n36654) );
  NANDN U20194 ( .A(n36648), .B(n36654), .Z(n54994) );
  NANDN U20195 ( .A(y[2780]), .B(x[2780]), .Z(n26768) );
  NANDN U20196 ( .A(y[2781]), .B(x[2781]), .Z(n26767) );
  AND U20197 ( .A(n26768), .B(n26767), .Z(n54992) );
  ANDN U20198 ( .B(y[2779]), .A(x[2779]), .Z(n36643) );
  ANDN U20199 ( .B(y[2780]), .A(x[2780]), .Z(n36649) );
  OR U20200 ( .A(n36643), .B(n36649), .Z(n54990) );
  NANDN U20201 ( .A(y[2778]), .B(x[2778]), .Z(n9957) );
  NANDN U20202 ( .A(y[2779]), .B(x[2779]), .Z(n26769) );
  AND U20203 ( .A(n9957), .B(n26769), .Z(n54988) );
  ANDN U20204 ( .B(y[2777]), .A(x[2777]), .Z(n54984) );
  XNOR U20205 ( .A(x[2778]), .B(y[2778]), .Z(n26771) );
  NANDN U20206 ( .A(y[2776]), .B(x[2776]), .Z(n9958) );
  NANDN U20207 ( .A(y[2777]), .B(x[2777]), .Z(n26770) );
  AND U20208 ( .A(n9958), .B(n26770), .Z(n54982) );
  NANDN U20209 ( .A(y[2774]), .B(x[2774]), .Z(n26775) );
  NANDN U20210 ( .A(y[2775]), .B(x[2775]), .Z(n26772) );
  AND U20211 ( .A(n26775), .B(n26772), .Z(n54976) );
  NANDN U20212 ( .A(x[2773]), .B(y[2773]), .Z(n36628) );
  NANDN U20213 ( .A(x[2774]), .B(y[2774]), .Z(n26774) );
  NAND U20214 ( .A(n36628), .B(n26774), .Z(n54974) );
  NANDN U20215 ( .A(y[2772]), .B(x[2772]), .Z(n26777) );
  NANDN U20216 ( .A(y[2773]), .B(x[2773]), .Z(n26776) );
  NAND U20217 ( .A(n26777), .B(n26776), .Z(n54972) );
  NANDN U20218 ( .A(x[2771]), .B(y[2771]), .Z(n36622) );
  NANDN U20219 ( .A(x[2772]), .B(y[2772]), .Z(n36629) );
  AND U20220 ( .A(n36622), .B(n36629), .Z(n54970) );
  NANDN U20221 ( .A(y[2770]), .B(x[2770]), .Z(n36619) );
  NANDN U20222 ( .A(y[2771]), .B(x[2771]), .Z(n26778) );
  NAND U20223 ( .A(n36619), .B(n26778), .Z(n54968) );
  NANDN U20224 ( .A(x[2769]), .B(y[2769]), .Z(n26779) );
  NANDN U20225 ( .A(x[2770]), .B(y[2770]), .Z(n36623) );
  AND U20226 ( .A(n26779), .B(n36623), .Z(n54966) );
  NANDN U20227 ( .A(y[2768]), .B(x[2768]), .Z(n9959) );
  NANDN U20228 ( .A(y[2769]), .B(x[2769]), .Z(n36620) );
  NAND U20229 ( .A(n9959), .B(n36620), .Z(n54964) );
  NANDN U20230 ( .A(x[2767]), .B(y[2767]), .Z(n54959) );
  NANDN U20231 ( .A(y[2766]), .B(x[2766]), .Z(n36607) );
  NANDN U20232 ( .A(y[2767]), .B(x[2767]), .Z(n36614) );
  AND U20233 ( .A(n36607), .B(n36614), .Z(n54957) );
  ANDN U20234 ( .B(y[2765]), .A(x[2765]), .Z(n36603) );
  NANDN U20235 ( .A(x[2766]), .B(y[2766]), .Z(n26780) );
  NANDN U20236 ( .A(n36603), .B(n26780), .Z(n54956) );
  NANDN U20237 ( .A(y[2764]), .B(x[2764]), .Z(n9960) );
  NANDN U20238 ( .A(y[2765]), .B(x[2765]), .Z(n36608) );
  AND U20239 ( .A(n9960), .B(n36608), .Z(n54955) );
  XNOR U20240 ( .A(y[2764]), .B(x[2764]), .Z(n36599) );
  NANDN U20241 ( .A(x[2763]), .B(y[2763]), .Z(n26781) );
  NAND U20242 ( .A(n36599), .B(n26781), .Z(n54954) );
  NANDN U20243 ( .A(y[2762]), .B(x[2762]), .Z(n36592) );
  NANDN U20244 ( .A(y[2763]), .B(x[2763]), .Z(n36601) );
  NAND U20245 ( .A(n36592), .B(n36601), .Z(n54953) );
  NANDN U20246 ( .A(x[2761]), .B(y[2761]), .Z(n26783) );
  NANDN U20247 ( .A(x[2762]), .B(y[2762]), .Z(n26782) );
  AND U20248 ( .A(n26783), .B(n26782), .Z(n52018) );
  XNOR U20249 ( .A(y[2760]), .B(x[2760]), .Z(n36587) );
  NANDN U20250 ( .A(x[2759]), .B(y[2759]), .Z(n36583) );
  AND U20251 ( .A(n36587), .B(n36583), .Z(n54951) );
  NANDN U20252 ( .A(y[2758]), .B(x[2758]), .Z(n26785) );
  NANDN U20253 ( .A(y[2759]), .B(x[2759]), .Z(n36586) );
  NAND U20254 ( .A(n26785), .B(n36586), .Z(n54950) );
  NANDN U20255 ( .A(x[2757]), .B(y[2757]), .Z(n36577) );
  NANDN U20256 ( .A(x[2758]), .B(y[2758]), .Z(n36584) );
  NAND U20257 ( .A(n36577), .B(n36584), .Z(n54949) );
  NANDN U20258 ( .A(y[2756]), .B(x[2756]), .Z(n26787) );
  NANDN U20259 ( .A(y[2757]), .B(x[2757]), .Z(n26786) );
  AND U20260 ( .A(n26787), .B(n26786), .Z(n54948) );
  NANDN U20261 ( .A(x[2755]), .B(y[2755]), .Z(n36571) );
  NANDN U20262 ( .A(x[2756]), .B(y[2756]), .Z(n36578) );
  NAND U20263 ( .A(n36571), .B(n36578), .Z(n54947) );
  NANDN U20264 ( .A(y[2754]), .B(x[2754]), .Z(n26789) );
  NANDN U20265 ( .A(y[2755]), .B(x[2755]), .Z(n26788) );
  AND U20266 ( .A(n26789), .B(n26788), .Z(n54946) );
  NANDN U20267 ( .A(x[2753]), .B(y[2753]), .Z(n36565) );
  NANDN U20268 ( .A(x[2754]), .B(y[2754]), .Z(n36572) );
  NAND U20269 ( .A(n36565), .B(n36572), .Z(n54945) );
  NANDN U20270 ( .A(y[2752]), .B(x[2752]), .Z(n26791) );
  NANDN U20271 ( .A(y[2753]), .B(x[2753]), .Z(n26790) );
  NAND U20272 ( .A(n26791), .B(n26790), .Z(n54944) );
  NANDN U20273 ( .A(x[2751]), .B(y[2751]), .Z(n36559) );
  NANDN U20274 ( .A(x[2752]), .B(y[2752]), .Z(n36566) );
  AND U20275 ( .A(n36559), .B(n36566), .Z(n54943) );
  NANDN U20276 ( .A(y[2750]), .B(x[2750]), .Z(n9961) );
  NANDN U20277 ( .A(y[2751]), .B(x[2751]), .Z(n26792) );
  NAND U20278 ( .A(n9961), .B(n26792), .Z(n54942) );
  NANDN U20279 ( .A(x[2749]), .B(y[2749]), .Z(n52019) );
  XNOR U20280 ( .A(x[2750]), .B(y[2750]), .Z(n36557) );
  AND U20281 ( .A(n52019), .B(n36557), .Z(n14361) );
  NANDN U20282 ( .A(y[2748]), .B(x[2748]), .Z(n26794) );
  ANDN U20283 ( .B(x[2749]), .A(y[2749]), .Z(n36556) );
  ANDN U20284 ( .B(n26794), .A(n36556), .Z(n54940) );
  NANDN U20285 ( .A(x[2747]), .B(y[2747]), .Z(n26796) );
  NANDN U20286 ( .A(x[2748]), .B(y[2748]), .Z(n26793) );
  NAND U20287 ( .A(n26796), .B(n26793), .Z(n54939) );
  NANDN U20288 ( .A(y[2747]), .B(x[2747]), .Z(n26795) );
  ANDN U20289 ( .B(x[2746]), .A(y[2746]), .Z(n36546) );
  ANDN U20290 ( .B(n26795), .A(n36546), .Z(n54938) );
  NANDN U20291 ( .A(x[2745]), .B(y[2745]), .Z(n26798) );
  NANDN U20292 ( .A(x[2746]), .B(y[2746]), .Z(n26797) );
  NAND U20293 ( .A(n26798), .B(n26797), .Z(n54937) );
  ANDN U20294 ( .B(x[2744]), .A(y[2744]), .Z(n36542) );
  ANDN U20295 ( .B(x[2745]), .A(y[2745]), .Z(n36547) );
  NOR U20296 ( .A(n36542), .B(n36547), .Z(n54936) );
  NANDN U20297 ( .A(x[2743]), .B(y[2743]), .Z(n36540) );
  NANDN U20298 ( .A(x[2744]), .B(y[2744]), .Z(n26799) );
  NAND U20299 ( .A(n36540), .B(n26799), .Z(n54935) );
  NANDN U20300 ( .A(x[2741]), .B(y[2741]), .Z(n9962) );
  ANDN U20301 ( .B(y[2742]), .A(x[2742]), .Z(n36535) );
  ANDN U20302 ( .B(n9962), .A(n36535), .Z(n54933) );
  NANDN U20303 ( .A(y[2740]), .B(x[2740]), .Z(n26801) );
  NANDN U20304 ( .A(y[2741]), .B(x[2741]), .Z(n36534) );
  NAND U20305 ( .A(n26801), .B(n36534), .Z(n54932) );
  NANDN U20306 ( .A(x[2740]), .B(y[2740]), .Z(n26800) );
  ANDN U20307 ( .B(y[2739]), .A(x[2739]), .Z(n36527) );
  ANDN U20308 ( .B(n26800), .A(n36527), .Z(n54931) );
  NANDN U20309 ( .A(x[2737]), .B(y[2737]), .Z(n26806) );
  NANDN U20310 ( .A(x[2738]), .B(y[2738]), .Z(n36528) );
  AND U20311 ( .A(n26806), .B(n36528), .Z(n14346) );
  ANDN U20312 ( .B(x[2737]), .A(y[2737]), .Z(n26803) );
  NANDN U20313 ( .A(x[2736]), .B(y[2736]), .Z(n26805) );
  NANDN U20314 ( .A(y[2734]), .B(x[2734]), .Z(n26809) );
  NANDN U20315 ( .A(y[2735]), .B(x[2735]), .Z(n26808) );
  NAND U20316 ( .A(n26809), .B(n26808), .Z(n54924) );
  NANDN U20317 ( .A(x[2733]), .B(y[2733]), .Z(n36512) );
  NANDN U20318 ( .A(x[2734]), .B(y[2734]), .Z(n36518) );
  AND U20319 ( .A(n36512), .B(n36518), .Z(n54922) );
  NANDN U20320 ( .A(y[2732]), .B(x[2732]), .Z(n26811) );
  NANDN U20321 ( .A(y[2733]), .B(x[2733]), .Z(n26810) );
  NAND U20322 ( .A(n26811), .B(n26810), .Z(n54920) );
  NANDN U20323 ( .A(x[2731]), .B(y[2731]), .Z(n36506) );
  NANDN U20324 ( .A(x[2732]), .B(y[2732]), .Z(n36513) );
  AND U20325 ( .A(n36506), .B(n36513), .Z(n54918) );
  NANDN U20326 ( .A(y[2730]), .B(x[2730]), .Z(n26813) );
  NANDN U20327 ( .A(y[2731]), .B(x[2731]), .Z(n26812) );
  NAND U20328 ( .A(n26813), .B(n26812), .Z(n54916) );
  NANDN U20329 ( .A(x[2729]), .B(y[2729]), .Z(n36500) );
  NANDN U20330 ( .A(x[2730]), .B(y[2730]), .Z(n36507) );
  NAND U20331 ( .A(n36500), .B(n36507), .Z(n54914) );
  NANDN U20332 ( .A(y[2728]), .B(x[2728]), .Z(n26815) );
  NANDN U20333 ( .A(y[2729]), .B(x[2729]), .Z(n26814) );
  AND U20334 ( .A(n26815), .B(n26814), .Z(n54912) );
  NANDN U20335 ( .A(x[2727]), .B(y[2727]), .Z(n36494) );
  NANDN U20336 ( .A(x[2728]), .B(y[2728]), .Z(n36501) );
  NAND U20337 ( .A(n36494), .B(n36501), .Z(n54910) );
  NANDN U20338 ( .A(y[2726]), .B(x[2726]), .Z(n26817) );
  NANDN U20339 ( .A(y[2727]), .B(x[2727]), .Z(n26816) );
  AND U20340 ( .A(n26817), .B(n26816), .Z(n54908) );
  NANDN U20341 ( .A(x[2725]), .B(y[2725]), .Z(n36488) );
  NANDN U20342 ( .A(x[2726]), .B(y[2726]), .Z(n36495) );
  NAND U20343 ( .A(n36488), .B(n36495), .Z(n54906) );
  NANDN U20344 ( .A(y[2724]), .B(x[2724]), .Z(n26819) );
  NANDN U20345 ( .A(y[2725]), .B(x[2725]), .Z(n26818) );
  NAND U20346 ( .A(n26819), .B(n26818), .Z(n54904) );
  NANDN U20347 ( .A(x[2723]), .B(y[2723]), .Z(n36482) );
  NANDN U20348 ( .A(x[2724]), .B(y[2724]), .Z(n36489) );
  AND U20349 ( .A(n36482), .B(n36489), .Z(n54902) );
  NANDN U20350 ( .A(y[2722]), .B(x[2722]), .Z(n26821) );
  NANDN U20351 ( .A(y[2723]), .B(x[2723]), .Z(n26820) );
  NAND U20352 ( .A(n26821), .B(n26820), .Z(n54900) );
  NANDN U20353 ( .A(x[2721]), .B(y[2721]), .Z(n36476) );
  NANDN U20354 ( .A(x[2722]), .B(y[2722]), .Z(n36483) );
  AND U20355 ( .A(n36476), .B(n36483), .Z(n54898) );
  NANDN U20356 ( .A(y[2720]), .B(x[2720]), .Z(n36473) );
  NANDN U20357 ( .A(y[2721]), .B(x[2721]), .Z(n26822) );
  NAND U20358 ( .A(n36473), .B(n26822), .Z(n54896) );
  NANDN U20359 ( .A(x[2719]), .B(y[2719]), .Z(n26823) );
  NANDN U20360 ( .A(x[2720]), .B(y[2720]), .Z(n36477) );
  NAND U20361 ( .A(n26823), .B(n36477), .Z(n54894) );
  NANDN U20362 ( .A(y[2718]), .B(x[2718]), .Z(n36467) );
  NANDN U20363 ( .A(y[2719]), .B(x[2719]), .Z(n36474) );
  AND U20364 ( .A(n36467), .B(n36474), .Z(n54892) );
  NANDN U20365 ( .A(x[2717]), .B(y[2717]), .Z(n26825) );
  NANDN U20366 ( .A(x[2718]), .B(y[2718]), .Z(n26824) );
  NAND U20367 ( .A(n26825), .B(n26824), .Z(n54890) );
  NANDN U20368 ( .A(y[2716]), .B(x[2716]), .Z(n9963) );
  NANDN U20369 ( .A(y[2717]), .B(x[2717]), .Z(n36468) );
  AND U20370 ( .A(n9963), .B(n36468), .Z(n54888) );
  ANDN U20371 ( .B(y[2715]), .A(x[2715]), .Z(n54883) );
  XNOR U20372 ( .A(x[2716]), .B(y[2716]), .Z(n36461) );
  NANDN U20373 ( .A(y[2714]), .B(x[2714]), .Z(n9964) );
  NANDN U20374 ( .A(y[2715]), .B(x[2715]), .Z(n36462) );
  AND U20375 ( .A(n9964), .B(n36462), .Z(n54882) );
  XNOR U20376 ( .A(x[2714]), .B(y[2714]), .Z(n26827) );
  ANDN U20377 ( .B(y[2713]), .A(x[2713]), .Z(n26828) );
  ANDN U20378 ( .B(n26827), .A(n26828), .Z(n14318) );
  NANDN U20379 ( .A(x[2712]), .B(y[2712]), .Z(n26829) );
  ANDN U20380 ( .B(y[2711]), .A(x[2711]), .Z(n36450) );
  ANDN U20381 ( .B(n26829), .A(n36450), .Z(n54878) );
  NANDN U20382 ( .A(y[2710]), .B(x[2710]), .Z(n9965) );
  NANDN U20383 ( .A(y[2711]), .B(x[2711]), .Z(n26831) );
  NAND U20384 ( .A(n9965), .B(n26831), .Z(n54877) );
  NANDN U20385 ( .A(x[2709]), .B(y[2709]), .Z(n52024) );
  NANDN U20386 ( .A(x[2707]), .B(y[2707]), .Z(n36437) );
  ANDN U20387 ( .B(y[2708]), .A(x[2708]), .Z(n36444) );
  ANDN U20388 ( .B(n36437), .A(n36444), .Z(n54875) );
  ANDN U20389 ( .B(x[2706]), .A(y[2706]), .Z(n36435) );
  NANDN U20390 ( .A(y[2707]), .B(x[2707]), .Z(n26833) );
  NANDN U20391 ( .A(n36435), .B(n26833), .Z(n54874) );
  NANDN U20392 ( .A(x[2705]), .B(y[2705]), .Z(n26834) );
  NANDN U20393 ( .A(x[2706]), .B(y[2706]), .Z(n36438) );
  NAND U20394 ( .A(n26834), .B(n36438), .Z(n54873) );
  NANDN U20395 ( .A(y[2704]), .B(x[2704]), .Z(n26836) );
  ANDN U20396 ( .B(x[2705]), .A(y[2705]), .Z(n36432) );
  ANDN U20397 ( .B(n26836), .A(n36432), .Z(n54872) );
  NANDN U20398 ( .A(x[2703]), .B(y[2703]), .Z(n36425) );
  NANDN U20399 ( .A(x[2704]), .B(y[2704]), .Z(n26835) );
  NAND U20400 ( .A(n36425), .B(n26835), .Z(n54871) );
  NANDN U20401 ( .A(y[2702]), .B(x[2702]), .Z(n9966) );
  NANDN U20402 ( .A(y[2703]), .B(x[2703]), .Z(n26837) );
  AND U20403 ( .A(n9966), .B(n26837), .Z(n54870) );
  XNOR U20404 ( .A(x[2702]), .B(y[2702]), .Z(n26839) );
  NANDN U20405 ( .A(y[2698]), .B(x[2698]), .Z(n26842) );
  NANDN U20406 ( .A(y[2699]), .B(x[2699]), .Z(n26841) );
  NAND U20407 ( .A(n26842), .B(n26841), .Z(n54863) );
  NANDN U20408 ( .A(x[2697]), .B(y[2697]), .Z(n36408) );
  NANDN U20409 ( .A(x[2698]), .B(y[2698]), .Z(n36415) );
  NAND U20410 ( .A(n36408), .B(n36415), .Z(n54862) );
  NANDN U20411 ( .A(y[2696]), .B(x[2696]), .Z(n36404) );
  NANDN U20412 ( .A(y[2697]), .B(x[2697]), .Z(n26843) );
  AND U20413 ( .A(n36404), .B(n26843), .Z(n54861) );
  NANDN U20414 ( .A(x[2695]), .B(y[2695]), .Z(n26844) );
  NANDN U20415 ( .A(x[2696]), .B(y[2696]), .Z(n36409) );
  NAND U20416 ( .A(n26844), .B(n36409), .Z(n54860) );
  NANDN U20417 ( .A(y[2694]), .B(x[2694]), .Z(n26846) );
  NANDN U20418 ( .A(y[2695]), .B(x[2695]), .Z(n36405) );
  AND U20419 ( .A(n26846), .B(n36405), .Z(n54859) );
  NANDN U20420 ( .A(x[2693]), .B(y[2693]), .Z(n26848) );
  NANDN U20421 ( .A(x[2694]), .B(y[2694]), .Z(n26845) );
  NAND U20422 ( .A(n26848), .B(n26845), .Z(n54858) );
  NANDN U20423 ( .A(y[2692]), .B(x[2692]), .Z(n26851) );
  NANDN U20424 ( .A(y[2693]), .B(x[2693]), .Z(n26847) );
  NAND U20425 ( .A(n26851), .B(n26847), .Z(n54857) );
  NANDN U20426 ( .A(x[2691]), .B(y[2691]), .Z(n26852) );
  XNOR U20427 ( .A(x[2692]), .B(y[2692]), .Z(n9967) );
  AND U20428 ( .A(n26852), .B(n9967), .Z(n54856) );
  NANDN U20429 ( .A(y[2690]), .B(x[2690]), .Z(n26854) );
  NANDN U20430 ( .A(y[2691]), .B(x[2691]), .Z(n26850) );
  NAND U20431 ( .A(n26854), .B(n26850), .Z(n54855) );
  NANDN U20432 ( .A(x[2689]), .B(y[2689]), .Z(n36388) );
  NANDN U20433 ( .A(x[2690]), .B(y[2690]), .Z(n26853) );
  AND U20434 ( .A(n36388), .B(n26853), .Z(n54854) );
  NANDN U20435 ( .A(x[2687]), .B(y[2687]), .Z(n36382) );
  XNOR U20436 ( .A(x[2688]), .B(y[2688]), .Z(n9968) );
  AND U20437 ( .A(n36382), .B(n9968), .Z(n54852) );
  NANDN U20438 ( .A(y[2686]), .B(x[2686]), .Z(n26858) );
  NANDN U20439 ( .A(y[2687]), .B(x[2687]), .Z(n26857) );
  NAND U20440 ( .A(n26858), .B(n26857), .Z(n54851) );
  NANDN U20441 ( .A(x[2685]), .B(y[2685]), .Z(n36376) );
  NANDN U20442 ( .A(x[2686]), .B(y[2686]), .Z(n36383) );
  NAND U20443 ( .A(n36376), .B(n36383), .Z(n52025) );
  NANDN U20444 ( .A(y[2684]), .B(x[2684]), .Z(n26860) );
  NANDN U20445 ( .A(y[2685]), .B(x[2685]), .Z(n26859) );
  AND U20446 ( .A(n26860), .B(n26859), .Z(n52026) );
  NANDN U20447 ( .A(x[2681]), .B(y[2681]), .Z(n36364) );
  NANDN U20448 ( .A(x[2682]), .B(y[2682]), .Z(n36371) );
  NAND U20449 ( .A(n36364), .B(n36371), .Z(n54848) );
  NANDN U20450 ( .A(y[2680]), .B(x[2680]), .Z(n26864) );
  NANDN U20451 ( .A(y[2681]), .B(x[2681]), .Z(n26863) );
  NAND U20452 ( .A(n26864), .B(n26863), .Z(n54847) );
  NANDN U20453 ( .A(x[2679]), .B(y[2679]), .Z(n36358) );
  NANDN U20454 ( .A(x[2680]), .B(y[2680]), .Z(n36365) );
  AND U20455 ( .A(n36358), .B(n36365), .Z(n54846) );
  NANDN U20456 ( .A(y[2678]), .B(x[2678]), .Z(n26866) );
  NANDN U20457 ( .A(y[2679]), .B(x[2679]), .Z(n26865) );
  NAND U20458 ( .A(n26866), .B(n26865), .Z(n54845) );
  NANDN U20459 ( .A(x[2677]), .B(y[2677]), .Z(n36352) );
  NANDN U20460 ( .A(x[2678]), .B(y[2678]), .Z(n36359) );
  AND U20461 ( .A(n36352), .B(n36359), .Z(n54844) );
  NANDN U20462 ( .A(y[2676]), .B(x[2676]), .Z(n36349) );
  NANDN U20463 ( .A(y[2677]), .B(x[2677]), .Z(n26867) );
  NAND U20464 ( .A(n36349), .B(n26867), .Z(n54843) );
  NANDN U20465 ( .A(x[2675]), .B(y[2675]), .Z(n26868) );
  NANDN U20466 ( .A(x[2676]), .B(y[2676]), .Z(n36353) );
  NAND U20467 ( .A(n26868), .B(n36353), .Z(n54842) );
  NANDN U20468 ( .A(y[2674]), .B(x[2674]), .Z(n36343) );
  NANDN U20469 ( .A(y[2675]), .B(x[2675]), .Z(n36350) );
  AND U20470 ( .A(n36343), .B(n36350), .Z(n54841) );
  NANDN U20471 ( .A(x[2673]), .B(y[2673]), .Z(n26870) );
  NANDN U20472 ( .A(x[2674]), .B(y[2674]), .Z(n26869) );
  NAND U20473 ( .A(n26870), .B(n26869), .Z(n54840) );
  NANDN U20474 ( .A(y[2672]), .B(x[2672]), .Z(n9969) );
  NANDN U20475 ( .A(y[2673]), .B(x[2673]), .Z(n36344) );
  AND U20476 ( .A(n9969), .B(n36344), .Z(n54839) );
  XNOR U20477 ( .A(x[2672]), .B(y[2672]), .Z(n36337) );
  NANDN U20478 ( .A(y[2670]), .B(x[2670]), .Z(n36330) );
  NANDN U20479 ( .A(y[2671]), .B(x[2671]), .Z(n36338) );
  AND U20480 ( .A(n36330), .B(n36338), .Z(n52028) );
  ANDN U20481 ( .B(y[2670]), .A(x[2670]), .Z(n36335) );
  NANDN U20482 ( .A(x[2669]), .B(y[2669]), .Z(n26871) );
  NANDN U20483 ( .A(n36335), .B(n26871), .Z(n52029) );
  NANDN U20484 ( .A(y[2668]), .B(x[2668]), .Z(n9970) );
  NANDN U20485 ( .A(y[2669]), .B(x[2669]), .Z(n36332) );
  AND U20486 ( .A(n9970), .B(n36332), .Z(n54833) );
  ANDN U20487 ( .B(y[2667]), .A(x[2667]), .Z(n26872) );
  XNOR U20488 ( .A(x[2668]), .B(y[2668]), .Z(n36324) );
  NANDN U20489 ( .A(y[2666]), .B(x[2666]), .Z(n36317) );
  NANDN U20490 ( .A(y[2667]), .B(x[2667]), .Z(n36323) );
  NAND U20491 ( .A(n36317), .B(n36323), .Z(n52032) );
  NANDN U20492 ( .A(x[2665]), .B(y[2665]), .Z(n26874) );
  NANDN U20493 ( .A(x[2666]), .B(y[2666]), .Z(n26873) );
  AND U20494 ( .A(n26874), .B(n26873), .Z(n52033) );
  NANDN U20495 ( .A(y[2662]), .B(x[2662]), .Z(n9971) );
  NANDN U20496 ( .A(y[2663]), .B(x[2663]), .Z(n36312) );
  NAND U20497 ( .A(n9971), .B(n36312), .Z(n54831) );
  XNOR U20498 ( .A(y[2662]), .B(x[2662]), .Z(n36306) );
  NANDN U20499 ( .A(x[2661]), .B(y[2661]), .Z(n26878) );
  NAND U20500 ( .A(n36306), .B(n26878), .Z(n54830) );
  NANDN U20501 ( .A(y[2660]), .B(x[2660]), .Z(n36299) );
  NANDN U20502 ( .A(y[2661]), .B(x[2661]), .Z(n36305) );
  AND U20503 ( .A(n36299), .B(n36305), .Z(n52035) );
  NANDN U20504 ( .A(x[2657]), .B(y[2657]), .Z(n36289) );
  NANDN U20505 ( .A(x[2658]), .B(y[2658]), .Z(n26881) );
  NAND U20506 ( .A(n36289), .B(n26881), .Z(n54826) );
  NANDN U20507 ( .A(y[2656]), .B(x[2656]), .Z(n26882) );
  NANDN U20508 ( .A(y[2657]), .B(x[2657]), .Z(n36294) );
  NAND U20509 ( .A(n26882), .B(n36294), .Z(n54825) );
  NANDN U20510 ( .A(x[2655]), .B(y[2655]), .Z(n26884) );
  NANDN U20511 ( .A(x[2656]), .B(y[2656]), .Z(n36290) );
  AND U20512 ( .A(n26884), .B(n36290), .Z(n52037) );
  NANDN U20513 ( .A(y[2650]), .B(x[2650]), .Z(n9972) );
  NANDN U20514 ( .A(y[2651]), .B(x[2651]), .Z(n26891) );
  NAND U20515 ( .A(n9972), .B(n26891), .Z(n54822) );
  XNOR U20516 ( .A(y[2650]), .B(x[2650]), .Z(n36274) );
  NANDN U20517 ( .A(x[2649]), .B(y[2649]), .Z(n26894) );
  NAND U20518 ( .A(n36274), .B(n26894), .Z(n52040) );
  NANDN U20519 ( .A(y[2648]), .B(x[2648]), .Z(n26896) );
  NANDN U20520 ( .A(y[2649]), .B(x[2649]), .Z(n36273) );
  AND U20521 ( .A(n26896), .B(n36273), .Z(n54820) );
  XNOR U20522 ( .A(y[2646]), .B(x[2646]), .Z(n26899) );
  NANDN U20523 ( .A(x[2645]), .B(y[2645]), .Z(n36260) );
  NAND U20524 ( .A(n26899), .B(n36260), .Z(n54816) );
  NANDN U20525 ( .A(y[2644]), .B(x[2644]), .Z(n9973) );
  NANDN U20526 ( .A(y[2645]), .B(x[2645]), .Z(n26898) );
  NAND U20527 ( .A(n9973), .B(n26898), .Z(n52042) );
  XNOR U20528 ( .A(y[2644]), .B(x[2644]), .Z(n26901) );
  NANDN U20529 ( .A(x[2643]), .B(y[2643]), .Z(n36254) );
  AND U20530 ( .A(n26901), .B(n36254), .Z(n54815) );
  NANDN U20531 ( .A(y[2640]), .B(x[2640]), .Z(n36246) );
  NANDN U20532 ( .A(y[2641]), .B(x[2641]), .Z(n26903) );
  NAND U20533 ( .A(n36246), .B(n26903), .Z(n54813) );
  ANDN U20534 ( .B(y[2639]), .A(x[2639]), .Z(n36242) );
  NANDN U20535 ( .A(x[2640]), .B(y[2640]), .Z(n26905) );
  NANDN U20536 ( .A(n36242), .B(n26905), .Z(n52044) );
  NANDN U20537 ( .A(y[2638]), .B(x[2638]), .Z(n9974) );
  NANDN U20538 ( .A(y[2639]), .B(x[2639]), .Z(n36247) );
  AND U20539 ( .A(n9974), .B(n36247), .Z(n54812) );
  NANDN U20540 ( .A(x[2635]), .B(y[2635]), .Z(n26910) );
  NANDN U20541 ( .A(x[2636]), .B(y[2636]), .Z(n26907) );
  NAND U20542 ( .A(n26910), .B(n26907), .Z(n54809) );
  ANDN U20543 ( .B(x[2634]), .A(y[2634]), .Z(n36227) );
  NANDN U20544 ( .A(y[2635]), .B(x[2635]), .Z(n26909) );
  NANDN U20545 ( .A(n36227), .B(n26909), .Z(n52046) );
  NANDN U20546 ( .A(x[2633]), .B(y[2633]), .Z(n36225) );
  NANDN U20547 ( .A(x[2634]), .B(y[2634]), .Z(n26911) );
  AND U20548 ( .A(n36225), .B(n26911), .Z(n54808) );
  NANDN U20549 ( .A(x[2631]), .B(y[2631]), .Z(n54806) );
  XOR U20550 ( .A(x[2632]), .B(y[2632]), .Z(n36221) );
  ANDN U20551 ( .B(n54806), .A(n36221), .Z(n14228) );
  ANDN U20552 ( .B(x[2631]), .A(y[2631]), .Z(n36223) );
  NANDN U20553 ( .A(y[2630]), .B(x[2630]), .Z(n9975) );
  NANDN U20554 ( .A(n36223), .B(n9975), .Z(n54805) );
  XNOR U20555 ( .A(y[2630]), .B(x[2630]), .Z(n14224) );
  NANDN U20556 ( .A(y[2628]), .B(x[2628]), .Z(n26914) );
  ANDN U20557 ( .B(x[2629]), .A(y[2629]), .Z(n26913) );
  ANDN U20558 ( .B(n26914), .A(n26913), .Z(n54804) );
  ANDN U20559 ( .B(y[2627]), .A(x[2627]), .Z(n36208) );
  ANDN U20560 ( .B(y[2628]), .A(x[2628]), .Z(n36214) );
  OR U20561 ( .A(n36208), .B(n36214), .Z(n54803) );
  NANDN U20562 ( .A(y[2626]), .B(x[2626]), .Z(n36204) );
  NANDN U20563 ( .A(y[2627]), .B(x[2627]), .Z(n26915) );
  AND U20564 ( .A(n36204), .B(n26915), .Z(n54802) );
  ANDN U20565 ( .B(y[2626]), .A(x[2626]), .Z(n36209) );
  NANDN U20566 ( .A(x[2625]), .B(y[2625]), .Z(n26916) );
  NANDN U20567 ( .A(n36209), .B(n26916), .Z(n54801) );
  NANDN U20568 ( .A(y[2624]), .B(x[2624]), .Z(n26918) );
  NANDN U20569 ( .A(y[2625]), .B(x[2625]), .Z(n36203) );
  AND U20570 ( .A(n26918), .B(n36203), .Z(n54800) );
  NANDN U20571 ( .A(x[2623]), .B(y[2623]), .Z(n26920) );
  NANDN U20572 ( .A(x[2624]), .B(y[2624]), .Z(n26917) );
  NAND U20573 ( .A(n26920), .B(n26917), .Z(n54799) );
  NANDN U20574 ( .A(y[2622]), .B(x[2622]), .Z(n26923) );
  NANDN U20575 ( .A(y[2623]), .B(x[2623]), .Z(n26919) );
  NAND U20576 ( .A(n26923), .B(n26919), .Z(n54798) );
  NANDN U20577 ( .A(x[2622]), .B(y[2622]), .Z(n26921) );
  ANDN U20578 ( .B(y[2621]), .A(x[2621]), .Z(n36193) );
  ANDN U20579 ( .B(n26921), .A(n36193), .Z(n54796) );
  NANDN U20580 ( .A(y[2620]), .B(x[2620]), .Z(n9976) );
  NANDN U20581 ( .A(y[2621]), .B(x[2621]), .Z(n26922) );
  NAND U20582 ( .A(n9976), .B(n26922), .Z(n54795) );
  XNOR U20583 ( .A(y[2620]), .B(x[2620]), .Z(n26925) );
  ANDN U20584 ( .B(y[2619]), .A(x[2619]), .Z(n36187) );
  ANDN U20585 ( .B(n26925), .A(n36187), .Z(n54794) );
  NANDN U20586 ( .A(y[2618]), .B(x[2618]), .Z(n9977) );
  NANDN U20587 ( .A(y[2619]), .B(x[2619]), .Z(n26924) );
  NAND U20588 ( .A(n9977), .B(n26924), .Z(n54793) );
  XNOR U20589 ( .A(x[2618]), .B(y[2618]), .Z(n36183) );
  NANDN U20590 ( .A(y[2616]), .B(x[2616]), .Z(n9978) );
  NANDN U20591 ( .A(y[2617]), .B(x[2617]), .Z(n36185) );
  NAND U20592 ( .A(n9978), .B(n36185), .Z(n54791) );
  NANDN U20593 ( .A(x[2613]), .B(y[2613]), .Z(n26926) );
  XOR U20594 ( .A(y[2614]), .B(x[2614]), .Z(n36170) );
  ANDN U20595 ( .B(n26926), .A(n36170), .Z(n54787) );
  ANDN U20596 ( .B(x[2613]), .A(y[2613]), .Z(n36172) );
  NANDN U20597 ( .A(y[2612]), .B(x[2612]), .Z(n36163) );
  NANDN U20598 ( .A(n36172), .B(n36163), .Z(n52051) );
  NANDN U20599 ( .A(y[2610]), .B(x[2610]), .Z(n36157) );
  NANDN U20600 ( .A(y[2611]), .B(x[2611]), .Z(n36164) );
  AND U20601 ( .A(n36157), .B(n36164), .Z(n54785) );
  NANDN U20602 ( .A(x[2609]), .B(y[2609]), .Z(n26930) );
  XNOR U20603 ( .A(x[2610]), .B(y[2610]), .Z(n9979) );
  NAND U20604 ( .A(n26930), .B(n9979), .Z(n54784) );
  NANDN U20605 ( .A(y[2608]), .B(x[2608]), .Z(n9980) );
  NANDN U20606 ( .A(y[2609]), .B(x[2609]), .Z(n36158) );
  AND U20607 ( .A(n9980), .B(n36158), .Z(n54782) );
  XNOR U20608 ( .A(y[2608]), .B(x[2608]), .Z(n36152) );
  NANDN U20609 ( .A(x[2607]), .B(y[2607]), .Z(n36148) );
  NAND U20610 ( .A(n36152), .B(n36148), .Z(n54781) );
  ANDN U20611 ( .B(x[2606]), .A(y[2606]), .Z(n36146) );
  ANDN U20612 ( .B(x[2607]), .A(y[2607]), .Z(n36153) );
  NOR U20613 ( .A(n36146), .B(n36153), .Z(n54780) );
  NANDN U20614 ( .A(x[2605]), .B(y[2605]), .Z(n26932) );
  XNOR U20615 ( .A(y[2606]), .B(x[2606]), .Z(n9981) );
  NAND U20616 ( .A(n26932), .B(n9981), .Z(n54779) );
  ANDN U20617 ( .B(x[2605]), .A(y[2605]), .Z(n36143) );
  NANDN U20618 ( .A(y[2604]), .B(x[2604]), .Z(n36137) );
  NANDN U20619 ( .A(n36143), .B(n36137), .Z(n54778) );
  NANDN U20620 ( .A(x[2603]), .B(y[2603]), .Z(n26934) );
  NANDN U20621 ( .A(x[2604]), .B(y[2604]), .Z(n26933) );
  AND U20622 ( .A(n26934), .B(n26933), .Z(n54777) );
  NANDN U20623 ( .A(y[2602]), .B(x[2602]), .Z(n36131) );
  NANDN U20624 ( .A(y[2603]), .B(x[2603]), .Z(n36138) );
  NAND U20625 ( .A(n36131), .B(n36138), .Z(n54776) );
  NANDN U20626 ( .A(x[2601]), .B(y[2601]), .Z(n26936) );
  NANDN U20627 ( .A(x[2602]), .B(y[2602]), .Z(n26935) );
  AND U20628 ( .A(n26936), .B(n26935), .Z(n54775) );
  NANDN U20629 ( .A(y[2600]), .B(x[2600]), .Z(n36125) );
  NANDN U20630 ( .A(y[2601]), .B(x[2601]), .Z(n36132) );
  NAND U20631 ( .A(n36125), .B(n36132), .Z(n54774) );
  NANDN U20632 ( .A(x[2599]), .B(y[2599]), .Z(n26938) );
  NANDN U20633 ( .A(x[2600]), .B(y[2600]), .Z(n26937) );
  NAND U20634 ( .A(n26938), .B(n26937), .Z(n54773) );
  NANDN U20635 ( .A(y[2598]), .B(x[2598]), .Z(n36119) );
  NANDN U20636 ( .A(y[2599]), .B(x[2599]), .Z(n36126) );
  AND U20637 ( .A(n36119), .B(n36126), .Z(n54772) );
  NANDN U20638 ( .A(x[2597]), .B(y[2597]), .Z(n36118) );
  NANDN U20639 ( .A(x[2598]), .B(y[2598]), .Z(n26939) );
  NAND U20640 ( .A(n36118), .B(n26939), .Z(n54771) );
  NANDN U20641 ( .A(y[2596]), .B(x[2596]), .Z(n9982) );
  NANDN U20642 ( .A(y[2597]), .B(x[2597]), .Z(n36120) );
  AND U20643 ( .A(n9982), .B(n36120), .Z(n54770) );
  NANDN U20644 ( .A(y[2594]), .B(x[2594]), .Z(n9983) );
  ANDN U20645 ( .B(x[2595]), .A(y[2595]), .Z(n36112) );
  ANDN U20646 ( .B(n9983), .A(n36112), .Z(n54768) );
  XOR U20647 ( .A(y[2594]), .B(x[2594]), .Z(n36108) );
  NANDN U20648 ( .A(x[2593]), .B(y[2593]), .Z(n36102) );
  NANDN U20649 ( .A(n36108), .B(n36102), .Z(n52052) );
  XNOR U20650 ( .A(y[2592]), .B(x[2592]), .Z(n26943) );
  ANDN U20651 ( .B(y[2591]), .A(x[2591]), .Z(n26945) );
  ANDN U20652 ( .B(n26943), .A(n26945), .Z(n54766) );
  ANDN U20653 ( .B(x[2588]), .A(y[2588]), .Z(n36088) );
  ANDN U20654 ( .B(x[2589]), .A(y[2589]), .Z(n36094) );
  OR U20655 ( .A(n36088), .B(n36094), .Z(n52054) );
  NANDN U20656 ( .A(y[2586]), .B(x[2586]), .Z(n9984) );
  ANDN U20657 ( .B(x[2587]), .A(y[2587]), .Z(n36089) );
  ANDN U20658 ( .B(n9984), .A(n36089), .Z(n54762) );
  XOR U20659 ( .A(y[2586]), .B(x[2586]), .Z(n36077) );
  NANDN U20660 ( .A(x[2585]), .B(y[2585]), .Z(n9985) );
  NANDN U20661 ( .A(n36077), .B(n9985), .Z(n54761) );
  ANDN U20662 ( .B(x[2584]), .A(y[2584]), .Z(n36072) );
  NANDN U20663 ( .A(y[2585]), .B(x[2585]), .Z(n9986) );
  NANDN U20664 ( .A(n36072), .B(n9986), .Z(n54760) );
  NANDN U20665 ( .A(x[2583]), .B(y[2583]), .Z(n36068) );
  NANDN U20666 ( .A(x[2584]), .B(y[2584]), .Z(n36076) );
  AND U20667 ( .A(n36068), .B(n36076), .Z(n54759) );
  ANDN U20668 ( .B(x[2582]), .A(y[2582]), .Z(n36067) );
  ANDN U20669 ( .B(x[2583]), .A(y[2583]), .Z(n36074) );
  OR U20670 ( .A(n36067), .B(n36074), .Z(n54758) );
  NANDN U20671 ( .A(x[2581]), .B(y[2581]), .Z(n26949) );
  NANDN U20672 ( .A(x[2582]), .B(y[2582]), .Z(n54757) );
  AND U20673 ( .A(n26949), .B(n54757), .Z(n14167) );
  NANDN U20674 ( .A(y[2580]), .B(x[2580]), .Z(n26950) );
  ANDN U20675 ( .B(y[2579]), .A(x[2579]), .Z(n26952) );
  NANDN U20676 ( .A(x[2578]), .B(y[2578]), .Z(n26953) );
  NANDN U20677 ( .A(x[2577]), .B(y[2577]), .Z(n26958) );
  AND U20678 ( .A(n26953), .B(n26958), .Z(n14159) );
  ANDN U20679 ( .B(x[2576]), .A(y[2576]), .Z(n54750) );
  NANDN U20680 ( .A(x[2576]), .B(y[2576]), .Z(n26957) );
  NANDN U20681 ( .A(y[2574]), .B(x[2574]), .Z(n36050) );
  NANDN U20682 ( .A(y[2575]), .B(x[2575]), .Z(n36057) );
  NAND U20683 ( .A(n36050), .B(n36057), .Z(n54747) );
  NANDN U20684 ( .A(x[2573]), .B(y[2573]), .Z(n26960) );
  XNOR U20685 ( .A(x[2574]), .B(y[2574]), .Z(n9987) );
  AND U20686 ( .A(n26960), .B(n9987), .Z(n54746) );
  NANDN U20687 ( .A(y[2572]), .B(x[2572]), .Z(n26961) );
  NANDN U20688 ( .A(y[2573]), .B(x[2573]), .Z(n36049) );
  NAND U20689 ( .A(n26961), .B(n36049), .Z(n54745) );
  ANDN U20690 ( .B(x[2570]), .A(y[2570]), .Z(n36040) );
  NANDN U20691 ( .A(y[2571]), .B(x[2571]), .Z(n26962) );
  NANDN U20692 ( .A(n36040), .B(n26962), .Z(n52056) );
  NANDN U20693 ( .A(x[2569]), .B(y[2569]), .Z(n26965) );
  NANDN U20694 ( .A(x[2570]), .B(y[2570]), .Z(n26963) );
  NAND U20695 ( .A(n26965), .B(n26963), .Z(n54744) );
  ANDN U20696 ( .B(x[2568]), .A(y[2568]), .Z(n36034) );
  ANDN U20697 ( .B(x[2569]), .A(y[2569]), .Z(n36041) );
  NOR U20698 ( .A(n36034), .B(n36041), .Z(n54743) );
  NANDN U20699 ( .A(x[2567]), .B(y[2567]), .Z(n36030) );
  NANDN U20700 ( .A(x[2568]), .B(y[2568]), .Z(n26966) );
  NAND U20701 ( .A(n36030), .B(n26966), .Z(n54742) );
  NANDN U20702 ( .A(y[2566]), .B(x[2566]), .Z(n26967) );
  ANDN U20703 ( .B(x[2567]), .A(y[2567]), .Z(n36035) );
  ANDN U20704 ( .B(n26967), .A(n36035), .Z(n54741) );
  NANDN U20705 ( .A(x[2566]), .B(y[2566]), .Z(n54740) );
  NANDN U20706 ( .A(y[2565]), .B(x[2565]), .Z(n54739) );
  ANDN U20707 ( .B(x[2564]), .A(y[2564]), .Z(n54737) );
  ANDN U20708 ( .B(n54739), .A(n54737), .Z(n14142) );
  NANDN U20709 ( .A(x[2564]), .B(y[2564]), .Z(n26969) );
  ANDN U20710 ( .B(x[2562]), .A(y[2562]), .Z(n36017) );
  ANDN U20711 ( .B(x[2563]), .A(y[2563]), .Z(n36025) );
  NOR U20712 ( .A(n36017), .B(n36025), .Z(n54736) );
  ANDN U20713 ( .B(x[2560]), .A(y[2560]), .Z(n36011) );
  ANDN U20714 ( .B(x[2561]), .A(y[2561]), .Z(n36020) );
  NOR U20715 ( .A(n36011), .B(n36020), .Z(n54734) );
  NANDN U20716 ( .A(x[2559]), .B(y[2559]), .Z(n26970) );
  NANDN U20717 ( .A(x[2560]), .B(y[2560]), .Z(n36015) );
  NAND U20718 ( .A(n26970), .B(n36015), .Z(n54732) );
  ANDN U20719 ( .B(x[2556]), .A(y[2556]), .Z(n54727) );
  XNOR U20720 ( .A(y[2556]), .B(x[2556]), .Z(n36000) );
  NANDN U20721 ( .A(x[2555]), .B(y[2555]), .Z(n35996) );
  AND U20722 ( .A(n36000), .B(n35996), .Z(n54726) );
  ANDN U20723 ( .B(x[2555]), .A(y[2555]), .Z(n36001) );
  NANDN U20724 ( .A(y[2554]), .B(x[2554]), .Z(n9988) );
  NANDN U20725 ( .A(n36001), .B(n9988), .Z(n54725) );
  NANDN U20726 ( .A(x[2553]), .B(y[2553]), .Z(n26972) );
  XOR U20727 ( .A(y[2554]), .B(x[2554]), .Z(n35992) );
  ANDN U20728 ( .B(n26972), .A(n35992), .Z(n54724) );
  ANDN U20729 ( .B(x[2553]), .A(y[2553]), .Z(n35994) );
  NANDN U20730 ( .A(y[2552]), .B(x[2552]), .Z(n9989) );
  NANDN U20731 ( .A(n35994), .B(n9989), .Z(n54723) );
  XNOR U20732 ( .A(y[2552]), .B(x[2552]), .Z(n26975) );
  NANDN U20733 ( .A(x[2551]), .B(y[2551]), .Z(n35984) );
  AND U20734 ( .A(n26975), .B(n35984), .Z(n54722) );
  NANDN U20735 ( .A(y[2550]), .B(x[2550]), .Z(n9990) );
  NANDN U20736 ( .A(y[2551]), .B(x[2551]), .Z(n26974) );
  NAND U20737 ( .A(n9990), .B(n26974), .Z(n54721) );
  NANDN U20738 ( .A(y[2548]), .B(x[2548]), .Z(n9991) );
  ANDN U20739 ( .B(x[2549]), .A(y[2549]), .Z(n35980) );
  ANDN U20740 ( .B(n9991), .A(n35980), .Z(n54719) );
  XNOR U20741 ( .A(y[2548]), .B(x[2548]), .Z(n35974) );
  NANDN U20742 ( .A(x[2547]), .B(y[2547]), .Z(n35970) );
  NAND U20743 ( .A(n35974), .B(n35970), .Z(n54718) );
  NANDN U20744 ( .A(y[2546]), .B(x[2546]), .Z(n9992) );
  NANDN U20745 ( .A(y[2547]), .B(x[2547]), .Z(n35973) );
  NAND U20746 ( .A(n9992), .B(n35973), .Z(n54717) );
  NANDN U20747 ( .A(x[2545]), .B(y[2545]), .Z(n35962) );
  XOR U20748 ( .A(y[2546]), .B(x[2546]), .Z(n35966) );
  ANDN U20749 ( .B(n35962), .A(n35966), .Z(n54716) );
  NANDN U20750 ( .A(x[2544]), .B(y[2544]), .Z(n35964) );
  ANDN U20751 ( .B(y[2543]), .A(x[2543]), .Z(n35956) );
  ANDN U20752 ( .B(n35964), .A(n35956), .Z(n54714) );
  ANDN U20753 ( .B(x[2543]), .A(y[2543]), .Z(n26976) );
  NANDN U20754 ( .A(y[2542]), .B(x[2542]), .Z(n26978) );
  NANDN U20755 ( .A(n26976), .B(n26978), .Z(n54713) );
  ANDN U20756 ( .B(y[2541]), .A(x[2541]), .Z(n35950) );
  XNOR U20757 ( .A(y[2542]), .B(x[2542]), .Z(n9993) );
  NANDN U20758 ( .A(n35950), .B(n9993), .Z(n52060) );
  NANDN U20759 ( .A(y[2540]), .B(x[2540]), .Z(n35946) );
  NANDN U20760 ( .A(y[2541]), .B(x[2541]), .Z(n26979) );
  AND U20761 ( .A(n35946), .B(n26979), .Z(n54712) );
  XNOR U20762 ( .A(x[2538]), .B(y[2538]), .Z(n52063) );
  NANDN U20763 ( .A(x[2536]), .B(y[2536]), .Z(n26984) );
  NANDN U20764 ( .A(x[2535]), .B(y[2535]), .Z(n54707) );
  AND U20765 ( .A(n26984), .B(n54707), .Z(n14104) );
  NANDN U20766 ( .A(y[2535]), .B(x[2535]), .Z(n26986) );
  ANDN U20767 ( .B(x[2534]), .A(y[2534]), .Z(n35933) );
  ANDN U20768 ( .B(n26986), .A(n35933), .Z(n54706) );
  NANDN U20769 ( .A(x[2533]), .B(y[2533]), .Z(n26988) );
  NANDN U20770 ( .A(x[2534]), .B(y[2534]), .Z(n26987) );
  NAND U20771 ( .A(n26988), .B(n26987), .Z(n54705) );
  ANDN U20772 ( .B(x[2532]), .A(y[2532]), .Z(n35927) );
  ANDN U20773 ( .B(x[2533]), .A(y[2533]), .Z(n35934) );
  OR U20774 ( .A(n35927), .B(n35934), .Z(n52064) );
  NANDN U20775 ( .A(x[2531]), .B(y[2531]), .Z(n35923) );
  NANDN U20776 ( .A(x[2532]), .B(y[2532]), .Z(n26989) );
  AND U20777 ( .A(n35923), .B(n26989), .Z(n54704) );
  NANDN U20778 ( .A(x[2529]), .B(y[2529]), .Z(n26992) );
  NANDN U20779 ( .A(x[2530]), .B(y[2530]), .Z(n54702) );
  AND U20780 ( .A(n26992), .B(n54702), .Z(n14097) );
  ANDN U20781 ( .B(x[2529]), .A(y[2529]), .Z(n26990) );
  NANDN U20782 ( .A(x[2528]), .B(y[2528]), .Z(n26993) );
  ANDN U20783 ( .B(x[2526]), .A(y[2526]), .Z(n35910) );
  ANDN U20784 ( .B(x[2527]), .A(y[2527]), .Z(n35918) );
  OR U20785 ( .A(n35910), .B(n35918), .Z(n52068) );
  NANDN U20786 ( .A(x[2525]), .B(y[2525]), .Z(n35907) );
  NANDN U20787 ( .A(x[2526]), .B(y[2526]), .Z(n35914) );
  AND U20788 ( .A(n35907), .B(n35914), .Z(n54699) );
  ANDN U20789 ( .B(x[2523]), .A(y[2523]), .Z(n35905) );
  NANDN U20790 ( .A(y[2522]), .B(x[2522]), .Z(n26994) );
  NANDN U20791 ( .A(n35905), .B(n26994), .Z(n54696) );
  NANDN U20792 ( .A(x[2521]), .B(y[2521]), .Z(n35893) );
  NANDN U20793 ( .A(x[2522]), .B(y[2522]), .Z(n35898) );
  AND U20794 ( .A(n35893), .B(n35898), .Z(n52069) );
  NANDN U20795 ( .A(y[2520]), .B(x[2520]), .Z(n9994) );
  NANDN U20796 ( .A(y[2521]), .B(x[2521]), .Z(n26995) );
  NAND U20797 ( .A(n9994), .B(n26995), .Z(n54695) );
  XOR U20798 ( .A(y[2520]), .B(x[2520]), .Z(n26996) );
  ANDN U20799 ( .B(y[2519]), .A(x[2519]), .Z(n35888) );
  NOR U20800 ( .A(n26996), .B(n35888), .Z(n54694) );
  ANDN U20801 ( .B(x[2519]), .A(y[2519]), .Z(n26997) );
  NANDN U20802 ( .A(y[2518]), .B(x[2518]), .Z(n35884) );
  NANDN U20803 ( .A(n26997), .B(n35884), .Z(n54693) );
  NANDN U20804 ( .A(y[2514]), .B(x[2514]), .Z(n27005) );
  NANDN U20805 ( .A(x[2514]), .B(y[2514]), .Z(n35880) );
  NANDN U20806 ( .A(x[2513]), .B(y[2513]), .Z(n27008) );
  AND U20807 ( .A(n35880), .B(n27008), .Z(n14074) );
  NANDN U20808 ( .A(y[2512]), .B(x[2512]), .Z(n54684) );
  ANDN U20809 ( .B(y[2511]), .A(x[2511]), .Z(n54683) );
  NANDN U20810 ( .A(y[2511]), .B(x[2511]), .Z(n27009) );
  ANDN U20811 ( .B(x[2510]), .A(y[2510]), .Z(n35870) );
  ANDN U20812 ( .B(n27009), .A(n35870), .Z(n54682) );
  NANDN U20813 ( .A(x[2509]), .B(y[2509]), .Z(n27011) );
  XNOR U20814 ( .A(x[2510]), .B(y[2510]), .Z(n9995) );
  NAND U20815 ( .A(n27011), .B(n9995), .Z(n54681) );
  ANDN U20816 ( .B(x[2508]), .A(y[2508]), .Z(n35864) );
  ANDN U20817 ( .B(x[2509]), .A(y[2509]), .Z(n35871) );
  NOR U20818 ( .A(n35864), .B(n35871), .Z(n54680) );
  NANDN U20819 ( .A(x[2507]), .B(y[2507]), .Z(n35860) );
  XNOR U20820 ( .A(x[2508]), .B(y[2508]), .Z(n9996) );
  NAND U20821 ( .A(n35860), .B(n9996), .Z(n54679) );
  ANDN U20822 ( .B(x[2506]), .A(y[2506]), .Z(n27014) );
  ANDN U20823 ( .B(x[2507]), .A(y[2507]), .Z(n35865) );
  NOR U20824 ( .A(n27014), .B(n35865), .Z(n54678) );
  ANDN U20825 ( .B(y[2505]), .A(x[2505]), .Z(n35854) );
  NANDN U20826 ( .A(x[2506]), .B(y[2506]), .Z(n35859) );
  NANDN U20827 ( .A(n35854), .B(n35859), .Z(n54677) );
  XNOR U20828 ( .A(y[2504]), .B(x[2504]), .Z(n9997) );
  ANDN U20829 ( .B(y[2503]), .A(x[2503]), .Z(n35848) );
  ANDN U20830 ( .B(n9997), .A(n35848), .Z(n54675) );
  NANDN U20831 ( .A(y[2502]), .B(x[2502]), .Z(n27017) );
  NANDN U20832 ( .A(y[2503]), .B(x[2503]), .Z(n27016) );
  NAND U20833 ( .A(n27017), .B(n27016), .Z(n54674) );
  NANDN U20834 ( .A(x[2501]), .B(y[2501]), .Z(n35842) );
  XNOR U20835 ( .A(x[2502]), .B(y[2502]), .Z(n9998) );
  AND U20836 ( .A(n35842), .B(n9998), .Z(n54673) );
  NANDN U20837 ( .A(y[2500]), .B(x[2500]), .Z(n9999) );
  NANDN U20838 ( .A(y[2501]), .B(x[2501]), .Z(n27018) );
  NAND U20839 ( .A(n9999), .B(n27018), .Z(n54672) );
  XNOR U20840 ( .A(y[2500]), .B(x[2500]), .Z(n35838) );
  NANDN U20841 ( .A(x[2499]), .B(y[2499]), .Z(n27019) );
  AND U20842 ( .A(n35838), .B(n27019), .Z(n54671) );
  NANDN U20843 ( .A(y[2498]), .B(x[2498]), .Z(n10000) );
  NANDN U20844 ( .A(y[2499]), .B(x[2499]), .Z(n35837) );
  NAND U20845 ( .A(n10000), .B(n35837), .Z(n54669) );
  ANDN U20846 ( .B(y[2497]), .A(x[2497]), .Z(n27020) );
  NANDN U20847 ( .A(y[2496]), .B(x[2496]), .Z(n10001) );
  NANDN U20848 ( .A(y[2497]), .B(x[2497]), .Z(n35831) );
  AND U20849 ( .A(n10001), .B(n35831), .Z(n54668) );
  XNOR U20850 ( .A(y[2496]), .B(x[2496]), .Z(n35826) );
  NANDN U20851 ( .A(x[2495]), .B(y[2495]), .Z(n35822) );
  NAND U20852 ( .A(n35826), .B(n35822), .Z(n54667) );
  NANDN U20853 ( .A(y[2494]), .B(x[2494]), .Z(n10002) );
  ANDN U20854 ( .B(x[2495]), .A(y[2495]), .Z(n35827) );
  ANDN U20855 ( .B(n10002), .A(n35827), .Z(n54666) );
  XOR U20856 ( .A(y[2494]), .B(x[2494]), .Z(n35818) );
  NANDN U20857 ( .A(x[2493]), .B(y[2493]), .Z(n27023) );
  NANDN U20858 ( .A(n35818), .B(n27023), .Z(n54665) );
  ANDN U20859 ( .B(x[2493]), .A(y[2493]), .Z(n35820) );
  NANDN U20860 ( .A(y[2492]), .B(x[2492]), .Z(n35812) );
  NANDN U20861 ( .A(n35820), .B(n35812), .Z(n54664) );
  NANDN U20862 ( .A(x[2492]), .B(y[2492]), .Z(n27022) );
  ANDN U20863 ( .B(y[2491]), .A(x[2491]), .Z(n35808) );
  ANDN U20864 ( .B(n27022), .A(n35808), .Z(n54663) );
  ANDN U20865 ( .B(x[2491]), .A(y[2491]), .Z(n35814) );
  NANDN U20866 ( .A(y[2490]), .B(x[2490]), .Z(n27024) );
  NANDN U20867 ( .A(n35814), .B(n27024), .Z(n54662) );
  ANDN U20868 ( .B(y[2489]), .A(x[2489]), .Z(n35802) );
  ANDN U20869 ( .B(y[2490]), .A(x[2490]), .Z(n35810) );
  NOR U20870 ( .A(n35802), .B(n35810), .Z(n54661) );
  NANDN U20871 ( .A(y[2488]), .B(x[2488]), .Z(n35798) );
  NANDN U20872 ( .A(y[2489]), .B(x[2489]), .Z(n27025) );
  NAND U20873 ( .A(n35798), .B(n27025), .Z(n54660) );
  NANDN U20874 ( .A(x[2487]), .B(y[2487]), .Z(n27027) );
  XNOR U20875 ( .A(x[2488]), .B(y[2488]), .Z(n10003) );
  NAND U20876 ( .A(n27027), .B(n10003), .Z(n54659) );
  NANDN U20877 ( .A(y[2486]), .B(x[2486]), .Z(n27028) );
  NANDN U20878 ( .A(y[2487]), .B(x[2487]), .Z(n35797) );
  AND U20879 ( .A(n27028), .B(n35797), .Z(n52072) );
  ANDN U20880 ( .B(y[2483]), .A(x[2483]), .Z(n27033) );
  XNOR U20881 ( .A(y[2484]), .B(x[2484]), .Z(n27031) );
  NANDN U20882 ( .A(n27033), .B(n27031), .Z(n52075) );
  ANDN U20883 ( .B(x[2482]), .A(y[2482]), .Z(n35782) );
  NANDN U20884 ( .A(y[2483]), .B(x[2483]), .Z(n27030) );
  NANDN U20885 ( .A(n35782), .B(n27030), .Z(n54656) );
  NANDN U20886 ( .A(x[2481]), .B(y[2481]), .Z(n27034) );
  ANDN U20887 ( .B(y[2482]), .A(x[2482]), .Z(n27032) );
  ANDN U20888 ( .B(n27034), .A(n27032), .Z(n54655) );
  ANDN U20889 ( .B(x[2480]), .A(y[2480]), .Z(n35776) );
  ANDN U20890 ( .B(x[2481]), .A(y[2481]), .Z(n35783) );
  OR U20891 ( .A(n35776), .B(n35783), .Z(n54654) );
  NANDN U20892 ( .A(x[2479]), .B(y[2479]), .Z(n35772) );
  NANDN U20893 ( .A(x[2480]), .B(y[2480]), .Z(n27035) );
  AND U20894 ( .A(n35772), .B(n27035), .Z(n54653) );
  ANDN U20895 ( .B(x[2479]), .A(y[2479]), .Z(n35777) );
  NANDN U20896 ( .A(y[2478]), .B(x[2478]), .Z(n27036) );
  NANDN U20897 ( .A(n35777), .B(n27036), .Z(n54652) );
  NANDN U20898 ( .A(x[2476]), .B(y[2476]), .Z(n54649) );
  NANDN U20899 ( .A(x[2477]), .B(y[2477]), .Z(n52077) );
  AND U20900 ( .A(n54649), .B(n52077), .Z(n35768) );
  NANDN U20901 ( .A(y[2476]), .B(x[2476]), .Z(n27037) );
  NANDN U20902 ( .A(x[2475]), .B(y[2475]), .Z(n54650) );
  ANDN U20903 ( .B(x[2475]), .A(y[2475]), .Z(n35765) );
  NANDN U20904 ( .A(y[2474]), .B(x[2474]), .Z(n10004) );
  NANDN U20905 ( .A(n35765), .B(n10004), .Z(n54648) );
  XNOR U20906 ( .A(y[2474]), .B(x[2474]), .Z(n27038) );
  NANDN U20907 ( .A(x[2473]), .B(y[2473]), .Z(n27040) );
  AND U20908 ( .A(n27038), .B(n27040), .Z(n54647) );
  NANDN U20909 ( .A(y[2472]), .B(x[2472]), .Z(n35753) );
  NANDN U20910 ( .A(y[2473]), .B(x[2473]), .Z(n27039) );
  NAND U20911 ( .A(n35753), .B(n27039), .Z(n54646) );
  NANDN U20912 ( .A(x[2471]), .B(y[2471]), .Z(n35750) );
  NANDN U20913 ( .A(x[2472]), .B(y[2472]), .Z(n27041) );
  AND U20914 ( .A(n35750), .B(n27041), .Z(n54645) );
  NANDN U20915 ( .A(y[2470]), .B(x[2470]), .Z(n10005) );
  NANDN U20916 ( .A(y[2471]), .B(x[2471]), .Z(n35754) );
  NAND U20917 ( .A(n10005), .B(n35754), .Z(n54644) );
  XNOR U20918 ( .A(y[2470]), .B(x[2470]), .Z(n27042) );
  NANDN U20919 ( .A(x[2469]), .B(y[2469]), .Z(n27044) );
  NAND U20920 ( .A(n27042), .B(n27044), .Z(n54641) );
  NANDN U20921 ( .A(y[2468]), .B(x[2468]), .Z(n35741) );
  NANDN U20922 ( .A(y[2469]), .B(x[2469]), .Z(n27043) );
  AND U20923 ( .A(n35741), .B(n27043), .Z(n52079) );
  NANDN U20924 ( .A(y[2466]), .B(x[2466]), .Z(n10006) );
  NANDN U20925 ( .A(y[2467]), .B(x[2467]), .Z(n35742) );
  AND U20926 ( .A(n10006), .B(n35742), .Z(n54639) );
  XOR U20927 ( .A(y[2466]), .B(x[2466]), .Z(n35731) );
  NANDN U20928 ( .A(x[2465]), .B(y[2465]), .Z(n10007) );
  NANDN U20929 ( .A(n35731), .B(n10007), .Z(n54638) );
  ANDN U20930 ( .B(x[2464]), .A(y[2464]), .Z(n35725) );
  NANDN U20931 ( .A(y[2465]), .B(x[2465]), .Z(n10008) );
  NANDN U20932 ( .A(n35725), .B(n10008), .Z(n54637) );
  NANDN U20933 ( .A(x[2463]), .B(y[2463]), .Z(n27046) );
  NANDN U20934 ( .A(x[2464]), .B(y[2464]), .Z(n35730) );
  AND U20935 ( .A(n27046), .B(n35730), .Z(n52080) );
  NANDN U20936 ( .A(x[2461]), .B(y[2461]), .Z(n27051) );
  NANDN U20937 ( .A(x[2462]), .B(y[2462]), .Z(n27047) );
  AND U20938 ( .A(n27051), .B(n27047), .Z(n54635) );
  NANDN U20939 ( .A(y[2460]), .B(x[2460]), .Z(n27052) );
  NANDN U20940 ( .A(y[2461]), .B(x[2461]), .Z(n27049) );
  NAND U20941 ( .A(n27052), .B(n27049), .Z(n54634) );
  ANDN U20942 ( .B(y[2460]), .A(x[2460]), .Z(n27050) );
  NANDN U20943 ( .A(x[2457]), .B(y[2457]), .Z(n27058) );
  NANDN U20944 ( .A(y[2456]), .B(x[2456]), .Z(n35711) );
  NANDN U20945 ( .A(x[2455]), .B(y[2455]), .Z(n27061) );
  NANDN U20946 ( .A(y[2455]), .B(x[2455]), .Z(n35712) );
  NANDN U20947 ( .A(x[2453]), .B(y[2453]), .Z(n54625) );
  ANDN U20948 ( .B(y[2454]), .A(x[2454]), .Z(n27059) );
  ANDN U20949 ( .B(n54625), .A(n27059), .Z(n14001) );
  NANDN U20950 ( .A(y[2450]), .B(x[2450]), .Z(n10009) );
  NANDN U20951 ( .A(y[2451]), .B(x[2451]), .Z(n27063) );
  NAND U20952 ( .A(n10009), .B(n27063), .Z(n52083) );
  NANDN U20953 ( .A(x[2449]), .B(y[2449]), .Z(n35692) );
  XOR U20954 ( .A(y[2450]), .B(x[2450]), .Z(n35697) );
  ANDN U20955 ( .B(n35692), .A(n35697), .Z(n54623) );
  XNOR U20956 ( .A(x[2448]), .B(y[2448]), .Z(n13993) );
  ANDN U20957 ( .B(y[2447]), .A(x[2447]), .Z(n35683) );
  NANDN U20958 ( .A(y[2446]), .B(x[2446]), .Z(n10010) );
  ANDN U20959 ( .B(x[2447]), .A(y[2447]), .Z(n35690) );
  ANDN U20960 ( .B(n10010), .A(n35690), .Z(n54619) );
  ANDN U20961 ( .B(y[2441]), .A(x[2441]), .Z(n35670) );
  NANDN U20962 ( .A(x[2443]), .B(y[2443]), .Z(n13985) );
  NANDN U20963 ( .A(x[2442]), .B(y[2442]), .Z(n10011) );
  AND U20964 ( .A(n13985), .B(n10011), .Z(n35676) );
  NANDN U20965 ( .A(n35670), .B(n35676), .Z(n54614) );
  NANDN U20966 ( .A(y[2440]), .B(x[2440]), .Z(n27071) );
  NANDN U20967 ( .A(y[2441]), .B(x[2441]), .Z(n35672) );
  AND U20968 ( .A(n27071), .B(n35672), .Z(n54613) );
  ANDN U20969 ( .B(y[2439]), .A(x[2439]), .Z(n35663) );
  ANDN U20970 ( .B(y[2440]), .A(x[2440]), .Z(n35667) );
  OR U20971 ( .A(n35663), .B(n35667), .Z(n54612) );
  NANDN U20972 ( .A(y[2438]), .B(x[2438]), .Z(n27072) );
  NANDN U20973 ( .A(y[2439]), .B(x[2439]), .Z(n27070) );
  AND U20974 ( .A(n27072), .B(n27070), .Z(n54611) );
  ANDN U20975 ( .B(y[2438]), .A(x[2438]), .Z(n54610) );
  NANDN U20976 ( .A(y[2437]), .B(x[2437]), .Z(n54609) );
  NANDN U20977 ( .A(x[2436]), .B(y[2436]), .Z(n10013) );
  NANDN U20978 ( .A(x[2437]), .B(y[2437]), .Z(n10012) );
  NAND U20979 ( .A(n10013), .B(n10012), .Z(n54608) );
  ANDN U20980 ( .B(y[2435]), .A(x[2435]), .Z(n54606) );
  NANDN U20981 ( .A(y[2432]), .B(x[2432]), .Z(n27077) );
  ANDN U20982 ( .B(x[2433]), .A(y[2433]), .Z(n35654) );
  ANDN U20983 ( .B(n27077), .A(n35654), .Z(n54603) );
  NANDN U20984 ( .A(x[2431]), .B(y[2431]), .Z(n35642) );
  NANDN U20985 ( .A(x[2432]), .B(y[2432]), .Z(n35648) );
  NAND U20986 ( .A(n35642), .B(n35648), .Z(n54602) );
  NANDN U20987 ( .A(y[2430]), .B(x[2430]), .Z(n10014) );
  NANDN U20988 ( .A(y[2431]), .B(x[2431]), .Z(n27076) );
  NAND U20989 ( .A(n10014), .B(n27076), .Z(n52086) );
  XNOR U20990 ( .A(y[2430]), .B(x[2430]), .Z(n35640) );
  NANDN U20991 ( .A(x[2429]), .B(y[2429]), .Z(n35635) );
  AND U20992 ( .A(n35640), .B(n35635), .Z(n54600) );
  NANDN U20993 ( .A(x[2427]), .B(y[2427]), .Z(n54595) );
  XOR U20994 ( .A(x[2428]), .B(y[2428]), .Z(n35634) );
  ANDN U20995 ( .B(n54595), .A(n35634), .Z(n13965) );
  NANDN U20996 ( .A(y[2426]), .B(x[2426]), .Z(n10015) );
  ANDN U20997 ( .B(x[2427]), .A(y[2427]), .Z(n35631) );
  ANDN U20998 ( .B(n10015), .A(n35631), .Z(n54594) );
  XOR U20999 ( .A(y[2426]), .B(x[2426]), .Z(n35625) );
  NANDN U21000 ( .A(x[2425]), .B(y[2425]), .Z(n35621) );
  NANDN U21001 ( .A(n35625), .B(n35621), .Z(n52087) );
  ANDN U21002 ( .B(x[2424]), .A(y[2424]), .Z(n35619) );
  ANDN U21003 ( .B(x[2425]), .A(y[2425]), .Z(n35627) );
  NOR U21004 ( .A(n35619), .B(n35627), .Z(n54593) );
  NANDN U21005 ( .A(y[2419]), .B(x[2419]), .Z(n10017) );
  NANDN U21006 ( .A(y[2418]), .B(x[2418]), .Z(n10016) );
  AND U21007 ( .A(n10017), .B(n10016), .Z(n54587) );
  NANDN U21008 ( .A(x[2417]), .B(y[2417]), .Z(n10019) );
  NANDN U21009 ( .A(x[2418]), .B(y[2418]), .Z(n10018) );
  NAND U21010 ( .A(n10019), .B(n10018), .Z(n54586) );
  NANDN U21011 ( .A(y[2417]), .B(x[2417]), .Z(n10021) );
  NANDN U21012 ( .A(y[2416]), .B(x[2416]), .Z(n10020) );
  AND U21013 ( .A(n10021), .B(n10020), .Z(n54585) );
  NANDN U21014 ( .A(x[2415]), .B(y[2415]), .Z(n10023) );
  NANDN U21015 ( .A(x[2416]), .B(y[2416]), .Z(n10022) );
  NAND U21016 ( .A(n10023), .B(n10022), .Z(n35605) );
  NANDN U21017 ( .A(y[2415]), .B(x[2415]), .Z(n35603) );
  NANDN U21018 ( .A(y[2414]), .B(x[2414]), .Z(n10024) );
  AND U21019 ( .A(n35603), .B(n10024), .Z(n54583) );
  NANDN U21020 ( .A(y[2413]), .B(x[2413]), .Z(n27078) );
  ANDN U21021 ( .B(x[2412]), .A(y[2412]), .Z(n35596) );
  ANDN U21022 ( .B(n27078), .A(n35596), .Z(n54581) );
  ANDN U21023 ( .B(y[2412]), .A(x[2412]), .Z(n27080) );
  NANDN U21024 ( .A(x[2411]), .B(y[2411]), .Z(n27081) );
  NANDN U21025 ( .A(n27080), .B(n27081), .Z(n54580) );
  ANDN U21026 ( .B(x[2410]), .A(y[2410]), .Z(n35590) );
  ANDN U21027 ( .B(x[2411]), .A(y[2411]), .Z(n35597) );
  OR U21028 ( .A(n35590), .B(n35597), .Z(n52088) );
  NANDN U21029 ( .A(x[2409]), .B(y[2409]), .Z(n35586) );
  NANDN U21030 ( .A(x[2410]), .B(y[2410]), .Z(n27082) );
  AND U21031 ( .A(n35586), .B(n27082), .Z(n54578) );
  NANDN U21032 ( .A(x[2407]), .B(y[2407]), .Z(n27084) );
  NANDN U21033 ( .A(x[2408]), .B(y[2408]), .Z(n52089) );
  AND U21034 ( .A(n27084), .B(n52089), .Z(n13935) );
  ANDN U21035 ( .B(x[2406]), .A(y[2406]), .Z(n27085) );
  ANDN U21036 ( .B(y[2406]), .A(x[2406]), .Z(n27083) );
  NANDN U21037 ( .A(x[2405]), .B(y[2405]), .Z(n27088) );
  NANDN U21038 ( .A(x[2404]), .B(y[2404]), .Z(n27087) );
  NANDN U21039 ( .A(x[2403]), .B(y[2403]), .Z(n35574) );
  AND U21040 ( .A(n27087), .B(n35574), .Z(n13927) );
  ANDN U21041 ( .B(x[2402]), .A(y[2402]), .Z(n54570) );
  NANDN U21042 ( .A(x[2402]), .B(y[2402]), .Z(n35575) );
  NANDN U21043 ( .A(y[2400]), .B(x[2400]), .Z(n35564) );
  NANDN U21044 ( .A(y[2401]), .B(x[2401]), .Z(n35572) );
  NAND U21045 ( .A(n35564), .B(n35572), .Z(n54566) );
  ANDN U21046 ( .B(y[2399]), .A(x[2399]), .Z(n35559) );
  ANDN U21047 ( .B(y[2400]), .A(x[2400]), .Z(n35568) );
  NOR U21048 ( .A(n35559), .B(n35568), .Z(n54565) );
  NANDN U21049 ( .A(y[2398]), .B(x[2398]), .Z(n35556) );
  NANDN U21050 ( .A(y[2399]), .B(x[2399]), .Z(n35563) );
  NAND U21051 ( .A(n35556), .B(n35563), .Z(n54564) );
  ANDN U21052 ( .B(y[2397]), .A(x[2397]), .Z(n35553) );
  ANDN U21053 ( .B(y[2398]), .A(x[2398]), .Z(n35562) );
  NOR U21054 ( .A(n35553), .B(n35562), .Z(n54563) );
  NANDN U21055 ( .A(y[2396]), .B(x[2396]), .Z(n27089) );
  NANDN U21056 ( .A(y[2397]), .B(x[2397]), .Z(n35557) );
  NAND U21057 ( .A(n27089), .B(n35557), .Z(n54562) );
  ANDN U21058 ( .B(x[2394]), .A(y[2394]), .Z(n27090) );
  NANDN U21059 ( .A(y[2393]), .B(x[2393]), .Z(n27091) );
  NANDN U21060 ( .A(x[2393]), .B(y[2393]), .Z(n10026) );
  NANDN U21061 ( .A(x[2392]), .B(y[2392]), .Z(n10025) );
  AND U21062 ( .A(n10026), .B(n10025), .Z(n35544) );
  NANDN U21063 ( .A(y[2388]), .B(x[2388]), .Z(n27097) );
  NANDN U21064 ( .A(x[2388]), .B(y[2388]), .Z(n35537) );
  NANDN U21065 ( .A(x[2387]), .B(y[2387]), .Z(n27099) );
  AND U21066 ( .A(n35537), .B(n27099), .Z(n13897) );
  ANDN U21067 ( .B(x[2386]), .A(y[2386]), .Z(n35532) );
  NANDN U21068 ( .A(x[2386]), .B(y[2386]), .Z(n27098) );
  ANDN U21069 ( .B(x[2384]), .A(y[2384]), .Z(n54547) );
  NANDN U21070 ( .A(x[2383]), .B(y[2383]), .Z(n35524) );
  NANDN U21071 ( .A(x[2384]), .B(y[2384]), .Z(n27100) );
  AND U21072 ( .A(n35524), .B(n27100), .Z(n52091) );
  XNOR U21073 ( .A(x[2382]), .B(y[2382]), .Z(n10027) );
  ANDN U21074 ( .B(y[2381]), .A(x[2381]), .Z(n35518) );
  ANDN U21075 ( .B(n10027), .A(n35518), .Z(n54546) );
  ANDN U21076 ( .B(x[2381]), .A(y[2381]), .Z(n35522) );
  NANDN U21077 ( .A(y[2380]), .B(x[2380]), .Z(n27101) );
  NANDN U21078 ( .A(n35522), .B(n27101), .Z(n54545) );
  ANDN U21079 ( .B(y[2380]), .A(x[2380]), .Z(n35515) );
  NANDN U21080 ( .A(x[2379]), .B(y[2379]), .Z(n35509) );
  NANDN U21081 ( .A(n35515), .B(n35509), .Z(n54544) );
  NANDN U21082 ( .A(y[2378]), .B(x[2378]), .Z(n27103) );
  NANDN U21083 ( .A(y[2379]), .B(x[2379]), .Z(n27102) );
  AND U21084 ( .A(n27103), .B(n27102), .Z(n54543) );
  NANDN U21085 ( .A(x[2377]), .B(y[2377]), .Z(n35503) );
  NANDN U21086 ( .A(x[2378]), .B(y[2378]), .Z(n35510) );
  NAND U21087 ( .A(n35503), .B(n35510), .Z(n54542) );
  NANDN U21088 ( .A(y[2376]), .B(x[2376]), .Z(n27105) );
  NANDN U21089 ( .A(y[2377]), .B(x[2377]), .Z(n27104) );
  AND U21090 ( .A(n27105), .B(n27104), .Z(n54541) );
  NANDN U21091 ( .A(x[2375]), .B(y[2375]), .Z(n35497) );
  NANDN U21092 ( .A(x[2376]), .B(y[2376]), .Z(n35504) );
  NAND U21093 ( .A(n35497), .B(n35504), .Z(n54540) );
  NANDN U21094 ( .A(y[2374]), .B(x[2374]), .Z(n27107) );
  NANDN U21095 ( .A(y[2375]), .B(x[2375]), .Z(n27106) );
  NAND U21096 ( .A(n27107), .B(n27106), .Z(n54539) );
  NANDN U21097 ( .A(x[2373]), .B(y[2373]), .Z(n35491) );
  NANDN U21098 ( .A(x[2374]), .B(y[2374]), .Z(n35498) );
  AND U21099 ( .A(n35491), .B(n35498), .Z(n54538) );
  NANDN U21100 ( .A(y[2372]), .B(x[2372]), .Z(n27109) );
  NANDN U21101 ( .A(y[2373]), .B(x[2373]), .Z(n27108) );
  NAND U21102 ( .A(n27109), .B(n27108), .Z(n54537) );
  NANDN U21103 ( .A(x[2371]), .B(y[2371]), .Z(n35485) );
  NANDN U21104 ( .A(x[2372]), .B(y[2372]), .Z(n35492) );
  AND U21105 ( .A(n35485), .B(n35492), .Z(n54536) );
  NANDN U21106 ( .A(y[2370]), .B(x[2370]), .Z(n27111) );
  NANDN U21107 ( .A(y[2371]), .B(x[2371]), .Z(n27110) );
  NAND U21108 ( .A(n27111), .B(n27110), .Z(n54535) );
  NANDN U21109 ( .A(x[2369]), .B(y[2369]), .Z(n35479) );
  NANDN U21110 ( .A(x[2370]), .B(y[2370]), .Z(n35486) );
  NAND U21111 ( .A(n35479), .B(n35486), .Z(n54534) );
  NANDN U21112 ( .A(y[2368]), .B(x[2368]), .Z(n35475) );
  NANDN U21113 ( .A(y[2369]), .B(x[2369]), .Z(n27112) );
  AND U21114 ( .A(n35475), .B(n27112), .Z(n54532) );
  NANDN U21115 ( .A(x[2367]), .B(y[2367]), .Z(n35474) );
  NANDN U21116 ( .A(x[2368]), .B(y[2368]), .Z(n35480) );
  NAND U21117 ( .A(n35474), .B(n35480), .Z(n54531) );
  NANDN U21118 ( .A(y[2367]), .B(x[2367]), .Z(n35476) );
  ANDN U21119 ( .B(x[2366]), .A(y[2366]), .Z(n35472) );
  ANDN U21120 ( .B(n35476), .A(n35472), .Z(n54530) );
  NANDN U21121 ( .A(x[2361]), .B(y[2361]), .Z(n10029) );
  NANDN U21122 ( .A(x[2362]), .B(y[2362]), .Z(n10028) );
  AND U21123 ( .A(n10029), .B(n10028), .Z(n54525) );
  NANDN U21124 ( .A(y[2361]), .B(x[2361]), .Z(n10031) );
  NANDN U21125 ( .A(y[2360]), .B(x[2360]), .Z(n10030) );
  NAND U21126 ( .A(n10031), .B(n10030), .Z(n54524) );
  NANDN U21127 ( .A(x[2359]), .B(y[2359]), .Z(n10033) );
  NANDN U21128 ( .A(x[2360]), .B(y[2360]), .Z(n10032) );
  AND U21129 ( .A(n10033), .B(n10032), .Z(n54523) );
  NANDN U21130 ( .A(y[2358]), .B(x[2358]), .Z(n10034) );
  ANDN U21131 ( .B(x[2359]), .A(y[2359]), .Z(n27115) );
  ANDN U21132 ( .B(n10034), .A(n27115), .Z(n54522) );
  NANDN U21133 ( .A(x[2357]), .B(y[2357]), .Z(n27118) );
  XNOR U21134 ( .A(x[2358]), .B(y[2358]), .Z(n10035) );
  NAND U21135 ( .A(n27118), .B(n10035), .Z(n54521) );
  NANDN U21136 ( .A(y[2356]), .B(x[2356]), .Z(n27120) );
  NANDN U21137 ( .A(y[2357]), .B(x[2357]), .Z(n27117) );
  AND U21138 ( .A(n27120), .B(n27117), .Z(n54520) );
  NANDN U21139 ( .A(x[2355]), .B(y[2355]), .Z(n35453) );
  NANDN U21140 ( .A(x[2356]), .B(y[2356]), .Z(n27119) );
  NAND U21141 ( .A(n35453), .B(n27119), .Z(n54519) );
  NANDN U21142 ( .A(y[2354]), .B(x[2354]), .Z(n27122) );
  NANDN U21143 ( .A(y[2355]), .B(x[2355]), .Z(n27121) );
  AND U21144 ( .A(n27122), .B(n27121), .Z(n54518) );
  NANDN U21145 ( .A(x[2353]), .B(y[2353]), .Z(n35447) );
  NANDN U21146 ( .A(x[2354]), .B(y[2354]), .Z(n35454) );
  NAND U21147 ( .A(n35447), .B(n35454), .Z(n54517) );
  NANDN U21148 ( .A(x[2351]), .B(y[2351]), .Z(n35440) );
  NANDN U21149 ( .A(x[2352]), .B(y[2352]), .Z(n35448) );
  NAND U21150 ( .A(n35440), .B(n35448), .Z(n52094) );
  NANDN U21151 ( .A(y[2350]), .B(x[2350]), .Z(n10036) );
  NANDN U21152 ( .A(y[2351]), .B(x[2351]), .Z(n35444) );
  NAND U21153 ( .A(n10036), .B(n35444), .Z(n54515) );
  XNOR U21154 ( .A(y[2350]), .B(x[2350]), .Z(n27125) );
  NANDN U21155 ( .A(x[2349]), .B(y[2349]), .Z(n27126) );
  AND U21156 ( .A(n27125), .B(n27126), .Z(n54514) );
  NANDN U21157 ( .A(y[2348]), .B(x[2348]), .Z(n27128) );
  NANDN U21158 ( .A(y[2349]), .B(x[2349]), .Z(n27124) );
  NAND U21159 ( .A(n27128), .B(n27124), .Z(n54513) );
  NANDN U21160 ( .A(y[2346]), .B(x[2346]), .Z(n27133) );
  NANDN U21161 ( .A(y[2347]), .B(x[2347]), .Z(n27129) );
  NAND U21162 ( .A(n27133), .B(n27129), .Z(n52096) );
  NANDN U21163 ( .A(x[2345]), .B(y[2345]), .Z(n27134) );
  NANDN U21164 ( .A(x[2346]), .B(y[2346]), .Z(n27131) );
  NAND U21165 ( .A(n27134), .B(n27131), .Z(n54512) );
  NANDN U21166 ( .A(y[2344]), .B(x[2344]), .Z(n35424) );
  NANDN U21167 ( .A(y[2345]), .B(x[2345]), .Z(n27132) );
  AND U21168 ( .A(n35424), .B(n27132), .Z(n54511) );
  NANDN U21169 ( .A(x[2343]), .B(y[2343]), .Z(n35419) );
  NANDN U21170 ( .A(x[2344]), .B(y[2344]), .Z(n27135) );
  NAND U21171 ( .A(n35419), .B(n27135), .Z(n54510) );
  NANDN U21172 ( .A(x[2341]), .B(y[2341]), .Z(n35413) );
  NANDN U21173 ( .A(x[2342]), .B(y[2342]), .Z(n35420) );
  NAND U21174 ( .A(n35413), .B(n35420), .Z(n52098) );
  NANDN U21175 ( .A(y[2340]), .B(x[2340]), .Z(n35409) );
  NANDN U21176 ( .A(y[2341]), .B(x[2341]), .Z(n27137) );
  NAND U21177 ( .A(n35409), .B(n27137), .Z(n54509) );
  NANDN U21178 ( .A(x[2339]), .B(y[2339]), .Z(n35407) );
  NANDN U21179 ( .A(x[2340]), .B(y[2340]), .Z(n35414) );
  AND U21180 ( .A(n35407), .B(n35414), .Z(n54508) );
  ANDN U21181 ( .B(x[2338]), .A(y[2338]), .Z(n35405) );
  NANDN U21182 ( .A(y[2339]), .B(x[2339]), .Z(n35410) );
  NANDN U21183 ( .A(n35405), .B(n35410), .Z(n54507) );
  NANDN U21184 ( .A(x[2337]), .B(y[2337]), .Z(n27138) );
  NANDN U21185 ( .A(x[2338]), .B(y[2338]), .Z(n54506) );
  AND U21186 ( .A(n27138), .B(n54506), .Z(n13835) );
  ANDN U21187 ( .B(x[2337]), .A(y[2337]), .Z(n54505) );
  NANDN U21188 ( .A(x[2336]), .B(y[2336]), .Z(n27139) );
  ANDN U21189 ( .B(x[2334]), .A(y[2334]), .Z(n35397) );
  NANDN U21190 ( .A(y[2333]), .B(x[2333]), .Z(n35398) );
  XNOR U21191 ( .A(y[2333]), .B(x[2333]), .Z(n13825) );
  ANDN U21192 ( .B(x[2332]), .A(y[2332]), .Z(n54499) );
  NANDN U21193 ( .A(x[2332]), .B(y[2332]), .Z(n35394) );
  NANDN U21194 ( .A(y[2330]), .B(x[2330]), .Z(n35385) );
  NANDN U21195 ( .A(y[2331]), .B(x[2331]), .Z(n35392) );
  NAND U21196 ( .A(n35385), .B(n35392), .Z(n52100) );
  NANDN U21197 ( .A(x[2329]), .B(y[2329]), .Z(n27145) );
  ANDN U21198 ( .B(y[2330]), .A(x[2330]), .Z(n35390) );
  ANDN U21199 ( .B(n27145), .A(n35390), .Z(n54497) );
  NANDN U21200 ( .A(y[2326]), .B(x[2326]), .Z(n35372) );
  NANDN U21201 ( .A(y[2327]), .B(x[2327]), .Z(n35379) );
  NAND U21202 ( .A(n35372), .B(n35379), .Z(n54495) );
  NANDN U21203 ( .A(x[2325]), .B(y[2325]), .Z(n27150) );
  NANDN U21204 ( .A(x[2326]), .B(y[2326]), .Z(n27148) );
  NAND U21205 ( .A(n27150), .B(n27148), .Z(n54494) );
  NANDN U21206 ( .A(y[2324]), .B(x[2324]), .Z(n35367) );
  NANDN U21207 ( .A(y[2325]), .B(x[2325]), .Z(n35373) );
  AND U21208 ( .A(n35367), .B(n35373), .Z(n52102) );
  NANDN U21209 ( .A(y[2322]), .B(x[2322]), .Z(n35361) );
  ANDN U21210 ( .B(x[2323]), .A(y[2323]), .Z(n35369) );
  ANDN U21211 ( .B(n35361), .A(n35369), .Z(n54491) );
  ANDN U21212 ( .B(x[2318]), .A(y[2318]), .Z(n27152) );
  NANDN U21213 ( .A(x[2319]), .B(y[2319]), .Z(n10040) );
  NAND U21214 ( .A(n27152), .B(n10040), .Z(n13806) );
  XNOR U21215 ( .A(x[2320]), .B(y[2320]), .Z(n10038) );
  NANDN U21216 ( .A(y[2319]), .B(x[2319]), .Z(n10037) );
  NAND U21217 ( .A(n10038), .B(n10037), .Z(n27156) );
  NANDN U21218 ( .A(x[2318]), .B(y[2318]), .Z(n10039) );
  AND U21219 ( .A(n10040), .B(n10039), .Z(n27154) );
  NANDN U21220 ( .A(x[2317]), .B(y[2317]), .Z(n10041) );
  AND U21221 ( .A(n27154), .B(n10041), .Z(n54485) );
  ANDN U21222 ( .B(x[2317]), .A(y[2317]), .Z(n27151) );
  ANDN U21223 ( .B(y[2316]), .A(x[2316]), .Z(n35355) );
  NANDN U21224 ( .A(x[2315]), .B(y[2315]), .Z(n27158) );
  NANDN U21225 ( .A(n35355), .B(n27158), .Z(n54487) );
  NANDN U21226 ( .A(x[2313]), .B(y[2313]), .Z(n35347) );
  NANDN U21227 ( .A(x[2314]), .B(y[2314]), .Z(n54482) );
  AND U21228 ( .A(n35347), .B(n54482), .Z(n54481) );
  ANDN U21229 ( .B(x[2312]), .A(y[2312]), .Z(n54480) );
  NANDN U21230 ( .A(x[2311]), .B(y[2311]), .Z(n35340) );
  ANDN U21231 ( .B(y[2312]), .A(x[2312]), .Z(n35349) );
  ANDN U21232 ( .B(n35340), .A(n35349), .Z(n54479) );
  ANDN U21233 ( .B(x[2310]), .A(y[2310]), .Z(n27162) );
  ANDN U21234 ( .B(x[2311]), .A(y[2311]), .Z(n35345) );
  OR U21235 ( .A(n27162), .B(n35345), .Z(n54477) );
  NANDN U21236 ( .A(x[2310]), .B(y[2310]), .Z(n35339) );
  ANDN U21237 ( .B(y[2309]), .A(x[2309]), .Z(n35334) );
  ANDN U21238 ( .B(n35339), .A(n35334), .Z(n54476) );
  ANDN U21239 ( .B(x[2309]), .A(y[2309]), .Z(n27161) );
  NANDN U21240 ( .A(y[2308]), .B(x[2308]), .Z(n27163) );
  NANDN U21241 ( .A(n27161), .B(n27163), .Z(n54475) );
  NANDN U21242 ( .A(x[2307]), .B(y[2307]), .Z(n35329) );
  ANDN U21243 ( .B(y[2308]), .A(x[2308]), .Z(n35335) );
  ANDN U21244 ( .B(n35329), .A(n35335), .Z(n54474) );
  NANDN U21245 ( .A(y[2306]), .B(x[2306]), .Z(n10042) );
  NANDN U21246 ( .A(y[2307]), .B(x[2307]), .Z(n27164) );
  NAND U21247 ( .A(n10042), .B(n27164), .Z(n54473) );
  XNOR U21248 ( .A(x[2306]), .B(y[2306]), .Z(n35325) );
  ANDN U21249 ( .B(x[2304]), .A(y[2304]), .Z(n35320) );
  NANDN U21250 ( .A(y[2305]), .B(x[2305]), .Z(n35324) );
  NANDN U21251 ( .A(n35320), .B(n35324), .Z(n52107) );
  NANDN U21252 ( .A(x[2303]), .B(y[2303]), .Z(n27165) );
  NANDN U21253 ( .A(x[2304]), .B(y[2304]), .Z(n35322) );
  AND U21254 ( .A(n27165), .B(n35322), .Z(n52108) );
  NANDN U21255 ( .A(y[2300]), .B(x[2300]), .Z(n10043) );
  NANDN U21256 ( .A(y[2301]), .B(x[2301]), .Z(n35312) );
  NAND U21257 ( .A(n10043), .B(n35312), .Z(n54471) );
  ANDN U21258 ( .B(x[2298]), .A(y[2298]), .Z(n35302) );
  ANDN U21259 ( .B(x[2299]), .A(y[2299]), .Z(n35307) );
  NOR U21260 ( .A(n35302), .B(n35307), .Z(n54467) );
  NANDN U21261 ( .A(x[2297]), .B(y[2297]), .Z(n27170) );
  NANDN U21262 ( .A(x[2298]), .B(y[2298]), .Z(n35304) );
  NAND U21263 ( .A(n27170), .B(n35304), .Z(n52110) );
  ANDN U21264 ( .B(x[2297]), .A(y[2297]), .Z(n35299) );
  NANDN U21265 ( .A(y[2296]), .B(x[2296]), .Z(n35294) );
  NANDN U21266 ( .A(n35299), .B(n35294), .Z(n54465) );
  NANDN U21267 ( .A(x[2296]), .B(y[2296]), .Z(n27169) );
  ANDN U21268 ( .B(y[2295]), .A(x[2295]), .Z(n35290) );
  ANDN U21269 ( .B(n27169), .A(n35290), .Z(n54464) );
  ANDN U21270 ( .B(x[2295]), .A(y[2295]), .Z(n35296) );
  NANDN U21271 ( .A(y[2294]), .B(x[2294]), .Z(n27172) );
  NANDN U21272 ( .A(n35296), .B(n27172), .Z(n54463) );
  NANDN U21273 ( .A(x[2293]), .B(y[2293]), .Z(n27174) );
  NANDN U21274 ( .A(x[2294]), .B(y[2294]), .Z(n35291) );
  AND U21275 ( .A(n27174), .B(n35291), .Z(n13774) );
  ANDN U21276 ( .B(x[2293]), .A(y[2293]), .Z(n27171) );
  NANDN U21277 ( .A(x[2292]), .B(y[2292]), .Z(n27173) );
  NANDN U21278 ( .A(y[2290]), .B(x[2290]), .Z(n27178) );
  NANDN U21279 ( .A(y[2291]), .B(x[2291]), .Z(n27176) );
  NAND U21280 ( .A(n27178), .B(n27176), .Z(n54457) );
  NANDN U21281 ( .A(x[2289]), .B(y[2289]), .Z(n27180) );
  ANDN U21282 ( .B(y[2290]), .A(x[2290]), .Z(n35283) );
  ANDN U21283 ( .B(n27180), .A(n35283), .Z(n54456) );
  NANDN U21284 ( .A(y[2288]), .B(x[2288]), .Z(n10044) );
  NANDN U21285 ( .A(y[2289]), .B(x[2289]), .Z(n27179) );
  NAND U21286 ( .A(n10044), .B(n27179), .Z(n54455) );
  XNOR U21287 ( .A(y[2288]), .B(x[2288]), .Z(n35274) );
  NANDN U21288 ( .A(x[2287]), .B(y[2287]), .Z(n35270) );
  AND U21289 ( .A(n35274), .B(n35270), .Z(n54454) );
  NANDN U21290 ( .A(y[2286]), .B(x[2286]), .Z(n27182) );
  NANDN U21291 ( .A(y[2287]), .B(x[2287]), .Z(n35275) );
  NAND U21292 ( .A(n27182), .B(n35275), .Z(n54453) );
  NANDN U21293 ( .A(x[2286]), .B(y[2286]), .Z(n54452) );
  NANDN U21294 ( .A(y[2285]), .B(x[2285]), .Z(n52111) );
  NANDN U21295 ( .A(y[2284]), .B(x[2284]), .Z(n10045) );
  NAND U21296 ( .A(n52111), .B(n10045), .Z(n13761) );
  NANDN U21297 ( .A(x[2284]), .B(y[2284]), .Z(n27184) );
  NANDN U21298 ( .A(x[2283]), .B(y[2283]), .Z(n35263) );
  AND U21299 ( .A(n27184), .B(n35263), .Z(n13759) );
  ANDN U21300 ( .B(x[2282]), .A(y[2282]), .Z(n13756) );
  XNOR U21301 ( .A(x[2282]), .B(y[2282]), .Z(n27190) );
  ANDN U21302 ( .B(y[2281]), .A(x[2281]), .Z(n54447) );
  ANDN U21303 ( .B(n27190), .A(n54447), .Z(n13754) );
  ANDN U21304 ( .B(x[2280]), .A(y[2280]), .Z(n54446) );
  NANDN U21305 ( .A(x[2279]), .B(y[2279]), .Z(n35253) );
  NANDN U21306 ( .A(x[2280]), .B(y[2280]), .Z(n35260) );
  AND U21307 ( .A(n35253), .B(n35260), .Z(n54445) );
  ANDN U21308 ( .B(x[2279]), .A(y[2279]), .Z(n35258) );
  NANDN U21309 ( .A(y[2278]), .B(x[2278]), .Z(n27192) );
  NANDN U21310 ( .A(n35258), .B(n27192), .Z(n54444) );
  NANDN U21311 ( .A(y[2276]), .B(x[2276]), .Z(n27196) );
  NANDN U21312 ( .A(y[2277]), .B(x[2277]), .Z(n27191) );
  NAND U21313 ( .A(n27196), .B(n27191), .Z(n52114) );
  NANDN U21314 ( .A(x[2276]), .B(y[2276]), .Z(n27194) );
  ANDN U21315 ( .B(y[2275]), .A(x[2275]), .Z(n35243) );
  ANDN U21316 ( .B(n27194), .A(n35243), .Z(n54443) );
  NANDN U21317 ( .A(x[2273]), .B(y[2273]), .Z(n27198) );
  NANDN U21318 ( .A(x[2274]), .B(y[2274]), .Z(n35244) );
  AND U21319 ( .A(n27198), .B(n35244), .Z(n13744) );
  ANDN U21320 ( .B(x[2272]), .A(y[2272]), .Z(n27200) );
  NANDN U21321 ( .A(y[2273]), .B(x[2273]), .Z(n54440) );
  ANDN U21322 ( .B(y[2271]), .A(x[2271]), .Z(n27202) );
  NANDN U21323 ( .A(y[2271]), .B(x[2271]), .Z(n27201) );
  XNOR U21324 ( .A(x[2270]), .B(y[2270]), .Z(n27205) );
  NANDN U21325 ( .A(x[2269]), .B(y[2269]), .Z(n27206) );
  AND U21326 ( .A(n27205), .B(n27206), .Z(n13735) );
  ANDN U21327 ( .B(x[2268]), .A(y[2268]), .Z(n35228) );
  NANDN U21328 ( .A(x[2268]), .B(y[2268]), .Z(n35233) );
  ANDN U21329 ( .B(y[2267]), .A(x[2267]), .Z(n35227) );
  ANDN U21330 ( .B(n35233), .A(n35227), .Z(n54432) );
  NANDN U21331 ( .A(x[2265]), .B(y[2265]), .Z(n35218) );
  ANDN U21332 ( .B(y[2266]), .A(x[2266]), .Z(n35224) );
  ANDN U21333 ( .B(n35218), .A(n35224), .Z(n54430) );
  NANDN U21334 ( .A(y[2264]), .B(x[2264]), .Z(n35214) );
  NANDN U21335 ( .A(y[2265]), .B(x[2265]), .Z(n27208) );
  NAND U21336 ( .A(n35214), .B(n27208), .Z(n54429) );
  NANDN U21337 ( .A(x[2263]), .B(y[2263]), .Z(n35211) );
  NANDN U21338 ( .A(x[2264]), .B(y[2264]), .Z(n35219) );
  NAND U21339 ( .A(n35211), .B(n35219), .Z(n52115) );
  NANDN U21340 ( .A(y[2262]), .B(x[2262]), .Z(n10046) );
  NANDN U21341 ( .A(y[2263]), .B(x[2263]), .Z(n35215) );
  AND U21342 ( .A(n10046), .B(n35215), .Z(n54428) );
  ANDN U21343 ( .B(x[2260]), .A(y[2260]), .Z(n35200) );
  ANDN U21344 ( .B(x[2261]), .A(y[2261]), .Z(n35207) );
  NOR U21345 ( .A(n35200), .B(n35207), .Z(n54426) );
  NANDN U21346 ( .A(x[2259]), .B(y[2259]), .Z(n35197) );
  NANDN U21347 ( .A(x[2260]), .B(y[2260]), .Z(n27210) );
  NAND U21348 ( .A(n35197), .B(n27210), .Z(n54425) );
  ANDN U21349 ( .B(x[2259]), .A(y[2259]), .Z(n35203) );
  NANDN U21350 ( .A(y[2258]), .B(x[2258]), .Z(n10047) );
  NANDN U21351 ( .A(n35203), .B(n10047), .Z(n52116) );
  XNOR U21352 ( .A(x[2258]), .B(y[2258]), .Z(n35193) );
  ANDN U21353 ( .B(y[2257]), .A(x[2257]), .Z(n35189) );
  ANDN U21354 ( .B(n35193), .A(n35189), .Z(n54424) );
  NANDN U21355 ( .A(x[2255]), .B(y[2255]), .Z(n27213) );
  NANDN U21356 ( .A(x[2256]), .B(y[2256]), .Z(n35190) );
  AND U21357 ( .A(n27213), .B(n35190), .Z(n13719) );
  ANDN U21358 ( .B(x[2255]), .A(y[2255]), .Z(n27211) );
  NANDN U21359 ( .A(x[2254]), .B(y[2254]), .Z(n27214) );
  ANDN U21360 ( .B(x[2252]), .A(y[2252]), .Z(n27217) );
  ANDN U21361 ( .B(x[2250]), .A(y[2250]), .Z(n35172) );
  NANDN U21362 ( .A(x[2249]), .B(y[2249]), .Z(n27220) );
  ANDN U21363 ( .B(y[2250]), .A(x[2250]), .Z(n35177) );
  ANDN U21364 ( .B(n27220), .A(n35177), .Z(n54412) );
  NANDN U21365 ( .A(y[2243]), .B(x[2243]), .Z(n54405) );
  NANDN U21366 ( .A(y[2244]), .B(x[2244]), .Z(n54408) );
  AND U21367 ( .A(n54405), .B(n54408), .Z(n35160) );
  NANDN U21368 ( .A(x[2242]), .B(y[2242]), .Z(n52123) );
  NANDN U21369 ( .A(x[2243]), .B(y[2243]), .Z(n52119) );
  NAND U21370 ( .A(n52123), .B(n52119), .Z(n35158) );
  NANDN U21371 ( .A(y[2241]), .B(x[2241]), .Z(n54403) );
  NANDN U21372 ( .A(y[2242]), .B(x[2242]), .Z(n52121) );
  AND U21373 ( .A(n54403), .B(n52121), .Z(n35155) );
  ANDN U21374 ( .B(x[2238]), .A(y[2238]), .Z(n35142) );
  ANDN U21375 ( .B(x[2239]), .A(y[2239]), .Z(n35152) );
  NOR U21376 ( .A(n35142), .B(n35152), .Z(n54400) );
  ANDN U21377 ( .B(x[2236]), .A(y[2236]), .Z(n35135) );
  ANDN U21378 ( .B(x[2237]), .A(y[2237]), .Z(n35145) );
  NOR U21379 ( .A(n35135), .B(n35145), .Z(n54399) );
  NANDN U21380 ( .A(x[2235]), .B(y[2235]), .Z(n35131) );
  NANDN U21381 ( .A(x[2236]), .B(y[2236]), .Z(n35140) );
  NAND U21382 ( .A(n35131), .B(n35140), .Z(n54397) );
  ANDN U21383 ( .B(x[2235]), .A(y[2235]), .Z(n35137) );
  NANDN U21384 ( .A(y[2234]), .B(x[2234]), .Z(n27225) );
  NANDN U21385 ( .A(n35137), .B(n27225), .Z(n54396) );
  NANDN U21386 ( .A(x[2233]), .B(y[2233]), .Z(n35125) );
  NANDN U21387 ( .A(x[2234]), .B(y[2234]), .Z(n35130) );
  AND U21388 ( .A(n35125), .B(n35130), .Z(n52125) );
  NANDN U21389 ( .A(y[2230]), .B(x[2230]), .Z(n10049) );
  NANDN U21390 ( .A(y[2231]), .B(x[2231]), .Z(n10048) );
  NAND U21391 ( .A(n10049), .B(n10048), .Z(n27227) );
  NANDN U21392 ( .A(x[2230]), .B(y[2230]), .Z(n10051) );
  NANDN U21393 ( .A(x[2229]), .B(y[2229]), .Z(n10050) );
  AND U21394 ( .A(n10051), .B(n10050), .Z(n27228) );
  NANDN U21395 ( .A(y[2228]), .B(x[2228]), .Z(n10053) );
  NANDN U21396 ( .A(y[2229]), .B(x[2229]), .Z(n10052) );
  NAND U21397 ( .A(n10053), .B(n10052), .Z(n27229) );
  NANDN U21398 ( .A(x[2227]), .B(y[2227]), .Z(n27230) );
  ANDN U21399 ( .B(y[2228]), .A(x[2228]), .Z(n35116) );
  ANDN U21400 ( .B(n27230), .A(n35116), .Z(n54390) );
  ANDN U21401 ( .B(x[2224]), .A(y[2224]), .Z(n35104) );
  NANDN U21402 ( .A(y[2225]), .B(x[2225]), .Z(n27232) );
  NANDN U21403 ( .A(n35104), .B(n27232), .Z(n54388) );
  NANDN U21404 ( .A(x[2223]), .B(y[2223]), .Z(n27236) );
  NANDN U21405 ( .A(x[2224]), .B(y[2224]), .Z(n27234) );
  NAND U21406 ( .A(n27236), .B(n27234), .Z(n54387) );
  ANDN U21407 ( .B(x[2222]), .A(y[2222]), .Z(n35100) );
  ANDN U21408 ( .B(x[2223]), .A(y[2223]), .Z(n35105) );
  NOR U21409 ( .A(n35100), .B(n35105), .Z(n54386) );
  NANDN U21410 ( .A(y[2219]), .B(x[2219]), .Z(n35093) );
  ANDN U21411 ( .B(x[2218]), .A(y[2218]), .Z(n35088) );
  ANDN U21412 ( .B(n35093), .A(n35088), .Z(n54382) );
  NANDN U21413 ( .A(x[2216]), .B(y[2216]), .Z(n10055) );
  NANDN U21414 ( .A(x[2217]), .B(y[2217]), .Z(n10054) );
  NAND U21415 ( .A(n10055), .B(n10054), .Z(n27239) );
  NANDN U21416 ( .A(y[2216]), .B(x[2216]), .Z(n10057) );
  NANDN U21417 ( .A(y[2215]), .B(x[2215]), .Z(n10056) );
  AND U21418 ( .A(n10057), .B(n10056), .Z(n35084) );
  NANDN U21419 ( .A(x[2214]), .B(y[2214]), .Z(n10059) );
  NANDN U21420 ( .A(x[2215]), .B(y[2215]), .Z(n10058) );
  NAND U21421 ( .A(n10059), .B(n10058), .Z(n35082) );
  NANDN U21422 ( .A(y[2214]), .B(x[2214]), .Z(n10061) );
  NANDN U21423 ( .A(y[2213]), .B(x[2213]), .Z(n10060) );
  NAND U21424 ( .A(n10061), .B(n10060), .Z(n54376) );
  XOR U21425 ( .A(x[2212]), .B(y[2212]), .Z(n13659) );
  NANDN U21426 ( .A(y[2210]), .B(x[2210]), .Z(n10062) );
  AND U21427 ( .A(n27242), .B(n10062), .Z(n54375) );
  ANDN U21428 ( .B(y[2209]), .A(x[2209]), .Z(n52130) );
  NANDN U21429 ( .A(y[2208]), .B(x[2208]), .Z(n10063) );
  ANDN U21430 ( .B(x[2209]), .A(y[2209]), .Z(n35079) );
  ANDN U21431 ( .B(n10063), .A(n35079), .Z(n54374) );
  XNOR U21432 ( .A(y[2208]), .B(x[2208]), .Z(n35071) );
  NANDN U21433 ( .A(x[2207]), .B(y[2207]), .Z(n27244) );
  NAND U21434 ( .A(n35071), .B(n27244), .Z(n52131) );
  NANDN U21435 ( .A(y[2206]), .B(x[2206]), .Z(n35064) );
  NANDN U21436 ( .A(y[2207]), .B(x[2207]), .Z(n35073) );
  AND U21437 ( .A(n35064), .B(n35073), .Z(n54372) );
  NANDN U21438 ( .A(x[2203]), .B(y[2203]), .Z(n35055) );
  NANDN U21439 ( .A(x[2204]), .B(y[2204]), .Z(n27246) );
  NAND U21440 ( .A(n35055), .B(n27246), .Z(n54368) );
  ANDN U21441 ( .B(x[2202]), .A(y[2202]), .Z(n35051) );
  ANDN U21442 ( .B(x[2203]), .A(y[2203]), .Z(n35061) );
  OR U21443 ( .A(n35051), .B(n35061), .Z(n52133) );
  NANDN U21444 ( .A(x[2201]), .B(y[2201]), .Z(n35047) );
  ANDN U21445 ( .B(y[2202]), .A(x[2202]), .Z(n35057) );
  ANDN U21446 ( .B(n35047), .A(n35057), .Z(n54367) );
  ANDN U21447 ( .B(x[2199]), .A(y[2199]), .Z(n54364) );
  NANDN U21448 ( .A(x[2199]), .B(y[2199]), .Z(n10065) );
  NANDN U21449 ( .A(x[2198]), .B(y[2198]), .Z(n10064) );
  AND U21450 ( .A(n10065), .B(n10064), .Z(n52134) );
  NANDN U21451 ( .A(y[2197]), .B(x[2197]), .Z(n10067) );
  NANDN U21452 ( .A(y[2198]), .B(x[2198]), .Z(n10066) );
  NAND U21453 ( .A(n10067), .B(n10066), .Z(n54363) );
  NANDN U21454 ( .A(x[2197]), .B(y[2197]), .Z(n10069) );
  NANDN U21455 ( .A(x[2196]), .B(y[2196]), .Z(n10068) );
  AND U21456 ( .A(n10069), .B(n10068), .Z(n54362) );
  NANDN U21457 ( .A(y[2195]), .B(x[2195]), .Z(n10071) );
  NANDN U21458 ( .A(y[2196]), .B(x[2196]), .Z(n10070) );
  NAND U21459 ( .A(n10071), .B(n10070), .Z(n54361) );
  NANDN U21460 ( .A(x[2195]), .B(y[2195]), .Z(n10073) );
  NANDN U21461 ( .A(x[2194]), .B(y[2194]), .Z(n10072) );
  AND U21462 ( .A(n10073), .B(n10072), .Z(n54360) );
  NANDN U21463 ( .A(y[2193]), .B(x[2193]), .Z(n10075) );
  NANDN U21464 ( .A(y[2194]), .B(x[2194]), .Z(n10074) );
  NAND U21465 ( .A(n10075), .B(n10074), .Z(n54358) );
  NANDN U21466 ( .A(x[2193]), .B(y[2193]), .Z(n10077) );
  NANDN U21467 ( .A(x[2192]), .B(y[2192]), .Z(n10076) );
  AND U21468 ( .A(n10077), .B(n10076), .Z(n54357) );
  NANDN U21469 ( .A(y[2192]), .B(x[2192]), .Z(n27249) );
  ANDN U21470 ( .B(y[2191]), .A(x[2191]), .Z(n35032) );
  NANDN U21471 ( .A(y[2191]), .B(x[2191]), .Z(n27248) );
  XNOR U21472 ( .A(y[2190]), .B(x[2190]), .Z(n35029) );
  NANDN U21473 ( .A(x[2189]), .B(y[2189]), .Z(n35025) );
  NAND U21474 ( .A(n35029), .B(n35025), .Z(n52136) );
  NANDN U21475 ( .A(y[2188]), .B(x[2188]), .Z(n10078) );
  NANDN U21476 ( .A(y[2189]), .B(x[2189]), .Z(n35028) );
  AND U21477 ( .A(n10078), .B(n35028), .Z(n52137) );
  NANDN U21478 ( .A(y[2186]), .B(x[2186]), .Z(n10079) );
  ANDN U21479 ( .B(x[2187]), .A(y[2187]), .Z(n35023) );
  ANDN U21480 ( .B(n10079), .A(n35023), .Z(n54354) );
  XOR U21481 ( .A(y[2186]), .B(x[2186]), .Z(n35015) );
  NANDN U21482 ( .A(x[2185]), .B(y[2185]), .Z(n35009) );
  NANDN U21483 ( .A(n35015), .B(n35009), .Z(n54353) );
  ANDN U21484 ( .B(x[2184]), .A(y[2184]), .Z(n35005) );
  ANDN U21485 ( .B(x[2185]), .A(y[2185]), .Z(n35012) );
  OR U21486 ( .A(n35005), .B(n35012), .Z(n54352) );
  NANDN U21487 ( .A(x[2183]), .B(y[2183]), .Z(n27250) );
  NANDN U21488 ( .A(x[2184]), .B(y[2184]), .Z(n35010) );
  AND U21489 ( .A(n27250), .B(n35010), .Z(n52139) );
  ANDN U21490 ( .B(x[2181]), .A(y[2181]), .Z(n35000) );
  NANDN U21491 ( .A(y[2180]), .B(x[2180]), .Z(n27252) );
  NANDN U21492 ( .A(n35000), .B(n27252), .Z(n54348) );
  NANDN U21493 ( .A(y[2179]), .B(x[2179]), .Z(n54346) );
  NANDN U21494 ( .A(x[2178]), .B(y[2178]), .Z(n52142) );
  NANDN U21495 ( .A(x[2179]), .B(y[2179]), .Z(n52141) );
  AND U21496 ( .A(n52142), .B(n52141), .Z(n34991) );
  ANDN U21497 ( .B(x[2178]), .A(y[2178]), .Z(n54345) );
  NANDN U21498 ( .A(x[2177]), .B(y[2177]), .Z(n52143) );
  ANDN U21499 ( .B(x[2176]), .A(y[2176]), .Z(n27254) );
  ANDN U21500 ( .B(x[2177]), .A(y[2177]), .Z(n34988) );
  OR U21501 ( .A(n27254), .B(n34988), .Z(n54344) );
  NANDN U21502 ( .A(x[2176]), .B(y[2176]), .Z(n34984) );
  ANDN U21503 ( .B(y[2175]), .A(x[2175]), .Z(n34979) );
  ANDN U21504 ( .B(n34984), .A(n34979), .Z(n54343) );
  ANDN U21505 ( .B(x[2175]), .A(y[2175]), .Z(n27253) );
  NANDN U21506 ( .A(y[2174]), .B(x[2174]), .Z(n27255) );
  NANDN U21507 ( .A(n27253), .B(n27255), .Z(n54342) );
  ANDN U21508 ( .B(y[2173]), .A(x[2173]), .Z(n34974) );
  ANDN U21509 ( .B(y[2174]), .A(x[2174]), .Z(n34980) );
  NOR U21510 ( .A(n34974), .B(n34980), .Z(n54341) );
  NANDN U21511 ( .A(y[2172]), .B(x[2172]), .Z(n34971) );
  NANDN U21512 ( .A(y[2173]), .B(x[2173]), .Z(n27256) );
  NAND U21513 ( .A(n34971), .B(n27256), .Z(n54340) );
  NANDN U21514 ( .A(y[2171]), .B(x[2171]), .Z(n54338) );
  NANDN U21515 ( .A(y[2170]), .B(x[2170]), .Z(n34966) );
  NAND U21516 ( .A(n54338), .B(n34966), .Z(n54336) );
  NANDN U21517 ( .A(x[2169]), .B(y[2169]), .Z(n54334) );
  ANDN U21518 ( .B(x[2168]), .A(y[2168]), .Z(n34961) );
  ANDN U21519 ( .B(x[2169]), .A(y[2169]), .Z(n34968) );
  OR U21520 ( .A(n34961), .B(n34968), .Z(n54333) );
  NANDN U21521 ( .A(x[2167]), .B(y[2167]), .Z(n27259) );
  ANDN U21522 ( .B(y[2168]), .A(x[2168]), .Z(n34964) );
  ANDN U21523 ( .B(n27259), .A(n34964), .Z(n54332) );
  ANDN U21524 ( .B(x[2167]), .A(y[2167]), .Z(n34958) );
  NANDN U21525 ( .A(y[2166]), .B(x[2166]), .Z(n34952) );
  NANDN U21526 ( .A(n34958), .B(n34952), .Z(n54331) );
  NANDN U21527 ( .A(x[2165]), .B(y[2165]), .Z(n27262) );
  NANDN U21528 ( .A(x[2166]), .B(y[2166]), .Z(n27260) );
  AND U21529 ( .A(n27262), .B(n27260), .Z(n54330) );
  ANDN U21530 ( .B(x[2164]), .A(y[2164]), .Z(n34947) );
  NANDN U21531 ( .A(y[2165]), .B(x[2165]), .Z(n34953) );
  NANDN U21532 ( .A(n34947), .B(n34953), .Z(n54329) );
  NANDN U21533 ( .A(x[2162]), .B(y[2162]), .Z(n10081) );
  NANDN U21534 ( .A(x[2163]), .B(y[2163]), .Z(n10080) );
  NAND U21535 ( .A(n10081), .B(n10080), .Z(n27263) );
  NANDN U21536 ( .A(y[2162]), .B(x[2162]), .Z(n10083) );
  NANDN U21537 ( .A(y[2161]), .B(x[2161]), .Z(n10082) );
  NAND U21538 ( .A(n10083), .B(n10082), .Z(n54325) );
  NANDN U21539 ( .A(x[2158]), .B(y[2158]), .Z(n10085) );
  NANDN U21540 ( .A(x[2159]), .B(y[2159]), .Z(n10084) );
  AND U21541 ( .A(n10085), .B(n10084), .Z(n54322) );
  XNOR U21542 ( .A(x[2158]), .B(y[2158]), .Z(n54321) );
  ANDN U21543 ( .B(y[2157]), .A(x[2157]), .Z(n54320) );
  NANDN U21544 ( .A(y[2156]), .B(x[2156]), .Z(n34932) );
  ANDN U21545 ( .B(x[2157]), .A(y[2157]), .Z(n34940) );
  ANDN U21546 ( .B(n34932), .A(n34940), .Z(n54319) );
  ANDN U21547 ( .B(y[2155]), .A(x[2155]), .Z(n34927) );
  ANDN U21548 ( .B(y[2156]), .A(x[2156]), .Z(n34936) );
  OR U21549 ( .A(n34927), .B(n34936), .Z(n54318) );
  NANDN U21550 ( .A(y[2154]), .B(x[2154]), .Z(n34924) );
  NANDN U21551 ( .A(y[2155]), .B(x[2155]), .Z(n34931) );
  NAND U21552 ( .A(n34924), .B(n34931), .Z(n54316) );
  ANDN U21553 ( .B(y[2153]), .A(x[2153]), .Z(n34921) );
  ANDN U21554 ( .B(y[2154]), .A(x[2154]), .Z(n34930) );
  NOR U21555 ( .A(n34921), .B(n34930), .Z(n54315) );
  NANDN U21556 ( .A(y[2152]), .B(x[2152]), .Z(n34918) );
  NANDN U21557 ( .A(y[2153]), .B(x[2153]), .Z(n34925) );
  NAND U21558 ( .A(n34918), .B(n34925), .Z(n54314) );
  NANDN U21559 ( .A(x[2151]), .B(y[2151]), .Z(n13579) );
  ANDN U21560 ( .B(x[2150]), .A(y[2150]), .Z(n34913) );
  NANDN U21561 ( .A(y[2151]), .B(x[2151]), .Z(n54312) );
  NANDN U21562 ( .A(n34913), .B(n54312), .Z(n10086) );
  AND U21563 ( .A(n13579), .B(n10086), .Z(n13582) );
  NANDN U21564 ( .A(y[2149]), .B(x[2149]), .Z(n34914) );
  NANDN U21565 ( .A(y[2148]), .B(x[2148]), .Z(n13575) );
  NANDN U21566 ( .A(x[2147]), .B(y[2147]), .Z(n54307) );
  XNOR U21567 ( .A(x[2148]), .B(y[2148]), .Z(n27267) );
  NAND U21568 ( .A(n54307), .B(n27267), .Z(n13573) );
  ANDN U21569 ( .B(x[2146]), .A(y[2146]), .Z(n54306) );
  NANDN U21570 ( .A(x[2145]), .B(y[2145]), .Z(n34903) );
  NANDN U21571 ( .A(x[2146]), .B(y[2146]), .Z(n27268) );
  AND U21572 ( .A(n34903), .B(n27268), .Z(n52144) );
  NANDN U21573 ( .A(y[2142]), .B(x[2142]), .Z(n27272) );
  NANDN U21574 ( .A(y[2143]), .B(x[2143]), .Z(n27270) );
  NAND U21575 ( .A(n27272), .B(n27270), .Z(n54302) );
  ANDN U21576 ( .B(y[2141]), .A(x[2141]), .Z(n34892) );
  NANDN U21577 ( .A(x[2142]), .B(y[2142]), .Z(n34897) );
  NANDN U21578 ( .A(n34892), .B(n34897), .Z(n54301) );
  NANDN U21579 ( .A(y[2140]), .B(x[2140]), .Z(n10087) );
  NANDN U21580 ( .A(y[2141]), .B(x[2141]), .Z(n27271) );
  AND U21581 ( .A(n10087), .B(n27271), .Z(n54300) );
  ANDN U21582 ( .B(y[2139]), .A(x[2139]), .Z(n34885) );
  XNOR U21583 ( .A(y[2140]), .B(x[2140]), .Z(n27274) );
  NANDN U21584 ( .A(n34885), .B(n27274), .Z(n54299) );
  NANDN U21585 ( .A(y[2138]), .B(x[2138]), .Z(n34881) );
  NANDN U21586 ( .A(y[2139]), .B(x[2139]), .Z(n27273) );
  AND U21587 ( .A(n34881), .B(n27273), .Z(n54298) );
  ANDN U21588 ( .B(y[2137]), .A(x[2137]), .Z(n34876) );
  ANDN U21589 ( .B(y[2138]), .A(x[2138]), .Z(n34886) );
  OR U21590 ( .A(n34876), .B(n34886), .Z(n54297) );
  NANDN U21591 ( .A(y[2136]), .B(x[2136]), .Z(n34873) );
  NANDN U21592 ( .A(y[2137]), .B(x[2137]), .Z(n34880) );
  NAND U21593 ( .A(n34873), .B(n34880), .Z(n54296) );
  ANDN U21594 ( .B(y[2135]), .A(x[2135]), .Z(n34869) );
  ANDN U21595 ( .B(y[2136]), .A(x[2136]), .Z(n34879) );
  NOR U21596 ( .A(n34869), .B(n34879), .Z(n54295) );
  NANDN U21597 ( .A(y[2134]), .B(x[2134]), .Z(n27275) );
  NANDN U21598 ( .A(y[2135]), .B(x[2135]), .Z(n34874) );
  NAND U21599 ( .A(n27275), .B(n34874), .Z(n54294) );
  ANDN U21600 ( .B(y[2133]), .A(x[2133]), .Z(n34863) );
  ANDN U21601 ( .B(y[2134]), .A(x[2134]), .Z(n34871) );
  NOR U21602 ( .A(n34863), .B(n34871), .Z(n54293) );
  NANDN U21603 ( .A(y[2132]), .B(x[2132]), .Z(n27277) );
  NANDN U21604 ( .A(y[2133]), .B(x[2133]), .Z(n27276) );
  NAND U21605 ( .A(n27277), .B(n27276), .Z(n54292) );
  ANDN U21606 ( .B(y[2131]), .A(x[2131]), .Z(n34858) );
  ANDN U21607 ( .B(y[2132]), .A(x[2132]), .Z(n34864) );
  OR U21608 ( .A(n34858), .B(n34864), .Z(n54291) );
  NANDN U21609 ( .A(y[2130]), .B(x[2130]), .Z(n34856) );
  NANDN U21610 ( .A(y[2131]), .B(x[2131]), .Z(n27278) );
  AND U21611 ( .A(n34856), .B(n27278), .Z(n54290) );
  NANDN U21612 ( .A(x[2129]), .B(y[2129]), .Z(n34851) );
  NANDN U21613 ( .A(x[2130]), .B(y[2130]), .Z(n10088) );
  NAND U21614 ( .A(n34851), .B(n10088), .Z(n54289) );
  ANDN U21615 ( .B(x[2128]), .A(y[2128]), .Z(n34849) );
  ANDN U21616 ( .B(x[2129]), .A(y[2129]), .Z(n34853) );
  NOR U21617 ( .A(n34849), .B(n34853), .Z(n54288) );
  NANDN U21618 ( .A(y[2126]), .B(x[2126]), .Z(n34840) );
  ANDN U21619 ( .B(x[2127]), .A(y[2127]), .Z(n34846) );
  ANDN U21620 ( .B(n34840), .A(n34846), .Z(n54286) );
  ANDN U21621 ( .B(y[2125]), .A(x[2125]), .Z(n34836) );
  NANDN U21622 ( .A(x[2126]), .B(y[2126]), .Z(n34844) );
  NANDN U21623 ( .A(n34836), .B(n34844), .Z(n54285) );
  ANDN U21624 ( .B(x[2125]), .A(y[2125]), .Z(n34842) );
  NANDN U21625 ( .A(y[2124]), .B(x[2124]), .Z(n27279) );
  NANDN U21626 ( .A(n34842), .B(n27279), .Z(n54284) );
  ANDN U21627 ( .B(y[2123]), .A(x[2123]), .Z(n34830) );
  ANDN U21628 ( .B(y[2124]), .A(x[2124]), .Z(n34838) );
  NOR U21629 ( .A(n34830), .B(n34838), .Z(n54283) );
  XNOR U21630 ( .A(y[2122]), .B(x[2122]), .Z(n34826) );
  ANDN U21631 ( .B(y[2121]), .A(x[2121]), .Z(n34821) );
  ANDN U21632 ( .B(n34826), .A(n34821), .Z(n54280) );
  NANDN U21633 ( .A(y[2120]), .B(x[2120]), .Z(n34818) );
  NANDN U21634 ( .A(y[2121]), .B(x[2121]), .Z(n34825) );
  NAND U21635 ( .A(n34818), .B(n34825), .Z(n54279) );
  ANDN U21636 ( .B(y[2119]), .A(x[2119]), .Z(n34814) );
  ANDN U21637 ( .B(y[2120]), .A(x[2120]), .Z(n34824) );
  OR U21638 ( .A(n34814), .B(n34824), .Z(n54278) );
  NANDN U21639 ( .A(y[2118]), .B(x[2118]), .Z(n27281) );
  NANDN U21640 ( .A(y[2119]), .B(x[2119]), .Z(n34819) );
  AND U21641 ( .A(n27281), .B(n34819), .Z(n54277) );
  ANDN U21642 ( .B(y[2117]), .A(x[2117]), .Z(n34810) );
  ANDN U21643 ( .B(y[2118]), .A(x[2118]), .Z(n34816) );
  OR U21644 ( .A(n34810), .B(n34816), .Z(n54276) );
  NANDN U21645 ( .A(y[2116]), .B(x[2116]), .Z(n34808) );
  NANDN U21646 ( .A(y[2117]), .B(x[2117]), .Z(n27282) );
  AND U21647 ( .A(n34808), .B(n27282), .Z(n54275) );
  NANDN U21648 ( .A(x[2115]), .B(y[2115]), .Z(n10090) );
  NANDN U21649 ( .A(x[2116]), .B(y[2116]), .Z(n10089) );
  NAND U21650 ( .A(n10090), .B(n10089), .Z(n54274) );
  NANDN U21651 ( .A(y[2114]), .B(x[2114]), .Z(n10092) );
  NANDN U21652 ( .A(y[2115]), .B(x[2115]), .Z(n10091) );
  NAND U21653 ( .A(n10092), .B(n10091), .Z(n27283) );
  NANDN U21654 ( .A(x[2114]), .B(y[2114]), .Z(n10094) );
  NANDN U21655 ( .A(x[2113]), .B(y[2113]), .Z(n10093) );
  AND U21656 ( .A(n10094), .B(n10093), .Z(n27284) );
  NANDN U21657 ( .A(y[2110]), .B(x[2110]), .Z(n10096) );
  NANDN U21658 ( .A(y[2111]), .B(x[2111]), .Z(n10095) );
  NAND U21659 ( .A(n10096), .B(n10095), .Z(n34799) );
  NANDN U21660 ( .A(x[2109]), .B(y[2109]), .Z(n10097) );
  ANDN U21661 ( .B(y[2110]), .A(x[2110]), .Z(n34793) );
  ANDN U21662 ( .B(n10097), .A(n34793), .Z(n54268) );
  ANDN U21663 ( .B(y[2107]), .A(x[2107]), .Z(n34783) );
  ANDN U21664 ( .B(y[2108]), .A(x[2108]), .Z(n34792) );
  NOR U21665 ( .A(n34783), .B(n34792), .Z(n54267) );
  NANDN U21666 ( .A(y[2106]), .B(x[2106]), .Z(n34780) );
  NANDN U21667 ( .A(y[2107]), .B(x[2107]), .Z(n34787) );
  NAND U21668 ( .A(n34780), .B(n34787), .Z(n52147) );
  ANDN U21669 ( .B(y[2105]), .A(x[2105]), .Z(n34776) );
  ANDN U21670 ( .B(y[2106]), .A(x[2106]), .Z(n34786) );
  NOR U21671 ( .A(n34776), .B(n34786), .Z(n54265) );
  ANDN U21672 ( .B(y[2103]), .A(x[2103]), .Z(n34770) );
  ANDN U21673 ( .B(y[2104]), .A(x[2104]), .Z(n34778) );
  NOR U21674 ( .A(n34770), .B(n34778), .Z(n54263) );
  NANDN U21675 ( .A(y[2102]), .B(x[2102]), .Z(n34766) );
  NANDN U21676 ( .A(y[2103]), .B(x[2103]), .Z(n27287) );
  NAND U21677 ( .A(n34766), .B(n27287), .Z(n54262) );
  ANDN U21678 ( .B(y[2101]), .A(x[2101]), .Z(n34761) );
  ANDN U21679 ( .B(y[2102]), .A(x[2102]), .Z(n34771) );
  NOR U21680 ( .A(n34761), .B(n34771), .Z(n54261) );
  NANDN U21681 ( .A(y[2100]), .B(x[2100]), .Z(n34758) );
  NANDN U21682 ( .A(y[2101]), .B(x[2101]), .Z(n34765) );
  NAND U21683 ( .A(n34758), .B(n34765), .Z(n54260) );
  ANDN U21684 ( .B(y[2099]), .A(x[2099]), .Z(n34754) );
  ANDN U21685 ( .B(y[2100]), .A(x[2100]), .Z(n34764) );
  NOR U21686 ( .A(n34754), .B(n34764), .Z(n54259) );
  NANDN U21687 ( .A(y[2098]), .B(x[2098]), .Z(n27288) );
  NANDN U21688 ( .A(y[2099]), .B(x[2099]), .Z(n34759) );
  NAND U21689 ( .A(n27288), .B(n34759), .Z(n54258) );
  ANDN U21690 ( .B(y[2097]), .A(x[2097]), .Z(n34748) );
  ANDN U21691 ( .B(y[2098]), .A(x[2098]), .Z(n34756) );
  NOR U21692 ( .A(n34748), .B(n34756), .Z(n54257) );
  NANDN U21693 ( .A(y[2096]), .B(x[2096]), .Z(n34744) );
  NANDN U21694 ( .A(y[2097]), .B(x[2097]), .Z(n27289) );
  NAND U21695 ( .A(n34744), .B(n27289), .Z(n52148) );
  ANDN U21696 ( .B(y[2095]), .A(x[2095]), .Z(n34740) );
  ANDN U21697 ( .B(y[2096]), .A(x[2096]), .Z(n34749) );
  NOR U21698 ( .A(n34740), .B(n34749), .Z(n54256) );
  NANDN U21699 ( .A(x[2093]), .B(y[2093]), .Z(n34735) );
  NANDN U21700 ( .A(x[2094]), .B(y[2094]), .Z(n27290) );
  AND U21701 ( .A(n34735), .B(n27290), .Z(n13508) );
  ANDN U21702 ( .B(x[2092]), .A(y[2092]), .Z(n13506) );
  NANDN U21703 ( .A(y[2093]), .B(x[2093]), .Z(n54253) );
  ANDN U21704 ( .B(y[2092]), .A(x[2092]), .Z(n34734) );
  NANDN U21705 ( .A(y[2091]), .B(x[2091]), .Z(n27292) );
  NANDN U21706 ( .A(x[2089]), .B(y[2089]), .Z(n54245) );
  NANDN U21707 ( .A(y[2088]), .B(x[2088]), .Z(n54244) );
  NANDN U21708 ( .A(x[2088]), .B(y[2088]), .Z(n27297) );
  ANDN U21709 ( .B(y[2087]), .A(x[2087]), .Z(n34726) );
  ANDN U21710 ( .B(n27297), .A(n34726), .Z(n54241) );
  NANDN U21711 ( .A(y[2086]), .B(x[2086]), .Z(n13491) );
  NANDN U21712 ( .A(y[2085]), .B(x[2085]), .Z(n10098) );
  AND U21713 ( .A(n13491), .B(n10098), .Z(n27301) );
  NANDN U21714 ( .A(y[2084]), .B(x[2084]), .Z(n10099) );
  NAND U21715 ( .A(n27301), .B(n10099), .Z(n34720) );
  ANDN U21716 ( .B(y[2083]), .A(x[2083]), .Z(n54233) );
  ANDN U21717 ( .B(y[2081]), .A(x[2081]), .Z(n34714) );
  ANDN U21718 ( .B(y[2082]), .A(x[2082]), .Z(n34717) );
  NOR U21719 ( .A(n34714), .B(n34717), .Z(n54230) );
  NANDN U21720 ( .A(y[2080]), .B(x[2080]), .Z(n10101) );
  NANDN U21721 ( .A(y[2081]), .B(x[2081]), .Z(n10100) );
  AND U21722 ( .A(n10101), .B(n10100), .Z(n54227) );
  NANDN U21723 ( .A(x[2080]), .B(y[2080]), .Z(n10103) );
  NANDN U21724 ( .A(x[2079]), .B(y[2079]), .Z(n10102) );
  AND U21725 ( .A(n10103), .B(n10102), .Z(n54226) );
  ANDN U21726 ( .B(x[2079]), .A(y[2079]), .Z(n10106) );
  NANDN U21727 ( .A(x[2078]), .B(y[2078]), .Z(n52150) );
  OR U21728 ( .A(n10106), .B(n52150), .Z(n10104) );
  NAND U21729 ( .A(n54226), .B(n10104), .Z(n34711) );
  NANDN U21730 ( .A(y[2078]), .B(x[2078]), .Z(n10105) );
  NANDN U21731 ( .A(n10106), .B(n10105), .Z(n27303) );
  ANDN U21732 ( .B(y[2077]), .A(x[2077]), .Z(n52149) );
  NANDN U21733 ( .A(y[2076]), .B(x[2076]), .Z(n27305) );
  NANDN U21734 ( .A(y[2077]), .B(x[2077]), .Z(n27304) );
  AND U21735 ( .A(n27305), .B(n27304), .Z(n54220) );
  ANDN U21736 ( .B(y[2075]), .A(x[2075]), .Z(n34700) );
  ANDN U21737 ( .B(y[2076]), .A(x[2076]), .Z(n34706) );
  OR U21738 ( .A(n34700), .B(n34706), .Z(n54217) );
  NANDN U21739 ( .A(y[2074]), .B(x[2074]), .Z(n34696) );
  NANDN U21740 ( .A(y[2075]), .B(x[2075]), .Z(n27306) );
  AND U21741 ( .A(n34696), .B(n27306), .Z(n54216) );
  ANDN U21742 ( .B(y[2074]), .A(x[2074]), .Z(n34701) );
  NANDN U21743 ( .A(x[2073]), .B(y[2073]), .Z(n27307) );
  NANDN U21744 ( .A(n34701), .B(n27307), .Z(n54214) );
  NANDN U21745 ( .A(y[2072]), .B(x[2072]), .Z(n27309) );
  NANDN U21746 ( .A(y[2073]), .B(x[2073]), .Z(n34695) );
  AND U21747 ( .A(n27309), .B(n34695), .Z(n54211) );
  NANDN U21748 ( .A(x[2071]), .B(y[2071]), .Z(n27311) );
  NANDN U21749 ( .A(x[2072]), .B(y[2072]), .Z(n27308) );
  NAND U21750 ( .A(n27311), .B(n27308), .Z(n54210) );
  NANDN U21751 ( .A(y[2070]), .B(x[2070]), .Z(n27314) );
  NANDN U21752 ( .A(y[2071]), .B(x[2071]), .Z(n27310) );
  NAND U21753 ( .A(n27314), .B(n27310), .Z(n54209) );
  NANDN U21754 ( .A(x[2070]), .B(y[2070]), .Z(n27312) );
  ANDN U21755 ( .B(y[2069]), .A(x[2069]), .Z(n34685) );
  ANDN U21756 ( .B(n27312), .A(n34685), .Z(n54208) );
  XNOR U21757 ( .A(y[2068]), .B(x[2068]), .Z(n27316) );
  ANDN U21758 ( .B(y[2067]), .A(x[2067]), .Z(n34678) );
  ANDN U21759 ( .B(n27316), .A(n34678), .Z(n54207) );
  NANDN U21760 ( .A(y[2066]), .B(x[2066]), .Z(n34674) );
  NANDN U21761 ( .A(y[2067]), .B(x[2067]), .Z(n27315) );
  NAND U21762 ( .A(n34674), .B(n27315), .Z(n54206) );
  ANDN U21763 ( .B(y[2065]), .A(x[2065]), .Z(n27318) );
  ANDN U21764 ( .B(y[2066]), .A(x[2066]), .Z(n34679) );
  OR U21765 ( .A(n27318), .B(n34679), .Z(n54205) );
  NANDN U21766 ( .A(y[2065]), .B(x[2065]), .Z(n34673) );
  ANDN U21767 ( .B(x[2064]), .A(y[2064]), .Z(n34668) );
  ANDN U21768 ( .B(n34673), .A(n34668), .Z(n54204) );
  ANDN U21769 ( .B(x[2062]), .A(y[2062]), .Z(n34662) );
  ANDN U21770 ( .B(x[2063]), .A(y[2063]), .Z(n34669) );
  NOR U21771 ( .A(n34662), .B(n34669), .Z(n54203) );
  ANDN U21772 ( .B(y[2061]), .A(x[2061]), .Z(n10109) );
  NANDN U21773 ( .A(y[2061]), .B(x[2061]), .Z(n34663) );
  NANDN U21774 ( .A(y[2060]), .B(x[2060]), .Z(n10107) );
  NAND U21775 ( .A(n34663), .B(n10107), .Z(n10108) );
  NANDN U21776 ( .A(n10109), .B(n10108), .Z(n13463) );
  NANDN U21777 ( .A(x[2060]), .B(y[2060]), .Z(n10110) );
  ANDN U21778 ( .B(n10110), .A(n10109), .Z(n54200) );
  ANDN U21779 ( .B(x[2057]), .A(y[2057]), .Z(n34652) );
  ANDN U21780 ( .B(x[2054]), .A(y[2054]), .Z(n34642) );
  ANDN U21781 ( .B(x[2055]), .A(y[2055]), .Z(n34647) );
  NOR U21782 ( .A(n34642), .B(n34647), .Z(n54193) );
  NANDN U21783 ( .A(x[2053]), .B(y[2053]), .Z(n34638) );
  NANDN U21784 ( .A(x[2054]), .B(y[2054]), .Z(n27323) );
  NAND U21785 ( .A(n34638), .B(n27323), .Z(n54192) );
  NANDN U21786 ( .A(x[2051]), .B(y[2051]), .Z(n54188) );
  ANDN U21787 ( .B(x[2050]), .A(y[2050]), .Z(n54187) );
  NANDN U21788 ( .A(y[2051]), .B(x[2051]), .Z(n27324) );
  NANDN U21789 ( .A(x[2049]), .B(y[2049]), .Z(n34629) );
  NANDN U21790 ( .A(x[2050]), .B(y[2050]), .Z(n27326) );
  NAND U21791 ( .A(n34629), .B(n27326), .Z(n54186) );
  ANDN U21792 ( .B(x[2049]), .A(y[2049]), .Z(n34633) );
  NANDN U21793 ( .A(y[2048]), .B(x[2048]), .Z(n10111) );
  NANDN U21794 ( .A(n34633), .B(n10111), .Z(n54185) );
  NANDN U21795 ( .A(x[2047]), .B(y[2047]), .Z(n34621) );
  XOR U21796 ( .A(y[2048]), .B(x[2048]), .Z(n34627) );
  ANDN U21797 ( .B(n34621), .A(n34627), .Z(n54184) );
  ANDN U21798 ( .B(x[2046]), .A(y[2046]), .Z(n34617) );
  ANDN U21799 ( .B(x[2047]), .A(y[2047]), .Z(n34624) );
  OR U21800 ( .A(n34617), .B(n34624), .Z(n54183) );
  NANDN U21801 ( .A(x[2045]), .B(y[2045]), .Z(n27327) );
  NANDN U21802 ( .A(x[2046]), .B(y[2046]), .Z(n34622) );
  AND U21803 ( .A(n27327), .B(n34622), .Z(n54182) );
  ANDN U21804 ( .B(x[2044]), .A(y[2044]), .Z(n34611) );
  ANDN U21805 ( .B(x[2045]), .A(y[2045]), .Z(n34619) );
  OR U21806 ( .A(n34611), .B(n34619), .Z(n54181) );
  NANDN U21807 ( .A(x[2043]), .B(y[2043]), .Z(n34607) );
  NANDN U21808 ( .A(x[2044]), .B(y[2044]), .Z(n27328) );
  AND U21809 ( .A(n34607), .B(n27328), .Z(n54180) );
  ANDN U21810 ( .B(x[2043]), .A(y[2043]), .Z(n34612) );
  NANDN U21811 ( .A(y[2042]), .B(x[2042]), .Z(n27329) );
  NANDN U21812 ( .A(n34612), .B(n27329), .Z(n54179) );
  NANDN U21813 ( .A(x[2041]), .B(y[2041]), .Z(n34600) );
  NANDN U21814 ( .A(x[2042]), .B(y[2042]), .Z(n34609) );
  AND U21815 ( .A(n34600), .B(n34609), .Z(n54178) );
  NANDN U21816 ( .A(y[2040]), .B(x[2040]), .Z(n27331) );
  NANDN U21817 ( .A(y[2041]), .B(x[2041]), .Z(n27330) );
  NAND U21818 ( .A(n27331), .B(n27330), .Z(n54176) );
  NANDN U21819 ( .A(x[2039]), .B(y[2039]), .Z(n34594) );
  NANDN U21820 ( .A(x[2040]), .B(y[2040]), .Z(n34601) );
  AND U21821 ( .A(n34594), .B(n34601), .Z(n54175) );
  NANDN U21822 ( .A(y[2038]), .B(x[2038]), .Z(n34590) );
  NANDN U21823 ( .A(y[2039]), .B(x[2039]), .Z(n27332) );
  NAND U21824 ( .A(n34590), .B(n27332), .Z(n54174) );
  NANDN U21825 ( .A(x[2037]), .B(y[2037]), .Z(n34587) );
  NANDN U21826 ( .A(x[2038]), .B(y[2038]), .Z(n34595) );
  AND U21827 ( .A(n34587), .B(n34595), .Z(n52153) );
  NANDN U21828 ( .A(y[2036]), .B(x[2036]), .Z(n10112) );
  NANDN U21829 ( .A(y[2037]), .B(x[2037]), .Z(n34591) );
  NAND U21830 ( .A(n10112), .B(n34591), .Z(n54173) );
  XNOR U21831 ( .A(y[2036]), .B(x[2036]), .Z(n27333) );
  NANDN U21832 ( .A(x[2035]), .B(y[2035]), .Z(n27335) );
  AND U21833 ( .A(n27333), .B(n27335), .Z(n54172) );
  NANDN U21834 ( .A(y[2034]), .B(x[2034]), .Z(n27337) );
  NANDN U21835 ( .A(y[2035]), .B(x[2035]), .Z(n27334) );
  NAND U21836 ( .A(n27337), .B(n27334), .Z(n54171) );
  NANDN U21837 ( .A(x[2033]), .B(y[2033]), .Z(n27339) );
  NANDN U21838 ( .A(x[2034]), .B(y[2034]), .Z(n27336) );
  NAND U21839 ( .A(n27339), .B(n27336), .Z(n54170) );
  NANDN U21840 ( .A(y[2032]), .B(x[2032]), .Z(n27341) );
  NANDN U21841 ( .A(y[2033]), .B(x[2033]), .Z(n27338) );
  AND U21842 ( .A(n27341), .B(n27338), .Z(n52154) );
  ANDN U21843 ( .B(y[2031]), .A(x[2031]), .Z(n34575) );
  NANDN U21844 ( .A(x[2032]), .B(y[2032]), .Z(n27340) );
  NANDN U21845 ( .A(n34575), .B(n27340), .Z(n54169) );
  NANDN U21846 ( .A(y[2030]), .B(x[2030]), .Z(n10113) );
  NANDN U21847 ( .A(y[2031]), .B(x[2031]), .Z(n27342) );
  AND U21848 ( .A(n10113), .B(n27342), .Z(n54168) );
  ANDN U21849 ( .B(y[2029]), .A(x[2029]), .Z(n34568) );
  XNOR U21850 ( .A(y[2030]), .B(x[2030]), .Z(n34570) );
  NANDN U21851 ( .A(n34568), .B(n34570), .Z(n54167) );
  NANDN U21852 ( .A(y[2029]), .B(x[2029]), .Z(n54164) );
  ANDN U21853 ( .B(y[2027]), .A(x[2027]), .Z(n34562) );
  ANDN U21854 ( .B(y[2028]), .A(x[2028]), .Z(n54165) );
  OR U21855 ( .A(n34562), .B(n54165), .Z(n54163) );
  NANDN U21856 ( .A(y[2026]), .B(x[2026]), .Z(n54161) );
  ANDN U21857 ( .B(y[2025]), .A(x[2025]), .Z(n34556) );
  ANDN U21858 ( .B(y[2026]), .A(x[2026]), .Z(n34563) );
  OR U21859 ( .A(n34556), .B(n34563), .Z(n54160) );
  NANDN U21860 ( .A(y[2024]), .B(x[2024]), .Z(n10114) );
  NANDN U21861 ( .A(y[2025]), .B(x[2025]), .Z(n27345) );
  AND U21862 ( .A(n10114), .B(n27345), .Z(n54159) );
  ANDN U21863 ( .B(y[2023]), .A(x[2023]), .Z(n34551) );
  XNOR U21864 ( .A(y[2024]), .B(x[2024]), .Z(n34552) );
  NANDN U21865 ( .A(n34551), .B(n34552), .Z(n54158) );
  NANDN U21866 ( .A(y[2022]), .B(x[2022]), .Z(n27347) );
  NANDN U21867 ( .A(y[2023]), .B(x[2023]), .Z(n54157) );
  AND U21868 ( .A(n27347), .B(n54157), .Z(n13413) );
  ANDN U21869 ( .B(y[2021]), .A(x[2021]), .Z(n27348) );
  NANDN U21870 ( .A(x[2019]), .B(y[2019]), .Z(n27354) );
  ANDN U21871 ( .B(x[2018]), .A(y[2018]), .Z(n27356) );
  NANDN U21872 ( .A(y[2016]), .B(x[2016]), .Z(n27358) );
  NANDN U21873 ( .A(y[2017]), .B(x[2017]), .Z(n27357) );
  AND U21874 ( .A(n27358), .B(n27357), .Z(n54149) );
  ANDN U21875 ( .B(y[2015]), .A(x[2015]), .Z(n34534) );
  ANDN U21876 ( .B(y[2016]), .A(x[2016]), .Z(n34540) );
  OR U21877 ( .A(n34534), .B(n34540), .Z(n54148) );
  NANDN U21878 ( .A(y[2014]), .B(x[2014]), .Z(n34530) );
  NANDN U21879 ( .A(y[2015]), .B(x[2015]), .Z(n27359) );
  NAND U21880 ( .A(n34530), .B(n27359), .Z(n52155) );
  ANDN U21881 ( .B(y[2013]), .A(x[2013]), .Z(n34526) );
  ANDN U21882 ( .B(y[2014]), .A(x[2014]), .Z(n34535) );
  NOR U21883 ( .A(n34526), .B(n34535), .Z(n54147) );
  NANDN U21884 ( .A(x[2011]), .B(y[2011]), .Z(n34520) );
  NANDN U21885 ( .A(x[2012]), .B(y[2012]), .Z(n27360) );
  AND U21886 ( .A(n34520), .B(n27360), .Z(n13396) );
  ANDN U21887 ( .B(x[2010]), .A(y[2010]), .Z(n13394) );
  NANDN U21888 ( .A(y[2011]), .B(x[2011]), .Z(n54143) );
  NANDN U21889 ( .A(y[2008]), .B(x[2008]), .Z(n54139) );
  NANDN U21890 ( .A(y[2006]), .B(x[2006]), .Z(n34506) );
  NANDN U21891 ( .A(y[2007]), .B(x[2007]), .Z(n34514) );
  AND U21892 ( .A(n34506), .B(n34514), .Z(n54137) );
  ANDN U21893 ( .B(y[2006]), .A(x[2006]), .Z(n34512) );
  NANDN U21894 ( .A(x[2005]), .B(y[2005]), .Z(n27364) );
  NANDN U21895 ( .A(n34512), .B(n27364), .Z(n54136) );
  NANDN U21896 ( .A(x[2003]), .B(y[2003]), .Z(n34500) );
  NANDN U21897 ( .A(x[2004]), .B(y[2004]), .Z(n54135) );
  NAND U21898 ( .A(n34500), .B(n54135), .Z(n52157) );
  NANDN U21899 ( .A(y[2003]), .B(x[2003]), .Z(n27366) );
  NANDN U21900 ( .A(y[2002]), .B(x[2002]), .Z(n27367) );
  AND U21901 ( .A(n27366), .B(n27367), .Z(n13381) );
  NANDN U21902 ( .A(y[2000]), .B(x[2000]), .Z(n34490) );
  ANDN U21903 ( .B(x[2001]), .A(y[2001]), .Z(n34498) );
  ANDN U21904 ( .B(n34490), .A(n34498), .Z(n54131) );
  ANDN U21905 ( .B(y[1999]), .A(x[1999]), .Z(n34488) );
  NANDN U21906 ( .A(x[2000]), .B(y[2000]), .Z(n27369) );
  NANDN U21907 ( .A(n34488), .B(n27369), .Z(n52158) );
  NANDN U21908 ( .A(y[1998]), .B(x[1998]), .Z(n10115) );
  NANDN U21909 ( .A(y[1999]), .B(x[1999]), .Z(n34491) );
  NAND U21910 ( .A(n10115), .B(n34491), .Z(n54128) );
  XNOR U21911 ( .A(y[1998]), .B(x[1998]), .Z(n27371) );
  NANDN U21912 ( .A(x[1997]), .B(y[1997]), .Z(n27372) );
  AND U21913 ( .A(n27371), .B(n27372), .Z(n54127) );
  NANDN U21914 ( .A(y[1996]), .B(x[1996]), .Z(n27374) );
  NANDN U21915 ( .A(y[1997]), .B(x[1997]), .Z(n27370) );
  NAND U21916 ( .A(n27374), .B(n27370), .Z(n54126) );
  NANDN U21917 ( .A(y[1994]), .B(x[1994]), .Z(n27378) );
  NANDN U21918 ( .A(y[1995]), .B(x[1995]), .Z(n27375) );
  NAND U21919 ( .A(n27378), .B(n27375), .Z(n52160) );
  ANDN U21920 ( .B(y[1993]), .A(x[1993]), .Z(n27381) );
  NANDN U21921 ( .A(x[1994]), .B(y[1994]), .Z(n27377) );
  NANDN U21922 ( .A(n27381), .B(n27377), .Z(n54125) );
  NANDN U21923 ( .A(y[1993]), .B(x[1993]), .Z(n27379) );
  ANDN U21924 ( .B(x[1992]), .A(y[1992]), .Z(n34471) );
  ANDN U21925 ( .B(n27379), .A(n34471), .Z(n54124) );
  ANDN U21926 ( .B(y[1992]), .A(x[1992]), .Z(n27380) );
  NANDN U21927 ( .A(x[1991]), .B(y[1991]), .Z(n27382) );
  NANDN U21928 ( .A(n27380), .B(n27382), .Z(n54123) );
  ANDN U21929 ( .B(x[1990]), .A(y[1990]), .Z(n34465) );
  ANDN U21930 ( .B(x[1991]), .A(y[1991]), .Z(n34472) );
  NOR U21931 ( .A(n34465), .B(n34472), .Z(n54122) );
  NANDN U21932 ( .A(x[1989]), .B(y[1989]), .Z(n34461) );
  NANDN U21933 ( .A(x[1990]), .B(y[1990]), .Z(n27383) );
  NAND U21934 ( .A(n34461), .B(n27383), .Z(n52161) );
  NANDN U21935 ( .A(x[1988]), .B(y[1988]), .Z(n54120) );
  ANDN U21936 ( .B(x[1986]), .A(y[1986]), .Z(n54117) );
  NANDN U21937 ( .A(y[1982]), .B(x[1982]), .Z(n27391) );
  NANDN U21938 ( .A(y[1983]), .B(x[1983]), .Z(n27387) );
  NAND U21939 ( .A(n27391), .B(n27387), .Z(n54112) );
  NANDN U21940 ( .A(x[1981]), .B(y[1981]), .Z(n34442) );
  NANDN U21941 ( .A(x[1982]), .B(y[1982]), .Z(n27390) );
  NAND U21942 ( .A(n34442), .B(n27390), .Z(n52163) );
  NANDN U21943 ( .A(y[1980]), .B(x[1980]), .Z(n27394) );
  NANDN U21944 ( .A(y[1981]), .B(x[1981]), .Z(n27392) );
  AND U21945 ( .A(n27394), .B(n27392), .Z(n54111) );
  ANDN U21946 ( .B(y[1978]), .A(x[1978]), .Z(n54109) );
  ANDN U21947 ( .B(y[1977]), .A(x[1977]), .Z(n13348) );
  NANDN U21948 ( .A(y[1977]), .B(x[1977]), .Z(n54108) );
  NANDN U21949 ( .A(y[1976]), .B(x[1976]), .Z(n54106) );
  NAND U21950 ( .A(n54108), .B(n54106), .Z(n10116) );
  NANDN U21951 ( .A(n13348), .B(n10116), .Z(n13351) );
  XNOR U21952 ( .A(y[1970]), .B(x[1970]), .Z(n34420) );
  ANDN U21953 ( .B(y[1969]), .A(x[1969]), .Z(n34419) );
  ANDN U21954 ( .B(n34420), .A(n34419), .Z(n54101) );
  ANDN U21955 ( .B(x[1969]), .A(y[1969]), .Z(n52171) );
  NANDN U21956 ( .A(x[1968]), .B(y[1968]), .Z(n27404) );
  ANDN U21957 ( .B(y[1967]), .A(x[1967]), .Z(n34418) );
  ANDN U21958 ( .B(n27404), .A(n34418), .Z(n54100) );
  ANDN U21959 ( .B(x[1966]), .A(y[1966]), .Z(n54099) );
  XNOR U21960 ( .A(y[1966]), .B(x[1966]), .Z(n10117) );
  NANDN U21961 ( .A(x[1965]), .B(y[1965]), .Z(n27407) );
  AND U21962 ( .A(n10117), .B(n27407), .Z(n54097) );
  ANDN U21963 ( .B(x[1962]), .A(y[1962]), .Z(n34410) );
  ANDN U21964 ( .B(x[1963]), .A(y[1963]), .Z(n34416) );
  OR U21965 ( .A(n34410), .B(n34416), .Z(n54093) );
  NANDN U21966 ( .A(x[1961]), .B(y[1961]), .Z(n34407) );
  NANDN U21967 ( .A(x[1962]), .B(y[1962]), .Z(n34413) );
  NAND U21968 ( .A(n34407), .B(n34413), .Z(n52173) );
  ANDN U21969 ( .B(x[1960]), .A(y[1960]), .Z(n34403) );
  ANDN U21970 ( .B(x[1961]), .A(y[1961]), .Z(n34412) );
  NOR U21971 ( .A(n34403), .B(n34412), .Z(n54092) );
  ANDN U21972 ( .B(x[1958]), .A(y[1958]), .Z(n34397) );
  ANDN U21973 ( .B(x[1959]), .A(y[1959]), .Z(n34405) );
  NOR U21974 ( .A(n34397), .B(n34405), .Z(n54090) );
  NANDN U21975 ( .A(x[1957]), .B(y[1957]), .Z(n34393) );
  XNOR U21976 ( .A(x[1958]), .B(y[1958]), .Z(n10118) );
  NAND U21977 ( .A(n34393), .B(n10118), .Z(n54089) );
  ANDN U21978 ( .B(x[1957]), .A(y[1957]), .Z(n34398) );
  NANDN U21979 ( .A(y[1956]), .B(x[1956]), .Z(n27412) );
  NANDN U21980 ( .A(n34398), .B(n27412), .Z(n52174) );
  NANDN U21981 ( .A(x[1955]), .B(y[1955]), .Z(n27413) );
  NANDN U21982 ( .A(x[1956]), .B(y[1956]), .Z(n34392) );
  AND U21983 ( .A(n27413), .B(n34392), .Z(n54088) );
  NANDN U21984 ( .A(y[1952]), .B(x[1952]), .Z(n27417) );
  NANDN U21985 ( .A(y[1953]), .B(x[1953]), .Z(n27416) );
  NAND U21986 ( .A(n27417), .B(n27416), .Z(n54086) );
  NANDN U21987 ( .A(x[1951]), .B(y[1951]), .Z(n34376) );
  NANDN U21988 ( .A(x[1952]), .B(y[1952]), .Z(n34383) );
  NAND U21989 ( .A(n34376), .B(n34383), .Z(n52176) );
  NANDN U21990 ( .A(y[1950]), .B(x[1950]), .Z(n27419) );
  NANDN U21991 ( .A(y[1951]), .B(x[1951]), .Z(n27418) );
  AND U21992 ( .A(n27419), .B(n27418), .Z(n54083) );
  NANDN U21993 ( .A(x[1947]), .B(y[1947]), .Z(n34364) );
  NANDN U21994 ( .A(x[1948]), .B(y[1948]), .Z(n34371) );
  NAND U21995 ( .A(n34364), .B(n34371), .Z(n54081) );
  NANDN U21996 ( .A(y[1946]), .B(x[1946]), .Z(n27423) );
  NANDN U21997 ( .A(y[1947]), .B(x[1947]), .Z(n27422) );
  AND U21998 ( .A(n27423), .B(n27422), .Z(n54080) );
  NANDN U21999 ( .A(x[1945]), .B(y[1945]), .Z(n34358) );
  NANDN U22000 ( .A(x[1946]), .B(y[1946]), .Z(n34365) );
  NAND U22001 ( .A(n34358), .B(n34365), .Z(n54079) );
  NANDN U22002 ( .A(y[1944]), .B(x[1944]), .Z(n27425) );
  NANDN U22003 ( .A(y[1945]), .B(x[1945]), .Z(n27424) );
  AND U22004 ( .A(n27425), .B(n27424), .Z(n54078) );
  NANDN U22005 ( .A(x[1943]), .B(y[1943]), .Z(n34352) );
  NANDN U22006 ( .A(x[1944]), .B(y[1944]), .Z(n34359) );
  NAND U22007 ( .A(n34352), .B(n34359), .Z(n54077) );
  NANDN U22008 ( .A(x[1941]), .B(y[1941]), .Z(n27427) );
  NANDN U22009 ( .A(x[1942]), .B(y[1942]), .Z(n34353) );
  NAND U22010 ( .A(n27427), .B(n34353), .Z(n52179) );
  NANDN U22011 ( .A(y[1940]), .B(x[1940]), .Z(n34344) );
  NANDN U22012 ( .A(y[1941]), .B(x[1941]), .Z(n34349) );
  AND U22013 ( .A(n34344), .B(n34349), .Z(n54076) );
  NANDN U22014 ( .A(y[1938]), .B(x[1938]), .Z(n27431) );
  NANDN U22015 ( .A(y[1939]), .B(x[1939]), .Z(n27429) );
  AND U22016 ( .A(n27431), .B(n27429), .Z(n13304) );
  ANDN U22017 ( .B(y[1937]), .A(x[1937]), .Z(n34336) );
  NANDN U22018 ( .A(x[1935]), .B(y[1935]), .Z(n27436) );
  NANDN U22019 ( .A(y[1934]), .B(x[1934]), .Z(n54067) );
  NANDN U22020 ( .A(y[1933]), .B(x[1933]), .Z(n27437) );
  ANDN U22021 ( .B(x[1932]), .A(y[1932]), .Z(n34329) );
  ANDN U22022 ( .B(n27437), .A(n34329), .Z(n54065) );
  NANDN U22023 ( .A(x[1931]), .B(y[1931]), .Z(n34327) );
  XNOR U22024 ( .A(x[1932]), .B(y[1932]), .Z(n10119) );
  NAND U22025 ( .A(n34327), .B(n10119), .Z(n54064) );
  NANDN U22026 ( .A(y[1930]), .B(x[1930]), .Z(n10121) );
  NANDN U22027 ( .A(y[1931]), .B(x[1931]), .Z(n10120) );
  NAND U22028 ( .A(n10121), .B(n10120), .Z(n54063) );
  NANDN U22029 ( .A(x[1930]), .B(y[1930]), .Z(n10123) );
  NANDN U22030 ( .A(x[1929]), .B(y[1929]), .Z(n10122) );
  AND U22031 ( .A(n10123), .B(n10122), .Z(n54062) );
  NANDN U22032 ( .A(x[1927]), .B(y[1927]), .Z(n27444) );
  NANDN U22033 ( .A(x[1928]), .B(y[1928]), .Z(n27439) );
  AND U22034 ( .A(n27444), .B(n27439), .Z(n54060) );
  ANDN U22035 ( .B(x[1926]), .A(y[1926]), .Z(n34315) );
  ANDN U22036 ( .B(x[1927]), .A(y[1927]), .Z(n34320) );
  OR U22037 ( .A(n34315), .B(n34320), .Z(n54059) );
  NANDN U22038 ( .A(x[1925]), .B(y[1925]), .Z(n27445) );
  NANDN U22039 ( .A(x[1926]), .B(y[1926]), .Z(n27443) );
  AND U22040 ( .A(n27445), .B(n27443), .Z(n52180) );
  NANDN U22041 ( .A(x[1922]), .B(y[1922]), .Z(n54056) );
  NANDN U22042 ( .A(y[1921]), .B(x[1921]), .Z(n54054) );
  NANDN U22043 ( .A(y[1922]), .B(x[1922]), .Z(n52183) );
  NAND U22044 ( .A(n54054), .B(n52183), .Z(n34301) );
  ANDN U22045 ( .B(y[1921]), .A(x[1921]), .Z(n13276) );
  NANDN U22046 ( .A(x[1919]), .B(y[1919]), .Z(n10124) );
  AND U22047 ( .A(n34305), .B(n10124), .Z(n54053) );
  NANDN U22048 ( .A(y[1919]), .B(x[1919]), .Z(n34302) );
  ANDN U22049 ( .B(y[1917]), .A(x[1917]), .Z(n34292) );
  NANDN U22050 ( .A(x[1918]), .B(y[1918]), .Z(n27448) );
  NANDN U22051 ( .A(n34292), .B(n27448), .Z(n54051) );
  NANDN U22052 ( .A(y[1916]), .B(x[1916]), .Z(n34288) );
  NANDN U22053 ( .A(y[1917]), .B(x[1917]), .Z(n34296) );
  AND U22054 ( .A(n34288), .B(n34296), .Z(n54050) );
  ANDN U22055 ( .B(y[1915]), .A(x[1915]), .Z(n34283) );
  ANDN U22056 ( .B(y[1916]), .A(x[1916]), .Z(n34294) );
  OR U22057 ( .A(n34283), .B(n34294), .Z(n54049) );
  NANDN U22058 ( .A(y[1914]), .B(x[1914]), .Z(n34280) );
  NANDN U22059 ( .A(y[1915]), .B(x[1915]), .Z(n34287) );
  AND U22060 ( .A(n34280), .B(n34287), .Z(n54048) );
  ANDN U22061 ( .B(y[1913]), .A(x[1913]), .Z(n34276) );
  ANDN U22062 ( .B(y[1914]), .A(x[1914]), .Z(n34286) );
  OR U22063 ( .A(n34276), .B(n34286), .Z(n52184) );
  NANDN U22064 ( .A(y[1912]), .B(x[1912]), .Z(n27449) );
  NANDN U22065 ( .A(y[1913]), .B(x[1913]), .Z(n34281) );
  NAND U22066 ( .A(n27449), .B(n34281), .Z(n54047) );
  ANDN U22067 ( .B(y[1911]), .A(x[1911]), .Z(n34271) );
  ANDN U22068 ( .B(y[1912]), .A(x[1912]), .Z(n34278) );
  NOR U22069 ( .A(n34271), .B(n34278), .Z(n54046) );
  NANDN U22070 ( .A(y[1910]), .B(x[1910]), .Z(n34267) );
  NANDN U22071 ( .A(y[1911]), .B(x[1911]), .Z(n27450) );
  NAND U22072 ( .A(n34267), .B(n27450), .Z(n54045) );
  NANDN U22073 ( .A(x[1909]), .B(y[1909]), .Z(n27452) );
  ANDN U22074 ( .B(y[1910]), .A(x[1910]), .Z(n54043) );
  ANDN U22075 ( .B(n27452), .A(n54043), .Z(n13264) );
  ANDN U22076 ( .B(x[1908]), .A(y[1908]), .Z(n27453) );
  ANDN U22077 ( .B(y[1907]), .A(x[1907]), .Z(n52186) );
  NANDN U22078 ( .A(y[1907]), .B(x[1907]), .Z(n27454) );
  NANDN U22079 ( .A(x[1906]), .B(y[1906]), .Z(n10126) );
  NANDN U22080 ( .A(x[1905]), .B(y[1905]), .Z(n10125) );
  NAND U22081 ( .A(n10126), .B(n10125), .Z(n54039) );
  NANDN U22082 ( .A(y[1905]), .B(x[1905]), .Z(n10128) );
  NANDN U22083 ( .A(y[1904]), .B(x[1904]), .Z(n10127) );
  AND U22084 ( .A(n10128), .B(n10127), .Z(n54038) );
  ANDN U22085 ( .B(y[1900]), .A(x[1900]), .Z(n34255) );
  NANDN U22086 ( .A(x[1899]), .B(y[1899]), .Z(n34249) );
  NANDN U22087 ( .A(n34255), .B(n34249), .Z(n52190) );
  ANDN U22088 ( .B(x[1898]), .A(y[1898]), .Z(n34245) );
  NANDN U22089 ( .A(y[1899]), .B(x[1899]), .Z(n27455) );
  NANDN U22090 ( .A(n34245), .B(n27455), .Z(n54035) );
  NANDN U22091 ( .A(x[1897]), .B(y[1897]), .Z(n34241) );
  ANDN U22092 ( .B(y[1898]), .A(x[1898]), .Z(n34251) );
  ANDN U22093 ( .B(n34241), .A(n34251), .Z(n54034) );
  ANDN U22094 ( .B(x[1897]), .A(y[1897]), .Z(n34247) );
  NANDN U22095 ( .A(y[1896]), .B(x[1896]), .Z(n27457) );
  NANDN U22096 ( .A(n34247), .B(n27457), .Z(n54033) );
  NANDN U22097 ( .A(x[1895]), .B(y[1895]), .Z(n34235) );
  NANDN U22098 ( .A(x[1896]), .B(y[1896]), .Z(n34240) );
  AND U22099 ( .A(n34235), .B(n34240), .Z(n54032) );
  NANDN U22100 ( .A(y[1894]), .B(x[1894]), .Z(n10129) );
  NANDN U22101 ( .A(y[1895]), .B(x[1895]), .Z(n27458) );
  NAND U22102 ( .A(n10129), .B(n27458), .Z(n54031) );
  XNOR U22103 ( .A(x[1894]), .B(y[1894]), .Z(n27459) );
  ANDN U22104 ( .B(x[1892]), .A(y[1892]), .Z(n13236) );
  XNOR U22105 ( .A(x[1892]), .B(y[1892]), .Z(n27463) );
  NANDN U22106 ( .A(x[1891]), .B(y[1891]), .Z(n27464) );
  ANDN U22107 ( .B(x[1890]), .A(y[1890]), .Z(n27466) );
  NANDN U22108 ( .A(x[1889]), .B(y[1889]), .Z(n54024) );
  XNOR U22109 ( .A(y[1888]), .B(x[1888]), .Z(n27468) );
  NANDN U22110 ( .A(x[1887]), .B(y[1887]), .Z(n27470) );
  NAND U22111 ( .A(n27468), .B(n27470), .Z(n54022) );
  NANDN U22112 ( .A(y[1886]), .B(x[1886]), .Z(n27472) );
  NANDN U22113 ( .A(y[1887]), .B(x[1887]), .Z(n27469) );
  AND U22114 ( .A(n27472), .B(n27469), .Z(n52191) );
  ANDN U22115 ( .B(y[1885]), .A(x[1885]), .Z(n34218) );
  NANDN U22116 ( .A(x[1886]), .B(y[1886]), .Z(n27471) );
  NANDN U22117 ( .A(n34218), .B(n27471), .Z(n54020) );
  NANDN U22118 ( .A(y[1884]), .B(x[1884]), .Z(n27474) );
  NANDN U22119 ( .A(y[1885]), .B(x[1885]), .Z(n54019) );
  AND U22120 ( .A(n27474), .B(n54019), .Z(n13222) );
  ANDN U22121 ( .B(y[1884]), .A(x[1884]), .Z(n54018) );
  NANDN U22122 ( .A(x[1882]), .B(y[1882]), .Z(n27475) );
  ANDN U22123 ( .B(y[1881]), .A(x[1881]), .Z(n34209) );
  ANDN U22124 ( .B(n27475), .A(n34209), .Z(n54014) );
  NANDN U22125 ( .A(y[1880]), .B(x[1880]), .Z(n27478) );
  NANDN U22126 ( .A(y[1881]), .B(x[1881]), .Z(n27477) );
  NAND U22127 ( .A(n27478), .B(n27477), .Z(n52192) );
  ANDN U22128 ( .B(y[1879]), .A(x[1879]), .Z(n34203) );
  ANDN U22129 ( .B(y[1880]), .A(x[1880]), .Z(n34210) );
  OR U22130 ( .A(n34203), .B(n34210), .Z(n54013) );
  NANDN U22131 ( .A(y[1878]), .B(x[1878]), .Z(n34199) );
  NANDN U22132 ( .A(y[1879]), .B(x[1879]), .Z(n27479) );
  AND U22133 ( .A(n34199), .B(n27479), .Z(n54012) );
  NANDN U22134 ( .A(x[1875]), .B(y[1875]), .Z(n27482) );
  NANDN U22135 ( .A(x[1876]), .B(y[1876]), .Z(n27481) );
  NAND U22136 ( .A(n27482), .B(n27481), .Z(n52195) );
  NANDN U22137 ( .A(y[1874]), .B(x[1874]), .Z(n34186) );
  NANDN U22138 ( .A(y[1875]), .B(x[1875]), .Z(n34193) );
  NAND U22139 ( .A(n34186), .B(n34193), .Z(n54011) );
  NANDN U22140 ( .A(x[1873]), .B(y[1873]), .Z(n27484) );
  NANDN U22141 ( .A(x[1874]), .B(y[1874]), .Z(n27483) );
  AND U22142 ( .A(n27484), .B(n27483), .Z(n54010) );
  NANDN U22143 ( .A(y[1872]), .B(x[1872]), .Z(n34180) );
  NANDN U22144 ( .A(y[1873]), .B(x[1873]), .Z(n34187) );
  NAND U22145 ( .A(n34180), .B(n34187), .Z(n54009) );
  NANDN U22146 ( .A(x[1871]), .B(y[1871]), .Z(n34176) );
  NANDN U22147 ( .A(x[1872]), .B(y[1872]), .Z(n27485) );
  AND U22148 ( .A(n34176), .B(n27485), .Z(n54007) );
  NANDN U22149 ( .A(y[1870]), .B(x[1870]), .Z(n34173) );
  NANDN U22150 ( .A(y[1871]), .B(x[1871]), .Z(n34181) );
  NAND U22151 ( .A(n34173), .B(n34181), .Z(n54006) );
  NANDN U22152 ( .A(x[1867]), .B(y[1867]), .Z(n27490) );
  NANDN U22153 ( .A(x[1868]), .B(y[1868]), .Z(n27487) );
  NAND U22154 ( .A(n27490), .B(n27487), .Z(n54003) );
  NANDN U22155 ( .A(y[1866]), .B(x[1866]), .Z(n27492) );
  NANDN U22156 ( .A(y[1867]), .B(x[1867]), .Z(n27489) );
  AND U22157 ( .A(n27492), .B(n27489), .Z(n52196) );
  NANDN U22158 ( .A(x[1865]), .B(y[1865]), .Z(n27495) );
  NANDN U22159 ( .A(x[1866]), .B(y[1866]), .Z(n27491) );
  AND U22160 ( .A(n27495), .B(n27491), .Z(n54002) );
  NANDN U22161 ( .A(y[1864]), .B(x[1864]), .Z(n27496) );
  NANDN U22162 ( .A(y[1865]), .B(x[1865]), .Z(n27493) );
  NAND U22163 ( .A(n27496), .B(n27493), .Z(n54001) );
  NANDN U22164 ( .A(x[1863]), .B(y[1863]), .Z(n27498) );
  NANDN U22165 ( .A(x[1864]), .B(y[1864]), .Z(n27494) );
  AND U22166 ( .A(n27498), .B(n27494), .Z(n54000) );
  NANDN U22167 ( .A(y[1862]), .B(x[1862]), .Z(n34156) );
  NANDN U22168 ( .A(y[1863]), .B(x[1863]), .Z(n27497) );
  NAND U22169 ( .A(n34156), .B(n27497), .Z(n53999) );
  NANDN U22170 ( .A(x[1861]), .B(y[1861]), .Z(n27499) );
  NANDN U22171 ( .A(x[1862]), .B(y[1862]), .Z(n53998) );
  AND U22172 ( .A(n27499), .B(n53998), .Z(n13196) );
  ANDN U22173 ( .B(x[1860]), .A(y[1860]), .Z(n13193) );
  XNOR U22174 ( .A(x[1860]), .B(y[1860]), .Z(n27502) );
  NANDN U22175 ( .A(x[1859]), .B(y[1859]), .Z(n27503) );
  AND U22176 ( .A(n27502), .B(n27503), .Z(n13191) );
  NANDN U22177 ( .A(y[1858]), .B(x[1858]), .Z(n27506) );
  NANDN U22178 ( .A(x[1858]), .B(y[1858]), .Z(n27504) );
  ANDN U22179 ( .B(x[1857]), .A(y[1857]), .Z(n27505) );
  ANDN U22180 ( .B(x[1855]), .A(y[1855]), .Z(n10130) );
  NAND U22181 ( .A(n10130), .B(x[1856]), .Z(n10133) );
  XOR U22182 ( .A(n10130), .B(x[1856]), .Z(n10131) );
  NANDN U22183 ( .A(y[1856]), .B(n10131), .Z(n10132) );
  NAND U22184 ( .A(n10133), .B(n10132), .Z(n53991) );
  NOR U22185 ( .A(n27505), .B(n53991), .Z(n13185) );
  NANDN U22186 ( .A(y[1852]), .B(x[1852]), .Z(n34142) );
  NANDN U22187 ( .A(x[1851]), .B(y[1851]), .Z(n27508) );
  XNOR U22188 ( .A(y[1851]), .B(x[1851]), .Z(n13170) );
  NANDN U22189 ( .A(y[1848]), .B(x[1848]), .Z(n34131) );
  NANDN U22190 ( .A(y[1849]), .B(x[1849]), .Z(n34138) );
  AND U22191 ( .A(n34131), .B(n34138), .Z(n53984) );
  ANDN U22192 ( .B(y[1847]), .A(x[1847]), .Z(n27510) );
  ANDN U22193 ( .B(y[1848]), .A(x[1848]), .Z(n34136) );
  OR U22194 ( .A(n27510), .B(n34136), .Z(n53983) );
  NANDN U22195 ( .A(y[1847]), .B(x[1847]), .Z(n34130) );
  ANDN U22196 ( .B(x[1846]), .A(y[1846]), .Z(n34125) );
  ANDN U22197 ( .B(n34130), .A(n34125), .Z(n53982) );
  NANDN U22198 ( .A(x[1845]), .B(y[1845]), .Z(n27511) );
  XNOR U22199 ( .A(x[1846]), .B(y[1846]), .Z(n10134) );
  NAND U22200 ( .A(n27511), .B(n10134), .Z(n53981) );
  ANDN U22201 ( .B(x[1844]), .A(y[1844]), .Z(n34120) );
  ANDN U22202 ( .B(x[1845]), .A(y[1845]), .Z(n34126) );
  NOR U22203 ( .A(n34120), .B(n34126), .Z(n53980) );
  NANDN U22204 ( .A(x[1843]), .B(y[1843]), .Z(n34118) );
  NANDN U22205 ( .A(x[1844]), .B(y[1844]), .Z(n27512) );
  NAND U22206 ( .A(n34118), .B(n27512), .Z(n53979) );
  NANDN U22207 ( .A(y[1842]), .B(x[1842]), .Z(n10135) );
  ANDN U22208 ( .B(x[1843]), .A(y[1843]), .Z(n53978) );
  ANDN U22209 ( .B(n10135), .A(n53978), .Z(n13159) );
  ANDN U22210 ( .B(y[1841]), .A(x[1841]), .Z(n53974) );
  ANDN U22211 ( .B(y[1839]), .A(x[1839]), .Z(n34104) );
  ANDN U22212 ( .B(y[1840]), .A(x[1840]), .Z(n34113) );
  NOR U22213 ( .A(n34104), .B(n34113), .Z(n53972) );
  ANDN U22214 ( .B(y[1837]), .A(x[1837]), .Z(n34099) );
  ANDN U22215 ( .B(y[1838]), .A(x[1838]), .Z(n34107) );
  NOR U22216 ( .A(n34099), .B(n34107), .Z(n53970) );
  ANDN U22217 ( .B(x[1836]), .A(y[1836]), .Z(n27515) );
  NANDN U22218 ( .A(y[1834]), .B(x[1834]), .Z(n53965) );
  NANDN U22219 ( .A(x[1833]), .B(y[1833]), .Z(n34090) );
  NANDN U22220 ( .A(x[1834]), .B(y[1834]), .Z(n27517) );
  AND U22221 ( .A(n34090), .B(n27517), .Z(n53964) );
  NANDN U22222 ( .A(y[1832]), .B(x[1832]), .Z(n10136) );
  NANDN U22223 ( .A(y[1833]), .B(x[1833]), .Z(n27518) );
  NAND U22224 ( .A(n10136), .B(n27518), .Z(n53963) );
  NANDN U22225 ( .A(x[1831]), .B(y[1831]), .Z(n34082) );
  XOR U22226 ( .A(y[1832]), .B(x[1832]), .Z(n34086) );
  ANDN U22227 ( .B(n34082), .A(n34086), .Z(n53962) );
  ANDN U22228 ( .B(x[1830]), .A(y[1830]), .Z(n34077) );
  ANDN U22229 ( .B(x[1831]), .A(y[1831]), .Z(n34088) );
  OR U22230 ( .A(n34077), .B(n34088), .Z(n53961) );
  NANDN U22231 ( .A(x[1829]), .B(y[1829]), .Z(n34074) );
  NANDN U22232 ( .A(x[1830]), .B(y[1830]), .Z(n34084) );
  AND U22233 ( .A(n34074), .B(n34084), .Z(n53960) );
  ANDN U22234 ( .B(x[1828]), .A(y[1828]), .Z(n34070) );
  ANDN U22235 ( .B(x[1829]), .A(y[1829]), .Z(n34080) );
  OR U22236 ( .A(n34070), .B(n34080), .Z(n53959) );
  NANDN U22237 ( .A(x[1827]), .B(y[1827]), .Z(n27519) );
  NANDN U22238 ( .A(x[1828]), .B(y[1828]), .Z(n34075) );
  AND U22239 ( .A(n27519), .B(n34075), .Z(n53958) );
  ANDN U22240 ( .B(x[1826]), .A(y[1826]), .Z(n34064) );
  ANDN U22241 ( .B(x[1827]), .A(y[1827]), .Z(n34072) );
  OR U22242 ( .A(n34064), .B(n34072), .Z(n53957) );
  NANDN U22243 ( .A(x[1825]), .B(y[1825]), .Z(n34060) );
  NANDN U22244 ( .A(x[1826]), .B(y[1826]), .Z(n27520) );
  AND U22245 ( .A(n34060), .B(n27520), .Z(n53955) );
  ANDN U22246 ( .B(x[1825]), .A(y[1825]), .Z(n34065) );
  NANDN U22247 ( .A(y[1824]), .B(x[1824]), .Z(n27521) );
  NANDN U22248 ( .A(n34065), .B(n27521), .Z(n53954) );
  NANDN U22249 ( .A(x[1823]), .B(y[1823]), .Z(n27523) );
  NANDN U22250 ( .A(x[1824]), .B(y[1824]), .Z(n53953) );
  AND U22251 ( .A(n27523), .B(n53953), .Z(n13134) );
  ANDN U22252 ( .B(x[1822]), .A(y[1822]), .Z(n27524) );
  ANDN U22253 ( .B(y[1821]), .A(x[1821]), .Z(n27526) );
  NANDN U22254 ( .A(y[1821]), .B(x[1821]), .Z(n27525) );
  NANDN U22255 ( .A(x[1820]), .B(y[1820]), .Z(n27528) );
  NANDN U22256 ( .A(x[1819]), .B(y[1819]), .Z(n34052) );
  AND U22257 ( .A(n27528), .B(n34052), .Z(n13126) );
  NANDN U22258 ( .A(y[1818]), .B(x[1818]), .Z(n53947) );
  ANDN U22259 ( .B(y[1815]), .A(x[1815]), .Z(n34039) );
  ANDN U22260 ( .B(y[1816]), .A(x[1816]), .Z(n34046) );
  OR U22261 ( .A(n34039), .B(n34046), .Z(n52202) );
  NANDN U22262 ( .A(y[1814]), .B(x[1814]), .Z(n34035) );
  NANDN U22263 ( .A(y[1815]), .B(x[1815]), .Z(n34044) );
  NAND U22264 ( .A(n34035), .B(n34044), .Z(n53946) );
  NANDN U22265 ( .A(x[1813]), .B(y[1813]), .Z(n27533) );
  ANDN U22266 ( .B(y[1814]), .A(x[1814]), .Z(n34041) );
  ANDN U22267 ( .B(n27533), .A(n34041), .Z(n53945) );
  NANDN U22268 ( .A(y[1812]), .B(x[1812]), .Z(n27535) );
  NANDN U22269 ( .A(y[1813]), .B(x[1813]), .Z(n34034) );
  NAND U22270 ( .A(n27535), .B(n34034), .Z(n53944) );
  NANDN U22271 ( .A(x[1811]), .B(y[1811]), .Z(n27537) );
  NANDN U22272 ( .A(x[1812]), .B(y[1812]), .Z(n27534) );
  AND U22273 ( .A(n27537), .B(n27534), .Z(n53942) );
  NANDN U22274 ( .A(y[1810]), .B(x[1810]), .Z(n27538) );
  NANDN U22275 ( .A(y[1811]), .B(x[1811]), .Z(n27536) );
  NAND U22276 ( .A(n27538), .B(n27536), .Z(n53941) );
  NANDN U22277 ( .A(x[1809]), .B(y[1809]), .Z(n27540) );
  ANDN U22278 ( .B(x[1808]), .A(y[1808]), .Z(n13111) );
  ANDN U22279 ( .B(y[1807]), .A(x[1807]), .Z(n27542) );
  NANDN U22280 ( .A(y[1807]), .B(x[1807]), .Z(n27541) );
  XOR U22281 ( .A(x[1806]), .B(y[1806]), .Z(n27545) );
  NANDN U22282 ( .A(x[1803]), .B(y[1803]), .Z(n34015) );
  NANDN U22283 ( .A(x[1804]), .B(y[1804]), .Z(n27549) );
  NAND U22284 ( .A(n34015), .B(n27549), .Z(n53932) );
  ANDN U22285 ( .B(x[1802]), .A(y[1802]), .Z(n34013) );
  ANDN U22286 ( .B(x[1803]), .A(y[1803]), .Z(n34017) );
  NOR U22287 ( .A(n34013), .B(n34017), .Z(n53931) );
  NANDN U22288 ( .A(x[1801]), .B(y[1801]), .Z(n10138) );
  NANDN U22289 ( .A(x[1802]), .B(y[1802]), .Z(n10137) );
  NAND U22290 ( .A(n10138), .B(n10137), .Z(n34010) );
  NANDN U22291 ( .A(y[1800]), .B(x[1800]), .Z(n52203) );
  ANDN U22292 ( .B(x[1801]), .A(y[1801]), .Z(n53929) );
  ANDN U22293 ( .B(n52203), .A(n53929), .Z(n34008) );
  NANDN U22294 ( .A(x[1800]), .B(y[1800]), .Z(n53928) );
  NANDN U22295 ( .A(x[1799]), .B(y[1799]), .Z(n53925) );
  AND U22296 ( .A(n53928), .B(n53925), .Z(n34007) );
  NANDN U22297 ( .A(y[1798]), .B(x[1798]), .Z(n53924) );
  NANDN U22298 ( .A(y[1799]), .B(x[1799]), .Z(n53927) );
  NAND U22299 ( .A(n53924), .B(n53927), .Z(n34005) );
  NANDN U22300 ( .A(x[1798]), .B(y[1798]), .Z(n10140) );
  NANDN U22301 ( .A(x[1797]), .B(y[1797]), .Z(n10139) );
  AND U22302 ( .A(n10140), .B(n10139), .Z(n53923) );
  NANDN U22303 ( .A(x[1795]), .B(y[1795]), .Z(n27554) );
  NANDN U22304 ( .A(x[1796]), .B(y[1796]), .Z(n27550) );
  AND U22305 ( .A(n27554), .B(n27550), .Z(n53921) );
  ANDN U22306 ( .B(x[1794]), .A(y[1794]), .Z(n33997) );
  NANDN U22307 ( .A(y[1795]), .B(x[1795]), .Z(n27553) );
  NANDN U22308 ( .A(n33997), .B(n27553), .Z(n53920) );
  NANDN U22309 ( .A(x[1793]), .B(y[1793]), .Z(n33995) );
  NANDN U22310 ( .A(x[1794]), .B(y[1794]), .Z(n27555) );
  AND U22311 ( .A(n33995), .B(n27555), .Z(n52204) );
  NANDN U22312 ( .A(y[1792]), .B(x[1792]), .Z(n10142) );
  NANDN U22313 ( .A(y[1793]), .B(x[1793]), .Z(n10141) );
  NAND U22314 ( .A(n10142), .B(n10141), .Z(n52205) );
  NANDN U22315 ( .A(x[1791]), .B(y[1791]), .Z(n10144) );
  ANDN U22316 ( .B(y[1792]), .A(x[1792]), .Z(n10143) );
  ANDN U22317 ( .B(n10144), .A(n10143), .Z(n53919) );
  NANDN U22318 ( .A(y[1790]), .B(x[1790]), .Z(n33989) );
  NANDN U22319 ( .A(y[1791]), .B(x[1791]), .Z(n10145) );
  AND U22320 ( .A(n33989), .B(n10145), .Z(n52206) );
  NANDN U22321 ( .A(x[1789]), .B(y[1789]), .Z(n10147) );
  NANDN U22322 ( .A(x[1790]), .B(y[1790]), .Z(n10146) );
  NAND U22323 ( .A(n10147), .B(n10146), .Z(n52207) );
  NANDN U22324 ( .A(y[1789]), .B(x[1789]), .Z(n10149) );
  NANDN U22325 ( .A(y[1788]), .B(x[1788]), .Z(n10148) );
  AND U22326 ( .A(n10149), .B(n10148), .Z(n53918) );
  ANDN U22327 ( .B(y[1786]), .A(x[1786]), .Z(n33983) );
  NANDN U22328 ( .A(x[1785]), .B(y[1785]), .Z(n27556) );
  NANDN U22329 ( .A(n33983), .B(n27556), .Z(n53912) );
  NANDN U22330 ( .A(y[1785]), .B(x[1785]), .Z(n33981) );
  NANDN U22331 ( .A(y[1784]), .B(x[1784]), .Z(n27559) );
  AND U22332 ( .A(n33981), .B(n27559), .Z(n52208) );
  ANDN U22333 ( .B(y[1783]), .A(x[1783]), .Z(n33973) );
  NANDN U22334 ( .A(x[1784]), .B(y[1784]), .Z(n27557) );
  NANDN U22335 ( .A(n33973), .B(n27557), .Z(n53911) );
  NANDN U22336 ( .A(y[1782]), .B(x[1782]), .Z(n10150) );
  NANDN U22337 ( .A(y[1783]), .B(x[1783]), .Z(n27558) );
  AND U22338 ( .A(n10150), .B(n27558), .Z(n53910) );
  XNOR U22339 ( .A(y[1782]), .B(x[1782]), .Z(n10151) );
  NANDN U22340 ( .A(x[1781]), .B(y[1781]), .Z(n27560) );
  NAND U22341 ( .A(n10151), .B(n27560), .Z(n53909) );
  ANDN U22342 ( .B(x[1780]), .A(y[1780]), .Z(n33970) );
  ANDN U22343 ( .B(x[1781]), .A(y[1781]), .Z(n33972) );
  NOR U22344 ( .A(n33970), .B(n33972), .Z(n53908) );
  NANDN U22345 ( .A(x[1779]), .B(y[1779]), .Z(n33969) );
  NANDN U22346 ( .A(x[1780]), .B(y[1780]), .Z(n27561) );
  NAND U22347 ( .A(n33969), .B(n27561), .Z(n53907) );
  ANDN U22348 ( .B(x[1778]), .A(y[1778]), .Z(n27563) );
  ANDN U22349 ( .B(x[1779]), .A(y[1779]), .Z(n33971) );
  NOR U22350 ( .A(n27563), .B(n33971), .Z(n53906) );
  ANDN U22351 ( .B(y[1777]), .A(x[1777]), .Z(n33967) );
  NANDN U22352 ( .A(x[1778]), .B(y[1778]), .Z(n33968) );
  NANDN U22353 ( .A(n33967), .B(n33968), .Z(n53905) );
  NANDN U22354 ( .A(y[1777]), .B(x[1777]), .Z(n27562) );
  ANDN U22355 ( .B(y[1776]), .A(x[1776]), .Z(n53903) );
  NANDN U22356 ( .A(x[1775]), .B(y[1775]), .Z(n53901) );
  NANDN U22357 ( .A(n53903), .B(n53901), .Z(n13065) );
  NANDN U22358 ( .A(x[1773]), .B(y[1773]), .Z(n33963) );
  NANDN U22359 ( .A(x[1774]), .B(y[1774]), .Z(n27566) );
  AND U22360 ( .A(n33963), .B(n27566), .Z(n53899) );
  ANDN U22361 ( .B(x[1772]), .A(y[1772]), .Z(n33960) );
  NANDN U22362 ( .A(y[1773]), .B(x[1773]), .Z(n27567) );
  NANDN U22363 ( .A(n33960), .B(n27567), .Z(n53898) );
  NANDN U22364 ( .A(x[1771]), .B(y[1771]), .Z(n27568) );
  ANDN U22365 ( .B(y[1772]), .A(x[1772]), .Z(n33965) );
  ANDN U22366 ( .B(n27568), .A(n33965), .Z(n53897) );
  ANDN U22367 ( .B(x[1771]), .A(y[1771]), .Z(n52209) );
  NANDN U22368 ( .A(x[1769]), .B(y[1769]), .Z(n33951) );
  ANDN U22369 ( .B(x[1769]), .A(y[1769]), .Z(n33954) );
  NANDN U22370 ( .A(x[1768]), .B(y[1768]), .Z(n33952) );
  NANDN U22371 ( .A(y[1767]), .B(x[1767]), .Z(n10153) );
  NANDN U22372 ( .A(y[1768]), .B(x[1768]), .Z(n10152) );
  NAND U22373 ( .A(n10153), .B(n10152), .Z(n53893) );
  NANDN U22374 ( .A(x[1767]), .B(y[1767]), .Z(n53892) );
  NANDN U22375 ( .A(x[1766]), .B(y[1766]), .Z(n52211) );
  AND U22376 ( .A(n53892), .B(n52211), .Z(n33949) );
  ANDN U22377 ( .B(x[1766]), .A(y[1766]), .Z(n53891) );
  NANDN U22378 ( .A(x[1765]), .B(y[1765]), .Z(n52212) );
  NANDN U22379 ( .A(y[1764]), .B(x[1764]), .Z(n27569) );
  ANDN U22380 ( .B(x[1765]), .A(y[1765]), .Z(n33946) );
  ANDN U22381 ( .B(n27569), .A(n33946), .Z(n53890) );
  NANDN U22382 ( .A(x[1763]), .B(y[1763]), .Z(n27571) );
  NANDN U22383 ( .A(x[1764]), .B(y[1764]), .Z(n33942) );
  NAND U22384 ( .A(n27571), .B(n33942), .Z(n53889) );
  NANDN U22385 ( .A(y[1762]), .B(x[1762]), .Z(n27573) );
  NANDN U22386 ( .A(y[1763]), .B(x[1763]), .Z(n27570) );
  AND U22387 ( .A(n27573), .B(n27570), .Z(n53888) );
  NANDN U22388 ( .A(x[1761]), .B(y[1761]), .Z(n27576) );
  NANDN U22389 ( .A(x[1762]), .B(y[1762]), .Z(n27572) );
  NAND U22390 ( .A(n27576), .B(n27572), .Z(n53887) );
  NANDN U22391 ( .A(y[1761]), .B(x[1761]), .Z(n27574) );
  ANDN U22392 ( .B(x[1760]), .A(y[1760]), .Z(n33931) );
  ANDN U22393 ( .B(n27574), .A(n33931), .Z(n53886) );
  NANDN U22394 ( .A(x[1759]), .B(y[1759]), .Z(n27577) );
  NANDN U22395 ( .A(x[1760]), .B(y[1760]), .Z(n27575) );
  NAND U22396 ( .A(n27577), .B(n27575), .Z(n53885) );
  ANDN U22397 ( .B(x[1756]), .A(y[1756]), .Z(n53879) );
  XNOR U22398 ( .A(y[1756]), .B(x[1756]), .Z(n27580) );
  NANDN U22399 ( .A(x[1755]), .B(y[1755]), .Z(n27582) );
  AND U22400 ( .A(n27580), .B(n27582), .Z(n53878) );
  NANDN U22401 ( .A(y[1754]), .B(x[1754]), .Z(n27585) );
  NANDN U22402 ( .A(y[1755]), .B(x[1755]), .Z(n27581) );
  NAND U22403 ( .A(n27585), .B(n27581), .Z(n53877) );
  NANDN U22404 ( .A(x[1753]), .B(y[1753]), .Z(n27586) );
  NANDN U22405 ( .A(x[1754]), .B(y[1754]), .Z(n27583) );
  AND U22406 ( .A(n27586), .B(n27583), .Z(n53876) );
  NANDN U22407 ( .A(y[1751]), .B(x[1751]), .Z(n10155) );
  NANDN U22408 ( .A(y[1750]), .B(x[1750]), .Z(n10154) );
  AND U22409 ( .A(n10155), .B(n10154), .Z(n10156) );
  NANDN U22410 ( .A(y[1752]), .B(x[1752]), .Z(n13031) );
  NAND U22411 ( .A(n10156), .B(n13031), .Z(n33914) );
  NANDN U22412 ( .A(y[1748]), .B(x[1748]), .Z(n10157) );
  ANDN U22413 ( .B(x[1749]), .A(y[1749]), .Z(n13022) );
  ANDN U22414 ( .B(n10157), .A(n13022), .Z(n53872) );
  ANDN U22415 ( .B(y[1747]), .A(x[1747]), .Z(n53871) );
  NANDN U22416 ( .A(y[1746]), .B(x[1746]), .Z(n33905) );
  NANDN U22417 ( .A(y[1747]), .B(x[1747]), .Z(n33910) );
  NAND U22418 ( .A(n33905), .B(n33910), .Z(n53869) );
  ANDN U22419 ( .B(y[1745]), .A(x[1745]), .Z(n33903) );
  ANDN U22420 ( .B(y[1746]), .A(x[1746]), .Z(n33908) );
  NOR U22421 ( .A(n33903), .B(n33908), .Z(n53868) );
  NANDN U22422 ( .A(y[1745]), .B(x[1745]), .Z(n10159) );
  NANDN U22423 ( .A(y[1744]), .B(x[1744]), .Z(n10158) );
  AND U22424 ( .A(n10159), .B(n10158), .Z(n52214) );
  NANDN U22425 ( .A(x[1743]), .B(y[1743]), .Z(n10161) );
  NANDN U22426 ( .A(x[1744]), .B(y[1744]), .Z(n10160) );
  NAND U22427 ( .A(n10161), .B(n10160), .Z(n52215) );
  NANDN U22428 ( .A(y[1743]), .B(x[1743]), .Z(n10163) );
  NANDN U22429 ( .A(y[1742]), .B(x[1742]), .Z(n10162) );
  AND U22430 ( .A(n10163), .B(n10162), .Z(n53865) );
  ANDN U22431 ( .B(y[1738]), .A(x[1738]), .Z(n52219) );
  NANDN U22432 ( .A(x[1737]), .B(y[1737]), .Z(n33888) );
  NANDN U22433 ( .A(y[1737]), .B(x[1737]), .Z(n53863) );
  NANDN U22434 ( .A(x[1736]), .B(y[1736]), .Z(n33889) );
  ANDN U22435 ( .B(x[1734]), .A(y[1734]), .Z(n27592) );
  NANDN U22436 ( .A(x[1731]), .B(y[1731]), .Z(n27596) );
  ANDN U22437 ( .B(y[1732]), .A(x[1732]), .Z(n27595) );
  ANDN U22438 ( .B(n27596), .A(n27595), .Z(n53855) );
  ANDN U22439 ( .B(x[1730]), .A(y[1730]), .Z(n33873) );
  ANDN U22440 ( .B(x[1731]), .A(y[1731]), .Z(n33880) );
  OR U22441 ( .A(n33873), .B(n33880), .Z(n53854) );
  NANDN U22442 ( .A(x[1729]), .B(y[1729]), .Z(n33870) );
  NANDN U22443 ( .A(x[1730]), .B(y[1730]), .Z(n27597) );
  AND U22444 ( .A(n33870), .B(n27597), .Z(n53853) );
  ANDN U22445 ( .B(x[1729]), .A(y[1729]), .Z(n33874) );
  NANDN U22446 ( .A(y[1728]), .B(x[1728]), .Z(n10164) );
  NANDN U22447 ( .A(n33874), .B(n10164), .Z(n53852) );
  ANDN U22448 ( .B(y[1727]), .A(x[1727]), .Z(n53850) );
  ANDN U22449 ( .B(x[1727]), .A(y[1727]), .Z(n27599) );
  NANDN U22450 ( .A(y[1726]), .B(x[1726]), .Z(n33862) );
  NANDN U22451 ( .A(n27599), .B(n33862), .Z(n53849) );
  ANDN U22452 ( .B(y[1726]), .A(x[1726]), .Z(n53848) );
  NANDN U22453 ( .A(y[1723]), .B(x[1723]), .Z(n10166) );
  NANDN U22454 ( .A(y[1724]), .B(x[1724]), .Z(n10165) );
  NAND U22455 ( .A(n10166), .B(n10165), .Z(n27603) );
  NANDN U22456 ( .A(x[1723]), .B(y[1723]), .Z(n12979) );
  NANDN U22457 ( .A(x[1722]), .B(y[1722]), .Z(n10167) );
  AND U22458 ( .A(n12979), .B(n10167), .Z(n27602) );
  NANDN U22459 ( .A(x[1721]), .B(y[1721]), .Z(n10168) );
  AND U22460 ( .A(n27602), .B(n10168), .Z(n27604) );
  ANDN U22461 ( .B(x[1720]), .A(y[1720]), .Z(n27605) );
  ANDN U22462 ( .B(y[1719]), .A(x[1719]), .Z(n33852) );
  ANDN U22463 ( .B(y[1720]), .A(x[1720]), .Z(n33858) );
  NOR U22464 ( .A(n33852), .B(n33858), .Z(n53842) );
  NANDN U22465 ( .A(y[1718]), .B(x[1718]), .Z(n10169) );
  NANDN U22466 ( .A(y[1719]), .B(x[1719]), .Z(n27606) );
  NAND U22467 ( .A(n10169), .B(n27606), .Z(n53840) );
  XNOR U22468 ( .A(y[1718]), .B(x[1718]), .Z(n33848) );
  NANDN U22469 ( .A(x[1717]), .B(y[1717]), .Z(n27607) );
  AND U22470 ( .A(n33848), .B(n27607), .Z(n53839) );
  NANDN U22471 ( .A(x[1715]), .B(y[1715]), .Z(n27610) );
  NANDN U22472 ( .A(x[1716]), .B(y[1716]), .Z(n52221) );
  NAND U22473 ( .A(n27610), .B(n52221), .Z(n12969) );
  NANDN U22474 ( .A(x[1713]), .B(y[1713]), .Z(n27611) );
  ANDN U22475 ( .B(y[1714]), .A(x[1714]), .Z(n33843) );
  ANDN U22476 ( .B(n27611), .A(n33843), .Z(n53835) );
  NANDN U22477 ( .A(y[1712]), .B(x[1712]), .Z(n33833) );
  NANDN U22478 ( .A(y[1713]), .B(x[1713]), .Z(n33840) );
  NAND U22479 ( .A(n33833), .B(n33840), .Z(n52222) );
  NANDN U22480 ( .A(x[1711]), .B(y[1711]), .Z(n27614) );
  NANDN U22481 ( .A(x[1712]), .B(y[1712]), .Z(n27612) );
  NAND U22482 ( .A(n27614), .B(n27612), .Z(n53834) );
  NANDN U22483 ( .A(y[1710]), .B(x[1710]), .Z(n33828) );
  NANDN U22484 ( .A(y[1711]), .B(x[1711]), .Z(n33834) );
  AND U22485 ( .A(n33828), .B(n33834), .Z(n53833) );
  NANDN U22486 ( .A(y[1708]), .B(x[1708]), .Z(n33820) );
  ANDN U22487 ( .B(x[1709]), .A(y[1709]), .Z(n33830) );
  ANDN U22488 ( .B(n33820), .A(n33830), .Z(n53832) );
  ANDN U22489 ( .B(y[1708]), .A(x[1708]), .Z(n33826) );
  NANDN U22490 ( .A(x[1707]), .B(y[1707]), .Z(n27615) );
  NANDN U22491 ( .A(n33826), .B(n27615), .Z(n52224) );
  NANDN U22492 ( .A(y[1706]), .B(x[1706]), .Z(n33816) );
  NANDN U22493 ( .A(y[1707]), .B(x[1707]), .Z(n33819) );
  AND U22494 ( .A(n33816), .B(n33819), .Z(n53829) );
  NANDN U22495 ( .A(x[1705]), .B(y[1705]), .Z(n27617) );
  NANDN U22496 ( .A(x[1706]), .B(y[1706]), .Z(n27616) );
  NAND U22497 ( .A(n27617), .B(n27616), .Z(n53828) );
  NANDN U22498 ( .A(y[1704]), .B(x[1704]), .Z(n33807) );
  ANDN U22499 ( .B(x[1705]), .A(y[1705]), .Z(n33814) );
  ANDN U22500 ( .B(n33807), .A(n33814), .Z(n53827) );
  NANDN U22501 ( .A(x[1701]), .B(y[1701]), .Z(n27621) );
  NANDN U22502 ( .A(x[1702]), .B(y[1702]), .Z(n27620) );
  NAND U22503 ( .A(n27621), .B(n27620), .Z(n52227) );
  NANDN U22504 ( .A(y[1700]), .B(x[1700]), .Z(n33795) );
  NANDN U22505 ( .A(y[1701]), .B(x[1701]), .Z(n33802) );
  AND U22506 ( .A(n33795), .B(n33802), .Z(n53826) );
  NANDN U22507 ( .A(x[1699]), .B(y[1699]), .Z(n27623) );
  NANDN U22508 ( .A(x[1700]), .B(y[1700]), .Z(n27622) );
  NAND U22509 ( .A(n27623), .B(n27622), .Z(n53825) );
  NANDN U22510 ( .A(y[1698]), .B(x[1698]), .Z(n33789) );
  NANDN U22511 ( .A(y[1699]), .B(x[1699]), .Z(n33796) );
  AND U22512 ( .A(n33789), .B(n33796), .Z(n52228) );
  NANDN U22513 ( .A(x[1695]), .B(y[1695]), .Z(n27627) );
  NANDN U22514 ( .A(x[1696]), .B(y[1696]), .Z(n27626) );
  NAND U22515 ( .A(n27627), .B(n27626), .Z(n52231) );
  NANDN U22516 ( .A(x[1693]), .B(y[1693]), .Z(n27629) );
  NANDN U22517 ( .A(x[1694]), .B(y[1694]), .Z(n27628) );
  AND U22518 ( .A(n27629), .B(n27628), .Z(n53821) );
  NANDN U22519 ( .A(y[1693]), .B(x[1693]), .Z(n53820) );
  NANDN U22520 ( .A(x[1691]), .B(y[1691]), .Z(n27633) );
  ANDN U22521 ( .B(x[1690]), .A(y[1690]), .Z(n27634) );
  NANDN U22522 ( .A(x[1690]), .B(y[1690]), .Z(n27632) );
  ANDN U22523 ( .B(x[1689]), .A(y[1689]), .Z(n27635) );
  NANDN U22524 ( .A(y[1687]), .B(x[1687]), .Z(n33769) );
  NANDN U22525 ( .A(y[1686]), .B(x[1686]), .Z(n27639) );
  AND U22526 ( .A(n33769), .B(n27639), .Z(n12933) );
  ANDN U22527 ( .B(y[1685]), .A(x[1685]), .Z(n27641) );
  NANDN U22528 ( .A(x[1686]), .B(y[1686]), .Z(n53814) );
  ANDN U22529 ( .B(x[1684]), .A(y[1684]), .Z(n53811) );
  NANDN U22530 ( .A(x[1683]), .B(y[1683]), .Z(n27642) );
  NANDN U22531 ( .A(x[1684]), .B(y[1684]), .Z(n33764) );
  AND U22532 ( .A(n27642), .B(n33764), .Z(n53810) );
  ANDN U22533 ( .B(x[1683]), .A(y[1683]), .Z(n33762) );
  NANDN U22534 ( .A(y[1682]), .B(x[1682]), .Z(n33754) );
  NANDN U22535 ( .A(n33762), .B(n33754), .Z(n53809) );
  NANDN U22536 ( .A(x[1682]), .B(y[1682]), .Z(n27643) );
  ANDN U22537 ( .B(y[1681]), .A(x[1681]), .Z(n33752) );
  ANDN U22538 ( .B(n27643), .A(n33752), .Z(n53808) );
  NANDN U22539 ( .A(y[1680]), .B(x[1680]), .Z(n10170) );
  NANDN U22540 ( .A(y[1681]), .B(x[1681]), .Z(n33755) );
  NAND U22541 ( .A(n10170), .B(n33755), .Z(n53806) );
  XNOR U22542 ( .A(y[1680]), .B(x[1680]), .Z(n27645) );
  ANDN U22543 ( .B(y[1679]), .A(x[1679]), .Z(n33744) );
  ANDN U22544 ( .B(n27645), .A(n33744), .Z(n53805) );
  NANDN U22545 ( .A(y[1678]), .B(x[1678]), .Z(n33741) );
  NANDN U22546 ( .A(y[1679]), .B(x[1679]), .Z(n27644) );
  NAND U22547 ( .A(n33741), .B(n27644), .Z(n53804) );
  ANDN U22548 ( .B(y[1677]), .A(x[1677]), .Z(n33738) );
  ANDN U22549 ( .B(y[1678]), .A(x[1678]), .Z(n33747) );
  NOR U22550 ( .A(n33738), .B(n33747), .Z(n53803) );
  NANDN U22551 ( .A(y[1676]), .B(x[1676]), .Z(n27646) );
  NANDN U22552 ( .A(y[1677]), .B(x[1677]), .Z(n33742) );
  NAND U22553 ( .A(n27646), .B(n33742), .Z(n53802) );
  NANDN U22554 ( .A(x[1675]), .B(y[1675]), .Z(n33733) );
  ANDN U22555 ( .B(y[1676]), .A(x[1676]), .Z(n53801) );
  ANDN U22556 ( .B(n33733), .A(n53801), .Z(n12919) );
  NANDN U22557 ( .A(y[1675]), .B(x[1675]), .Z(n53800) );
  NANDN U22558 ( .A(x[1674]), .B(y[1674]), .Z(n33732) );
  NANDN U22559 ( .A(y[1672]), .B(x[1672]), .Z(n53797) );
  ANDN U22560 ( .B(y[1672]), .A(x[1672]), .Z(n27650) );
  NANDN U22561 ( .A(x[1671]), .B(y[1671]), .Z(n10171) );
  NANDN U22562 ( .A(n27650), .B(n10171), .Z(n33725) );
  IV U22563 ( .A(n33725), .Z(n53796) );
  NANDN U22564 ( .A(y[1670]), .B(x[1670]), .Z(n27652) );
  NANDN U22565 ( .A(y[1671]), .B(x[1671]), .Z(n27649) );
  NAND U22566 ( .A(n27652), .B(n27649), .Z(n53795) );
  NANDN U22567 ( .A(x[1669]), .B(y[1669]), .Z(n33718) );
  ANDN U22568 ( .B(y[1670]), .A(x[1670]), .Z(n33727) );
  ANDN U22569 ( .B(n33718), .A(n33727), .Z(n53794) );
  NANDN U22570 ( .A(y[1668]), .B(x[1668]), .Z(n27655) );
  NANDN U22571 ( .A(y[1669]), .B(x[1669]), .Z(n27653) );
  NAND U22572 ( .A(n27655), .B(n27653), .Z(n53793) );
  NANDN U22573 ( .A(x[1668]), .B(y[1668]), .Z(n33719) );
  ANDN U22574 ( .B(y[1667]), .A(x[1667]), .Z(n33713) );
  ANDN U22575 ( .B(n33719), .A(n33713), .Z(n53792) );
  NANDN U22576 ( .A(y[1666]), .B(x[1666]), .Z(n27656) );
  NANDN U22577 ( .A(y[1667]), .B(x[1667]), .Z(n27654) );
  NAND U22578 ( .A(n27656), .B(n27654), .Z(n53791) );
  ANDN U22579 ( .B(y[1665]), .A(x[1665]), .Z(n33708) );
  ANDN U22580 ( .B(y[1666]), .A(x[1666]), .Z(n33714) );
  NOR U22581 ( .A(n33708), .B(n33714), .Z(n53790) );
  NANDN U22582 ( .A(y[1664]), .B(x[1664]), .Z(n33704) );
  NANDN U22583 ( .A(y[1665]), .B(x[1665]), .Z(n27657) );
  NAND U22584 ( .A(n33704), .B(n27657), .Z(n53788) );
  ANDN U22585 ( .B(y[1664]), .A(x[1664]), .Z(n53783) );
  NANDN U22586 ( .A(x[1659]), .B(y[1659]), .Z(n27660) );
  ANDN U22587 ( .B(y[1660]), .A(x[1660]), .Z(n33698) );
  ANDN U22588 ( .B(n27660), .A(n33698), .Z(n53774) );
  NANDN U22589 ( .A(y[1658]), .B(x[1658]), .Z(n27661) );
  NANDN U22590 ( .A(y[1659]), .B(x[1659]), .Z(n33693) );
  NAND U22591 ( .A(n27661), .B(n33693), .Z(n53772) );
  NANDN U22592 ( .A(x[1657]), .B(y[1657]), .Z(n27663) );
  NANDN U22593 ( .A(x[1658]), .B(y[1658]), .Z(n27659) );
  AND U22594 ( .A(n27663), .B(n27659), .Z(n53770) );
  NANDN U22595 ( .A(y[1656]), .B(x[1656]), .Z(n27665) );
  NANDN U22596 ( .A(y[1657]), .B(x[1657]), .Z(n27662) );
  NAND U22597 ( .A(n27665), .B(n27662), .Z(n53768) );
  NANDN U22598 ( .A(x[1655]), .B(y[1655]), .Z(n27667) );
  NANDN U22599 ( .A(x[1656]), .B(y[1656]), .Z(n27664) );
  AND U22600 ( .A(n27667), .B(n27664), .Z(n53766) );
  NANDN U22601 ( .A(y[1654]), .B(x[1654]), .Z(n10172) );
  NANDN U22602 ( .A(y[1655]), .B(x[1655]), .Z(n27666) );
  NAND U22603 ( .A(n10172), .B(n27666), .Z(n53764) );
  XNOR U22604 ( .A(y[1654]), .B(x[1654]), .Z(n27670) );
  NANDN U22605 ( .A(x[1653]), .B(y[1653]), .Z(n27671) );
  AND U22606 ( .A(n27670), .B(n27671), .Z(n53762) );
  NANDN U22607 ( .A(y[1652]), .B(x[1652]), .Z(n33675) );
  NANDN U22608 ( .A(y[1653]), .B(x[1653]), .Z(n27669) );
  NAND U22609 ( .A(n33675), .B(n27669), .Z(n53760) );
  NANDN U22610 ( .A(x[1651]), .B(y[1651]), .Z(n27673) );
  NANDN U22611 ( .A(x[1652]), .B(y[1652]), .Z(n27672) );
  AND U22612 ( .A(n27673), .B(n27672), .Z(n53758) );
  NANDN U22613 ( .A(y[1650]), .B(x[1650]), .Z(n33671) );
  NANDN U22614 ( .A(y[1651]), .B(x[1651]), .Z(n33676) );
  NAND U22615 ( .A(n33671), .B(n33676), .Z(n53756) );
  NANDN U22616 ( .A(x[1650]), .B(y[1650]), .Z(n53754) );
  ANDN U22617 ( .B(x[1649]), .A(y[1649]), .Z(n53752) );
  NANDN U22618 ( .A(y[1644]), .B(x[1644]), .Z(n27677) );
  NANDN U22619 ( .A(y[1645]), .B(x[1645]), .Z(n33661) );
  NAND U22620 ( .A(n27677), .B(n33661), .Z(n52240) );
  NANDN U22621 ( .A(x[1643]), .B(y[1643]), .Z(n27678) );
  NANDN U22622 ( .A(x[1644]), .B(y[1644]), .Z(n27675) );
  AND U22623 ( .A(n27678), .B(n27675), .Z(n53749) );
  NANDN U22624 ( .A(y[1642]), .B(x[1642]), .Z(n27680) );
  NANDN U22625 ( .A(y[1643]), .B(x[1643]), .Z(n27676) );
  NAND U22626 ( .A(n27680), .B(n27676), .Z(n53748) );
  NANDN U22627 ( .A(x[1642]), .B(y[1642]), .Z(n52241) );
  ANDN U22628 ( .B(x[1640]), .A(y[1640]), .Z(n27683) );
  NANDN U22629 ( .A(x[1639]), .B(y[1639]), .Z(n27686) );
  ANDN U22630 ( .B(x[1638]), .A(y[1638]), .Z(n33647) );
  NANDN U22631 ( .A(x[1638]), .B(y[1638]), .Z(n27685) );
  ANDN U22632 ( .B(x[1636]), .A(y[1636]), .Z(n52244) );
  NANDN U22633 ( .A(x[1636]), .B(y[1636]), .Z(n27687) );
  ANDN U22634 ( .B(y[1635]), .A(x[1635]), .Z(n33639) );
  ANDN U22635 ( .B(n27687), .A(n33639), .Z(n53742) );
  NANDN U22636 ( .A(y[1634]), .B(x[1634]), .Z(n10173) );
  NANDN U22637 ( .A(y[1635]), .B(x[1635]), .Z(n33643) );
  NAND U22638 ( .A(n10173), .B(n33643), .Z(n52245) );
  XNOR U22639 ( .A(y[1634]), .B(x[1634]), .Z(n33635) );
  NANDN U22640 ( .A(x[1633]), .B(y[1633]), .Z(n27688) );
  AND U22641 ( .A(n33635), .B(n27688), .Z(n53741) );
  ANDN U22642 ( .B(x[1632]), .A(y[1632]), .Z(n27690) );
  NANDN U22643 ( .A(y[1633]), .B(x[1633]), .Z(n53738) );
  NANDN U22644 ( .A(y[1631]), .B(x[1631]), .Z(n27691) );
  NANDN U22645 ( .A(y[1630]), .B(x[1630]), .Z(n53736) );
  AND U22646 ( .A(n27691), .B(n53736), .Z(n12853) );
  ANDN U22647 ( .B(y[1629]), .A(x[1629]), .Z(n33624) );
  ANDN U22648 ( .B(y[1630]), .A(x[1630]), .Z(n33630) );
  NOR U22649 ( .A(n33624), .B(n33630), .Z(n53735) );
  NANDN U22650 ( .A(y[1628]), .B(x[1628]), .Z(n10174) );
  NANDN U22651 ( .A(y[1629]), .B(x[1629]), .Z(n33625) );
  NAND U22652 ( .A(n10174), .B(n33625), .Z(n53734) );
  XNOR U22653 ( .A(y[1628]), .B(x[1628]), .Z(n33618) );
  ANDN U22654 ( .B(y[1627]), .A(x[1627]), .Z(n33614) );
  ANDN U22655 ( .B(n33618), .A(n33614), .Z(n53733) );
  NANDN U22656 ( .A(y[1626]), .B(x[1626]), .Z(n27692) );
  NANDN U22657 ( .A(y[1627]), .B(x[1627]), .Z(n33619) );
  NAND U22658 ( .A(n27692), .B(n33619), .Z(n53732) );
  ANDN U22659 ( .B(y[1625]), .A(x[1625]), .Z(n33608) );
  ANDN U22660 ( .B(y[1626]), .A(x[1626]), .Z(n33616) );
  NOR U22661 ( .A(n33608), .B(n33616), .Z(n53731) );
  NANDN U22662 ( .A(y[1624]), .B(x[1624]), .Z(n33604) );
  NANDN U22663 ( .A(y[1625]), .B(x[1625]), .Z(n27693) );
  NAND U22664 ( .A(n33604), .B(n27693), .Z(n53730) );
  ANDN U22665 ( .B(y[1623]), .A(x[1623]), .Z(n33599) );
  ANDN U22666 ( .B(y[1624]), .A(x[1624]), .Z(n33609) );
  NOR U22667 ( .A(n33599), .B(n33609), .Z(n53728) );
  NANDN U22668 ( .A(y[1622]), .B(x[1622]), .Z(n33596) );
  NANDN U22669 ( .A(y[1623]), .B(x[1623]), .Z(n33603) );
  NAND U22670 ( .A(n33596), .B(n33603), .Z(n53727) );
  ANDN U22671 ( .B(y[1621]), .A(x[1621]), .Z(n33592) );
  ANDN U22672 ( .B(y[1622]), .A(x[1622]), .Z(n33602) );
  NOR U22673 ( .A(n33592), .B(n33602), .Z(n53726) );
  NANDN U22674 ( .A(y[1620]), .B(x[1620]), .Z(n27694) );
  NANDN U22675 ( .A(y[1621]), .B(x[1621]), .Z(n33597) );
  NAND U22676 ( .A(n27694), .B(n33597), .Z(n53725) );
  ANDN U22677 ( .B(y[1619]), .A(x[1619]), .Z(n33586) );
  ANDN U22678 ( .B(y[1620]), .A(x[1620]), .Z(n33594) );
  NOR U22679 ( .A(n33586), .B(n33594), .Z(n53724) );
  NANDN U22680 ( .A(y[1618]), .B(x[1618]), .Z(n33582) );
  NANDN U22681 ( .A(y[1619]), .B(x[1619]), .Z(n27695) );
  NAND U22682 ( .A(n33582), .B(n27695), .Z(n53723) );
  ANDN U22683 ( .B(y[1617]), .A(x[1617]), .Z(n33577) );
  ANDN U22684 ( .B(y[1618]), .A(x[1618]), .Z(n33587) );
  NOR U22685 ( .A(n33577), .B(n33587), .Z(n53722) );
  NANDN U22686 ( .A(y[1616]), .B(x[1616]), .Z(n33574) );
  NANDN U22687 ( .A(y[1617]), .B(x[1617]), .Z(n33581) );
  NAND U22688 ( .A(n33574), .B(n33581), .Z(n53721) );
  ANDN U22689 ( .B(y[1615]), .A(x[1615]), .Z(n33570) );
  ANDN U22690 ( .B(y[1616]), .A(x[1616]), .Z(n33580) );
  NOR U22691 ( .A(n33570), .B(n33580), .Z(n53720) );
  NANDN U22692 ( .A(y[1614]), .B(x[1614]), .Z(n27696) );
  NANDN U22693 ( .A(y[1615]), .B(x[1615]), .Z(n33575) );
  NAND U22694 ( .A(n27696), .B(n33575), .Z(n53719) );
  ANDN U22695 ( .B(y[1613]), .A(x[1613]), .Z(n33564) );
  ANDN U22696 ( .B(y[1614]), .A(x[1614]), .Z(n33572) );
  NOR U22697 ( .A(n33564), .B(n33572), .Z(n53718) );
  NANDN U22698 ( .A(y[1612]), .B(x[1612]), .Z(n33560) );
  NANDN U22699 ( .A(y[1613]), .B(x[1613]), .Z(n27697) );
  NAND U22700 ( .A(n33560), .B(n27697), .Z(n53717) );
  ANDN U22701 ( .B(y[1611]), .A(x[1611]), .Z(n33556) );
  ANDN U22702 ( .B(y[1612]), .A(x[1612]), .Z(n33565) );
  NOR U22703 ( .A(n33556), .B(n33565), .Z(n53716) );
  NANDN U22704 ( .A(y[1610]), .B(x[1610]), .Z(n33554) );
  NANDN U22705 ( .A(y[1611]), .B(x[1611]), .Z(n33559) );
  NAND U22706 ( .A(n33554), .B(n33559), .Z(n53715) );
  ANDN U22707 ( .B(y[1610]), .A(x[1610]), .Z(n53714) );
  NANDN U22708 ( .A(y[1609]), .B(x[1609]), .Z(n53713) );
  ANDN U22709 ( .B(y[1607]), .A(x[1607]), .Z(n53710) );
  XNOR U22710 ( .A(x[1608]), .B(y[1608]), .Z(n27699) );
  NANDN U22711 ( .A(y[1606]), .B(x[1606]), .Z(n53708) );
  ANDN U22712 ( .B(y[1605]), .A(x[1605]), .Z(n33540) );
  ANDN U22713 ( .B(y[1606]), .A(x[1606]), .Z(n33546) );
  NOR U22714 ( .A(n33540), .B(n33546), .Z(n53707) );
  NANDN U22715 ( .A(y[1604]), .B(x[1604]), .Z(n33536) );
  NANDN U22716 ( .A(y[1605]), .B(x[1605]), .Z(n33544) );
  NAND U22717 ( .A(n33536), .B(n33544), .Z(n53706) );
  ANDN U22718 ( .B(y[1603]), .A(x[1603]), .Z(n33535) );
  ANDN U22719 ( .B(y[1604]), .A(x[1604]), .Z(n33542) );
  NOR U22720 ( .A(n33535), .B(n33542), .Z(n53705) );
  NANDN U22721 ( .A(y[1603]), .B(x[1603]), .Z(n53704) );
  NANDN U22722 ( .A(x[1601]), .B(y[1601]), .Z(n27703) );
  NANDN U22723 ( .A(y[1601]), .B(x[1601]), .Z(n27701) );
  NANDN U22724 ( .A(y[1600]), .B(x[1600]), .Z(n27706) );
  AND U22725 ( .A(n27701), .B(n27706), .Z(n12815) );
  ANDN U22726 ( .B(y[1600]), .A(x[1600]), .Z(n27702) );
  NANDN U22727 ( .A(x[1599]), .B(y[1599]), .Z(n33528) );
  NANDN U22728 ( .A(y[1598]), .B(x[1598]), .Z(n53699) );
  NANDN U22729 ( .A(x[1598]), .B(y[1598]), .Z(n33527) );
  NANDN U22730 ( .A(y[1596]), .B(x[1596]), .Z(n27708) );
  NANDN U22731 ( .A(y[1597]), .B(x[1597]), .Z(n27707) );
  NAND U22732 ( .A(n27708), .B(n27707), .Z(n53697) );
  ANDN U22733 ( .B(y[1595]), .A(x[1595]), .Z(n33519) );
  ANDN U22734 ( .B(y[1596]), .A(x[1596]), .Z(n33523) );
  NOR U22735 ( .A(n33519), .B(n33523), .Z(n53696) );
  NANDN U22736 ( .A(y[1594]), .B(x[1594]), .Z(n33517) );
  NANDN U22737 ( .A(y[1595]), .B(x[1595]), .Z(n27709) );
  NAND U22738 ( .A(n33517), .B(n27709), .Z(n53695) );
  NANDN U22739 ( .A(y[1592]), .B(x[1592]), .Z(n10176) );
  NANDN U22740 ( .A(y[1593]), .B(x[1593]), .Z(n10175) );
  NAND U22741 ( .A(n10176), .B(n10175), .Z(n33513) );
  NANDN U22742 ( .A(x[1592]), .B(y[1592]), .Z(n10178) );
  NANDN U22743 ( .A(x[1591]), .B(y[1591]), .Z(n10177) );
  AND U22744 ( .A(n10178), .B(n10177), .Z(n53691) );
  NANDN U22745 ( .A(y[1591]), .B(x[1591]), .Z(n53690) );
  NANDN U22746 ( .A(y[1590]), .B(x[1590]), .Z(n53687) );
  NAND U22747 ( .A(n53690), .B(n53687), .Z(n33510) );
  NANDN U22748 ( .A(x[1590]), .B(y[1590]), .Z(n53688) );
  NANDN U22749 ( .A(x[1589]), .B(y[1589]), .Z(n52248) );
  AND U22750 ( .A(n53688), .B(n52248), .Z(n33509) );
  NANDN U22751 ( .A(x[1588]), .B(y[1588]), .Z(n33506) );
  ANDN U22752 ( .B(y[1587]), .A(x[1587]), .Z(n33498) );
  ANDN U22753 ( .B(n33506), .A(n33498), .Z(n53685) );
  NANDN U22754 ( .A(y[1586]), .B(x[1586]), .Z(n33494) );
  NANDN U22755 ( .A(y[1587]), .B(x[1587]), .Z(n33502) );
  NAND U22756 ( .A(n33494), .B(n33502), .Z(n52249) );
  ANDN U22757 ( .B(y[1585]), .A(x[1585]), .Z(n27714) );
  ANDN U22758 ( .B(y[1586]), .A(x[1586]), .Z(n33500) );
  OR U22759 ( .A(n27714), .B(n33500), .Z(n53684) );
  NANDN U22760 ( .A(y[1585]), .B(x[1585]), .Z(n53681) );
  NANDN U22761 ( .A(y[1584]), .B(x[1584]), .Z(n10181) );
  NANDN U22762 ( .A(x[1583]), .B(y[1583]), .Z(n10179) );
  ANDN U22763 ( .B(y[1584]), .A(x[1584]), .Z(n53682) );
  ANDN U22764 ( .B(n10179), .A(n53682), .Z(n53680) );
  ANDN U22765 ( .B(n10181), .A(n53680), .Z(n27711) );
  NANDN U22766 ( .A(y[1583]), .B(x[1583]), .Z(n10180) );
  AND U22767 ( .A(n10181), .B(n10180), .Z(n53683) );
  NANDN U22768 ( .A(y[1582]), .B(x[1582]), .Z(n53679) );
  AND U22769 ( .A(n53683), .B(n53679), .Z(n33489) );
  ANDN U22770 ( .B(y[1581]), .A(x[1581]), .Z(n27716) );
  ANDN U22771 ( .B(y[1582]), .A(x[1582]), .Z(n27710) );
  NOR U22772 ( .A(n27716), .B(n27710), .Z(n53678) );
  ANDN U22773 ( .B(x[1580]), .A(y[1580]), .Z(n33483) );
  NANDN U22774 ( .A(y[1581]), .B(x[1581]), .Z(n33488) );
  NANDN U22775 ( .A(n33483), .B(n33488), .Z(n53677) );
  NANDN U22776 ( .A(x[1579]), .B(y[1579]), .Z(n27717) );
  ANDN U22777 ( .B(y[1580]), .A(x[1580]), .Z(n27715) );
  ANDN U22778 ( .B(n27717), .A(n27715), .Z(n53676) );
  ANDN U22779 ( .B(x[1578]), .A(y[1578]), .Z(n33477) );
  ANDN U22780 ( .B(x[1579]), .A(y[1579]), .Z(n33484) );
  OR U22781 ( .A(n33477), .B(n33484), .Z(n53675) );
  NANDN U22782 ( .A(x[1577]), .B(y[1577]), .Z(n33473) );
  NANDN U22783 ( .A(x[1578]), .B(y[1578]), .Z(n27718) );
  AND U22784 ( .A(n33473), .B(n27718), .Z(n53673) );
  ANDN U22785 ( .B(x[1577]), .A(y[1577]), .Z(n33478) );
  NANDN U22786 ( .A(y[1576]), .B(x[1576]), .Z(n10182) );
  NANDN U22787 ( .A(n33478), .B(n10182), .Z(n53671) );
  XNOR U22788 ( .A(y[1576]), .B(x[1576]), .Z(n27720) );
  NANDN U22789 ( .A(x[1575]), .B(y[1575]), .Z(n27721) );
  AND U22790 ( .A(n27720), .B(n27721), .Z(n53669) );
  NANDN U22791 ( .A(y[1574]), .B(x[1574]), .Z(n27723) );
  NANDN U22792 ( .A(y[1575]), .B(x[1575]), .Z(n27719) );
  NAND U22793 ( .A(n27723), .B(n27719), .Z(n53667) );
  NANDN U22794 ( .A(x[1573]), .B(y[1573]), .Z(n27726) );
  NANDN U22795 ( .A(x[1574]), .B(y[1574]), .Z(n27722) );
  AND U22796 ( .A(n27726), .B(n27722), .Z(n53665) );
  ANDN U22797 ( .B(x[1572]), .A(y[1572]), .Z(n33461) );
  NANDN U22798 ( .A(y[1573]), .B(x[1573]), .Z(n27724) );
  NANDN U22799 ( .A(n33461), .B(n27724), .Z(n53663) );
  NANDN U22800 ( .A(x[1571]), .B(y[1571]), .Z(n27727) );
  NANDN U22801 ( .A(x[1572]), .B(y[1572]), .Z(n27725) );
  AND U22802 ( .A(n27727), .B(n27725), .Z(n53661) );
  ANDN U22803 ( .B(x[1570]), .A(y[1570]), .Z(n33455) );
  ANDN U22804 ( .B(x[1571]), .A(y[1571]), .Z(n33462) );
  OR U22805 ( .A(n33455), .B(n33462), .Z(n53659) );
  NANDN U22806 ( .A(x[1569]), .B(y[1569]), .Z(n33451) );
  NANDN U22807 ( .A(x[1570]), .B(y[1570]), .Z(n27728) );
  AND U22808 ( .A(n33451), .B(n27728), .Z(n53657) );
  ANDN U22809 ( .B(x[1569]), .A(y[1569]), .Z(n33456) );
  NANDN U22810 ( .A(y[1568]), .B(x[1568]), .Z(n27729) );
  NANDN U22811 ( .A(n33456), .B(n27729), .Z(n53655) );
  NANDN U22812 ( .A(x[1567]), .B(y[1567]), .Z(n27730) );
  NANDN U22813 ( .A(x[1568]), .B(y[1568]), .Z(n53653) );
  AND U22814 ( .A(n27730), .B(n53653), .Z(n12775) );
  NANDN U22815 ( .A(y[1567]), .B(x[1567]), .Z(n53650) );
  NANDN U22816 ( .A(x[1566]), .B(y[1566]), .Z(n27731) );
  ANDN U22817 ( .B(x[1565]), .A(y[1565]), .Z(n33446) );
  NANDN U22818 ( .A(y[1564]), .B(x[1564]), .Z(n10183) );
  NANDN U22819 ( .A(n33446), .B(n10183), .Z(n53642) );
  XOR U22820 ( .A(y[1564]), .B(x[1564]), .Z(n27732) );
  ANDN U22821 ( .B(y[1563]), .A(x[1563]), .Z(n33437) );
  NOR U22822 ( .A(n27732), .B(n33437), .Z(n53641) );
  ANDN U22823 ( .B(x[1563]), .A(y[1563]), .Z(n27733) );
  NANDN U22824 ( .A(y[1562]), .B(x[1562]), .Z(n27734) );
  NANDN U22825 ( .A(n27733), .B(n27734), .Z(n53639) );
  ANDN U22826 ( .B(y[1561]), .A(x[1561]), .Z(n33432) );
  ANDN U22827 ( .B(y[1562]), .A(x[1562]), .Z(n33438) );
  NOR U22828 ( .A(n33432), .B(n33438), .Z(n53637) );
  NANDN U22829 ( .A(y[1560]), .B(x[1560]), .Z(n33429) );
  NANDN U22830 ( .A(y[1561]), .B(x[1561]), .Z(n27735) );
  NAND U22831 ( .A(n33429), .B(n27735), .Z(n53635) );
  ANDN U22832 ( .B(y[1560]), .A(x[1560]), .Z(n53633) );
  NANDN U22833 ( .A(y[1559]), .B(x[1559]), .Z(n52250) );
  NANDN U22834 ( .A(x[1558]), .B(y[1558]), .Z(n53631) );
  NANDN U22835 ( .A(x[1559]), .B(y[1559]), .Z(n53632) );
  AND U22836 ( .A(n53631), .B(n53632), .Z(n33427) );
  ANDN U22837 ( .B(x[1556]), .A(y[1556]), .Z(n27738) );
  ANDN U22838 ( .B(y[1555]), .A(x[1555]), .Z(n33420) );
  NANDN U22839 ( .A(y[1555]), .B(x[1555]), .Z(n27739) );
  ANDN U22840 ( .B(y[1553]), .A(x[1553]), .Z(n52253) );
  NANDN U22841 ( .A(x[1549]), .B(y[1549]), .Z(n27744) );
  NANDN U22842 ( .A(x[1550]), .B(y[1550]), .Z(n27741) );
  NAND U22843 ( .A(n27744), .B(n27741), .Z(n53624) );
  NANDN U22844 ( .A(y[1548]), .B(x[1548]), .Z(n27745) );
  NANDN U22845 ( .A(y[1549]), .B(x[1549]), .Z(n27743) );
  AND U22846 ( .A(n27745), .B(n27743), .Z(n53620) );
  NANDN U22847 ( .A(x[1548]), .B(y[1548]), .Z(n53621) );
  NANDN U22848 ( .A(x[1547]), .B(y[1547]), .Z(n33399) );
  NAND U22849 ( .A(n53621), .B(n33399), .Z(n53619) );
  NANDN U22850 ( .A(x[1545]), .B(y[1545]), .Z(n33392) );
  ANDN U22851 ( .B(y[1546]), .A(x[1546]), .Z(n33401) );
  ANDN U22852 ( .B(n33392), .A(n33401), .Z(n53618) );
  ANDN U22853 ( .B(x[1545]), .A(y[1545]), .Z(n33397) );
  NANDN U22854 ( .A(y[1544]), .B(x[1544]), .Z(n27747) );
  NANDN U22855 ( .A(n33397), .B(n27747), .Z(n52256) );
  NANDN U22856 ( .A(x[1543]), .B(y[1543]), .Z(n27748) );
  NANDN U22857 ( .A(x[1544]), .B(y[1544]), .Z(n33391) );
  NAND U22858 ( .A(n27748), .B(n33391), .Z(n53617) );
  NANDN U22859 ( .A(y[1542]), .B(x[1542]), .Z(n33383) );
  NANDN U22860 ( .A(y[1543]), .B(x[1543]), .Z(n27746) );
  AND U22861 ( .A(n33383), .B(n27746), .Z(n53616) );
  NANDN U22862 ( .A(x[1541]), .B(y[1541]), .Z(n33380) );
  NANDN U22863 ( .A(x[1542]), .B(y[1542]), .Z(n27749) );
  NAND U22864 ( .A(n33380), .B(n27749), .Z(n53615) );
  NANDN U22865 ( .A(y[1540]), .B(x[1540]), .Z(n27750) );
  NANDN U22866 ( .A(y[1541]), .B(x[1541]), .Z(n33384) );
  AND U22867 ( .A(n27750), .B(n33384), .Z(n53614) );
  NANDN U22868 ( .A(x[1539]), .B(y[1539]), .Z(n27752) );
  NANDN U22869 ( .A(x[1540]), .B(y[1540]), .Z(n33382) );
  NAND U22870 ( .A(n27752), .B(n33382), .Z(n53613) );
  NANDN U22871 ( .A(y[1538]), .B(x[1538]), .Z(n27754) );
  NANDN U22872 ( .A(y[1539]), .B(x[1539]), .Z(n27751) );
  AND U22873 ( .A(n27754), .B(n27751), .Z(n53612) );
  NANDN U22874 ( .A(x[1537]), .B(y[1537]), .Z(n27757) );
  NANDN U22875 ( .A(x[1538]), .B(y[1538]), .Z(n27753) );
  NAND U22876 ( .A(n27757), .B(n27753), .Z(n53611) );
  NANDN U22877 ( .A(y[1537]), .B(x[1537]), .Z(n27755) );
  ANDN U22878 ( .B(x[1536]), .A(y[1536]), .Z(n33370) );
  ANDN U22879 ( .B(n27755), .A(n33370), .Z(n53610) );
  NANDN U22880 ( .A(x[1535]), .B(y[1535]), .Z(n33368) );
  XNOR U22881 ( .A(y[1536]), .B(x[1536]), .Z(n10184) );
  NAND U22882 ( .A(n33368), .B(n10184), .Z(n53609) );
  NANDN U22883 ( .A(x[1533]), .B(y[1533]), .Z(n10186) );
  NANDN U22884 ( .A(x[1534]), .B(y[1534]), .Z(n10185) );
  AND U22885 ( .A(n10186), .B(n10185), .Z(n53607) );
  NANDN U22886 ( .A(y[1532]), .B(x[1532]), .Z(n10187) );
  ANDN U22887 ( .B(x[1533]), .A(y[1533]), .Z(n33359) );
  ANDN U22888 ( .B(n10187), .A(n33359), .Z(n53605) );
  NANDN U22889 ( .A(x[1531]), .B(y[1531]), .Z(n27758) );
  NANDN U22890 ( .A(x[1532]), .B(y[1532]), .Z(n10188) );
  NAND U22891 ( .A(n27758), .B(n10188), .Z(n53604) );
  ANDN U22892 ( .B(x[1530]), .A(y[1530]), .Z(n33352) );
  ANDN U22893 ( .B(x[1531]), .A(y[1531]), .Z(n33358) );
  NOR U22894 ( .A(n33352), .B(n33358), .Z(n53603) );
  NANDN U22895 ( .A(x[1529]), .B(y[1529]), .Z(n27760) );
  XNOR U22896 ( .A(y[1530]), .B(x[1530]), .Z(n10189) );
  NAND U22897 ( .A(n27760), .B(n10189), .Z(n53602) );
  NANDN U22898 ( .A(y[1528]), .B(x[1528]), .Z(n33347) );
  ANDN U22899 ( .B(x[1529]), .A(y[1529]), .Z(n33353) );
  ANDN U22900 ( .B(n33347), .A(n33353), .Z(n53601) );
  ANDN U22901 ( .B(y[1527]), .A(x[1527]), .Z(n33344) );
  NANDN U22902 ( .A(x[1528]), .B(y[1528]), .Z(n27761) );
  NANDN U22903 ( .A(n33344), .B(n27761), .Z(n53600) );
  NANDN U22904 ( .A(y[1525]), .B(x[1525]), .Z(n27762) );
  NANDN U22905 ( .A(y[1524]), .B(x[1524]), .Z(n33339) );
  AND U22906 ( .A(n27762), .B(n33339), .Z(n12716) );
  ANDN U22907 ( .B(y[1523]), .A(x[1523]), .Z(n52258) );
  NANDN U22908 ( .A(y[1523]), .B(x[1523]), .Z(n33338) );
  ANDN U22909 ( .B(y[1521]), .A(x[1521]), .Z(n27767) );
  ANDN U22910 ( .B(y[1522]), .A(x[1522]), .Z(n33336) );
  OR U22911 ( .A(n27767), .B(n33336), .Z(n53594) );
  NANDN U22912 ( .A(y[1521]), .B(x[1521]), .Z(n33332) );
  ANDN U22913 ( .B(x[1520]), .A(y[1520]), .Z(n33328) );
  ANDN U22914 ( .B(n33332), .A(n33328), .Z(n53593) );
  ANDN U22915 ( .B(y[1520]), .A(x[1520]), .Z(n27766) );
  NANDN U22916 ( .A(x[1519]), .B(y[1519]), .Z(n33324) );
  NANDN U22917 ( .A(n27766), .B(n33324), .Z(n53592) );
  NANDN U22918 ( .A(y[1518]), .B(x[1518]), .Z(n27768) );
  ANDN U22919 ( .B(x[1519]), .A(y[1519]), .Z(n53590) );
  ANDN U22920 ( .B(n27768), .A(n53590), .Z(n12707) );
  ANDN U22921 ( .B(y[1517]), .A(x[1517]), .Z(n27770) );
  NANDN U22922 ( .A(y[1517]), .B(x[1517]), .Z(n27769) );
  NANDN U22923 ( .A(y[1516]), .B(x[1516]), .Z(n33320) );
  AND U22924 ( .A(n27769), .B(n33320), .Z(n12703) );
  ANDN U22925 ( .B(y[1515]), .A(x[1515]), .Z(n27772) );
  NANDN U22926 ( .A(y[1515]), .B(x[1515]), .Z(n33319) );
  ANDN U22927 ( .B(y[1513]), .A(x[1513]), .Z(n53584) );
  NANDN U22928 ( .A(y[1512]), .B(x[1512]), .Z(n33309) );
  NANDN U22929 ( .A(y[1513]), .B(x[1513]), .Z(n33316) );
  AND U22930 ( .A(n33309), .B(n33316), .Z(n53583) );
  NANDN U22931 ( .A(x[1511]), .B(y[1511]), .Z(n27775) );
  XNOR U22932 ( .A(y[1512]), .B(x[1512]), .Z(n10190) );
  NAND U22933 ( .A(n27775), .B(n10190), .Z(n53582) );
  NANDN U22934 ( .A(y[1510]), .B(x[1510]), .Z(n27776) );
  NANDN U22935 ( .A(y[1511]), .B(x[1511]), .Z(n33308) );
  AND U22936 ( .A(n27776), .B(n33308), .Z(n52260) );
  NANDN U22937 ( .A(y[1509]), .B(x[1509]), .Z(n27777) );
  ANDN U22938 ( .B(x[1508]), .A(y[1508]), .Z(n33299) );
  ANDN U22939 ( .B(n27777), .A(n33299), .Z(n53581) );
  NANDN U22940 ( .A(x[1507]), .B(y[1507]), .Z(n27781) );
  NANDN U22941 ( .A(x[1508]), .B(y[1508]), .Z(n27778) );
  NAND U22942 ( .A(n27781), .B(n27778), .Z(n53580) );
  NANDN U22943 ( .A(y[1505]), .B(x[1505]), .Z(n27782) );
  NANDN U22944 ( .A(y[1504]), .B(x[1504]), .Z(n27785) );
  AND U22945 ( .A(n27782), .B(n27785), .Z(n12685) );
  NANDN U22946 ( .A(x[1504]), .B(y[1504]), .Z(n27784) );
  ANDN U22947 ( .B(y[1503]), .A(x[1503]), .Z(n33287) );
  ANDN U22948 ( .B(n27784), .A(n33287), .Z(n53573) );
  NANDN U22949 ( .A(y[1502]), .B(x[1502]), .Z(n33283) );
  NANDN U22950 ( .A(y[1503]), .B(x[1503]), .Z(n33291) );
  NAND U22951 ( .A(n33283), .B(n33291), .Z(n53572) );
  NANDN U22952 ( .A(x[1501]), .B(y[1501]), .Z(n27786) );
  ANDN U22953 ( .B(y[1502]), .A(x[1502]), .Z(n33289) );
  ANDN U22954 ( .B(n27786), .A(n33289), .Z(n53571) );
  NANDN U22955 ( .A(y[1501]), .B(x[1501]), .Z(n53570) );
  NANDN U22956 ( .A(x[1499]), .B(y[1499]), .Z(n53567) );
  NANDN U22957 ( .A(x[1500]), .B(y[1500]), .Z(n53569) );
  AND U22958 ( .A(n53567), .B(n53569), .Z(n12678) );
  ANDN U22959 ( .B(x[1498]), .A(y[1498]), .Z(n52262) );
  NANDN U22960 ( .A(y[1499]), .B(x[1499]), .Z(n27788) );
  ANDN U22961 ( .B(y[1498]), .A(x[1498]), .Z(n33279) );
  NANDN U22962 ( .A(x[1497]), .B(y[1497]), .Z(n27789) );
  NANDN U22963 ( .A(n33279), .B(n27789), .Z(n53566) );
  ANDN U22964 ( .B(x[1497]), .A(y[1497]), .Z(n33276) );
  NANDN U22965 ( .A(y[1496]), .B(x[1496]), .Z(n33268) );
  NANDN U22966 ( .A(n33276), .B(n33268), .Z(n52263) );
  NANDN U22967 ( .A(x[1495]), .B(y[1495]), .Z(n27791) );
  NANDN U22968 ( .A(x[1496]), .B(y[1496]), .Z(n27790) );
  AND U22969 ( .A(n27791), .B(n27790), .Z(n53565) );
  NANDN U22970 ( .A(y[1494]), .B(x[1494]), .Z(n33262) );
  NANDN U22971 ( .A(y[1495]), .B(x[1495]), .Z(n33269) );
  NAND U22972 ( .A(n33262), .B(n33269), .Z(n53564) );
  NANDN U22973 ( .A(x[1493]), .B(y[1493]), .Z(n27793) );
  NANDN U22974 ( .A(x[1494]), .B(y[1494]), .Z(n27792) );
  AND U22975 ( .A(n27793), .B(n27792), .Z(n53563) );
  NANDN U22976 ( .A(y[1492]), .B(x[1492]), .Z(n33256) );
  NANDN U22977 ( .A(y[1493]), .B(x[1493]), .Z(n33263) );
  NAND U22978 ( .A(n33256), .B(n33263), .Z(n53562) );
  NANDN U22979 ( .A(x[1491]), .B(y[1491]), .Z(n27796) );
  NANDN U22980 ( .A(x[1492]), .B(y[1492]), .Z(n27794) );
  AND U22981 ( .A(n27796), .B(n27794), .Z(n53560) );
  ANDN U22982 ( .B(x[1490]), .A(y[1490]), .Z(n33251) );
  NANDN U22983 ( .A(y[1491]), .B(x[1491]), .Z(n33257) );
  NANDN U22984 ( .A(n33251), .B(n33257), .Z(n53559) );
  NANDN U22985 ( .A(x[1489]), .B(y[1489]), .Z(n27797) );
  XNOR U22986 ( .A(y[1490]), .B(x[1490]), .Z(n10191) );
  AND U22987 ( .A(n27797), .B(n10191), .Z(n53558) );
  ANDN U22988 ( .B(x[1488]), .A(y[1488]), .Z(n33245) );
  ANDN U22989 ( .B(x[1489]), .A(y[1489]), .Z(n33252) );
  NOR U22990 ( .A(n33245), .B(n33252), .Z(n53557) );
  NANDN U22991 ( .A(x[1487]), .B(y[1487]), .Z(n33241) );
  NANDN U22992 ( .A(x[1488]), .B(y[1488]), .Z(n27798) );
  NAND U22993 ( .A(n33241), .B(n27798), .Z(n52264) );
  ANDN U22994 ( .B(x[1486]), .A(y[1486]), .Z(n27800) );
  ANDN U22995 ( .B(x[1487]), .A(y[1487]), .Z(n33246) );
  NOR U22996 ( .A(n27800), .B(n33246), .Z(n53556) );
  NANDN U22997 ( .A(y[1484]), .B(x[1484]), .Z(n27801) );
  ANDN U22998 ( .B(x[1485]), .A(y[1485]), .Z(n27799) );
  ANDN U22999 ( .B(n27801), .A(n27799), .Z(n53554) );
  NANDN U23000 ( .A(y[1482]), .B(x[1482]), .Z(n53552) );
  NANDN U23001 ( .A(y[1483]), .B(x[1483]), .Z(n52266) );
  AND U23002 ( .A(n53552), .B(n52266), .Z(n12658) );
  NANDN U23003 ( .A(y[1481]), .B(x[1481]), .Z(n27802) );
  NANDN U23004 ( .A(y[1480]), .B(x[1480]), .Z(n10192) );
  AND U23005 ( .A(n27802), .B(n10192), .Z(n53550) );
  NANDN U23006 ( .A(x[1479]), .B(y[1479]), .Z(n33220) );
  ANDN U23007 ( .B(y[1480]), .A(x[1480]), .Z(n27803) );
  ANDN U23008 ( .B(n33220), .A(n27803), .Z(n53549) );
  ANDN U23009 ( .B(x[1478]), .A(y[1478]), .Z(n33216) );
  NANDN U23010 ( .A(y[1479]), .B(x[1479]), .Z(n33224) );
  NANDN U23011 ( .A(n33216), .B(n33224), .Z(n53547) );
  NANDN U23012 ( .A(x[1477]), .B(y[1477]), .Z(n33212) );
  ANDN U23013 ( .B(y[1478]), .A(x[1478]), .Z(n33222) );
  ANDN U23014 ( .B(n33212), .A(n33222), .Z(n53546) );
  ANDN U23015 ( .B(x[1476]), .A(y[1476]), .Z(n33207) );
  ANDN U23016 ( .B(x[1477]), .A(y[1477]), .Z(n33218) );
  OR U23017 ( .A(n33207), .B(n33218), .Z(n53545) );
  NANDN U23018 ( .A(x[1475]), .B(y[1475]), .Z(n33205) );
  NANDN U23019 ( .A(x[1476]), .B(y[1476]), .Z(n33211) );
  AND U23020 ( .A(n33205), .B(n33211), .Z(n53544) );
  ANDN U23021 ( .B(x[1474]), .A(y[1474]), .Z(n33202) );
  ANDN U23022 ( .B(x[1475]), .A(y[1475]), .Z(n33210) );
  OR U23023 ( .A(n33202), .B(n33210), .Z(n53543) );
  NANDN U23024 ( .A(x[1474]), .B(y[1474]), .Z(n53542) );
  ANDN U23025 ( .B(x[1473]), .A(y[1473]), .Z(n53541) );
  NANDN U23026 ( .A(x[1473]), .B(y[1473]), .Z(n10194) );
  NANDN U23027 ( .A(x[1472]), .B(y[1472]), .Z(n10193) );
  AND U23028 ( .A(n10194), .B(n10193), .Z(n53540) );
  NANDN U23029 ( .A(y[1471]), .B(x[1471]), .Z(n10196) );
  NANDN U23030 ( .A(y[1472]), .B(x[1472]), .Z(n10195) );
  NAND U23031 ( .A(n10196), .B(n10195), .Z(n27809) );
  NANDN U23032 ( .A(x[1471]), .B(y[1471]), .Z(n12642) );
  NANDN U23033 ( .A(x[1470]), .B(y[1470]), .Z(n10197) );
  AND U23034 ( .A(n12642), .B(n10197), .Z(n27807) );
  NANDN U23035 ( .A(x[1469]), .B(y[1469]), .Z(n10198) );
  AND U23036 ( .A(n27807), .B(n10198), .Z(n53538) );
  NANDN U23037 ( .A(x[1468]), .B(y[1468]), .Z(n27810) );
  ANDN U23038 ( .B(y[1467]), .A(x[1467]), .Z(n33191) );
  ANDN U23039 ( .B(n27810), .A(n33191), .Z(n53536) );
  NANDN U23040 ( .A(y[1466]), .B(x[1466]), .Z(n33187) );
  NANDN U23041 ( .A(y[1467]), .B(x[1467]), .Z(n33195) );
  NAND U23042 ( .A(n33187), .B(n33195), .Z(n53535) );
  ANDN U23043 ( .B(y[1466]), .A(x[1466]), .Z(n33193) );
  NANDN U23044 ( .A(x[1465]), .B(y[1465]), .Z(n27812) );
  NANDN U23045 ( .A(n33193), .B(n27812), .Z(n52267) );
  NANDN U23046 ( .A(x[1464]), .B(y[1464]), .Z(n53533) );
  NANDN U23047 ( .A(x[1463]), .B(y[1463]), .Z(n27815) );
  AND U23048 ( .A(n53533), .B(n27815), .Z(n12632) );
  ANDN U23049 ( .B(x[1462]), .A(y[1462]), .Z(n33177) );
  ANDN U23050 ( .B(y[1461]), .A(x[1461]), .Z(n33173) );
  ANDN U23051 ( .B(y[1462]), .A(x[1462]), .Z(n33182) );
  NOR U23052 ( .A(n33173), .B(n33182), .Z(n53528) );
  ANDN U23053 ( .B(y[1459]), .A(x[1459]), .Z(n33166) );
  ANDN U23054 ( .B(y[1460]), .A(x[1460]), .Z(n33176) );
  NOR U23055 ( .A(n33166), .B(n33176), .Z(n53527) );
  NANDN U23056 ( .A(y[1458]), .B(x[1458]), .Z(n27816) );
  NANDN U23057 ( .A(y[1459]), .B(x[1459]), .Z(n33171) );
  NAND U23058 ( .A(n27816), .B(n33171), .Z(n53526) );
  ANDN U23059 ( .B(y[1457]), .A(x[1457]), .Z(n33160) );
  ANDN U23060 ( .B(y[1458]), .A(x[1458]), .Z(n33168) );
  NOR U23061 ( .A(n33160), .B(n33168), .Z(n53525) );
  NANDN U23062 ( .A(y[1456]), .B(x[1456]), .Z(n33156) );
  NANDN U23063 ( .A(y[1457]), .B(x[1457]), .Z(n27817) );
  NAND U23064 ( .A(n33156), .B(n27817), .Z(n52269) );
  NANDN U23065 ( .A(x[1455]), .B(y[1455]), .Z(n27818) );
  XNOR U23066 ( .A(y[1456]), .B(x[1456]), .Z(n10199) );
  AND U23067 ( .A(n27818), .B(n10199), .Z(n52270) );
  NANDN U23068 ( .A(y[1452]), .B(x[1452]), .Z(n27824) );
  NANDN U23069 ( .A(y[1453]), .B(x[1453]), .Z(n27821) );
  NAND U23070 ( .A(n27824), .B(n27821), .Z(n53523) );
  NANDN U23071 ( .A(x[1452]), .B(y[1452]), .Z(n27823) );
  ANDN U23072 ( .B(y[1451]), .A(x[1451]), .Z(n33143) );
  ANDN U23073 ( .B(n27823), .A(n33143), .Z(n53522) );
  NANDN U23074 ( .A(y[1450]), .B(x[1450]), .Z(n33140) );
  NANDN U23075 ( .A(y[1451]), .B(x[1451]), .Z(n27825) );
  NAND U23076 ( .A(n33140), .B(n27825), .Z(n52272) );
  ANDN U23077 ( .B(y[1449]), .A(x[1449]), .Z(n33136) );
  ANDN U23078 ( .B(y[1450]), .A(x[1450]), .Z(n33146) );
  NOR U23079 ( .A(n33136), .B(n33146), .Z(n53520) );
  ANDN U23080 ( .B(y[1447]), .A(x[1447]), .Z(n33130) );
  ANDN U23081 ( .B(y[1448]), .A(x[1448]), .Z(n33138) );
  NOR U23082 ( .A(n33130), .B(n33138), .Z(n53519) );
  NANDN U23083 ( .A(y[1446]), .B(x[1446]), .Z(n33128) );
  NANDN U23084 ( .A(y[1447]), .B(x[1447]), .Z(n33131) );
  NAND U23085 ( .A(n33128), .B(n33131), .Z(n53518) );
  NANDN U23086 ( .A(x[1446]), .B(y[1446]), .Z(n10201) );
  NANDN U23087 ( .A(x[1445]), .B(y[1445]), .Z(n10200) );
  AND U23088 ( .A(n10201), .B(n10200), .Z(n33125) );
  NANDN U23089 ( .A(y[1444]), .B(x[1444]), .Z(n10203) );
  NANDN U23090 ( .A(y[1445]), .B(x[1445]), .Z(n10202) );
  AND U23091 ( .A(n10203), .B(n10202), .Z(n27829) );
  NANDN U23092 ( .A(x[1443]), .B(y[1443]), .Z(n10204) );
  ANDN U23093 ( .B(y[1444]), .A(x[1444]), .Z(n27827) );
  ANDN U23094 ( .B(n10204), .A(n27827), .Z(n12608) );
  NANDN U23095 ( .A(y[1442]), .B(x[1442]), .Z(n27831) );
  NANDN U23096 ( .A(y[1443]), .B(x[1443]), .Z(n27826) );
  NAND U23097 ( .A(n27831), .B(n27826), .Z(n10205) );
  NAND U23098 ( .A(n12608), .B(n10205), .Z(n10206) );
  NAND U23099 ( .A(n27829), .B(n10206), .Z(n52274) );
  NANDN U23100 ( .A(x[1441]), .B(y[1441]), .Z(n33117) );
  ANDN U23101 ( .B(x[1441]), .A(y[1441]), .Z(n27830) );
  ANDN U23102 ( .B(y[1439]), .A(x[1439]), .Z(n53513) );
  NANDN U23103 ( .A(x[1440]), .B(y[1440]), .Z(n33118) );
  ANDN U23104 ( .B(x[1438]), .A(y[1438]), .Z(n53512) );
  NANDN U23105 ( .A(x[1437]), .B(y[1437]), .Z(n33107) );
  NANDN U23106 ( .A(x[1438]), .B(y[1438]), .Z(n33114) );
  AND U23107 ( .A(n33107), .B(n33114), .Z(n53511) );
  ANDN U23108 ( .B(x[1436]), .A(y[1436]), .Z(n33103) );
  ANDN U23109 ( .B(x[1437]), .A(y[1437]), .Z(n33111) );
  OR U23110 ( .A(n33103), .B(n33111), .Z(n53510) );
  ANDN U23111 ( .B(x[1435]), .A(y[1435]), .Z(n52277) );
  NANDN U23112 ( .A(x[1433]), .B(y[1433]), .Z(n27836) );
  NANDN U23113 ( .A(y[1432]), .B(x[1432]), .Z(n27837) );
  ANDN U23114 ( .B(x[1433]), .A(y[1433]), .Z(n33098) );
  ANDN U23115 ( .B(n27837), .A(n33098), .Z(n12593) );
  NANDN U23116 ( .A(x[1431]), .B(y[1431]), .Z(n27841) );
  NANDN U23117 ( .A(y[1431]), .B(x[1431]), .Z(n27838) );
  NANDN U23118 ( .A(x[1429]), .B(y[1429]), .Z(n53502) );
  NANDN U23119 ( .A(y[1428]), .B(x[1428]), .Z(n10207) );
  ANDN U23120 ( .B(x[1429]), .A(y[1429]), .Z(n33089) );
  ANDN U23121 ( .B(n10207), .A(n33089), .Z(n53501) );
  ANDN U23122 ( .B(y[1427]), .A(x[1427]), .Z(n33083) );
  ANDN U23123 ( .B(y[1428]), .A(x[1428]), .Z(n33088) );
  OR U23124 ( .A(n33083), .B(n33088), .Z(n53500) );
  NANDN U23125 ( .A(y[1426]), .B(x[1426]), .Z(n33079) );
  ANDN U23126 ( .B(x[1427]), .A(y[1427]), .Z(n33087) );
  ANDN U23127 ( .B(n33079), .A(n33087), .Z(n53499) );
  ANDN U23128 ( .B(y[1425]), .A(x[1425]), .Z(n27843) );
  NANDN U23129 ( .A(y[1424]), .B(x[1424]), .Z(n27844) );
  NANDN U23130 ( .A(y[1425]), .B(x[1425]), .Z(n53498) );
  AND U23131 ( .A(n27844), .B(n53498), .Z(n12580) );
  ANDN U23132 ( .B(y[1423]), .A(x[1423]), .Z(n33075) );
  NANDN U23133 ( .A(y[1423]), .B(x[1423]), .Z(n27845) );
  XOR U23134 ( .A(x[1422]), .B(y[1422]), .Z(n27846) );
  NANDN U23135 ( .A(y[1419]), .B(x[1419]), .Z(n33068) );
  ANDN U23136 ( .B(x[1418]), .A(y[1418]), .Z(n33063) );
  ANDN U23137 ( .B(n33068), .A(n33063), .Z(n53491) );
  ANDN U23138 ( .B(y[1418]), .A(x[1418]), .Z(n27849) );
  NANDN U23139 ( .A(x[1417]), .B(y[1417]), .Z(n27851) );
  NANDN U23140 ( .A(n27849), .B(n27851), .Z(n53490) );
  NANDN U23141 ( .A(y[1417]), .B(x[1417]), .Z(n33064) );
  NANDN U23142 ( .A(y[1416]), .B(x[1416]), .Z(n27852) );
  NANDN U23143 ( .A(y[1415]), .B(x[1415]), .Z(n27853) );
  NANDN U23144 ( .A(y[1414]), .B(x[1414]), .Z(n27855) );
  AND U23145 ( .A(n27853), .B(n27855), .Z(n12562) );
  ANDN U23146 ( .B(y[1411]), .A(x[1411]), .Z(n33047) );
  ANDN U23147 ( .B(y[1412]), .A(x[1412]), .Z(n33053) );
  OR U23148 ( .A(n33047), .B(n33053), .Z(n53480) );
  NANDN U23149 ( .A(y[1410]), .B(x[1410]), .Z(n27859) );
  NANDN U23150 ( .A(y[1411]), .B(x[1411]), .Z(n27857) );
  NAND U23151 ( .A(n27859), .B(n27857), .Z(n53479) );
  NANDN U23152 ( .A(x[1409]), .B(y[1409]), .Z(n10208) );
  ANDN U23153 ( .B(y[1410]), .A(x[1410]), .Z(n27861) );
  ANDN U23154 ( .B(n10208), .A(n27861), .Z(n53478) );
  NANDN U23155 ( .A(y[1409]), .B(x[1409]), .Z(n27858) );
  ANDN U23156 ( .B(x[1408]), .A(y[1408]), .Z(n33037) );
  ANDN U23157 ( .B(n27858), .A(n33037), .Z(n53477) );
  NANDN U23158 ( .A(x[1408]), .B(y[1408]), .Z(n33040) );
  NANDN U23159 ( .A(x[1407]), .B(y[1407]), .Z(n10209) );
  NAND U23160 ( .A(n33040), .B(n10209), .Z(n27862) );
  NANDN U23161 ( .A(y[1406]), .B(x[1406]), .Z(n33031) );
  ANDN U23162 ( .B(x[1407]), .A(y[1407]), .Z(n33038) );
  ANDN U23163 ( .B(n33031), .A(n33038), .Z(n53475) );
  NANDN U23164 ( .A(x[1403]), .B(y[1403]), .Z(n33023) );
  NANDN U23165 ( .A(x[1404]), .B(y[1404]), .Z(n33028) );
  NAND U23166 ( .A(n33023), .B(n33028), .Z(n53473) );
  NANDN U23167 ( .A(y[1403]), .B(x[1403]), .Z(n27865) );
  ANDN U23168 ( .B(x[1402]), .A(y[1402]), .Z(n33019) );
  ANDN U23169 ( .B(n27865), .A(n33019), .Z(n53472) );
  ANDN U23170 ( .B(y[1402]), .A(x[1402]), .Z(n53471) );
  NANDN U23171 ( .A(x[1401]), .B(y[1401]), .Z(n27867) );
  NANDN U23172 ( .A(n53471), .B(n27867), .Z(n12548) );
  NANDN U23173 ( .A(y[1400]), .B(x[1400]), .Z(n27868) );
  NANDN U23174 ( .A(y[1401]), .B(x[1401]), .Z(n33020) );
  AND U23175 ( .A(n27868), .B(n33020), .Z(n12546) );
  NANDN U23176 ( .A(x[1399]), .B(y[1399]), .Z(n27871) );
  NANDN U23177 ( .A(y[1396]), .B(x[1396]), .Z(n27873) );
  ANDN U23178 ( .B(x[1397]), .A(y[1397]), .Z(n33012) );
  ANDN U23179 ( .B(n27873), .A(n33012), .Z(n53464) );
  NANDN U23180 ( .A(x[1395]), .B(y[1395]), .Z(n27874) );
  NANDN U23181 ( .A(x[1396]), .B(y[1396]), .Z(n33008) );
  NAND U23182 ( .A(n27874), .B(n33008), .Z(n52283) );
  NANDN U23183 ( .A(y[1394]), .B(x[1394]), .Z(n33000) );
  NANDN U23184 ( .A(y[1395]), .B(x[1395]), .Z(n27872) );
  NAND U23185 ( .A(n33000), .B(n27872), .Z(n53462) );
  NANDN U23186 ( .A(x[1393]), .B(y[1393]), .Z(n32995) );
  NANDN U23187 ( .A(x[1394]), .B(y[1394]), .Z(n27875) );
  AND U23188 ( .A(n32995), .B(n27875), .Z(n53461) );
  NANDN U23189 ( .A(y[1392]), .B(x[1392]), .Z(n27876) );
  NANDN U23190 ( .A(y[1393]), .B(x[1393]), .Z(n33001) );
  NAND U23191 ( .A(n27876), .B(n33001), .Z(n53460) );
  NANDN U23192 ( .A(x[1391]), .B(y[1391]), .Z(n32990) );
  NANDN U23193 ( .A(x[1392]), .B(y[1392]), .Z(n32996) );
  AND U23194 ( .A(n32990), .B(n32996), .Z(n53459) );
  NANDN U23195 ( .A(y[1390]), .B(x[1390]), .Z(n27878) );
  NANDN U23196 ( .A(y[1391]), .B(x[1391]), .Z(n27877) );
  NAND U23197 ( .A(n27878), .B(n27877), .Z(n53458) );
  NANDN U23198 ( .A(x[1389]), .B(y[1389]), .Z(n27880) );
  ANDN U23199 ( .B(x[1388]), .A(y[1388]), .Z(n27881) );
  ANDN U23200 ( .B(y[1387]), .A(x[1387]), .Z(n27884) );
  NANDN U23201 ( .A(y[1387]), .B(x[1387]), .Z(n27882) );
  ANDN U23202 ( .B(y[1385]), .A(x[1385]), .Z(n52285) );
  NANDN U23203 ( .A(x[1381]), .B(y[1381]), .Z(n10211) );
  NANDN U23204 ( .A(x[1382]), .B(y[1382]), .Z(n10210) );
  NAND U23205 ( .A(n10211), .B(n10210), .Z(n53447) );
  NANDN U23206 ( .A(y[1381]), .B(x[1381]), .Z(n10213) );
  NANDN U23207 ( .A(y[1380]), .B(x[1380]), .Z(n10212) );
  AND U23208 ( .A(n10213), .B(n10212), .Z(n27892) );
  NANDN U23209 ( .A(x[1379]), .B(y[1379]), .Z(n10214) );
  NANDN U23210 ( .A(x[1380]), .B(y[1380]), .Z(n27888) );
  AND U23211 ( .A(n10214), .B(n27888), .Z(n53445) );
  NANDN U23212 ( .A(y[1378]), .B(x[1378]), .Z(n32973) );
  NANDN U23213 ( .A(x[1377]), .B(y[1377]), .Z(n32968) );
  NANDN U23214 ( .A(x[1378]), .B(y[1378]), .Z(n32976) );
  NAND U23215 ( .A(n32968), .B(n32976), .Z(n52286) );
  ANDN U23216 ( .B(x[1376]), .A(y[1376]), .Z(n32963) );
  ANDN U23217 ( .B(x[1377]), .A(y[1377]), .Z(n32972) );
  NOR U23218 ( .A(n32963), .B(n32972), .Z(n53443) );
  NANDN U23219 ( .A(x[1375]), .B(y[1375]), .Z(n32960) );
  NANDN U23220 ( .A(x[1376]), .B(y[1376]), .Z(n32967) );
  AND U23221 ( .A(n32960), .B(n32967), .Z(n53442) );
  ANDN U23222 ( .B(x[1374]), .A(y[1374]), .Z(n32956) );
  ANDN U23223 ( .B(x[1375]), .A(y[1375]), .Z(n32966) );
  OR U23224 ( .A(n32956), .B(n32966), .Z(n53441) );
  NANDN U23225 ( .A(x[1373]), .B(y[1373]), .Z(n27893) );
  NANDN U23226 ( .A(x[1374]), .B(y[1374]), .Z(n32961) );
  AND U23227 ( .A(n27893), .B(n32961), .Z(n52287) );
  ANDN U23228 ( .B(x[1371]), .A(y[1371]), .Z(n32951) );
  NANDN U23229 ( .A(y[1370]), .B(x[1370]), .Z(n27896) );
  NANDN U23230 ( .A(n32951), .B(n27896), .Z(n53438) );
  NANDN U23231 ( .A(x[1369]), .B(y[1369]), .Z(n27897) );
  NANDN U23232 ( .A(x[1370]), .B(y[1370]), .Z(n32945) );
  AND U23233 ( .A(n27897), .B(n32945), .Z(n52289) );
  NANDN U23234 ( .A(y[1368]), .B(x[1368]), .Z(n27900) );
  NANDN U23235 ( .A(y[1369]), .B(x[1369]), .Z(n27895) );
  NAND U23236 ( .A(n27900), .B(n27895), .Z(n52290) );
  NANDN U23237 ( .A(x[1367]), .B(y[1367]), .Z(n32936) );
  NANDN U23238 ( .A(x[1368]), .B(y[1368]), .Z(n27898) );
  AND U23239 ( .A(n32936), .B(n27898), .Z(n52291) );
  NANDN U23240 ( .A(x[1365]), .B(y[1365]), .Z(n27901) );
  ANDN U23241 ( .B(y[1366]), .A(x[1366]), .Z(n32938) );
  ANDN U23242 ( .B(n27901), .A(n32938), .Z(n53435) );
  ANDN U23243 ( .B(x[1364]), .A(y[1364]), .Z(n32926) );
  ANDN U23244 ( .B(x[1365]), .A(y[1365]), .Z(n32934) );
  OR U23245 ( .A(n32926), .B(n32934), .Z(n53434) );
  NANDN U23246 ( .A(x[1363]), .B(y[1363]), .Z(n32922) );
  NANDN U23247 ( .A(x[1364]), .B(y[1364]), .Z(n27902) );
  AND U23248 ( .A(n32922), .B(n27902), .Z(n52293) );
  ANDN U23249 ( .B(x[1363]), .A(y[1363]), .Z(n32927) );
  NANDN U23250 ( .A(y[1362]), .B(x[1362]), .Z(n27903) );
  NANDN U23251 ( .A(n32927), .B(n27903), .Z(n52294) );
  NANDN U23252 ( .A(x[1361]), .B(y[1361]), .Z(n32915) );
  NANDN U23253 ( .A(x[1362]), .B(y[1362]), .Z(n32924) );
  AND U23254 ( .A(n32915), .B(n32924), .Z(n52295) );
  NANDN U23255 ( .A(y[1358]), .B(x[1358]), .Z(n27907) );
  NANDN U23256 ( .A(y[1359]), .B(x[1359]), .Z(n27906) );
  NAND U23257 ( .A(n27907), .B(n27906), .Z(n53430) );
  NANDN U23258 ( .A(x[1357]), .B(y[1357]), .Z(n32903) );
  NANDN U23259 ( .A(x[1358]), .B(y[1358]), .Z(n32910) );
  AND U23260 ( .A(n32903), .B(n32910), .Z(n52297) );
  NANDN U23261 ( .A(y[1356]), .B(x[1356]), .Z(n27910) );
  NANDN U23262 ( .A(y[1357]), .B(x[1357]), .Z(n27908) );
  NAND U23263 ( .A(n27910), .B(n27908), .Z(n52298) );
  NANDN U23264 ( .A(x[1356]), .B(y[1356]), .Z(n32904) );
  ANDN U23265 ( .B(y[1355]), .A(x[1355]), .Z(n32898) );
  ANDN U23266 ( .B(n32904), .A(n32898), .Z(n53429) );
  ANDN U23267 ( .B(y[1353]), .A(x[1353]), .Z(n32893) );
  ANDN U23268 ( .B(y[1354]), .A(x[1354]), .Z(n32899) );
  NOR U23269 ( .A(n32893), .B(n32899), .Z(n53428) );
  NANDN U23270 ( .A(y[1352]), .B(x[1352]), .Z(n32889) );
  NANDN U23271 ( .A(y[1353]), .B(x[1353]), .Z(n27912) );
  NAND U23272 ( .A(n32889), .B(n27912), .Z(n53427) );
  ANDN U23273 ( .B(y[1352]), .A(x[1352]), .Z(n53425) );
  NANDN U23274 ( .A(y[1351]), .B(x[1351]), .Z(n52300) );
  NANDN U23275 ( .A(x[1350]), .B(y[1350]), .Z(n53424) );
  NANDN U23276 ( .A(x[1351]), .B(y[1351]), .Z(n53426) );
  NAND U23277 ( .A(n53424), .B(n53426), .Z(n32888) );
  NANDN U23278 ( .A(y[1348]), .B(x[1348]), .Z(n32879) );
  NANDN U23279 ( .A(y[1349]), .B(x[1349]), .Z(n27914) );
  NAND U23280 ( .A(n32879), .B(n27914), .Z(n53422) );
  ANDN U23281 ( .B(y[1347]), .A(x[1347]), .Z(n32874) );
  ANDN U23282 ( .B(y[1348]), .A(x[1348]), .Z(n32883) );
  NOR U23283 ( .A(n32874), .B(n32883), .Z(n53421) );
  NANDN U23284 ( .A(y[1346]), .B(x[1346]), .Z(n32871) );
  NANDN U23285 ( .A(y[1347]), .B(x[1347]), .Z(n32878) );
  NAND U23286 ( .A(n32871), .B(n32878), .Z(n53420) );
  ANDN U23287 ( .B(y[1345]), .A(x[1345]), .Z(n32867) );
  ANDN U23288 ( .B(y[1346]), .A(x[1346]), .Z(n32877) );
  NOR U23289 ( .A(n32867), .B(n32877), .Z(n53419) );
  NANDN U23290 ( .A(y[1344]), .B(x[1344]), .Z(n27915) );
  NANDN U23291 ( .A(y[1345]), .B(x[1345]), .Z(n32872) );
  NAND U23292 ( .A(n27915), .B(n32872), .Z(n53417) );
  ANDN U23293 ( .B(y[1343]), .A(x[1343]), .Z(n32861) );
  ANDN U23294 ( .B(y[1344]), .A(x[1344]), .Z(n32869) );
  NOR U23295 ( .A(n32861), .B(n32869), .Z(n53416) );
  NANDN U23296 ( .A(y[1342]), .B(x[1342]), .Z(n32857) );
  NANDN U23297 ( .A(y[1343]), .B(x[1343]), .Z(n27916) );
  NAND U23298 ( .A(n32857), .B(n27916), .Z(n53415) );
  XNOR U23299 ( .A(x[1342]), .B(y[1342]), .Z(n10215) );
  ANDN U23300 ( .B(y[1341]), .A(x[1341]), .Z(n27918) );
  ANDN U23301 ( .B(n10215), .A(n27918), .Z(n53414) );
  NANDN U23302 ( .A(x[1339]), .B(y[1339]), .Z(n27919) );
  ANDN U23303 ( .B(y[1340]), .A(x[1340]), .Z(n27917) );
  ANDN U23304 ( .B(n27919), .A(n27917), .Z(n53413) );
  NANDN U23305 ( .A(x[1338]), .B(y[1338]), .Z(n53412) );
  NANDN U23306 ( .A(x[1337]), .B(y[1337]), .Z(n27921) );
  NAND U23307 ( .A(n53412), .B(n27921), .Z(n53409) );
  ANDN U23308 ( .B(x[1336]), .A(y[1336]), .Z(n53408) );
  NANDN U23309 ( .A(x[1335]), .B(y[1335]), .Z(n27922) );
  NANDN U23310 ( .A(x[1336]), .B(y[1336]), .Z(n27920) );
  NAND U23311 ( .A(n27922), .B(n27920), .Z(n52303) );
  ANDN U23312 ( .B(x[1334]), .A(y[1334]), .Z(n32836) );
  ANDN U23313 ( .B(x[1335]), .A(y[1335]), .Z(n32842) );
  NOR U23314 ( .A(n32836), .B(n32842), .Z(n53407) );
  NANDN U23315 ( .A(x[1333]), .B(y[1333]), .Z(n32832) );
  XNOR U23316 ( .A(x[1334]), .B(y[1334]), .Z(n10216) );
  AND U23317 ( .A(n32832), .B(n10216), .Z(n53406) );
  ANDN U23318 ( .B(x[1333]), .A(y[1333]), .Z(n32837) );
  NANDN U23319 ( .A(y[1332]), .B(x[1332]), .Z(n27924) );
  NANDN U23320 ( .A(n32837), .B(n27924), .Z(n53405) );
  NANDN U23321 ( .A(x[1331]), .B(y[1331]), .Z(n27926) );
  NANDN U23322 ( .A(x[1332]), .B(y[1332]), .Z(n32831) );
  AND U23323 ( .A(n27926), .B(n32831), .Z(n53404) );
  NANDN U23324 ( .A(y[1330]), .B(x[1330]), .Z(n27928) );
  NANDN U23325 ( .A(y[1331]), .B(x[1331]), .Z(n27925) );
  NAND U23326 ( .A(n27928), .B(n27925), .Z(n53402) );
  NANDN U23327 ( .A(x[1329]), .B(y[1329]), .Z(n27931) );
  NANDN U23328 ( .A(x[1330]), .B(y[1330]), .Z(n27927) );
  AND U23329 ( .A(n27931), .B(n27927), .Z(n53400) );
  ANDN U23330 ( .B(x[1328]), .A(y[1328]), .Z(n32820) );
  NANDN U23331 ( .A(y[1329]), .B(x[1329]), .Z(n27929) );
  NANDN U23332 ( .A(n32820), .B(n27929), .Z(n53398) );
  NANDN U23333 ( .A(x[1327]), .B(y[1327]), .Z(n27932) );
  NANDN U23334 ( .A(x[1328]), .B(y[1328]), .Z(n27930) );
  AND U23335 ( .A(n27932), .B(n27930), .Z(n53396) );
  ANDN U23336 ( .B(x[1326]), .A(y[1326]), .Z(n32814) );
  ANDN U23337 ( .B(x[1327]), .A(y[1327]), .Z(n32821) );
  OR U23338 ( .A(n32814), .B(n32821), .Z(n53394) );
  NANDN U23339 ( .A(x[1325]), .B(y[1325]), .Z(n32810) );
  NANDN U23340 ( .A(x[1326]), .B(y[1326]), .Z(n27933) );
  AND U23341 ( .A(n32810), .B(n27933), .Z(n53392) );
  ANDN U23342 ( .B(x[1324]), .A(y[1324]), .Z(n27935) );
  ANDN U23343 ( .B(x[1325]), .A(y[1325]), .Z(n32815) );
  OR U23344 ( .A(n27935), .B(n32815), .Z(n53390) );
  NANDN U23345 ( .A(x[1324]), .B(y[1324]), .Z(n32809) );
  ANDN U23346 ( .B(y[1323]), .A(x[1323]), .Z(n32805) );
  ANDN U23347 ( .B(n32809), .A(n32805), .Z(n53388) );
  ANDN U23348 ( .B(x[1323]), .A(y[1323]), .Z(n27934) );
  NANDN U23349 ( .A(y[1322]), .B(x[1322]), .Z(n10217) );
  NANDN U23350 ( .A(n27934), .B(n10217), .Z(n53386) );
  XNOR U23351 ( .A(y[1322]), .B(x[1322]), .Z(n32800) );
  ANDN U23352 ( .B(y[1321]), .A(x[1321]), .Z(n32795) );
  ANDN U23353 ( .B(n32800), .A(n32795), .Z(n53384) );
  NANDN U23354 ( .A(y[1320]), .B(x[1320]), .Z(n32792) );
  NANDN U23355 ( .A(y[1321]), .B(x[1321]), .Z(n32799) );
  NAND U23356 ( .A(n32792), .B(n32799), .Z(n53382) );
  NANDN U23357 ( .A(x[1319]), .B(y[1319]), .Z(n32787) );
  ANDN U23358 ( .B(y[1320]), .A(x[1320]), .Z(n32798) );
  ANDN U23359 ( .B(n32787), .A(n32798), .Z(n53380) );
  NANDN U23360 ( .A(y[1318]), .B(x[1318]), .Z(n27937) );
  NANDN U23361 ( .A(y[1319]), .B(x[1319]), .Z(n32793) );
  NAND U23362 ( .A(n27937), .B(n32793), .Z(n53378) );
  NANDN U23363 ( .A(x[1318]), .B(y[1318]), .Z(n32788) );
  ANDN U23364 ( .B(y[1317]), .A(x[1317]), .Z(n32782) );
  ANDN U23365 ( .B(n32788), .A(n32782), .Z(n53376) );
  NANDN U23366 ( .A(y[1316]), .B(x[1316]), .Z(n32778) );
  NANDN U23367 ( .A(y[1317]), .B(x[1317]), .Z(n27936) );
  NAND U23368 ( .A(n32778), .B(n27936), .Z(n53374) );
  ANDN U23369 ( .B(y[1315]), .A(x[1315]), .Z(n32773) );
  ANDN U23370 ( .B(y[1316]), .A(x[1316]), .Z(n32783) );
  NOR U23371 ( .A(n32773), .B(n32783), .Z(n53372) );
  NANDN U23372 ( .A(y[1314]), .B(x[1314]), .Z(n32770) );
  NANDN U23373 ( .A(y[1315]), .B(x[1315]), .Z(n32777) );
  NAND U23374 ( .A(n32770), .B(n32777), .Z(n53370) );
  ANDN U23375 ( .B(y[1313]), .A(x[1313]), .Z(n32768) );
  ANDN U23376 ( .B(y[1314]), .A(x[1314]), .Z(n32776) );
  NOR U23377 ( .A(n32768), .B(n32776), .Z(n53368) );
  NANDN U23378 ( .A(y[1312]), .B(x[1312]), .Z(n32766) );
  NANDN U23379 ( .A(y[1313]), .B(x[1313]), .Z(n32771) );
  NAND U23380 ( .A(n32766), .B(n32771), .Z(n53366) );
  NANDN U23381 ( .A(y[1310]), .B(x[1310]), .Z(n10219) );
  NANDN U23382 ( .A(y[1311]), .B(x[1311]), .Z(n10218) );
  AND U23383 ( .A(n10219), .B(n10218), .Z(n27941) );
  NANDN U23384 ( .A(x[1309]), .B(y[1309]), .Z(n10220) );
  ANDN U23385 ( .B(y[1310]), .A(x[1310]), .Z(n27939) );
  ANDN U23386 ( .B(n10220), .A(n27939), .Z(n10224) );
  ANDN U23387 ( .B(x[1308]), .A(y[1308]), .Z(n32759) );
  NANDN U23388 ( .A(y[1309]), .B(x[1309]), .Z(n27938) );
  NANDN U23389 ( .A(n32759), .B(n27938), .Z(n10221) );
  NAND U23390 ( .A(n10224), .B(n10221), .Z(n10222) );
  NAND U23391 ( .A(n27941), .B(n10222), .Z(n53362) );
  NANDN U23392 ( .A(x[1308]), .B(y[1308]), .Z(n10223) );
  AND U23393 ( .A(n10224), .B(n10223), .Z(n53360) );
  NANDN U23394 ( .A(y[1307]), .B(x[1307]), .Z(n52304) );
  NANDN U23395 ( .A(x[1306]), .B(y[1306]), .Z(n53359) );
  NANDN U23396 ( .A(x[1307]), .B(y[1307]), .Z(n53361) );
  AND U23397 ( .A(n53359), .B(n53361), .Z(n32757) );
  NANDN U23398 ( .A(y[1305]), .B(x[1305]), .Z(n53358) );
  ANDN U23399 ( .B(x[1306]), .A(y[1306]), .Z(n12447) );
  IV U23400 ( .A(n12447), .Z(n52305) );
  AND U23401 ( .A(n53358), .B(n52305), .Z(n32755) );
  NANDN U23402 ( .A(y[1302]), .B(x[1302]), .Z(n32743) );
  NANDN U23403 ( .A(y[1303]), .B(x[1303]), .Z(n32750) );
  AND U23404 ( .A(n32743), .B(n32750), .Z(n53354) );
  ANDN U23405 ( .B(y[1302]), .A(x[1302]), .Z(n32746) );
  NANDN U23406 ( .A(x[1301]), .B(y[1301]), .Z(n32739) );
  NANDN U23407 ( .A(n32746), .B(n32739), .Z(n53353) );
  ANDN U23408 ( .B(x[1300]), .A(y[1300]), .Z(n32735) );
  NANDN U23409 ( .A(y[1301]), .B(x[1301]), .Z(n32744) );
  NANDN U23410 ( .A(n32735), .B(n32744), .Z(n52306) );
  NANDN U23411 ( .A(x[1299]), .B(y[1299]), .Z(n32731) );
  ANDN U23412 ( .B(y[1300]), .A(x[1300]), .Z(n32741) );
  ANDN U23413 ( .B(n32731), .A(n32741), .Z(n53352) );
  NANDN U23414 ( .A(x[1295]), .B(y[1295]), .Z(n53348) );
  NANDN U23415 ( .A(x[1296]), .B(y[1296]), .Z(n52308) );
  NAND U23416 ( .A(n53348), .B(n52308), .Z(n12433) );
  ANDN U23417 ( .B(x[1294]), .A(y[1294]), .Z(n53347) );
  NANDN U23418 ( .A(x[1293]), .B(y[1293]), .Z(n27946) );
  NANDN U23419 ( .A(x[1294]), .B(y[1294]), .Z(n32721) );
  NAND U23420 ( .A(n27946), .B(n32721), .Z(n52310) );
  NANDN U23421 ( .A(y[1292]), .B(x[1292]), .Z(n32712) );
  ANDN U23422 ( .B(x[1293]), .A(y[1293]), .Z(n32719) );
  ANDN U23423 ( .B(n32712), .A(n32719), .Z(n53346) );
  NANDN U23424 ( .A(x[1292]), .B(y[1292]), .Z(n27947) );
  ANDN U23425 ( .B(y[1291]), .A(x[1291]), .Z(n32708) );
  ANDN U23426 ( .B(n27947), .A(n32708), .Z(n53345) );
  ANDN U23427 ( .B(x[1291]), .A(y[1291]), .Z(n32714) );
  NANDN U23428 ( .A(y[1290]), .B(x[1290]), .Z(n32704) );
  NANDN U23429 ( .A(n32714), .B(n32704), .Z(n53344) );
  NANDN U23430 ( .A(x[1289]), .B(y[1289]), .Z(n27948) );
  ANDN U23431 ( .B(y[1290]), .A(x[1290]), .Z(n32710) );
  ANDN U23432 ( .B(n27948), .A(n32710), .Z(n53343) );
  NANDN U23433 ( .A(y[1288]), .B(x[1288]), .Z(n27950) );
  NANDN U23434 ( .A(y[1289]), .B(x[1289]), .Z(n32703) );
  NAND U23435 ( .A(n27950), .B(n32703), .Z(n53342) );
  NANDN U23436 ( .A(x[1288]), .B(y[1288]), .Z(n27949) );
  ANDN U23437 ( .B(y[1287]), .A(x[1287]), .Z(n32696) );
  ANDN U23438 ( .B(n27949), .A(n32696), .Z(n53341) );
  NANDN U23439 ( .A(y[1286]), .B(x[1286]), .Z(n32692) );
  NANDN U23440 ( .A(y[1287]), .B(x[1287]), .Z(n27951) );
  NAND U23441 ( .A(n32692), .B(n27951), .Z(n53340) );
  NANDN U23442 ( .A(x[1285]), .B(y[1285]), .Z(n27952) );
  ANDN U23443 ( .B(y[1286]), .A(x[1286]), .Z(n32697) );
  ANDN U23444 ( .B(n27952), .A(n32697), .Z(n53339) );
  NANDN U23445 ( .A(y[1284]), .B(x[1284]), .Z(n27954) );
  NANDN U23446 ( .A(y[1285]), .B(x[1285]), .Z(n32691) );
  NAND U23447 ( .A(n27954), .B(n32691), .Z(n53338) );
  NANDN U23448 ( .A(x[1284]), .B(y[1284]), .Z(n27953) );
  ANDN U23449 ( .B(y[1283]), .A(x[1283]), .Z(n32684) );
  ANDN U23450 ( .B(n27953), .A(n32684), .Z(n53337) );
  NANDN U23451 ( .A(y[1282]), .B(x[1282]), .Z(n32680) );
  NANDN U23452 ( .A(y[1283]), .B(x[1283]), .Z(n27955) );
  NAND U23453 ( .A(n32680), .B(n27955), .Z(n53336) );
  ANDN U23454 ( .B(y[1281]), .A(x[1281]), .Z(n27957) );
  ANDN U23455 ( .B(y[1282]), .A(x[1282]), .Z(n32685) );
  NOR U23456 ( .A(n27957), .B(n32685), .Z(n53334) );
  ANDN U23457 ( .B(x[1280]), .A(y[1280]), .Z(n32674) );
  NANDN U23458 ( .A(y[1281]), .B(x[1281]), .Z(n32679) );
  NANDN U23459 ( .A(n32674), .B(n32679), .Z(n53333) );
  NANDN U23460 ( .A(x[1279]), .B(y[1279]), .Z(n32670) );
  ANDN U23461 ( .B(y[1280]), .A(x[1280]), .Z(n27956) );
  ANDN U23462 ( .B(n32670), .A(n27956), .Z(n53332) );
  ANDN U23463 ( .B(x[1278]), .A(y[1278]), .Z(n32669) );
  ANDN U23464 ( .B(x[1279]), .A(y[1279]), .Z(n32675) );
  OR U23465 ( .A(n32669), .B(n32675), .Z(n53331) );
  NANDN U23466 ( .A(x[1278]), .B(y[1278]), .Z(n53330) );
  ANDN U23467 ( .B(x[1277]), .A(y[1277]), .Z(n53329) );
  NANDN U23468 ( .A(x[1276]), .B(y[1276]), .Z(n27959) );
  ANDN U23469 ( .B(x[1274]), .A(y[1274]), .Z(n53325) );
  NANDN U23470 ( .A(x[1274]), .B(y[1274]), .Z(n32662) );
  NANDN U23471 ( .A(x[1273]), .B(y[1273]), .Z(n10225) );
  AND U23472 ( .A(n32662), .B(n10225), .Z(n53324) );
  NANDN U23473 ( .A(y[1272]), .B(x[1272]), .Z(n32652) );
  NANDN U23474 ( .A(y[1273]), .B(x[1273]), .Z(n32660) );
  AND U23475 ( .A(n32652), .B(n32660), .Z(n53323) );
  ANDN U23476 ( .B(y[1271]), .A(x[1271]), .Z(n32650) );
  NANDN U23477 ( .A(x[1272]), .B(y[1272]), .Z(n32655) );
  NANDN U23478 ( .A(n32650), .B(n32655), .Z(n53322) );
  NANDN U23479 ( .A(y[1270]), .B(x[1270]), .Z(n32645) );
  NANDN U23480 ( .A(y[1271]), .B(x[1271]), .Z(n32653) );
  AND U23481 ( .A(n32645), .B(n32653), .Z(n52311) );
  ANDN U23482 ( .B(y[1270]), .A(x[1270]), .Z(n53321) );
  NANDN U23483 ( .A(y[1269]), .B(x[1269]), .Z(n53320) );
  NANDN U23484 ( .A(y[1268]), .B(x[1268]), .Z(n27965) );
  NANDN U23485 ( .A(x[1267]), .B(y[1267]), .Z(n27967) );
  XNOR U23486 ( .A(y[1267]), .B(x[1267]), .Z(n12395) );
  NANDN U23487 ( .A(y[1266]), .B(x[1266]), .Z(n27969) );
  NANDN U23488 ( .A(y[1265]), .B(x[1265]), .Z(n27968) );
  NANDN U23489 ( .A(y[1264]), .B(x[1264]), .Z(n53313) );
  AND U23490 ( .A(n27968), .B(n53313), .Z(n12390) );
  NANDN U23491 ( .A(x[1263]), .B(y[1263]), .Z(n32633) );
  ANDN U23492 ( .B(y[1264]), .A(x[1264]), .Z(n32640) );
  ANDN U23493 ( .B(n32633), .A(n32640), .Z(n53312) );
  ANDN U23494 ( .B(x[1262]), .A(y[1262]), .Z(n32629) );
  NANDN U23495 ( .A(y[1263]), .B(x[1263]), .Z(n27970) );
  NANDN U23496 ( .A(n32629), .B(n27970), .Z(n53311) );
  NANDN U23497 ( .A(x[1261]), .B(y[1261]), .Z(n32625) );
  ANDN U23498 ( .B(y[1262]), .A(x[1262]), .Z(n32635) );
  ANDN U23499 ( .B(n32625), .A(n32635), .Z(n53310) );
  ANDN U23500 ( .B(x[1261]), .A(y[1261]), .Z(n32631) );
  NANDN U23501 ( .A(y[1260]), .B(x[1260]), .Z(n27971) );
  NANDN U23502 ( .A(n32631), .B(n27971), .Z(n53309) );
  NANDN U23503 ( .A(x[1259]), .B(y[1259]), .Z(n27973) );
  NANDN U23504 ( .A(x[1260]), .B(y[1260]), .Z(n32624) );
  AND U23505 ( .A(n27973), .B(n32624), .Z(n53308) );
  ANDN U23506 ( .B(x[1258]), .A(y[1258]), .Z(n32617) );
  NANDN U23507 ( .A(y[1259]), .B(x[1259]), .Z(n27972) );
  NANDN U23508 ( .A(n32617), .B(n27972), .Z(n53307) );
  NANDN U23509 ( .A(x[1257]), .B(y[1257]), .Z(n32613) );
  NANDN U23510 ( .A(x[1258]), .B(y[1258]), .Z(n27974) );
  AND U23511 ( .A(n32613), .B(n27974), .Z(n53306) );
  ANDN U23512 ( .B(x[1256]), .A(y[1256]), .Z(n27976) );
  ANDN U23513 ( .B(x[1257]), .A(y[1257]), .Z(n32618) );
  OR U23514 ( .A(n27976), .B(n32618), .Z(n53305) );
  NANDN U23515 ( .A(x[1256]), .B(y[1256]), .Z(n32612) );
  ANDN U23516 ( .B(y[1255]), .A(x[1255]), .Z(n32607) );
  ANDN U23517 ( .B(n32612), .A(n32607), .Z(n53304) );
  ANDN U23518 ( .B(y[1253]), .A(x[1253]), .Z(n32599) );
  ANDN U23519 ( .B(y[1254]), .A(x[1254]), .Z(n32608) );
  NOR U23520 ( .A(n32599), .B(n32608), .Z(n53303) );
  NANDN U23521 ( .A(y[1252]), .B(x[1252]), .Z(n32597) );
  NANDN U23522 ( .A(y[1253]), .B(x[1253]), .Z(n32602) );
  NAND U23523 ( .A(n32597), .B(n32602), .Z(n52313) );
  NANDN U23524 ( .A(x[1252]), .B(y[1252]), .Z(n27977) );
  NANDN U23525 ( .A(x[1251]), .B(y[1251]), .Z(n27978) );
  NANDN U23526 ( .A(y[1250]), .B(x[1250]), .Z(n53298) );
  NANDN U23527 ( .A(y[1251]), .B(x[1251]), .Z(n53300) );
  NAND U23528 ( .A(n53298), .B(n53300), .Z(n12374) );
  NANDN U23529 ( .A(y[1248]), .B(x[1248]), .Z(n32588) );
  NANDN U23530 ( .A(y[1249]), .B(x[1249]), .Z(n32593) );
  NAND U23531 ( .A(n32588), .B(n32593), .Z(n53296) );
  ANDN U23532 ( .B(y[1247]), .A(x[1247]), .Z(n32586) );
  ANDN U23533 ( .B(y[1248]), .A(x[1248]), .Z(n32591) );
  NOR U23534 ( .A(n32586), .B(n32591), .Z(n53295) );
  NANDN U23535 ( .A(y[1247]), .B(x[1247]), .Z(n10227) );
  NANDN U23536 ( .A(y[1246]), .B(x[1246]), .Z(n10226) );
  AND U23537 ( .A(n10227), .B(n10226), .Z(n53294) );
  NANDN U23538 ( .A(y[1245]), .B(x[1245]), .Z(n32580) );
  NANDN U23539 ( .A(y[1244]), .B(x[1244]), .Z(n10228) );
  AND U23540 ( .A(n32580), .B(n10228), .Z(n12365) );
  ANDN U23541 ( .B(y[1244]), .A(x[1244]), .Z(n32581) );
  NANDN U23542 ( .A(x[1243]), .B(y[1243]), .Z(n27980) );
  NANDN U23543 ( .A(n32581), .B(n27980), .Z(n10229) );
  NAND U23544 ( .A(n12365), .B(n10229), .Z(n10232) );
  NANDN U23545 ( .A(x[1246]), .B(y[1246]), .Z(n10231) );
  NANDN U23546 ( .A(x[1245]), .B(y[1245]), .Z(n10230) );
  NAND U23547 ( .A(n10231), .B(n10230), .Z(n32579) );
  ANDN U23548 ( .B(n10232), .A(n32579), .Z(n53293) );
  NANDN U23549 ( .A(y[1242]), .B(x[1242]), .Z(n27982) );
  NANDN U23550 ( .A(x[1241]), .B(y[1241]), .Z(n32571) );
  NANDN U23551 ( .A(y[1240]), .B(x[1240]), .Z(n27984) );
  NANDN U23552 ( .A(x[1239]), .B(y[1239]), .Z(n32568) );
  NANDN U23553 ( .A(x[1240]), .B(y[1240]), .Z(n32572) );
  ANDN U23554 ( .B(x[1238]), .A(y[1238]), .Z(n32562) );
  ANDN U23555 ( .B(y[1237]), .A(x[1237]), .Z(n32558) );
  ANDN U23556 ( .B(y[1238]), .A(x[1238]), .Z(n32567) );
  NOR U23557 ( .A(n32558), .B(n32567), .Z(n53285) );
  XNOR U23558 ( .A(x[1236]), .B(y[1236]), .Z(n10233) );
  ANDN U23559 ( .B(y[1235]), .A(x[1235]), .Z(n32551) );
  ANDN U23560 ( .B(n10233), .A(n32551), .Z(n53283) );
  NANDN U23561 ( .A(y[1234]), .B(x[1234]), .Z(n32547) );
  NANDN U23562 ( .A(y[1235]), .B(x[1235]), .Z(n32556) );
  NAND U23563 ( .A(n32547), .B(n32556), .Z(n52314) );
  NANDN U23564 ( .A(x[1233]), .B(y[1233]), .Z(n27985) );
  ANDN U23565 ( .B(y[1234]), .A(x[1234]), .Z(n32553) );
  ANDN U23566 ( .B(n27985), .A(n32553), .Z(n53281) );
  NANDN U23567 ( .A(y[1232]), .B(x[1232]), .Z(n27987) );
  NANDN U23568 ( .A(y[1233]), .B(x[1233]), .Z(n32546) );
  NAND U23569 ( .A(n27987), .B(n32546), .Z(n52315) );
  NANDN U23570 ( .A(x[1232]), .B(y[1232]), .Z(n27986) );
  ANDN U23571 ( .B(y[1231]), .A(x[1231]), .Z(n32539) );
  ANDN U23572 ( .B(n27986), .A(n32539), .Z(n53280) );
  NANDN U23573 ( .A(x[1229]), .B(y[1229]), .Z(n27989) );
  ANDN U23574 ( .B(y[1230]), .A(x[1230]), .Z(n32540) );
  ANDN U23575 ( .B(n27989), .A(n32540), .Z(n53278) );
  NANDN U23576 ( .A(y[1228]), .B(x[1228]), .Z(n32529) );
  NANDN U23577 ( .A(y[1229]), .B(x[1229]), .Z(n32537) );
  NAND U23578 ( .A(n32529), .B(n32537), .Z(n53277) );
  NANDN U23579 ( .A(x[1228]), .B(y[1228]), .Z(n27990) );
  ANDN U23580 ( .B(y[1227]), .A(x[1227]), .Z(n32527) );
  ANDN U23581 ( .B(n27990), .A(n32527), .Z(n53276) );
  ANDN U23582 ( .B(x[1227]), .A(y[1227]), .Z(n32531) );
  NANDN U23583 ( .A(y[1226]), .B(x[1226]), .Z(n32522) );
  NANDN U23584 ( .A(n32531), .B(n32522), .Z(n53275) );
  ANDN U23585 ( .B(y[1226]), .A(x[1226]), .Z(n53274) );
  NANDN U23586 ( .A(y[1224]), .B(x[1224]), .Z(n53272) );
  NANDN U23587 ( .A(y[1225]), .B(x[1225]), .Z(n52316) );
  NAND U23588 ( .A(n53272), .B(n52316), .Z(n12340) );
  ANDN U23589 ( .B(y[1223]), .A(x[1223]), .Z(n53270) );
  ANDN U23590 ( .B(x[1222]), .A(y[1222]), .Z(n32513) );
  NANDN U23591 ( .A(y[1223]), .B(x[1223]), .Z(n27993) );
  NANDN U23592 ( .A(n32513), .B(n27993), .Z(n53269) );
  NANDN U23593 ( .A(x[1221]), .B(y[1221]), .Z(n32509) );
  NANDN U23594 ( .A(x[1222]), .B(y[1222]), .Z(n32517) );
  AND U23595 ( .A(n32509), .B(n32517), .Z(n53268) );
  ANDN U23596 ( .B(x[1220]), .A(y[1220]), .Z(n32504) );
  ANDN U23597 ( .B(x[1221]), .A(y[1221]), .Z(n32515) );
  OR U23598 ( .A(n32504), .B(n32515), .Z(n53267) );
  NANDN U23599 ( .A(x[1219]), .B(y[1219]), .Z(n32502) );
  NANDN U23600 ( .A(x[1220]), .B(y[1220]), .Z(n32508) );
  AND U23601 ( .A(n32502), .B(n32508), .Z(n53266) );
  ANDN U23602 ( .B(x[1218]), .A(y[1218]), .Z(n32499) );
  ANDN U23603 ( .B(x[1219]), .A(y[1219]), .Z(n32507) );
  OR U23604 ( .A(n32499), .B(n32507), .Z(n53265) );
  NANDN U23605 ( .A(x[1218]), .B(y[1218]), .Z(n53264) );
  ANDN U23606 ( .B(x[1217]), .A(y[1217]), .Z(n53263) );
  NANDN U23607 ( .A(x[1216]), .B(y[1216]), .Z(n27995) );
  NANDN U23608 ( .A(y[1215]), .B(x[1215]), .Z(n27997) );
  ANDN U23609 ( .B(x[1214]), .A(y[1214]), .Z(n28000) );
  ANDN U23610 ( .B(n27997), .A(n28000), .Z(n12325) );
  ANDN U23611 ( .B(y[1213]), .A(x[1213]), .Z(n28003) );
  NANDN U23612 ( .A(y[1213]), .B(x[1213]), .Z(n28001) );
  NANDN U23613 ( .A(x[1211]), .B(y[1211]), .Z(n32484) );
  NANDN U23614 ( .A(x[1212]), .B(y[1212]), .Z(n32492) );
  NAND U23615 ( .A(n32484), .B(n32492), .Z(n53256) );
  ANDN U23616 ( .B(x[1210]), .A(y[1210]), .Z(n32479) );
  ANDN U23617 ( .B(x[1211]), .A(y[1211]), .Z(n32488) );
  NOR U23618 ( .A(n32479), .B(n32488), .Z(n53255) );
  ANDN U23619 ( .B(x[1208]), .A(y[1208]), .Z(n32472) );
  ANDN U23620 ( .B(x[1209]), .A(y[1209]), .Z(n32482) );
  NOR U23621 ( .A(n32472), .B(n32482), .Z(n53254) );
  NANDN U23622 ( .A(x[1207]), .B(y[1207]), .Z(n32468) );
  XNOR U23623 ( .A(x[1208]), .B(y[1208]), .Z(n10234) );
  NAND U23624 ( .A(n32468), .B(n10234), .Z(n52319) );
  ANDN U23625 ( .B(x[1206]), .A(y[1206]), .Z(n28005) );
  ANDN U23626 ( .B(x[1207]), .A(y[1207]), .Z(n32474) );
  NOR U23627 ( .A(n28005), .B(n32474), .Z(n53251) );
  ANDN U23628 ( .B(y[1205]), .A(x[1205]), .Z(n32462) );
  NANDN U23629 ( .A(x[1206]), .B(y[1206]), .Z(n32467) );
  NANDN U23630 ( .A(n32462), .B(n32467), .Z(n53250) );
  NANDN U23631 ( .A(y[1204]), .B(x[1204]), .Z(n32458) );
  ANDN U23632 ( .B(x[1205]), .A(y[1205]), .Z(n28004) );
  ANDN U23633 ( .B(n32458), .A(n28004), .Z(n53249) );
  ANDN U23634 ( .B(y[1203]), .A(x[1203]), .Z(n32456) );
  ANDN U23635 ( .B(y[1204]), .A(x[1204]), .Z(n32463) );
  NOR U23636 ( .A(n32456), .B(n32463), .Z(n53248) );
  NANDN U23637 ( .A(y[1202]), .B(x[1202]), .Z(n10235) );
  NANDN U23638 ( .A(y[1203]), .B(x[1203]), .Z(n32457) );
  NAND U23639 ( .A(n10235), .B(n32457), .Z(n53247) );
  NANDN U23640 ( .A(y[1200]), .B(x[1200]), .Z(n32446) );
  NANDN U23641 ( .A(y[1201]), .B(x[1201]), .Z(n32452) );
  NAND U23642 ( .A(n32446), .B(n32452), .Z(n53244) );
  ANDN U23643 ( .B(y[1199]), .A(x[1199]), .Z(n32443) );
  ANDN U23644 ( .B(y[1200]), .A(x[1200]), .Z(n32449) );
  NOR U23645 ( .A(n32443), .B(n32449), .Z(n53243) );
  NANDN U23646 ( .A(y[1199]), .B(x[1199]), .Z(n28006) );
  NANDN U23647 ( .A(y[1198]), .B(x[1198]), .Z(n10236) );
  AND U23648 ( .A(n28006), .B(n10236), .Z(n52321) );
  NANDN U23649 ( .A(y[1196]), .B(x[1196]), .Z(n10237) );
  NANDN U23650 ( .A(y[1197]), .B(x[1197]), .Z(n28008) );
  AND U23651 ( .A(n10237), .B(n28008), .Z(n53242) );
  ANDN U23652 ( .B(y[1195]), .A(x[1195]), .Z(n28010) );
  XNOR U23653 ( .A(y[1196]), .B(x[1196]), .Z(n32434) );
  NANDN U23654 ( .A(n28010), .B(n32434), .Z(n53241) );
  ANDN U23655 ( .B(x[1194]), .A(y[1194]), .Z(n32428) );
  NANDN U23656 ( .A(y[1195]), .B(x[1195]), .Z(n32433) );
  NANDN U23657 ( .A(n32428), .B(n32433), .Z(n52323) );
  NANDN U23658 ( .A(x[1193]), .B(y[1193]), .Z(n32424) );
  ANDN U23659 ( .B(y[1194]), .A(x[1194]), .Z(n28009) );
  ANDN U23660 ( .B(n32424), .A(n28009), .Z(n53238) );
  NANDN U23661 ( .A(x[1189]), .B(y[1189]), .Z(n28012) );
  NANDN U23662 ( .A(x[1190]), .B(y[1190]), .Z(n52325) );
  AND U23663 ( .A(n28012), .B(n52325), .Z(n12293) );
  ANDN U23664 ( .B(x[1189]), .A(y[1189]), .Z(n32413) );
  NANDN U23665 ( .A(y[1188]), .B(x[1188]), .Z(n28013) );
  NANDN U23666 ( .A(x[1187]), .B(y[1187]), .Z(n53232) );
  NANDN U23667 ( .A(y[1187]), .B(x[1187]), .Z(n28014) );
  ANDN U23668 ( .B(y[1185]), .A(x[1185]), .Z(n32404) );
  NANDN U23669 ( .A(x[1186]), .B(y[1186]), .Z(n32409) );
  NANDN U23670 ( .A(n32404), .B(n32409), .Z(n53230) );
  NANDN U23671 ( .A(y[1184]), .B(x[1184]), .Z(n28015) );
  NANDN U23672 ( .A(y[1185]), .B(x[1185]), .Z(n32406) );
  AND U23673 ( .A(n28015), .B(n32406), .Z(n53229) );
  NANDN U23674 ( .A(x[1183]), .B(y[1183]), .Z(n32396) );
  ANDN U23675 ( .B(y[1184]), .A(x[1184]), .Z(n32401) );
  ANDN U23676 ( .B(n32396), .A(n32401), .Z(n53228) );
  ANDN U23677 ( .B(x[1182]), .A(y[1182]), .Z(n32392) );
  NANDN U23678 ( .A(y[1183]), .B(x[1183]), .Z(n28016) );
  NANDN U23679 ( .A(n32392), .B(n28016), .Z(n52326) );
  NANDN U23680 ( .A(x[1181]), .B(y[1181]), .Z(n32388) );
  ANDN U23681 ( .B(y[1182]), .A(x[1182]), .Z(n32398) );
  ANDN U23682 ( .B(n32388), .A(n32398), .Z(n53227) );
  ANDN U23683 ( .B(x[1181]), .A(y[1181]), .Z(n32394) );
  NANDN U23684 ( .A(y[1180]), .B(x[1180]), .Z(n10238) );
  NANDN U23685 ( .A(n32394), .B(n10238), .Z(n53225) );
  XNOR U23686 ( .A(y[1180]), .B(x[1180]), .Z(n28018) );
  NANDN U23687 ( .A(x[1179]), .B(y[1179]), .Z(n28019) );
  AND U23688 ( .A(n28018), .B(n28019), .Z(n53224) );
  ANDN U23689 ( .B(x[1178]), .A(y[1178]), .Z(n32380) );
  NANDN U23690 ( .A(y[1179]), .B(x[1179]), .Z(n28017) );
  NANDN U23691 ( .A(n32380), .B(n28017), .Z(n53223) );
  NANDN U23692 ( .A(x[1177]), .B(y[1177]), .Z(n32376) );
  NANDN U23693 ( .A(x[1178]), .B(y[1178]), .Z(n28020) );
  AND U23694 ( .A(n32376), .B(n28020), .Z(n53222) );
  ANDN U23695 ( .B(x[1177]), .A(y[1177]), .Z(n32381) );
  NANDN U23696 ( .A(y[1176]), .B(x[1176]), .Z(n28022) );
  NANDN U23697 ( .A(n32381), .B(n28022), .Z(n53221) );
  NANDN U23698 ( .A(x[1176]), .B(y[1176]), .Z(n32375) );
  ANDN U23699 ( .B(y[1175]), .A(x[1175]), .Z(n32371) );
  ANDN U23700 ( .B(n32375), .A(n32371), .Z(n53220) );
  NANDN U23701 ( .A(y[1174]), .B(x[1174]), .Z(n32367) );
  NANDN U23702 ( .A(y[1175]), .B(x[1175]), .Z(n28021) );
  NAND U23703 ( .A(n32367), .B(n28021), .Z(n53219) );
  NANDN U23704 ( .A(x[1173]), .B(y[1173]), .Z(n28023) );
  ANDN U23705 ( .B(y[1174]), .A(x[1174]), .Z(n53218) );
  ANDN U23706 ( .B(n28023), .A(n53218), .Z(n12273) );
  NANDN U23707 ( .A(y[1173]), .B(x[1173]), .Z(n53217) );
  NANDN U23708 ( .A(x[1172]), .B(y[1172]), .Z(n28024) );
  NANDN U23709 ( .A(y[1170]), .B(x[1170]), .Z(n32358) );
  NANDN U23710 ( .A(y[1171]), .B(x[1171]), .Z(n28025) );
  NAND U23711 ( .A(n32358), .B(n28025), .Z(n53213) );
  XNOR U23712 ( .A(x[1170]), .B(y[1170]), .Z(n10239) );
  ANDN U23713 ( .B(y[1169]), .A(x[1169]), .Z(n28027) );
  ANDN U23714 ( .B(n10239), .A(n28027), .Z(n53212) );
  NANDN U23715 ( .A(y[1169]), .B(x[1169]), .Z(n32357) );
  ANDN U23716 ( .B(x[1168]), .A(y[1168]), .Z(n32352) );
  ANDN U23717 ( .B(n32357), .A(n32352), .Z(n53211) );
  ANDN U23718 ( .B(y[1168]), .A(x[1168]), .Z(n28026) );
  NANDN U23719 ( .A(x[1167]), .B(y[1167]), .Z(n32348) );
  NANDN U23720 ( .A(n28026), .B(n32348), .Z(n52327) );
  ANDN U23721 ( .B(x[1166]), .A(y[1166]), .Z(n32344) );
  ANDN U23722 ( .B(x[1167]), .A(y[1167]), .Z(n32353) );
  NOR U23723 ( .A(n32344), .B(n32353), .Z(n53210) );
  NANDN U23724 ( .A(y[1164]), .B(x[1164]), .Z(n28030) );
  NANDN U23725 ( .A(y[1165]), .B(x[1165]), .Z(n28028) );
  AND U23726 ( .A(n28030), .B(n28028), .Z(n12260) );
  ANDN U23727 ( .B(y[1163]), .A(x[1163]), .Z(n28031) );
  NANDN U23728 ( .A(x[1164]), .B(y[1164]), .Z(n53206) );
  ANDN U23729 ( .B(x[1162]), .A(y[1162]), .Z(n53203) );
  ANDN U23730 ( .B(x[1160]), .A(y[1160]), .Z(n32330) );
  ANDN U23731 ( .B(x[1161]), .A(y[1161]), .Z(n32336) );
  NOR U23732 ( .A(n32330), .B(n32336), .Z(n53201) );
  NANDN U23733 ( .A(x[1159]), .B(y[1159]), .Z(n32326) );
  NANDN U23734 ( .A(x[1160]), .B(y[1160]), .Z(n32334) );
  NAND U23735 ( .A(n32326), .B(n32334), .Z(n52329) );
  ANDN U23736 ( .B(x[1159]), .A(y[1159]), .Z(n32332) );
  NANDN U23737 ( .A(y[1158]), .B(x[1158]), .Z(n28034) );
  NANDN U23738 ( .A(n32332), .B(n28034), .Z(n53200) );
  NANDN U23739 ( .A(x[1157]), .B(y[1157]), .Z(n28036) );
  NANDN U23740 ( .A(x[1158]), .B(y[1158]), .Z(n32325) );
  AND U23741 ( .A(n28036), .B(n32325), .Z(n53199) );
  ANDN U23742 ( .B(x[1156]), .A(y[1156]), .Z(n32318) );
  NANDN U23743 ( .A(y[1157]), .B(x[1157]), .Z(n28035) );
  NANDN U23744 ( .A(n32318), .B(n28035), .Z(n53198) );
  NANDN U23745 ( .A(x[1155]), .B(y[1155]), .Z(n32314) );
  NANDN U23746 ( .A(x[1156]), .B(y[1156]), .Z(n28037) );
  AND U23747 ( .A(n32314), .B(n28037), .Z(n53197) );
  ANDN U23748 ( .B(x[1155]), .A(y[1155]), .Z(n32319) );
  NANDN U23749 ( .A(y[1154]), .B(x[1154]), .Z(n28038) );
  NANDN U23750 ( .A(n32319), .B(n28038), .Z(n53196) );
  NANDN U23751 ( .A(x[1153]), .B(y[1153]), .Z(n28040) );
  NANDN U23752 ( .A(x[1154]), .B(y[1154]), .Z(n32313) );
  AND U23753 ( .A(n28040), .B(n32313), .Z(n53195) );
  ANDN U23754 ( .B(x[1152]), .A(y[1152]), .Z(n32306) );
  NANDN U23755 ( .A(y[1153]), .B(x[1153]), .Z(n28039) );
  NANDN U23756 ( .A(n32306), .B(n28039), .Z(n53194) );
  NANDN U23757 ( .A(x[1151]), .B(y[1151]), .Z(n32302) );
  NANDN U23758 ( .A(x[1152]), .B(y[1152]), .Z(n28041) );
  AND U23759 ( .A(n32302), .B(n28041), .Z(n53193) );
  ANDN U23760 ( .B(x[1151]), .A(y[1151]), .Z(n32307) );
  NANDN U23761 ( .A(y[1150]), .B(x[1150]), .Z(n28043) );
  NANDN U23762 ( .A(n32307), .B(n28043), .Z(n53192) );
  NANDN U23763 ( .A(x[1150]), .B(y[1150]), .Z(n32301) );
  ANDN U23764 ( .B(y[1149]), .A(x[1149]), .Z(n32297) );
  ANDN U23765 ( .B(n32301), .A(n32297), .Z(n53191) );
  NANDN U23766 ( .A(y[1148]), .B(x[1148]), .Z(n32293) );
  NANDN U23767 ( .A(y[1149]), .B(x[1149]), .Z(n28042) );
  NAND U23768 ( .A(n32293), .B(n28042), .Z(n53190) );
  NANDN U23769 ( .A(x[1146]), .B(y[1146]), .Z(n28045) );
  ANDN U23770 ( .B(y[1145]), .A(x[1145]), .Z(n53184) );
  ANDN U23771 ( .B(n28045), .A(n53184), .Z(n12235) );
  NANDN U23772 ( .A(y[1144]), .B(x[1144]), .Z(n32283) );
  NANDN U23773 ( .A(y[1145]), .B(x[1145]), .Z(n32289) );
  AND U23774 ( .A(n32283), .B(n32289), .Z(n53183) );
  ANDN U23775 ( .B(y[1143]), .A(x[1143]), .Z(n32279) );
  ANDN U23776 ( .B(y[1144]), .A(x[1144]), .Z(n32286) );
  OR U23777 ( .A(n32279), .B(n32286), .Z(n53182) );
  NANDN U23778 ( .A(y[1142]), .B(x[1142]), .Z(n10240) );
  NANDN U23779 ( .A(y[1143]), .B(x[1143]), .Z(n32284) );
  AND U23780 ( .A(n10240), .B(n32284), .Z(n52330) );
  XNOR U23781 ( .A(y[1140]), .B(x[1140]), .Z(n32269) );
  NANDN U23782 ( .A(x[1139]), .B(y[1139]), .Z(n32265) );
  NAND U23783 ( .A(n32269), .B(n32265), .Z(n52333) );
  NANDN U23784 ( .A(y[1139]), .B(x[1139]), .Z(n32268) );
  ANDN U23785 ( .B(x[1138]), .A(y[1138]), .Z(n32263) );
  ANDN U23786 ( .B(n32268), .A(n32263), .Z(n53181) );
  NANDN U23787 ( .A(x[1137]), .B(y[1137]), .Z(n28048) );
  NANDN U23788 ( .A(x[1138]), .B(y[1138]), .Z(n32266) );
  NAND U23789 ( .A(n28048), .B(n32266), .Z(n53178) );
  NANDN U23790 ( .A(y[1136]), .B(x[1136]), .Z(n32255) );
  ANDN U23791 ( .B(x[1137]), .A(y[1137]), .Z(n32260) );
  ANDN U23792 ( .B(n32255), .A(n32260), .Z(n53177) );
  NANDN U23793 ( .A(y[1134]), .B(x[1134]), .Z(n32247) );
  ANDN U23794 ( .B(x[1135]), .A(y[1135]), .Z(n32257) );
  ANDN U23795 ( .B(n32247), .A(n32257), .Z(n53176) );
  ANDN U23796 ( .B(y[1134]), .A(x[1134]), .Z(n32253) );
  NANDN U23797 ( .A(x[1133]), .B(y[1133]), .Z(n28050) );
  NANDN U23798 ( .A(n32253), .B(n28050), .Z(n52335) );
  NANDN U23799 ( .A(y[1132]), .B(x[1132]), .Z(n28052) );
  NANDN U23800 ( .A(y[1133]), .B(x[1133]), .Z(n32246) );
  AND U23801 ( .A(n28052), .B(n32246), .Z(n53175) );
  ANDN U23802 ( .B(y[1131]), .A(x[1131]), .Z(n32239) );
  NANDN U23803 ( .A(x[1132]), .B(y[1132]), .Z(n28051) );
  NANDN U23804 ( .A(n32239), .B(n28051), .Z(n53174) );
  NANDN U23805 ( .A(y[1130]), .B(x[1130]), .Z(n32235) );
  NANDN U23806 ( .A(y[1131]), .B(x[1131]), .Z(n28053) );
  AND U23807 ( .A(n32235), .B(n28053), .Z(n52336) );
  ANDN U23808 ( .B(y[1127]), .A(x[1127]), .Z(n32227) );
  NANDN U23809 ( .A(x[1128]), .B(y[1128]), .Z(n28055) );
  NANDN U23810 ( .A(n32227), .B(n28055), .Z(n52339) );
  NANDN U23811 ( .A(y[1126]), .B(x[1126]), .Z(n32223) );
  NANDN U23812 ( .A(y[1127]), .B(x[1127]), .Z(n28057) );
  AND U23813 ( .A(n32223), .B(n28057), .Z(n53172) );
  ANDN U23814 ( .B(y[1126]), .A(x[1126]), .Z(n32228) );
  NANDN U23815 ( .A(x[1125]), .B(y[1125]), .Z(n28058) );
  NANDN U23816 ( .A(n32228), .B(n28058), .Z(n53169) );
  NANDN U23817 ( .A(y[1124]), .B(x[1124]), .Z(n32217) );
  NANDN U23818 ( .A(y[1125]), .B(x[1125]), .Z(n32225) );
  AND U23819 ( .A(n32217), .B(n32225), .Z(n52340) );
  NANDN U23820 ( .A(y[1122]), .B(x[1122]), .Z(n32209) );
  ANDN U23821 ( .B(x[1123]), .A(y[1123]), .Z(n32219) );
  ANDN U23822 ( .B(n32209), .A(n32219), .Z(n53168) );
  NANDN U23823 ( .A(y[1121]), .B(x[1121]), .Z(n53166) );
  NANDN U23824 ( .A(y[1120]), .B(x[1120]), .Z(n53164) );
  AND U23825 ( .A(n53166), .B(n53164), .Z(n12207) );
  ANDN U23826 ( .B(y[1119]), .A(x[1119]), .Z(n53163) );
  NANDN U23827 ( .A(y[1118]), .B(x[1118]), .Z(n32200) );
  NANDN U23828 ( .A(y[1119]), .B(x[1119]), .Z(n28062) );
  AND U23829 ( .A(n32200), .B(n28062), .Z(n52342) );
  ANDN U23830 ( .B(y[1115]), .A(x[1115]), .Z(n32188) );
  XNOR U23831 ( .A(y[1116]), .B(x[1116]), .Z(n10241) );
  NANDN U23832 ( .A(n32188), .B(n10241), .Z(n52345) );
  NANDN U23833 ( .A(y[1114]), .B(x[1114]), .Z(n32184) );
  NANDN U23834 ( .A(y[1115]), .B(x[1115]), .Z(n32192) );
  AND U23835 ( .A(n32184), .B(n32192), .Z(n53160) );
  ANDN U23836 ( .B(y[1113]), .A(x[1113]), .Z(n32183) );
  ANDN U23837 ( .B(y[1114]), .A(x[1114]), .Z(n32190) );
  OR U23838 ( .A(n32183), .B(n32190), .Z(n53158) );
  NANDN U23839 ( .A(y[1113]), .B(x[1113]), .Z(n53156) );
  XOR U23840 ( .A(x[1112]), .B(y[1112]), .Z(n28063) );
  NANDN U23841 ( .A(y[1111]), .B(x[1111]), .Z(n28064) );
  ANDN U23842 ( .B(y[1109]), .A(x[1109]), .Z(n53146) );
  NANDN U23843 ( .A(y[1108]), .B(x[1108]), .Z(n32171) );
  NANDN U23844 ( .A(y[1109]), .B(x[1109]), .Z(n28067) );
  AND U23845 ( .A(n32171), .B(n28067), .Z(n53144) );
  ANDN U23846 ( .B(y[1107]), .A(x[1107]), .Z(n32166) );
  ANDN U23847 ( .B(y[1108]), .A(x[1108]), .Z(n32175) );
  OR U23848 ( .A(n32166), .B(n32175), .Z(n53142) );
  NANDN U23849 ( .A(y[1106]), .B(x[1106]), .Z(n32163) );
  NANDN U23850 ( .A(y[1107]), .B(x[1107]), .Z(n32170) );
  AND U23851 ( .A(n32163), .B(n32170), .Z(n53140) );
  ANDN U23852 ( .B(y[1106]), .A(x[1106]), .Z(n32169) );
  NANDN U23853 ( .A(x[1105]), .B(y[1105]), .Z(n32158) );
  NANDN U23854 ( .A(n32169), .B(n32158), .Z(n53138) );
  NANDN U23855 ( .A(y[1104]), .B(x[1104]), .Z(n28069) );
  NANDN U23856 ( .A(y[1105]), .B(x[1105]), .Z(n32164) );
  AND U23857 ( .A(n28069), .B(n32164), .Z(n53136) );
  ANDN U23858 ( .B(y[1103]), .A(x[1103]), .Z(n32153) );
  NANDN U23859 ( .A(x[1104]), .B(y[1104]), .Z(n32159) );
  NANDN U23860 ( .A(n32153), .B(n32159), .Z(n53134) );
  NANDN U23861 ( .A(y[1102]), .B(x[1102]), .Z(n32149) );
  NANDN U23862 ( .A(y[1103]), .B(x[1103]), .Z(n28068) );
  AND U23863 ( .A(n32149), .B(n28068), .Z(n53132) );
  ANDN U23864 ( .B(y[1101]), .A(x[1101]), .Z(n32144) );
  ANDN U23865 ( .B(y[1102]), .A(x[1102]), .Z(n32154) );
  OR U23866 ( .A(n32144), .B(n32154), .Z(n53130) );
  NANDN U23867 ( .A(y[1100]), .B(x[1100]), .Z(n32141) );
  NANDN U23868 ( .A(y[1101]), .B(x[1101]), .Z(n32148) );
  AND U23869 ( .A(n32141), .B(n32148), .Z(n53128) );
  ANDN U23870 ( .B(y[1100]), .A(x[1100]), .Z(n32147) );
  NANDN U23871 ( .A(x[1099]), .B(y[1099]), .Z(n32137) );
  NANDN U23872 ( .A(n32147), .B(n32137), .Z(n53126) );
  NANDN U23873 ( .A(y[1099]), .B(x[1099]), .Z(n32142) );
  ANDN U23874 ( .B(x[1098]), .A(y[1098]), .Z(n32133) );
  ANDN U23875 ( .B(n32142), .A(n32133), .Z(n53124) );
  ANDN U23876 ( .B(y[1098]), .A(x[1098]), .Z(n32139) );
  NANDN U23877 ( .A(x[1097]), .B(y[1097]), .Z(n32129) );
  NANDN U23878 ( .A(n32139), .B(n32129), .Z(n53122) );
  ANDN U23879 ( .B(x[1096]), .A(y[1096]), .Z(n32125) );
  ANDN U23880 ( .B(x[1097]), .A(y[1097]), .Z(n32135) );
  NOR U23881 ( .A(n32125), .B(n32135), .Z(n53120) );
  NANDN U23882 ( .A(x[1095]), .B(y[1095]), .Z(n32123) );
  NANDN U23883 ( .A(x[1096]), .B(y[1096]), .Z(n32128) );
  AND U23884 ( .A(n32123), .B(n32128), .Z(n53119) );
  ANDN U23885 ( .B(x[1094]), .A(y[1094]), .Z(n53117) );
  ANDN U23886 ( .B(x[1095]), .A(y[1095]), .Z(n53118) );
  OR U23887 ( .A(n53117), .B(n53118), .Z(n12174) );
  NANDN U23888 ( .A(x[1094]), .B(y[1094]), .Z(n52346) );
  NANDN U23889 ( .A(y[1092]), .B(x[1092]), .Z(n28070) );
  ANDN U23890 ( .B(x[1093]), .A(y[1093]), .Z(n32121) );
  ANDN U23891 ( .B(n28070), .A(n32121), .Z(n53115) );
  NANDN U23892 ( .A(x[1091]), .B(y[1091]), .Z(n28072) );
  NANDN U23893 ( .A(x[1092]), .B(y[1092]), .Z(n32116) );
  NAND U23894 ( .A(n28072), .B(n32116), .Z(n53114) );
  NANDN U23895 ( .A(y[1091]), .B(x[1091]), .Z(n28071) );
  ANDN U23896 ( .B(x[1090]), .A(y[1090]), .Z(n32109) );
  ANDN U23897 ( .B(n28071), .A(n32109), .Z(n53113) );
  NANDN U23898 ( .A(x[1089]), .B(y[1089]), .Z(n32105) );
  NANDN U23899 ( .A(x[1090]), .B(y[1090]), .Z(n28073) );
  AND U23900 ( .A(n32105), .B(n28073), .Z(n53112) );
  ANDN U23901 ( .B(x[1089]), .A(y[1089]), .Z(n32110) );
  NANDN U23902 ( .A(y[1088]), .B(x[1088]), .Z(n28074) );
  NANDN U23903 ( .A(n32110), .B(n28074), .Z(n53111) );
  NANDN U23904 ( .A(x[1087]), .B(y[1087]), .Z(n28076) );
  NANDN U23905 ( .A(x[1088]), .B(y[1088]), .Z(n32104) );
  AND U23906 ( .A(n28076), .B(n32104), .Z(n53110) );
  ANDN U23907 ( .B(x[1086]), .A(y[1086]), .Z(n32097) );
  NANDN U23908 ( .A(y[1087]), .B(x[1087]), .Z(n28075) );
  NANDN U23909 ( .A(n32097), .B(n28075), .Z(n53109) );
  NANDN U23910 ( .A(x[1085]), .B(y[1085]), .Z(n32093) );
  NANDN U23911 ( .A(x[1086]), .B(y[1086]), .Z(n28077) );
  AND U23912 ( .A(n32093), .B(n28077), .Z(n53108) );
  ANDN U23913 ( .B(x[1085]), .A(y[1085]), .Z(n32098) );
  NANDN U23914 ( .A(y[1084]), .B(x[1084]), .Z(n28078) );
  NANDN U23915 ( .A(n32098), .B(n28078), .Z(n53107) );
  NANDN U23916 ( .A(x[1083]), .B(y[1083]), .Z(n28080) );
  NANDN U23917 ( .A(x[1084]), .B(y[1084]), .Z(n32092) );
  AND U23918 ( .A(n28080), .B(n32092), .Z(n53106) );
  ANDN U23919 ( .B(x[1082]), .A(y[1082]), .Z(n32085) );
  NANDN U23920 ( .A(y[1083]), .B(x[1083]), .Z(n28079) );
  NANDN U23921 ( .A(n32085), .B(n28079), .Z(n53105) );
  NANDN U23922 ( .A(x[1081]), .B(y[1081]), .Z(n32081) );
  NANDN U23923 ( .A(x[1082]), .B(y[1082]), .Z(n28081) );
  AND U23924 ( .A(n32081), .B(n28081), .Z(n53104) );
  ANDN U23925 ( .B(x[1081]), .A(y[1081]), .Z(n32086) );
  NANDN U23926 ( .A(y[1080]), .B(x[1080]), .Z(n28082) );
  NANDN U23927 ( .A(n32086), .B(n28082), .Z(n53102) );
  NANDN U23928 ( .A(x[1079]), .B(y[1079]), .Z(n28084) );
  NANDN U23929 ( .A(x[1080]), .B(y[1080]), .Z(n32080) );
  AND U23930 ( .A(n28084), .B(n32080), .Z(n53101) );
  ANDN U23931 ( .B(x[1078]), .A(y[1078]), .Z(n32073) );
  NANDN U23932 ( .A(y[1079]), .B(x[1079]), .Z(n28083) );
  NANDN U23933 ( .A(n32073), .B(n28083), .Z(n53100) );
  NANDN U23934 ( .A(x[1077]), .B(y[1077]), .Z(n32069) );
  NANDN U23935 ( .A(x[1078]), .B(y[1078]), .Z(n28085) );
  AND U23936 ( .A(n32069), .B(n28085), .Z(n53099) );
  ANDN U23937 ( .B(x[1076]), .A(y[1076]), .Z(n28087) );
  ANDN U23938 ( .B(x[1077]), .A(y[1077]), .Z(n32074) );
  OR U23939 ( .A(n28087), .B(n32074), .Z(n53098) );
  NANDN U23940 ( .A(x[1076]), .B(y[1076]), .Z(n32068) );
  ANDN U23941 ( .B(y[1075]), .A(x[1075]), .Z(n32063) );
  ANDN U23942 ( .B(n32068), .A(n32063), .Z(n53097) );
  ANDN U23943 ( .B(x[1075]), .A(y[1075]), .Z(n28086) );
  NANDN U23944 ( .A(y[1074]), .B(x[1074]), .Z(n32059) );
  NANDN U23945 ( .A(n28086), .B(n32059), .Z(n53096) );
  ANDN U23946 ( .B(y[1073]), .A(x[1073]), .Z(n32055) );
  ANDN U23947 ( .B(y[1074]), .A(x[1074]), .Z(n32064) );
  NOR U23948 ( .A(n32055), .B(n32064), .Z(n53095) );
  NANDN U23949 ( .A(y[1072]), .B(x[1072]), .Z(n32053) );
  NANDN U23950 ( .A(y[1073]), .B(x[1073]), .Z(n32058) );
  NAND U23951 ( .A(n32053), .B(n32058), .Z(n53094) );
  NANDN U23952 ( .A(x[1070]), .B(y[1070]), .Z(n32050) );
  NANDN U23953 ( .A(x[1069]), .B(y[1069]), .Z(n28090) );
  AND U23954 ( .A(n32050), .B(n28090), .Z(n12145) );
  ANDN U23955 ( .B(x[1068]), .A(y[1068]), .Z(n28092) );
  NANDN U23956 ( .A(x[1068]), .B(y[1068]), .Z(n28091) );
  NANDN U23957 ( .A(y[1066]), .B(x[1066]), .Z(n32038) );
  NANDN U23958 ( .A(y[1067]), .B(x[1067]), .Z(n32045) );
  NAND U23959 ( .A(n32038), .B(n32045), .Z(n53086) );
  NANDN U23960 ( .A(x[1066]), .B(y[1066]), .Z(n28093) );
  NANDN U23961 ( .A(y[1064]), .B(x[1064]), .Z(n53081) );
  NANDN U23962 ( .A(y[1065]), .B(x[1065]), .Z(n53083) );
  NAND U23963 ( .A(n53081), .B(n53083), .Z(n12136) );
  ANDN U23964 ( .B(y[1063]), .A(x[1063]), .Z(n53080) );
  NANDN U23965 ( .A(y[1063]), .B(x[1063]), .Z(n28096) );
  ANDN U23966 ( .B(x[1062]), .A(y[1062]), .Z(n32029) );
  ANDN U23967 ( .B(n28096), .A(n32029), .Z(n53079) );
  NANDN U23968 ( .A(x[1061]), .B(y[1061]), .Z(n32025) );
  NANDN U23969 ( .A(x[1062]), .B(y[1062]), .Z(n32033) );
  NAND U23970 ( .A(n32025), .B(n32033), .Z(n52347) );
  ANDN U23971 ( .B(x[1060]), .A(y[1060]), .Z(n32020) );
  ANDN U23972 ( .B(x[1061]), .A(y[1061]), .Z(n32031) );
  NOR U23973 ( .A(n32020), .B(n32031), .Z(n53078) );
  NANDN U23974 ( .A(y[1058]), .B(x[1058]), .Z(n32012) );
  ANDN U23975 ( .B(x[1059]), .A(y[1059]), .Z(n32023) );
  ANDN U23976 ( .B(n32012), .A(n32023), .Z(n53076) );
  NANDN U23977 ( .A(x[1057]), .B(y[1057]), .Z(n28098) );
  NANDN U23978 ( .A(x[1058]), .B(y[1058]), .Z(n32018) );
  NAND U23979 ( .A(n28098), .B(n32018), .Z(n52348) );
  NANDN U23980 ( .A(y[1057]), .B(x[1057]), .Z(n32013) );
  ANDN U23981 ( .B(x[1056]), .A(y[1056]), .Z(n32007) );
  ANDN U23982 ( .B(n32013), .A(n32007), .Z(n53075) );
  NANDN U23983 ( .A(x[1055]), .B(y[1055]), .Z(n32003) );
  NANDN U23984 ( .A(x[1056]), .B(y[1056]), .Z(n28097) );
  NAND U23985 ( .A(n32003), .B(n28097), .Z(n52349) );
  ANDN U23986 ( .B(x[1054]), .A(y[1054]), .Z(n31998) );
  ANDN U23987 ( .B(x[1055]), .A(y[1055]), .Z(n32008) );
  NOR U23988 ( .A(n31998), .B(n32008), .Z(n53074) );
  NANDN U23989 ( .A(y[1052]), .B(x[1052]), .Z(n31991) );
  ANDN U23990 ( .B(x[1053]), .A(y[1053]), .Z(n32001) );
  ANDN U23991 ( .B(n31991), .A(n32001), .Z(n53071) );
  ANDN U23992 ( .B(y[1051]), .A(x[1051]), .Z(n31987) );
  NANDN U23993 ( .A(x[1052]), .B(y[1052]), .Z(n31996) );
  NANDN U23994 ( .A(n31987), .B(n31996), .Z(n52350) );
  XNOR U23995 ( .A(x[1050]), .B(y[1050]), .Z(n10242) );
  ANDN U23996 ( .B(y[1049]), .A(x[1049]), .Z(n31978) );
  ANDN U23997 ( .B(n10242), .A(n31978), .Z(n53068) );
  NANDN U23998 ( .A(y[1048]), .B(x[1048]), .Z(n31976) );
  NANDN U23999 ( .A(y[1049]), .B(x[1049]), .Z(n31982) );
  NAND U24000 ( .A(n31976), .B(n31982), .Z(n53067) );
  NANDN U24001 ( .A(x[1047]), .B(y[1047]), .Z(n31971) );
  XNOR U24002 ( .A(x[1048]), .B(y[1048]), .Z(n10243) );
  NAND U24003 ( .A(n31971), .B(n10243), .Z(n53066) );
  NANDN U24004 ( .A(y[1046]), .B(x[1046]), .Z(n10244) );
  NANDN U24005 ( .A(y[1047]), .B(x[1047]), .Z(n31975) );
  AND U24006 ( .A(n10244), .B(n31975), .Z(n52351) );
  NANDN U24007 ( .A(x[1045]), .B(y[1045]), .Z(n31964) );
  XOR U24008 ( .A(y[1046]), .B(x[1046]), .Z(n31968) );
  ANDN U24009 ( .B(n31964), .A(n31968), .Z(n53065) );
  NANDN U24010 ( .A(y[1044]), .B(x[1044]), .Z(n31960) );
  NANDN U24011 ( .A(y[1045]), .B(x[1045]), .Z(n53064) );
  NAND U24012 ( .A(n31960), .B(n53064), .Z(n12114) );
  NANDN U24013 ( .A(x[1044]), .B(y[1044]), .Z(n53063) );
  ANDN U24014 ( .B(x[1042]), .A(y[1042]), .Z(n31954) );
  ANDN U24015 ( .B(x[1043]), .A(y[1043]), .Z(n31963) );
  OR U24016 ( .A(n31954), .B(n31963), .Z(n53060) );
  NANDN U24017 ( .A(x[1041]), .B(y[1041]), .Z(n31950) );
  NANDN U24018 ( .A(x[1042]), .B(y[1042]), .Z(n31958) );
  AND U24019 ( .A(n31950), .B(n31958), .Z(n53059) );
  ANDN U24020 ( .B(x[1040]), .A(y[1040]), .Z(n28100) );
  ANDN U24021 ( .B(x[1041]), .A(y[1041]), .Z(n31956) );
  OR U24022 ( .A(n28100), .B(n31956), .Z(n53058) );
  NANDN U24023 ( .A(x[1040]), .B(y[1040]), .Z(n31949) );
  ANDN U24024 ( .B(y[1039]), .A(x[1039]), .Z(n31944) );
  ANDN U24025 ( .B(n31949), .A(n31944), .Z(n53057) );
  ANDN U24026 ( .B(x[1039]), .A(y[1039]), .Z(n28099) );
  NANDN U24027 ( .A(y[1038]), .B(x[1038]), .Z(n31940) );
  NANDN U24028 ( .A(n28099), .B(n31940), .Z(n53056) );
  ANDN U24029 ( .B(y[1037]), .A(x[1037]), .Z(n31938) );
  ANDN U24030 ( .B(y[1038]), .A(x[1038]), .Z(n31945) );
  NOR U24031 ( .A(n31938), .B(n31945), .Z(n53055) );
  NANDN U24032 ( .A(y[1036]), .B(x[1036]), .Z(n10245) );
  NANDN U24033 ( .A(y[1037]), .B(x[1037]), .Z(n31939) );
  NAND U24034 ( .A(n10245), .B(n31939), .Z(n53053) );
  NANDN U24035 ( .A(x[1035]), .B(y[1035]), .Z(n31930) );
  XNOR U24036 ( .A(y[1036]), .B(x[1036]), .Z(n53052) );
  NANDN U24037 ( .A(y[1034]), .B(x[1034]), .Z(n53049) );
  NANDN U24038 ( .A(y[1035]), .B(x[1035]), .Z(n53051) );
  NAND U24039 ( .A(n53049), .B(n53051), .Z(n12101) );
  ANDN U24040 ( .B(y[1033]), .A(x[1033]), .Z(n53048) );
  NANDN U24041 ( .A(y[1032]), .B(x[1032]), .Z(n28102) );
  NANDN U24042 ( .A(y[1033]), .B(x[1033]), .Z(n28101) );
  NAND U24043 ( .A(n28102), .B(n28101), .Z(n53047) );
  NANDN U24044 ( .A(x[1031]), .B(y[1031]), .Z(n31920) );
  XNOR U24045 ( .A(y[1032]), .B(x[1032]), .Z(n10246) );
  AND U24046 ( .A(n31920), .B(n10246), .Z(n53046) );
  ANDN U24047 ( .B(x[1030]), .A(y[1030]), .Z(n31918) );
  NANDN U24048 ( .A(y[1031]), .B(x[1031]), .Z(n28103) );
  NANDN U24049 ( .A(n31918), .B(n28103), .Z(n53045) );
  NANDN U24050 ( .A(x[1029]), .B(y[1029]), .Z(n28104) );
  ANDN U24051 ( .B(y[1030]), .A(x[1030]), .Z(n31922) );
  ANDN U24052 ( .B(n28104), .A(n31922), .Z(n53044) );
  ANDN U24053 ( .B(x[1029]), .A(y[1029]), .Z(n31915) );
  NANDN U24054 ( .A(y[1028]), .B(x[1028]), .Z(n31910) );
  NANDN U24055 ( .A(n31915), .B(n31910), .Z(n53043) );
  NANDN U24056 ( .A(x[1028]), .B(y[1028]), .Z(n28105) );
  ANDN U24057 ( .B(y[1027]), .A(x[1027]), .Z(n31908) );
  ANDN U24058 ( .B(n28105), .A(n31908), .Z(n53042) );
  ANDN U24059 ( .B(x[1027]), .A(y[1027]), .Z(n31912) );
  NANDN U24060 ( .A(y[1026]), .B(x[1026]), .Z(n31903) );
  NANDN U24061 ( .A(n31912), .B(n31903), .Z(n53041) );
  ANDN U24062 ( .B(y[1026]), .A(x[1026]), .Z(n53040) );
  NANDN U24063 ( .A(y[1024]), .B(x[1024]), .Z(n53037) );
  NANDN U24064 ( .A(y[1022]), .B(x[1022]), .Z(n31894) );
  NANDN U24065 ( .A(y[1023]), .B(x[1023]), .Z(n28108) );
  NAND U24066 ( .A(n31894), .B(n28108), .Z(n53035) );
  ANDN U24067 ( .B(y[1021]), .A(x[1021]), .Z(n28110) );
  ANDN U24068 ( .B(y[1022]), .A(x[1022]), .Z(n31898) );
  NOR U24069 ( .A(n28110), .B(n31898), .Z(n53033) );
  ANDN U24070 ( .B(x[1020]), .A(y[1020]), .Z(n31888) );
  NANDN U24071 ( .A(y[1021]), .B(x[1021]), .Z(n31893) );
  NANDN U24072 ( .A(n31888), .B(n31893), .Z(n53032) );
  NANDN U24073 ( .A(x[1019]), .B(y[1019]), .Z(n31884) );
  ANDN U24074 ( .B(y[1020]), .A(x[1020]), .Z(n28109) );
  ANDN U24075 ( .B(n31884), .A(n28109), .Z(n53031) );
  ANDN U24076 ( .B(x[1018]), .A(y[1018]), .Z(n31879) );
  ANDN U24077 ( .B(x[1019]), .A(y[1019]), .Z(n31889) );
  NOR U24078 ( .A(n31879), .B(n31889), .Z(n53030) );
  NANDN U24079 ( .A(x[1017]), .B(y[1017]), .Z(n31877) );
  NANDN U24080 ( .A(x[1018]), .B(y[1018]), .Z(n31883) );
  NAND U24081 ( .A(n31877), .B(n31883), .Z(n52352) );
  ANDN U24082 ( .B(x[1016]), .A(y[1016]), .Z(n31875) );
  ANDN U24083 ( .B(x[1017]), .A(y[1017]), .Z(n31882) );
  NOR U24084 ( .A(n31875), .B(n31882), .Z(n53029) );
  ANDN U24085 ( .B(y[1016]), .A(x[1016]), .Z(n28111) );
  NANDN U24086 ( .A(y[1014]), .B(x[1014]), .Z(n31870) );
  NANDN U24087 ( .A(x[1014]), .B(y[1014]), .Z(n28114) );
  ANDN U24088 ( .B(y[1013]), .A(x[1013]), .Z(n28115) );
  ANDN U24089 ( .B(n28114), .A(n28115), .Z(n12073) );
  NANDN U24090 ( .A(x[1012]), .B(y[1012]), .Z(n10248) );
  NANDN U24091 ( .A(x[1011]), .B(y[1011]), .Z(n10247) );
  AND U24092 ( .A(n10248), .B(n10247), .Z(n53022) );
  NANDN U24093 ( .A(x[1010]), .B(y[1010]), .Z(n10250) );
  NANDN U24094 ( .A(x[1009]), .B(y[1009]), .Z(n10249) );
  AND U24095 ( .A(n10250), .B(n10249), .Z(n53020) );
  NANDN U24096 ( .A(y[1008]), .B(x[1008]), .Z(n10252) );
  NANDN U24097 ( .A(y[1009]), .B(x[1009]), .Z(n10251) );
  NAND U24098 ( .A(n10252), .B(n10251), .Z(n53019) );
  NANDN U24099 ( .A(x[1008]), .B(y[1008]), .Z(n31860) );
  NANDN U24100 ( .A(x[1007]), .B(y[1007]), .Z(n10253) );
  AND U24101 ( .A(n31860), .B(n10253), .Z(n53018) );
  ANDN U24102 ( .B(x[1006]), .A(y[1006]), .Z(n31850) );
  NANDN U24103 ( .A(y[1007]), .B(x[1007]), .Z(n31858) );
  NANDN U24104 ( .A(n31850), .B(n31858), .Z(n53017) );
  NANDN U24105 ( .A(x[1005]), .B(y[1005]), .Z(n31846) );
  NANDN U24106 ( .A(x[1006]), .B(y[1006]), .Z(n31854) );
  AND U24107 ( .A(n31846), .B(n31854), .Z(n53016) );
  ANDN U24108 ( .B(x[1005]), .A(y[1005]), .Z(n31852) );
  NANDN U24109 ( .A(y[1004]), .B(x[1004]), .Z(n28116) );
  NANDN U24110 ( .A(n31852), .B(n28116), .Z(n53014) );
  NANDN U24111 ( .A(x[1003]), .B(y[1003]), .Z(n28118) );
  NANDN U24112 ( .A(x[1004]), .B(y[1004]), .Z(n31845) );
  AND U24113 ( .A(n28118), .B(n31845), .Z(n53013) );
  ANDN U24114 ( .B(x[1002]), .A(y[1002]), .Z(n31838) );
  NANDN U24115 ( .A(y[1003]), .B(x[1003]), .Z(n28117) );
  NANDN U24116 ( .A(n31838), .B(n28117), .Z(n53012) );
  NANDN U24117 ( .A(x[1001]), .B(y[1001]), .Z(n31834) );
  NANDN U24118 ( .A(x[1002]), .B(y[1002]), .Z(n28119) );
  AND U24119 ( .A(n31834), .B(n28119), .Z(n53011) );
  ANDN U24120 ( .B(x[1000]), .A(y[1000]), .Z(n28121) );
  ANDN U24121 ( .B(x[1001]), .A(y[1001]), .Z(n31839) );
  OR U24122 ( .A(n28121), .B(n31839), .Z(n53010) );
  NANDN U24123 ( .A(x[1000]), .B(y[1000]), .Z(n31833) );
  ANDN U24124 ( .B(y[999]), .A(x[999]), .Z(n31828) );
  ANDN U24125 ( .B(n31833), .A(n31828), .Z(n53009) );
  ANDN U24126 ( .B(x[999]), .A(y[999]), .Z(n28120) );
  NANDN U24127 ( .A(y[998]), .B(x[998]), .Z(n31824) );
  NANDN U24128 ( .A(n28120), .B(n31824), .Z(n53008) );
  ANDN U24129 ( .B(y[997]), .A(x[997]), .Z(n31822) );
  ANDN U24130 ( .B(y[998]), .A(x[998]), .Z(n31829) );
  NOR U24131 ( .A(n31822), .B(n31829), .Z(n53007) );
  NANDN U24132 ( .A(y[996]), .B(x[996]), .Z(n10254) );
  NANDN U24133 ( .A(y[997]), .B(x[997]), .Z(n31823) );
  NAND U24134 ( .A(n10254), .B(n31823), .Z(n53006) );
  XNOR U24135 ( .A(y[996]), .B(x[996]), .Z(n53005) );
  NANDN U24136 ( .A(y[994]), .B(x[994]), .Z(n53004) );
  NANDN U24137 ( .A(y[995]), .B(x[995]), .Z(n52353) );
  NAND U24138 ( .A(n53004), .B(n52353), .Z(n12050) );
  NANDN U24139 ( .A(y[992]), .B(x[992]), .Z(n31806) );
  NANDN U24140 ( .A(y[993]), .B(x[993]), .Z(n28122) );
  NAND U24141 ( .A(n31806), .B(n28122), .Z(n53002) );
  ANDN U24142 ( .B(y[991]), .A(x[991]), .Z(n31801) );
  ANDN U24143 ( .B(y[992]), .A(x[992]), .Z(n31810) );
  NOR U24144 ( .A(n31801), .B(n31810), .Z(n53001) );
  NANDN U24145 ( .A(y[990]), .B(x[990]), .Z(n31798) );
  NANDN U24146 ( .A(y[991]), .B(x[991]), .Z(n31805) );
  NAND U24147 ( .A(n31798), .B(n31805), .Z(n53000) );
  NANDN U24148 ( .A(x[989]), .B(y[989]), .Z(n31794) );
  ANDN U24149 ( .B(y[990]), .A(x[990]), .Z(n31804) );
  ANDN U24150 ( .B(n31794), .A(n31804), .Z(n52998) );
  ANDN U24151 ( .B(x[988]), .A(y[988]), .Z(n31790) );
  NANDN U24152 ( .A(y[989]), .B(x[989]), .Z(n31799) );
  NANDN U24153 ( .A(n31790), .B(n31799), .Z(n52997) );
  NANDN U24154 ( .A(x[987]), .B(y[987]), .Z(n31786) );
  ANDN U24155 ( .B(y[988]), .A(x[988]), .Z(n31796) );
  ANDN U24156 ( .B(n31786), .A(n31796), .Z(n52996) );
  ANDN U24157 ( .B(x[986]), .A(y[986]), .Z(n31782) );
  ANDN U24158 ( .B(x[987]), .A(y[987]), .Z(n31792) );
  OR U24159 ( .A(n31782), .B(n31792), .Z(n52995) );
  NANDN U24160 ( .A(x[985]), .B(y[985]), .Z(n31780) );
  NANDN U24161 ( .A(x[986]), .B(y[986]), .Z(n31785) );
  AND U24162 ( .A(n31780), .B(n31785), .Z(n52994) );
  NANDN U24163 ( .A(y[984]), .B(x[984]), .Z(n52991) );
  NANDN U24164 ( .A(y[985]), .B(x[985]), .Z(n52993) );
  NAND U24165 ( .A(n52991), .B(n52993), .Z(n12038) );
  NANDN U24166 ( .A(x[984]), .B(y[984]), .Z(n52992) );
  ANDN U24167 ( .B(x[983]), .A(y[983]), .Z(n31778) );
  NANDN U24168 ( .A(y[982]), .B(x[982]), .Z(n10255) );
  NANDN U24169 ( .A(n31778), .B(n10255), .Z(n52989) );
  XNOR U24170 ( .A(y[982]), .B(x[982]), .Z(n31770) );
  ANDN U24171 ( .B(y[981]), .A(x[981]), .Z(n28124) );
  ANDN U24172 ( .B(n31770), .A(n28124), .Z(n52988) );
  ANDN U24173 ( .B(x[980]), .A(y[980]), .Z(n31764) );
  NANDN U24174 ( .A(y[981]), .B(x[981]), .Z(n31769) );
  NANDN U24175 ( .A(n31764), .B(n31769), .Z(n52987) );
  NANDN U24176 ( .A(x[979]), .B(y[979]), .Z(n31760) );
  ANDN U24177 ( .B(y[980]), .A(x[980]), .Z(n28123) );
  ANDN U24178 ( .B(n31760), .A(n28123), .Z(n52986) );
  NANDN U24179 ( .A(x[977]), .B(y[977]), .Z(n31753) );
  NANDN U24180 ( .A(x[978]), .B(y[978]), .Z(n31759) );
  AND U24181 ( .A(n31753), .B(n31759), .Z(n52984) );
  ANDN U24182 ( .B(x[976]), .A(y[976]), .Z(n31751) );
  ANDN U24183 ( .B(x[977]), .A(y[977]), .Z(n31758) );
  OR U24184 ( .A(n31751), .B(n31758), .Z(n52983) );
  NANDN U24185 ( .A(x[976]), .B(y[976]), .Z(n52982) );
  NANDN U24186 ( .A(y[974]), .B(x[974]), .Z(n52978) );
  NANDN U24187 ( .A(y[975]), .B(x[975]), .Z(n52981) );
  NAND U24188 ( .A(n52978), .B(n52981), .Z(n12025) );
  NANDN U24189 ( .A(x[973]), .B(y[973]), .Z(n52977) );
  ANDN U24190 ( .B(x[972]), .A(y[972]), .Z(n31742) );
  NANDN U24191 ( .A(y[973]), .B(x[973]), .Z(n28127) );
  NANDN U24192 ( .A(n31742), .B(n28127), .Z(n52976) );
  NANDN U24193 ( .A(x[971]), .B(y[971]), .Z(n28129) );
  XNOR U24194 ( .A(x[972]), .B(y[972]), .Z(n10256) );
  AND U24195 ( .A(n28129), .B(n10256), .Z(n52975) );
  ANDN U24196 ( .B(x[970]), .A(y[970]), .Z(n31734) );
  ANDN U24197 ( .B(x[971]), .A(y[971]), .Z(n31739) );
  OR U24198 ( .A(n31734), .B(n31739), .Z(n52974) );
  NANDN U24199 ( .A(x[969]), .B(y[969]), .Z(n31730) );
  XNOR U24200 ( .A(x[970]), .B(y[970]), .Z(n10257) );
  AND U24201 ( .A(n31730), .B(n10257), .Z(n52973) );
  ANDN U24202 ( .B(x[968]), .A(y[968]), .Z(n31725) );
  ANDN U24203 ( .B(x[969]), .A(y[969]), .Z(n31735) );
  OR U24204 ( .A(n31725), .B(n31735), .Z(n52972) );
  NANDN U24205 ( .A(x[967]), .B(y[967]), .Z(n31722) );
  NANDN U24206 ( .A(x[968]), .B(y[968]), .Z(n31729) );
  AND U24207 ( .A(n31722), .B(n31729), .Z(n52971) );
  ANDN U24208 ( .B(x[967]), .A(y[967]), .Z(n31728) );
  NANDN U24209 ( .A(y[966]), .B(x[966]), .Z(n10258) );
  NANDN U24210 ( .A(n31728), .B(n10258), .Z(n52970) );
  XNOR U24211 ( .A(y[966]), .B(x[966]), .Z(n52969) );
  ANDN U24212 ( .B(x[964]), .A(y[964]), .Z(n52967) );
  NANDN U24213 ( .A(y[965]), .B(x[965]), .Z(n52968) );
  NANDN U24214 ( .A(n52967), .B(n52968), .Z(n12012) );
  NANDN U24215 ( .A(x[963]), .B(y[963]), .Z(n52966) );
  ANDN U24216 ( .B(x[963]), .A(y[963]), .Z(n31715) );
  NANDN U24217 ( .A(y[962]), .B(x[962]), .Z(n28130) );
  NANDN U24218 ( .A(n31715), .B(n28130), .Z(n52965) );
  NANDN U24219 ( .A(x[961]), .B(y[961]), .Z(n28132) );
  NANDN U24220 ( .A(x[962]), .B(y[962]), .Z(n31710) );
  AND U24221 ( .A(n28132), .B(n31710), .Z(n52964) );
  ANDN U24222 ( .B(x[960]), .A(y[960]), .Z(n31703) );
  NANDN U24223 ( .A(y[961]), .B(x[961]), .Z(n28131) );
  NANDN U24224 ( .A(n31703), .B(n28131), .Z(n52963) );
  NANDN U24225 ( .A(x[959]), .B(y[959]), .Z(n31699) );
  NANDN U24226 ( .A(x[960]), .B(y[960]), .Z(n28133) );
  AND U24227 ( .A(n31699), .B(n28133), .Z(n52962) );
  ANDN U24228 ( .B(x[959]), .A(y[959]), .Z(n31704) );
  NANDN U24229 ( .A(y[958]), .B(x[958]), .Z(n28134) );
  NANDN U24230 ( .A(n31704), .B(n28134), .Z(n52960) );
  NANDN U24231 ( .A(x[957]), .B(y[957]), .Z(n28136) );
  NANDN U24232 ( .A(x[958]), .B(y[958]), .Z(n31698) );
  AND U24233 ( .A(n28136), .B(n31698), .Z(n52959) );
  ANDN U24234 ( .B(x[956]), .A(y[956]), .Z(n31691) );
  NANDN U24235 ( .A(y[957]), .B(x[957]), .Z(n28135) );
  NANDN U24236 ( .A(n31691), .B(n28135), .Z(n52958) );
  NANDN U24237 ( .A(x[955]), .B(y[955]), .Z(n31687) );
  NANDN U24238 ( .A(x[956]), .B(y[956]), .Z(n28137) );
  AND U24239 ( .A(n31687), .B(n28137), .Z(n52957) );
  ANDN U24240 ( .B(x[955]), .A(y[955]), .Z(n31692) );
  NANDN U24241 ( .A(y[954]), .B(x[954]), .Z(n28138) );
  NANDN U24242 ( .A(n31692), .B(n28138), .Z(n52956) );
  NANDN U24243 ( .A(x[953]), .B(y[953]), .Z(n28140) );
  NANDN U24244 ( .A(x[954]), .B(y[954]), .Z(n31686) );
  AND U24245 ( .A(n28140), .B(n31686), .Z(n52955) );
  ANDN U24246 ( .B(x[952]), .A(y[952]), .Z(n31679) );
  NANDN U24247 ( .A(y[953]), .B(x[953]), .Z(n28139) );
  NANDN U24248 ( .A(n31679), .B(n28139), .Z(n52954) );
  NANDN U24249 ( .A(x[951]), .B(y[951]), .Z(n31675) );
  NANDN U24250 ( .A(x[952]), .B(y[952]), .Z(n28141) );
  AND U24251 ( .A(n31675), .B(n28141), .Z(n52953) );
  ANDN U24252 ( .B(x[950]), .A(y[950]), .Z(n28143) );
  ANDN U24253 ( .B(x[951]), .A(y[951]), .Z(n31680) );
  OR U24254 ( .A(n28143), .B(n31680), .Z(n52952) );
  NANDN U24255 ( .A(x[950]), .B(y[950]), .Z(n31674) );
  ANDN U24256 ( .B(y[949]), .A(x[949]), .Z(n31669) );
  ANDN U24257 ( .B(n31674), .A(n31669), .Z(n52951) );
  ANDN U24258 ( .B(x[949]), .A(y[949]), .Z(n28142) );
  NANDN U24259 ( .A(y[948]), .B(x[948]), .Z(n31665) );
  NANDN U24260 ( .A(n28142), .B(n31665), .Z(n52950) );
  ANDN U24261 ( .B(y[947]), .A(x[947]), .Z(n31661) );
  ANDN U24262 ( .B(y[948]), .A(x[948]), .Z(n31670) );
  NOR U24263 ( .A(n31661), .B(n31670), .Z(n52949) );
  NANDN U24264 ( .A(y[946]), .B(x[946]), .Z(n31659) );
  NANDN U24265 ( .A(y[947]), .B(x[947]), .Z(n31664) );
  NAND U24266 ( .A(n31659), .B(n31664), .Z(n52948) );
  NANDN U24267 ( .A(x[945]), .B(y[945]), .Z(n31655) );
  ANDN U24268 ( .B(y[946]), .A(x[946]), .Z(n52947) );
  ANDN U24269 ( .B(n31655), .A(n52947), .Z(n11991) );
  NANDN U24270 ( .A(y[944]), .B(x[944]), .Z(n52945) );
  NANDN U24271 ( .A(y[945]), .B(x[945]), .Z(n52356) );
  NAND U24272 ( .A(n52945), .B(n52356), .Z(n11989) );
  NANDN U24273 ( .A(x[944]), .B(y[944]), .Z(n31656) );
  ANDN U24274 ( .B(y[943]), .A(x[943]), .Z(n52943) );
  ANDN U24275 ( .B(n31656), .A(n52943), .Z(n11987) );
  NANDN U24276 ( .A(y[942]), .B(x[942]), .Z(n31647) );
  NANDN U24277 ( .A(y[943]), .B(x[943]), .Z(n28144) );
  NAND U24278 ( .A(n31647), .B(n28144), .Z(n52942) );
  ANDN U24279 ( .B(y[941]), .A(x[941]), .Z(n31642) );
  ANDN U24280 ( .B(y[942]), .A(x[942]), .Z(n31651) );
  NOR U24281 ( .A(n31642), .B(n31651), .Z(n52941) );
  NANDN U24282 ( .A(y[940]), .B(x[940]), .Z(n31639) );
  NANDN U24283 ( .A(y[941]), .B(x[941]), .Z(n31646) );
  NAND U24284 ( .A(n31639), .B(n31646), .Z(n52940) );
  NANDN U24285 ( .A(x[939]), .B(y[939]), .Z(n31634) );
  ANDN U24286 ( .B(y[940]), .A(x[940]), .Z(n31645) );
  ANDN U24287 ( .B(n31634), .A(n31645), .Z(n52939) );
  NANDN U24288 ( .A(y[938]), .B(x[938]), .Z(n28146) );
  NANDN U24289 ( .A(y[939]), .B(x[939]), .Z(n31640) );
  NAND U24290 ( .A(n28146), .B(n31640), .Z(n52938) );
  NANDN U24291 ( .A(x[938]), .B(y[938]), .Z(n31635) );
  ANDN U24292 ( .B(y[937]), .A(x[937]), .Z(n31630) );
  ANDN U24293 ( .B(n31635), .A(n31630), .Z(n52937) );
  NANDN U24294 ( .A(y[936]), .B(x[936]), .Z(n31626) );
  NANDN U24295 ( .A(y[937]), .B(x[937]), .Z(n28145) );
  NAND U24296 ( .A(n31626), .B(n28145), .Z(n52936) );
  NANDN U24297 ( .A(x[935]), .B(y[935]), .Z(n28148) );
  ANDN U24298 ( .B(y[936]), .A(x[936]), .Z(n52358) );
  ANDN U24299 ( .B(n28148), .A(n52358), .Z(n11978) );
  NANDN U24300 ( .A(y[934]), .B(x[934]), .Z(n52934) );
  NANDN U24301 ( .A(y[932]), .B(x[932]), .Z(n10259) );
  ANDN U24302 ( .B(x[933]), .A(y[933]), .Z(n31620) );
  ANDN U24303 ( .B(n10259), .A(n31620), .Z(n52932) );
  ANDN U24304 ( .B(y[931]), .A(x[931]), .Z(n31616) );
  NANDN U24305 ( .A(x[932]), .B(y[932]), .Z(n31618) );
  NANDN U24306 ( .A(n31616), .B(n31618), .Z(n52360) );
  NANDN U24307 ( .A(y[931]), .B(x[931]), .Z(n10261) );
  NANDN U24308 ( .A(y[930]), .B(x[930]), .Z(n10260) );
  AND U24309 ( .A(n10261), .B(n10260), .Z(n28149) );
  NANDN U24310 ( .A(x[929]), .B(y[929]), .Z(n10263) );
  NANDN U24311 ( .A(x[930]), .B(y[930]), .Z(n10262) );
  NAND U24312 ( .A(n10263), .B(n10262), .Z(n28150) );
  NANDN U24313 ( .A(y[929]), .B(x[929]), .Z(n10265) );
  NANDN U24314 ( .A(y[928]), .B(x[928]), .Z(n10264) );
  AND U24315 ( .A(n10265), .B(n10264), .Z(n31611) );
  ANDN U24316 ( .B(x[927]), .A(y[927]), .Z(n31608) );
  ANDN U24317 ( .B(x[926]), .A(y[926]), .Z(n31605) );
  NOR U24318 ( .A(n31608), .B(n31605), .Z(n52926) );
  NANDN U24319 ( .A(y[924]), .B(x[924]), .Z(n52922) );
  NANDN U24320 ( .A(y[925]), .B(x[925]), .Z(n28151) );
  AND U24321 ( .A(n52922), .B(n28151), .Z(n11961) );
  NANDN U24322 ( .A(y[922]), .B(x[922]), .Z(n31593) );
  ANDN U24323 ( .B(x[923]), .A(y[923]), .Z(n31601) );
  ANDN U24324 ( .B(n31593), .A(n31601), .Z(n52920) );
  ANDN U24325 ( .B(y[921]), .A(x[921]), .Z(n28155) );
  ANDN U24326 ( .B(y[922]), .A(x[922]), .Z(n31597) );
  OR U24327 ( .A(n28155), .B(n31597), .Z(n52361) );
  NANDN U24328 ( .A(y[921]), .B(x[921]), .Z(n31592) );
  ANDN U24329 ( .B(x[920]), .A(y[920]), .Z(n31587) );
  ANDN U24330 ( .B(n31592), .A(n31587), .Z(n52919) );
  ANDN U24331 ( .B(y[920]), .A(x[920]), .Z(n28154) );
  NANDN U24332 ( .A(x[919]), .B(y[919]), .Z(n31583) );
  NANDN U24333 ( .A(n28154), .B(n31583), .Z(n52362) );
  ANDN U24334 ( .B(x[918]), .A(y[918]), .Z(n31578) );
  ANDN U24335 ( .B(x[919]), .A(y[919]), .Z(n31588) );
  NOR U24336 ( .A(n31578), .B(n31588), .Z(n52918) );
  ANDN U24337 ( .B(x[916]), .A(y[916]), .Z(n31572) );
  ANDN U24338 ( .B(x[917]), .A(y[917]), .Z(n31581) );
  NOR U24339 ( .A(n31572), .B(n31581), .Z(n52916) );
  NANDN U24340 ( .A(y[914]), .B(x[914]), .Z(n52911) );
  NANDN U24341 ( .A(y[915]), .B(x[915]), .Z(n31571) );
  AND U24342 ( .A(n52911), .B(n31571), .Z(n11948) );
  NANDN U24343 ( .A(y[913]), .B(x[913]), .Z(n31566) );
  ANDN U24344 ( .B(x[912]), .A(y[912]), .Z(n31561) );
  ANDN U24345 ( .B(n31566), .A(n31561), .Z(n52909) );
  NANDN U24346 ( .A(x[911]), .B(y[911]), .Z(n28160) );
  XNOR U24347 ( .A(y[912]), .B(x[912]), .Z(n10266) );
  NAND U24348 ( .A(n28160), .B(n10266), .Z(n52363) );
  NANDN U24349 ( .A(y[910]), .B(x[910]), .Z(n31555) );
  ANDN U24350 ( .B(x[911]), .A(y[911]), .Z(n31562) );
  ANDN U24351 ( .B(n31555), .A(n31562), .Z(n52908) );
  ANDN U24352 ( .B(y[909]), .A(x[909]), .Z(n31553) );
  NANDN U24353 ( .A(x[910]), .B(y[910]), .Z(n28161) );
  NANDN U24354 ( .A(n31553), .B(n28161), .Z(n52907) );
  NANDN U24355 ( .A(y[908]), .B(x[908]), .Z(n28162) );
  ANDN U24356 ( .B(x[909]), .A(y[909]), .Z(n31557) );
  ANDN U24357 ( .B(n28162), .A(n31557), .Z(n52906) );
  NANDN U24358 ( .A(y[907]), .B(x[907]), .Z(n28163) );
  ANDN U24359 ( .B(x[906]), .A(y[906]), .Z(n31541) );
  ANDN U24360 ( .B(n28163), .A(n31541), .Z(n52905) );
  ANDN U24361 ( .B(y[906]), .A(x[906]), .Z(n31547) );
  NANDN U24362 ( .A(x[905]), .B(y[905]), .Z(n31537) );
  NANDN U24363 ( .A(n31547), .B(n31537), .Z(n52365) );
  NANDN U24364 ( .A(y[904]), .B(x[904]), .Z(n28164) );
  ANDN U24365 ( .B(x[905]), .A(y[905]), .Z(n31543) );
  ANDN U24366 ( .B(n28164), .A(n31543), .Z(n52904) );
  NANDN U24367 ( .A(x[903]), .B(y[903]), .Z(n28166) );
  NANDN U24368 ( .A(x[904]), .B(y[904]), .Z(n31536) );
  NAND U24369 ( .A(n28166), .B(n31536), .Z(n52901) );
  NANDN U24370 ( .A(y[902]), .B(x[902]), .Z(n31529) );
  NANDN U24371 ( .A(y[903]), .B(x[903]), .Z(n28165) );
  AND U24372 ( .A(n31529), .B(n28165), .Z(n52366) );
  NANDN U24373 ( .A(y[900]), .B(x[900]), .Z(n28168) );
  ANDN U24374 ( .B(x[901]), .A(y[901]), .Z(n31531) );
  ANDN U24375 ( .B(n28168), .A(n31531), .Z(n52900) );
  ANDN U24376 ( .B(y[900]), .A(x[900]), .Z(n31524) );
  NANDN U24377 ( .A(x[899]), .B(y[899]), .Z(n31519) );
  NANDN U24378 ( .A(n31524), .B(n31519), .Z(n52368) );
  NANDN U24379 ( .A(y[899]), .B(x[899]), .Z(n28169) );
  ANDN U24380 ( .B(x[898]), .A(y[898]), .Z(n31515) );
  ANDN U24381 ( .B(n28169), .A(n31515), .Z(n52899) );
  ANDN U24382 ( .B(y[898]), .A(x[898]), .Z(n31521) );
  NANDN U24383 ( .A(x[897]), .B(y[897]), .Z(n31511) );
  NANDN U24384 ( .A(n31521), .B(n31511), .Z(n52898) );
  NANDN U24385 ( .A(y[896]), .B(x[896]), .Z(n10267) );
  ANDN U24386 ( .B(x[897]), .A(y[897]), .Z(n31517) );
  ANDN U24387 ( .B(n10267), .A(n31517), .Z(n52897) );
  NANDN U24388 ( .A(y[895]), .B(x[895]), .Z(n28170) );
  ANDN U24389 ( .B(x[894]), .A(y[894]), .Z(n31503) );
  ANDN U24390 ( .B(n28170), .A(n31503), .Z(n52896) );
  NANDN U24391 ( .A(x[893]), .B(y[893]), .Z(n31499) );
  NANDN U24392 ( .A(x[894]), .B(y[894]), .Z(n28173) );
  NAND U24393 ( .A(n31499), .B(n28173), .Z(n52370) );
  NANDN U24394 ( .A(y[892]), .B(x[892]), .Z(n31497) );
  ANDN U24395 ( .B(x[893]), .A(y[893]), .Z(n31504) );
  ANDN U24396 ( .B(n31497), .A(n31504), .Z(n52895) );
  ANDN U24397 ( .B(y[891]), .A(x[891]), .Z(n31495) );
  XNOR U24398 ( .A(x[892]), .B(y[892]), .Z(n10268) );
  NANDN U24399 ( .A(n31495), .B(n10268), .Z(n52894) );
  NANDN U24400 ( .A(y[891]), .B(x[891]), .Z(n10270) );
  NANDN U24401 ( .A(y[890]), .B(x[890]), .Z(n10269) );
  AND U24402 ( .A(n10270), .B(n10269), .Z(n52371) );
  NANDN U24403 ( .A(x[887]), .B(y[887]), .Z(n10271) );
  ANDN U24404 ( .B(y[888]), .A(x[888]), .Z(n31487) );
  ANDN U24405 ( .B(n10271), .A(n31487), .Z(n11916) );
  NANDN U24406 ( .A(x[886]), .B(y[886]), .Z(n10272) );
  AND U24407 ( .A(n11916), .B(n10272), .Z(n52891) );
  ANDN U24408 ( .B(y[885]), .A(x[885]), .Z(n31479) );
  NANDN U24409 ( .A(y[885]), .B(x[885]), .Z(n52890) );
  NANDN U24410 ( .A(y[884]), .B(x[884]), .Z(n52374) );
  AND U24411 ( .A(n52890), .B(n52374), .Z(n11910) );
  ANDN U24412 ( .B(y[883]), .A(x[883]), .Z(n52375) );
  NANDN U24413 ( .A(y[882]), .B(x[882]), .Z(n10273) );
  ANDN U24414 ( .B(x[883]), .A(y[883]), .Z(n28175) );
  ANDN U24415 ( .B(n10273), .A(n28175), .Z(n52888) );
  ANDN U24416 ( .B(y[879]), .A(x[879]), .Z(n31464) );
  NANDN U24417 ( .A(x[880]), .B(y[880]), .Z(n31470) );
  NANDN U24418 ( .A(n31464), .B(n31470), .Z(n52886) );
  NANDN U24419 ( .A(y[878]), .B(x[878]), .Z(n31460) );
  NANDN U24420 ( .A(y[879]), .B(x[879]), .Z(n28177) );
  AND U24421 ( .A(n31460), .B(n28177), .Z(n52377) );
  ANDN U24422 ( .B(y[877]), .A(x[877]), .Z(n31456) );
  ANDN U24423 ( .B(y[878]), .A(x[878]), .Z(n31465) );
  OR U24424 ( .A(n31456), .B(n31465), .Z(n52378) );
  NANDN U24425 ( .A(y[876]), .B(x[876]), .Z(n31454) );
  NANDN U24426 ( .A(y[877]), .B(x[877]), .Z(n31459) );
  AND U24427 ( .A(n31454), .B(n31459), .Z(n52379) );
  ANDN U24428 ( .B(y[875]), .A(x[875]), .Z(n28179) );
  ANDN U24429 ( .B(y[873]), .A(x[873]), .Z(n31445) );
  ANDN U24430 ( .B(x[872]), .A(y[872]), .Z(n31441) );
  ANDN U24431 ( .B(x[873]), .A(y[873]), .Z(n31450) );
  NOR U24432 ( .A(n31441), .B(n31450), .Z(n52879) );
  NANDN U24433 ( .A(x[871]), .B(y[871]), .Z(n31438) );
  NANDN U24434 ( .A(x[872]), .B(y[872]), .Z(n31446) );
  NAND U24435 ( .A(n31438), .B(n31446), .Z(n52380) );
  NANDN U24436 ( .A(y[870]), .B(x[870]), .Z(n31434) );
  ANDN U24437 ( .B(x[871]), .A(y[871]), .Z(n31444) );
  ANDN U24438 ( .B(n31434), .A(n31444), .Z(n52878) );
  NANDN U24439 ( .A(y[868]), .B(x[868]), .Z(n31426) );
  ANDN U24440 ( .B(x[869]), .A(y[869]), .Z(n31436) );
  ANDN U24441 ( .B(n31426), .A(n31436), .Z(n52876) );
  ANDN U24442 ( .B(y[867]), .A(x[867]), .Z(n31422) );
  ANDN U24443 ( .B(y[868]), .A(x[868]), .Z(n31432) );
  OR U24444 ( .A(n31422), .B(n31432), .Z(n52381) );
  NANDN U24445 ( .A(y[866]), .B(x[866]), .Z(n31420) );
  NANDN U24446 ( .A(y[867]), .B(x[867]), .Z(n31425) );
  AND U24447 ( .A(n31420), .B(n31425), .Z(n52382) );
  ANDN U24448 ( .B(y[866]), .A(x[866]), .Z(n52383) );
  NANDN U24449 ( .A(y[864]), .B(x[864]), .Z(n52384) );
  ANDN U24450 ( .B(y[861]), .A(x[861]), .Z(n31404) );
  ANDN U24451 ( .B(y[862]), .A(x[862]), .Z(n31413) );
  OR U24452 ( .A(n31404), .B(n31413), .Z(n52387) );
  NANDN U24453 ( .A(y[860]), .B(x[860]), .Z(n31401) );
  NANDN U24454 ( .A(y[861]), .B(x[861]), .Z(n31408) );
  AND U24455 ( .A(n31401), .B(n31408), .Z(n52871) );
  ANDN U24456 ( .B(y[860]), .A(x[860]), .Z(n31407) );
  NANDN U24457 ( .A(x[859]), .B(y[859]), .Z(n31396) );
  NANDN U24458 ( .A(n31407), .B(n31396), .Z(n52870) );
  NANDN U24459 ( .A(y[858]), .B(x[858]), .Z(n28184) );
  NANDN U24460 ( .A(y[859]), .B(x[859]), .Z(n31402) );
  AND U24461 ( .A(n28184), .B(n31402), .Z(n52388) );
  ANDN U24462 ( .B(y[855]), .A(x[855]), .Z(n31382) );
  ANDN U24463 ( .B(y[856]), .A(x[856]), .Z(n31392) );
  OR U24464 ( .A(n31382), .B(n31392), .Z(n52391) );
  NANDN U24465 ( .A(y[854]), .B(x[854]), .Z(n31379) );
  NANDN U24466 ( .A(y[855]), .B(x[855]), .Z(n31386) );
  AND U24467 ( .A(n31379), .B(n31386), .Z(n52867) );
  ANDN U24468 ( .B(y[853]), .A(x[853]), .Z(n31375) );
  ANDN U24469 ( .B(y[854]), .A(x[854]), .Z(n31385) );
  OR U24470 ( .A(n31375), .B(n31385), .Z(n52866) );
  NANDN U24471 ( .A(y[852]), .B(x[852]), .Z(n31371) );
  NANDN U24472 ( .A(y[853]), .B(x[853]), .Z(n31380) );
  AND U24473 ( .A(n31371), .B(n31380), .Z(n52392) );
  NANDN U24474 ( .A(x[849]), .B(y[849]), .Z(n31363) );
  NANDN U24475 ( .A(x[850]), .B(y[850]), .Z(n28186) );
  NAND U24476 ( .A(n31363), .B(n28186), .Z(n52395) );
  NANDN U24477 ( .A(y[849]), .B(x[849]), .Z(n28188) );
  ANDN U24478 ( .B(x[848]), .A(y[848]), .Z(n31361) );
  ANDN U24479 ( .B(n28188), .A(n31361), .Z(n52865) );
  ANDN U24480 ( .B(y[848]), .A(x[848]), .Z(n31365) );
  NANDN U24481 ( .A(x[847]), .B(y[847]), .Z(n28189) );
  NANDN U24482 ( .A(n31365), .B(n28189), .Z(n52864) );
  NANDN U24483 ( .A(y[846]), .B(x[846]), .Z(n31354) );
  ANDN U24484 ( .B(x[847]), .A(y[847]), .Z(n31358) );
  ANDN U24485 ( .B(n31354), .A(n31358), .Z(n52863) );
  NANDN U24486 ( .A(y[844]), .B(x[844]), .Z(n52859) );
  NANDN U24487 ( .A(y[845]), .B(x[845]), .Z(n28191) );
  AND U24488 ( .A(n52859), .B(n28191), .Z(n11861) );
  NANDN U24489 ( .A(y[842]), .B(x[842]), .Z(n31342) );
  NANDN U24490 ( .A(y[843]), .B(x[843]), .Z(n28192) );
  NAND U24491 ( .A(n31342), .B(n28192), .Z(n52857) );
  NANDN U24492 ( .A(x[841]), .B(y[841]), .Z(n28193) );
  XNOR U24493 ( .A(y[842]), .B(x[842]), .Z(n10274) );
  AND U24494 ( .A(n28193), .B(n10274), .Z(n52856) );
  NANDN U24495 ( .A(y[840]), .B(x[840]), .Z(n28195) );
  NANDN U24496 ( .A(y[841]), .B(x[841]), .Z(n31341) );
  NAND U24497 ( .A(n28195), .B(n31341), .Z(n52855) );
  NANDN U24498 ( .A(x[840]), .B(y[840]), .Z(n28194) );
  ANDN U24499 ( .B(y[839]), .A(x[839]), .Z(n31336) );
  ANDN U24500 ( .B(n28194), .A(n31336), .Z(n52854) );
  NANDN U24501 ( .A(y[838]), .B(x[838]), .Z(n31334) );
  NANDN U24502 ( .A(y[839]), .B(x[839]), .Z(n28196) );
  NAND U24503 ( .A(n31334), .B(n28196), .Z(n52853) );
  NANDN U24504 ( .A(x[838]), .B(y[838]), .Z(n10276) );
  NANDN U24505 ( .A(x[837]), .B(y[837]), .Z(n10275) );
  NAND U24506 ( .A(n10276), .B(n10275), .Z(n52852) );
  NANDN U24507 ( .A(y[837]), .B(x[837]), .Z(n31330) );
  NANDN U24508 ( .A(y[836]), .B(x[836]), .Z(n31326) );
  NAND U24509 ( .A(n31330), .B(n31326), .Z(n52851) );
  NANDN U24510 ( .A(x[835]), .B(y[835]), .Z(n28198) );
  NANDN U24511 ( .A(y[834]), .B(x[834]), .Z(n52848) );
  NANDN U24512 ( .A(y[832]), .B(x[832]), .Z(n31316) );
  NANDN U24513 ( .A(y[833]), .B(x[833]), .Z(n31322) );
  NAND U24514 ( .A(n31316), .B(n31322), .Z(n52845) );
  XNOR U24515 ( .A(y[832]), .B(x[832]), .Z(n10277) );
  ANDN U24516 ( .B(y[831]), .A(x[831]), .Z(n31312) );
  ANDN U24517 ( .B(n10277), .A(n31312), .Z(n52843) );
  NANDN U24518 ( .A(y[830]), .B(x[830]), .Z(n31308) );
  NANDN U24519 ( .A(y[831]), .B(x[831]), .Z(n31317) );
  NAND U24520 ( .A(n31308), .B(n31317), .Z(n52841) );
  NANDN U24521 ( .A(x[829]), .B(y[829]), .Z(n28200) );
  ANDN U24522 ( .B(y[830]), .A(x[830]), .Z(n31314) );
  ANDN U24523 ( .B(n28200), .A(n31314), .Z(n52839) );
  ANDN U24524 ( .B(x[828]), .A(y[828]), .Z(n31302) );
  NANDN U24525 ( .A(y[829]), .B(x[829]), .Z(n31307) );
  NANDN U24526 ( .A(n31302), .B(n31307), .Z(n52837) );
  NANDN U24527 ( .A(x[827]), .B(y[827]), .Z(n31300) );
  XNOR U24528 ( .A(x[828]), .B(y[828]), .Z(n10278) );
  AND U24529 ( .A(n31300), .B(n10278), .Z(n52835) );
  ANDN U24530 ( .B(x[826]), .A(y[826]), .Z(n31298) );
  ANDN U24531 ( .B(x[827]), .A(y[827]), .Z(n31303) );
  OR U24532 ( .A(n31298), .B(n31303), .Z(n52833) );
  NANDN U24533 ( .A(x[825]), .B(y[825]), .Z(n31290) );
  XNOR U24534 ( .A(x[826]), .B(y[826]), .Z(n10279) );
  AND U24535 ( .A(n31290), .B(n10279), .Z(n52831) );
  ANDN U24536 ( .B(x[825]), .A(y[825]), .Z(n31294) );
  ANDN U24537 ( .B(x[824]), .A(y[824]), .Z(n31286) );
  OR U24538 ( .A(n31294), .B(n31286), .Z(n52829) );
  NANDN U24539 ( .A(x[823]), .B(y[823]), .Z(n31282) );
  NANDN U24540 ( .A(x[824]), .B(y[824]), .Z(n31291) );
  AND U24541 ( .A(n31282), .B(n31291), .Z(n52827) );
  ANDN U24542 ( .B(x[823]), .A(y[823]), .Z(n31288) );
  NANDN U24543 ( .A(y[822]), .B(x[822]), .Z(n28201) );
  NANDN U24544 ( .A(n31288), .B(n28201), .Z(n52825) );
  NANDN U24545 ( .A(x[821]), .B(y[821]), .Z(n28203) );
  NANDN U24546 ( .A(x[822]), .B(y[822]), .Z(n31281) );
  AND U24547 ( .A(n28203), .B(n31281), .Z(n52823) );
  ANDN U24548 ( .B(x[820]), .A(y[820]), .Z(n31274) );
  NANDN U24549 ( .A(y[821]), .B(x[821]), .Z(n28202) );
  NANDN U24550 ( .A(n31274), .B(n28202), .Z(n52821) );
  NANDN U24551 ( .A(x[819]), .B(y[819]), .Z(n31270) );
  NANDN U24552 ( .A(x[820]), .B(y[820]), .Z(n28204) );
  AND U24553 ( .A(n31270), .B(n28204), .Z(n52819) );
  ANDN U24554 ( .B(x[819]), .A(y[819]), .Z(n31275) );
  NANDN U24555 ( .A(y[818]), .B(x[818]), .Z(n28206) );
  NANDN U24556 ( .A(n31275), .B(n28206), .Z(n52817) );
  NANDN U24557 ( .A(x[818]), .B(y[818]), .Z(n31269) );
  ANDN U24558 ( .B(y[817]), .A(x[817]), .Z(n31264) );
  ANDN U24559 ( .B(n31269), .A(n31264), .Z(n52815) );
  NANDN U24560 ( .A(y[816]), .B(x[816]), .Z(n10280) );
  NANDN U24561 ( .A(y[817]), .B(x[817]), .Z(n28205) );
  NAND U24562 ( .A(n10280), .B(n28205), .Z(n52813) );
  NANDN U24563 ( .A(x[815]), .B(y[815]), .Z(n28207) );
  XNOR U24564 ( .A(y[816]), .B(x[816]), .Z(n52811) );
  AND U24565 ( .A(n28207), .B(n52811), .Z(n11827) );
  NANDN U24566 ( .A(y[815]), .B(x[815]), .Z(n52808) );
  NANDN U24567 ( .A(x[814]), .B(y[814]), .Z(n28208) );
  NANDN U24568 ( .A(y[812]), .B(x[812]), .Z(n31252) );
  NANDN U24569 ( .A(y[813]), .B(x[813]), .Z(n28209) );
  NAND U24570 ( .A(n31252), .B(n28209), .Z(n52800) );
  NANDN U24571 ( .A(x[811]), .B(y[811]), .Z(n28210) );
  ANDN U24572 ( .B(y[812]), .A(x[812]), .Z(n31256) );
  ANDN U24573 ( .B(n28210), .A(n31256), .Z(n52798) );
  NANDN U24574 ( .A(y[810]), .B(x[810]), .Z(n28212) );
  NANDN U24575 ( .A(y[811]), .B(x[811]), .Z(n31251) );
  NAND U24576 ( .A(n28212), .B(n31251), .Z(n52796) );
  NANDN U24577 ( .A(x[810]), .B(y[810]), .Z(n28211) );
  ANDN U24578 ( .B(y[809]), .A(x[809]), .Z(n31244) );
  ANDN U24579 ( .B(n28211), .A(n31244), .Z(n52794) );
  NANDN U24580 ( .A(y[808]), .B(x[808]), .Z(n31240) );
  NANDN U24581 ( .A(y[809]), .B(x[809]), .Z(n28213) );
  NAND U24582 ( .A(n31240), .B(n28213), .Z(n52792) );
  ANDN U24583 ( .B(y[807]), .A(x[807]), .Z(n28214) );
  ANDN U24584 ( .B(y[808]), .A(x[808]), .Z(n31245) );
  NOR U24585 ( .A(n28214), .B(n31245), .Z(n52790) );
  NANDN U24586 ( .A(y[806]), .B(x[806]), .Z(n10281) );
  NANDN U24587 ( .A(y[807]), .B(x[807]), .Z(n31239) );
  NAND U24588 ( .A(n10281), .B(n31239), .Z(n52788) );
  XNOR U24589 ( .A(y[806]), .B(x[806]), .Z(n31234) );
  NANDN U24590 ( .A(x[805]), .B(y[805]), .Z(n31230) );
  AND U24591 ( .A(n31234), .B(n31230), .Z(n52786) );
  ANDN U24592 ( .B(x[804]), .A(y[804]), .Z(n31228) );
  NANDN U24593 ( .A(y[805]), .B(x[805]), .Z(n31233) );
  NANDN U24594 ( .A(n31228), .B(n31233), .Z(n52784) );
  NANDN U24595 ( .A(x[803]), .B(y[803]), .Z(n28216) );
  NANDN U24596 ( .A(x[804]), .B(y[804]), .Z(n31231) );
  AND U24597 ( .A(n28216), .B(n31231), .Z(n52782) );
  ANDN U24598 ( .B(x[803]), .A(y[803]), .Z(n31225) );
  NANDN U24599 ( .A(y[802]), .B(x[802]), .Z(n31220) );
  NANDN U24600 ( .A(n31225), .B(n31220), .Z(n52780) );
  NANDN U24601 ( .A(x[802]), .B(y[802]), .Z(n28217) );
  ANDN U24602 ( .B(y[801]), .A(x[801]), .Z(n31216) );
  ANDN U24603 ( .B(n28217), .A(n31216), .Z(n52778) );
  ANDN U24604 ( .B(x[801]), .A(y[801]), .Z(n31222) );
  NANDN U24605 ( .A(y[800]), .B(x[800]), .Z(n31212) );
  NANDN U24606 ( .A(n31222), .B(n31212), .Z(n52776) );
  NANDN U24607 ( .A(x[799]), .B(y[799]), .Z(n28218) );
  ANDN U24608 ( .B(y[800]), .A(x[800]), .Z(n31218) );
  ANDN U24609 ( .B(n28218), .A(n31218), .Z(n52774) );
  NANDN U24610 ( .A(y[798]), .B(x[798]), .Z(n31206) );
  NANDN U24611 ( .A(y[799]), .B(x[799]), .Z(n31214) );
  NAND U24612 ( .A(n31206), .B(n31214), .Z(n52772) );
  NANDN U24613 ( .A(x[798]), .B(y[798]), .Z(n28219) );
  ANDN U24614 ( .B(y[797]), .A(x[797]), .Z(n31204) );
  ANDN U24615 ( .B(n28219), .A(n31204), .Z(n52770) );
  ANDN U24616 ( .B(x[797]), .A(y[797]), .Z(n31208) );
  NANDN U24617 ( .A(y[796]), .B(x[796]), .Z(n31199) );
  NANDN U24618 ( .A(n31208), .B(n31199), .Z(n52768) );
  NANDN U24619 ( .A(y[794]), .B(x[794]), .Z(n52764) );
  NANDN U24620 ( .A(y[795]), .B(x[795]), .Z(n52398) );
  NAND U24621 ( .A(n52764), .B(n52398), .Z(n11802) );
  NANDN U24622 ( .A(y[792]), .B(x[792]), .Z(n31190) );
  NANDN U24623 ( .A(y[793]), .B(x[793]), .Z(n28222) );
  NAND U24624 ( .A(n31190), .B(n28222), .Z(n52762) );
  ANDN U24625 ( .B(y[791]), .A(x[791]), .Z(n28224) );
  ANDN U24626 ( .B(y[792]), .A(x[792]), .Z(n31194) );
  NOR U24627 ( .A(n28224), .B(n31194), .Z(n52761) );
  ANDN U24628 ( .B(x[790]), .A(y[790]), .Z(n31184) );
  NANDN U24629 ( .A(y[791]), .B(x[791]), .Z(n31189) );
  NANDN U24630 ( .A(n31184), .B(n31189), .Z(n52760) );
  NANDN U24631 ( .A(x[789]), .B(y[789]), .Z(n31180) );
  ANDN U24632 ( .B(y[790]), .A(x[790]), .Z(n28223) );
  ANDN U24633 ( .B(n31180), .A(n28223), .Z(n52759) );
  ANDN U24634 ( .B(x[788]), .A(y[788]), .Z(n31175) );
  ANDN U24635 ( .B(x[789]), .A(y[789]), .Z(n31185) );
  OR U24636 ( .A(n31175), .B(n31185), .Z(n52758) );
  NANDN U24637 ( .A(x[787]), .B(y[787]), .Z(n31172) );
  NANDN U24638 ( .A(x[788]), .B(y[788]), .Z(n31179) );
  AND U24639 ( .A(n31172), .B(n31179), .Z(n52757) );
  ANDN U24640 ( .B(x[787]), .A(y[787]), .Z(n31178) );
  NANDN U24641 ( .A(y[786]), .B(x[786]), .Z(n10282) );
  NANDN U24642 ( .A(n31178), .B(n10282), .Z(n52756) );
  XNOR U24643 ( .A(y[786]), .B(x[786]), .Z(n52755) );
  NANDN U24644 ( .A(y[784]), .B(x[784]), .Z(n31166) );
  NANDN U24645 ( .A(y[785]), .B(x[785]), .Z(n52400) );
  NAND U24646 ( .A(n31166), .B(n52400), .Z(n11789) );
  NANDN U24647 ( .A(x[783]), .B(y[783]), .Z(n52752) );
  NANDN U24648 ( .A(y[783]), .B(x[783]), .Z(n10284) );
  NANDN U24649 ( .A(y[782]), .B(x[782]), .Z(n10283) );
  NAND U24650 ( .A(n10284), .B(n10283), .Z(n52750) );
  NANDN U24651 ( .A(x[782]), .B(y[782]), .Z(n10286) );
  NANDN U24652 ( .A(x[781]), .B(y[781]), .Z(n10285) );
  AND U24653 ( .A(n10286), .B(n10285), .Z(n52749) );
  NANDN U24654 ( .A(y[780]), .B(x[780]), .Z(n10287) );
  ANDN U24655 ( .B(x[781]), .A(y[781]), .Z(n31157) );
  ANDN U24656 ( .B(n10287), .A(n31157), .Z(n52748) );
  NANDN U24657 ( .A(x[779]), .B(y[779]), .Z(n28227) );
  NANDN U24658 ( .A(x[780]), .B(y[780]), .Z(n10288) );
  AND U24659 ( .A(n28227), .B(n10288), .Z(n52401) );
  ANDN U24660 ( .B(x[777]), .A(y[777]), .Z(n31151) );
  NANDN U24661 ( .A(y[776]), .B(x[776]), .Z(n31143) );
  NANDN U24662 ( .A(n31151), .B(n31143), .Z(n52404) );
  NANDN U24663 ( .A(x[775]), .B(y[775]), .Z(n31141) );
  XNOR U24664 ( .A(y[776]), .B(x[776]), .Z(n10289) );
  AND U24665 ( .A(n31141), .B(n10289), .Z(n52747) );
  NANDN U24666 ( .A(y[775]), .B(x[775]), .Z(n52746) );
  ANDN U24667 ( .B(x[774]), .A(y[774]), .Z(n52745) );
  ANDN U24668 ( .B(n52746), .A(n52745), .Z(n11777) );
  NANDN U24669 ( .A(x[774]), .B(y[774]), .Z(n52405) );
  ANDN U24670 ( .B(x[772]), .A(y[772]), .Z(n28230) );
  ANDN U24671 ( .B(x[773]), .A(y[773]), .Z(n31138) );
  OR U24672 ( .A(n28230), .B(n31138), .Z(n52407) );
  NANDN U24673 ( .A(x[772]), .B(y[772]), .Z(n31133) );
  ANDN U24674 ( .B(y[771]), .A(x[771]), .Z(n31128) );
  ANDN U24675 ( .B(n31133), .A(n31128), .Z(n52742) );
  ANDN U24676 ( .B(y[769]), .A(x[769]), .Z(n31119) );
  ANDN U24677 ( .B(y[770]), .A(x[770]), .Z(n31129) );
  NOR U24678 ( .A(n31119), .B(n31129), .Z(n52740) );
  NANDN U24679 ( .A(y[768]), .B(x[768]), .Z(n31116) );
  NANDN U24680 ( .A(y[769]), .B(x[769]), .Z(n31123) );
  NAND U24681 ( .A(n31116), .B(n31123), .Z(n52408) );
  ANDN U24682 ( .B(y[767]), .A(x[767]), .Z(n31112) );
  ANDN U24683 ( .B(y[768]), .A(x[768]), .Z(n31122) );
  NOR U24684 ( .A(n31112), .B(n31122), .Z(n52739) );
  NANDN U24685 ( .A(y[766]), .B(x[766]), .Z(n31108) );
  NANDN U24686 ( .A(y[767]), .B(x[767]), .Z(n31117) );
  NAND U24687 ( .A(n31108), .B(n31117), .Z(n52409) );
  NANDN U24688 ( .A(x[766]), .B(y[766]), .Z(n31113) );
  NANDN U24689 ( .A(y[764]), .B(x[764]), .Z(n52735) );
  NANDN U24690 ( .A(y[765]), .B(x[765]), .Z(n52737) );
  NAND U24691 ( .A(n52735), .B(n52737), .Z(n11764) );
  ANDN U24692 ( .B(y[763]), .A(x[763]), .Z(n52734) );
  NANDN U24693 ( .A(y[762]), .B(x[762]), .Z(n31099) );
  NANDN U24694 ( .A(y[763]), .B(x[763]), .Z(n28233) );
  NAND U24695 ( .A(n31099), .B(n28233), .Z(n52733) );
  NANDN U24696 ( .A(x[761]), .B(y[761]), .Z(n28234) );
  ANDN U24697 ( .B(y[762]), .A(x[762]), .Z(n31103) );
  ANDN U24698 ( .B(n28234), .A(n31103), .Z(n52732) );
  NANDN U24699 ( .A(y[760]), .B(x[760]), .Z(n28236) );
  NANDN U24700 ( .A(y[761]), .B(x[761]), .Z(n31098) );
  NAND U24701 ( .A(n28236), .B(n31098), .Z(n52731) );
  NANDN U24702 ( .A(x[760]), .B(y[760]), .Z(n28235) );
  ANDN U24703 ( .B(y[759]), .A(x[759]), .Z(n31091) );
  ANDN U24704 ( .B(n28235), .A(n31091), .Z(n52730) );
  NANDN U24705 ( .A(y[758]), .B(x[758]), .Z(n31087) );
  NANDN U24706 ( .A(y[759]), .B(x[759]), .Z(n28237) );
  NAND U24707 ( .A(n31087), .B(n28237), .Z(n52729) );
  NANDN U24708 ( .A(x[757]), .B(y[757]), .Z(n28238) );
  ANDN U24709 ( .B(y[758]), .A(x[758]), .Z(n31092) );
  ANDN U24710 ( .B(n28238), .A(n31092), .Z(n52728) );
  NANDN U24711 ( .A(y[756]), .B(x[756]), .Z(n28240) );
  NANDN U24712 ( .A(y[757]), .B(x[757]), .Z(n31086) );
  NAND U24713 ( .A(n28240), .B(n31086), .Z(n52726) );
  NANDN U24714 ( .A(x[756]), .B(y[756]), .Z(n28239) );
  ANDN U24715 ( .B(y[755]), .A(x[755]), .Z(n31079) );
  ANDN U24716 ( .B(n28239), .A(n31079), .Z(n52724) );
  NANDN U24717 ( .A(y[754]), .B(x[754]), .Z(n31075) );
  NANDN U24718 ( .A(y[755]), .B(x[755]), .Z(n28241) );
  NAND U24719 ( .A(n31075), .B(n28241), .Z(n52722) );
  NANDN U24720 ( .A(x[753]), .B(y[753]), .Z(n28242) );
  ANDN U24721 ( .B(y[754]), .A(x[754]), .Z(n31080) );
  ANDN U24722 ( .B(n28242), .A(n31080), .Z(n52720) );
  NANDN U24723 ( .A(y[752]), .B(x[752]), .Z(n28244) );
  NANDN U24724 ( .A(y[753]), .B(x[753]), .Z(n31074) );
  NAND U24725 ( .A(n28244), .B(n31074), .Z(n52718) );
  NANDN U24726 ( .A(x[752]), .B(y[752]), .Z(n28243) );
  ANDN U24727 ( .B(y[751]), .A(x[751]), .Z(n31067) );
  ANDN U24728 ( .B(n28243), .A(n31067), .Z(n52716) );
  NANDN U24729 ( .A(y[750]), .B(x[750]), .Z(n31063) );
  NANDN U24730 ( .A(y[751]), .B(x[751]), .Z(n28245) );
  NAND U24731 ( .A(n31063), .B(n28245), .Z(n52714) );
  ANDN U24732 ( .B(y[749]), .A(x[749]), .Z(n28247) );
  ANDN U24733 ( .B(y[750]), .A(x[750]), .Z(n31068) );
  NOR U24734 ( .A(n28247), .B(n31068), .Z(n52712) );
  ANDN U24735 ( .B(x[748]), .A(y[748]), .Z(n31057) );
  NANDN U24736 ( .A(y[749]), .B(x[749]), .Z(n31062) );
  NANDN U24737 ( .A(n31057), .B(n31062), .Z(n52710) );
  NANDN U24738 ( .A(x[747]), .B(y[747]), .Z(n31053) );
  ANDN U24739 ( .B(y[748]), .A(x[748]), .Z(n28246) );
  ANDN U24740 ( .B(n31053), .A(n28246), .Z(n52708) );
  ANDN U24741 ( .B(x[746]), .A(y[746]), .Z(n31049) );
  ANDN U24742 ( .B(x[747]), .A(y[747]), .Z(n31058) );
  OR U24743 ( .A(n31049), .B(n31058), .Z(n52706) );
  NANDN U24744 ( .A(x[745]), .B(y[745]), .Z(n31047) );
  NANDN U24745 ( .A(x[746]), .B(y[746]), .Z(n31052) );
  AND U24746 ( .A(n31047), .B(n31052), .Z(n52704) );
  NANDN U24747 ( .A(y[744]), .B(x[744]), .Z(n52697) );
  NANDN U24748 ( .A(y[745]), .B(x[745]), .Z(n28248) );
  AND U24749 ( .A(n52697), .B(n28248), .Z(n11742) );
  NANDN U24750 ( .A(x[744]), .B(y[744]), .Z(n52700) );
  ANDN U24751 ( .B(x[742]), .A(y[742]), .Z(n28250) );
  ANDN U24752 ( .B(x[743]), .A(y[743]), .Z(n31045) );
  OR U24753 ( .A(n28250), .B(n31045), .Z(n52694) );
  NANDN U24754 ( .A(x[742]), .B(y[742]), .Z(n31040) );
  ANDN U24755 ( .B(y[741]), .A(x[741]), .Z(n31035) );
  ANDN U24756 ( .B(n31040), .A(n31035), .Z(n52692) );
  ANDN U24757 ( .B(x[741]), .A(y[741]), .Z(n28249) );
  NANDN U24758 ( .A(y[740]), .B(x[740]), .Z(n31031) );
  NANDN U24759 ( .A(n28249), .B(n31031), .Z(n52690) );
  ANDN U24760 ( .B(y[739]), .A(x[739]), .Z(n31026) );
  ANDN U24761 ( .B(y[740]), .A(x[740]), .Z(n31036) );
  NOR U24762 ( .A(n31026), .B(n31036), .Z(n52688) );
  NANDN U24763 ( .A(y[738]), .B(x[738]), .Z(n31023) );
  NANDN U24764 ( .A(y[739]), .B(x[739]), .Z(n31030) );
  NAND U24765 ( .A(n31023), .B(n31030), .Z(n52686) );
  NANDN U24766 ( .A(x[737]), .B(y[737]), .Z(n31019) );
  ANDN U24767 ( .B(y[738]), .A(x[738]), .Z(n31029) );
  ANDN U24768 ( .B(n31019), .A(n31029), .Z(n52685) );
  ANDN U24769 ( .B(x[736]), .A(y[736]), .Z(n31016) );
  NANDN U24770 ( .A(y[737]), .B(x[737]), .Z(n31024) );
  NANDN U24771 ( .A(n31016), .B(n31024), .Z(n52684) );
  NANDN U24772 ( .A(x[735]), .B(y[735]), .Z(n31012) );
  ANDN U24773 ( .B(y[736]), .A(x[736]), .Z(n31021) );
  ANDN U24774 ( .B(n31012), .A(n31021), .Z(n52683) );
  NANDN U24775 ( .A(y[734]), .B(x[734]), .Z(n31008) );
  NANDN U24776 ( .A(y[735]), .B(x[735]), .Z(n52682) );
  NAND U24777 ( .A(n31008), .B(n52682), .Z(n11730) );
  NANDN U24778 ( .A(x[733]), .B(y[733]), .Z(n52679) );
  NANDN U24779 ( .A(x[734]), .B(y[734]), .Z(n52681) );
  AND U24780 ( .A(n52679), .B(n52681), .Z(n11728) );
  ANDN U24781 ( .B(x[732]), .A(y[732]), .Z(n31002) );
  ANDN U24782 ( .B(x[733]), .A(y[733]), .Z(n31011) );
  OR U24783 ( .A(n31002), .B(n31011), .Z(n52678) );
  NANDN U24784 ( .A(x[731]), .B(y[731]), .Z(n30998) );
  NANDN U24785 ( .A(x[732]), .B(y[732]), .Z(n31006) );
  AND U24786 ( .A(n30998), .B(n31006), .Z(n52677) );
  ANDN U24787 ( .B(x[730]), .A(y[730]), .Z(n28252) );
  ANDN U24788 ( .B(x[731]), .A(y[731]), .Z(n31004) );
  OR U24789 ( .A(n28252), .B(n31004), .Z(n52676) );
  NANDN U24790 ( .A(x[730]), .B(y[730]), .Z(n30997) );
  ANDN U24791 ( .B(y[729]), .A(x[729]), .Z(n30992) );
  ANDN U24792 ( .B(n30997), .A(n30992), .Z(n52675) );
  ANDN U24793 ( .B(x[729]), .A(y[729]), .Z(n28251) );
  NANDN U24794 ( .A(y[728]), .B(x[728]), .Z(n28253) );
  NANDN U24795 ( .A(n28251), .B(n28253), .Z(n52674) );
  XNOR U24796 ( .A(y[728]), .B(x[728]), .Z(n10290) );
  ANDN U24797 ( .B(y[727]), .A(x[727]), .Z(n30986) );
  ANDN U24798 ( .B(n10290), .A(n30986), .Z(n52673) );
  NANDN U24799 ( .A(y[726]), .B(x[726]), .Z(n10291) );
  NANDN U24800 ( .A(y[727]), .B(x[727]), .Z(n28254) );
  NAND U24801 ( .A(n10291), .B(n28254), .Z(n52672) );
  NANDN U24802 ( .A(x[725]), .B(y[725]), .Z(n28255) );
  XNOR U24803 ( .A(y[726]), .B(x[726]), .Z(n52671) );
  AND U24804 ( .A(n28255), .B(n52671), .Z(n11719) );
  NANDN U24805 ( .A(y[724]), .B(x[724]), .Z(n52669) );
  NANDN U24806 ( .A(y[725]), .B(x[725]), .Z(n52410) );
  NAND U24807 ( .A(n52669), .B(n52410), .Z(n11717) );
  NANDN U24808 ( .A(x[724]), .B(y[724]), .Z(n28256) );
  ANDN U24809 ( .B(y[723]), .A(x[723]), .Z(n52668) );
  ANDN U24810 ( .B(n28256), .A(n52668), .Z(n11715) );
  NANDN U24811 ( .A(y[722]), .B(x[722]), .Z(n30974) );
  NANDN U24812 ( .A(y[723]), .B(x[723]), .Z(n28257) );
  NAND U24813 ( .A(n30974), .B(n28257), .Z(n52667) );
  ANDN U24814 ( .B(y[721]), .A(x[721]), .Z(n28259) );
  ANDN U24815 ( .B(y[722]), .A(x[722]), .Z(n30978) );
  NOR U24816 ( .A(n28259), .B(n30978), .Z(n52666) );
  ANDN U24817 ( .B(x[720]), .A(y[720]), .Z(n30968) );
  NANDN U24818 ( .A(y[721]), .B(x[721]), .Z(n30973) );
  NANDN U24819 ( .A(n30968), .B(n30973), .Z(n52665) );
  NANDN U24820 ( .A(x[719]), .B(y[719]), .Z(n30964) );
  ANDN U24821 ( .B(y[720]), .A(x[720]), .Z(n28258) );
  ANDN U24822 ( .B(n30964), .A(n28258), .Z(n52664) );
  ANDN U24823 ( .B(x[718]), .A(y[718]), .Z(n30959) );
  ANDN U24824 ( .B(x[719]), .A(y[719]), .Z(n30969) );
  OR U24825 ( .A(n30959), .B(n30969), .Z(n52663) );
  NANDN U24826 ( .A(x[717]), .B(y[717]), .Z(n30957) );
  NANDN U24827 ( .A(x[718]), .B(y[718]), .Z(n30963) );
  AND U24828 ( .A(n30957), .B(n30963), .Z(n52662) );
  ANDN U24829 ( .B(x[716]), .A(y[716]), .Z(n30954) );
  ANDN U24830 ( .B(x[717]), .A(y[717]), .Z(n30962) );
  OR U24831 ( .A(n30954), .B(n30962), .Z(n52661) );
  NANDN U24832 ( .A(x[715]), .B(y[715]), .Z(n28260) );
  NANDN U24833 ( .A(x[716]), .B(y[716]), .Z(n52660) );
  AND U24834 ( .A(n28260), .B(n52660), .Z(n11706) );
  NANDN U24835 ( .A(y[714]), .B(x[714]), .Z(n28262) );
  NANDN U24836 ( .A(y[715]), .B(x[715]), .Z(n52659) );
  NAND U24837 ( .A(n28262), .B(n52659), .Z(n11704) );
  NANDN U24838 ( .A(x[714]), .B(y[714]), .Z(n28261) );
  NANDN U24839 ( .A(x[713]), .B(y[713]), .Z(n52656) );
  AND U24840 ( .A(n28261), .B(n52656), .Z(n11702) );
  ANDN U24841 ( .B(x[712]), .A(y[712]), .Z(n30945) );
  ANDN U24842 ( .B(x[713]), .A(y[713]), .Z(n30950) );
  OR U24843 ( .A(n30945), .B(n30950), .Z(n52655) );
  NANDN U24844 ( .A(x[711]), .B(y[711]), .Z(n30943) );
  NANDN U24845 ( .A(x[712]), .B(y[712]), .Z(n30946) );
  AND U24846 ( .A(n30943), .B(n30946), .Z(n52654) );
  NANDN U24847 ( .A(y[710]), .B(x[710]), .Z(n10293) );
  NANDN U24848 ( .A(y[711]), .B(x[711]), .Z(n10292) );
  NAND U24849 ( .A(n10293), .B(n10292), .Z(n52653) );
  NANDN U24850 ( .A(x[710]), .B(y[710]), .Z(n10295) );
  NANDN U24851 ( .A(x[709]), .B(y[709]), .Z(n10294) );
  AND U24852 ( .A(n10295), .B(n10294), .Z(n52652) );
  NANDN U24853 ( .A(y[708]), .B(x[708]), .Z(n10297) );
  NANDN U24854 ( .A(y[709]), .B(x[709]), .Z(n10296) );
  NAND U24855 ( .A(n10297), .B(n10296), .Z(n52651) );
  NANDN U24856 ( .A(x[708]), .B(y[708]), .Z(n10299) );
  NANDN U24857 ( .A(x[707]), .B(y[707]), .Z(n10298) );
  AND U24858 ( .A(n10299), .B(n10298), .Z(n52649) );
  NANDN U24859 ( .A(y[706]), .B(x[706]), .Z(n10301) );
  NANDN U24860 ( .A(y[707]), .B(x[707]), .Z(n10300) );
  NAND U24861 ( .A(n10301), .B(n10300), .Z(n52647) );
  NANDN U24862 ( .A(x[706]), .B(y[706]), .Z(n30936) );
  NANDN U24863 ( .A(x[705]), .B(y[705]), .Z(n10302) );
  AND U24864 ( .A(n30936), .B(n10302), .Z(n52645) );
  ANDN U24865 ( .B(x[704]), .A(y[704]), .Z(n30926) );
  NANDN U24866 ( .A(y[705]), .B(x[705]), .Z(n30934) );
  NANDN U24867 ( .A(n30926), .B(n30934), .Z(n52643) );
  NANDN U24868 ( .A(x[703]), .B(y[703]), .Z(n30922) );
  NANDN U24869 ( .A(x[704]), .B(y[704]), .Z(n30930) );
  AND U24870 ( .A(n30922), .B(n30930), .Z(n52641) );
  ANDN U24871 ( .B(x[702]), .A(y[702]), .Z(n30917) );
  ANDN U24872 ( .B(x[703]), .A(y[703]), .Z(n30928) );
  OR U24873 ( .A(n30917), .B(n30928), .Z(n52639) );
  NANDN U24874 ( .A(x[701]), .B(y[701]), .Z(n30914) );
  NANDN U24875 ( .A(x[702]), .B(y[702]), .Z(n30921) );
  AND U24876 ( .A(n30914), .B(n30921), .Z(n52637) );
  ANDN U24877 ( .B(x[701]), .A(y[701]), .Z(n30920) );
  NANDN U24878 ( .A(y[700]), .B(x[700]), .Z(n30910) );
  NANDN U24879 ( .A(n30920), .B(n30910), .Z(n52635) );
  NANDN U24880 ( .A(x[700]), .B(y[700]), .Z(n30915) );
  ANDN U24881 ( .B(y[699]), .A(x[699]), .Z(n30906) );
  ANDN U24882 ( .B(n30915), .A(n30906), .Z(n52633) );
  ANDN U24883 ( .B(x[699]), .A(y[699]), .Z(n30912) );
  NANDN U24884 ( .A(y[698]), .B(x[698]), .Z(n30902) );
  NANDN U24885 ( .A(n30912), .B(n30902), .Z(n52631) );
  ANDN U24886 ( .B(y[697]), .A(x[697]), .Z(n28264) );
  ANDN U24887 ( .B(y[698]), .A(x[698]), .Z(n30908) );
  NOR U24888 ( .A(n28264), .B(n30908), .Z(n52629) );
  NANDN U24889 ( .A(y[696]), .B(x[696]), .Z(n10303) );
  NANDN U24890 ( .A(y[697]), .B(x[697]), .Z(n30901) );
  NAND U24891 ( .A(n10303), .B(n30901), .Z(n52627) );
  XNOR U24892 ( .A(y[696]), .B(x[696]), .Z(n30897) );
  NANDN U24893 ( .A(x[695]), .B(y[695]), .Z(n30892) );
  AND U24894 ( .A(n30897), .B(n30892), .Z(n52625) );
  ANDN U24895 ( .B(x[694]), .A(y[694]), .Z(n30887) );
  ANDN U24896 ( .B(x[695]), .A(y[695]), .Z(n30896) );
  OR U24897 ( .A(n30887), .B(n30896), .Z(n52623) );
  NANDN U24898 ( .A(x[693]), .B(y[693]), .Z(n30884) );
  NANDN U24899 ( .A(x[694]), .B(y[694]), .Z(n30891) );
  AND U24900 ( .A(n30884), .B(n30891), .Z(n52621) );
  ANDN U24901 ( .B(x[693]), .A(y[693]), .Z(n30890) );
  NANDN U24902 ( .A(y[692]), .B(x[692]), .Z(n30879) );
  NANDN U24903 ( .A(n30890), .B(n30879), .Z(n52619) );
  NANDN U24904 ( .A(x[691]), .B(y[691]), .Z(n28266) );
  NANDN U24905 ( .A(x[692]), .B(y[692]), .Z(n30885) );
  AND U24906 ( .A(n28266), .B(n30885), .Z(n52617) );
  ANDN U24907 ( .B(x[690]), .A(y[690]), .Z(n30874) );
  NANDN U24908 ( .A(y[691]), .B(x[691]), .Z(n30880) );
  NANDN U24909 ( .A(n30874), .B(n30880), .Z(n52615) );
  NANDN U24910 ( .A(x[689]), .B(y[689]), .Z(n30870) );
  NANDN U24911 ( .A(x[690]), .B(y[690]), .Z(n28265) );
  AND U24912 ( .A(n30870), .B(n28265), .Z(n52613) );
  ANDN U24913 ( .B(x[688]), .A(y[688]), .Z(n30865) );
  ANDN U24914 ( .B(x[689]), .A(y[689]), .Z(n30875) );
  OR U24915 ( .A(n30865), .B(n30875), .Z(n52611) );
  NANDN U24916 ( .A(x[687]), .B(y[687]), .Z(n30862) );
  NANDN U24917 ( .A(x[688]), .B(y[688]), .Z(n30869) );
  AND U24918 ( .A(n30862), .B(n30869), .Z(n52609) );
  ANDN U24919 ( .B(x[687]), .A(y[687]), .Z(n30868) );
  NANDN U24920 ( .A(y[686]), .B(x[686]), .Z(n10304) );
  NANDN U24921 ( .A(n30868), .B(n10304), .Z(n52608) );
  XNOR U24922 ( .A(y[686]), .B(x[686]), .Z(n52607) );
  ANDN U24923 ( .B(y[683]), .A(x[683]), .Z(n30851) );
  ANDN U24924 ( .B(x[682]), .A(y[682]), .Z(n28270) );
  ANDN U24925 ( .B(x[683]), .A(y[683]), .Z(n30856) );
  NOR U24926 ( .A(n28270), .B(n30856), .Z(n52602) );
  ANDN U24927 ( .B(y[681]), .A(x[681]), .Z(n30846) );
  NANDN U24928 ( .A(x[682]), .B(y[682]), .Z(n30852) );
  NANDN U24929 ( .A(n30846), .B(n30852), .Z(n52412) );
  NANDN U24930 ( .A(y[680]), .B(x[680]), .Z(n30842) );
  ANDN U24931 ( .B(x[681]), .A(y[681]), .Z(n28269) );
  ANDN U24932 ( .B(n30842), .A(n28269), .Z(n52601) );
  ANDN U24933 ( .B(y[677]), .A(x[677]), .Z(n30831) );
  ANDN U24934 ( .B(y[678]), .A(x[678]), .Z(n30840) );
  OR U24935 ( .A(n30831), .B(n30840), .Z(n52414) );
  NANDN U24936 ( .A(y[676]), .B(x[676]), .Z(n30827) );
  NANDN U24937 ( .A(y[677]), .B(x[677]), .Z(n30835) );
  AND U24938 ( .A(n30827), .B(n30835), .Z(n52415) );
  ANDN U24939 ( .B(y[676]), .A(x[676]), .Z(n52416) );
  NANDN U24940 ( .A(y[674]), .B(x[674]), .Z(n52417) );
  ANDN U24941 ( .B(y[671]), .A(x[671]), .Z(n30814) );
  ANDN U24942 ( .B(y[672]), .A(x[672]), .Z(n30819) );
  OR U24943 ( .A(n30814), .B(n30819), .Z(n52419) );
  NANDN U24944 ( .A(y[670]), .B(x[670]), .Z(n28274) );
  NANDN U24945 ( .A(y[671]), .B(x[671]), .Z(n30817) );
  AND U24946 ( .A(n28274), .B(n30817), .Z(n52595) );
  ANDN U24947 ( .B(y[669]), .A(x[669]), .Z(n30806) );
  ANDN U24948 ( .B(y[670]), .A(x[670]), .Z(n30811) );
  OR U24949 ( .A(n30806), .B(n30811), .Z(n52594) );
  NANDN U24950 ( .A(y[668]), .B(x[668]), .Z(n30802) );
  NANDN U24951 ( .A(y[669]), .B(x[669]), .Z(n28273) );
  AND U24952 ( .A(n30802), .B(n28273), .Z(n52420) );
  NANDN U24953 ( .A(y[665]), .B(x[665]), .Z(n52592) );
  NANDN U24954 ( .A(y[664]), .B(x[664]), .Z(n52424) );
  AND U24955 ( .A(n52592), .B(n52424), .Z(n11645) );
  ANDN U24956 ( .B(y[663]), .A(x[663]), .Z(n52425) );
  NANDN U24957 ( .A(y[662]), .B(x[662]), .Z(n10306) );
  NANDN U24958 ( .A(y[663]), .B(x[663]), .Z(n10305) );
  AND U24959 ( .A(n10306), .B(n10305), .Z(n52426) );
  NANDN U24960 ( .A(x[662]), .B(y[662]), .Z(n10308) );
  NANDN U24961 ( .A(x[661]), .B(y[661]), .Z(n10307) );
  NAND U24962 ( .A(n10308), .B(n10307), .Z(n52590) );
  NANDN U24963 ( .A(y[660]), .B(x[660]), .Z(n10310) );
  NANDN U24964 ( .A(y[661]), .B(x[661]), .Z(n10309) );
  AND U24965 ( .A(n10310), .B(n10309), .Z(n52589) );
  NANDN U24966 ( .A(x[660]), .B(y[660]), .Z(n10312) );
  NANDN U24967 ( .A(x[659]), .B(y[659]), .Z(n10311) );
  NAND U24968 ( .A(n10312), .B(n10311), .Z(n52588) );
  NANDN U24969 ( .A(x[657]), .B(y[657]), .Z(n10313) );
  ANDN U24970 ( .B(y[658]), .A(x[658]), .Z(n30781) );
  ANDN U24971 ( .B(n10313), .A(n30781), .Z(n52586) );
  NANDN U24972 ( .A(y[656]), .B(x[656]), .Z(n30776) );
  NANDN U24973 ( .A(y[657]), .B(x[657]), .Z(n10314) );
  NAND U24974 ( .A(n30776), .B(n10314), .Z(n52585) );
  ANDN U24975 ( .B(y[655]), .A(x[655]), .Z(n30771) );
  ANDN U24976 ( .B(y[656]), .A(x[656]), .Z(n30780) );
  NOR U24977 ( .A(n30771), .B(n30780), .Z(n52584) );
  NANDN U24978 ( .A(y[654]), .B(x[654]), .Z(n30768) );
  NANDN U24979 ( .A(y[655]), .B(x[655]), .Z(n30775) );
  NAND U24980 ( .A(n30768), .B(n30775), .Z(n52582) );
  ANDN U24981 ( .B(y[653]), .A(x[653]), .Z(n30764) );
  ANDN U24982 ( .B(y[654]), .A(x[654]), .Z(n30774) );
  NOR U24983 ( .A(n30764), .B(n30774), .Z(n52581) );
  NANDN U24984 ( .A(y[652]), .B(x[652]), .Z(n30760) );
  NANDN U24985 ( .A(y[653]), .B(x[653]), .Z(n30769) );
  NAND U24986 ( .A(n30760), .B(n30769), .Z(n52580) );
  XNOR U24987 ( .A(y[652]), .B(x[652]), .Z(n10315) );
  ANDN U24988 ( .B(y[651]), .A(x[651]), .Z(n30755) );
  ANDN U24989 ( .B(n10315), .A(n30755), .Z(n52579) );
  NANDN U24990 ( .A(y[650]), .B(x[650]), .Z(n30752) );
  NANDN U24991 ( .A(y[651]), .B(x[651]), .Z(n30759) );
  NAND U24992 ( .A(n30752), .B(n30759), .Z(n52578) );
  ANDN U24993 ( .B(y[649]), .A(x[649]), .Z(n30750) );
  ANDN U24994 ( .B(y[650]), .A(x[650]), .Z(n30758) );
  NOR U24995 ( .A(n30750), .B(n30758), .Z(n52577) );
  NANDN U24996 ( .A(y[648]), .B(x[648]), .Z(n28278) );
  NANDN U24997 ( .A(y[649]), .B(x[649]), .Z(n30753) );
  NAND U24998 ( .A(n28278), .B(n30753), .Z(n52576) );
  ANDN U24999 ( .B(y[647]), .A(x[647]), .Z(n30743) );
  ANDN U25000 ( .B(y[648]), .A(x[648]), .Z(n30747) );
  NOR U25001 ( .A(n30743), .B(n30747), .Z(n52575) );
  NANDN U25002 ( .A(y[646]), .B(x[646]), .Z(n30739) );
  NANDN U25003 ( .A(y[647]), .B(x[647]), .Z(n28277) );
  NAND U25004 ( .A(n30739), .B(n28277), .Z(n52574) );
  NANDN U25005 ( .A(x[645]), .B(y[645]), .Z(n28279) );
  ANDN U25006 ( .B(y[646]), .A(x[646]), .Z(n52573) );
  ANDN U25007 ( .B(n28279), .A(n52573), .Z(n11622) );
  NANDN U25008 ( .A(y[644]), .B(x[644]), .Z(n52572) );
  NANDN U25009 ( .A(y[645]), .B(x[645]), .Z(n52427) );
  NAND U25010 ( .A(n52572), .B(n52427), .Z(n11620) );
  NANDN U25011 ( .A(x[644]), .B(y[644]), .Z(n28280) );
  ANDN U25012 ( .B(y[643]), .A(x[643]), .Z(n52571) );
  ANDN U25013 ( .B(n28280), .A(n52571), .Z(n11618) );
  NANDN U25014 ( .A(y[642]), .B(x[642]), .Z(n10316) );
  NANDN U25015 ( .A(y[643]), .B(x[643]), .Z(n30735) );
  NAND U25016 ( .A(n10316), .B(n30735), .Z(n52570) );
  XNOR U25017 ( .A(y[642]), .B(x[642]), .Z(n30729) );
  ANDN U25018 ( .B(y[641]), .A(x[641]), .Z(n30727) );
  ANDN U25019 ( .B(n30729), .A(n30727), .Z(n52569) );
  NANDN U25020 ( .A(y[640]), .B(x[640]), .Z(n28282) );
  NANDN U25021 ( .A(y[641]), .B(x[641]), .Z(n30730) );
  NAND U25022 ( .A(n28282), .B(n30730), .Z(n52568) );
  ANDN U25023 ( .B(y[639]), .A(x[639]), .Z(n30719) );
  ANDN U25024 ( .B(y[640]), .A(x[640]), .Z(n30724) );
  NOR U25025 ( .A(n30719), .B(n30724), .Z(n52566) );
  NANDN U25026 ( .A(y[638]), .B(x[638]), .Z(n30715) );
  NANDN U25027 ( .A(y[639]), .B(x[639]), .Z(n28281) );
  NAND U25028 ( .A(n30715), .B(n28281), .Z(n52564) );
  ANDN U25029 ( .B(y[637]), .A(x[637]), .Z(n30710) );
  ANDN U25030 ( .B(y[638]), .A(x[638]), .Z(n30720) );
  NOR U25031 ( .A(n30710), .B(n30720), .Z(n52562) );
  NANDN U25032 ( .A(y[636]), .B(x[636]), .Z(n30707) );
  NANDN U25033 ( .A(y[637]), .B(x[637]), .Z(n30714) );
  NAND U25034 ( .A(n30707), .B(n30714), .Z(n52560) );
  ANDN U25035 ( .B(y[635]), .A(x[635]), .Z(n30705) );
  ANDN U25036 ( .B(y[636]), .A(x[636]), .Z(n30713) );
  NOR U25037 ( .A(n30705), .B(n30713), .Z(n52558) );
  NANDN U25038 ( .A(y[634]), .B(x[634]), .Z(n28284) );
  NANDN U25039 ( .A(y[635]), .B(x[635]), .Z(n30708) );
  NAND U25040 ( .A(n28284), .B(n30708), .Z(n52556) );
  ANDN U25041 ( .B(y[633]), .A(x[633]), .Z(n30697) );
  ANDN U25042 ( .B(y[634]), .A(x[634]), .Z(n30702) );
  NOR U25043 ( .A(n30697), .B(n30702), .Z(n52554) );
  NANDN U25044 ( .A(y[632]), .B(x[632]), .Z(n30693) );
  NANDN U25045 ( .A(y[633]), .B(x[633]), .Z(n28283) );
  NAND U25046 ( .A(n30693), .B(n28283), .Z(n52552) );
  ANDN U25047 ( .B(y[631]), .A(x[631]), .Z(n30688) );
  ANDN U25048 ( .B(y[632]), .A(x[632]), .Z(n30698) );
  NOR U25049 ( .A(n30688), .B(n30698), .Z(n52550) );
  NANDN U25050 ( .A(y[630]), .B(x[630]), .Z(n30685) );
  NANDN U25051 ( .A(y[631]), .B(x[631]), .Z(n30692) );
  NAND U25052 ( .A(n30685), .B(n30692), .Z(n52548) );
  XNOR U25053 ( .A(x[630]), .B(y[630]), .Z(n10317) );
  ANDN U25054 ( .B(y[629]), .A(x[629]), .Z(n30683) );
  ANDN U25055 ( .B(n10317), .A(n30683), .Z(n52546) );
  NANDN U25056 ( .A(y[628]), .B(x[628]), .Z(n28286) );
  NANDN U25057 ( .A(y[629]), .B(x[629]), .Z(n30686) );
  NAND U25058 ( .A(n28286), .B(n30686), .Z(n52544) );
  XNOR U25059 ( .A(y[628]), .B(x[628]), .Z(n10318) );
  ANDN U25060 ( .B(y[627]), .A(x[627]), .Z(n30675) );
  ANDN U25061 ( .B(n10318), .A(n30675), .Z(n52542) );
  NANDN U25062 ( .A(y[626]), .B(x[626]), .Z(n30671) );
  NANDN U25063 ( .A(y[627]), .B(x[627]), .Z(n28285) );
  NAND U25064 ( .A(n30671), .B(n28285), .Z(n52540) );
  ANDN U25065 ( .B(y[625]), .A(x[625]), .Z(n30666) );
  ANDN U25066 ( .B(y[626]), .A(x[626]), .Z(n30676) );
  NOR U25067 ( .A(n30666), .B(n30676), .Z(n52538) );
  NANDN U25068 ( .A(y[624]), .B(x[624]), .Z(n30663) );
  NANDN U25069 ( .A(y[625]), .B(x[625]), .Z(n30670) );
  NAND U25070 ( .A(n30663), .B(n30670), .Z(n52536) );
  ANDN U25071 ( .B(y[623]), .A(x[623]), .Z(n30661) );
  ANDN U25072 ( .B(y[624]), .A(x[624]), .Z(n30669) );
  NOR U25073 ( .A(n30661), .B(n30669), .Z(n52534) );
  NANDN U25074 ( .A(y[622]), .B(x[622]), .Z(n28288) );
  NANDN U25075 ( .A(y[623]), .B(x[623]), .Z(n30664) );
  NAND U25076 ( .A(n28288), .B(n30664), .Z(n52532) );
  NANDN U25077 ( .A(x[621]), .B(y[621]), .Z(n30653) );
  XNOR U25078 ( .A(x[622]), .B(y[622]), .Z(n10319) );
  AND U25079 ( .A(n30653), .B(n10319), .Z(n52530) );
  NANDN U25080 ( .A(y[620]), .B(x[620]), .Z(n30651) );
  NANDN U25081 ( .A(y[621]), .B(x[621]), .Z(n28287) );
  NAND U25082 ( .A(n30651), .B(n28287), .Z(n52528) );
  XNOR U25083 ( .A(y[620]), .B(x[620]), .Z(n10320) );
  ANDN U25084 ( .B(y[619]), .A(x[619]), .Z(n30648) );
  ANDN U25085 ( .B(n10320), .A(n30648), .Z(n52526) );
  NANDN U25086 ( .A(y[619]), .B(x[619]), .Z(n52525) );
  NANDN U25087 ( .A(x[617]), .B(y[617]), .Z(n28291) );
  NANDN U25088 ( .A(y[616]), .B(x[616]), .Z(n28294) );
  NANDN U25089 ( .A(x[614]), .B(y[614]), .Z(n30641) );
  ANDN U25090 ( .B(y[613]), .A(x[613]), .Z(n30637) );
  ANDN U25091 ( .B(n30641), .A(n30637), .Z(n52518) );
  NANDN U25092 ( .A(x[611]), .B(y[611]), .Z(n28297) );
  ANDN U25093 ( .B(y[612]), .A(x[612]), .Z(n52516) );
  ANDN U25094 ( .B(n28297), .A(n52516), .Z(n11579) );
  ANDN U25095 ( .B(x[610]), .A(y[610]), .Z(n11576) );
  ANDN U25096 ( .B(y[609]), .A(x[609]), .Z(n52513) );
  XNOR U25097 ( .A(x[610]), .B(y[610]), .Z(n28301) );
  ANDN U25098 ( .B(x[608]), .A(y[608]), .Z(n52512) );
  XNOR U25099 ( .A(y[608]), .B(x[608]), .Z(n30626) );
  ANDN U25100 ( .B(y[607]), .A(x[607]), .Z(n30625) );
  ANDN U25101 ( .B(n30626), .A(n30625), .Z(n52511) );
  NANDN U25102 ( .A(y[607]), .B(x[607]), .Z(n52510) );
  NANDN U25103 ( .A(x[604]), .B(y[604]), .Z(n28305) );
  ANDN U25104 ( .B(y[603]), .A(x[603]), .Z(n52505) );
  ANDN U25105 ( .B(n28305), .A(n52505), .Z(n11563) );
  NANDN U25106 ( .A(y[602]), .B(x[602]), .Z(n52504) );
  XNOR U25107 ( .A(y[602]), .B(x[602]), .Z(n10321) );
  ANDN U25108 ( .B(y[601]), .A(x[601]), .Z(n30614) );
  ANDN U25109 ( .B(n10321), .A(n30614), .Z(n52503) );
  NANDN U25110 ( .A(y[601]), .B(x[601]), .Z(n52502) );
  NANDN U25111 ( .A(x[599]), .B(y[599]), .Z(n28313) );
  ANDN U25112 ( .B(x[598]), .A(y[598]), .Z(n28314) );
  ANDN U25113 ( .B(y[595]), .A(x[595]), .Z(n30602) );
  ANDN U25114 ( .B(y[596]), .A(x[596]), .Z(n30607) );
  NOR U25115 ( .A(n30602), .B(n30607), .Z(n52495) );
  NANDN U25116 ( .A(x[593]), .B(y[593]), .Z(n30597) );
  ANDN U25117 ( .B(y[594]), .A(x[594]), .Z(n52493) );
  ANDN U25118 ( .B(n30597), .A(n52493), .Z(n11545) );
  ANDN U25119 ( .B(x[592]), .A(y[592]), .Z(n28319) );
  NANDN U25120 ( .A(x[592]), .B(y[592]), .Z(n30598) );
  NANDN U25121 ( .A(y[590]), .B(x[590]), .Z(n52488) );
  NANDN U25122 ( .A(x[589]), .B(y[589]), .Z(n30589) );
  ANDN U25123 ( .B(y[590]), .A(x[590]), .Z(n30595) );
  ANDN U25124 ( .B(n30589), .A(n30595), .Z(n52487) );
  ANDN U25125 ( .B(x[589]), .A(y[589]), .Z(n52486) );
  NANDN U25126 ( .A(x[588]), .B(y[588]), .Z(n52485) );
  NANDN U25127 ( .A(x[586]), .B(y[586]), .Z(n28325) );
  NANDN U25128 ( .A(x[585]), .B(y[585]), .Z(n52481) );
  AND U25129 ( .A(n28325), .B(n52481), .Z(n11530) );
  NANDN U25130 ( .A(y[584]), .B(x[584]), .Z(n52480) );
  NANDN U25131 ( .A(x[584]), .B(y[584]), .Z(n30583) );
  ANDN U25132 ( .B(y[583]), .A(x[583]), .Z(n30579) );
  ANDN U25133 ( .B(n30583), .A(n30579), .Z(n52479) );
  ANDN U25134 ( .B(x[582]), .A(y[582]), .Z(n28329) );
  NANDN U25135 ( .A(x[581]), .B(y[581]), .Z(n28332) );
  ANDN U25136 ( .B(x[580]), .A(y[580]), .Z(n28334) );
  XNOR U25137 ( .A(y[578]), .B(x[578]), .Z(n30569) );
  ANDN U25138 ( .B(y[577]), .A(x[577]), .Z(n30567) );
  ANDN U25139 ( .B(n30569), .A(n30567), .Z(n52471) );
  NANDN U25140 ( .A(x[575]), .B(y[575]), .Z(n28339) );
  ANDN U25141 ( .B(y[576]), .A(x[576]), .Z(n52469) );
  ANDN U25142 ( .B(n28339), .A(n52469), .Z(n11512) );
  NANDN U25143 ( .A(y[574]), .B(x[574]), .Z(n28342) );
  NANDN U25144 ( .A(x[574]), .B(y[574]), .Z(n28340) );
  ANDN U25145 ( .B(x[573]), .A(y[573]), .Z(n28341) );
  NANDN U25146 ( .A(x[572]), .B(y[572]), .Z(n28344) );
  ANDN U25147 ( .B(y[571]), .A(x[571]), .Z(n30558) );
  NANDN U25148 ( .A(y[572]), .B(x[572]), .Z(n10323) );
  NAND U25149 ( .A(n30558), .B(n10323), .Z(n52435) );
  ANDN U25150 ( .B(x[570]), .A(y[570]), .Z(n28345) );
  NANDN U25151 ( .A(y[571]), .B(x[571]), .Z(n10322) );
  AND U25152 ( .A(n10323), .B(n10322), .Z(n52466) );
  NANDN U25153 ( .A(x[568]), .B(y[568]), .Z(n30553) );
  ANDN U25154 ( .B(y[567]), .A(x[567]), .Z(n52462) );
  ANDN U25155 ( .B(n30553), .A(n52462), .Z(n11497) );
  NANDN U25156 ( .A(y[566]), .B(x[566]), .Z(n52460) );
  XNOR U25157 ( .A(y[566]), .B(x[566]), .Z(n10324) );
  ANDN U25158 ( .B(y[565]), .A(x[565]), .Z(n30545) );
  ANDN U25159 ( .B(n10324), .A(n30545), .Z(n52459) );
  NANDN U25160 ( .A(y[565]), .B(x[565]), .Z(n52458) );
  NANDN U25161 ( .A(x[563]), .B(y[563]), .Z(n30541) );
  ANDN U25162 ( .B(x[562]), .A(y[562]), .Z(n28353) );
  XNOR U25163 ( .A(y[560]), .B(x[560]), .Z(n10325) );
  ANDN U25164 ( .B(y[559]), .A(x[559]), .Z(n30532) );
  ANDN U25165 ( .B(n10325), .A(n30532), .Z(n52452) );
  NANDN U25166 ( .A(x[557]), .B(y[557]), .Z(n30527) );
  ANDN U25167 ( .B(y[558]), .A(x[558]), .Z(n52450) );
  ANDN U25168 ( .B(n30527), .A(n52450), .Z(n11479) );
  ANDN U25169 ( .B(x[556]), .A(y[556]), .Z(n11476) );
  ANDN U25170 ( .B(y[555]), .A(x[555]), .Z(n52446) );
  XNOR U25171 ( .A(x[556]), .B(y[556]), .Z(n28359) );
  NANDN U25172 ( .A(y[554]), .B(x[554]), .Z(n52445) );
  ANDN U25173 ( .B(y[553]), .A(x[553]), .Z(n30520) );
  ANDN U25174 ( .B(y[554]), .A(x[554]), .Z(n30525) );
  NOR U25175 ( .A(n30520), .B(n30525), .Z(n52444) );
  NANDN U25176 ( .A(y[552]), .B(x[552]), .Z(n28361) );
  ANDN U25177 ( .B(x[551]), .A(y[551]), .Z(n28360) );
  NANDN U25178 ( .A(y[550]), .B(x[550]), .Z(n10327) );
  NANDN U25179 ( .A(y[549]), .B(x[549]), .Z(n10326) );
  AND U25180 ( .A(n10327), .B(n10326), .Z(n30514) );
  NANDN U25181 ( .A(x[547]), .B(y[547]), .Z(n28367) );
  ANDN U25182 ( .B(x[546]), .A(y[546]), .Z(n30503) );
  NANDN U25183 ( .A(x[545]), .B(y[545]), .Z(n30499) );
  ANDN U25184 ( .B(x[544]), .A(y[544]), .Z(n30494) );
  NANDN U25185 ( .A(x[544]), .B(y[544]), .Z(n30498) );
  NANDN U25186 ( .A(y[542]), .B(x[542]), .Z(n11449) );
  XOR U25187 ( .A(y[542]), .B(x[542]), .Z(n30487) );
  ANDN U25188 ( .B(x[540]), .A(y[540]), .Z(n30481) );
  ANDN U25189 ( .B(x[538]), .A(y[538]), .Z(n30475) );
  ANDN U25190 ( .B(x[539]), .A(y[539]), .Z(n30482) );
  NOR U25191 ( .A(n30475), .B(n30482), .Z(n11440) );
  NANDN U25192 ( .A(x[538]), .B(y[538]), .Z(n30476) );
  NANDN U25193 ( .A(y[537]), .B(x[537]), .Z(n10329) );
  NANDN U25194 ( .A(y[536]), .B(x[536]), .Z(n10328) );
  NAND U25195 ( .A(n10329), .B(n10328), .Z(n30471) );
  NANDN U25196 ( .A(x[533]), .B(y[533]), .Z(n10331) );
  NANDN U25197 ( .A(x[534]), .B(y[534]), .Z(n10330) );
  AND U25198 ( .A(n10331), .B(n10330), .Z(n30465) );
  NANDN U25199 ( .A(y[533]), .B(x[533]), .Z(n10333) );
  NANDN U25200 ( .A(y[532]), .B(x[532]), .Z(n10332) );
  NAND U25201 ( .A(n10333), .B(n10332), .Z(n30463) );
  NANDN U25202 ( .A(x[531]), .B(y[531]), .Z(n10335) );
  NANDN U25203 ( .A(x[532]), .B(y[532]), .Z(n10334) );
  AND U25204 ( .A(n10335), .B(n10334), .Z(n30461) );
  NANDN U25205 ( .A(y[531]), .B(x[531]), .Z(n10337) );
  NANDN U25206 ( .A(y[530]), .B(x[530]), .Z(n10336) );
  NAND U25207 ( .A(n10337), .B(n10336), .Z(n30459) );
  NANDN U25208 ( .A(x[527]), .B(y[527]), .Z(n10339) );
  NANDN U25209 ( .A(x[528]), .B(y[528]), .Z(n10338) );
  AND U25210 ( .A(n10339), .B(n10338), .Z(n30453) );
  NANDN U25211 ( .A(y[526]), .B(x[526]), .Z(n10340) );
  ANDN U25212 ( .B(x[527]), .A(y[527]), .Z(n30446) );
  ANDN U25213 ( .B(n10340), .A(n30446), .Z(n11418) );
  NANDN U25214 ( .A(x[525]), .B(y[525]), .Z(n30441) );
  ANDN U25215 ( .B(x[524]), .A(y[524]), .Z(n30436) );
  ANDN U25216 ( .B(x[523]), .A(y[523]), .Z(n30439) );
  ANDN U25217 ( .B(x[522]), .A(y[522]), .Z(n30431) );
  NOR U25218 ( .A(n30439), .B(n30431), .Z(n11409) );
  NANDN U25219 ( .A(x[522]), .B(y[522]), .Z(n30434) );
  ANDN U25220 ( .B(x[520]), .A(y[520]), .Z(n30423) );
  NANDN U25221 ( .A(x[519]), .B(y[519]), .Z(n30419) );
  ANDN U25222 ( .B(x[518]), .A(y[518]), .Z(n30414) );
  ANDN U25223 ( .B(x[517]), .A(y[517]), .Z(n30417) );
  ANDN U25224 ( .B(x[516]), .A(y[516]), .Z(n30409) );
  NOR U25225 ( .A(n30417), .B(n30409), .Z(n11397) );
  NANDN U25226 ( .A(x[516]), .B(y[516]), .Z(n30412) );
  ANDN U25227 ( .B(x[514]), .A(y[514]), .Z(n30401) );
  NANDN U25228 ( .A(x[513]), .B(y[513]), .Z(n30397) );
  ANDN U25229 ( .B(x[512]), .A(y[512]), .Z(n30392) );
  ANDN U25230 ( .B(x[511]), .A(y[511]), .Z(n30395) );
  ANDN U25231 ( .B(x[510]), .A(y[510]), .Z(n30387) );
  NOR U25232 ( .A(n30395), .B(n30387), .Z(n11385) );
  NANDN U25233 ( .A(x[510]), .B(y[510]), .Z(n30390) );
  ANDN U25234 ( .B(x[508]), .A(y[508]), .Z(n30379) );
  NANDN U25235 ( .A(x[507]), .B(y[507]), .Z(n30375) );
  ANDN U25236 ( .B(x[506]), .A(y[506]), .Z(n30370) );
  ANDN U25237 ( .B(x[505]), .A(y[505]), .Z(n30373) );
  ANDN U25238 ( .B(x[504]), .A(y[504]), .Z(n30365) );
  NOR U25239 ( .A(n30373), .B(n30365), .Z(n11373) );
  NANDN U25240 ( .A(x[504]), .B(y[504]), .Z(n30368) );
  ANDN U25241 ( .B(x[502]), .A(y[502]), .Z(n30357) );
  NANDN U25242 ( .A(x[501]), .B(y[501]), .Z(n30353) );
  ANDN U25243 ( .B(x[500]), .A(y[500]), .Z(n30348) );
  ANDN U25244 ( .B(x[499]), .A(y[499]), .Z(n30351) );
  ANDN U25245 ( .B(x[498]), .A(y[498]), .Z(n30343) );
  NOR U25246 ( .A(n30351), .B(n30343), .Z(n11361) );
  NANDN U25247 ( .A(x[498]), .B(y[498]), .Z(n30346) );
  ANDN U25248 ( .B(x[496]), .A(y[496]), .Z(n30335) );
  NANDN U25249 ( .A(x[495]), .B(y[495]), .Z(n30331) );
  ANDN U25250 ( .B(x[494]), .A(y[494]), .Z(n30326) );
  ANDN U25251 ( .B(x[493]), .A(y[493]), .Z(n30329) );
  ANDN U25252 ( .B(x[492]), .A(y[492]), .Z(n30321) );
  NOR U25253 ( .A(n30329), .B(n30321), .Z(n11349) );
  NANDN U25254 ( .A(x[492]), .B(y[492]), .Z(n30324) );
  ANDN U25255 ( .B(x[490]), .A(y[490]), .Z(n30313) );
  NANDN U25256 ( .A(x[489]), .B(y[489]), .Z(n30309) );
  ANDN U25257 ( .B(x[488]), .A(y[488]), .Z(n30304) );
  ANDN U25258 ( .B(x[487]), .A(y[487]), .Z(n30307) );
  ANDN U25259 ( .B(x[486]), .A(y[486]), .Z(n30299) );
  NOR U25260 ( .A(n30307), .B(n30299), .Z(n11337) );
  NANDN U25261 ( .A(x[486]), .B(y[486]), .Z(n30302) );
  ANDN U25262 ( .B(x[484]), .A(y[484]), .Z(n30291) );
  NANDN U25263 ( .A(x[483]), .B(y[483]), .Z(n30287) );
  ANDN U25264 ( .B(x[482]), .A(y[482]), .Z(n30282) );
  ANDN U25265 ( .B(x[481]), .A(y[481]), .Z(n30285) );
  ANDN U25266 ( .B(x[480]), .A(y[480]), .Z(n30277) );
  NOR U25267 ( .A(n30285), .B(n30277), .Z(n11325) );
  NANDN U25268 ( .A(x[480]), .B(y[480]), .Z(n30280) );
  ANDN U25269 ( .B(x[478]), .A(y[478]), .Z(n30269) );
  NANDN U25270 ( .A(x[477]), .B(y[477]), .Z(n30265) );
  ANDN U25271 ( .B(x[476]), .A(y[476]), .Z(n30260) );
  ANDN U25272 ( .B(x[475]), .A(y[475]), .Z(n30263) );
  ANDN U25273 ( .B(x[474]), .A(y[474]), .Z(n30255) );
  NOR U25274 ( .A(n30263), .B(n30255), .Z(n11313) );
  NANDN U25275 ( .A(x[474]), .B(y[474]), .Z(n30258) );
  ANDN U25276 ( .B(x[472]), .A(y[472]), .Z(n30247) );
  NANDN U25277 ( .A(x[471]), .B(y[471]), .Z(n30243) );
  ANDN U25278 ( .B(x[470]), .A(y[470]), .Z(n30238) );
  ANDN U25279 ( .B(x[469]), .A(y[469]), .Z(n30241) );
  ANDN U25280 ( .B(x[468]), .A(y[468]), .Z(n30233) );
  NOR U25281 ( .A(n30241), .B(n30233), .Z(n11301) );
  NANDN U25282 ( .A(x[468]), .B(y[468]), .Z(n30236) );
  ANDN U25283 ( .B(x[466]), .A(y[466]), .Z(n30225) );
  NANDN U25284 ( .A(x[465]), .B(y[465]), .Z(n30221) );
  ANDN U25285 ( .B(x[464]), .A(y[464]), .Z(n30216) );
  ANDN U25286 ( .B(x[463]), .A(y[463]), .Z(n30219) );
  ANDN U25287 ( .B(x[462]), .A(y[462]), .Z(n30211) );
  NOR U25288 ( .A(n30219), .B(n30211), .Z(n11289) );
  NANDN U25289 ( .A(x[462]), .B(y[462]), .Z(n30214) );
  ANDN U25290 ( .B(x[460]), .A(y[460]), .Z(n30203) );
  NANDN U25291 ( .A(x[459]), .B(y[459]), .Z(n30199) );
  ANDN U25292 ( .B(x[458]), .A(y[458]), .Z(n30194) );
  ANDN U25293 ( .B(x[457]), .A(y[457]), .Z(n30197) );
  ANDN U25294 ( .B(x[456]), .A(y[456]), .Z(n30189) );
  NOR U25295 ( .A(n30197), .B(n30189), .Z(n11277) );
  NANDN U25296 ( .A(x[456]), .B(y[456]), .Z(n30192) );
  ANDN U25297 ( .B(x[454]), .A(y[454]), .Z(n30181) );
  NANDN U25298 ( .A(x[453]), .B(y[453]), .Z(n30177) );
  ANDN U25299 ( .B(x[452]), .A(y[452]), .Z(n30172) );
  ANDN U25300 ( .B(x[451]), .A(y[451]), .Z(n30175) );
  ANDN U25301 ( .B(x[450]), .A(y[450]), .Z(n30167) );
  NOR U25302 ( .A(n30175), .B(n30167), .Z(n11265) );
  NANDN U25303 ( .A(x[450]), .B(y[450]), .Z(n30170) );
  ANDN U25304 ( .B(x[448]), .A(y[448]), .Z(n30159) );
  NANDN U25305 ( .A(x[447]), .B(y[447]), .Z(n30155) );
  ANDN U25306 ( .B(x[446]), .A(y[446]), .Z(n30150) );
  ANDN U25307 ( .B(x[445]), .A(y[445]), .Z(n30153) );
  ANDN U25308 ( .B(x[444]), .A(y[444]), .Z(n30145) );
  NOR U25309 ( .A(n30153), .B(n30145), .Z(n11253) );
  NANDN U25310 ( .A(x[444]), .B(y[444]), .Z(n30148) );
  ANDN U25311 ( .B(x[442]), .A(y[442]), .Z(n30137) );
  NANDN U25312 ( .A(x[441]), .B(y[441]), .Z(n30133) );
  ANDN U25313 ( .B(x[440]), .A(y[440]), .Z(n30128) );
  ANDN U25314 ( .B(x[439]), .A(y[439]), .Z(n30131) );
  ANDN U25315 ( .B(x[438]), .A(y[438]), .Z(n30123) );
  NOR U25316 ( .A(n30131), .B(n30123), .Z(n11241) );
  NANDN U25317 ( .A(x[438]), .B(y[438]), .Z(n30126) );
  ANDN U25318 ( .B(x[436]), .A(y[436]), .Z(n30115) );
  NANDN U25319 ( .A(x[435]), .B(y[435]), .Z(n30111) );
  ANDN U25320 ( .B(x[434]), .A(y[434]), .Z(n30106) );
  NANDN U25321 ( .A(y[432]), .B(x[432]), .Z(n10341) );
  ANDN U25322 ( .B(x[433]), .A(y[433]), .Z(n30109) );
  ANDN U25323 ( .B(n10341), .A(n30109), .Z(n11229) );
  XOR U25324 ( .A(y[432]), .B(x[432]), .Z(n30099) );
  ANDN U25325 ( .B(x[431]), .A(y[431]), .Z(n30101) );
  NANDN U25326 ( .A(x[429]), .B(y[429]), .Z(n30089) );
  ANDN U25327 ( .B(x[428]), .A(y[428]), .Z(n30084) );
  ANDN U25328 ( .B(x[427]), .A(y[427]), .Z(n30087) );
  ANDN U25329 ( .B(x[426]), .A(y[426]), .Z(n30079) );
  NOR U25330 ( .A(n30087), .B(n30079), .Z(n11217) );
  NANDN U25331 ( .A(x[426]), .B(y[426]), .Z(n30082) );
  ANDN U25332 ( .B(x[424]), .A(y[424]), .Z(n30071) );
  NANDN U25333 ( .A(x[423]), .B(y[423]), .Z(n30067) );
  ANDN U25334 ( .B(x[422]), .A(y[422]), .Z(n30062) );
  ANDN U25335 ( .B(x[421]), .A(y[421]), .Z(n30065) );
  ANDN U25336 ( .B(x[420]), .A(y[420]), .Z(n30057) );
  NOR U25337 ( .A(n30065), .B(n30057), .Z(n11205) );
  NANDN U25338 ( .A(x[420]), .B(y[420]), .Z(n30060) );
  ANDN U25339 ( .B(x[418]), .A(y[418]), .Z(n30049) );
  NANDN U25340 ( .A(x[417]), .B(y[417]), .Z(n30045) );
  ANDN U25341 ( .B(x[416]), .A(y[416]), .Z(n30040) );
  ANDN U25342 ( .B(x[415]), .A(y[415]), .Z(n30043) );
  ANDN U25343 ( .B(x[414]), .A(y[414]), .Z(n30035) );
  NOR U25344 ( .A(n30043), .B(n30035), .Z(n11193) );
  NANDN U25345 ( .A(x[414]), .B(y[414]), .Z(n30038) );
  ANDN U25346 ( .B(x[412]), .A(y[412]), .Z(n30027) );
  NANDN U25347 ( .A(x[411]), .B(y[411]), .Z(n30023) );
  ANDN U25348 ( .B(x[410]), .A(y[410]), .Z(n30018) );
  ANDN U25349 ( .B(x[409]), .A(y[409]), .Z(n30021) );
  ANDN U25350 ( .B(x[408]), .A(y[408]), .Z(n30013) );
  NOR U25351 ( .A(n30021), .B(n30013), .Z(n11181) );
  NANDN U25352 ( .A(x[408]), .B(y[408]), .Z(n30016) );
  ANDN U25353 ( .B(x[406]), .A(y[406]), .Z(n30005) );
  NANDN U25354 ( .A(x[405]), .B(y[405]), .Z(n30001) );
  ANDN U25355 ( .B(x[404]), .A(y[404]), .Z(n29996) );
  ANDN U25356 ( .B(x[403]), .A(y[403]), .Z(n29999) );
  ANDN U25357 ( .B(x[402]), .A(y[402]), .Z(n29991) );
  NOR U25358 ( .A(n29999), .B(n29991), .Z(n11169) );
  NANDN U25359 ( .A(x[402]), .B(y[402]), .Z(n29994) );
  ANDN U25360 ( .B(x[400]), .A(y[400]), .Z(n29983) );
  NANDN U25361 ( .A(x[399]), .B(y[399]), .Z(n29979) );
  ANDN U25362 ( .B(x[398]), .A(y[398]), .Z(n29974) );
  ANDN U25363 ( .B(x[397]), .A(y[397]), .Z(n29977) );
  ANDN U25364 ( .B(x[396]), .A(y[396]), .Z(n29969) );
  NOR U25365 ( .A(n29977), .B(n29969), .Z(n11157) );
  NANDN U25366 ( .A(x[396]), .B(y[396]), .Z(n29972) );
  ANDN U25367 ( .B(x[394]), .A(y[394]), .Z(n29961) );
  NANDN U25368 ( .A(x[393]), .B(y[393]), .Z(n29957) );
  ANDN U25369 ( .B(x[392]), .A(y[392]), .Z(n29952) );
  ANDN U25370 ( .B(x[391]), .A(y[391]), .Z(n29955) );
  ANDN U25371 ( .B(x[390]), .A(y[390]), .Z(n29947) );
  NOR U25372 ( .A(n29955), .B(n29947), .Z(n11145) );
  NANDN U25373 ( .A(x[390]), .B(y[390]), .Z(n29950) );
  ANDN U25374 ( .B(x[388]), .A(y[388]), .Z(n29939) );
  NANDN U25375 ( .A(x[387]), .B(y[387]), .Z(n29935) );
  ANDN U25376 ( .B(x[386]), .A(y[386]), .Z(n29930) );
  ANDN U25377 ( .B(x[385]), .A(y[385]), .Z(n29933) );
  ANDN U25378 ( .B(x[384]), .A(y[384]), .Z(n29925) );
  NOR U25379 ( .A(n29933), .B(n29925), .Z(n11133) );
  NANDN U25380 ( .A(x[384]), .B(y[384]), .Z(n29928) );
  ANDN U25381 ( .B(x[382]), .A(y[382]), .Z(n29917) );
  NANDN U25382 ( .A(x[381]), .B(y[381]), .Z(n29913) );
  ANDN U25383 ( .B(x[380]), .A(y[380]), .Z(n29908) );
  ANDN U25384 ( .B(x[379]), .A(y[379]), .Z(n29911) );
  ANDN U25385 ( .B(x[378]), .A(y[378]), .Z(n29903) );
  NOR U25386 ( .A(n29911), .B(n29903), .Z(n11121) );
  NANDN U25387 ( .A(x[378]), .B(y[378]), .Z(n29906) );
  ANDN U25388 ( .B(x[376]), .A(y[376]), .Z(n29895) );
  NANDN U25389 ( .A(x[375]), .B(y[375]), .Z(n29891) );
  ANDN U25390 ( .B(x[374]), .A(y[374]), .Z(n29886) );
  ANDN U25391 ( .B(x[373]), .A(y[373]), .Z(n29889) );
  ANDN U25392 ( .B(x[372]), .A(y[372]), .Z(n29881) );
  NOR U25393 ( .A(n29889), .B(n29881), .Z(n11109) );
  NANDN U25394 ( .A(x[372]), .B(y[372]), .Z(n29884) );
  ANDN U25395 ( .B(x[370]), .A(y[370]), .Z(n29873) );
  NANDN U25396 ( .A(x[369]), .B(y[369]), .Z(n29869) );
  ANDN U25397 ( .B(x[368]), .A(y[368]), .Z(n29864) );
  ANDN U25398 ( .B(x[367]), .A(y[367]), .Z(n29867) );
  ANDN U25399 ( .B(x[366]), .A(y[366]), .Z(n29859) );
  NOR U25400 ( .A(n29867), .B(n29859), .Z(n11097) );
  NANDN U25401 ( .A(x[366]), .B(y[366]), .Z(n29862) );
  NANDN U25402 ( .A(y[364]), .B(x[364]), .Z(n11093) );
  XOR U25403 ( .A(y[364]), .B(x[364]), .Z(n29851) );
  ANDN U25404 ( .B(x[362]), .A(y[362]), .Z(n29842) );
  ANDN U25405 ( .B(x[361]), .A(y[361]), .Z(n29845) );
  ANDN U25406 ( .B(x[360]), .A(y[360]), .Z(n29837) );
  NOR U25407 ( .A(n29845), .B(n29837), .Z(n11084) );
  NANDN U25408 ( .A(x[360]), .B(y[360]), .Z(n29840) );
  ANDN U25409 ( .B(x[358]), .A(y[358]), .Z(n29829) );
  NANDN U25410 ( .A(x[357]), .B(y[357]), .Z(n29825) );
  ANDN U25411 ( .B(x[356]), .A(y[356]), .Z(n29820) );
  ANDN U25412 ( .B(x[355]), .A(y[355]), .Z(n29823) );
  ANDN U25413 ( .B(x[354]), .A(y[354]), .Z(n29815) );
  NOR U25414 ( .A(n29823), .B(n29815), .Z(n11072) );
  NANDN U25415 ( .A(x[354]), .B(y[354]), .Z(n29818) );
  ANDN U25416 ( .B(x[352]), .A(y[352]), .Z(n29807) );
  NANDN U25417 ( .A(x[351]), .B(y[351]), .Z(n29803) );
  ANDN U25418 ( .B(x[349]), .A(y[349]), .Z(n29798) );
  ANDN U25419 ( .B(x[348]), .A(y[348]), .Z(n29793) );
  NOR U25420 ( .A(n29798), .B(n29793), .Z(n11059) );
  NANDN U25421 ( .A(x[348]), .B(y[348]), .Z(n29796) );
  ANDN U25422 ( .B(x[346]), .A(y[346]), .Z(n29785) );
  NANDN U25423 ( .A(x[345]), .B(y[345]), .Z(n29781) );
  ANDN U25424 ( .B(x[344]), .A(y[344]), .Z(n29776) );
  ANDN U25425 ( .B(x[343]), .A(y[343]), .Z(n29779) );
  ANDN U25426 ( .B(x[342]), .A(y[342]), .Z(n29771) );
  NOR U25427 ( .A(n29779), .B(n29771), .Z(n11047) );
  NANDN U25428 ( .A(x[342]), .B(y[342]), .Z(n29774) );
  ANDN U25429 ( .B(x[340]), .A(y[340]), .Z(n29763) );
  NANDN U25430 ( .A(x[339]), .B(y[339]), .Z(n29759) );
  ANDN U25431 ( .B(x[337]), .A(y[337]), .Z(n29754) );
  ANDN U25432 ( .B(x[336]), .A(y[336]), .Z(n29749) );
  NOR U25433 ( .A(n29754), .B(n29749), .Z(n11034) );
  NANDN U25434 ( .A(x[336]), .B(y[336]), .Z(n29752) );
  ANDN U25435 ( .B(x[334]), .A(y[334]), .Z(n29741) );
  NANDN U25436 ( .A(x[333]), .B(y[333]), .Z(n29737) );
  ANDN U25437 ( .B(x[332]), .A(y[332]), .Z(n29732) );
  ANDN U25438 ( .B(x[331]), .A(y[331]), .Z(n29735) );
  ANDN U25439 ( .B(x[330]), .A(y[330]), .Z(n29727) );
  NOR U25440 ( .A(n29735), .B(n29727), .Z(n11022) );
  NANDN U25441 ( .A(x[330]), .B(y[330]), .Z(n29730) );
  ANDN U25442 ( .B(x[328]), .A(y[328]), .Z(n29719) );
  NANDN U25443 ( .A(x[327]), .B(y[327]), .Z(n29715) );
  ANDN U25444 ( .B(x[326]), .A(y[326]), .Z(n29710) );
  ANDN U25445 ( .B(x[325]), .A(y[325]), .Z(n29713) );
  ANDN U25446 ( .B(x[324]), .A(y[324]), .Z(n29705) );
  NOR U25447 ( .A(n29713), .B(n29705), .Z(n11010) );
  NANDN U25448 ( .A(x[324]), .B(y[324]), .Z(n29708) );
  ANDN U25449 ( .B(x[322]), .A(y[322]), .Z(n29697) );
  NANDN U25450 ( .A(x[321]), .B(y[321]), .Z(n29693) );
  ANDN U25451 ( .B(x[320]), .A(y[320]), .Z(n29688) );
  ANDN U25452 ( .B(x[319]), .A(y[319]), .Z(n29691) );
  ANDN U25453 ( .B(x[318]), .A(y[318]), .Z(n29683) );
  NOR U25454 ( .A(n29691), .B(n29683), .Z(n10998) );
  NANDN U25455 ( .A(x[318]), .B(y[318]), .Z(n29686) );
  ANDN U25456 ( .B(x[316]), .A(y[316]), .Z(n29675) );
  NANDN U25457 ( .A(x[315]), .B(y[315]), .Z(n29671) );
  ANDN U25458 ( .B(x[314]), .A(y[314]), .Z(n29666) );
  ANDN U25459 ( .B(x[313]), .A(y[313]), .Z(n29669) );
  ANDN U25460 ( .B(x[312]), .A(y[312]), .Z(n29661) );
  NOR U25461 ( .A(n29669), .B(n29661), .Z(n10986) );
  NANDN U25462 ( .A(x[312]), .B(y[312]), .Z(n29664) );
  ANDN U25463 ( .B(x[310]), .A(y[310]), .Z(n29653) );
  NANDN U25464 ( .A(x[309]), .B(y[309]), .Z(n29649) );
  ANDN U25465 ( .B(x[308]), .A(y[308]), .Z(n29644) );
  ANDN U25466 ( .B(x[307]), .A(y[307]), .Z(n29647) );
  ANDN U25467 ( .B(x[306]), .A(y[306]), .Z(n29639) );
  NOR U25468 ( .A(n29647), .B(n29639), .Z(n10974) );
  NANDN U25469 ( .A(x[306]), .B(y[306]), .Z(n29642) );
  ANDN U25470 ( .B(x[304]), .A(y[304]), .Z(n29631) );
  NANDN U25471 ( .A(x[303]), .B(y[303]), .Z(n29627) );
  ANDN U25472 ( .B(x[302]), .A(y[302]), .Z(n29622) );
  ANDN U25473 ( .B(x[301]), .A(y[301]), .Z(n29625) );
  ANDN U25474 ( .B(x[300]), .A(y[300]), .Z(n29617) );
  NOR U25475 ( .A(n29625), .B(n29617), .Z(n10962) );
  NANDN U25476 ( .A(x[300]), .B(y[300]), .Z(n29620) );
  ANDN U25477 ( .B(x[298]), .A(y[298]), .Z(n29609) );
  NANDN U25478 ( .A(x[297]), .B(y[297]), .Z(n29605) );
  ANDN U25479 ( .B(x[296]), .A(y[296]), .Z(n29600) );
  ANDN U25480 ( .B(x[295]), .A(y[295]), .Z(n29603) );
  ANDN U25481 ( .B(x[294]), .A(y[294]), .Z(n29595) );
  NOR U25482 ( .A(n29603), .B(n29595), .Z(n10950) );
  NANDN U25483 ( .A(x[294]), .B(y[294]), .Z(n29598) );
  ANDN U25484 ( .B(x[292]), .A(y[292]), .Z(n29587) );
  NANDN U25485 ( .A(x[291]), .B(y[291]), .Z(n29583) );
  ANDN U25486 ( .B(x[290]), .A(y[290]), .Z(n29578) );
  ANDN U25487 ( .B(x[289]), .A(y[289]), .Z(n29581) );
  ANDN U25488 ( .B(x[288]), .A(y[288]), .Z(n29573) );
  NOR U25489 ( .A(n29581), .B(n29573), .Z(n10938) );
  NANDN U25490 ( .A(x[288]), .B(y[288]), .Z(n29576) );
  ANDN U25491 ( .B(x[286]), .A(y[286]), .Z(n29565) );
  NANDN U25492 ( .A(x[285]), .B(y[285]), .Z(n29561) );
  ANDN U25493 ( .B(x[284]), .A(y[284]), .Z(n29556) );
  ANDN U25494 ( .B(x[283]), .A(y[283]), .Z(n29559) );
  ANDN U25495 ( .B(x[282]), .A(y[282]), .Z(n29551) );
  NOR U25496 ( .A(n29559), .B(n29551), .Z(n10926) );
  NANDN U25497 ( .A(x[282]), .B(y[282]), .Z(n29554) );
  ANDN U25498 ( .B(x[280]), .A(y[280]), .Z(n29543) );
  NANDN U25499 ( .A(x[279]), .B(y[279]), .Z(n29539) );
  ANDN U25500 ( .B(x[278]), .A(y[278]), .Z(n29534) );
  NANDN U25501 ( .A(x[276]), .B(y[276]), .Z(n29532) );
  NANDN U25502 ( .A(y[276]), .B(x[276]), .Z(n10343) );
  NANDN U25503 ( .A(y[275]), .B(x[275]), .Z(n10342) );
  NAND U25504 ( .A(n10343), .B(n10342), .Z(n29529) );
  NANDN U25505 ( .A(x[273]), .B(y[273]), .Z(n29519) );
  ANDN U25506 ( .B(x[272]), .A(y[272]), .Z(n29517) );
  NANDN U25507 ( .A(x[272]), .B(y[272]), .Z(n29520) );
  NANDN U25508 ( .A(y[271]), .B(x[271]), .Z(n10345) );
  NANDN U25509 ( .A(y[270]), .B(x[270]), .Z(n10344) );
  NAND U25510 ( .A(n10345), .B(n10344), .Z(n29513) );
  NANDN U25511 ( .A(x[269]), .B(y[269]), .Z(n10347) );
  NANDN U25512 ( .A(x[270]), .B(y[270]), .Z(n10346) );
  AND U25513 ( .A(n10347), .B(n10346), .Z(n29511) );
  NANDN U25514 ( .A(y[269]), .B(x[269]), .Z(n10349) );
  NANDN U25515 ( .A(y[268]), .B(x[268]), .Z(n10348) );
  NAND U25516 ( .A(n10349), .B(n10348), .Z(n29509) );
  NANDN U25517 ( .A(x[265]), .B(y[265]), .Z(n10351) );
  NANDN U25518 ( .A(x[266]), .B(y[266]), .Z(n10350) );
  AND U25519 ( .A(n10351), .B(n10350), .Z(n29503) );
  NANDN U25520 ( .A(y[264]), .B(x[264]), .Z(n10352) );
  ANDN U25521 ( .B(x[265]), .A(y[265]), .Z(n29496) );
  ANDN U25522 ( .B(n10352), .A(n29496), .Z(n10891) );
  NANDN U25523 ( .A(x[263]), .B(y[263]), .Z(n29491) );
  ANDN U25524 ( .B(x[262]), .A(y[262]), .Z(n29486) );
  ANDN U25525 ( .B(x[261]), .A(y[261]), .Z(n29489) );
  ANDN U25526 ( .B(x[260]), .A(y[260]), .Z(n29481) );
  NOR U25527 ( .A(n29489), .B(n29481), .Z(n10882) );
  NANDN U25528 ( .A(x[260]), .B(y[260]), .Z(n29484) );
  ANDN U25529 ( .B(x[258]), .A(y[258]), .Z(n29473) );
  NANDN U25530 ( .A(x[257]), .B(y[257]), .Z(n29469) );
  ANDN U25531 ( .B(x[256]), .A(y[256]), .Z(n29464) );
  ANDN U25532 ( .B(x[255]), .A(y[255]), .Z(n29467) );
  ANDN U25533 ( .B(x[254]), .A(y[254]), .Z(n29459) );
  NOR U25534 ( .A(n29467), .B(n29459), .Z(n10870) );
  NANDN U25535 ( .A(x[254]), .B(y[254]), .Z(n29462) );
  ANDN U25536 ( .B(x[252]), .A(y[252]), .Z(n29451) );
  NANDN U25537 ( .A(x[251]), .B(y[251]), .Z(n29447) );
  ANDN U25538 ( .B(x[250]), .A(y[250]), .Z(n29442) );
  ANDN U25539 ( .B(x[249]), .A(y[249]), .Z(n29445) );
  ANDN U25540 ( .B(x[248]), .A(y[248]), .Z(n29437) );
  NOR U25541 ( .A(n29445), .B(n29437), .Z(n10858) );
  NANDN U25542 ( .A(x[248]), .B(y[248]), .Z(n29440) );
  ANDN U25543 ( .B(x[246]), .A(y[246]), .Z(n29429) );
  NANDN U25544 ( .A(x[245]), .B(y[245]), .Z(n29425) );
  ANDN U25545 ( .B(x[244]), .A(y[244]), .Z(n29420) );
  ANDN U25546 ( .B(x[243]), .A(y[243]), .Z(n29423) );
  ANDN U25547 ( .B(x[242]), .A(y[242]), .Z(n29415) );
  NOR U25548 ( .A(n29423), .B(n29415), .Z(n10846) );
  NANDN U25549 ( .A(x[242]), .B(y[242]), .Z(n29418) );
  ANDN U25550 ( .B(x[240]), .A(y[240]), .Z(n29407) );
  NANDN U25551 ( .A(x[239]), .B(y[239]), .Z(n29403) );
  ANDN U25552 ( .B(x[238]), .A(y[238]), .Z(n29398) );
  ANDN U25553 ( .B(x[237]), .A(y[237]), .Z(n29401) );
  ANDN U25554 ( .B(x[236]), .A(y[236]), .Z(n29393) );
  NOR U25555 ( .A(n29401), .B(n29393), .Z(n10834) );
  NANDN U25556 ( .A(x[236]), .B(y[236]), .Z(n29396) );
  ANDN U25557 ( .B(x[234]), .A(y[234]), .Z(n29385) );
  NANDN U25558 ( .A(x[233]), .B(y[233]), .Z(n29381) );
  ANDN U25559 ( .B(x[232]), .A(y[232]), .Z(n29376) );
  ANDN U25560 ( .B(x[231]), .A(y[231]), .Z(n29379) );
  ANDN U25561 ( .B(x[230]), .A(y[230]), .Z(n29371) );
  NOR U25562 ( .A(n29379), .B(n29371), .Z(n10822) );
  NANDN U25563 ( .A(x[230]), .B(y[230]), .Z(n29374) );
  NANDN U25564 ( .A(y[228]), .B(x[228]), .Z(n10818) );
  XOR U25565 ( .A(y[228]), .B(x[228]), .Z(n29363) );
  ANDN U25566 ( .B(x[226]), .A(y[226]), .Z(n29354) );
  ANDN U25567 ( .B(x[225]), .A(y[225]), .Z(n29357) );
  ANDN U25568 ( .B(x[224]), .A(y[224]), .Z(n29349) );
  NOR U25569 ( .A(n29357), .B(n29349), .Z(n10809) );
  NANDN U25570 ( .A(x[224]), .B(y[224]), .Z(n29352) );
  ANDN U25571 ( .B(x[222]), .A(y[222]), .Z(n29341) );
  NANDN U25572 ( .A(x[221]), .B(y[221]), .Z(n29337) );
  ANDN U25573 ( .B(x[220]), .A(y[220]), .Z(n29332) );
  ANDN U25574 ( .B(x[219]), .A(y[219]), .Z(n29335) );
  ANDN U25575 ( .B(x[218]), .A(y[218]), .Z(n29327) );
  NOR U25576 ( .A(n29335), .B(n29327), .Z(n10797) );
  NANDN U25577 ( .A(x[218]), .B(y[218]), .Z(n29330) );
  ANDN U25578 ( .B(x[216]), .A(y[216]), .Z(n29319) );
  NANDN U25579 ( .A(x[215]), .B(y[215]), .Z(n29315) );
  ANDN U25580 ( .B(x[214]), .A(y[214]), .Z(n29310) );
  ANDN U25581 ( .B(x[213]), .A(y[213]), .Z(n29313) );
  ANDN U25582 ( .B(x[212]), .A(y[212]), .Z(n29305) );
  NOR U25583 ( .A(n29313), .B(n29305), .Z(n10785) );
  NANDN U25584 ( .A(x[212]), .B(y[212]), .Z(n29308) );
  ANDN U25585 ( .B(x[210]), .A(y[210]), .Z(n29297) );
  NANDN U25586 ( .A(x[209]), .B(y[209]), .Z(n29293) );
  ANDN U25587 ( .B(x[208]), .A(y[208]), .Z(n29288) );
  ANDN U25588 ( .B(x[207]), .A(y[207]), .Z(n29291) );
  ANDN U25589 ( .B(x[206]), .A(y[206]), .Z(n29283) );
  NOR U25590 ( .A(n29291), .B(n29283), .Z(n10773) );
  NANDN U25591 ( .A(x[206]), .B(y[206]), .Z(n29286) );
  ANDN U25592 ( .B(x[204]), .A(y[204]), .Z(n29275) );
  NANDN U25593 ( .A(x[203]), .B(y[203]), .Z(n29271) );
  ANDN U25594 ( .B(x[202]), .A(y[202]), .Z(n29266) );
  ANDN U25595 ( .B(x[201]), .A(y[201]), .Z(n29269) );
  ANDN U25596 ( .B(x[200]), .A(y[200]), .Z(n29261) );
  NOR U25597 ( .A(n29269), .B(n29261), .Z(n10761) );
  NANDN U25598 ( .A(x[200]), .B(y[200]), .Z(n29264) );
  ANDN U25599 ( .B(x[198]), .A(y[198]), .Z(n29253) );
  NANDN U25600 ( .A(x[197]), .B(y[197]), .Z(n29249) );
  ANDN U25601 ( .B(x[196]), .A(y[196]), .Z(n29244) );
  NANDN U25602 ( .A(x[194]), .B(y[194]), .Z(n29242) );
  NANDN U25603 ( .A(y[194]), .B(x[194]), .Z(n10354) );
  NANDN U25604 ( .A(y[193]), .B(x[193]), .Z(n10353) );
  NAND U25605 ( .A(n10354), .B(n10353), .Z(n29239) );
  NANDN U25606 ( .A(x[193]), .B(y[193]), .Z(n29236) );
  ANDN U25607 ( .B(x[192]), .A(y[192]), .Z(n29235) );
  NANDN U25608 ( .A(x[190]), .B(y[190]), .Z(n29229) );
  NANDN U25609 ( .A(x[189]), .B(y[189]), .Z(n10355) );
  AND U25610 ( .A(n29229), .B(n10355), .Z(n10738) );
  ANDN U25611 ( .B(x[188]), .A(y[188]), .Z(n29221) );
  NANDN U25612 ( .A(y[189]), .B(x[189]), .Z(n29227) );
  ANDN U25613 ( .B(x[187]), .A(y[187]), .Z(n29218) );
  ANDN U25614 ( .B(x[186]), .A(y[186]), .Z(n29213) );
  NOR U25615 ( .A(n29218), .B(n29213), .Z(n10732) );
  NANDN U25616 ( .A(x[186]), .B(y[186]), .Z(n28476) );
  ANDN U25617 ( .B(x[184]), .A(y[184]), .Z(n29204) );
  NANDN U25618 ( .A(x[183]), .B(y[183]), .Z(n29201) );
  ANDN U25619 ( .B(x[182]), .A(y[182]), .Z(n29199) );
  ANDN U25620 ( .B(x[181]), .A(y[181]), .Z(n29196) );
  ANDN U25621 ( .B(x[180]), .A(y[180]), .Z(n29191) );
  NOR U25622 ( .A(n29196), .B(n29191), .Z(n10720) );
  NANDN U25623 ( .A(x[180]), .B(y[180]), .Z(n28478) );
  ANDN U25624 ( .B(x[178]), .A(y[178]), .Z(n29182) );
  NANDN U25625 ( .A(x[177]), .B(y[177]), .Z(n29179) );
  ANDN U25626 ( .B(x[176]), .A(y[176]), .Z(n29177) );
  ANDN U25627 ( .B(x[175]), .A(y[175]), .Z(n29174) );
  ANDN U25628 ( .B(x[174]), .A(y[174]), .Z(n29169) );
  NOR U25629 ( .A(n29174), .B(n29169), .Z(n10708) );
  NANDN U25630 ( .A(x[174]), .B(y[174]), .Z(n28480) );
  NANDN U25631 ( .A(y[172]), .B(x[172]), .Z(n10704) );
  XOR U25632 ( .A(y[172]), .B(x[172]), .Z(n29163) );
  ANDN U25633 ( .B(x[170]), .A(y[170]), .Z(n29155) );
  ANDN U25634 ( .B(x[169]), .A(y[169]), .Z(n29152) );
  ANDN U25635 ( .B(x[168]), .A(y[168]), .Z(n29147) );
  NOR U25636 ( .A(n29152), .B(n29147), .Z(n10695) );
  NANDN U25637 ( .A(x[168]), .B(y[168]), .Z(n28482) );
  ANDN U25638 ( .B(x[166]), .A(y[166]), .Z(n29138) );
  NANDN U25639 ( .A(x[165]), .B(y[165]), .Z(n29135) );
  ANDN U25640 ( .B(x[164]), .A(y[164]), .Z(n29133) );
  ANDN U25641 ( .B(x[163]), .A(y[163]), .Z(n29130) );
  ANDN U25642 ( .B(x[162]), .A(y[162]), .Z(n29125) );
  NOR U25643 ( .A(n29130), .B(n29125), .Z(n10683) );
  NANDN U25644 ( .A(x[162]), .B(y[162]), .Z(n28484) );
  ANDN U25645 ( .B(x[160]), .A(y[160]), .Z(n29116) );
  NANDN U25646 ( .A(x[159]), .B(y[159]), .Z(n29113) );
  ANDN U25647 ( .B(x[158]), .A(y[158]), .Z(n29111) );
  ANDN U25648 ( .B(x[157]), .A(y[157]), .Z(n29108) );
  ANDN U25649 ( .B(x[156]), .A(y[156]), .Z(n29103) );
  NOR U25650 ( .A(n29108), .B(n29103), .Z(n10671) );
  NANDN U25651 ( .A(x[156]), .B(y[156]), .Z(n28486) );
  ANDN U25652 ( .B(x[154]), .A(y[154]), .Z(n29094) );
  NANDN U25653 ( .A(x[153]), .B(y[153]), .Z(n29091) );
  ANDN U25654 ( .B(x[152]), .A(y[152]), .Z(n29089) );
  ANDN U25655 ( .B(x[150]), .A(y[150]), .Z(n29083) );
  ANDN U25656 ( .B(x[151]), .A(y[151]), .Z(n29086) );
  NOR U25657 ( .A(n29083), .B(n29086), .Z(n10659) );
  NANDN U25658 ( .A(x[150]), .B(y[150]), .Z(n28488) );
  NANDN U25659 ( .A(y[149]), .B(x[149]), .Z(n10357) );
  NANDN U25660 ( .A(y[148]), .B(x[148]), .Z(n10356) );
  NAND U25661 ( .A(n10357), .B(n10356), .Z(n29079) );
  NANDN U25662 ( .A(x[147]), .B(y[147]), .Z(n29071) );
  ANDN U25663 ( .B(x[147]), .A(y[147]), .Z(n29075) );
  NANDN U25664 ( .A(x[145]), .B(y[145]), .Z(n29063) );
  ANDN U25665 ( .B(x[144]), .A(y[144]), .Z(n29061) );
  ANDN U25666 ( .B(x[143]), .A(y[143]), .Z(n29058) );
  ANDN U25667 ( .B(x[142]), .A(y[142]), .Z(n29053) );
  NOR U25668 ( .A(n29058), .B(n29053), .Z(n10644) );
  NANDN U25669 ( .A(x[142]), .B(y[142]), .Z(n28490) );
  ANDN U25670 ( .B(x[140]), .A(y[140]), .Z(n29044) );
  NANDN U25671 ( .A(x[139]), .B(y[139]), .Z(n29041) );
  ANDN U25672 ( .B(x[138]), .A(y[138]), .Z(n29039) );
  ANDN U25673 ( .B(x[137]), .A(y[137]), .Z(n29036) );
  ANDN U25674 ( .B(x[136]), .A(y[136]), .Z(n29031) );
  NOR U25675 ( .A(n29036), .B(n29031), .Z(n10632) );
  NANDN U25676 ( .A(x[136]), .B(y[136]), .Z(n28492) );
  ANDN U25677 ( .B(x[134]), .A(y[134]), .Z(n29022) );
  NANDN U25678 ( .A(x[133]), .B(y[133]), .Z(n29019) );
  ANDN U25679 ( .B(x[132]), .A(y[132]), .Z(n29017) );
  ANDN U25680 ( .B(x[131]), .A(y[131]), .Z(n29014) );
  ANDN U25681 ( .B(x[130]), .A(y[130]), .Z(n29009) );
  NOR U25682 ( .A(n29014), .B(n29009), .Z(n10620) );
  NANDN U25683 ( .A(x[130]), .B(y[130]), .Z(n28494) );
  ANDN U25684 ( .B(x[128]), .A(y[128]), .Z(n29000) );
  NANDN U25685 ( .A(x[127]), .B(y[127]), .Z(n28997) );
  ANDN U25686 ( .B(x[126]), .A(y[126]), .Z(n28995) );
  ANDN U25687 ( .B(x[125]), .A(y[125]), .Z(n28992) );
  ANDN U25688 ( .B(x[124]), .A(y[124]), .Z(n28987) );
  NOR U25689 ( .A(n28992), .B(n28987), .Z(n10608) );
  NANDN U25690 ( .A(x[124]), .B(y[124]), .Z(n28496) );
  ANDN U25691 ( .B(x[122]), .A(y[122]), .Z(n28978) );
  NANDN U25692 ( .A(x[121]), .B(y[121]), .Z(n28975) );
  ANDN U25693 ( .B(x[120]), .A(y[120]), .Z(n28973) );
  ANDN U25694 ( .B(x[119]), .A(y[119]), .Z(n28970) );
  ANDN U25695 ( .B(x[118]), .A(y[118]), .Z(n28965) );
  NOR U25696 ( .A(n28970), .B(n28965), .Z(n10596) );
  NANDN U25697 ( .A(x[118]), .B(y[118]), .Z(n28498) );
  ANDN U25698 ( .B(x[116]), .A(y[116]), .Z(n28956) );
  NANDN U25699 ( .A(x[115]), .B(y[115]), .Z(n28953) );
  ANDN U25700 ( .B(x[114]), .A(y[114]), .Z(n28951) );
  ANDN U25701 ( .B(x[113]), .A(y[113]), .Z(n28948) );
  ANDN U25702 ( .B(x[112]), .A(y[112]), .Z(n28943) );
  NOR U25703 ( .A(n28948), .B(n28943), .Z(n10584) );
  NANDN U25704 ( .A(x[112]), .B(y[112]), .Z(n28500) );
  ANDN U25705 ( .B(x[110]), .A(y[110]), .Z(n28934) );
  NANDN U25706 ( .A(x[109]), .B(y[109]), .Z(n28931) );
  ANDN U25707 ( .B(x[108]), .A(y[108]), .Z(n28929) );
  ANDN U25708 ( .B(x[107]), .A(y[107]), .Z(n28926) );
  ANDN U25709 ( .B(x[106]), .A(y[106]), .Z(n28921) );
  NOR U25710 ( .A(n28926), .B(n28921), .Z(n10572) );
  NANDN U25711 ( .A(x[106]), .B(y[106]), .Z(n28502) );
  ANDN U25712 ( .B(x[104]), .A(y[104]), .Z(n28912) );
  NANDN U25713 ( .A(x[103]), .B(y[103]), .Z(n28909) );
  ANDN U25714 ( .B(x[102]), .A(y[102]), .Z(n28907) );
  ANDN U25715 ( .B(x[101]), .A(y[101]), .Z(n28904) );
  ANDN U25716 ( .B(x[100]), .A(y[100]), .Z(n28899) );
  NOR U25717 ( .A(n28904), .B(n28899), .Z(n10560) );
  NANDN U25718 ( .A(x[100]), .B(y[100]), .Z(n28504) );
  ANDN U25719 ( .B(x[98]), .A(y[98]), .Z(n28890) );
  NANDN U25720 ( .A(x[97]), .B(y[97]), .Z(n28887) );
  ANDN U25721 ( .B(x[96]), .A(y[96]), .Z(n28885) );
  ANDN U25722 ( .B(x[95]), .A(y[95]), .Z(n28882) );
  ANDN U25723 ( .B(x[94]), .A(y[94]), .Z(n28877) );
  NOR U25724 ( .A(n28882), .B(n28877), .Z(n10548) );
  NANDN U25725 ( .A(x[94]), .B(y[94]), .Z(n28506) );
  ANDN U25726 ( .B(x[92]), .A(y[92]), .Z(n28868) );
  NANDN U25727 ( .A(x[91]), .B(y[91]), .Z(n28865) );
  ANDN U25728 ( .B(x[90]), .A(y[90]), .Z(n28863) );
  ANDN U25729 ( .B(x[89]), .A(y[89]), .Z(n28860) );
  ANDN U25730 ( .B(x[88]), .A(y[88]), .Z(n28855) );
  NOR U25731 ( .A(n28860), .B(n28855), .Z(n10536) );
  NANDN U25732 ( .A(x[88]), .B(y[88]), .Z(n28508) );
  ANDN U25733 ( .B(x[86]), .A(y[86]), .Z(n28846) );
  NANDN U25734 ( .A(x[85]), .B(y[85]), .Z(n28843) );
  ANDN U25735 ( .B(x[84]), .A(y[84]), .Z(n28841) );
  ANDN U25736 ( .B(x[83]), .A(y[83]), .Z(n28838) );
  ANDN U25737 ( .B(x[82]), .A(y[82]), .Z(n28833) );
  NOR U25738 ( .A(n28838), .B(n28833), .Z(n10524) );
  NANDN U25739 ( .A(x[82]), .B(y[82]), .Z(n28510) );
  ANDN U25740 ( .B(x[80]), .A(y[80]), .Z(n28824) );
  NANDN U25741 ( .A(x[79]), .B(y[79]), .Z(n28821) );
  ANDN U25742 ( .B(x[78]), .A(y[78]), .Z(n28819) );
  ANDN U25743 ( .B(x[77]), .A(y[77]), .Z(n28816) );
  ANDN U25744 ( .B(x[76]), .A(y[76]), .Z(n28811) );
  NOR U25745 ( .A(n28816), .B(n28811), .Z(n10512) );
  NANDN U25746 ( .A(x[76]), .B(y[76]), .Z(n28512) );
  ANDN U25747 ( .B(x[74]), .A(y[74]), .Z(n28802) );
  NANDN U25748 ( .A(x[73]), .B(y[73]), .Z(n28799) );
  ANDN U25749 ( .B(x[72]), .A(y[72]), .Z(n28797) );
  ANDN U25750 ( .B(x[71]), .A(y[71]), .Z(n28794) );
  ANDN U25751 ( .B(x[70]), .A(y[70]), .Z(n28789) );
  NOR U25752 ( .A(n28794), .B(n28789), .Z(n10500) );
  NANDN U25753 ( .A(x[70]), .B(y[70]), .Z(n28514) );
  ANDN U25754 ( .B(x[68]), .A(y[68]), .Z(n28780) );
  NANDN U25755 ( .A(x[67]), .B(y[67]), .Z(n28777) );
  ANDN U25756 ( .B(x[66]), .A(y[66]), .Z(n28775) );
  ANDN U25757 ( .B(x[65]), .A(y[65]), .Z(n28772) );
  ANDN U25758 ( .B(x[64]), .A(y[64]), .Z(n28767) );
  NOR U25759 ( .A(n28772), .B(n28767), .Z(n10488) );
  NANDN U25760 ( .A(x[64]), .B(y[64]), .Z(n28516) );
  ANDN U25761 ( .B(x[62]), .A(y[62]), .Z(n28758) );
  NANDN U25762 ( .A(x[61]), .B(y[61]), .Z(n28755) );
  ANDN U25763 ( .B(x[60]), .A(y[60]), .Z(n28753) );
  ANDN U25764 ( .B(x[59]), .A(y[59]), .Z(n28750) );
  ANDN U25765 ( .B(x[58]), .A(y[58]), .Z(n28745) );
  NOR U25766 ( .A(n28750), .B(n28745), .Z(n10476) );
  NANDN U25767 ( .A(x[58]), .B(y[58]), .Z(n28518) );
  ANDN U25768 ( .B(x[56]), .A(y[56]), .Z(n28736) );
  NANDN U25769 ( .A(x[55]), .B(y[55]), .Z(n28733) );
  ANDN U25770 ( .B(x[54]), .A(y[54]), .Z(n28731) );
  ANDN U25771 ( .B(x[53]), .A(y[53]), .Z(n28728) );
  ANDN U25772 ( .B(x[52]), .A(y[52]), .Z(n28723) );
  NOR U25773 ( .A(n28728), .B(n28723), .Z(n10464) );
  NANDN U25774 ( .A(x[52]), .B(y[52]), .Z(n28520) );
  ANDN U25775 ( .B(x[50]), .A(y[50]), .Z(n28714) );
  NANDN U25776 ( .A(x[49]), .B(y[49]), .Z(n28711) );
  ANDN U25777 ( .B(x[48]), .A(y[48]), .Z(n28709) );
  ANDN U25778 ( .B(x[47]), .A(y[47]), .Z(n28706) );
  ANDN U25779 ( .B(x[46]), .A(y[46]), .Z(n28701) );
  NOR U25780 ( .A(n28706), .B(n28701), .Z(n10452) );
  NANDN U25781 ( .A(x[46]), .B(y[46]), .Z(n28522) );
  ANDN U25782 ( .B(x[44]), .A(y[44]), .Z(n28692) );
  NANDN U25783 ( .A(x[43]), .B(y[43]), .Z(n28689) );
  ANDN U25784 ( .B(x[42]), .A(y[42]), .Z(n28687) );
  ANDN U25785 ( .B(x[40]), .A(y[40]), .Z(n28679) );
  ANDN U25786 ( .B(x[41]), .A(y[41]), .Z(n28684) );
  NOR U25787 ( .A(n28679), .B(n28684), .Z(n10440) );
  NANDN U25788 ( .A(x[38]), .B(y[38]), .Z(n10359) );
  NANDN U25789 ( .A(x[39]), .B(y[39]), .Z(n10358) );
  AND U25790 ( .A(n10359), .B(n10358), .Z(n28677) );
  ANDN U25791 ( .B(x[38]), .A(y[38]), .Z(n28674) );
  NANDN U25792 ( .A(x[37]), .B(y[37]), .Z(n28668) );
  ANDN U25793 ( .B(x[36]), .A(y[36]), .Z(n28664) );
  NANDN U25794 ( .A(x[35]), .B(y[35]), .Z(n28661) );
  ANDN U25795 ( .B(x[34]), .A(y[34]), .Z(n28659) );
  ANDN U25796 ( .B(x[33]), .A(y[33]), .Z(n28656) );
  ANDN U25797 ( .B(x[32]), .A(y[32]), .Z(n28651) );
  NOR U25798 ( .A(n28656), .B(n28651), .Z(n10425) );
  NANDN U25799 ( .A(x[32]), .B(y[32]), .Z(n28526) );
  ANDN U25800 ( .B(x[30]), .A(y[30]), .Z(n28642) );
  NANDN U25801 ( .A(x[29]), .B(y[29]), .Z(n28639) );
  ANDN U25802 ( .B(x[28]), .A(y[28]), .Z(n28637) );
  ANDN U25803 ( .B(x[27]), .A(y[27]), .Z(n28634) );
  ANDN U25804 ( .B(x[26]), .A(y[26]), .Z(n28629) );
  NOR U25805 ( .A(n28634), .B(n28629), .Z(n10413) );
  NANDN U25806 ( .A(x[26]), .B(y[26]), .Z(n28528) );
  ANDN U25807 ( .B(x[24]), .A(y[24]), .Z(n28620) );
  NANDN U25808 ( .A(x[23]), .B(y[23]), .Z(n28617) );
  ANDN U25809 ( .B(x[22]), .A(y[22]), .Z(n28615) );
  NANDN U25810 ( .A(y[20]), .B(x[20]), .Z(n10360) );
  ANDN U25811 ( .B(x[21]), .A(y[21]), .Z(n28612) );
  ANDN U25812 ( .B(n10360), .A(n28612), .Z(n10401) );
  XOR U25813 ( .A(y[20]), .B(x[20]), .Z(n28607) );
  ANDN U25814 ( .B(x[19]), .A(y[19]), .Z(n28608) );
  NANDN U25815 ( .A(x[17]), .B(y[17]), .Z(n28595) );
  ANDN U25816 ( .B(x[16]), .A(y[16]), .Z(n28593) );
  ANDN U25817 ( .B(x[15]), .A(y[15]), .Z(n28590) );
  ANDN U25818 ( .B(x[14]), .A(y[14]), .Z(n28585) );
  NOR U25819 ( .A(n28590), .B(n28585), .Z(n10389) );
  NANDN U25820 ( .A(x[14]), .B(y[14]), .Z(n28532) );
  ANDN U25821 ( .B(x[12]), .A(y[12]), .Z(n28576) );
  NANDN U25822 ( .A(x[11]), .B(y[11]), .Z(n28573) );
  ANDN U25823 ( .B(x[10]), .A(y[10]), .Z(n28571) );
  ANDN U25824 ( .B(x[9]), .A(y[9]), .Z(n28568) );
  ANDN U25825 ( .B(x[8]), .A(y[8]), .Z(n28563) );
  NOR U25826 ( .A(n28568), .B(n28563), .Z(n10377) );
  NANDN U25827 ( .A(x[8]), .B(y[8]), .Z(n28534) );
  ANDN U25828 ( .B(x[6]), .A(y[6]), .Z(n28554) );
  NANDN U25829 ( .A(x[5]), .B(y[5]), .Z(n28551) );
  ANDN U25830 ( .B(x[4]), .A(y[4]), .Z(n28549) );
  ANDN U25831 ( .B(x[3]), .A(y[3]), .Z(n28546) );
  ANDN U25832 ( .B(x[2]), .A(y[2]), .Z(n28541) );
  NOR U25833 ( .A(n28546), .B(n28541), .Z(n10365) );
  NANDN U25834 ( .A(x[2]), .B(y[2]), .Z(n28536) );
  ANDN U25835 ( .B(x[1]), .A(y[1]), .Z(n28542) );
  NANDN U25836 ( .A(y[0]), .B(x[0]), .Z(n10361) );
  NANDN U25837 ( .A(n28542), .B(n10361), .Z(n10362) );
  NAND U25838 ( .A(n28536), .B(n10362), .Z(n10363) );
  NANDN U25839 ( .A(x[1]), .B(y[1]), .Z(n28539) );
  NANDN U25840 ( .A(n10363), .B(n28539), .Z(n10364) );
  AND U25841 ( .A(n10365), .B(n10364), .Z(n10367) );
  NANDN U25842 ( .A(x[3]), .B(y[3]), .Z(n28537) );
  NANDN U25843 ( .A(x[4]), .B(y[4]), .Z(n28552) );
  AND U25844 ( .A(n28537), .B(n28552), .Z(n10366) );
  NANDN U25845 ( .A(n10367), .B(n10366), .Z(n10368) );
  ANDN U25846 ( .B(x[5]), .A(y[5]), .Z(n28557) );
  ANDN U25847 ( .B(n10368), .A(n28557), .Z(n10369) );
  NANDN U25848 ( .A(n28549), .B(n10369), .Z(n10370) );
  NANDN U25849 ( .A(x[6]), .B(y[6]), .Z(n28558) );
  AND U25850 ( .A(n10370), .B(n28558), .Z(n10371) );
  NAND U25851 ( .A(n28551), .B(n10371), .Z(n10372) );
  ANDN U25852 ( .B(x[7]), .A(y[7]), .Z(n28564) );
  ANDN U25853 ( .B(n10372), .A(n28564), .Z(n10373) );
  NANDN U25854 ( .A(n28554), .B(n10373), .Z(n10374) );
  NAND U25855 ( .A(n28534), .B(n10374), .Z(n10375) );
  NANDN U25856 ( .A(x[7]), .B(y[7]), .Z(n28559) );
  NANDN U25857 ( .A(n10375), .B(n28559), .Z(n10376) );
  AND U25858 ( .A(n10377), .B(n10376), .Z(n10379) );
  NANDN U25859 ( .A(x[9]), .B(y[9]), .Z(n28535) );
  NANDN U25860 ( .A(x[10]), .B(y[10]), .Z(n28574) );
  AND U25861 ( .A(n28535), .B(n28574), .Z(n10378) );
  NANDN U25862 ( .A(n10379), .B(n10378), .Z(n10380) );
  ANDN U25863 ( .B(x[11]), .A(y[11]), .Z(n28579) );
  ANDN U25864 ( .B(n10380), .A(n28579), .Z(n10381) );
  NANDN U25865 ( .A(n28571), .B(n10381), .Z(n10382) );
  NANDN U25866 ( .A(x[12]), .B(y[12]), .Z(n28580) );
  AND U25867 ( .A(n10382), .B(n28580), .Z(n10383) );
  NAND U25868 ( .A(n28573), .B(n10383), .Z(n10384) );
  ANDN U25869 ( .B(x[13]), .A(y[13]), .Z(n28586) );
  ANDN U25870 ( .B(n10384), .A(n28586), .Z(n10385) );
  NANDN U25871 ( .A(n28576), .B(n10385), .Z(n10386) );
  NAND U25872 ( .A(n28532), .B(n10386), .Z(n10387) );
  NANDN U25873 ( .A(x[13]), .B(y[13]), .Z(n28581) );
  NANDN U25874 ( .A(n10387), .B(n28581), .Z(n10388) );
  AND U25875 ( .A(n10389), .B(n10388), .Z(n10391) );
  NANDN U25876 ( .A(x[15]), .B(y[15]), .Z(n28533) );
  NANDN U25877 ( .A(x[16]), .B(y[16]), .Z(n28596) );
  AND U25878 ( .A(n28533), .B(n28596), .Z(n10390) );
  NANDN U25879 ( .A(n10391), .B(n10390), .Z(n10392) );
  ANDN U25880 ( .B(x[17]), .A(y[17]), .Z(n28601) );
  ANDN U25881 ( .B(n10392), .A(n28601), .Z(n10393) );
  NANDN U25882 ( .A(n28593), .B(n10393), .Z(n10394) );
  NANDN U25883 ( .A(x[18]), .B(y[18]), .Z(n28605) );
  AND U25884 ( .A(n10394), .B(n28605), .Z(n10395) );
  NAND U25885 ( .A(n28595), .B(n10395), .Z(n10396) );
  ANDN U25886 ( .B(x[18]), .A(y[18]), .Z(n28598) );
  ANDN U25887 ( .B(n10396), .A(n28598), .Z(n10397) );
  NANDN U25888 ( .A(n28608), .B(n10397), .Z(n10398) );
  NANDN U25889 ( .A(n28607), .B(n10398), .Z(n10399) );
  NANDN U25890 ( .A(x[19]), .B(y[19]), .Z(n28603) );
  NANDN U25891 ( .A(n10399), .B(n28603), .Z(n10400) );
  AND U25892 ( .A(n10401), .B(n10400), .Z(n10403) );
  NANDN U25893 ( .A(x[21]), .B(y[21]), .Z(n28530) );
  NANDN U25894 ( .A(x[22]), .B(y[22]), .Z(n28618) );
  AND U25895 ( .A(n28530), .B(n28618), .Z(n10402) );
  NANDN U25896 ( .A(n10403), .B(n10402), .Z(n10404) );
  ANDN U25897 ( .B(x[23]), .A(y[23]), .Z(n28623) );
  ANDN U25898 ( .B(n10404), .A(n28623), .Z(n10405) );
  NANDN U25899 ( .A(n28615), .B(n10405), .Z(n10406) );
  NANDN U25900 ( .A(x[24]), .B(y[24]), .Z(n28624) );
  AND U25901 ( .A(n10406), .B(n28624), .Z(n10407) );
  NAND U25902 ( .A(n28617), .B(n10407), .Z(n10408) );
  ANDN U25903 ( .B(x[25]), .A(y[25]), .Z(n28630) );
  ANDN U25904 ( .B(n10408), .A(n28630), .Z(n10409) );
  NANDN U25905 ( .A(n28620), .B(n10409), .Z(n10410) );
  NAND U25906 ( .A(n28528), .B(n10410), .Z(n10411) );
  NANDN U25907 ( .A(x[25]), .B(y[25]), .Z(n28625) );
  NANDN U25908 ( .A(n10411), .B(n28625), .Z(n10412) );
  AND U25909 ( .A(n10413), .B(n10412), .Z(n10415) );
  NANDN U25910 ( .A(x[27]), .B(y[27]), .Z(n28529) );
  NANDN U25911 ( .A(x[28]), .B(y[28]), .Z(n28640) );
  AND U25912 ( .A(n28529), .B(n28640), .Z(n10414) );
  NANDN U25913 ( .A(n10415), .B(n10414), .Z(n10416) );
  ANDN U25914 ( .B(x[29]), .A(y[29]), .Z(n28645) );
  ANDN U25915 ( .B(n10416), .A(n28645), .Z(n10417) );
  NANDN U25916 ( .A(n28637), .B(n10417), .Z(n10418) );
  NANDN U25917 ( .A(x[30]), .B(y[30]), .Z(n28646) );
  AND U25918 ( .A(n10418), .B(n28646), .Z(n10419) );
  NAND U25919 ( .A(n28639), .B(n10419), .Z(n10420) );
  ANDN U25920 ( .B(x[31]), .A(y[31]), .Z(n28652) );
  ANDN U25921 ( .B(n10420), .A(n28652), .Z(n10421) );
  NANDN U25922 ( .A(n28642), .B(n10421), .Z(n10422) );
  NAND U25923 ( .A(n28526), .B(n10422), .Z(n10423) );
  NANDN U25924 ( .A(x[31]), .B(y[31]), .Z(n28647) );
  NANDN U25925 ( .A(n10423), .B(n28647), .Z(n10424) );
  AND U25926 ( .A(n10425), .B(n10424), .Z(n10427) );
  NANDN U25927 ( .A(x[33]), .B(y[33]), .Z(n28527) );
  NANDN U25928 ( .A(x[34]), .B(y[34]), .Z(n28662) );
  AND U25929 ( .A(n28527), .B(n28662), .Z(n10426) );
  NANDN U25930 ( .A(n10427), .B(n10426), .Z(n10428) );
  ANDN U25931 ( .B(x[35]), .A(y[35]), .Z(n28667) );
  ANDN U25932 ( .B(n10428), .A(n28667), .Z(n10429) );
  NANDN U25933 ( .A(n28659), .B(n10429), .Z(n10430) );
  NANDN U25934 ( .A(x[36]), .B(y[36]), .Z(n28669) );
  AND U25935 ( .A(n10430), .B(n28669), .Z(n10431) );
  NAND U25936 ( .A(n28661), .B(n10431), .Z(n10432) );
  ANDN U25937 ( .B(x[37]), .A(y[37]), .Z(n28673) );
  ANDN U25938 ( .B(n10432), .A(n28673), .Z(n10433) );
  NANDN U25939 ( .A(n28664), .B(n10433), .Z(n10434) );
  NAND U25940 ( .A(n28668), .B(n10434), .Z(n10435) );
  NANDN U25941 ( .A(n28674), .B(n10435), .Z(n10436) );
  NAND U25942 ( .A(n28677), .B(n10436), .Z(n10437) );
  ANDN U25943 ( .B(x[39]), .A(y[39]), .Z(n28680) );
  ANDN U25944 ( .B(n10437), .A(n28680), .Z(n10438) );
  NANDN U25945 ( .A(x[40]), .B(y[40]), .Z(n28524) );
  NANDN U25946 ( .A(n10438), .B(n28524), .Z(n10439) );
  AND U25947 ( .A(n10440), .B(n10439), .Z(n10442) );
  NANDN U25948 ( .A(x[41]), .B(y[41]), .Z(n28525) );
  NANDN U25949 ( .A(x[42]), .B(y[42]), .Z(n28690) );
  AND U25950 ( .A(n28525), .B(n28690), .Z(n10441) );
  NANDN U25951 ( .A(n10442), .B(n10441), .Z(n10443) );
  ANDN U25952 ( .B(x[43]), .A(y[43]), .Z(n28695) );
  ANDN U25953 ( .B(n10443), .A(n28695), .Z(n10444) );
  NANDN U25954 ( .A(n28687), .B(n10444), .Z(n10445) );
  NANDN U25955 ( .A(x[44]), .B(y[44]), .Z(n28696) );
  AND U25956 ( .A(n10445), .B(n28696), .Z(n10446) );
  NAND U25957 ( .A(n28689), .B(n10446), .Z(n10447) );
  ANDN U25958 ( .B(x[45]), .A(y[45]), .Z(n28702) );
  ANDN U25959 ( .B(n10447), .A(n28702), .Z(n10448) );
  NANDN U25960 ( .A(n28692), .B(n10448), .Z(n10449) );
  NAND U25961 ( .A(n28522), .B(n10449), .Z(n10450) );
  NANDN U25962 ( .A(x[45]), .B(y[45]), .Z(n28697) );
  NANDN U25963 ( .A(n10450), .B(n28697), .Z(n10451) );
  AND U25964 ( .A(n10452), .B(n10451), .Z(n10454) );
  NANDN U25965 ( .A(x[47]), .B(y[47]), .Z(n28523) );
  NANDN U25966 ( .A(x[48]), .B(y[48]), .Z(n28712) );
  AND U25967 ( .A(n28523), .B(n28712), .Z(n10453) );
  NANDN U25968 ( .A(n10454), .B(n10453), .Z(n10455) );
  ANDN U25969 ( .B(x[49]), .A(y[49]), .Z(n28717) );
  ANDN U25970 ( .B(n10455), .A(n28717), .Z(n10456) );
  NANDN U25971 ( .A(n28709), .B(n10456), .Z(n10457) );
  NANDN U25972 ( .A(x[50]), .B(y[50]), .Z(n28718) );
  AND U25973 ( .A(n10457), .B(n28718), .Z(n10458) );
  NAND U25974 ( .A(n28711), .B(n10458), .Z(n10459) );
  ANDN U25975 ( .B(x[51]), .A(y[51]), .Z(n28724) );
  ANDN U25976 ( .B(n10459), .A(n28724), .Z(n10460) );
  NANDN U25977 ( .A(n28714), .B(n10460), .Z(n10461) );
  NAND U25978 ( .A(n28520), .B(n10461), .Z(n10462) );
  NANDN U25979 ( .A(x[51]), .B(y[51]), .Z(n28719) );
  NANDN U25980 ( .A(n10462), .B(n28719), .Z(n10463) );
  AND U25981 ( .A(n10464), .B(n10463), .Z(n10466) );
  NANDN U25982 ( .A(x[53]), .B(y[53]), .Z(n28521) );
  NANDN U25983 ( .A(x[54]), .B(y[54]), .Z(n28734) );
  AND U25984 ( .A(n28521), .B(n28734), .Z(n10465) );
  NANDN U25985 ( .A(n10466), .B(n10465), .Z(n10467) );
  ANDN U25986 ( .B(x[55]), .A(y[55]), .Z(n28739) );
  ANDN U25987 ( .B(n10467), .A(n28739), .Z(n10468) );
  NANDN U25988 ( .A(n28731), .B(n10468), .Z(n10469) );
  NANDN U25989 ( .A(x[56]), .B(y[56]), .Z(n28740) );
  AND U25990 ( .A(n10469), .B(n28740), .Z(n10470) );
  NAND U25991 ( .A(n28733), .B(n10470), .Z(n10471) );
  ANDN U25992 ( .B(x[57]), .A(y[57]), .Z(n28746) );
  ANDN U25993 ( .B(n10471), .A(n28746), .Z(n10472) );
  NANDN U25994 ( .A(n28736), .B(n10472), .Z(n10473) );
  NAND U25995 ( .A(n28518), .B(n10473), .Z(n10474) );
  NANDN U25996 ( .A(x[57]), .B(y[57]), .Z(n28741) );
  NANDN U25997 ( .A(n10474), .B(n28741), .Z(n10475) );
  AND U25998 ( .A(n10476), .B(n10475), .Z(n10478) );
  NANDN U25999 ( .A(x[59]), .B(y[59]), .Z(n28519) );
  NANDN U26000 ( .A(x[60]), .B(y[60]), .Z(n28756) );
  AND U26001 ( .A(n28519), .B(n28756), .Z(n10477) );
  NANDN U26002 ( .A(n10478), .B(n10477), .Z(n10479) );
  ANDN U26003 ( .B(x[61]), .A(y[61]), .Z(n28761) );
  ANDN U26004 ( .B(n10479), .A(n28761), .Z(n10480) );
  NANDN U26005 ( .A(n28753), .B(n10480), .Z(n10481) );
  NANDN U26006 ( .A(x[62]), .B(y[62]), .Z(n28762) );
  AND U26007 ( .A(n10481), .B(n28762), .Z(n10482) );
  NAND U26008 ( .A(n28755), .B(n10482), .Z(n10483) );
  ANDN U26009 ( .B(x[63]), .A(y[63]), .Z(n28768) );
  ANDN U26010 ( .B(n10483), .A(n28768), .Z(n10484) );
  NANDN U26011 ( .A(n28758), .B(n10484), .Z(n10485) );
  NAND U26012 ( .A(n28516), .B(n10485), .Z(n10486) );
  NANDN U26013 ( .A(x[63]), .B(y[63]), .Z(n28763) );
  NANDN U26014 ( .A(n10486), .B(n28763), .Z(n10487) );
  AND U26015 ( .A(n10488), .B(n10487), .Z(n10490) );
  NANDN U26016 ( .A(x[65]), .B(y[65]), .Z(n28517) );
  NANDN U26017 ( .A(x[66]), .B(y[66]), .Z(n28778) );
  AND U26018 ( .A(n28517), .B(n28778), .Z(n10489) );
  NANDN U26019 ( .A(n10490), .B(n10489), .Z(n10491) );
  ANDN U26020 ( .B(x[67]), .A(y[67]), .Z(n28783) );
  ANDN U26021 ( .B(n10491), .A(n28783), .Z(n10492) );
  NANDN U26022 ( .A(n28775), .B(n10492), .Z(n10493) );
  NANDN U26023 ( .A(x[68]), .B(y[68]), .Z(n28784) );
  AND U26024 ( .A(n10493), .B(n28784), .Z(n10494) );
  NAND U26025 ( .A(n28777), .B(n10494), .Z(n10495) );
  ANDN U26026 ( .B(x[69]), .A(y[69]), .Z(n28790) );
  ANDN U26027 ( .B(n10495), .A(n28790), .Z(n10496) );
  NANDN U26028 ( .A(n28780), .B(n10496), .Z(n10497) );
  NAND U26029 ( .A(n28514), .B(n10497), .Z(n10498) );
  NANDN U26030 ( .A(x[69]), .B(y[69]), .Z(n28785) );
  NANDN U26031 ( .A(n10498), .B(n28785), .Z(n10499) );
  AND U26032 ( .A(n10500), .B(n10499), .Z(n10502) );
  NANDN U26033 ( .A(x[71]), .B(y[71]), .Z(n28515) );
  NANDN U26034 ( .A(x[72]), .B(y[72]), .Z(n28800) );
  AND U26035 ( .A(n28515), .B(n28800), .Z(n10501) );
  NANDN U26036 ( .A(n10502), .B(n10501), .Z(n10503) );
  ANDN U26037 ( .B(x[73]), .A(y[73]), .Z(n28805) );
  ANDN U26038 ( .B(n10503), .A(n28805), .Z(n10504) );
  NANDN U26039 ( .A(n28797), .B(n10504), .Z(n10505) );
  NANDN U26040 ( .A(x[74]), .B(y[74]), .Z(n28806) );
  AND U26041 ( .A(n10505), .B(n28806), .Z(n10506) );
  NAND U26042 ( .A(n28799), .B(n10506), .Z(n10507) );
  ANDN U26043 ( .B(x[75]), .A(y[75]), .Z(n28812) );
  ANDN U26044 ( .B(n10507), .A(n28812), .Z(n10508) );
  NANDN U26045 ( .A(n28802), .B(n10508), .Z(n10509) );
  NAND U26046 ( .A(n28512), .B(n10509), .Z(n10510) );
  NANDN U26047 ( .A(x[75]), .B(y[75]), .Z(n28807) );
  NANDN U26048 ( .A(n10510), .B(n28807), .Z(n10511) );
  AND U26049 ( .A(n10512), .B(n10511), .Z(n10514) );
  NANDN U26050 ( .A(x[77]), .B(y[77]), .Z(n28513) );
  NANDN U26051 ( .A(x[78]), .B(y[78]), .Z(n28822) );
  AND U26052 ( .A(n28513), .B(n28822), .Z(n10513) );
  NANDN U26053 ( .A(n10514), .B(n10513), .Z(n10515) );
  ANDN U26054 ( .B(x[79]), .A(y[79]), .Z(n28827) );
  ANDN U26055 ( .B(n10515), .A(n28827), .Z(n10516) );
  NANDN U26056 ( .A(n28819), .B(n10516), .Z(n10517) );
  NANDN U26057 ( .A(x[80]), .B(y[80]), .Z(n28828) );
  AND U26058 ( .A(n10517), .B(n28828), .Z(n10518) );
  NAND U26059 ( .A(n28821), .B(n10518), .Z(n10519) );
  ANDN U26060 ( .B(x[81]), .A(y[81]), .Z(n28834) );
  ANDN U26061 ( .B(n10519), .A(n28834), .Z(n10520) );
  NANDN U26062 ( .A(n28824), .B(n10520), .Z(n10521) );
  NAND U26063 ( .A(n28510), .B(n10521), .Z(n10522) );
  NANDN U26064 ( .A(x[81]), .B(y[81]), .Z(n28829) );
  NANDN U26065 ( .A(n10522), .B(n28829), .Z(n10523) );
  AND U26066 ( .A(n10524), .B(n10523), .Z(n10526) );
  NANDN U26067 ( .A(x[83]), .B(y[83]), .Z(n28511) );
  NANDN U26068 ( .A(x[84]), .B(y[84]), .Z(n28844) );
  AND U26069 ( .A(n28511), .B(n28844), .Z(n10525) );
  NANDN U26070 ( .A(n10526), .B(n10525), .Z(n10527) );
  ANDN U26071 ( .B(x[85]), .A(y[85]), .Z(n28849) );
  ANDN U26072 ( .B(n10527), .A(n28849), .Z(n10528) );
  NANDN U26073 ( .A(n28841), .B(n10528), .Z(n10529) );
  NANDN U26074 ( .A(x[86]), .B(y[86]), .Z(n28850) );
  AND U26075 ( .A(n10529), .B(n28850), .Z(n10530) );
  NAND U26076 ( .A(n28843), .B(n10530), .Z(n10531) );
  ANDN U26077 ( .B(x[87]), .A(y[87]), .Z(n28856) );
  ANDN U26078 ( .B(n10531), .A(n28856), .Z(n10532) );
  NANDN U26079 ( .A(n28846), .B(n10532), .Z(n10533) );
  NAND U26080 ( .A(n28508), .B(n10533), .Z(n10534) );
  NANDN U26081 ( .A(x[87]), .B(y[87]), .Z(n28851) );
  NANDN U26082 ( .A(n10534), .B(n28851), .Z(n10535) );
  AND U26083 ( .A(n10536), .B(n10535), .Z(n10538) );
  NANDN U26084 ( .A(x[89]), .B(y[89]), .Z(n28509) );
  NANDN U26085 ( .A(x[90]), .B(y[90]), .Z(n28866) );
  AND U26086 ( .A(n28509), .B(n28866), .Z(n10537) );
  NANDN U26087 ( .A(n10538), .B(n10537), .Z(n10539) );
  ANDN U26088 ( .B(x[91]), .A(y[91]), .Z(n28871) );
  ANDN U26089 ( .B(n10539), .A(n28871), .Z(n10540) );
  NANDN U26090 ( .A(n28863), .B(n10540), .Z(n10541) );
  NANDN U26091 ( .A(x[92]), .B(y[92]), .Z(n28872) );
  AND U26092 ( .A(n10541), .B(n28872), .Z(n10542) );
  NAND U26093 ( .A(n28865), .B(n10542), .Z(n10543) );
  ANDN U26094 ( .B(x[93]), .A(y[93]), .Z(n28878) );
  ANDN U26095 ( .B(n10543), .A(n28878), .Z(n10544) );
  NANDN U26096 ( .A(n28868), .B(n10544), .Z(n10545) );
  NAND U26097 ( .A(n28506), .B(n10545), .Z(n10546) );
  NANDN U26098 ( .A(x[93]), .B(y[93]), .Z(n28873) );
  NANDN U26099 ( .A(n10546), .B(n28873), .Z(n10547) );
  AND U26100 ( .A(n10548), .B(n10547), .Z(n10550) );
  NANDN U26101 ( .A(x[95]), .B(y[95]), .Z(n28507) );
  NANDN U26102 ( .A(x[96]), .B(y[96]), .Z(n28888) );
  AND U26103 ( .A(n28507), .B(n28888), .Z(n10549) );
  NANDN U26104 ( .A(n10550), .B(n10549), .Z(n10551) );
  ANDN U26105 ( .B(x[97]), .A(y[97]), .Z(n28893) );
  ANDN U26106 ( .B(n10551), .A(n28893), .Z(n10552) );
  NANDN U26107 ( .A(n28885), .B(n10552), .Z(n10553) );
  NANDN U26108 ( .A(x[98]), .B(y[98]), .Z(n28894) );
  AND U26109 ( .A(n10553), .B(n28894), .Z(n10554) );
  NAND U26110 ( .A(n28887), .B(n10554), .Z(n10555) );
  ANDN U26111 ( .B(x[99]), .A(y[99]), .Z(n28900) );
  ANDN U26112 ( .B(n10555), .A(n28900), .Z(n10556) );
  NANDN U26113 ( .A(n28890), .B(n10556), .Z(n10557) );
  NAND U26114 ( .A(n28504), .B(n10557), .Z(n10558) );
  NANDN U26115 ( .A(x[99]), .B(y[99]), .Z(n28895) );
  NANDN U26116 ( .A(n10558), .B(n28895), .Z(n10559) );
  AND U26117 ( .A(n10560), .B(n10559), .Z(n10562) );
  NANDN U26118 ( .A(x[101]), .B(y[101]), .Z(n28505) );
  NANDN U26119 ( .A(x[102]), .B(y[102]), .Z(n28910) );
  AND U26120 ( .A(n28505), .B(n28910), .Z(n10561) );
  NANDN U26121 ( .A(n10562), .B(n10561), .Z(n10563) );
  ANDN U26122 ( .B(x[103]), .A(y[103]), .Z(n28915) );
  ANDN U26123 ( .B(n10563), .A(n28915), .Z(n10564) );
  NANDN U26124 ( .A(n28907), .B(n10564), .Z(n10565) );
  NANDN U26125 ( .A(x[104]), .B(y[104]), .Z(n28916) );
  AND U26126 ( .A(n10565), .B(n28916), .Z(n10566) );
  NAND U26127 ( .A(n28909), .B(n10566), .Z(n10567) );
  ANDN U26128 ( .B(x[105]), .A(y[105]), .Z(n28922) );
  ANDN U26129 ( .B(n10567), .A(n28922), .Z(n10568) );
  NANDN U26130 ( .A(n28912), .B(n10568), .Z(n10569) );
  NAND U26131 ( .A(n28502), .B(n10569), .Z(n10570) );
  NANDN U26132 ( .A(x[105]), .B(y[105]), .Z(n28917) );
  NANDN U26133 ( .A(n10570), .B(n28917), .Z(n10571) );
  AND U26134 ( .A(n10572), .B(n10571), .Z(n10574) );
  NANDN U26135 ( .A(x[107]), .B(y[107]), .Z(n28503) );
  NANDN U26136 ( .A(x[108]), .B(y[108]), .Z(n28932) );
  AND U26137 ( .A(n28503), .B(n28932), .Z(n10573) );
  NANDN U26138 ( .A(n10574), .B(n10573), .Z(n10575) );
  ANDN U26139 ( .B(x[109]), .A(y[109]), .Z(n28937) );
  ANDN U26140 ( .B(n10575), .A(n28937), .Z(n10576) );
  NANDN U26141 ( .A(n28929), .B(n10576), .Z(n10577) );
  NANDN U26142 ( .A(x[110]), .B(y[110]), .Z(n28938) );
  AND U26143 ( .A(n10577), .B(n28938), .Z(n10578) );
  NAND U26144 ( .A(n28931), .B(n10578), .Z(n10579) );
  ANDN U26145 ( .B(x[111]), .A(y[111]), .Z(n28944) );
  ANDN U26146 ( .B(n10579), .A(n28944), .Z(n10580) );
  NANDN U26147 ( .A(n28934), .B(n10580), .Z(n10581) );
  NAND U26148 ( .A(n28500), .B(n10581), .Z(n10582) );
  NANDN U26149 ( .A(x[111]), .B(y[111]), .Z(n28939) );
  NANDN U26150 ( .A(n10582), .B(n28939), .Z(n10583) );
  AND U26151 ( .A(n10584), .B(n10583), .Z(n10586) );
  NANDN U26152 ( .A(x[113]), .B(y[113]), .Z(n28501) );
  NANDN U26153 ( .A(x[114]), .B(y[114]), .Z(n28954) );
  AND U26154 ( .A(n28501), .B(n28954), .Z(n10585) );
  NANDN U26155 ( .A(n10586), .B(n10585), .Z(n10587) );
  ANDN U26156 ( .B(x[115]), .A(y[115]), .Z(n28959) );
  ANDN U26157 ( .B(n10587), .A(n28959), .Z(n10588) );
  NANDN U26158 ( .A(n28951), .B(n10588), .Z(n10589) );
  NANDN U26159 ( .A(x[116]), .B(y[116]), .Z(n28960) );
  AND U26160 ( .A(n10589), .B(n28960), .Z(n10590) );
  NAND U26161 ( .A(n28953), .B(n10590), .Z(n10591) );
  ANDN U26162 ( .B(x[117]), .A(y[117]), .Z(n28966) );
  ANDN U26163 ( .B(n10591), .A(n28966), .Z(n10592) );
  NANDN U26164 ( .A(n28956), .B(n10592), .Z(n10593) );
  NAND U26165 ( .A(n28498), .B(n10593), .Z(n10594) );
  NANDN U26166 ( .A(x[117]), .B(y[117]), .Z(n28961) );
  NANDN U26167 ( .A(n10594), .B(n28961), .Z(n10595) );
  AND U26168 ( .A(n10596), .B(n10595), .Z(n10598) );
  NANDN U26169 ( .A(x[119]), .B(y[119]), .Z(n28499) );
  NANDN U26170 ( .A(x[120]), .B(y[120]), .Z(n28976) );
  AND U26171 ( .A(n28499), .B(n28976), .Z(n10597) );
  NANDN U26172 ( .A(n10598), .B(n10597), .Z(n10599) );
  ANDN U26173 ( .B(x[121]), .A(y[121]), .Z(n28981) );
  ANDN U26174 ( .B(n10599), .A(n28981), .Z(n10600) );
  NANDN U26175 ( .A(n28973), .B(n10600), .Z(n10601) );
  NANDN U26176 ( .A(x[122]), .B(y[122]), .Z(n28982) );
  AND U26177 ( .A(n10601), .B(n28982), .Z(n10602) );
  NAND U26178 ( .A(n28975), .B(n10602), .Z(n10603) );
  ANDN U26179 ( .B(x[123]), .A(y[123]), .Z(n28988) );
  ANDN U26180 ( .B(n10603), .A(n28988), .Z(n10604) );
  NANDN U26181 ( .A(n28978), .B(n10604), .Z(n10605) );
  NAND U26182 ( .A(n28496), .B(n10605), .Z(n10606) );
  NANDN U26183 ( .A(x[123]), .B(y[123]), .Z(n28983) );
  NANDN U26184 ( .A(n10606), .B(n28983), .Z(n10607) );
  AND U26185 ( .A(n10608), .B(n10607), .Z(n10610) );
  NANDN U26186 ( .A(x[125]), .B(y[125]), .Z(n28497) );
  NANDN U26187 ( .A(x[126]), .B(y[126]), .Z(n28998) );
  AND U26188 ( .A(n28497), .B(n28998), .Z(n10609) );
  NANDN U26189 ( .A(n10610), .B(n10609), .Z(n10611) );
  ANDN U26190 ( .B(x[127]), .A(y[127]), .Z(n29003) );
  ANDN U26191 ( .B(n10611), .A(n29003), .Z(n10612) );
  NANDN U26192 ( .A(n28995), .B(n10612), .Z(n10613) );
  NANDN U26193 ( .A(x[128]), .B(y[128]), .Z(n29004) );
  AND U26194 ( .A(n10613), .B(n29004), .Z(n10614) );
  NAND U26195 ( .A(n28997), .B(n10614), .Z(n10615) );
  ANDN U26196 ( .B(x[129]), .A(y[129]), .Z(n29010) );
  ANDN U26197 ( .B(n10615), .A(n29010), .Z(n10616) );
  NANDN U26198 ( .A(n29000), .B(n10616), .Z(n10617) );
  NAND U26199 ( .A(n28494), .B(n10617), .Z(n10618) );
  NANDN U26200 ( .A(x[129]), .B(y[129]), .Z(n29005) );
  NANDN U26201 ( .A(n10618), .B(n29005), .Z(n10619) );
  AND U26202 ( .A(n10620), .B(n10619), .Z(n10622) );
  NANDN U26203 ( .A(x[131]), .B(y[131]), .Z(n28495) );
  NANDN U26204 ( .A(x[132]), .B(y[132]), .Z(n29020) );
  AND U26205 ( .A(n28495), .B(n29020), .Z(n10621) );
  NANDN U26206 ( .A(n10622), .B(n10621), .Z(n10623) );
  ANDN U26207 ( .B(x[133]), .A(y[133]), .Z(n29025) );
  ANDN U26208 ( .B(n10623), .A(n29025), .Z(n10624) );
  NANDN U26209 ( .A(n29017), .B(n10624), .Z(n10625) );
  NANDN U26210 ( .A(x[134]), .B(y[134]), .Z(n29026) );
  AND U26211 ( .A(n10625), .B(n29026), .Z(n10626) );
  NAND U26212 ( .A(n29019), .B(n10626), .Z(n10627) );
  ANDN U26213 ( .B(x[135]), .A(y[135]), .Z(n29032) );
  ANDN U26214 ( .B(n10627), .A(n29032), .Z(n10628) );
  NANDN U26215 ( .A(n29022), .B(n10628), .Z(n10629) );
  NAND U26216 ( .A(n28492), .B(n10629), .Z(n10630) );
  NANDN U26217 ( .A(x[135]), .B(y[135]), .Z(n29027) );
  NANDN U26218 ( .A(n10630), .B(n29027), .Z(n10631) );
  AND U26219 ( .A(n10632), .B(n10631), .Z(n10634) );
  NANDN U26220 ( .A(x[137]), .B(y[137]), .Z(n28493) );
  NANDN U26221 ( .A(x[138]), .B(y[138]), .Z(n29042) );
  AND U26222 ( .A(n28493), .B(n29042), .Z(n10633) );
  NANDN U26223 ( .A(n10634), .B(n10633), .Z(n10635) );
  ANDN U26224 ( .B(x[139]), .A(y[139]), .Z(n29047) );
  ANDN U26225 ( .B(n10635), .A(n29047), .Z(n10636) );
  NANDN U26226 ( .A(n29039), .B(n10636), .Z(n10637) );
  NANDN U26227 ( .A(x[140]), .B(y[140]), .Z(n29048) );
  AND U26228 ( .A(n10637), .B(n29048), .Z(n10638) );
  NAND U26229 ( .A(n29041), .B(n10638), .Z(n10639) );
  ANDN U26230 ( .B(x[141]), .A(y[141]), .Z(n29054) );
  ANDN U26231 ( .B(n10639), .A(n29054), .Z(n10640) );
  NANDN U26232 ( .A(n29044), .B(n10640), .Z(n10641) );
  NAND U26233 ( .A(n28490), .B(n10641), .Z(n10642) );
  NANDN U26234 ( .A(x[141]), .B(y[141]), .Z(n29049) );
  NANDN U26235 ( .A(n10642), .B(n29049), .Z(n10643) );
  AND U26236 ( .A(n10644), .B(n10643), .Z(n10646) );
  NANDN U26237 ( .A(x[143]), .B(y[143]), .Z(n28491) );
  NANDN U26238 ( .A(x[144]), .B(y[144]), .Z(n29064) );
  AND U26239 ( .A(n28491), .B(n29064), .Z(n10645) );
  NANDN U26240 ( .A(n10646), .B(n10645), .Z(n10647) );
  ANDN U26241 ( .B(x[145]), .A(y[145]), .Z(n29069) );
  ANDN U26242 ( .B(n10647), .A(n29069), .Z(n10648) );
  NANDN U26243 ( .A(n29061), .B(n10648), .Z(n10649) );
  NANDN U26244 ( .A(x[146]), .B(y[146]), .Z(n29070) );
  AND U26245 ( .A(n10649), .B(n29070), .Z(n10650) );
  NAND U26246 ( .A(n29063), .B(n10650), .Z(n10651) );
  ANDN U26247 ( .B(x[146]), .A(y[146]), .Z(n29066) );
  ANDN U26248 ( .B(n10651), .A(n29066), .Z(n10652) );
  NANDN U26249 ( .A(n29075), .B(n10652), .Z(n10653) );
  NAND U26250 ( .A(n29071), .B(n10653), .Z(n10654) );
  NANDN U26251 ( .A(x[148]), .B(y[148]), .Z(n29076) );
  NANDN U26252 ( .A(n10654), .B(n29076), .Z(n10655) );
  NANDN U26253 ( .A(n29079), .B(n10655), .Z(n10656) );
  NAND U26254 ( .A(n28488), .B(n10656), .Z(n10657) );
  NANDN U26255 ( .A(x[149]), .B(y[149]), .Z(n29081) );
  NANDN U26256 ( .A(n10657), .B(n29081), .Z(n10658) );
  AND U26257 ( .A(n10659), .B(n10658), .Z(n10661) );
  NANDN U26258 ( .A(x[151]), .B(y[151]), .Z(n28489) );
  NANDN U26259 ( .A(x[152]), .B(y[152]), .Z(n29092) );
  AND U26260 ( .A(n28489), .B(n29092), .Z(n10660) );
  NANDN U26261 ( .A(n10661), .B(n10660), .Z(n10662) );
  ANDN U26262 ( .B(x[153]), .A(y[153]), .Z(n29097) );
  ANDN U26263 ( .B(n10662), .A(n29097), .Z(n10663) );
  NANDN U26264 ( .A(n29089), .B(n10663), .Z(n10664) );
  NANDN U26265 ( .A(x[154]), .B(y[154]), .Z(n29098) );
  AND U26266 ( .A(n10664), .B(n29098), .Z(n10665) );
  NAND U26267 ( .A(n29091), .B(n10665), .Z(n10666) );
  ANDN U26268 ( .B(x[155]), .A(y[155]), .Z(n29104) );
  ANDN U26269 ( .B(n10666), .A(n29104), .Z(n10667) );
  NANDN U26270 ( .A(n29094), .B(n10667), .Z(n10668) );
  NAND U26271 ( .A(n28486), .B(n10668), .Z(n10669) );
  NANDN U26272 ( .A(x[155]), .B(y[155]), .Z(n29099) );
  NANDN U26273 ( .A(n10669), .B(n29099), .Z(n10670) );
  AND U26274 ( .A(n10671), .B(n10670), .Z(n10673) );
  NANDN U26275 ( .A(x[157]), .B(y[157]), .Z(n28487) );
  NANDN U26276 ( .A(x[158]), .B(y[158]), .Z(n29114) );
  AND U26277 ( .A(n28487), .B(n29114), .Z(n10672) );
  NANDN U26278 ( .A(n10673), .B(n10672), .Z(n10674) );
  ANDN U26279 ( .B(x[159]), .A(y[159]), .Z(n29119) );
  ANDN U26280 ( .B(n10674), .A(n29119), .Z(n10675) );
  NANDN U26281 ( .A(n29111), .B(n10675), .Z(n10676) );
  NANDN U26282 ( .A(x[160]), .B(y[160]), .Z(n29120) );
  AND U26283 ( .A(n10676), .B(n29120), .Z(n10677) );
  NAND U26284 ( .A(n29113), .B(n10677), .Z(n10678) );
  ANDN U26285 ( .B(x[161]), .A(y[161]), .Z(n29126) );
  ANDN U26286 ( .B(n10678), .A(n29126), .Z(n10679) );
  NANDN U26287 ( .A(n29116), .B(n10679), .Z(n10680) );
  NAND U26288 ( .A(n28484), .B(n10680), .Z(n10681) );
  NANDN U26289 ( .A(x[161]), .B(y[161]), .Z(n29121) );
  NANDN U26290 ( .A(n10681), .B(n29121), .Z(n10682) );
  AND U26291 ( .A(n10683), .B(n10682), .Z(n10685) );
  NANDN U26292 ( .A(x[163]), .B(y[163]), .Z(n28485) );
  NANDN U26293 ( .A(x[164]), .B(y[164]), .Z(n29136) );
  AND U26294 ( .A(n28485), .B(n29136), .Z(n10684) );
  NANDN U26295 ( .A(n10685), .B(n10684), .Z(n10686) );
  ANDN U26296 ( .B(x[165]), .A(y[165]), .Z(n29141) );
  ANDN U26297 ( .B(n10686), .A(n29141), .Z(n10687) );
  NANDN U26298 ( .A(n29133), .B(n10687), .Z(n10688) );
  NANDN U26299 ( .A(x[166]), .B(y[166]), .Z(n29142) );
  AND U26300 ( .A(n10688), .B(n29142), .Z(n10689) );
  NAND U26301 ( .A(n29135), .B(n10689), .Z(n10690) );
  ANDN U26302 ( .B(x[167]), .A(y[167]), .Z(n29148) );
  ANDN U26303 ( .B(n10690), .A(n29148), .Z(n10691) );
  NANDN U26304 ( .A(n29138), .B(n10691), .Z(n10692) );
  NAND U26305 ( .A(n28482), .B(n10692), .Z(n10693) );
  NANDN U26306 ( .A(x[167]), .B(y[167]), .Z(n29143) );
  NANDN U26307 ( .A(n10693), .B(n29143), .Z(n10694) );
  AND U26308 ( .A(n10695), .B(n10694), .Z(n10697) );
  NANDN U26309 ( .A(x[169]), .B(y[169]), .Z(n28483) );
  NANDN U26310 ( .A(x[170]), .B(y[170]), .Z(n29158) );
  AND U26311 ( .A(n28483), .B(n29158), .Z(n10696) );
  NANDN U26312 ( .A(n10697), .B(n10696), .Z(n10698) );
  ANDN U26313 ( .B(x[171]), .A(y[171]), .Z(n29160) );
  ANDN U26314 ( .B(n10698), .A(n29160), .Z(n10699) );
  NANDN U26315 ( .A(n29155), .B(n10699), .Z(n10700) );
  NANDN U26316 ( .A(x[171]), .B(y[171]), .Z(n29157) );
  AND U26317 ( .A(n10700), .B(n29157), .Z(n10701) );
  NANDN U26318 ( .A(n29163), .B(n10701), .Z(n10702) );
  ANDN U26319 ( .B(x[173]), .A(y[173]), .Z(n29170) );
  ANDN U26320 ( .B(n10702), .A(n29170), .Z(n10703) );
  NAND U26321 ( .A(n10704), .B(n10703), .Z(n10705) );
  NAND U26322 ( .A(n28480), .B(n10705), .Z(n10706) );
  NANDN U26323 ( .A(x[173]), .B(y[173]), .Z(n29165) );
  NANDN U26324 ( .A(n10706), .B(n29165), .Z(n10707) );
  AND U26325 ( .A(n10708), .B(n10707), .Z(n10710) );
  NANDN U26326 ( .A(x[175]), .B(y[175]), .Z(n28481) );
  NANDN U26327 ( .A(x[176]), .B(y[176]), .Z(n29180) );
  AND U26328 ( .A(n28481), .B(n29180), .Z(n10709) );
  NANDN U26329 ( .A(n10710), .B(n10709), .Z(n10711) );
  ANDN U26330 ( .B(x[177]), .A(y[177]), .Z(n29185) );
  ANDN U26331 ( .B(n10711), .A(n29185), .Z(n10712) );
  NANDN U26332 ( .A(n29177), .B(n10712), .Z(n10713) );
  NANDN U26333 ( .A(x[178]), .B(y[178]), .Z(n29186) );
  AND U26334 ( .A(n10713), .B(n29186), .Z(n10714) );
  NAND U26335 ( .A(n29179), .B(n10714), .Z(n10715) );
  ANDN U26336 ( .B(x[179]), .A(y[179]), .Z(n29192) );
  ANDN U26337 ( .B(n10715), .A(n29192), .Z(n10716) );
  NANDN U26338 ( .A(n29182), .B(n10716), .Z(n10717) );
  NAND U26339 ( .A(n28478), .B(n10717), .Z(n10718) );
  NANDN U26340 ( .A(x[179]), .B(y[179]), .Z(n29187) );
  NANDN U26341 ( .A(n10718), .B(n29187), .Z(n10719) );
  AND U26342 ( .A(n10720), .B(n10719), .Z(n10722) );
  NANDN U26343 ( .A(x[181]), .B(y[181]), .Z(n28479) );
  NANDN U26344 ( .A(x[182]), .B(y[182]), .Z(n29202) );
  AND U26345 ( .A(n28479), .B(n29202), .Z(n10721) );
  NANDN U26346 ( .A(n10722), .B(n10721), .Z(n10723) );
  ANDN U26347 ( .B(x[183]), .A(y[183]), .Z(n29207) );
  ANDN U26348 ( .B(n10723), .A(n29207), .Z(n10724) );
  NANDN U26349 ( .A(n29199), .B(n10724), .Z(n10725) );
  NANDN U26350 ( .A(x[184]), .B(y[184]), .Z(n29208) );
  AND U26351 ( .A(n10725), .B(n29208), .Z(n10726) );
  NAND U26352 ( .A(n29201), .B(n10726), .Z(n10727) );
  ANDN U26353 ( .B(x[185]), .A(y[185]), .Z(n29214) );
  ANDN U26354 ( .B(n10727), .A(n29214), .Z(n10728) );
  NANDN U26355 ( .A(n29204), .B(n10728), .Z(n10729) );
  NAND U26356 ( .A(n28476), .B(n10729), .Z(n10730) );
  NANDN U26357 ( .A(x[185]), .B(y[185]), .Z(n29209) );
  NANDN U26358 ( .A(n10730), .B(n29209), .Z(n10731) );
  AND U26359 ( .A(n10732), .B(n10731), .Z(n10734) );
  NANDN U26360 ( .A(x[187]), .B(y[187]), .Z(n28477) );
  NANDN U26361 ( .A(x[188]), .B(y[188]), .Z(n29223) );
  AND U26362 ( .A(n28477), .B(n29223), .Z(n10733) );
  NANDN U26363 ( .A(n10734), .B(n10733), .Z(n10735) );
  AND U26364 ( .A(n29227), .B(n10735), .Z(n10736) );
  NANDN U26365 ( .A(n29221), .B(n10736), .Z(n10737) );
  NAND U26366 ( .A(n10738), .B(n10737), .Z(n10741) );
  NANDN U26367 ( .A(y[191]), .B(x[191]), .Z(n10740) );
  NANDN U26368 ( .A(y[190]), .B(x[190]), .Z(n10739) );
  NAND U26369 ( .A(n10740), .B(n10739), .Z(n29230) );
  ANDN U26370 ( .B(n10741), .A(n29230), .Z(n10744) );
  NANDN U26371 ( .A(x[192]), .B(y[192]), .Z(n10743) );
  NANDN U26372 ( .A(x[191]), .B(y[191]), .Z(n10742) );
  AND U26373 ( .A(n10743), .B(n10742), .Z(n29233) );
  NANDN U26374 ( .A(n10744), .B(n29233), .Z(n10745) );
  NANDN U26375 ( .A(n29235), .B(n10745), .Z(n10746) );
  NAND U26376 ( .A(n29236), .B(n10746), .Z(n10747) );
  NANDN U26377 ( .A(n29239), .B(n10747), .Z(n10748) );
  NAND U26378 ( .A(n29242), .B(n10748), .Z(n10749) );
  ANDN U26379 ( .B(x[195]), .A(y[195]), .Z(n29247) );
  ANDN U26380 ( .B(n10749), .A(n29247), .Z(n10751) );
  NANDN U26381 ( .A(x[195]), .B(y[195]), .Z(n29241) );
  NANDN U26382 ( .A(x[196]), .B(y[196]), .Z(n29248) );
  AND U26383 ( .A(n29241), .B(n29248), .Z(n10750) );
  NANDN U26384 ( .A(n10751), .B(n10750), .Z(n10752) );
  ANDN U26385 ( .B(x[197]), .A(y[197]), .Z(n29254) );
  ANDN U26386 ( .B(n10752), .A(n29254), .Z(n10753) );
  NANDN U26387 ( .A(n29244), .B(n10753), .Z(n10754) );
  NANDN U26388 ( .A(x[198]), .B(y[198]), .Z(n28474) );
  AND U26389 ( .A(n10754), .B(n28474), .Z(n10755) );
  NAND U26390 ( .A(n29249), .B(n10755), .Z(n10756) );
  ANDN U26391 ( .B(x[199]), .A(y[199]), .Z(n29258) );
  ANDN U26392 ( .B(n10756), .A(n29258), .Z(n10757) );
  NANDN U26393 ( .A(n29253), .B(n10757), .Z(n10758) );
  NAND U26394 ( .A(n29264), .B(n10758), .Z(n10759) );
  NANDN U26395 ( .A(x[199]), .B(y[199]), .Z(n28475) );
  NANDN U26396 ( .A(n10759), .B(n28475), .Z(n10760) );
  AND U26397 ( .A(n10761), .B(n10760), .Z(n10763) );
  NANDN U26398 ( .A(x[201]), .B(y[201]), .Z(n29263) );
  NANDN U26399 ( .A(x[202]), .B(y[202]), .Z(n29270) );
  AND U26400 ( .A(n29263), .B(n29270), .Z(n10762) );
  NANDN U26401 ( .A(n10763), .B(n10762), .Z(n10764) );
  ANDN U26402 ( .B(x[203]), .A(y[203]), .Z(n29276) );
  ANDN U26403 ( .B(n10764), .A(n29276), .Z(n10765) );
  NANDN U26404 ( .A(n29266), .B(n10765), .Z(n10766) );
  NANDN U26405 ( .A(x[204]), .B(y[204]), .Z(n28472) );
  AND U26406 ( .A(n10766), .B(n28472), .Z(n10767) );
  NAND U26407 ( .A(n29271), .B(n10767), .Z(n10768) );
  ANDN U26408 ( .B(x[205]), .A(y[205]), .Z(n29280) );
  ANDN U26409 ( .B(n10768), .A(n29280), .Z(n10769) );
  NANDN U26410 ( .A(n29275), .B(n10769), .Z(n10770) );
  NAND U26411 ( .A(n29286), .B(n10770), .Z(n10771) );
  NANDN U26412 ( .A(x[205]), .B(y[205]), .Z(n28473) );
  NANDN U26413 ( .A(n10771), .B(n28473), .Z(n10772) );
  AND U26414 ( .A(n10773), .B(n10772), .Z(n10775) );
  NANDN U26415 ( .A(x[207]), .B(y[207]), .Z(n29285) );
  NANDN U26416 ( .A(x[208]), .B(y[208]), .Z(n29292) );
  AND U26417 ( .A(n29285), .B(n29292), .Z(n10774) );
  NANDN U26418 ( .A(n10775), .B(n10774), .Z(n10776) );
  ANDN U26419 ( .B(x[209]), .A(y[209]), .Z(n29298) );
  ANDN U26420 ( .B(n10776), .A(n29298), .Z(n10777) );
  NANDN U26421 ( .A(n29288), .B(n10777), .Z(n10778) );
  NANDN U26422 ( .A(x[210]), .B(y[210]), .Z(n28470) );
  AND U26423 ( .A(n10778), .B(n28470), .Z(n10779) );
  NAND U26424 ( .A(n29293), .B(n10779), .Z(n10780) );
  ANDN U26425 ( .B(x[211]), .A(y[211]), .Z(n29302) );
  ANDN U26426 ( .B(n10780), .A(n29302), .Z(n10781) );
  NANDN U26427 ( .A(n29297), .B(n10781), .Z(n10782) );
  NAND U26428 ( .A(n29308), .B(n10782), .Z(n10783) );
  NANDN U26429 ( .A(x[211]), .B(y[211]), .Z(n28471) );
  NANDN U26430 ( .A(n10783), .B(n28471), .Z(n10784) );
  AND U26431 ( .A(n10785), .B(n10784), .Z(n10787) );
  NANDN U26432 ( .A(x[213]), .B(y[213]), .Z(n29307) );
  NANDN U26433 ( .A(x[214]), .B(y[214]), .Z(n29314) );
  AND U26434 ( .A(n29307), .B(n29314), .Z(n10786) );
  NANDN U26435 ( .A(n10787), .B(n10786), .Z(n10788) );
  ANDN U26436 ( .B(x[215]), .A(y[215]), .Z(n29320) );
  ANDN U26437 ( .B(n10788), .A(n29320), .Z(n10789) );
  NANDN U26438 ( .A(n29310), .B(n10789), .Z(n10790) );
  NANDN U26439 ( .A(x[216]), .B(y[216]), .Z(n28468) );
  AND U26440 ( .A(n10790), .B(n28468), .Z(n10791) );
  NAND U26441 ( .A(n29315), .B(n10791), .Z(n10792) );
  ANDN U26442 ( .B(x[217]), .A(y[217]), .Z(n29324) );
  ANDN U26443 ( .B(n10792), .A(n29324), .Z(n10793) );
  NANDN U26444 ( .A(n29319), .B(n10793), .Z(n10794) );
  NAND U26445 ( .A(n29330), .B(n10794), .Z(n10795) );
  NANDN U26446 ( .A(x[217]), .B(y[217]), .Z(n28469) );
  NANDN U26447 ( .A(n10795), .B(n28469), .Z(n10796) );
  AND U26448 ( .A(n10797), .B(n10796), .Z(n10799) );
  NANDN U26449 ( .A(x[219]), .B(y[219]), .Z(n29329) );
  NANDN U26450 ( .A(x[220]), .B(y[220]), .Z(n29336) );
  AND U26451 ( .A(n29329), .B(n29336), .Z(n10798) );
  NANDN U26452 ( .A(n10799), .B(n10798), .Z(n10800) );
  ANDN U26453 ( .B(x[221]), .A(y[221]), .Z(n29342) );
  ANDN U26454 ( .B(n10800), .A(n29342), .Z(n10801) );
  NANDN U26455 ( .A(n29332), .B(n10801), .Z(n10802) );
  NANDN U26456 ( .A(x[222]), .B(y[222]), .Z(n28466) );
  AND U26457 ( .A(n10802), .B(n28466), .Z(n10803) );
  NAND U26458 ( .A(n29337), .B(n10803), .Z(n10804) );
  ANDN U26459 ( .B(x[223]), .A(y[223]), .Z(n29346) );
  ANDN U26460 ( .B(n10804), .A(n29346), .Z(n10805) );
  NANDN U26461 ( .A(n29341), .B(n10805), .Z(n10806) );
  NAND U26462 ( .A(n29352), .B(n10806), .Z(n10807) );
  NANDN U26463 ( .A(x[223]), .B(y[223]), .Z(n28467) );
  NANDN U26464 ( .A(n10807), .B(n28467), .Z(n10808) );
  AND U26465 ( .A(n10809), .B(n10808), .Z(n10811) );
  NANDN U26466 ( .A(x[225]), .B(y[225]), .Z(n29351) );
  NANDN U26467 ( .A(x[226]), .B(y[226]), .Z(n29361) );
  AND U26468 ( .A(n29351), .B(n29361), .Z(n10810) );
  NANDN U26469 ( .A(n10811), .B(n10810), .Z(n10812) );
  ANDN U26470 ( .B(x[227]), .A(y[227]), .Z(n29364) );
  ANDN U26471 ( .B(n10812), .A(n29364), .Z(n10813) );
  NANDN U26472 ( .A(n29354), .B(n10813), .Z(n10814) );
  NANDN U26473 ( .A(x[227]), .B(y[227]), .Z(n29359) );
  AND U26474 ( .A(n10814), .B(n29359), .Z(n10815) );
  NANDN U26475 ( .A(n29363), .B(n10815), .Z(n10816) );
  ANDN U26476 ( .B(x[229]), .A(y[229]), .Z(n29368) );
  ANDN U26477 ( .B(n10816), .A(n29368), .Z(n10817) );
  NAND U26478 ( .A(n10818), .B(n10817), .Z(n10819) );
  NAND U26479 ( .A(n29374), .B(n10819), .Z(n10820) );
  NANDN U26480 ( .A(x[229]), .B(y[229]), .Z(n28464) );
  NANDN U26481 ( .A(n10820), .B(n28464), .Z(n10821) );
  AND U26482 ( .A(n10822), .B(n10821), .Z(n10824) );
  NANDN U26483 ( .A(x[231]), .B(y[231]), .Z(n29373) );
  NANDN U26484 ( .A(x[232]), .B(y[232]), .Z(n29380) );
  AND U26485 ( .A(n29373), .B(n29380), .Z(n10823) );
  NANDN U26486 ( .A(n10824), .B(n10823), .Z(n10825) );
  ANDN U26487 ( .B(x[233]), .A(y[233]), .Z(n29386) );
  ANDN U26488 ( .B(n10825), .A(n29386), .Z(n10826) );
  NANDN U26489 ( .A(n29376), .B(n10826), .Z(n10827) );
  NANDN U26490 ( .A(x[234]), .B(y[234]), .Z(n28462) );
  AND U26491 ( .A(n10827), .B(n28462), .Z(n10828) );
  NAND U26492 ( .A(n29381), .B(n10828), .Z(n10829) );
  ANDN U26493 ( .B(x[235]), .A(y[235]), .Z(n29390) );
  ANDN U26494 ( .B(n10829), .A(n29390), .Z(n10830) );
  NANDN U26495 ( .A(n29385), .B(n10830), .Z(n10831) );
  NAND U26496 ( .A(n29396), .B(n10831), .Z(n10832) );
  NANDN U26497 ( .A(x[235]), .B(y[235]), .Z(n28463) );
  NANDN U26498 ( .A(n10832), .B(n28463), .Z(n10833) );
  AND U26499 ( .A(n10834), .B(n10833), .Z(n10836) );
  NANDN U26500 ( .A(x[237]), .B(y[237]), .Z(n29395) );
  NANDN U26501 ( .A(x[238]), .B(y[238]), .Z(n29402) );
  AND U26502 ( .A(n29395), .B(n29402), .Z(n10835) );
  NANDN U26503 ( .A(n10836), .B(n10835), .Z(n10837) );
  ANDN U26504 ( .B(x[239]), .A(y[239]), .Z(n29408) );
  ANDN U26505 ( .B(n10837), .A(n29408), .Z(n10838) );
  NANDN U26506 ( .A(n29398), .B(n10838), .Z(n10839) );
  NANDN U26507 ( .A(x[240]), .B(y[240]), .Z(n28460) );
  AND U26508 ( .A(n10839), .B(n28460), .Z(n10840) );
  NAND U26509 ( .A(n29403), .B(n10840), .Z(n10841) );
  ANDN U26510 ( .B(x[241]), .A(y[241]), .Z(n29412) );
  ANDN U26511 ( .B(n10841), .A(n29412), .Z(n10842) );
  NANDN U26512 ( .A(n29407), .B(n10842), .Z(n10843) );
  NAND U26513 ( .A(n29418), .B(n10843), .Z(n10844) );
  NANDN U26514 ( .A(x[241]), .B(y[241]), .Z(n28461) );
  NANDN U26515 ( .A(n10844), .B(n28461), .Z(n10845) );
  AND U26516 ( .A(n10846), .B(n10845), .Z(n10848) );
  NANDN U26517 ( .A(x[243]), .B(y[243]), .Z(n29417) );
  NANDN U26518 ( .A(x[244]), .B(y[244]), .Z(n29424) );
  AND U26519 ( .A(n29417), .B(n29424), .Z(n10847) );
  NANDN U26520 ( .A(n10848), .B(n10847), .Z(n10849) );
  ANDN U26521 ( .B(x[245]), .A(y[245]), .Z(n29430) );
  ANDN U26522 ( .B(n10849), .A(n29430), .Z(n10850) );
  NANDN U26523 ( .A(n29420), .B(n10850), .Z(n10851) );
  NANDN U26524 ( .A(x[246]), .B(y[246]), .Z(n28458) );
  AND U26525 ( .A(n10851), .B(n28458), .Z(n10852) );
  NAND U26526 ( .A(n29425), .B(n10852), .Z(n10853) );
  ANDN U26527 ( .B(x[247]), .A(y[247]), .Z(n29434) );
  ANDN U26528 ( .B(n10853), .A(n29434), .Z(n10854) );
  NANDN U26529 ( .A(n29429), .B(n10854), .Z(n10855) );
  NAND U26530 ( .A(n29440), .B(n10855), .Z(n10856) );
  NANDN U26531 ( .A(x[247]), .B(y[247]), .Z(n28459) );
  NANDN U26532 ( .A(n10856), .B(n28459), .Z(n10857) );
  AND U26533 ( .A(n10858), .B(n10857), .Z(n10860) );
  NANDN U26534 ( .A(x[249]), .B(y[249]), .Z(n29439) );
  NANDN U26535 ( .A(x[250]), .B(y[250]), .Z(n29446) );
  AND U26536 ( .A(n29439), .B(n29446), .Z(n10859) );
  NANDN U26537 ( .A(n10860), .B(n10859), .Z(n10861) );
  ANDN U26538 ( .B(x[251]), .A(y[251]), .Z(n29452) );
  ANDN U26539 ( .B(n10861), .A(n29452), .Z(n10862) );
  NANDN U26540 ( .A(n29442), .B(n10862), .Z(n10863) );
  NANDN U26541 ( .A(x[252]), .B(y[252]), .Z(n28456) );
  AND U26542 ( .A(n10863), .B(n28456), .Z(n10864) );
  NAND U26543 ( .A(n29447), .B(n10864), .Z(n10865) );
  ANDN U26544 ( .B(x[253]), .A(y[253]), .Z(n29456) );
  ANDN U26545 ( .B(n10865), .A(n29456), .Z(n10866) );
  NANDN U26546 ( .A(n29451), .B(n10866), .Z(n10867) );
  NAND U26547 ( .A(n29462), .B(n10867), .Z(n10868) );
  NANDN U26548 ( .A(x[253]), .B(y[253]), .Z(n28457) );
  NANDN U26549 ( .A(n10868), .B(n28457), .Z(n10869) );
  AND U26550 ( .A(n10870), .B(n10869), .Z(n10872) );
  NANDN U26551 ( .A(x[255]), .B(y[255]), .Z(n29461) );
  NANDN U26552 ( .A(x[256]), .B(y[256]), .Z(n29468) );
  AND U26553 ( .A(n29461), .B(n29468), .Z(n10871) );
  NANDN U26554 ( .A(n10872), .B(n10871), .Z(n10873) );
  ANDN U26555 ( .B(x[257]), .A(y[257]), .Z(n29474) );
  ANDN U26556 ( .B(n10873), .A(n29474), .Z(n10874) );
  NANDN U26557 ( .A(n29464), .B(n10874), .Z(n10875) );
  NANDN U26558 ( .A(x[258]), .B(y[258]), .Z(n28454) );
  AND U26559 ( .A(n10875), .B(n28454), .Z(n10876) );
  NAND U26560 ( .A(n29469), .B(n10876), .Z(n10877) );
  ANDN U26561 ( .B(x[259]), .A(y[259]), .Z(n29478) );
  ANDN U26562 ( .B(n10877), .A(n29478), .Z(n10878) );
  NANDN U26563 ( .A(n29473), .B(n10878), .Z(n10879) );
  NAND U26564 ( .A(n29484), .B(n10879), .Z(n10880) );
  NANDN U26565 ( .A(x[259]), .B(y[259]), .Z(n28455) );
  NANDN U26566 ( .A(n10880), .B(n28455), .Z(n10881) );
  AND U26567 ( .A(n10882), .B(n10881), .Z(n10884) );
  NANDN U26568 ( .A(x[261]), .B(y[261]), .Z(n29483) );
  NANDN U26569 ( .A(x[262]), .B(y[262]), .Z(n29490) );
  AND U26570 ( .A(n29483), .B(n29490), .Z(n10883) );
  NANDN U26571 ( .A(n10884), .B(n10883), .Z(n10885) );
  ANDN U26572 ( .B(x[263]), .A(y[263]), .Z(n29495) );
  ANDN U26573 ( .B(n10885), .A(n29495), .Z(n10886) );
  NANDN U26574 ( .A(n29486), .B(n10886), .Z(n10888) );
  ANDN U26575 ( .B(y[264]), .A(x[264]), .Z(n10887) );
  ANDN U26576 ( .B(n10888), .A(n10887), .Z(n10889) );
  NAND U26577 ( .A(n29491), .B(n10889), .Z(n10890) );
  NAND U26578 ( .A(n10891), .B(n10890), .Z(n10892) );
  NAND U26579 ( .A(n29503), .B(n10892), .Z(n10895) );
  NANDN U26580 ( .A(y[267]), .B(x[267]), .Z(n10894) );
  NANDN U26581 ( .A(y[266]), .B(x[266]), .Z(n10893) );
  NAND U26582 ( .A(n10894), .B(n10893), .Z(n29505) );
  ANDN U26583 ( .B(n10895), .A(n29505), .Z(n10898) );
  NANDN U26584 ( .A(x[267]), .B(y[267]), .Z(n10897) );
  NANDN U26585 ( .A(x[268]), .B(y[268]), .Z(n10896) );
  AND U26586 ( .A(n10897), .B(n10896), .Z(n29507) );
  NANDN U26587 ( .A(n10898), .B(n29507), .Z(n10899) );
  NANDN U26588 ( .A(n29509), .B(n10899), .Z(n10900) );
  NAND U26589 ( .A(n29511), .B(n10900), .Z(n10901) );
  NANDN U26590 ( .A(n29513), .B(n10901), .Z(n10902) );
  NANDN U26591 ( .A(x[271]), .B(y[271]), .Z(n29514) );
  AND U26592 ( .A(n10902), .B(n29514), .Z(n10903) );
  NAND U26593 ( .A(n29520), .B(n10903), .Z(n10904) );
  ANDN U26594 ( .B(x[273]), .A(y[273]), .Z(n29525) );
  ANDN U26595 ( .B(n10904), .A(n29525), .Z(n10905) );
  NANDN U26596 ( .A(n29517), .B(n10905), .Z(n10906) );
  NAND U26597 ( .A(n29519), .B(n10906), .Z(n10908) );
  NANDN U26598 ( .A(x[274]), .B(n10908), .Z(n10907) );
  NANDN U26599 ( .A(x[275]), .B(y[275]), .Z(n28453) );
  AND U26600 ( .A(n10907), .B(n28453), .Z(n10911) );
  XNOR U26601 ( .A(n10908), .B(x[274]), .Z(n10909) );
  NAND U26602 ( .A(n10909), .B(y[274]), .Z(n10910) );
  NAND U26603 ( .A(n10911), .B(n10910), .Z(n10912) );
  NANDN U26604 ( .A(n29529), .B(n10912), .Z(n10913) );
  NAND U26605 ( .A(n29532), .B(n10913), .Z(n10914) );
  ANDN U26606 ( .B(x[277]), .A(y[277]), .Z(n29537) );
  ANDN U26607 ( .B(n10914), .A(n29537), .Z(n10916) );
  NANDN U26608 ( .A(x[277]), .B(y[277]), .Z(n29531) );
  NANDN U26609 ( .A(x[278]), .B(y[278]), .Z(n29538) );
  AND U26610 ( .A(n29531), .B(n29538), .Z(n10915) );
  NANDN U26611 ( .A(n10916), .B(n10915), .Z(n10917) );
  ANDN U26612 ( .B(x[279]), .A(y[279]), .Z(n29544) );
  ANDN U26613 ( .B(n10917), .A(n29544), .Z(n10918) );
  NANDN U26614 ( .A(n29534), .B(n10918), .Z(n10919) );
  NANDN U26615 ( .A(x[280]), .B(y[280]), .Z(n28450) );
  AND U26616 ( .A(n10919), .B(n28450), .Z(n10920) );
  NAND U26617 ( .A(n29539), .B(n10920), .Z(n10921) );
  ANDN U26618 ( .B(x[281]), .A(y[281]), .Z(n29548) );
  ANDN U26619 ( .B(n10921), .A(n29548), .Z(n10922) );
  NANDN U26620 ( .A(n29543), .B(n10922), .Z(n10923) );
  NAND U26621 ( .A(n29554), .B(n10923), .Z(n10924) );
  NANDN U26622 ( .A(x[281]), .B(y[281]), .Z(n28451) );
  NANDN U26623 ( .A(n10924), .B(n28451), .Z(n10925) );
  AND U26624 ( .A(n10926), .B(n10925), .Z(n10928) );
  NANDN U26625 ( .A(x[283]), .B(y[283]), .Z(n29553) );
  NANDN U26626 ( .A(x[284]), .B(y[284]), .Z(n29560) );
  AND U26627 ( .A(n29553), .B(n29560), .Z(n10927) );
  NANDN U26628 ( .A(n10928), .B(n10927), .Z(n10929) );
  ANDN U26629 ( .B(x[285]), .A(y[285]), .Z(n29566) );
  ANDN U26630 ( .B(n10929), .A(n29566), .Z(n10930) );
  NANDN U26631 ( .A(n29556), .B(n10930), .Z(n10931) );
  NANDN U26632 ( .A(x[286]), .B(y[286]), .Z(n28448) );
  AND U26633 ( .A(n10931), .B(n28448), .Z(n10932) );
  NAND U26634 ( .A(n29561), .B(n10932), .Z(n10933) );
  ANDN U26635 ( .B(x[287]), .A(y[287]), .Z(n29570) );
  ANDN U26636 ( .B(n10933), .A(n29570), .Z(n10934) );
  NANDN U26637 ( .A(n29565), .B(n10934), .Z(n10935) );
  NAND U26638 ( .A(n29576), .B(n10935), .Z(n10936) );
  NANDN U26639 ( .A(x[287]), .B(y[287]), .Z(n28449) );
  NANDN U26640 ( .A(n10936), .B(n28449), .Z(n10937) );
  AND U26641 ( .A(n10938), .B(n10937), .Z(n10940) );
  NANDN U26642 ( .A(x[289]), .B(y[289]), .Z(n29575) );
  NANDN U26643 ( .A(x[290]), .B(y[290]), .Z(n29582) );
  AND U26644 ( .A(n29575), .B(n29582), .Z(n10939) );
  NANDN U26645 ( .A(n10940), .B(n10939), .Z(n10941) );
  ANDN U26646 ( .B(x[291]), .A(y[291]), .Z(n29588) );
  ANDN U26647 ( .B(n10941), .A(n29588), .Z(n10942) );
  NANDN U26648 ( .A(n29578), .B(n10942), .Z(n10943) );
  NANDN U26649 ( .A(x[292]), .B(y[292]), .Z(n28446) );
  AND U26650 ( .A(n10943), .B(n28446), .Z(n10944) );
  NAND U26651 ( .A(n29583), .B(n10944), .Z(n10945) );
  ANDN U26652 ( .B(x[293]), .A(y[293]), .Z(n29592) );
  ANDN U26653 ( .B(n10945), .A(n29592), .Z(n10946) );
  NANDN U26654 ( .A(n29587), .B(n10946), .Z(n10947) );
  NAND U26655 ( .A(n29598), .B(n10947), .Z(n10948) );
  NANDN U26656 ( .A(x[293]), .B(y[293]), .Z(n28447) );
  NANDN U26657 ( .A(n10948), .B(n28447), .Z(n10949) );
  AND U26658 ( .A(n10950), .B(n10949), .Z(n10952) );
  NANDN U26659 ( .A(x[295]), .B(y[295]), .Z(n29597) );
  NANDN U26660 ( .A(x[296]), .B(y[296]), .Z(n29604) );
  AND U26661 ( .A(n29597), .B(n29604), .Z(n10951) );
  NANDN U26662 ( .A(n10952), .B(n10951), .Z(n10953) );
  ANDN U26663 ( .B(x[297]), .A(y[297]), .Z(n29610) );
  ANDN U26664 ( .B(n10953), .A(n29610), .Z(n10954) );
  NANDN U26665 ( .A(n29600), .B(n10954), .Z(n10955) );
  NANDN U26666 ( .A(x[298]), .B(y[298]), .Z(n28444) );
  AND U26667 ( .A(n10955), .B(n28444), .Z(n10956) );
  NAND U26668 ( .A(n29605), .B(n10956), .Z(n10957) );
  ANDN U26669 ( .B(x[299]), .A(y[299]), .Z(n29614) );
  ANDN U26670 ( .B(n10957), .A(n29614), .Z(n10958) );
  NANDN U26671 ( .A(n29609), .B(n10958), .Z(n10959) );
  NAND U26672 ( .A(n29620), .B(n10959), .Z(n10960) );
  NANDN U26673 ( .A(x[299]), .B(y[299]), .Z(n28445) );
  NANDN U26674 ( .A(n10960), .B(n28445), .Z(n10961) );
  AND U26675 ( .A(n10962), .B(n10961), .Z(n10964) );
  NANDN U26676 ( .A(x[301]), .B(y[301]), .Z(n29619) );
  NANDN U26677 ( .A(x[302]), .B(y[302]), .Z(n29626) );
  AND U26678 ( .A(n29619), .B(n29626), .Z(n10963) );
  NANDN U26679 ( .A(n10964), .B(n10963), .Z(n10965) );
  ANDN U26680 ( .B(x[303]), .A(y[303]), .Z(n29632) );
  ANDN U26681 ( .B(n10965), .A(n29632), .Z(n10966) );
  NANDN U26682 ( .A(n29622), .B(n10966), .Z(n10967) );
  NANDN U26683 ( .A(x[304]), .B(y[304]), .Z(n28442) );
  AND U26684 ( .A(n10967), .B(n28442), .Z(n10968) );
  NAND U26685 ( .A(n29627), .B(n10968), .Z(n10969) );
  ANDN U26686 ( .B(x[305]), .A(y[305]), .Z(n29636) );
  ANDN U26687 ( .B(n10969), .A(n29636), .Z(n10970) );
  NANDN U26688 ( .A(n29631), .B(n10970), .Z(n10971) );
  NAND U26689 ( .A(n29642), .B(n10971), .Z(n10972) );
  NANDN U26690 ( .A(x[305]), .B(y[305]), .Z(n28443) );
  NANDN U26691 ( .A(n10972), .B(n28443), .Z(n10973) );
  AND U26692 ( .A(n10974), .B(n10973), .Z(n10976) );
  NANDN U26693 ( .A(x[307]), .B(y[307]), .Z(n29641) );
  NANDN U26694 ( .A(x[308]), .B(y[308]), .Z(n29648) );
  AND U26695 ( .A(n29641), .B(n29648), .Z(n10975) );
  NANDN U26696 ( .A(n10976), .B(n10975), .Z(n10977) );
  ANDN U26697 ( .B(x[309]), .A(y[309]), .Z(n29654) );
  ANDN U26698 ( .B(n10977), .A(n29654), .Z(n10978) );
  NANDN U26699 ( .A(n29644), .B(n10978), .Z(n10979) );
  NANDN U26700 ( .A(x[310]), .B(y[310]), .Z(n28440) );
  AND U26701 ( .A(n10979), .B(n28440), .Z(n10980) );
  NAND U26702 ( .A(n29649), .B(n10980), .Z(n10981) );
  ANDN U26703 ( .B(x[311]), .A(y[311]), .Z(n29658) );
  ANDN U26704 ( .B(n10981), .A(n29658), .Z(n10982) );
  NANDN U26705 ( .A(n29653), .B(n10982), .Z(n10983) );
  NAND U26706 ( .A(n29664), .B(n10983), .Z(n10984) );
  NANDN U26707 ( .A(x[311]), .B(y[311]), .Z(n28441) );
  NANDN U26708 ( .A(n10984), .B(n28441), .Z(n10985) );
  AND U26709 ( .A(n10986), .B(n10985), .Z(n10988) );
  NANDN U26710 ( .A(x[313]), .B(y[313]), .Z(n29663) );
  NANDN U26711 ( .A(x[314]), .B(y[314]), .Z(n29670) );
  AND U26712 ( .A(n29663), .B(n29670), .Z(n10987) );
  NANDN U26713 ( .A(n10988), .B(n10987), .Z(n10989) );
  ANDN U26714 ( .B(x[315]), .A(y[315]), .Z(n29676) );
  ANDN U26715 ( .B(n10989), .A(n29676), .Z(n10990) );
  NANDN U26716 ( .A(n29666), .B(n10990), .Z(n10991) );
  NANDN U26717 ( .A(x[316]), .B(y[316]), .Z(n28438) );
  AND U26718 ( .A(n10991), .B(n28438), .Z(n10992) );
  NAND U26719 ( .A(n29671), .B(n10992), .Z(n10993) );
  ANDN U26720 ( .B(x[317]), .A(y[317]), .Z(n29680) );
  ANDN U26721 ( .B(n10993), .A(n29680), .Z(n10994) );
  NANDN U26722 ( .A(n29675), .B(n10994), .Z(n10995) );
  NAND U26723 ( .A(n29686), .B(n10995), .Z(n10996) );
  NANDN U26724 ( .A(x[317]), .B(y[317]), .Z(n28439) );
  NANDN U26725 ( .A(n10996), .B(n28439), .Z(n10997) );
  AND U26726 ( .A(n10998), .B(n10997), .Z(n11000) );
  NANDN U26727 ( .A(x[319]), .B(y[319]), .Z(n29685) );
  NANDN U26728 ( .A(x[320]), .B(y[320]), .Z(n29692) );
  AND U26729 ( .A(n29685), .B(n29692), .Z(n10999) );
  NANDN U26730 ( .A(n11000), .B(n10999), .Z(n11001) );
  ANDN U26731 ( .B(x[321]), .A(y[321]), .Z(n29698) );
  ANDN U26732 ( .B(n11001), .A(n29698), .Z(n11002) );
  NANDN U26733 ( .A(n29688), .B(n11002), .Z(n11003) );
  NANDN U26734 ( .A(x[322]), .B(y[322]), .Z(n28436) );
  AND U26735 ( .A(n11003), .B(n28436), .Z(n11004) );
  NAND U26736 ( .A(n29693), .B(n11004), .Z(n11005) );
  ANDN U26737 ( .B(x[323]), .A(y[323]), .Z(n29702) );
  ANDN U26738 ( .B(n11005), .A(n29702), .Z(n11006) );
  NANDN U26739 ( .A(n29697), .B(n11006), .Z(n11007) );
  NAND U26740 ( .A(n29708), .B(n11007), .Z(n11008) );
  NANDN U26741 ( .A(x[323]), .B(y[323]), .Z(n28437) );
  NANDN U26742 ( .A(n11008), .B(n28437), .Z(n11009) );
  AND U26743 ( .A(n11010), .B(n11009), .Z(n11012) );
  NANDN U26744 ( .A(x[325]), .B(y[325]), .Z(n29707) );
  NANDN U26745 ( .A(x[326]), .B(y[326]), .Z(n29714) );
  AND U26746 ( .A(n29707), .B(n29714), .Z(n11011) );
  NANDN U26747 ( .A(n11012), .B(n11011), .Z(n11013) );
  ANDN U26748 ( .B(x[327]), .A(y[327]), .Z(n29720) );
  ANDN U26749 ( .B(n11013), .A(n29720), .Z(n11014) );
  NANDN U26750 ( .A(n29710), .B(n11014), .Z(n11015) );
  NANDN U26751 ( .A(x[328]), .B(y[328]), .Z(n28434) );
  AND U26752 ( .A(n11015), .B(n28434), .Z(n11016) );
  NAND U26753 ( .A(n29715), .B(n11016), .Z(n11017) );
  ANDN U26754 ( .B(x[329]), .A(y[329]), .Z(n29724) );
  ANDN U26755 ( .B(n11017), .A(n29724), .Z(n11018) );
  NANDN U26756 ( .A(n29719), .B(n11018), .Z(n11019) );
  NAND U26757 ( .A(n29730), .B(n11019), .Z(n11020) );
  NANDN U26758 ( .A(x[329]), .B(y[329]), .Z(n28435) );
  NANDN U26759 ( .A(n11020), .B(n28435), .Z(n11021) );
  AND U26760 ( .A(n11022), .B(n11021), .Z(n11024) );
  NANDN U26761 ( .A(x[331]), .B(y[331]), .Z(n29729) );
  NANDN U26762 ( .A(x[332]), .B(y[332]), .Z(n29736) );
  AND U26763 ( .A(n29729), .B(n29736), .Z(n11023) );
  NANDN U26764 ( .A(n11024), .B(n11023), .Z(n11025) );
  ANDN U26765 ( .B(x[333]), .A(y[333]), .Z(n29742) );
  ANDN U26766 ( .B(n11025), .A(n29742), .Z(n11026) );
  NANDN U26767 ( .A(n29732), .B(n11026), .Z(n11027) );
  NANDN U26768 ( .A(x[334]), .B(y[334]), .Z(n28432) );
  AND U26769 ( .A(n11027), .B(n28432), .Z(n11028) );
  NAND U26770 ( .A(n29737), .B(n11028), .Z(n11029) );
  ANDN U26771 ( .B(x[335]), .A(y[335]), .Z(n29746) );
  ANDN U26772 ( .B(n11029), .A(n29746), .Z(n11030) );
  NANDN U26773 ( .A(n29741), .B(n11030), .Z(n11031) );
  NAND U26774 ( .A(n29752), .B(n11031), .Z(n11032) );
  NANDN U26775 ( .A(x[335]), .B(y[335]), .Z(n28433) );
  NANDN U26776 ( .A(n11032), .B(n28433), .Z(n11033) );
  AND U26777 ( .A(n11034), .B(n11033), .Z(n11036) );
  NANDN U26778 ( .A(x[337]), .B(y[337]), .Z(n29751) );
  XOR U26779 ( .A(y[338]), .B(x[338]), .Z(n29757) );
  ANDN U26780 ( .B(n29751), .A(n29757), .Z(n11035) );
  NANDN U26781 ( .A(n11036), .B(n11035), .Z(n11037) );
  ANDN U26782 ( .B(x[339]), .A(y[339]), .Z(n29764) );
  ANDN U26783 ( .B(n11037), .A(n29764), .Z(n11039) );
  NANDN U26784 ( .A(y[338]), .B(x[338]), .Z(n11038) );
  NAND U26785 ( .A(n11039), .B(n11038), .Z(n11040) );
  NANDN U26786 ( .A(x[340]), .B(y[340]), .Z(n28430) );
  AND U26787 ( .A(n11040), .B(n28430), .Z(n11041) );
  NAND U26788 ( .A(n29759), .B(n11041), .Z(n11042) );
  ANDN U26789 ( .B(x[341]), .A(y[341]), .Z(n29768) );
  ANDN U26790 ( .B(n11042), .A(n29768), .Z(n11043) );
  NANDN U26791 ( .A(n29763), .B(n11043), .Z(n11044) );
  NAND U26792 ( .A(n29774), .B(n11044), .Z(n11045) );
  NANDN U26793 ( .A(x[341]), .B(y[341]), .Z(n28431) );
  NANDN U26794 ( .A(n11045), .B(n28431), .Z(n11046) );
  AND U26795 ( .A(n11047), .B(n11046), .Z(n11049) );
  NANDN U26796 ( .A(x[343]), .B(y[343]), .Z(n29773) );
  NANDN U26797 ( .A(x[344]), .B(y[344]), .Z(n29780) );
  AND U26798 ( .A(n29773), .B(n29780), .Z(n11048) );
  NANDN U26799 ( .A(n11049), .B(n11048), .Z(n11050) );
  ANDN U26800 ( .B(x[345]), .A(y[345]), .Z(n29786) );
  ANDN U26801 ( .B(n11050), .A(n29786), .Z(n11051) );
  NANDN U26802 ( .A(n29776), .B(n11051), .Z(n11052) );
  NANDN U26803 ( .A(x[346]), .B(y[346]), .Z(n28428) );
  AND U26804 ( .A(n11052), .B(n28428), .Z(n11053) );
  NAND U26805 ( .A(n29781), .B(n11053), .Z(n11054) );
  ANDN U26806 ( .B(x[347]), .A(y[347]), .Z(n29790) );
  ANDN U26807 ( .B(n11054), .A(n29790), .Z(n11055) );
  NANDN U26808 ( .A(n29785), .B(n11055), .Z(n11056) );
  NAND U26809 ( .A(n29796), .B(n11056), .Z(n11057) );
  NANDN U26810 ( .A(x[347]), .B(y[347]), .Z(n28429) );
  NANDN U26811 ( .A(n11057), .B(n28429), .Z(n11058) );
  AND U26812 ( .A(n11059), .B(n11058), .Z(n11061) );
  NANDN U26813 ( .A(x[349]), .B(y[349]), .Z(n29795) );
  XOR U26814 ( .A(y[350]), .B(x[350]), .Z(n29801) );
  ANDN U26815 ( .B(n29795), .A(n29801), .Z(n11060) );
  NANDN U26816 ( .A(n11061), .B(n11060), .Z(n11062) );
  ANDN U26817 ( .B(x[351]), .A(y[351]), .Z(n29808) );
  ANDN U26818 ( .B(n11062), .A(n29808), .Z(n11064) );
  NANDN U26819 ( .A(y[350]), .B(x[350]), .Z(n11063) );
  NAND U26820 ( .A(n11064), .B(n11063), .Z(n11065) );
  NANDN U26821 ( .A(x[352]), .B(y[352]), .Z(n28426) );
  AND U26822 ( .A(n11065), .B(n28426), .Z(n11066) );
  NAND U26823 ( .A(n29803), .B(n11066), .Z(n11067) );
  ANDN U26824 ( .B(x[353]), .A(y[353]), .Z(n29812) );
  ANDN U26825 ( .B(n11067), .A(n29812), .Z(n11068) );
  NANDN U26826 ( .A(n29807), .B(n11068), .Z(n11069) );
  NAND U26827 ( .A(n29818), .B(n11069), .Z(n11070) );
  NANDN U26828 ( .A(x[353]), .B(y[353]), .Z(n28427) );
  NANDN U26829 ( .A(n11070), .B(n28427), .Z(n11071) );
  AND U26830 ( .A(n11072), .B(n11071), .Z(n11074) );
  NANDN U26831 ( .A(x[355]), .B(y[355]), .Z(n29817) );
  NANDN U26832 ( .A(x[356]), .B(y[356]), .Z(n29824) );
  AND U26833 ( .A(n29817), .B(n29824), .Z(n11073) );
  NANDN U26834 ( .A(n11074), .B(n11073), .Z(n11075) );
  ANDN U26835 ( .B(x[357]), .A(y[357]), .Z(n29830) );
  ANDN U26836 ( .B(n11075), .A(n29830), .Z(n11076) );
  NANDN U26837 ( .A(n29820), .B(n11076), .Z(n11077) );
  NANDN U26838 ( .A(x[358]), .B(y[358]), .Z(n28424) );
  AND U26839 ( .A(n11077), .B(n28424), .Z(n11078) );
  NAND U26840 ( .A(n29825), .B(n11078), .Z(n11079) );
  ANDN U26841 ( .B(x[359]), .A(y[359]), .Z(n29834) );
  ANDN U26842 ( .B(n11079), .A(n29834), .Z(n11080) );
  NANDN U26843 ( .A(n29829), .B(n11080), .Z(n11081) );
  NAND U26844 ( .A(n29840), .B(n11081), .Z(n11082) );
  NANDN U26845 ( .A(x[359]), .B(y[359]), .Z(n28425) );
  NANDN U26846 ( .A(n11082), .B(n28425), .Z(n11083) );
  AND U26847 ( .A(n11084), .B(n11083), .Z(n11086) );
  NANDN U26848 ( .A(x[361]), .B(y[361]), .Z(n29839) );
  NANDN U26849 ( .A(x[362]), .B(y[362]), .Z(n29849) );
  AND U26850 ( .A(n29839), .B(n29849), .Z(n11085) );
  NANDN U26851 ( .A(n11086), .B(n11085), .Z(n11087) );
  ANDN U26852 ( .B(x[363]), .A(y[363]), .Z(n29852) );
  ANDN U26853 ( .B(n11087), .A(n29852), .Z(n11088) );
  NANDN U26854 ( .A(n29842), .B(n11088), .Z(n11089) );
  NANDN U26855 ( .A(x[363]), .B(y[363]), .Z(n29847) );
  AND U26856 ( .A(n11089), .B(n29847), .Z(n11090) );
  NANDN U26857 ( .A(n29851), .B(n11090), .Z(n11091) );
  ANDN U26858 ( .B(x[365]), .A(y[365]), .Z(n29856) );
  ANDN U26859 ( .B(n11091), .A(n29856), .Z(n11092) );
  NAND U26860 ( .A(n11093), .B(n11092), .Z(n11094) );
  NAND U26861 ( .A(n29862), .B(n11094), .Z(n11095) );
  NANDN U26862 ( .A(x[365]), .B(y[365]), .Z(n28422) );
  NANDN U26863 ( .A(n11095), .B(n28422), .Z(n11096) );
  AND U26864 ( .A(n11097), .B(n11096), .Z(n11099) );
  NANDN U26865 ( .A(x[367]), .B(y[367]), .Z(n29861) );
  NANDN U26866 ( .A(x[368]), .B(y[368]), .Z(n29868) );
  AND U26867 ( .A(n29861), .B(n29868), .Z(n11098) );
  NANDN U26868 ( .A(n11099), .B(n11098), .Z(n11100) );
  ANDN U26869 ( .B(x[369]), .A(y[369]), .Z(n29874) );
  ANDN U26870 ( .B(n11100), .A(n29874), .Z(n11101) );
  NANDN U26871 ( .A(n29864), .B(n11101), .Z(n11102) );
  NANDN U26872 ( .A(x[370]), .B(y[370]), .Z(n28420) );
  AND U26873 ( .A(n11102), .B(n28420), .Z(n11103) );
  NAND U26874 ( .A(n29869), .B(n11103), .Z(n11104) );
  ANDN U26875 ( .B(x[371]), .A(y[371]), .Z(n29878) );
  ANDN U26876 ( .B(n11104), .A(n29878), .Z(n11105) );
  NANDN U26877 ( .A(n29873), .B(n11105), .Z(n11106) );
  NAND U26878 ( .A(n29884), .B(n11106), .Z(n11107) );
  NANDN U26879 ( .A(x[371]), .B(y[371]), .Z(n28421) );
  NANDN U26880 ( .A(n11107), .B(n28421), .Z(n11108) );
  AND U26881 ( .A(n11109), .B(n11108), .Z(n11111) );
  NANDN U26882 ( .A(x[373]), .B(y[373]), .Z(n29883) );
  NANDN U26883 ( .A(x[374]), .B(y[374]), .Z(n29890) );
  AND U26884 ( .A(n29883), .B(n29890), .Z(n11110) );
  NANDN U26885 ( .A(n11111), .B(n11110), .Z(n11112) );
  ANDN U26886 ( .B(x[375]), .A(y[375]), .Z(n29896) );
  ANDN U26887 ( .B(n11112), .A(n29896), .Z(n11113) );
  NANDN U26888 ( .A(n29886), .B(n11113), .Z(n11114) );
  NANDN U26889 ( .A(x[376]), .B(y[376]), .Z(n28418) );
  AND U26890 ( .A(n11114), .B(n28418), .Z(n11115) );
  NAND U26891 ( .A(n29891), .B(n11115), .Z(n11116) );
  ANDN U26892 ( .B(x[377]), .A(y[377]), .Z(n29900) );
  ANDN U26893 ( .B(n11116), .A(n29900), .Z(n11117) );
  NANDN U26894 ( .A(n29895), .B(n11117), .Z(n11118) );
  NAND U26895 ( .A(n29906), .B(n11118), .Z(n11119) );
  NANDN U26896 ( .A(x[377]), .B(y[377]), .Z(n28419) );
  NANDN U26897 ( .A(n11119), .B(n28419), .Z(n11120) );
  AND U26898 ( .A(n11121), .B(n11120), .Z(n11123) );
  NANDN U26899 ( .A(x[379]), .B(y[379]), .Z(n29905) );
  NANDN U26900 ( .A(x[380]), .B(y[380]), .Z(n29912) );
  AND U26901 ( .A(n29905), .B(n29912), .Z(n11122) );
  NANDN U26902 ( .A(n11123), .B(n11122), .Z(n11124) );
  ANDN U26903 ( .B(x[381]), .A(y[381]), .Z(n29918) );
  ANDN U26904 ( .B(n11124), .A(n29918), .Z(n11125) );
  NANDN U26905 ( .A(n29908), .B(n11125), .Z(n11126) );
  NANDN U26906 ( .A(x[382]), .B(y[382]), .Z(n28416) );
  AND U26907 ( .A(n11126), .B(n28416), .Z(n11127) );
  NAND U26908 ( .A(n29913), .B(n11127), .Z(n11128) );
  ANDN U26909 ( .B(x[383]), .A(y[383]), .Z(n29922) );
  ANDN U26910 ( .B(n11128), .A(n29922), .Z(n11129) );
  NANDN U26911 ( .A(n29917), .B(n11129), .Z(n11130) );
  NAND U26912 ( .A(n29928), .B(n11130), .Z(n11131) );
  NANDN U26913 ( .A(x[383]), .B(y[383]), .Z(n28417) );
  NANDN U26914 ( .A(n11131), .B(n28417), .Z(n11132) );
  AND U26915 ( .A(n11133), .B(n11132), .Z(n11135) );
  NANDN U26916 ( .A(x[385]), .B(y[385]), .Z(n29927) );
  NANDN U26917 ( .A(x[386]), .B(y[386]), .Z(n29934) );
  AND U26918 ( .A(n29927), .B(n29934), .Z(n11134) );
  NANDN U26919 ( .A(n11135), .B(n11134), .Z(n11136) );
  ANDN U26920 ( .B(x[387]), .A(y[387]), .Z(n29940) );
  ANDN U26921 ( .B(n11136), .A(n29940), .Z(n11137) );
  NANDN U26922 ( .A(n29930), .B(n11137), .Z(n11138) );
  NANDN U26923 ( .A(x[388]), .B(y[388]), .Z(n28414) );
  AND U26924 ( .A(n11138), .B(n28414), .Z(n11139) );
  NAND U26925 ( .A(n29935), .B(n11139), .Z(n11140) );
  ANDN U26926 ( .B(x[389]), .A(y[389]), .Z(n29944) );
  ANDN U26927 ( .B(n11140), .A(n29944), .Z(n11141) );
  NANDN U26928 ( .A(n29939), .B(n11141), .Z(n11142) );
  NAND U26929 ( .A(n29950), .B(n11142), .Z(n11143) );
  NANDN U26930 ( .A(x[389]), .B(y[389]), .Z(n28415) );
  NANDN U26931 ( .A(n11143), .B(n28415), .Z(n11144) );
  AND U26932 ( .A(n11145), .B(n11144), .Z(n11147) );
  NANDN U26933 ( .A(x[391]), .B(y[391]), .Z(n29949) );
  NANDN U26934 ( .A(x[392]), .B(y[392]), .Z(n29956) );
  AND U26935 ( .A(n29949), .B(n29956), .Z(n11146) );
  NANDN U26936 ( .A(n11147), .B(n11146), .Z(n11148) );
  ANDN U26937 ( .B(x[393]), .A(y[393]), .Z(n29962) );
  ANDN U26938 ( .B(n11148), .A(n29962), .Z(n11149) );
  NANDN U26939 ( .A(n29952), .B(n11149), .Z(n11150) );
  NANDN U26940 ( .A(x[394]), .B(y[394]), .Z(n28412) );
  AND U26941 ( .A(n11150), .B(n28412), .Z(n11151) );
  NAND U26942 ( .A(n29957), .B(n11151), .Z(n11152) );
  ANDN U26943 ( .B(x[395]), .A(y[395]), .Z(n29966) );
  ANDN U26944 ( .B(n11152), .A(n29966), .Z(n11153) );
  NANDN U26945 ( .A(n29961), .B(n11153), .Z(n11154) );
  NAND U26946 ( .A(n29972), .B(n11154), .Z(n11155) );
  NANDN U26947 ( .A(x[395]), .B(y[395]), .Z(n28413) );
  NANDN U26948 ( .A(n11155), .B(n28413), .Z(n11156) );
  AND U26949 ( .A(n11157), .B(n11156), .Z(n11159) );
  NANDN U26950 ( .A(x[397]), .B(y[397]), .Z(n29971) );
  NANDN U26951 ( .A(x[398]), .B(y[398]), .Z(n29978) );
  AND U26952 ( .A(n29971), .B(n29978), .Z(n11158) );
  NANDN U26953 ( .A(n11159), .B(n11158), .Z(n11160) );
  ANDN U26954 ( .B(x[399]), .A(y[399]), .Z(n29984) );
  ANDN U26955 ( .B(n11160), .A(n29984), .Z(n11161) );
  NANDN U26956 ( .A(n29974), .B(n11161), .Z(n11162) );
  NANDN U26957 ( .A(x[400]), .B(y[400]), .Z(n28410) );
  AND U26958 ( .A(n11162), .B(n28410), .Z(n11163) );
  NAND U26959 ( .A(n29979), .B(n11163), .Z(n11164) );
  ANDN U26960 ( .B(x[401]), .A(y[401]), .Z(n29988) );
  ANDN U26961 ( .B(n11164), .A(n29988), .Z(n11165) );
  NANDN U26962 ( .A(n29983), .B(n11165), .Z(n11166) );
  NAND U26963 ( .A(n29994), .B(n11166), .Z(n11167) );
  NANDN U26964 ( .A(x[401]), .B(y[401]), .Z(n28411) );
  NANDN U26965 ( .A(n11167), .B(n28411), .Z(n11168) );
  AND U26966 ( .A(n11169), .B(n11168), .Z(n11171) );
  NANDN U26967 ( .A(x[403]), .B(y[403]), .Z(n29993) );
  NANDN U26968 ( .A(x[404]), .B(y[404]), .Z(n30000) );
  AND U26969 ( .A(n29993), .B(n30000), .Z(n11170) );
  NANDN U26970 ( .A(n11171), .B(n11170), .Z(n11172) );
  ANDN U26971 ( .B(x[405]), .A(y[405]), .Z(n30006) );
  ANDN U26972 ( .B(n11172), .A(n30006), .Z(n11173) );
  NANDN U26973 ( .A(n29996), .B(n11173), .Z(n11174) );
  NANDN U26974 ( .A(x[406]), .B(y[406]), .Z(n28408) );
  AND U26975 ( .A(n11174), .B(n28408), .Z(n11175) );
  NAND U26976 ( .A(n30001), .B(n11175), .Z(n11176) );
  ANDN U26977 ( .B(x[407]), .A(y[407]), .Z(n30010) );
  ANDN U26978 ( .B(n11176), .A(n30010), .Z(n11177) );
  NANDN U26979 ( .A(n30005), .B(n11177), .Z(n11178) );
  NAND U26980 ( .A(n30016), .B(n11178), .Z(n11179) );
  NANDN U26981 ( .A(x[407]), .B(y[407]), .Z(n28409) );
  NANDN U26982 ( .A(n11179), .B(n28409), .Z(n11180) );
  AND U26983 ( .A(n11181), .B(n11180), .Z(n11183) );
  NANDN U26984 ( .A(x[409]), .B(y[409]), .Z(n30015) );
  NANDN U26985 ( .A(x[410]), .B(y[410]), .Z(n30022) );
  AND U26986 ( .A(n30015), .B(n30022), .Z(n11182) );
  NANDN U26987 ( .A(n11183), .B(n11182), .Z(n11184) );
  ANDN U26988 ( .B(x[411]), .A(y[411]), .Z(n30028) );
  ANDN U26989 ( .B(n11184), .A(n30028), .Z(n11185) );
  NANDN U26990 ( .A(n30018), .B(n11185), .Z(n11186) );
  NANDN U26991 ( .A(x[412]), .B(y[412]), .Z(n28406) );
  AND U26992 ( .A(n11186), .B(n28406), .Z(n11187) );
  NAND U26993 ( .A(n30023), .B(n11187), .Z(n11188) );
  ANDN U26994 ( .B(x[413]), .A(y[413]), .Z(n30032) );
  ANDN U26995 ( .B(n11188), .A(n30032), .Z(n11189) );
  NANDN U26996 ( .A(n30027), .B(n11189), .Z(n11190) );
  NAND U26997 ( .A(n30038), .B(n11190), .Z(n11191) );
  NANDN U26998 ( .A(x[413]), .B(y[413]), .Z(n28407) );
  NANDN U26999 ( .A(n11191), .B(n28407), .Z(n11192) );
  AND U27000 ( .A(n11193), .B(n11192), .Z(n11195) );
  NANDN U27001 ( .A(x[415]), .B(y[415]), .Z(n30037) );
  NANDN U27002 ( .A(x[416]), .B(y[416]), .Z(n30044) );
  AND U27003 ( .A(n30037), .B(n30044), .Z(n11194) );
  NANDN U27004 ( .A(n11195), .B(n11194), .Z(n11196) );
  ANDN U27005 ( .B(x[417]), .A(y[417]), .Z(n30050) );
  ANDN U27006 ( .B(n11196), .A(n30050), .Z(n11197) );
  NANDN U27007 ( .A(n30040), .B(n11197), .Z(n11198) );
  NANDN U27008 ( .A(x[418]), .B(y[418]), .Z(n28404) );
  AND U27009 ( .A(n11198), .B(n28404), .Z(n11199) );
  NAND U27010 ( .A(n30045), .B(n11199), .Z(n11200) );
  ANDN U27011 ( .B(x[419]), .A(y[419]), .Z(n30054) );
  ANDN U27012 ( .B(n11200), .A(n30054), .Z(n11201) );
  NANDN U27013 ( .A(n30049), .B(n11201), .Z(n11202) );
  NAND U27014 ( .A(n30060), .B(n11202), .Z(n11203) );
  NANDN U27015 ( .A(x[419]), .B(y[419]), .Z(n28405) );
  NANDN U27016 ( .A(n11203), .B(n28405), .Z(n11204) );
  AND U27017 ( .A(n11205), .B(n11204), .Z(n11207) );
  NANDN U27018 ( .A(x[421]), .B(y[421]), .Z(n30059) );
  NANDN U27019 ( .A(x[422]), .B(y[422]), .Z(n30066) );
  AND U27020 ( .A(n30059), .B(n30066), .Z(n11206) );
  NANDN U27021 ( .A(n11207), .B(n11206), .Z(n11208) );
  ANDN U27022 ( .B(x[423]), .A(y[423]), .Z(n30072) );
  ANDN U27023 ( .B(n11208), .A(n30072), .Z(n11209) );
  NANDN U27024 ( .A(n30062), .B(n11209), .Z(n11210) );
  NANDN U27025 ( .A(x[424]), .B(y[424]), .Z(n28402) );
  AND U27026 ( .A(n11210), .B(n28402), .Z(n11211) );
  NAND U27027 ( .A(n30067), .B(n11211), .Z(n11212) );
  ANDN U27028 ( .B(x[425]), .A(y[425]), .Z(n30076) );
  ANDN U27029 ( .B(n11212), .A(n30076), .Z(n11213) );
  NANDN U27030 ( .A(n30071), .B(n11213), .Z(n11214) );
  NAND U27031 ( .A(n30082), .B(n11214), .Z(n11215) );
  NANDN U27032 ( .A(x[425]), .B(y[425]), .Z(n28403) );
  NANDN U27033 ( .A(n11215), .B(n28403), .Z(n11216) );
  AND U27034 ( .A(n11217), .B(n11216), .Z(n11219) );
  NANDN U27035 ( .A(x[427]), .B(y[427]), .Z(n30081) );
  NANDN U27036 ( .A(x[428]), .B(y[428]), .Z(n30088) );
  AND U27037 ( .A(n30081), .B(n30088), .Z(n11218) );
  NANDN U27038 ( .A(n11219), .B(n11218), .Z(n11220) );
  ANDN U27039 ( .B(x[429]), .A(y[429]), .Z(n30094) );
  ANDN U27040 ( .B(n11220), .A(n30094), .Z(n11221) );
  NANDN U27041 ( .A(n30084), .B(n11221), .Z(n11222) );
  NANDN U27042 ( .A(x[430]), .B(y[430]), .Z(n28400) );
  AND U27043 ( .A(n11222), .B(n28400), .Z(n11223) );
  NAND U27044 ( .A(n30089), .B(n11223), .Z(n11224) );
  ANDN U27045 ( .B(x[430]), .A(y[430]), .Z(n30093) );
  ANDN U27046 ( .B(n11224), .A(n30093), .Z(n11225) );
  NANDN U27047 ( .A(n30101), .B(n11225), .Z(n11226) );
  NANDN U27048 ( .A(n30099), .B(n11226), .Z(n11227) );
  NANDN U27049 ( .A(x[431]), .B(y[431]), .Z(n28401) );
  NANDN U27050 ( .A(n11227), .B(n28401), .Z(n11228) );
  AND U27051 ( .A(n11229), .B(n11228), .Z(n11231) );
  NANDN U27052 ( .A(x[433]), .B(y[433]), .Z(n30103) );
  NANDN U27053 ( .A(x[434]), .B(y[434]), .Z(n30110) );
  AND U27054 ( .A(n30103), .B(n30110), .Z(n11230) );
  NANDN U27055 ( .A(n11231), .B(n11230), .Z(n11232) );
  ANDN U27056 ( .B(x[435]), .A(y[435]), .Z(n30116) );
  ANDN U27057 ( .B(n11232), .A(n30116), .Z(n11233) );
  NANDN U27058 ( .A(n30106), .B(n11233), .Z(n11234) );
  NANDN U27059 ( .A(x[436]), .B(y[436]), .Z(n28398) );
  AND U27060 ( .A(n11234), .B(n28398), .Z(n11235) );
  NAND U27061 ( .A(n30111), .B(n11235), .Z(n11236) );
  ANDN U27062 ( .B(x[437]), .A(y[437]), .Z(n30120) );
  ANDN U27063 ( .B(n11236), .A(n30120), .Z(n11237) );
  NANDN U27064 ( .A(n30115), .B(n11237), .Z(n11238) );
  NAND U27065 ( .A(n30126), .B(n11238), .Z(n11239) );
  NANDN U27066 ( .A(x[437]), .B(y[437]), .Z(n28399) );
  NANDN U27067 ( .A(n11239), .B(n28399), .Z(n11240) );
  AND U27068 ( .A(n11241), .B(n11240), .Z(n11243) );
  NANDN U27069 ( .A(x[439]), .B(y[439]), .Z(n30125) );
  NANDN U27070 ( .A(x[440]), .B(y[440]), .Z(n30132) );
  AND U27071 ( .A(n30125), .B(n30132), .Z(n11242) );
  NANDN U27072 ( .A(n11243), .B(n11242), .Z(n11244) );
  ANDN U27073 ( .B(x[441]), .A(y[441]), .Z(n30138) );
  ANDN U27074 ( .B(n11244), .A(n30138), .Z(n11245) );
  NANDN U27075 ( .A(n30128), .B(n11245), .Z(n11246) );
  NANDN U27076 ( .A(x[442]), .B(y[442]), .Z(n28396) );
  AND U27077 ( .A(n11246), .B(n28396), .Z(n11247) );
  NAND U27078 ( .A(n30133), .B(n11247), .Z(n11248) );
  ANDN U27079 ( .B(x[443]), .A(y[443]), .Z(n30142) );
  ANDN U27080 ( .B(n11248), .A(n30142), .Z(n11249) );
  NANDN U27081 ( .A(n30137), .B(n11249), .Z(n11250) );
  NAND U27082 ( .A(n30148), .B(n11250), .Z(n11251) );
  NANDN U27083 ( .A(x[443]), .B(y[443]), .Z(n28397) );
  NANDN U27084 ( .A(n11251), .B(n28397), .Z(n11252) );
  AND U27085 ( .A(n11253), .B(n11252), .Z(n11255) );
  NANDN U27086 ( .A(x[445]), .B(y[445]), .Z(n30147) );
  NANDN U27087 ( .A(x[446]), .B(y[446]), .Z(n30154) );
  AND U27088 ( .A(n30147), .B(n30154), .Z(n11254) );
  NANDN U27089 ( .A(n11255), .B(n11254), .Z(n11256) );
  ANDN U27090 ( .B(x[447]), .A(y[447]), .Z(n30160) );
  ANDN U27091 ( .B(n11256), .A(n30160), .Z(n11257) );
  NANDN U27092 ( .A(n30150), .B(n11257), .Z(n11258) );
  NANDN U27093 ( .A(x[448]), .B(y[448]), .Z(n28394) );
  AND U27094 ( .A(n11258), .B(n28394), .Z(n11259) );
  NAND U27095 ( .A(n30155), .B(n11259), .Z(n11260) );
  ANDN U27096 ( .B(x[449]), .A(y[449]), .Z(n30164) );
  ANDN U27097 ( .B(n11260), .A(n30164), .Z(n11261) );
  NANDN U27098 ( .A(n30159), .B(n11261), .Z(n11262) );
  NAND U27099 ( .A(n30170), .B(n11262), .Z(n11263) );
  NANDN U27100 ( .A(x[449]), .B(y[449]), .Z(n28395) );
  NANDN U27101 ( .A(n11263), .B(n28395), .Z(n11264) );
  AND U27102 ( .A(n11265), .B(n11264), .Z(n11267) );
  NANDN U27103 ( .A(x[451]), .B(y[451]), .Z(n30169) );
  NANDN U27104 ( .A(x[452]), .B(y[452]), .Z(n30176) );
  AND U27105 ( .A(n30169), .B(n30176), .Z(n11266) );
  NANDN U27106 ( .A(n11267), .B(n11266), .Z(n11268) );
  ANDN U27107 ( .B(x[453]), .A(y[453]), .Z(n30182) );
  ANDN U27108 ( .B(n11268), .A(n30182), .Z(n11269) );
  NANDN U27109 ( .A(n30172), .B(n11269), .Z(n11270) );
  NANDN U27110 ( .A(x[454]), .B(y[454]), .Z(n28392) );
  AND U27111 ( .A(n11270), .B(n28392), .Z(n11271) );
  NAND U27112 ( .A(n30177), .B(n11271), .Z(n11272) );
  ANDN U27113 ( .B(x[455]), .A(y[455]), .Z(n30186) );
  ANDN U27114 ( .B(n11272), .A(n30186), .Z(n11273) );
  NANDN U27115 ( .A(n30181), .B(n11273), .Z(n11274) );
  NAND U27116 ( .A(n30192), .B(n11274), .Z(n11275) );
  NANDN U27117 ( .A(x[455]), .B(y[455]), .Z(n28393) );
  NANDN U27118 ( .A(n11275), .B(n28393), .Z(n11276) );
  AND U27119 ( .A(n11277), .B(n11276), .Z(n11279) );
  NANDN U27120 ( .A(x[457]), .B(y[457]), .Z(n30191) );
  NANDN U27121 ( .A(x[458]), .B(y[458]), .Z(n30198) );
  AND U27122 ( .A(n30191), .B(n30198), .Z(n11278) );
  NANDN U27123 ( .A(n11279), .B(n11278), .Z(n11280) );
  ANDN U27124 ( .B(x[459]), .A(y[459]), .Z(n30204) );
  ANDN U27125 ( .B(n11280), .A(n30204), .Z(n11281) );
  NANDN U27126 ( .A(n30194), .B(n11281), .Z(n11282) );
  NANDN U27127 ( .A(x[460]), .B(y[460]), .Z(n28390) );
  AND U27128 ( .A(n11282), .B(n28390), .Z(n11283) );
  NAND U27129 ( .A(n30199), .B(n11283), .Z(n11284) );
  ANDN U27130 ( .B(x[461]), .A(y[461]), .Z(n30208) );
  ANDN U27131 ( .B(n11284), .A(n30208), .Z(n11285) );
  NANDN U27132 ( .A(n30203), .B(n11285), .Z(n11286) );
  NAND U27133 ( .A(n30214), .B(n11286), .Z(n11287) );
  NANDN U27134 ( .A(x[461]), .B(y[461]), .Z(n28391) );
  NANDN U27135 ( .A(n11287), .B(n28391), .Z(n11288) );
  AND U27136 ( .A(n11289), .B(n11288), .Z(n11291) );
  NANDN U27137 ( .A(x[463]), .B(y[463]), .Z(n30213) );
  NANDN U27138 ( .A(x[464]), .B(y[464]), .Z(n30220) );
  AND U27139 ( .A(n30213), .B(n30220), .Z(n11290) );
  NANDN U27140 ( .A(n11291), .B(n11290), .Z(n11292) );
  ANDN U27141 ( .B(x[465]), .A(y[465]), .Z(n30226) );
  ANDN U27142 ( .B(n11292), .A(n30226), .Z(n11293) );
  NANDN U27143 ( .A(n30216), .B(n11293), .Z(n11294) );
  NANDN U27144 ( .A(x[466]), .B(y[466]), .Z(n28388) );
  AND U27145 ( .A(n11294), .B(n28388), .Z(n11295) );
  NAND U27146 ( .A(n30221), .B(n11295), .Z(n11296) );
  ANDN U27147 ( .B(x[467]), .A(y[467]), .Z(n30230) );
  ANDN U27148 ( .B(n11296), .A(n30230), .Z(n11297) );
  NANDN U27149 ( .A(n30225), .B(n11297), .Z(n11298) );
  NAND U27150 ( .A(n30236), .B(n11298), .Z(n11299) );
  NANDN U27151 ( .A(x[467]), .B(y[467]), .Z(n28389) );
  NANDN U27152 ( .A(n11299), .B(n28389), .Z(n11300) );
  AND U27153 ( .A(n11301), .B(n11300), .Z(n11303) );
  NANDN U27154 ( .A(x[469]), .B(y[469]), .Z(n30235) );
  NANDN U27155 ( .A(x[470]), .B(y[470]), .Z(n30242) );
  AND U27156 ( .A(n30235), .B(n30242), .Z(n11302) );
  NANDN U27157 ( .A(n11303), .B(n11302), .Z(n11304) );
  ANDN U27158 ( .B(x[471]), .A(y[471]), .Z(n30248) );
  ANDN U27159 ( .B(n11304), .A(n30248), .Z(n11305) );
  NANDN U27160 ( .A(n30238), .B(n11305), .Z(n11306) );
  NANDN U27161 ( .A(x[472]), .B(y[472]), .Z(n28386) );
  AND U27162 ( .A(n11306), .B(n28386), .Z(n11307) );
  NAND U27163 ( .A(n30243), .B(n11307), .Z(n11308) );
  ANDN U27164 ( .B(x[473]), .A(y[473]), .Z(n30252) );
  ANDN U27165 ( .B(n11308), .A(n30252), .Z(n11309) );
  NANDN U27166 ( .A(n30247), .B(n11309), .Z(n11310) );
  NAND U27167 ( .A(n30258), .B(n11310), .Z(n11311) );
  NANDN U27168 ( .A(x[473]), .B(y[473]), .Z(n28387) );
  NANDN U27169 ( .A(n11311), .B(n28387), .Z(n11312) );
  AND U27170 ( .A(n11313), .B(n11312), .Z(n11315) );
  NANDN U27171 ( .A(x[475]), .B(y[475]), .Z(n30257) );
  NANDN U27172 ( .A(x[476]), .B(y[476]), .Z(n30264) );
  AND U27173 ( .A(n30257), .B(n30264), .Z(n11314) );
  NANDN U27174 ( .A(n11315), .B(n11314), .Z(n11316) );
  ANDN U27175 ( .B(x[477]), .A(y[477]), .Z(n30270) );
  ANDN U27176 ( .B(n11316), .A(n30270), .Z(n11317) );
  NANDN U27177 ( .A(n30260), .B(n11317), .Z(n11318) );
  NANDN U27178 ( .A(x[478]), .B(y[478]), .Z(n28384) );
  AND U27179 ( .A(n11318), .B(n28384), .Z(n11319) );
  NAND U27180 ( .A(n30265), .B(n11319), .Z(n11320) );
  ANDN U27181 ( .B(x[479]), .A(y[479]), .Z(n30274) );
  ANDN U27182 ( .B(n11320), .A(n30274), .Z(n11321) );
  NANDN U27183 ( .A(n30269), .B(n11321), .Z(n11322) );
  NAND U27184 ( .A(n30280), .B(n11322), .Z(n11323) );
  NANDN U27185 ( .A(x[479]), .B(y[479]), .Z(n28385) );
  NANDN U27186 ( .A(n11323), .B(n28385), .Z(n11324) );
  AND U27187 ( .A(n11325), .B(n11324), .Z(n11327) );
  NANDN U27188 ( .A(x[481]), .B(y[481]), .Z(n30279) );
  NANDN U27189 ( .A(x[482]), .B(y[482]), .Z(n30286) );
  AND U27190 ( .A(n30279), .B(n30286), .Z(n11326) );
  NANDN U27191 ( .A(n11327), .B(n11326), .Z(n11328) );
  ANDN U27192 ( .B(x[483]), .A(y[483]), .Z(n30292) );
  ANDN U27193 ( .B(n11328), .A(n30292), .Z(n11329) );
  NANDN U27194 ( .A(n30282), .B(n11329), .Z(n11330) );
  NANDN U27195 ( .A(x[484]), .B(y[484]), .Z(n28382) );
  AND U27196 ( .A(n11330), .B(n28382), .Z(n11331) );
  NAND U27197 ( .A(n30287), .B(n11331), .Z(n11332) );
  ANDN U27198 ( .B(x[485]), .A(y[485]), .Z(n30296) );
  ANDN U27199 ( .B(n11332), .A(n30296), .Z(n11333) );
  NANDN U27200 ( .A(n30291), .B(n11333), .Z(n11334) );
  NAND U27201 ( .A(n30302), .B(n11334), .Z(n11335) );
  NANDN U27202 ( .A(x[485]), .B(y[485]), .Z(n28383) );
  NANDN U27203 ( .A(n11335), .B(n28383), .Z(n11336) );
  AND U27204 ( .A(n11337), .B(n11336), .Z(n11339) );
  NANDN U27205 ( .A(x[487]), .B(y[487]), .Z(n30301) );
  NANDN U27206 ( .A(x[488]), .B(y[488]), .Z(n30308) );
  AND U27207 ( .A(n30301), .B(n30308), .Z(n11338) );
  NANDN U27208 ( .A(n11339), .B(n11338), .Z(n11340) );
  ANDN U27209 ( .B(x[489]), .A(y[489]), .Z(n30314) );
  ANDN U27210 ( .B(n11340), .A(n30314), .Z(n11341) );
  NANDN U27211 ( .A(n30304), .B(n11341), .Z(n11342) );
  NANDN U27212 ( .A(x[490]), .B(y[490]), .Z(n28380) );
  AND U27213 ( .A(n11342), .B(n28380), .Z(n11343) );
  NAND U27214 ( .A(n30309), .B(n11343), .Z(n11344) );
  ANDN U27215 ( .B(x[491]), .A(y[491]), .Z(n30318) );
  ANDN U27216 ( .B(n11344), .A(n30318), .Z(n11345) );
  NANDN U27217 ( .A(n30313), .B(n11345), .Z(n11346) );
  NAND U27218 ( .A(n30324), .B(n11346), .Z(n11347) );
  NANDN U27219 ( .A(x[491]), .B(y[491]), .Z(n28381) );
  NANDN U27220 ( .A(n11347), .B(n28381), .Z(n11348) );
  AND U27221 ( .A(n11349), .B(n11348), .Z(n11351) );
  NANDN U27222 ( .A(x[493]), .B(y[493]), .Z(n30323) );
  NANDN U27223 ( .A(x[494]), .B(y[494]), .Z(n30330) );
  AND U27224 ( .A(n30323), .B(n30330), .Z(n11350) );
  NANDN U27225 ( .A(n11351), .B(n11350), .Z(n11352) );
  ANDN U27226 ( .B(x[495]), .A(y[495]), .Z(n30336) );
  ANDN U27227 ( .B(n11352), .A(n30336), .Z(n11353) );
  NANDN U27228 ( .A(n30326), .B(n11353), .Z(n11354) );
  NANDN U27229 ( .A(x[496]), .B(y[496]), .Z(n28378) );
  AND U27230 ( .A(n11354), .B(n28378), .Z(n11355) );
  NAND U27231 ( .A(n30331), .B(n11355), .Z(n11356) );
  ANDN U27232 ( .B(x[497]), .A(y[497]), .Z(n30340) );
  ANDN U27233 ( .B(n11356), .A(n30340), .Z(n11357) );
  NANDN U27234 ( .A(n30335), .B(n11357), .Z(n11358) );
  NAND U27235 ( .A(n30346), .B(n11358), .Z(n11359) );
  NANDN U27236 ( .A(x[497]), .B(y[497]), .Z(n28379) );
  NANDN U27237 ( .A(n11359), .B(n28379), .Z(n11360) );
  AND U27238 ( .A(n11361), .B(n11360), .Z(n11363) );
  NANDN U27239 ( .A(x[499]), .B(y[499]), .Z(n30345) );
  NANDN U27240 ( .A(x[500]), .B(y[500]), .Z(n30352) );
  AND U27241 ( .A(n30345), .B(n30352), .Z(n11362) );
  NANDN U27242 ( .A(n11363), .B(n11362), .Z(n11364) );
  ANDN U27243 ( .B(x[501]), .A(y[501]), .Z(n30358) );
  ANDN U27244 ( .B(n11364), .A(n30358), .Z(n11365) );
  NANDN U27245 ( .A(n30348), .B(n11365), .Z(n11366) );
  NANDN U27246 ( .A(x[502]), .B(y[502]), .Z(n28376) );
  AND U27247 ( .A(n11366), .B(n28376), .Z(n11367) );
  NAND U27248 ( .A(n30353), .B(n11367), .Z(n11368) );
  ANDN U27249 ( .B(x[503]), .A(y[503]), .Z(n30362) );
  ANDN U27250 ( .B(n11368), .A(n30362), .Z(n11369) );
  NANDN U27251 ( .A(n30357), .B(n11369), .Z(n11370) );
  NAND U27252 ( .A(n30368), .B(n11370), .Z(n11371) );
  NANDN U27253 ( .A(x[503]), .B(y[503]), .Z(n28377) );
  NANDN U27254 ( .A(n11371), .B(n28377), .Z(n11372) );
  AND U27255 ( .A(n11373), .B(n11372), .Z(n11375) );
  NANDN U27256 ( .A(x[505]), .B(y[505]), .Z(n30367) );
  NANDN U27257 ( .A(x[506]), .B(y[506]), .Z(n30374) );
  AND U27258 ( .A(n30367), .B(n30374), .Z(n11374) );
  NANDN U27259 ( .A(n11375), .B(n11374), .Z(n11376) );
  ANDN U27260 ( .B(x[507]), .A(y[507]), .Z(n30380) );
  ANDN U27261 ( .B(n11376), .A(n30380), .Z(n11377) );
  NANDN U27262 ( .A(n30370), .B(n11377), .Z(n11378) );
  NANDN U27263 ( .A(x[508]), .B(y[508]), .Z(n28374) );
  AND U27264 ( .A(n11378), .B(n28374), .Z(n11379) );
  NAND U27265 ( .A(n30375), .B(n11379), .Z(n11380) );
  ANDN U27266 ( .B(x[509]), .A(y[509]), .Z(n30384) );
  ANDN U27267 ( .B(n11380), .A(n30384), .Z(n11381) );
  NANDN U27268 ( .A(n30379), .B(n11381), .Z(n11382) );
  NAND U27269 ( .A(n30390), .B(n11382), .Z(n11383) );
  NANDN U27270 ( .A(x[509]), .B(y[509]), .Z(n28375) );
  NANDN U27271 ( .A(n11383), .B(n28375), .Z(n11384) );
  AND U27272 ( .A(n11385), .B(n11384), .Z(n11387) );
  NANDN U27273 ( .A(x[511]), .B(y[511]), .Z(n30389) );
  NANDN U27274 ( .A(x[512]), .B(y[512]), .Z(n30396) );
  AND U27275 ( .A(n30389), .B(n30396), .Z(n11386) );
  NANDN U27276 ( .A(n11387), .B(n11386), .Z(n11388) );
  ANDN U27277 ( .B(x[513]), .A(y[513]), .Z(n30402) );
  ANDN U27278 ( .B(n11388), .A(n30402), .Z(n11389) );
  NANDN U27279 ( .A(n30392), .B(n11389), .Z(n11390) );
  NANDN U27280 ( .A(x[514]), .B(y[514]), .Z(n28372) );
  AND U27281 ( .A(n11390), .B(n28372), .Z(n11391) );
  NAND U27282 ( .A(n30397), .B(n11391), .Z(n11392) );
  ANDN U27283 ( .B(x[515]), .A(y[515]), .Z(n30406) );
  ANDN U27284 ( .B(n11392), .A(n30406), .Z(n11393) );
  NANDN U27285 ( .A(n30401), .B(n11393), .Z(n11394) );
  NAND U27286 ( .A(n30412), .B(n11394), .Z(n11395) );
  NANDN U27287 ( .A(x[515]), .B(y[515]), .Z(n28373) );
  NANDN U27288 ( .A(n11395), .B(n28373), .Z(n11396) );
  AND U27289 ( .A(n11397), .B(n11396), .Z(n11399) );
  NANDN U27290 ( .A(x[517]), .B(y[517]), .Z(n30411) );
  NANDN U27291 ( .A(x[518]), .B(y[518]), .Z(n30418) );
  AND U27292 ( .A(n30411), .B(n30418), .Z(n11398) );
  NANDN U27293 ( .A(n11399), .B(n11398), .Z(n11400) );
  ANDN U27294 ( .B(x[519]), .A(y[519]), .Z(n30424) );
  ANDN U27295 ( .B(n11400), .A(n30424), .Z(n11401) );
  NANDN U27296 ( .A(n30414), .B(n11401), .Z(n11402) );
  NANDN U27297 ( .A(x[520]), .B(y[520]), .Z(n28370) );
  AND U27298 ( .A(n11402), .B(n28370), .Z(n11403) );
  NAND U27299 ( .A(n30419), .B(n11403), .Z(n11404) );
  ANDN U27300 ( .B(x[521]), .A(y[521]), .Z(n30428) );
  ANDN U27301 ( .B(n11404), .A(n30428), .Z(n11405) );
  NANDN U27302 ( .A(n30423), .B(n11405), .Z(n11406) );
  NAND U27303 ( .A(n30434), .B(n11406), .Z(n11407) );
  NANDN U27304 ( .A(x[521]), .B(y[521]), .Z(n28371) );
  NANDN U27305 ( .A(n11407), .B(n28371), .Z(n11408) );
  AND U27306 ( .A(n11409), .B(n11408), .Z(n11411) );
  NANDN U27307 ( .A(x[523]), .B(y[523]), .Z(n30433) );
  NANDN U27308 ( .A(x[524]), .B(y[524]), .Z(n30440) );
  AND U27309 ( .A(n30433), .B(n30440), .Z(n11410) );
  NANDN U27310 ( .A(n11411), .B(n11410), .Z(n11412) );
  ANDN U27311 ( .B(x[525]), .A(y[525]), .Z(n30445) );
  ANDN U27312 ( .B(n11412), .A(n30445), .Z(n11413) );
  NANDN U27313 ( .A(n30436), .B(n11413), .Z(n11415) );
  ANDN U27314 ( .B(y[526]), .A(x[526]), .Z(n11414) );
  ANDN U27315 ( .B(n11415), .A(n11414), .Z(n11416) );
  NAND U27316 ( .A(n30441), .B(n11416), .Z(n11417) );
  NAND U27317 ( .A(n11418), .B(n11417), .Z(n11419) );
  NAND U27318 ( .A(n30453), .B(n11419), .Z(n11422) );
  NANDN U27319 ( .A(y[529]), .B(x[529]), .Z(n11421) );
  NANDN U27320 ( .A(y[528]), .B(x[528]), .Z(n11420) );
  NAND U27321 ( .A(n11421), .B(n11420), .Z(n30455) );
  ANDN U27322 ( .B(n11422), .A(n30455), .Z(n11425) );
  NANDN U27323 ( .A(x[529]), .B(y[529]), .Z(n11424) );
  NANDN U27324 ( .A(x[530]), .B(y[530]), .Z(n11423) );
  AND U27325 ( .A(n11424), .B(n11423), .Z(n30457) );
  NANDN U27326 ( .A(n11425), .B(n30457), .Z(n11426) );
  NANDN U27327 ( .A(n30459), .B(n11426), .Z(n11427) );
  NAND U27328 ( .A(n30461), .B(n11427), .Z(n11428) );
  NANDN U27329 ( .A(n30463), .B(n11428), .Z(n11429) );
  NAND U27330 ( .A(n30465), .B(n11429), .Z(n11432) );
  NANDN U27331 ( .A(y[535]), .B(x[535]), .Z(n11431) );
  NANDN U27332 ( .A(y[534]), .B(x[534]), .Z(n11430) );
  NAND U27333 ( .A(n11431), .B(n11430), .Z(n30467) );
  ANDN U27334 ( .B(n11432), .A(n30467), .Z(n11435) );
  NANDN U27335 ( .A(x[535]), .B(y[535]), .Z(n11434) );
  NANDN U27336 ( .A(x[536]), .B(y[536]), .Z(n11433) );
  AND U27337 ( .A(n11434), .B(n11433), .Z(n30469) );
  NANDN U27338 ( .A(n11435), .B(n30469), .Z(n11436) );
  NANDN U27339 ( .A(n30471), .B(n11436), .Z(n11437) );
  NAND U27340 ( .A(n30476), .B(n11437), .Z(n11438) );
  NANDN U27341 ( .A(x[537]), .B(y[537]), .Z(n30473) );
  NANDN U27342 ( .A(n11438), .B(n30473), .Z(n11439) );
  AND U27343 ( .A(n11440), .B(n11439), .Z(n11442) );
  NANDN U27344 ( .A(x[539]), .B(y[539]), .Z(n30477) );
  NANDN U27345 ( .A(x[540]), .B(y[540]), .Z(n28368) );
  AND U27346 ( .A(n30477), .B(n28368), .Z(n11441) );
  NANDN U27347 ( .A(n11442), .B(n11441), .Z(n11443) );
  ANDN U27348 ( .B(x[541]), .A(y[541]), .Z(n30489) );
  ANDN U27349 ( .B(n11443), .A(n30489), .Z(n11444) );
  NANDN U27350 ( .A(n30481), .B(n11444), .Z(n11445) );
  NANDN U27351 ( .A(x[541]), .B(y[541]), .Z(n28369) );
  AND U27352 ( .A(n11445), .B(n28369), .Z(n11446) );
  NANDN U27353 ( .A(n30487), .B(n11446), .Z(n11447) );
  ANDN U27354 ( .B(x[543]), .A(y[543]), .Z(n30497) );
  ANDN U27355 ( .B(n11447), .A(n30497), .Z(n11448) );
  NAND U27356 ( .A(n11449), .B(n11448), .Z(n11450) );
  NAND U27357 ( .A(n30498), .B(n11450), .Z(n11451) );
  NANDN U27358 ( .A(x[543]), .B(y[543]), .Z(n30491) );
  NANDN U27359 ( .A(n11451), .B(n30491), .Z(n11452) );
  ANDN U27360 ( .B(x[545]), .A(y[545]), .Z(n30504) );
  ANDN U27361 ( .B(n11452), .A(n30504), .Z(n11453) );
  NANDN U27362 ( .A(n30494), .B(n11453), .Z(n11454) );
  NANDN U27363 ( .A(x[546]), .B(y[546]), .Z(n28366) );
  AND U27364 ( .A(n11454), .B(n28366), .Z(n11455) );
  NAND U27365 ( .A(n30499), .B(n11455), .Z(n11456) );
  ANDN U27366 ( .B(x[547]), .A(y[547]), .Z(n30509) );
  ANDN U27367 ( .B(n11456), .A(n30509), .Z(n11457) );
  NANDN U27368 ( .A(n30503), .B(n11457), .Z(n11458) );
  NAND U27369 ( .A(n28367), .B(n11458), .Z(n11460) );
  NANDN U27370 ( .A(x[548]), .B(n11460), .Z(n11459) );
  NANDN U27371 ( .A(x[549]), .B(y[549]), .Z(n28365) );
  AND U27372 ( .A(n11459), .B(n28365), .Z(n11463) );
  XNOR U27373 ( .A(x[548]), .B(n11460), .Z(n11461) );
  NAND U27374 ( .A(n11461), .B(y[548]), .Z(n11462) );
  NAND U27375 ( .A(n11463), .B(n11462), .Z(n11464) );
  NAND U27376 ( .A(n30514), .B(n11464), .Z(n52439) );
  NANDN U27377 ( .A(x[550]), .B(y[550]), .Z(n28363) );
  NAND U27378 ( .A(n52439), .B(n28363), .Z(n11465) );
  NANDN U27379 ( .A(n28360), .B(n11465), .Z(n11466) );
  ANDN U27380 ( .B(y[552]), .A(x[552]), .Z(n52441) );
  ANDN U27381 ( .B(n11466), .A(n52441), .Z(n11467) );
  NANDN U27382 ( .A(x[551]), .B(y[551]), .Z(n28362) );
  NAND U27383 ( .A(n11467), .B(n28362), .Z(n11468) );
  NANDN U27384 ( .A(y[553]), .B(x[553]), .Z(n52442) );
  AND U27385 ( .A(n11468), .B(n52442), .Z(n11469) );
  NAND U27386 ( .A(n28361), .B(n11469), .Z(n11470) );
  NAND U27387 ( .A(n52444), .B(n11470), .Z(n11471) );
  ANDN U27388 ( .B(x[555]), .A(y[555]), .Z(n28358) );
  ANDN U27389 ( .B(n11471), .A(n28358), .Z(n11472) );
  NAND U27390 ( .A(n52445), .B(n11472), .Z(n11473) );
  AND U27391 ( .A(n28359), .B(n11473), .Z(n11474) );
  NANDN U27392 ( .A(n52446), .B(n11474), .Z(n11475) );
  NANDN U27393 ( .A(n11476), .B(n11475), .Z(n11477) );
  ANDN U27394 ( .B(x[557]), .A(y[557]), .Z(n28356) );
  OR U27395 ( .A(n11477), .B(n28356), .Z(n11478) );
  AND U27396 ( .A(n11479), .B(n11478), .Z(n11481) );
  NANDN U27397 ( .A(y[559]), .B(x[559]), .Z(n52451) );
  NANDN U27398 ( .A(y[558]), .B(x[558]), .Z(n28357) );
  AND U27399 ( .A(n52451), .B(n28357), .Z(n11480) );
  NANDN U27400 ( .A(n11481), .B(n11480), .Z(n11482) );
  AND U27401 ( .A(n52452), .B(n11482), .Z(n11484) );
  NANDN U27402 ( .A(y[560]), .B(x[560]), .Z(n52453) );
  NANDN U27403 ( .A(y[561]), .B(x[561]), .Z(n28355) );
  AND U27404 ( .A(n52453), .B(n28355), .Z(n11483) );
  NANDN U27405 ( .A(n11484), .B(n11483), .Z(n11485) );
  ANDN U27406 ( .B(y[561]), .A(x[561]), .Z(n52454) );
  ANDN U27407 ( .B(n11485), .A(n52454), .Z(n11486) );
  NANDN U27408 ( .A(x[562]), .B(y[562]), .Z(n30540) );
  NAND U27409 ( .A(n11486), .B(n30540), .Z(n11487) );
  ANDN U27410 ( .B(x[563]), .A(y[563]), .Z(n28350) );
  ANDN U27411 ( .B(n11487), .A(n28350), .Z(n11488) );
  NANDN U27412 ( .A(n28353), .B(n11488), .Z(n11489) );
  ANDN U27413 ( .B(y[564]), .A(x[564]), .Z(n52457) );
  ANDN U27414 ( .B(n11489), .A(n52457), .Z(n11490) );
  NAND U27415 ( .A(n30541), .B(n11490), .Z(n11491) );
  NAND U27416 ( .A(n52458), .B(n11491), .Z(n11492) );
  NANDN U27417 ( .A(y[564]), .B(x[564]), .Z(n28352) );
  NANDN U27418 ( .A(n11492), .B(n28352), .Z(n11493) );
  NAND U27419 ( .A(n52459), .B(n11493), .Z(n11494) );
  NAND U27420 ( .A(n52460), .B(n11494), .Z(n11495) );
  NANDN U27421 ( .A(y[567]), .B(x[567]), .Z(n28349) );
  NANDN U27422 ( .A(n11495), .B(n28349), .Z(n11496) );
  AND U27423 ( .A(n11497), .B(n11496), .Z(n11499) );
  NANDN U27424 ( .A(y[569]), .B(x[569]), .Z(n28346) );
  ANDN U27425 ( .B(x[568]), .A(y[568]), .Z(n28347) );
  ANDN U27426 ( .B(n28346), .A(n28347), .Z(n11498) );
  NANDN U27427 ( .A(n11499), .B(n11498), .Z(n11500) );
  ANDN U27428 ( .B(y[570]), .A(x[570]), .Z(n52465) );
  ANDN U27429 ( .B(n11500), .A(n52465), .Z(n11501) );
  NANDN U27430 ( .A(x[569]), .B(y[569]), .Z(n30554) );
  NAND U27431 ( .A(n11501), .B(n30554), .Z(n11502) );
  AND U27432 ( .A(n52466), .B(n11502), .Z(n11503) );
  NANDN U27433 ( .A(n28345), .B(n11503), .Z(n11504) );
  AND U27434 ( .A(n52435), .B(n11504), .Z(n11505) );
  NAND U27435 ( .A(n28344), .B(n11505), .Z(n11506) );
  NANDN U27436 ( .A(n28341), .B(n11506), .Z(n11507) );
  NANDN U27437 ( .A(x[573]), .B(y[573]), .Z(n28343) );
  AND U27438 ( .A(n11507), .B(n28343), .Z(n11508) );
  NAND U27439 ( .A(n28340), .B(n11508), .Z(n11509) );
  NAND U27440 ( .A(n28342), .B(n11509), .Z(n11510) );
  NANDN U27441 ( .A(y[575]), .B(x[575]), .Z(n28338) );
  NANDN U27442 ( .A(n11510), .B(n28338), .Z(n11511) );
  AND U27443 ( .A(n11512), .B(n11511), .Z(n11514) );
  NANDN U27444 ( .A(y[577]), .B(x[577]), .Z(n52470) );
  ANDN U27445 ( .B(x[576]), .A(y[576]), .Z(n28336) );
  ANDN U27446 ( .B(n52470), .A(n28336), .Z(n11513) );
  NANDN U27447 ( .A(n11514), .B(n11513), .Z(n11515) );
  AND U27448 ( .A(n52471), .B(n11515), .Z(n11517) );
  NANDN U27449 ( .A(y[579]), .B(x[579]), .Z(n28335) );
  ANDN U27450 ( .B(x[578]), .A(y[578]), .Z(n52472) );
  ANDN U27451 ( .B(n28335), .A(n52472), .Z(n11516) );
  NANDN U27452 ( .A(n11517), .B(n11516), .Z(n11518) );
  ANDN U27453 ( .B(y[579]), .A(x[579]), .Z(n52473) );
  ANDN U27454 ( .B(n11518), .A(n52473), .Z(n11519) );
  NANDN U27455 ( .A(x[580]), .B(y[580]), .Z(n28333) );
  NAND U27456 ( .A(n11519), .B(n28333), .Z(n11520) );
  NANDN U27457 ( .A(y[581]), .B(x[581]), .Z(n28331) );
  AND U27458 ( .A(n11520), .B(n28331), .Z(n11521) );
  NANDN U27459 ( .A(n28334), .B(n11521), .Z(n11522) );
  ANDN U27460 ( .B(y[582]), .A(x[582]), .Z(n52477) );
  ANDN U27461 ( .B(n11522), .A(n52477), .Z(n11523) );
  NAND U27462 ( .A(n28332), .B(n11523), .Z(n11524) );
  NANDN U27463 ( .A(n28329), .B(n11524), .Z(n11525) );
  NANDN U27464 ( .A(y[583]), .B(x[583]), .Z(n52478) );
  NANDN U27465 ( .A(n11525), .B(n52478), .Z(n11526) );
  NAND U27466 ( .A(n52479), .B(n11526), .Z(n11527) );
  NAND U27467 ( .A(n52480), .B(n11527), .Z(n11528) );
  ANDN U27468 ( .B(x[585]), .A(y[585]), .Z(n28327) );
  OR U27469 ( .A(n11528), .B(n28327), .Z(n11529) );
  AND U27470 ( .A(n11530), .B(n11529), .Z(n11532) );
  NANDN U27471 ( .A(y[586]), .B(x[586]), .Z(n28328) );
  ANDN U27472 ( .B(x[587]), .A(y[587]), .Z(n28322) );
  ANDN U27473 ( .B(n28328), .A(n28322), .Z(n11531) );
  NANDN U27474 ( .A(n11532), .B(n11531), .Z(n11533) );
  AND U27475 ( .A(n52485), .B(n11533), .Z(n11534) );
  NANDN U27476 ( .A(x[587]), .B(y[587]), .Z(n28326) );
  NAND U27477 ( .A(n11534), .B(n28326), .Z(n11535) );
  NANDN U27478 ( .A(y[588]), .B(x[588]), .Z(n28323) );
  AND U27479 ( .A(n11535), .B(n28323), .Z(n11536) );
  NANDN U27480 ( .A(n52486), .B(n11536), .Z(n11537) );
  NAND U27481 ( .A(n52487), .B(n11537), .Z(n11538) );
  NANDN U27482 ( .A(y[591]), .B(x[591]), .Z(n28321) );
  AND U27483 ( .A(n11538), .B(n28321), .Z(n11539) );
  NAND U27484 ( .A(n52488), .B(n11539), .Z(n11540) );
  ANDN U27485 ( .B(y[591]), .A(x[591]), .Z(n52489) );
  ANDN U27486 ( .B(n11540), .A(n52489), .Z(n11541) );
  NAND U27487 ( .A(n30598), .B(n11541), .Z(n11542) );
  NANDN U27488 ( .A(n28319), .B(n11542), .Z(n11543) );
  NANDN U27489 ( .A(y[593]), .B(x[593]), .Z(n28318) );
  NANDN U27490 ( .A(n11543), .B(n28318), .Z(n11544) );
  AND U27491 ( .A(n11545), .B(n11544), .Z(n11547) );
  NANDN U27492 ( .A(y[595]), .B(x[595]), .Z(n52494) );
  ANDN U27493 ( .B(x[594]), .A(y[594]), .Z(n28317) );
  ANDN U27494 ( .B(n52494), .A(n28317), .Z(n11546) );
  NANDN U27495 ( .A(n11547), .B(n11546), .Z(n11548) );
  AND U27496 ( .A(n52495), .B(n11548), .Z(n11550) );
  NANDN U27497 ( .A(y[596]), .B(x[596]), .Z(n52496) );
  NANDN U27498 ( .A(y[597]), .B(x[597]), .Z(n28316) );
  AND U27499 ( .A(n52496), .B(n28316), .Z(n11549) );
  NANDN U27500 ( .A(n11550), .B(n11549), .Z(n11551) );
  ANDN U27501 ( .B(y[597]), .A(x[597]), .Z(n52497) );
  ANDN U27502 ( .B(n11551), .A(n52497), .Z(n11552) );
  NANDN U27503 ( .A(x[598]), .B(y[598]), .Z(n28312) );
  NAND U27504 ( .A(n11552), .B(n28312), .Z(n11553) );
  NANDN U27505 ( .A(y[599]), .B(x[599]), .Z(n28311) );
  AND U27506 ( .A(n11553), .B(n28311), .Z(n11554) );
  NANDN U27507 ( .A(n28314), .B(n11554), .Z(n11555) );
  ANDN U27508 ( .B(y[600]), .A(x[600]), .Z(n52501) );
  ANDN U27509 ( .B(n11555), .A(n52501), .Z(n11556) );
  NAND U27510 ( .A(n28313), .B(n11556), .Z(n11557) );
  NAND U27511 ( .A(n52502), .B(n11557), .Z(n11558) );
  ANDN U27512 ( .B(x[600]), .A(y[600]), .Z(n28310) );
  OR U27513 ( .A(n11558), .B(n28310), .Z(n11559) );
  NAND U27514 ( .A(n52503), .B(n11559), .Z(n11560) );
  NAND U27515 ( .A(n52504), .B(n11560), .Z(n11561) );
  NANDN U27516 ( .A(y[603]), .B(x[603]), .Z(n28309) );
  NANDN U27517 ( .A(n11561), .B(n28309), .Z(n11562) );
  AND U27518 ( .A(n11563), .B(n11562), .Z(n11565) );
  NANDN U27519 ( .A(y[605]), .B(x[605]), .Z(n28304) );
  ANDN U27520 ( .B(x[604]), .A(y[604]), .Z(n28307) );
  ANDN U27521 ( .B(n28304), .A(n28307), .Z(n11564) );
  NANDN U27522 ( .A(n11565), .B(n11564), .Z(n11566) );
  ANDN U27523 ( .B(y[606]), .A(x[606]), .Z(n52508) );
  ANDN U27524 ( .B(n11566), .A(n52508), .Z(n11567) );
  NANDN U27525 ( .A(x[605]), .B(y[605]), .Z(n28306) );
  NAND U27526 ( .A(n11567), .B(n28306), .Z(n11568) );
  ANDN U27527 ( .B(x[606]), .A(y[606]), .Z(n28302) );
  ANDN U27528 ( .B(n11568), .A(n28302), .Z(n11569) );
  NAND U27529 ( .A(n52510), .B(n11569), .Z(n11570) );
  NAND U27530 ( .A(n52511), .B(n11570), .Z(n11571) );
  ANDN U27531 ( .B(x[609]), .A(y[609]), .Z(n28299) );
  ANDN U27532 ( .B(n11571), .A(n28299), .Z(n11572) );
  NANDN U27533 ( .A(n52512), .B(n11572), .Z(n11573) );
  AND U27534 ( .A(n28301), .B(n11573), .Z(n11574) );
  NANDN U27535 ( .A(n52513), .B(n11574), .Z(n11575) );
  NANDN U27536 ( .A(n11576), .B(n11575), .Z(n11577) );
  NANDN U27537 ( .A(y[611]), .B(x[611]), .Z(n28296) );
  NANDN U27538 ( .A(n11577), .B(n28296), .Z(n11578) );
  AND U27539 ( .A(n11579), .B(n11578), .Z(n11581) );
  NANDN U27540 ( .A(y[613]), .B(x[613]), .Z(n52517) );
  ANDN U27541 ( .B(x[612]), .A(y[612]), .Z(n28295) );
  ANDN U27542 ( .B(n52517), .A(n28295), .Z(n11580) );
  NANDN U27543 ( .A(n11581), .B(n11580), .Z(n11582) );
  AND U27544 ( .A(n52518), .B(n11582), .Z(n11584) );
  NANDN U27545 ( .A(y[614]), .B(x[614]), .Z(n52519) );
  ANDN U27546 ( .B(x[615]), .A(y[615]), .Z(n28293) );
  ANDN U27547 ( .B(n52519), .A(n28293), .Z(n11583) );
  NANDN U27548 ( .A(n11584), .B(n11583), .Z(n11585) );
  ANDN U27549 ( .B(y[615]), .A(x[615]), .Z(n52520) );
  ANDN U27550 ( .B(n11585), .A(n52520), .Z(n11586) );
  NANDN U27551 ( .A(x[616]), .B(y[616]), .Z(n28292) );
  NAND U27552 ( .A(n11586), .B(n28292), .Z(n11587) );
  ANDN U27553 ( .B(x[617]), .A(y[617]), .Z(n28289) );
  ANDN U27554 ( .B(n11587), .A(n28289), .Z(n11588) );
  NAND U27555 ( .A(n28294), .B(n11588), .Z(n11589) );
  ANDN U27556 ( .B(y[618]), .A(x[618]), .Z(n52524) );
  ANDN U27557 ( .B(n11589), .A(n52524), .Z(n11590) );
  NAND U27558 ( .A(n28291), .B(n11590), .Z(n11591) );
  NAND U27559 ( .A(n52525), .B(n11591), .Z(n11592) );
  NANDN U27560 ( .A(y[618]), .B(x[618]), .Z(n28290) );
  NANDN U27561 ( .A(n11592), .B(n28290), .Z(n11593) );
  NAND U27562 ( .A(n52526), .B(n11593), .Z(n11594) );
  NANDN U27563 ( .A(n52528), .B(n11594), .Z(n11595) );
  NAND U27564 ( .A(n52530), .B(n11595), .Z(n11596) );
  NANDN U27565 ( .A(n52532), .B(n11596), .Z(n11597) );
  AND U27566 ( .A(n52534), .B(n11597), .Z(n11598) );
  OR U27567 ( .A(n52536), .B(n11598), .Z(n11599) );
  NAND U27568 ( .A(n52538), .B(n11599), .Z(n11600) );
  NANDN U27569 ( .A(n52540), .B(n11600), .Z(n11601) );
  NAND U27570 ( .A(n52542), .B(n11601), .Z(n11602) );
  NANDN U27571 ( .A(n52544), .B(n11602), .Z(n11603) );
  AND U27572 ( .A(n52546), .B(n11603), .Z(n11604) );
  OR U27573 ( .A(n52548), .B(n11604), .Z(n11605) );
  NAND U27574 ( .A(n52550), .B(n11605), .Z(n11606) );
  NANDN U27575 ( .A(n52552), .B(n11606), .Z(n11607) );
  NAND U27576 ( .A(n52554), .B(n11607), .Z(n11608) );
  NANDN U27577 ( .A(n52556), .B(n11608), .Z(n11609) );
  AND U27578 ( .A(n52558), .B(n11609), .Z(n11610) );
  OR U27579 ( .A(n52560), .B(n11610), .Z(n11611) );
  NAND U27580 ( .A(n52562), .B(n11611), .Z(n11612) );
  NANDN U27581 ( .A(n52564), .B(n11612), .Z(n11613) );
  NAND U27582 ( .A(n52566), .B(n11613), .Z(n11614) );
  NANDN U27583 ( .A(n52568), .B(n11614), .Z(n11615) );
  AND U27584 ( .A(n52569), .B(n11615), .Z(n11616) );
  OR U27585 ( .A(n52570), .B(n11616), .Z(n11617) );
  AND U27586 ( .A(n11618), .B(n11617), .Z(n11619) );
  OR U27587 ( .A(n11620), .B(n11619), .Z(n11621) );
  AND U27588 ( .A(n11622), .B(n11621), .Z(n11623) );
  OR U27589 ( .A(n52574), .B(n11623), .Z(n11624) );
  NAND U27590 ( .A(n52575), .B(n11624), .Z(n11625) );
  NANDN U27591 ( .A(n52576), .B(n11625), .Z(n11626) );
  NAND U27592 ( .A(n52577), .B(n11626), .Z(n11627) );
  NANDN U27593 ( .A(n52578), .B(n11627), .Z(n11628) );
  AND U27594 ( .A(n52579), .B(n11628), .Z(n11629) );
  OR U27595 ( .A(n52580), .B(n11629), .Z(n11630) );
  NAND U27596 ( .A(n52581), .B(n11630), .Z(n11631) );
  NANDN U27597 ( .A(n52582), .B(n11631), .Z(n11632) );
  NAND U27598 ( .A(n52584), .B(n11632), .Z(n11633) );
  NANDN U27599 ( .A(n52585), .B(n11633), .Z(n11634) );
  AND U27600 ( .A(n52586), .B(n11634), .Z(n11637) );
  NANDN U27601 ( .A(y[658]), .B(x[658]), .Z(n11636) );
  NANDN U27602 ( .A(y[659]), .B(x[659]), .Z(n11635) );
  AND U27603 ( .A(n11636), .B(n11635), .Z(n52587) );
  NANDN U27604 ( .A(n11637), .B(n52587), .Z(n11638) );
  NANDN U27605 ( .A(n52588), .B(n11638), .Z(n11639) );
  NAND U27606 ( .A(n52589), .B(n11639), .Z(n11640) );
  NANDN U27607 ( .A(n52590), .B(n11640), .Z(n11641) );
  NAND U27608 ( .A(n52426), .B(n11641), .Z(n11642) );
  NANDN U27609 ( .A(n52425), .B(n11642), .Z(n11643) );
  ANDN U27610 ( .B(y[664]), .A(x[664]), .Z(n28275) );
  OR U27611 ( .A(n11643), .B(n28275), .Z(n11644) );
  AND U27612 ( .A(n11645), .B(n11644), .Z(n11647) );
  NANDN U27613 ( .A(x[665]), .B(y[665]), .Z(n28276) );
  ANDN U27614 ( .B(y[666]), .A(x[666]), .Z(n52423) );
  ANDN U27615 ( .B(n28276), .A(n52423), .Z(n11646) );
  NANDN U27616 ( .A(n11647), .B(n11646), .Z(n11648) );
  NANDN U27617 ( .A(y[666]), .B(x[666]), .Z(n30796) );
  NANDN U27618 ( .A(y[667]), .B(x[667]), .Z(n30801) );
  AND U27619 ( .A(n30796), .B(n30801), .Z(n52422) );
  AND U27620 ( .A(n11648), .B(n52422), .Z(n11649) );
  ANDN U27621 ( .B(y[667]), .A(x[667]), .Z(n30798) );
  ANDN U27622 ( .B(y[668]), .A(x[668]), .Z(n30807) );
  OR U27623 ( .A(n30798), .B(n30807), .Z(n52421) );
  OR U27624 ( .A(n11649), .B(n52421), .Z(n11650) );
  NAND U27625 ( .A(n52420), .B(n11650), .Z(n11651) );
  NANDN U27626 ( .A(n52594), .B(n11651), .Z(n11652) );
  NAND U27627 ( .A(n52595), .B(n11652), .Z(n11653) );
  NANDN U27628 ( .A(n52419), .B(n11653), .Z(n11654) );
  NANDN U27629 ( .A(y[672]), .B(x[672]), .Z(n30816) );
  NANDN U27630 ( .A(y[673]), .B(x[673]), .Z(n30823) );
  AND U27631 ( .A(n30816), .B(n30823), .Z(n52418) );
  AND U27632 ( .A(n11654), .B(n52418), .Z(n11656) );
  ANDN U27633 ( .B(y[673]), .A(x[673]), .Z(n30822) );
  IV U27634 ( .A(n30822), .Z(n52596) );
  ANDN U27635 ( .B(y[674]), .A(x[674]), .Z(n28272) );
  ANDN U27636 ( .B(n52596), .A(n28272), .Z(n11655) );
  NANDN U27637 ( .A(n11656), .B(n11655), .Z(n11657) );
  NANDN U27638 ( .A(y[675]), .B(x[675]), .Z(n52598) );
  AND U27639 ( .A(n11657), .B(n52598), .Z(n11658) );
  NAND U27640 ( .A(n52417), .B(n11658), .Z(n11659) );
  ANDN U27641 ( .B(y[675]), .A(x[675]), .Z(n28271) );
  ANDN U27642 ( .B(n11659), .A(n28271), .Z(n11660) );
  NANDN U27643 ( .A(n52416), .B(n11660), .Z(n11661) );
  NAND U27644 ( .A(n52415), .B(n11661), .Z(n11662) );
  NANDN U27645 ( .A(n52414), .B(n11662), .Z(n11663) );
  NANDN U27646 ( .A(y[678]), .B(x[678]), .Z(n30834) );
  NANDN U27647 ( .A(y[679]), .B(x[679]), .Z(n30841) );
  AND U27648 ( .A(n30834), .B(n30841), .Z(n52413) );
  AND U27649 ( .A(n11663), .B(n52413), .Z(n11664) );
  ANDN U27650 ( .B(y[679]), .A(x[679]), .Z(n30837) );
  ANDN U27651 ( .B(y[680]), .A(x[680]), .Z(n30847) );
  OR U27652 ( .A(n30837), .B(n30847), .Z(n52600) );
  OR U27653 ( .A(n11664), .B(n52600), .Z(n11665) );
  NAND U27654 ( .A(n52601), .B(n11665), .Z(n11666) );
  NANDN U27655 ( .A(n52412), .B(n11666), .Z(n11667) );
  NAND U27656 ( .A(n52602), .B(n11667), .Z(n11668) );
  ANDN U27657 ( .B(y[684]), .A(x[684]), .Z(n28267) );
  ANDN U27658 ( .B(n11668), .A(n28267), .Z(n11669) );
  NANDN U27659 ( .A(n30851), .B(n11669), .Z(n11671) );
  NANDN U27660 ( .A(y[684]), .B(x[684]), .Z(n52604) );
  NANDN U27661 ( .A(y[685]), .B(x[685]), .Z(n52606) );
  AND U27662 ( .A(n52604), .B(n52606), .Z(n11670) );
  NAND U27663 ( .A(n11671), .B(n11670), .Z(n11672) );
  AND U27664 ( .A(n52607), .B(n11672), .Z(n11673) );
  NANDN U27665 ( .A(x[685]), .B(y[685]), .Z(n28268) );
  NAND U27666 ( .A(n11673), .B(n28268), .Z(n11674) );
  NANDN U27667 ( .A(n52608), .B(n11674), .Z(n11675) );
  AND U27668 ( .A(n52609), .B(n11675), .Z(n11676) );
  OR U27669 ( .A(n52611), .B(n11676), .Z(n11677) );
  NAND U27670 ( .A(n52613), .B(n11677), .Z(n11678) );
  NANDN U27671 ( .A(n52615), .B(n11678), .Z(n11679) );
  NAND U27672 ( .A(n52617), .B(n11679), .Z(n11680) );
  NANDN U27673 ( .A(n52619), .B(n11680), .Z(n11681) );
  AND U27674 ( .A(n52621), .B(n11681), .Z(n11682) );
  OR U27675 ( .A(n52623), .B(n11682), .Z(n11683) );
  NAND U27676 ( .A(n52625), .B(n11683), .Z(n11684) );
  NANDN U27677 ( .A(n52627), .B(n11684), .Z(n11685) );
  NAND U27678 ( .A(n52629), .B(n11685), .Z(n11686) );
  NANDN U27679 ( .A(n52631), .B(n11686), .Z(n11687) );
  AND U27680 ( .A(n52633), .B(n11687), .Z(n11688) );
  OR U27681 ( .A(n52635), .B(n11688), .Z(n11689) );
  NAND U27682 ( .A(n52637), .B(n11689), .Z(n11690) );
  NANDN U27683 ( .A(n52639), .B(n11690), .Z(n11691) );
  NAND U27684 ( .A(n52641), .B(n11691), .Z(n11692) );
  NANDN U27685 ( .A(n52643), .B(n11692), .Z(n11693) );
  AND U27686 ( .A(n52645), .B(n11693), .Z(n11694) );
  OR U27687 ( .A(n52647), .B(n11694), .Z(n11695) );
  NAND U27688 ( .A(n52649), .B(n11695), .Z(n11696) );
  NANDN U27689 ( .A(n52651), .B(n11696), .Z(n11697) );
  NAND U27690 ( .A(n52652), .B(n11697), .Z(n11698) );
  NANDN U27691 ( .A(n52653), .B(n11698), .Z(n11699) );
  AND U27692 ( .A(n52654), .B(n11699), .Z(n11700) );
  OR U27693 ( .A(n52655), .B(n11700), .Z(n11701) );
  AND U27694 ( .A(n11702), .B(n11701), .Z(n11703) );
  OR U27695 ( .A(n11704), .B(n11703), .Z(n11705) );
  AND U27696 ( .A(n11706), .B(n11705), .Z(n11707) );
  OR U27697 ( .A(n52661), .B(n11707), .Z(n11708) );
  NAND U27698 ( .A(n52662), .B(n11708), .Z(n11709) );
  NANDN U27699 ( .A(n52663), .B(n11709), .Z(n11710) );
  NAND U27700 ( .A(n52664), .B(n11710), .Z(n11711) );
  NANDN U27701 ( .A(n52665), .B(n11711), .Z(n11712) );
  AND U27702 ( .A(n52666), .B(n11712), .Z(n11713) );
  OR U27703 ( .A(n52667), .B(n11713), .Z(n11714) );
  AND U27704 ( .A(n11715), .B(n11714), .Z(n11716) );
  OR U27705 ( .A(n11717), .B(n11716), .Z(n11718) );
  AND U27706 ( .A(n11719), .B(n11718), .Z(n11720) );
  OR U27707 ( .A(n52672), .B(n11720), .Z(n11721) );
  NAND U27708 ( .A(n52673), .B(n11721), .Z(n11722) );
  NANDN U27709 ( .A(n52674), .B(n11722), .Z(n11723) );
  NAND U27710 ( .A(n52675), .B(n11723), .Z(n11724) );
  NANDN U27711 ( .A(n52676), .B(n11724), .Z(n11725) );
  AND U27712 ( .A(n52677), .B(n11725), .Z(n11726) );
  OR U27713 ( .A(n52678), .B(n11726), .Z(n11727) );
  AND U27714 ( .A(n11728), .B(n11727), .Z(n11729) );
  OR U27715 ( .A(n11730), .B(n11729), .Z(n11731) );
  NAND U27716 ( .A(n52683), .B(n11731), .Z(n11732) );
  NANDN U27717 ( .A(n52684), .B(n11732), .Z(n11733) );
  NAND U27718 ( .A(n52685), .B(n11733), .Z(n11734) );
  NANDN U27719 ( .A(n52686), .B(n11734), .Z(n11735) );
  AND U27720 ( .A(n52688), .B(n11735), .Z(n11736) );
  OR U27721 ( .A(n52690), .B(n11736), .Z(n11737) );
  NAND U27722 ( .A(n52692), .B(n11737), .Z(n11738) );
  NANDN U27723 ( .A(n52694), .B(n11738), .Z(n11739) );
  NANDN U27724 ( .A(x[743]), .B(y[743]), .Z(n52696) );
  AND U27725 ( .A(n11739), .B(n52696), .Z(n11740) );
  NAND U27726 ( .A(n52700), .B(n11740), .Z(n11741) );
  NAND U27727 ( .A(n11742), .B(n11741), .Z(n11743) );
  NAND U27728 ( .A(n52704), .B(n11743), .Z(n11744) );
  NANDN U27729 ( .A(n52706), .B(n11744), .Z(n11745) );
  AND U27730 ( .A(n52708), .B(n11745), .Z(n11746) );
  OR U27731 ( .A(n52710), .B(n11746), .Z(n11747) );
  NAND U27732 ( .A(n52712), .B(n11747), .Z(n11748) );
  NANDN U27733 ( .A(n52714), .B(n11748), .Z(n11749) );
  NAND U27734 ( .A(n52716), .B(n11749), .Z(n11750) );
  NANDN U27735 ( .A(n52718), .B(n11750), .Z(n11751) );
  AND U27736 ( .A(n52720), .B(n11751), .Z(n11752) );
  OR U27737 ( .A(n52722), .B(n11752), .Z(n11753) );
  NAND U27738 ( .A(n52724), .B(n11753), .Z(n11754) );
  NANDN U27739 ( .A(n52726), .B(n11754), .Z(n11755) );
  NAND U27740 ( .A(n52728), .B(n11755), .Z(n11756) );
  NANDN U27741 ( .A(n52729), .B(n11756), .Z(n11757) );
  AND U27742 ( .A(n52730), .B(n11757), .Z(n11758) );
  OR U27743 ( .A(n52731), .B(n11758), .Z(n11759) );
  NAND U27744 ( .A(n52732), .B(n11759), .Z(n11760) );
  NANDN U27745 ( .A(n52733), .B(n11760), .Z(n11761) );
  NANDN U27746 ( .A(x[764]), .B(y[764]), .Z(n28232) );
  AND U27747 ( .A(n11761), .B(n28232), .Z(n11762) );
  NANDN U27748 ( .A(n52734), .B(n11762), .Z(n11763) );
  NANDN U27749 ( .A(n11764), .B(n11763), .Z(n11765) );
  NANDN U27750 ( .A(x[765]), .B(y[765]), .Z(n28231) );
  AND U27751 ( .A(n11765), .B(n28231), .Z(n11766) );
  NAND U27752 ( .A(n31113), .B(n11766), .Z(n11767) );
  NANDN U27753 ( .A(n52409), .B(n11767), .Z(n11768) );
  NAND U27754 ( .A(n52739), .B(n11768), .Z(n11769) );
  NANDN U27755 ( .A(n52408), .B(n11769), .Z(n11770) );
  AND U27756 ( .A(n52740), .B(n11770), .Z(n11771) );
  ANDN U27757 ( .B(x[771]), .A(y[771]), .Z(n28229) );
  NANDN U27758 ( .A(y[770]), .B(x[770]), .Z(n31124) );
  NANDN U27759 ( .A(n28229), .B(n31124), .Z(n52741) );
  OR U27760 ( .A(n11771), .B(n52741), .Z(n11772) );
  NAND U27761 ( .A(n52742), .B(n11772), .Z(n11773) );
  NANDN U27762 ( .A(n52407), .B(n11773), .Z(n11774) );
  NANDN U27763 ( .A(x[773]), .B(y[773]), .Z(n52406) );
  AND U27764 ( .A(n11774), .B(n52406), .Z(n11775) );
  NAND U27765 ( .A(n52405), .B(n11775), .Z(n11776) );
  NAND U27766 ( .A(n11777), .B(n11776), .Z(n11778) );
  NAND U27767 ( .A(n52747), .B(n11778), .Z(n11779) );
  NANDN U27768 ( .A(n52404), .B(n11779), .Z(n11780) );
  NANDN U27769 ( .A(x[777]), .B(y[777]), .Z(n31146) );
  NANDN U27770 ( .A(x[778]), .B(y[778]), .Z(n28228) );
  AND U27771 ( .A(n31146), .B(n28228), .Z(n52403) );
  AND U27772 ( .A(n11780), .B(n52403), .Z(n11781) );
  ANDN U27773 ( .B(x[778]), .A(y[778]), .Z(n31150) );
  ANDN U27774 ( .B(x[779]), .A(y[779]), .Z(n31156) );
  OR U27775 ( .A(n31150), .B(n31156), .Z(n52402) );
  OR U27776 ( .A(n11781), .B(n52402), .Z(n11782) );
  NAND U27777 ( .A(n52401), .B(n11782), .Z(n11783) );
  NAND U27778 ( .A(n52748), .B(n11783), .Z(n11784) );
  NAND U27779 ( .A(n52749), .B(n11784), .Z(n11785) );
  NANDN U27780 ( .A(n52750), .B(n11785), .Z(n11786) );
  AND U27781 ( .A(n52752), .B(n11786), .Z(n11787) );
  NANDN U27782 ( .A(x[784]), .B(y[784]), .Z(n28226) );
  NAND U27783 ( .A(n11787), .B(n28226), .Z(n11788) );
  NANDN U27784 ( .A(n11789), .B(n11788), .Z(n11790) );
  AND U27785 ( .A(n52755), .B(n11790), .Z(n11791) );
  NANDN U27786 ( .A(x[785]), .B(y[785]), .Z(n28225) );
  NAND U27787 ( .A(n11791), .B(n28225), .Z(n11792) );
  NANDN U27788 ( .A(n52756), .B(n11792), .Z(n11793) );
  AND U27789 ( .A(n52757), .B(n11793), .Z(n11794) );
  OR U27790 ( .A(n52758), .B(n11794), .Z(n11795) );
  NAND U27791 ( .A(n52759), .B(n11795), .Z(n11796) );
  NANDN U27792 ( .A(n52760), .B(n11796), .Z(n11797) );
  NAND U27793 ( .A(n52761), .B(n11797), .Z(n11798) );
  NANDN U27794 ( .A(n52762), .B(n11798), .Z(n11799) );
  ANDN U27795 ( .B(y[793]), .A(x[793]), .Z(n52763) );
  ANDN U27796 ( .B(n11799), .A(n52763), .Z(n11800) );
  NANDN U27797 ( .A(x[794]), .B(y[794]), .Z(n28221) );
  NAND U27798 ( .A(n11800), .B(n28221), .Z(n11801) );
  NANDN U27799 ( .A(n11802), .B(n11801), .Z(n11803) );
  ANDN U27800 ( .B(y[796]), .A(x[796]), .Z(n52766) );
  ANDN U27801 ( .B(n11803), .A(n52766), .Z(n11804) );
  NANDN U27802 ( .A(x[795]), .B(y[795]), .Z(n28220) );
  NAND U27803 ( .A(n11804), .B(n28220), .Z(n11805) );
  NANDN U27804 ( .A(n52768), .B(n11805), .Z(n11806) );
  AND U27805 ( .A(n52770), .B(n11806), .Z(n11807) );
  OR U27806 ( .A(n52772), .B(n11807), .Z(n11808) );
  NAND U27807 ( .A(n52774), .B(n11808), .Z(n11809) );
  NANDN U27808 ( .A(n52776), .B(n11809), .Z(n11810) );
  NAND U27809 ( .A(n52778), .B(n11810), .Z(n11811) );
  NANDN U27810 ( .A(n52780), .B(n11811), .Z(n11812) );
  AND U27811 ( .A(n52782), .B(n11812), .Z(n11813) );
  OR U27812 ( .A(n52784), .B(n11813), .Z(n11814) );
  NAND U27813 ( .A(n52786), .B(n11814), .Z(n11815) );
  NANDN U27814 ( .A(n52788), .B(n11815), .Z(n11816) );
  NAND U27815 ( .A(n52790), .B(n11816), .Z(n11817) );
  NANDN U27816 ( .A(n52792), .B(n11817), .Z(n11818) );
  AND U27817 ( .A(n52794), .B(n11818), .Z(n11819) );
  OR U27818 ( .A(n52796), .B(n11819), .Z(n11820) );
  NAND U27819 ( .A(n52798), .B(n11820), .Z(n11821) );
  NANDN U27820 ( .A(n52800), .B(n11821), .Z(n11822) );
  ANDN U27821 ( .B(y[813]), .A(x[813]), .Z(n52802) );
  ANDN U27822 ( .B(n11822), .A(n52802), .Z(n11823) );
  NAND U27823 ( .A(n28208), .B(n11823), .Z(n11824) );
  NAND U27824 ( .A(n52808), .B(n11824), .Z(n11825) );
  NANDN U27825 ( .A(y[814]), .B(x[814]), .Z(n52804) );
  NANDN U27826 ( .A(n11825), .B(n52804), .Z(n11826) );
  AND U27827 ( .A(n11827), .B(n11826), .Z(n11828) );
  OR U27828 ( .A(n52813), .B(n11828), .Z(n11829) );
  NAND U27829 ( .A(n52815), .B(n11829), .Z(n11830) );
  NANDN U27830 ( .A(n52817), .B(n11830), .Z(n11831) );
  NAND U27831 ( .A(n52819), .B(n11831), .Z(n11832) );
  NANDN U27832 ( .A(n52821), .B(n11832), .Z(n11833) );
  AND U27833 ( .A(n52823), .B(n11833), .Z(n11834) );
  OR U27834 ( .A(n52825), .B(n11834), .Z(n11835) );
  NAND U27835 ( .A(n52827), .B(n11835), .Z(n11836) );
  NANDN U27836 ( .A(n52829), .B(n11836), .Z(n11837) );
  NAND U27837 ( .A(n52831), .B(n11837), .Z(n11838) );
  NANDN U27838 ( .A(n52833), .B(n11838), .Z(n11839) );
  AND U27839 ( .A(n52835), .B(n11839), .Z(n11840) );
  OR U27840 ( .A(n52837), .B(n11840), .Z(n11841) );
  NAND U27841 ( .A(n52839), .B(n11841), .Z(n11842) );
  NANDN U27842 ( .A(n52841), .B(n11842), .Z(n11843) );
  NAND U27843 ( .A(n52843), .B(n11843), .Z(n11844) );
  NANDN U27844 ( .A(n52845), .B(n11844), .Z(n11845) );
  ANDN U27845 ( .B(y[833]), .A(x[833]), .Z(n52847) );
  ANDN U27846 ( .B(n11845), .A(n52847), .Z(n11846) );
  NANDN U27847 ( .A(x[834]), .B(y[834]), .Z(n28197) );
  NAND U27848 ( .A(n11846), .B(n28197), .Z(n11847) );
  NANDN U27849 ( .A(y[835]), .B(x[835]), .Z(n52849) );
  AND U27850 ( .A(n11847), .B(n52849), .Z(n11848) );
  NAND U27851 ( .A(n52848), .B(n11848), .Z(n11849) );
  ANDN U27852 ( .B(y[836]), .A(x[836]), .Z(n52850) );
  ANDN U27853 ( .B(n11849), .A(n52850), .Z(n11850) );
  NAND U27854 ( .A(n28198), .B(n11850), .Z(n11851) );
  NANDN U27855 ( .A(n52851), .B(n11851), .Z(n11852) );
  NANDN U27856 ( .A(n52852), .B(n11852), .Z(n11853) );
  NANDN U27857 ( .A(n52853), .B(n11853), .Z(n11854) );
  AND U27858 ( .A(n52854), .B(n11854), .Z(n11855) );
  OR U27859 ( .A(n52855), .B(n11855), .Z(n11856) );
  NAND U27860 ( .A(n52856), .B(n11856), .Z(n11857) );
  NANDN U27861 ( .A(n52857), .B(n11857), .Z(n11859) );
  ANDN U27862 ( .B(y[843]), .A(x[843]), .Z(n52858) );
  ANDN U27863 ( .B(y[844]), .A(x[844]), .Z(n52860) );
  NOR U27864 ( .A(n52858), .B(n52860), .Z(n11858) );
  NAND U27865 ( .A(n11859), .B(n11858), .Z(n11860) );
  AND U27866 ( .A(n11861), .B(n11860), .Z(n11862) );
  ANDN U27867 ( .B(y[845]), .A(x[845]), .Z(n31352) );
  NANDN U27868 ( .A(x[846]), .B(y[846]), .Z(n28190) );
  NANDN U27869 ( .A(n31352), .B(n28190), .Z(n52396) );
  OR U27870 ( .A(n11862), .B(n52396), .Z(n11863) );
  NAND U27871 ( .A(n52863), .B(n11863), .Z(n11864) );
  NANDN U27872 ( .A(n52864), .B(n11864), .Z(n11865) );
  NAND U27873 ( .A(n52865), .B(n11865), .Z(n11866) );
  NANDN U27874 ( .A(n52395), .B(n11866), .Z(n11867) );
  NANDN U27875 ( .A(y[850]), .B(x[850]), .Z(n28187) );
  NANDN U27876 ( .A(y[851]), .B(x[851]), .Z(n31370) );
  AND U27877 ( .A(n28187), .B(n31370), .Z(n52394) );
  AND U27878 ( .A(n11867), .B(n52394), .Z(n11869) );
  NANDN U27879 ( .A(x[851]), .B(y[851]), .Z(n28185) );
  XNOR U27880 ( .A(x[852]), .B(y[852]), .Z(n11868) );
  NAND U27881 ( .A(n28185), .B(n11868), .Z(n52393) );
  OR U27882 ( .A(n11869), .B(n52393), .Z(n11870) );
  NAND U27883 ( .A(n52392), .B(n11870), .Z(n11871) );
  NANDN U27884 ( .A(n52866), .B(n11871), .Z(n11872) );
  NAND U27885 ( .A(n52867), .B(n11872), .Z(n11873) );
  NANDN U27886 ( .A(n52391), .B(n11873), .Z(n11874) );
  NANDN U27887 ( .A(y[856]), .B(x[856]), .Z(n31387) );
  NANDN U27888 ( .A(y[857]), .B(x[857]), .Z(n28183) );
  AND U27889 ( .A(n31387), .B(n28183), .Z(n52390) );
  AND U27890 ( .A(n11874), .B(n52390), .Z(n11875) );
  ANDN U27891 ( .B(y[857]), .A(x[857]), .Z(n31391) );
  NANDN U27892 ( .A(x[858]), .B(y[858]), .Z(n31397) );
  NANDN U27893 ( .A(n31391), .B(n31397), .Z(n52389) );
  OR U27894 ( .A(n11875), .B(n52389), .Z(n11876) );
  NAND U27895 ( .A(n52388), .B(n11876), .Z(n11877) );
  NANDN U27896 ( .A(n52870), .B(n11877), .Z(n11878) );
  NAND U27897 ( .A(n52871), .B(n11878), .Z(n11879) );
  NANDN U27898 ( .A(n52387), .B(n11879), .Z(n11880) );
  NANDN U27899 ( .A(y[862]), .B(x[862]), .Z(n31409) );
  NANDN U27900 ( .A(y[863]), .B(x[863]), .Z(n31416) );
  AND U27901 ( .A(n31409), .B(n31416), .Z(n52386) );
  AND U27902 ( .A(n11880), .B(n52386), .Z(n11882) );
  NANDN U27903 ( .A(x[864]), .B(y[864]), .Z(n28182) );
  ANDN U27904 ( .B(y[863]), .A(x[863]), .Z(n52385) );
  ANDN U27905 ( .B(n28182), .A(n52385), .Z(n11881) );
  NANDN U27906 ( .A(n11882), .B(n11881), .Z(n11883) );
  NANDN U27907 ( .A(y[865]), .B(x[865]), .Z(n52873) );
  AND U27908 ( .A(n11883), .B(n52873), .Z(n11884) );
  NAND U27909 ( .A(n52384), .B(n11884), .Z(n11885) );
  ANDN U27910 ( .B(y[865]), .A(x[865]), .Z(n28181) );
  ANDN U27911 ( .B(n11885), .A(n28181), .Z(n11886) );
  NANDN U27912 ( .A(n52383), .B(n11886), .Z(n11887) );
  NAND U27913 ( .A(n52382), .B(n11887), .Z(n11888) );
  NANDN U27914 ( .A(n52381), .B(n11888), .Z(n11889) );
  AND U27915 ( .A(n52876), .B(n11889), .Z(n11890) );
  ANDN U27916 ( .B(y[869]), .A(x[869]), .Z(n31430) );
  NANDN U27917 ( .A(x[870]), .B(y[870]), .Z(n31439) );
  NANDN U27918 ( .A(n31430), .B(n31439), .Z(n52877) );
  OR U27919 ( .A(n11890), .B(n52877), .Z(n11891) );
  NAND U27920 ( .A(n52878), .B(n11891), .Z(n11892) );
  NANDN U27921 ( .A(n52380), .B(n11892), .Z(n11893) );
  NAND U27922 ( .A(n52879), .B(n11893), .Z(n11894) );
  ANDN U27923 ( .B(y[874]), .A(x[874]), .Z(n28180) );
  ANDN U27924 ( .B(n11894), .A(n28180), .Z(n11895) );
  NANDN U27925 ( .A(n31445), .B(n11895), .Z(n11897) );
  NANDN U27926 ( .A(y[874]), .B(x[874]), .Z(n52881) );
  NANDN U27927 ( .A(y[875]), .B(x[875]), .Z(n52883) );
  AND U27928 ( .A(n52881), .B(n52883), .Z(n11896) );
  NAND U27929 ( .A(n11897), .B(n11896), .Z(n11898) );
  ANDN U27930 ( .B(y[876]), .A(x[876]), .Z(n52884) );
  ANDN U27931 ( .B(n11898), .A(n52884), .Z(n11899) );
  NANDN U27932 ( .A(n28179), .B(n11899), .Z(n11900) );
  NAND U27933 ( .A(n52379), .B(n11900), .Z(n11901) );
  NANDN U27934 ( .A(n52378), .B(n11901), .Z(n11902) );
  NAND U27935 ( .A(n52377), .B(n11902), .Z(n11903) );
  NANDN U27936 ( .A(n52886), .B(n11903), .Z(n11904) );
  NANDN U27937 ( .A(y[880]), .B(x[880]), .Z(n28178) );
  NANDN U27938 ( .A(y[881]), .B(x[881]), .Z(n31474) );
  AND U27939 ( .A(n28178), .B(n31474), .Z(n52887) );
  AND U27940 ( .A(n11904), .B(n52887), .Z(n11905) );
  NANDN U27941 ( .A(x[881]), .B(y[881]), .Z(n31469) );
  NANDN U27942 ( .A(x[882]), .B(y[882]), .Z(n28174) );
  NAND U27943 ( .A(n31469), .B(n28174), .Z(n52376) );
  OR U27944 ( .A(n11905), .B(n52376), .Z(n11906) );
  NAND U27945 ( .A(n52888), .B(n11906), .Z(n11907) );
  NANDN U27946 ( .A(n52375), .B(n11907), .Z(n11908) );
  ANDN U27947 ( .B(y[884]), .A(x[884]), .Z(n31480) );
  OR U27948 ( .A(n11908), .B(n31480), .Z(n11909) );
  AND U27949 ( .A(n11910), .B(n11909), .Z(n11911) );
  NOR U27950 ( .A(n31479), .B(n11911), .Z(n11912) );
  NAND U27951 ( .A(n52891), .B(n11912), .Z(n11918) );
  NANDN U27952 ( .A(y[889]), .B(x[889]), .Z(n11914) );
  NANDN U27953 ( .A(y[888]), .B(x[888]), .Z(n11913) );
  AND U27954 ( .A(n11914), .B(n11913), .Z(n31489) );
  NANDN U27955 ( .A(y[887]), .B(x[887]), .Z(n31486) );
  NANDN U27956 ( .A(y[886]), .B(x[886]), .Z(n31483) );
  NAND U27957 ( .A(n31486), .B(n31483), .Z(n11915) );
  NAND U27958 ( .A(n11916), .B(n11915), .Z(n11917) );
  AND U27959 ( .A(n31489), .B(n11917), .Z(n52373) );
  AND U27960 ( .A(n11918), .B(n52373), .Z(n11921) );
  NANDN U27961 ( .A(x[889]), .B(y[889]), .Z(n11920) );
  NANDN U27962 ( .A(x[890]), .B(y[890]), .Z(n11919) );
  NAND U27963 ( .A(n11920), .B(n11919), .Z(n52372) );
  OR U27964 ( .A(n11921), .B(n52372), .Z(n11922) );
  NAND U27965 ( .A(n52371), .B(n11922), .Z(n11923) );
  NANDN U27966 ( .A(n52894), .B(n11923), .Z(n11924) );
  NAND U27967 ( .A(n52895), .B(n11924), .Z(n11925) );
  NANDN U27968 ( .A(n52370), .B(n11925), .Z(n11926) );
  AND U27969 ( .A(n52896), .B(n11926), .Z(n11927) );
  XNOR U27970 ( .A(y[896]), .B(x[896]), .Z(n28171) );
  NANDN U27971 ( .A(x[895]), .B(y[895]), .Z(n28172) );
  NAND U27972 ( .A(n28171), .B(n28172), .Z(n52369) );
  OR U27973 ( .A(n11927), .B(n52369), .Z(n11928) );
  NAND U27974 ( .A(n52897), .B(n11928), .Z(n11929) );
  NANDN U27975 ( .A(n52898), .B(n11929), .Z(n11930) );
  NAND U27976 ( .A(n52899), .B(n11930), .Z(n11931) );
  NANDN U27977 ( .A(n52368), .B(n11931), .Z(n11932) );
  AND U27978 ( .A(n52900), .B(n11932), .Z(n11933) );
  ANDN U27979 ( .B(y[901]), .A(x[901]), .Z(n31527) );
  NANDN U27980 ( .A(x[902]), .B(y[902]), .Z(n28167) );
  NANDN U27981 ( .A(n31527), .B(n28167), .Z(n52367) );
  OR U27982 ( .A(n11933), .B(n52367), .Z(n11934) );
  NAND U27983 ( .A(n52366), .B(n11934), .Z(n11935) );
  NANDN U27984 ( .A(n52901), .B(n11935), .Z(n11936) );
  NAND U27985 ( .A(n52904), .B(n11936), .Z(n11937) );
  NANDN U27986 ( .A(n52365), .B(n11937), .Z(n11938) );
  AND U27987 ( .A(n52905), .B(n11938), .Z(n11939) );
  ANDN U27988 ( .B(y[908]), .A(x[908]), .Z(n31550) );
  NANDN U27989 ( .A(x[907]), .B(y[907]), .Z(n31545) );
  NANDN U27990 ( .A(n31550), .B(n31545), .Z(n52364) );
  OR U27991 ( .A(n11939), .B(n52364), .Z(n11940) );
  NAND U27992 ( .A(n52906), .B(n11940), .Z(n11941) );
  NANDN U27993 ( .A(n52907), .B(n11941), .Z(n11942) );
  NAND U27994 ( .A(n52908), .B(n11942), .Z(n11943) );
  NANDN U27995 ( .A(n52363), .B(n11943), .Z(n11944) );
  AND U27996 ( .A(n52909), .B(n11944), .Z(n11946) );
  XNOR U27997 ( .A(y[914]), .B(x[914]), .Z(n31567) );
  ANDN U27998 ( .B(y[913]), .A(x[913]), .Z(n52910) );
  ANDN U27999 ( .B(n31567), .A(n52910), .Z(n11945) );
  NANDN U28000 ( .A(n11946), .B(n11945), .Z(n11947) );
  AND U28001 ( .A(n11948), .B(n11947), .Z(n11950) );
  NANDN U28002 ( .A(x[915]), .B(y[915]), .Z(n28157) );
  ANDN U28003 ( .B(y[916]), .A(x[916]), .Z(n28156) );
  ANDN U28004 ( .B(n28157), .A(n28156), .Z(n11949) );
  NANDN U28005 ( .A(n11950), .B(n11949), .Z(n11951) );
  AND U28006 ( .A(n52916), .B(n11951), .Z(n11952) );
  NANDN U28007 ( .A(x[917]), .B(y[917]), .Z(n31576) );
  NANDN U28008 ( .A(x[918]), .B(y[918]), .Z(n31582) );
  NAND U28009 ( .A(n31576), .B(n31582), .Z(n52917) );
  OR U28010 ( .A(n11952), .B(n52917), .Z(n11953) );
  NAND U28011 ( .A(n52918), .B(n11953), .Z(n11954) );
  NANDN U28012 ( .A(n52362), .B(n11954), .Z(n11955) );
  NAND U28013 ( .A(n52919), .B(n11955), .Z(n11956) );
  NANDN U28014 ( .A(n52361), .B(n11956), .Z(n11957) );
  AND U28015 ( .A(n52920), .B(n11957), .Z(n11959) );
  NANDN U28016 ( .A(x[924]), .B(y[924]), .Z(n28153) );
  ANDN U28017 ( .B(y[923]), .A(x[923]), .Z(n52921) );
  ANDN U28018 ( .B(n28153), .A(n52921), .Z(n11958) );
  NANDN U28019 ( .A(n11959), .B(n11958), .Z(n11960) );
  AND U28020 ( .A(n11961), .B(n11960), .Z(n11963) );
  NANDN U28021 ( .A(x[926]), .B(y[926]), .Z(n52925) );
  ANDN U28022 ( .B(y[925]), .A(x[925]), .Z(n28152) );
  ANDN U28023 ( .B(n52925), .A(n28152), .Z(n11962) );
  NANDN U28024 ( .A(n11963), .B(n11962), .Z(n11964) );
  AND U28025 ( .A(n52926), .B(n11964), .Z(n11967) );
  NANDN U28026 ( .A(x[927]), .B(y[927]), .Z(n11966) );
  NANDN U28027 ( .A(x[928]), .B(y[928]), .Z(n11965) );
  NAND U28028 ( .A(n11966), .B(n11965), .Z(n31609) );
  OR U28029 ( .A(n11967), .B(n31609), .Z(n11968) );
  NAND U28030 ( .A(n31611), .B(n11968), .Z(n11969) );
  NANDN U28031 ( .A(n28150), .B(n11969), .Z(n11970) );
  NAND U28032 ( .A(n28149), .B(n11970), .Z(n11971) );
  NANDN U28033 ( .A(n52360), .B(n11971), .Z(n11972) );
  AND U28034 ( .A(n52932), .B(n11972), .Z(n11974) );
  ANDN U28035 ( .B(y[933]), .A(x[933]), .Z(n31619) );
  IV U28036 ( .A(n31619), .Z(n52933) );
  ANDN U28037 ( .B(y[934]), .A(x[934]), .Z(n28147) );
  ANDN U28038 ( .B(n52933), .A(n28147), .Z(n11973) );
  NANDN U28039 ( .A(n11974), .B(n11973), .Z(n11975) );
  NANDN U28040 ( .A(y[935]), .B(x[935]), .Z(n52359) );
  AND U28041 ( .A(n11975), .B(n52359), .Z(n11976) );
  NAND U28042 ( .A(n52934), .B(n11976), .Z(n11977) );
  AND U28043 ( .A(n11978), .B(n11977), .Z(n11979) );
  OR U28044 ( .A(n52936), .B(n11979), .Z(n11980) );
  NAND U28045 ( .A(n52937), .B(n11980), .Z(n11981) );
  NANDN U28046 ( .A(n52938), .B(n11981), .Z(n11982) );
  NAND U28047 ( .A(n52939), .B(n11982), .Z(n11983) );
  NANDN U28048 ( .A(n52940), .B(n11983), .Z(n11984) );
  AND U28049 ( .A(n52941), .B(n11984), .Z(n11985) );
  OR U28050 ( .A(n52942), .B(n11985), .Z(n11986) );
  AND U28051 ( .A(n11987), .B(n11986), .Z(n11988) );
  OR U28052 ( .A(n11989), .B(n11988), .Z(n11990) );
  AND U28053 ( .A(n11991), .B(n11990), .Z(n11992) );
  OR U28054 ( .A(n52948), .B(n11992), .Z(n11993) );
  NAND U28055 ( .A(n52949), .B(n11993), .Z(n11994) );
  NANDN U28056 ( .A(n52950), .B(n11994), .Z(n11995) );
  NAND U28057 ( .A(n52951), .B(n11995), .Z(n11996) );
  NANDN U28058 ( .A(n52952), .B(n11996), .Z(n11997) );
  AND U28059 ( .A(n52953), .B(n11997), .Z(n11998) );
  OR U28060 ( .A(n52954), .B(n11998), .Z(n11999) );
  NAND U28061 ( .A(n52955), .B(n11999), .Z(n12000) );
  NANDN U28062 ( .A(n52956), .B(n12000), .Z(n12001) );
  NAND U28063 ( .A(n52957), .B(n12001), .Z(n12002) );
  NANDN U28064 ( .A(n52958), .B(n12002), .Z(n12003) );
  AND U28065 ( .A(n52959), .B(n12003), .Z(n12004) );
  OR U28066 ( .A(n52960), .B(n12004), .Z(n12005) );
  NAND U28067 ( .A(n52962), .B(n12005), .Z(n12006) );
  NANDN U28068 ( .A(n52963), .B(n12006), .Z(n12007) );
  NAND U28069 ( .A(n52964), .B(n12007), .Z(n12008) );
  NANDN U28070 ( .A(n52965), .B(n12008), .Z(n12009) );
  AND U28071 ( .A(n52966), .B(n12009), .Z(n12010) );
  NANDN U28072 ( .A(x[964]), .B(y[964]), .Z(n31717) );
  NAND U28073 ( .A(n12010), .B(n31717), .Z(n12011) );
  NANDN U28074 ( .A(n12012), .B(n12011), .Z(n12013) );
  AND U28075 ( .A(n52969), .B(n12013), .Z(n12014) );
  NANDN U28076 ( .A(x[965]), .B(y[965]), .Z(n31716) );
  NAND U28077 ( .A(n12014), .B(n31716), .Z(n12015) );
  NANDN U28078 ( .A(n52970), .B(n12015), .Z(n12016) );
  AND U28079 ( .A(n52971), .B(n12016), .Z(n12017) );
  OR U28080 ( .A(n52972), .B(n12017), .Z(n12018) );
  NAND U28081 ( .A(n52973), .B(n12018), .Z(n12019) );
  NANDN U28082 ( .A(n52974), .B(n12019), .Z(n12020) );
  NAND U28083 ( .A(n52975), .B(n12020), .Z(n12021) );
  NANDN U28084 ( .A(n52976), .B(n12021), .Z(n12022) );
  AND U28085 ( .A(n52977), .B(n12022), .Z(n12023) );
  NANDN U28086 ( .A(x[974]), .B(y[974]), .Z(n28126) );
  NAND U28087 ( .A(n12023), .B(n28126), .Z(n12024) );
  NANDN U28088 ( .A(n12025), .B(n12024), .Z(n12026) );
  AND U28089 ( .A(n52982), .B(n12026), .Z(n12027) );
  NANDN U28090 ( .A(x[975]), .B(y[975]), .Z(n28125) );
  NAND U28091 ( .A(n12027), .B(n28125), .Z(n12028) );
  NANDN U28092 ( .A(n52983), .B(n12028), .Z(n12029) );
  AND U28093 ( .A(n52984), .B(n12029), .Z(n12030) );
  ANDN U28094 ( .B(x[978]), .A(y[978]), .Z(n31755) );
  ANDN U28095 ( .B(x[979]), .A(y[979]), .Z(n31765) );
  OR U28096 ( .A(n31755), .B(n31765), .Z(n52985) );
  OR U28097 ( .A(n12030), .B(n52985), .Z(n12031) );
  AND U28098 ( .A(n52986), .B(n12031), .Z(n12032) );
  OR U28099 ( .A(n52987), .B(n12032), .Z(n12033) );
  NAND U28100 ( .A(n52988), .B(n12033), .Z(n12034) );
  NANDN U28101 ( .A(n52989), .B(n12034), .Z(n12035) );
  ANDN U28102 ( .B(y[983]), .A(x[983]), .Z(n52990) );
  ANDN U28103 ( .B(n12035), .A(n52990), .Z(n12036) );
  NAND U28104 ( .A(n52992), .B(n12036), .Z(n12037) );
  NANDN U28105 ( .A(n12038), .B(n12037), .Z(n12039) );
  NAND U28106 ( .A(n52994), .B(n12039), .Z(n12040) );
  NANDN U28107 ( .A(n52995), .B(n12040), .Z(n12041) );
  AND U28108 ( .A(n52996), .B(n12041), .Z(n12042) );
  OR U28109 ( .A(n52997), .B(n12042), .Z(n12043) );
  NAND U28110 ( .A(n52998), .B(n12043), .Z(n12044) );
  NANDN U28111 ( .A(n53000), .B(n12044), .Z(n12045) );
  NAND U28112 ( .A(n53001), .B(n12045), .Z(n12046) );
  NANDN U28113 ( .A(n53002), .B(n12046), .Z(n12047) );
  ANDN U28114 ( .B(y[993]), .A(x[993]), .Z(n53003) );
  ANDN U28115 ( .B(n12047), .A(n53003), .Z(n12048) );
  NANDN U28116 ( .A(x[994]), .B(y[994]), .Z(n31815) );
  NAND U28117 ( .A(n12048), .B(n31815), .Z(n12049) );
  NANDN U28118 ( .A(n12050), .B(n12049), .Z(n12051) );
  AND U28119 ( .A(n53005), .B(n12051), .Z(n12052) );
  NANDN U28120 ( .A(x[995]), .B(y[995]), .Z(n31814) );
  NAND U28121 ( .A(n12052), .B(n31814), .Z(n12053) );
  NANDN U28122 ( .A(n53006), .B(n12053), .Z(n12054) );
  AND U28123 ( .A(n53007), .B(n12054), .Z(n12055) );
  OR U28124 ( .A(n53008), .B(n12055), .Z(n12056) );
  NAND U28125 ( .A(n53009), .B(n12056), .Z(n12057) );
  NANDN U28126 ( .A(n53010), .B(n12057), .Z(n12058) );
  NAND U28127 ( .A(n53011), .B(n12058), .Z(n12059) );
  NANDN U28128 ( .A(n53012), .B(n12059), .Z(n12060) );
  AND U28129 ( .A(n53013), .B(n12060), .Z(n12061) );
  OR U28130 ( .A(n53014), .B(n12061), .Z(n12062) );
  NAND U28131 ( .A(n53016), .B(n12062), .Z(n12063) );
  NANDN U28132 ( .A(n53017), .B(n12063), .Z(n12064) );
  NAND U28133 ( .A(n53018), .B(n12064), .Z(n12065) );
  NANDN U28134 ( .A(n53019), .B(n12065), .Z(n12066) );
  AND U28135 ( .A(n53020), .B(n12066), .Z(n12069) );
  NANDN U28136 ( .A(y[1010]), .B(x[1010]), .Z(n12068) );
  NANDN U28137 ( .A(y[1011]), .B(x[1011]), .Z(n12067) );
  NAND U28138 ( .A(n12068), .B(n12067), .Z(n53021) );
  OR U28139 ( .A(n12069), .B(n53021), .Z(n12070) );
  AND U28140 ( .A(n53022), .B(n12070), .Z(n12071) );
  ANDN U28141 ( .B(x[1012]), .A(y[1012]), .Z(n31866) );
  ANDN U28142 ( .B(x[1013]), .A(y[1013]), .Z(n31869) );
  NOR U28143 ( .A(n31866), .B(n31869), .Z(n53023) );
  NANDN U28144 ( .A(n12071), .B(n53023), .Z(n12072) );
  NAND U28145 ( .A(n12073), .B(n12072), .Z(n12074) );
  NANDN U28146 ( .A(y[1015]), .B(x[1015]), .Z(n28112) );
  AND U28147 ( .A(n12074), .B(n28112), .Z(n12075) );
  NAND U28148 ( .A(n31870), .B(n12075), .Z(n12076) );
  NANDN U28149 ( .A(n28111), .B(n12076), .Z(n12077) );
  ANDN U28150 ( .B(y[1015]), .A(x[1015]), .Z(n28113) );
  OR U28151 ( .A(n12077), .B(n28113), .Z(n12078) );
  NAND U28152 ( .A(n53029), .B(n12078), .Z(n12079) );
  NANDN U28153 ( .A(n52352), .B(n12079), .Z(n12080) );
  NAND U28154 ( .A(n53030), .B(n12080), .Z(n12081) );
  NAND U28155 ( .A(n53031), .B(n12081), .Z(n12082) );
  NANDN U28156 ( .A(n53032), .B(n12082), .Z(n12083) );
  NAND U28157 ( .A(n53033), .B(n12083), .Z(n12084) );
  NANDN U28158 ( .A(n53035), .B(n12084), .Z(n12085) );
  ANDN U28159 ( .B(y[1023]), .A(x[1023]), .Z(n53036) );
  ANDN U28160 ( .B(n12085), .A(n53036), .Z(n12086) );
  NANDN U28161 ( .A(x[1024]), .B(y[1024]), .Z(n28107) );
  NAND U28162 ( .A(n12086), .B(n28107), .Z(n12087) );
  NANDN U28163 ( .A(y[1025]), .B(x[1025]), .Z(n53039) );
  AND U28164 ( .A(n12087), .B(n53039), .Z(n12088) );
  NAND U28165 ( .A(n53037), .B(n12088), .Z(n12089) );
  NANDN U28166 ( .A(x[1025]), .B(y[1025]), .Z(n28106) );
  AND U28167 ( .A(n12089), .B(n28106), .Z(n12090) );
  NANDN U28168 ( .A(n53040), .B(n12090), .Z(n12091) );
  NANDN U28169 ( .A(n53041), .B(n12091), .Z(n12092) );
  NAND U28170 ( .A(n53042), .B(n12092), .Z(n12093) );
  NANDN U28171 ( .A(n53043), .B(n12093), .Z(n12094) );
  AND U28172 ( .A(n53044), .B(n12094), .Z(n12095) );
  OR U28173 ( .A(n53045), .B(n12095), .Z(n12096) );
  NAND U28174 ( .A(n53046), .B(n12096), .Z(n12097) );
  NANDN U28175 ( .A(n53047), .B(n12097), .Z(n12098) );
  NANDN U28176 ( .A(x[1034]), .B(y[1034]), .Z(n31931) );
  AND U28177 ( .A(n12098), .B(n31931), .Z(n12099) );
  NANDN U28178 ( .A(n53048), .B(n12099), .Z(n12100) );
  NANDN U28179 ( .A(n12101), .B(n12100), .Z(n12102) );
  AND U28180 ( .A(n53052), .B(n12102), .Z(n12103) );
  NAND U28181 ( .A(n31930), .B(n12103), .Z(n12104) );
  NANDN U28182 ( .A(n53053), .B(n12104), .Z(n12105) );
  NAND U28183 ( .A(n53055), .B(n12105), .Z(n12106) );
  NANDN U28184 ( .A(n53056), .B(n12106), .Z(n12107) );
  AND U28185 ( .A(n53057), .B(n12107), .Z(n12108) );
  OR U28186 ( .A(n53058), .B(n12108), .Z(n12109) );
  NAND U28187 ( .A(n53059), .B(n12109), .Z(n12110) );
  NANDN U28188 ( .A(n53060), .B(n12110), .Z(n12111) );
  NANDN U28189 ( .A(x[1043]), .B(y[1043]), .Z(n53061) );
  AND U28190 ( .A(n12111), .B(n53061), .Z(n12112) );
  NAND U28191 ( .A(n53063), .B(n12112), .Z(n12113) );
  NANDN U28192 ( .A(n12114), .B(n12113), .Z(n12115) );
  NAND U28193 ( .A(n53065), .B(n12115), .Z(n12116) );
  NAND U28194 ( .A(n52351), .B(n12116), .Z(n12117) );
  NANDN U28195 ( .A(n53066), .B(n12117), .Z(n12118) );
  NANDN U28196 ( .A(n53067), .B(n12118), .Z(n12119) );
  AND U28197 ( .A(n53068), .B(n12119), .Z(n12120) );
  NANDN U28198 ( .A(y[1050]), .B(x[1050]), .Z(n31983) );
  ANDN U28199 ( .B(x[1051]), .A(y[1051]), .Z(n31993) );
  ANDN U28200 ( .B(n31983), .A(n31993), .Z(n53069) );
  NANDN U28201 ( .A(n12120), .B(n53069), .Z(n12121) );
  NANDN U28202 ( .A(n52350), .B(n12121), .Z(n12122) );
  AND U28203 ( .A(n53071), .B(n12122), .Z(n12123) );
  NANDN U28204 ( .A(x[1053]), .B(y[1053]), .Z(n31995) );
  NANDN U28205 ( .A(x[1054]), .B(y[1054]), .Z(n32002) );
  NAND U28206 ( .A(n31995), .B(n32002), .Z(n53072) );
  OR U28207 ( .A(n12123), .B(n53072), .Z(n12124) );
  NAND U28208 ( .A(n53074), .B(n12124), .Z(n12125) );
  NANDN U28209 ( .A(n52349), .B(n12125), .Z(n12126) );
  NAND U28210 ( .A(n53075), .B(n12126), .Z(n12127) );
  NANDN U28211 ( .A(n52348), .B(n12127), .Z(n12128) );
  AND U28212 ( .A(n53076), .B(n12128), .Z(n12129) );
  NANDN U28213 ( .A(x[1059]), .B(y[1059]), .Z(n32017) );
  NANDN U28214 ( .A(x[1060]), .B(y[1060]), .Z(n32024) );
  NAND U28215 ( .A(n32017), .B(n32024), .Z(n53077) );
  OR U28216 ( .A(n12129), .B(n53077), .Z(n12130) );
  NAND U28217 ( .A(n53078), .B(n12130), .Z(n12131) );
  NANDN U28218 ( .A(n52347), .B(n12131), .Z(n12132) );
  NAND U28219 ( .A(n53079), .B(n12132), .Z(n12133) );
  NANDN U28220 ( .A(x[1064]), .B(y[1064]), .Z(n28095) );
  AND U28221 ( .A(n12133), .B(n28095), .Z(n12134) );
  NANDN U28222 ( .A(n53080), .B(n12134), .Z(n12135) );
  NANDN U28223 ( .A(n12136), .B(n12135), .Z(n12137) );
  NANDN U28224 ( .A(x[1065]), .B(y[1065]), .Z(n28094) );
  AND U28225 ( .A(n12137), .B(n28094), .Z(n12138) );
  NAND U28226 ( .A(n28093), .B(n12138), .Z(n12139) );
  NANDN U28227 ( .A(n53086), .B(n12139), .Z(n12140) );
  NANDN U28228 ( .A(x[1067]), .B(y[1067]), .Z(n32042) );
  AND U28229 ( .A(n12140), .B(n32042), .Z(n12141) );
  NAND U28230 ( .A(n28091), .B(n12141), .Z(n12142) );
  NANDN U28231 ( .A(n28092), .B(n12142), .Z(n12143) );
  ANDN U28232 ( .B(x[1069]), .A(y[1069]), .Z(n28088) );
  OR U28233 ( .A(n12143), .B(n28088), .Z(n12144) );
  AND U28234 ( .A(n12145), .B(n12144), .Z(n12147) );
  NANDN U28235 ( .A(y[1071]), .B(x[1071]), .Z(n53092) );
  NANDN U28236 ( .A(y[1070]), .B(x[1070]), .Z(n28089) );
  AND U28237 ( .A(n53092), .B(n28089), .Z(n12146) );
  NANDN U28238 ( .A(n12147), .B(n12146), .Z(n12148) );
  ANDN U28239 ( .B(y[1072]), .A(x[1072]), .Z(n53093) );
  ANDN U28240 ( .B(n12148), .A(n53093), .Z(n12149) );
  NANDN U28241 ( .A(x[1071]), .B(y[1071]), .Z(n32049) );
  NAND U28242 ( .A(n12149), .B(n32049), .Z(n12150) );
  NANDN U28243 ( .A(n53094), .B(n12150), .Z(n12151) );
  AND U28244 ( .A(n53095), .B(n12151), .Z(n12152) );
  OR U28245 ( .A(n53096), .B(n12152), .Z(n12153) );
  NAND U28246 ( .A(n53097), .B(n12153), .Z(n12154) );
  NANDN U28247 ( .A(n53098), .B(n12154), .Z(n12155) );
  NAND U28248 ( .A(n53099), .B(n12155), .Z(n12156) );
  NANDN U28249 ( .A(n53100), .B(n12156), .Z(n12157) );
  AND U28250 ( .A(n53101), .B(n12157), .Z(n12158) );
  OR U28251 ( .A(n53102), .B(n12158), .Z(n12159) );
  NAND U28252 ( .A(n53104), .B(n12159), .Z(n12160) );
  NANDN U28253 ( .A(n53105), .B(n12160), .Z(n12161) );
  NAND U28254 ( .A(n53106), .B(n12161), .Z(n12162) );
  NANDN U28255 ( .A(n53107), .B(n12162), .Z(n12163) );
  AND U28256 ( .A(n53108), .B(n12163), .Z(n12164) );
  OR U28257 ( .A(n53109), .B(n12164), .Z(n12165) );
  NAND U28258 ( .A(n53110), .B(n12165), .Z(n12166) );
  NANDN U28259 ( .A(n53111), .B(n12166), .Z(n12167) );
  NAND U28260 ( .A(n53112), .B(n12167), .Z(n12168) );
  NAND U28261 ( .A(n53113), .B(n12168), .Z(n12169) );
  NANDN U28262 ( .A(n53114), .B(n12169), .Z(n12170) );
  NAND U28263 ( .A(n53115), .B(n12170), .Z(n12171) );
  NANDN U28264 ( .A(x[1093]), .B(y[1093]), .Z(n53116) );
  AND U28265 ( .A(n12171), .B(n53116), .Z(n12172) );
  NAND U28266 ( .A(n52346), .B(n12172), .Z(n12173) );
  NANDN U28267 ( .A(n12174), .B(n12173), .Z(n12175) );
  NAND U28268 ( .A(n53119), .B(n12175), .Z(n12176) );
  NAND U28269 ( .A(n53120), .B(n12176), .Z(n12177) );
  NANDN U28270 ( .A(n53122), .B(n12177), .Z(n12178) );
  NAND U28271 ( .A(n53124), .B(n12178), .Z(n12179) );
  NANDN U28272 ( .A(n53126), .B(n12179), .Z(n12180) );
  AND U28273 ( .A(n53128), .B(n12180), .Z(n12181) );
  OR U28274 ( .A(n53130), .B(n12181), .Z(n12182) );
  NAND U28275 ( .A(n53132), .B(n12182), .Z(n12183) );
  NANDN U28276 ( .A(n53134), .B(n12183), .Z(n12184) );
  NAND U28277 ( .A(n53136), .B(n12184), .Z(n12185) );
  NANDN U28278 ( .A(n53138), .B(n12185), .Z(n12186) );
  AND U28279 ( .A(n53140), .B(n12186), .Z(n12187) );
  OR U28280 ( .A(n53142), .B(n12187), .Z(n12188) );
  NAND U28281 ( .A(n53144), .B(n12188), .Z(n12189) );
  NANDN U28282 ( .A(n53146), .B(n12189), .Z(n12190) );
  NANDN U28283 ( .A(x[1110]), .B(y[1110]), .Z(n28066) );
  NANDN U28284 ( .A(n12190), .B(n28066), .Z(n12191) );
  AND U28285 ( .A(n28064), .B(n12191), .Z(n12192) );
  NANDN U28286 ( .A(y[1110]), .B(x[1110]), .Z(n53147) );
  NAND U28287 ( .A(n12192), .B(n53147), .Z(n12193) );
  ANDN U28288 ( .B(y[1111]), .A(x[1111]), .Z(n28065) );
  ANDN U28289 ( .B(n12193), .A(n28065), .Z(n12194) );
  NANDN U28290 ( .A(n28063), .B(n12194), .Z(n12196) );
  NANDN U28291 ( .A(y[1112]), .B(x[1112]), .Z(n12195) );
  AND U28292 ( .A(n12196), .B(n12195), .Z(n12197) );
  NAND U28293 ( .A(n53156), .B(n12197), .Z(n12198) );
  NANDN U28294 ( .A(n53158), .B(n12198), .Z(n12199) );
  NAND U28295 ( .A(n53160), .B(n12199), .Z(n12200) );
  NANDN U28296 ( .A(n52345), .B(n12200), .Z(n12201) );
  NANDN U28297 ( .A(y[1116]), .B(x[1116]), .Z(n32193) );
  NANDN U28298 ( .A(y[1117]), .B(x[1117]), .Z(n32199) );
  AND U28299 ( .A(n32193), .B(n32199), .Z(n52344) );
  AND U28300 ( .A(n12201), .B(n52344), .Z(n12202) );
  ANDN U28301 ( .B(y[1117]), .A(x[1117]), .Z(n32195) );
  ANDN U28302 ( .B(y[1118]), .A(x[1118]), .Z(n32204) );
  OR U28303 ( .A(n32195), .B(n32204), .Z(n52343) );
  OR U28304 ( .A(n12202), .B(n52343), .Z(n12203) );
  NAND U28305 ( .A(n52342), .B(n12203), .Z(n12204) );
  NANDN U28306 ( .A(n53163), .B(n12204), .Z(n12205) );
  ANDN U28307 ( .B(y[1120]), .A(x[1120]), .Z(n28060) );
  OR U28308 ( .A(n12205), .B(n28060), .Z(n12206) );
  AND U28309 ( .A(n12207), .B(n12206), .Z(n12209) );
  ANDN U28310 ( .B(y[1122]), .A(x[1122]), .Z(n32213) );
  IV U28311 ( .A(n32213), .Z(n53167) );
  ANDN U28312 ( .B(y[1121]), .A(x[1121]), .Z(n28061) );
  ANDN U28313 ( .B(n53167), .A(n28061), .Z(n12208) );
  NANDN U28314 ( .A(n12209), .B(n12208), .Z(n12210) );
  AND U28315 ( .A(n53168), .B(n12210), .Z(n12211) );
  ANDN U28316 ( .B(y[1123]), .A(x[1123]), .Z(n32215) );
  NANDN U28317 ( .A(x[1124]), .B(y[1124]), .Z(n28059) );
  NANDN U28318 ( .A(n32215), .B(n28059), .Z(n52341) );
  OR U28319 ( .A(n12211), .B(n52341), .Z(n12212) );
  NAND U28320 ( .A(n52340), .B(n12212), .Z(n12213) );
  NANDN U28321 ( .A(n53169), .B(n12213), .Z(n12214) );
  NAND U28322 ( .A(n53172), .B(n12214), .Z(n12215) );
  NANDN U28323 ( .A(n52339), .B(n12215), .Z(n12216) );
  NANDN U28324 ( .A(y[1128]), .B(x[1128]), .Z(n28056) );
  NANDN U28325 ( .A(y[1129]), .B(x[1129]), .Z(n32234) );
  AND U28326 ( .A(n28056), .B(n32234), .Z(n52338) );
  AND U28327 ( .A(n12216), .B(n52338), .Z(n12217) );
  ANDN U28328 ( .B(y[1130]), .A(x[1130]), .Z(n32240) );
  NANDN U28329 ( .A(x[1129]), .B(y[1129]), .Z(n28054) );
  NANDN U28330 ( .A(n32240), .B(n28054), .Z(n52337) );
  OR U28331 ( .A(n12217), .B(n52337), .Z(n12218) );
  NAND U28332 ( .A(n52336), .B(n12218), .Z(n12219) );
  NANDN U28333 ( .A(n53174), .B(n12219), .Z(n12220) );
  NAND U28334 ( .A(n53175), .B(n12220), .Z(n12221) );
  NANDN U28335 ( .A(n52335), .B(n12221), .Z(n12222) );
  AND U28336 ( .A(n53176), .B(n12222), .Z(n12223) );
  ANDN U28337 ( .B(y[1135]), .A(x[1135]), .Z(n32251) );
  NANDN U28338 ( .A(x[1136]), .B(y[1136]), .Z(n28049) );
  NANDN U28339 ( .A(n32251), .B(n28049), .Z(n52334) );
  OR U28340 ( .A(n12223), .B(n52334), .Z(n12224) );
  NAND U28341 ( .A(n53177), .B(n12224), .Z(n12225) );
  NANDN U28342 ( .A(n53178), .B(n12225), .Z(n12226) );
  NAND U28343 ( .A(n53181), .B(n12226), .Z(n12227) );
  NANDN U28344 ( .A(n52333), .B(n12227), .Z(n12229) );
  NANDN U28345 ( .A(y[1140]), .B(x[1140]), .Z(n12228) );
  NANDN U28346 ( .A(y[1141]), .B(x[1141]), .Z(n32274) );
  AND U28347 ( .A(n12228), .B(n32274), .Z(n52332) );
  AND U28348 ( .A(n12229), .B(n52332), .Z(n12230) );
  ANDN U28349 ( .B(y[1141]), .A(x[1141]), .Z(n28046) );
  XNOR U28350 ( .A(y[1142]), .B(x[1142]), .Z(n32275) );
  NANDN U28351 ( .A(n28046), .B(n32275), .Z(n52331) );
  OR U28352 ( .A(n12230), .B(n52331), .Z(n12231) );
  NAND U28353 ( .A(n52330), .B(n12231), .Z(n12232) );
  NANDN U28354 ( .A(n53182), .B(n12232), .Z(n12233) );
  NAND U28355 ( .A(n53183), .B(n12233), .Z(n12234) );
  AND U28356 ( .A(n12235), .B(n12234), .Z(n12237) );
  NANDN U28357 ( .A(y[1146]), .B(x[1146]), .Z(n53185) );
  NANDN U28358 ( .A(y[1147]), .B(x[1147]), .Z(n53187) );
  AND U28359 ( .A(n53185), .B(n53187), .Z(n12236) );
  NANDN U28360 ( .A(n12237), .B(n12236), .Z(n12238) );
  ANDN U28361 ( .B(y[1148]), .A(x[1148]), .Z(n53188) );
  ANDN U28362 ( .B(n12238), .A(n53188), .Z(n12239) );
  NANDN U28363 ( .A(x[1147]), .B(y[1147]), .Z(n28044) );
  NAND U28364 ( .A(n12239), .B(n28044), .Z(n12240) );
  NANDN U28365 ( .A(n53190), .B(n12240), .Z(n12241) );
  AND U28366 ( .A(n53191), .B(n12241), .Z(n12242) );
  OR U28367 ( .A(n53192), .B(n12242), .Z(n12243) );
  NAND U28368 ( .A(n53193), .B(n12243), .Z(n12244) );
  NANDN U28369 ( .A(n53194), .B(n12244), .Z(n12245) );
  NAND U28370 ( .A(n53195), .B(n12245), .Z(n12246) );
  NANDN U28371 ( .A(n53196), .B(n12246), .Z(n12247) );
  AND U28372 ( .A(n53197), .B(n12247), .Z(n12248) );
  OR U28373 ( .A(n53198), .B(n12248), .Z(n12249) );
  NAND U28374 ( .A(n53199), .B(n12249), .Z(n12250) );
  NANDN U28375 ( .A(n53200), .B(n12250), .Z(n12251) );
  NANDN U28376 ( .A(n52329), .B(n12251), .Z(n12252) );
  AND U28377 ( .A(n53201), .B(n12252), .Z(n12254) );
  NANDN U28378 ( .A(x[1162]), .B(y[1162]), .Z(n28032) );
  ANDN U28379 ( .B(y[1161]), .A(x[1161]), .Z(n28033) );
  ANDN U28380 ( .B(n28032), .A(n28033), .Z(n12253) );
  NANDN U28381 ( .A(n12254), .B(n12253), .Z(n12255) );
  NANDN U28382 ( .A(n53203), .B(n12255), .Z(n12256) );
  ANDN U28383 ( .B(x[1163]), .A(y[1163]), .Z(n28029) );
  OR U28384 ( .A(n12256), .B(n28029), .Z(n12257) );
  AND U28385 ( .A(n53206), .B(n12257), .Z(n12258) );
  NANDN U28386 ( .A(n28031), .B(n12258), .Z(n12259) );
  AND U28387 ( .A(n12260), .B(n12259), .Z(n12262) );
  NANDN U28388 ( .A(x[1165]), .B(y[1165]), .Z(n32342) );
  XNOR U28389 ( .A(x[1166]), .B(y[1166]), .Z(n12261) );
  NAND U28390 ( .A(n32342), .B(n12261), .Z(n52328) );
  OR U28391 ( .A(n12262), .B(n52328), .Z(n12263) );
  NAND U28392 ( .A(n53210), .B(n12263), .Z(n12264) );
  NANDN U28393 ( .A(n52327), .B(n12264), .Z(n12265) );
  NAND U28394 ( .A(n53211), .B(n12265), .Z(n12266) );
  NAND U28395 ( .A(n53212), .B(n12266), .Z(n12267) );
  NANDN U28396 ( .A(n53213), .B(n12267), .Z(n12268) );
  ANDN U28397 ( .B(y[1171]), .A(x[1171]), .Z(n53214) );
  ANDN U28398 ( .B(n12268), .A(n53214), .Z(n12269) );
  NAND U28399 ( .A(n28024), .B(n12269), .Z(n12270) );
  NAND U28400 ( .A(n53217), .B(n12270), .Z(n12271) );
  NANDN U28401 ( .A(y[1172]), .B(x[1172]), .Z(n53215) );
  NANDN U28402 ( .A(n12271), .B(n53215), .Z(n12272) );
  AND U28403 ( .A(n12273), .B(n12272), .Z(n12274) );
  OR U28404 ( .A(n53219), .B(n12274), .Z(n12275) );
  NAND U28405 ( .A(n53220), .B(n12275), .Z(n12276) );
  NANDN U28406 ( .A(n53221), .B(n12276), .Z(n12277) );
  NAND U28407 ( .A(n53222), .B(n12277), .Z(n12278) );
  NANDN U28408 ( .A(n53223), .B(n12278), .Z(n12279) );
  AND U28409 ( .A(n53224), .B(n12279), .Z(n12280) );
  OR U28410 ( .A(n53225), .B(n12280), .Z(n12281) );
  NAND U28411 ( .A(n53227), .B(n12281), .Z(n12282) );
  NANDN U28412 ( .A(n52326), .B(n12282), .Z(n12283) );
  NAND U28413 ( .A(n53228), .B(n12283), .Z(n12284) );
  NAND U28414 ( .A(n53229), .B(n12284), .Z(n12285) );
  NANDN U28415 ( .A(n53230), .B(n12285), .Z(n12286) );
  ANDN U28416 ( .B(x[1186]), .A(y[1186]), .Z(n53231) );
  ANDN U28417 ( .B(n12286), .A(n53231), .Z(n12287) );
  NAND U28418 ( .A(n28014), .B(n12287), .Z(n12288) );
  NAND U28419 ( .A(n53232), .B(n12288), .Z(n12289) );
  ANDN U28420 ( .B(y[1188]), .A(x[1188]), .Z(n28011) );
  OR U28421 ( .A(n12289), .B(n28011), .Z(n12290) );
  AND U28422 ( .A(n28013), .B(n12290), .Z(n12291) );
  NANDN U28423 ( .A(n32413), .B(n12291), .Z(n12292) );
  AND U28424 ( .A(n12293), .B(n12292), .Z(n12295) );
  ANDN U28425 ( .B(x[1191]), .A(y[1191]), .Z(n32422) );
  IV U28426 ( .A(n32422), .Z(n53236) );
  ANDN U28427 ( .B(x[1190]), .A(y[1190]), .Z(n32414) );
  ANDN U28428 ( .B(n53236), .A(n32414), .Z(n12294) );
  NANDN U28429 ( .A(n12295), .B(n12294), .Z(n12296) );
  NANDN U28430 ( .A(x[1191]), .B(y[1191]), .Z(n32417) );
  NANDN U28431 ( .A(x[1192]), .B(y[1192]), .Z(n32423) );
  AND U28432 ( .A(n32417), .B(n32423), .Z(n52324) );
  AND U28433 ( .A(n12296), .B(n52324), .Z(n12297) );
  ANDN U28434 ( .B(x[1192]), .A(y[1192]), .Z(n32419) );
  ANDN U28435 ( .B(x[1193]), .A(y[1193]), .Z(n32429) );
  OR U28436 ( .A(n32419), .B(n32429), .Z(n53237) );
  OR U28437 ( .A(n12297), .B(n53237), .Z(n12298) );
  NAND U28438 ( .A(n53238), .B(n12298), .Z(n12299) );
  NANDN U28439 ( .A(n52323), .B(n12299), .Z(n12300) );
  NANDN U28440 ( .A(n53241), .B(n12300), .Z(n12301) );
  AND U28441 ( .A(n53242), .B(n12301), .Z(n12303) );
  ANDN U28442 ( .B(y[1197]), .A(x[1197]), .Z(n52322) );
  ANDN U28443 ( .B(y[1198]), .A(x[1198]), .Z(n28007) );
  NOR U28444 ( .A(n52322), .B(n28007), .Z(n12302) );
  NANDN U28445 ( .A(n12303), .B(n12302), .Z(n12304) );
  NAND U28446 ( .A(n52321), .B(n12304), .Z(n12305) );
  NAND U28447 ( .A(n53243), .B(n12305), .Z(n12306) );
  NANDN U28448 ( .A(n53244), .B(n12306), .Z(n12307) );
  ANDN U28449 ( .B(y[1201]), .A(x[1201]), .Z(n53246) );
  ANDN U28450 ( .B(n12307), .A(n53246), .Z(n12308) );
  XNOR U28451 ( .A(x[1202]), .B(y[1202]), .Z(n32451) );
  NAND U28452 ( .A(n12308), .B(n32451), .Z(n12309) );
  NANDN U28453 ( .A(n53247), .B(n12309), .Z(n12310) );
  NAND U28454 ( .A(n53248), .B(n12310), .Z(n12311) );
  NAND U28455 ( .A(n53249), .B(n12311), .Z(n12312) );
  NANDN U28456 ( .A(n53250), .B(n12312), .Z(n12313) );
  NAND U28457 ( .A(n53251), .B(n12313), .Z(n12314) );
  NANDN U28458 ( .A(n52319), .B(n12314), .Z(n12315) );
  AND U28459 ( .A(n53254), .B(n12315), .Z(n12317) );
  NANDN U28460 ( .A(x[1209]), .B(y[1209]), .Z(n32476) );
  XNOR U28461 ( .A(x[1210]), .B(y[1210]), .Z(n12316) );
  NAND U28462 ( .A(n32476), .B(n12316), .Z(n52318) );
  OR U28463 ( .A(n12317), .B(n52318), .Z(n12318) );
  NAND U28464 ( .A(n53255), .B(n12318), .Z(n12319) );
  NANDN U28465 ( .A(n53256), .B(n12319), .Z(n12320) );
  NANDN U28466 ( .A(y[1212]), .B(x[1212]), .Z(n32489) );
  AND U28467 ( .A(n12320), .B(n32489), .Z(n12321) );
  NAND U28468 ( .A(n28001), .B(n12321), .Z(n12322) );
  NANDN U28469 ( .A(n28003), .B(n12322), .Z(n12323) );
  ANDN U28470 ( .B(y[1214]), .A(x[1214]), .Z(n27998) );
  OR U28471 ( .A(n12323), .B(n27998), .Z(n12324) );
  NAND U28472 ( .A(n12325), .B(n12324), .Z(n12326) );
  NANDN U28473 ( .A(x[1215]), .B(y[1215]), .Z(n27999) );
  AND U28474 ( .A(n12326), .B(n27999), .Z(n12327) );
  NAND U28475 ( .A(n27995), .B(n12327), .Z(n12328) );
  NANDN U28476 ( .A(n53263), .B(n12328), .Z(n12329) );
  ANDN U28477 ( .B(x[1216]), .A(y[1216]), .Z(n27996) );
  OR U28478 ( .A(n12329), .B(n27996), .Z(n12330) );
  AND U28479 ( .A(n53264), .B(n12330), .Z(n12331) );
  NANDN U28480 ( .A(x[1217]), .B(y[1217]), .Z(n27994) );
  NAND U28481 ( .A(n12331), .B(n27994), .Z(n12332) );
  NANDN U28482 ( .A(n53265), .B(n12332), .Z(n12333) );
  AND U28483 ( .A(n53266), .B(n12333), .Z(n12334) );
  OR U28484 ( .A(n53267), .B(n12334), .Z(n12335) );
  NAND U28485 ( .A(n53268), .B(n12335), .Z(n12336) );
  NANDN U28486 ( .A(n53269), .B(n12336), .Z(n12337) );
  NANDN U28487 ( .A(x[1224]), .B(y[1224]), .Z(n27992) );
  AND U28488 ( .A(n12337), .B(n27992), .Z(n12338) );
  NANDN U28489 ( .A(n53270), .B(n12338), .Z(n12339) );
  NANDN U28490 ( .A(n12340), .B(n12339), .Z(n12341) );
  NANDN U28491 ( .A(x[1225]), .B(y[1225]), .Z(n27991) );
  AND U28492 ( .A(n12341), .B(n27991), .Z(n12342) );
  NANDN U28493 ( .A(n53274), .B(n12342), .Z(n12343) );
  NANDN U28494 ( .A(n53275), .B(n12343), .Z(n12344) );
  NAND U28495 ( .A(n53276), .B(n12344), .Z(n12345) );
  NANDN U28496 ( .A(n53277), .B(n12345), .Z(n12346) );
  AND U28497 ( .A(n53278), .B(n12346), .Z(n12347) );
  NANDN U28498 ( .A(y[1230]), .B(x[1230]), .Z(n32535) );
  NANDN U28499 ( .A(y[1231]), .B(x[1231]), .Z(n27988) );
  NAND U28500 ( .A(n32535), .B(n27988), .Z(n53279) );
  OR U28501 ( .A(n12347), .B(n53279), .Z(n12348) );
  NAND U28502 ( .A(n53280), .B(n12348), .Z(n12349) );
  NANDN U28503 ( .A(n52315), .B(n12349), .Z(n12350) );
  NAND U28504 ( .A(n53281), .B(n12350), .Z(n12351) );
  NANDN U28505 ( .A(n52314), .B(n12351), .Z(n12352) );
  AND U28506 ( .A(n53283), .B(n12352), .Z(n12353) );
  NANDN U28507 ( .A(y[1236]), .B(x[1236]), .Z(n32555) );
  NANDN U28508 ( .A(y[1237]), .B(x[1237]), .Z(n32563) );
  NAND U28509 ( .A(n32555), .B(n32563), .Z(n53284) );
  OR U28510 ( .A(n12353), .B(n53284), .Z(n12354) );
  NAND U28511 ( .A(n53285), .B(n12354), .Z(n12355) );
  NANDN U28512 ( .A(n32562), .B(n12355), .Z(n12356) );
  ANDN U28513 ( .B(x[1239]), .A(y[1239]), .Z(n27983) );
  OR U28514 ( .A(n12356), .B(n27983), .Z(n12357) );
  AND U28515 ( .A(n32572), .B(n12357), .Z(n12358) );
  NAND U28516 ( .A(n32568), .B(n12358), .Z(n12359) );
  ANDN U28517 ( .B(x[1241]), .A(y[1241]), .Z(n27981) );
  ANDN U28518 ( .B(n12359), .A(n27981), .Z(n12360) );
  NAND U28519 ( .A(n27984), .B(n12360), .Z(n12361) );
  NANDN U28520 ( .A(x[1242]), .B(y[1242]), .Z(n53291) );
  AND U28521 ( .A(n12361), .B(n53291), .Z(n12362) );
  NAND U28522 ( .A(n32571), .B(n12362), .Z(n12363) );
  NAND U28523 ( .A(n27982), .B(n12363), .Z(n12366) );
  NANDN U28524 ( .A(y[1243]), .B(x[1243]), .Z(n12364) );
  AND U28525 ( .A(n12365), .B(n12364), .Z(n53292) );
  NANDN U28526 ( .A(n12366), .B(n53292), .Z(n12367) );
  NAND U28527 ( .A(n53293), .B(n12367), .Z(n12368) );
  NAND U28528 ( .A(n53294), .B(n12368), .Z(n12369) );
  NAND U28529 ( .A(n53295), .B(n12369), .Z(n12370) );
  NANDN U28530 ( .A(n53296), .B(n12370), .Z(n12371) );
  ANDN U28531 ( .B(y[1249]), .A(x[1249]), .Z(n53297) );
  ANDN U28532 ( .B(n12371), .A(n53297), .Z(n12372) );
  NANDN U28533 ( .A(x[1250]), .B(y[1250]), .Z(n27979) );
  NAND U28534 ( .A(n12372), .B(n27979), .Z(n12373) );
  NANDN U28535 ( .A(n12374), .B(n12373), .Z(n12375) );
  AND U28536 ( .A(n27978), .B(n12375), .Z(n12376) );
  NAND U28537 ( .A(n27977), .B(n12376), .Z(n12377) );
  NANDN U28538 ( .A(n52313), .B(n12377), .Z(n12378) );
  AND U28539 ( .A(n53303), .B(n12378), .Z(n12379) );
  ANDN U28540 ( .B(x[1255]), .A(y[1255]), .Z(n27975) );
  NANDN U28541 ( .A(y[1254]), .B(x[1254]), .Z(n32603) );
  NANDN U28542 ( .A(n27975), .B(n32603), .Z(n52312) );
  OR U28543 ( .A(n12379), .B(n52312), .Z(n12380) );
  NAND U28544 ( .A(n53304), .B(n12380), .Z(n12381) );
  NANDN U28545 ( .A(n53305), .B(n12381), .Z(n12382) );
  NAND U28546 ( .A(n53306), .B(n12382), .Z(n12383) );
  NANDN U28547 ( .A(n53307), .B(n12383), .Z(n12384) );
  AND U28548 ( .A(n53308), .B(n12384), .Z(n12385) );
  OR U28549 ( .A(n53309), .B(n12385), .Z(n12386) );
  NAND U28550 ( .A(n53310), .B(n12386), .Z(n12387) );
  NANDN U28551 ( .A(n53311), .B(n12387), .Z(n12388) );
  NAND U28552 ( .A(n53312), .B(n12388), .Z(n12389) );
  AND U28553 ( .A(n12390), .B(n12389), .Z(n12392) );
  ANDN U28554 ( .B(y[1266]), .A(x[1266]), .Z(n27966) );
  ANDN U28555 ( .B(y[1265]), .A(x[1265]), .Z(n53314) );
  NOR U28556 ( .A(n27966), .B(n53314), .Z(n12391) );
  NANDN U28557 ( .A(n12392), .B(n12391), .Z(n12393) );
  AND U28558 ( .A(n27969), .B(n12393), .Z(n12394) );
  NAND U28559 ( .A(n12395), .B(n12394), .Z(n12396) );
  NAND U28560 ( .A(n27967), .B(n12396), .Z(n12397) );
  AND U28561 ( .A(n27965), .B(n12397), .Z(n12398) );
  ANDN U28562 ( .B(y[1268]), .A(x[1268]), .Z(n27962) );
  OR U28563 ( .A(n12398), .B(n27962), .Z(n12399) );
  NAND U28564 ( .A(n53320), .B(n12399), .Z(n12400) );
  NANDN U28565 ( .A(n53321), .B(n12400), .Z(n12401) );
  NANDN U28566 ( .A(x[1269]), .B(y[1269]), .Z(n27963) );
  NANDN U28567 ( .A(n12401), .B(n27963), .Z(n12402) );
  NAND U28568 ( .A(n52311), .B(n12402), .Z(n12403) );
  NANDN U28569 ( .A(n53322), .B(n12403), .Z(n12404) );
  NAND U28570 ( .A(n53323), .B(n12404), .Z(n12405) );
  NAND U28571 ( .A(n53324), .B(n12405), .Z(n12406) );
  NANDN U28572 ( .A(n53325), .B(n12406), .Z(n12407) );
  ANDN U28573 ( .B(x[1275]), .A(y[1275]), .Z(n27960) );
  OR U28574 ( .A(n12407), .B(n27960), .Z(n12408) );
  AND U28575 ( .A(n27959), .B(n12408), .Z(n12409) );
  NANDN U28576 ( .A(x[1275]), .B(y[1275]), .Z(n53326) );
  NAND U28577 ( .A(n12409), .B(n53326), .Z(n12410) );
  NANDN U28578 ( .A(y[1276]), .B(x[1276]), .Z(n27961) );
  AND U28579 ( .A(n12410), .B(n27961), .Z(n12411) );
  NANDN U28580 ( .A(n53329), .B(n12411), .Z(n12412) );
  NANDN U28581 ( .A(x[1277]), .B(y[1277]), .Z(n27958) );
  AND U28582 ( .A(n12412), .B(n27958), .Z(n12413) );
  NAND U28583 ( .A(n53330), .B(n12413), .Z(n12414) );
  NANDN U28584 ( .A(n53331), .B(n12414), .Z(n12415) );
  NAND U28585 ( .A(n53332), .B(n12415), .Z(n12416) );
  NANDN U28586 ( .A(n53333), .B(n12416), .Z(n12417) );
  AND U28587 ( .A(n53334), .B(n12417), .Z(n12418) );
  OR U28588 ( .A(n53336), .B(n12418), .Z(n12419) );
  NAND U28589 ( .A(n53337), .B(n12419), .Z(n12420) );
  NANDN U28590 ( .A(n53338), .B(n12420), .Z(n12421) );
  NAND U28591 ( .A(n53339), .B(n12421), .Z(n12422) );
  NANDN U28592 ( .A(n53340), .B(n12422), .Z(n12423) );
  AND U28593 ( .A(n53341), .B(n12423), .Z(n12424) );
  OR U28594 ( .A(n53342), .B(n12424), .Z(n12425) );
  NAND U28595 ( .A(n53343), .B(n12425), .Z(n12426) );
  NANDN U28596 ( .A(n53344), .B(n12426), .Z(n12427) );
  NAND U28597 ( .A(n53345), .B(n12427), .Z(n12428) );
  NAND U28598 ( .A(n53346), .B(n12428), .Z(n12429) );
  NANDN U28599 ( .A(n52310), .B(n12429), .Z(n12430) );
  NANDN U28600 ( .A(y[1295]), .B(x[1295]), .Z(n27945) );
  AND U28601 ( .A(n12430), .B(n27945), .Z(n12431) );
  NANDN U28602 ( .A(n53347), .B(n12431), .Z(n12432) );
  NANDN U28603 ( .A(n12433), .B(n12432), .Z(n12435) );
  NANDN U28604 ( .A(y[1296]), .B(x[1296]), .Z(n27944) );
  ANDN U28605 ( .B(x[1297]), .A(y[1297]), .Z(n53350) );
  ANDN U28606 ( .B(n27944), .A(n53350), .Z(n12434) );
  NAND U28607 ( .A(n12435), .B(n12434), .Z(n12436) );
  NANDN U28608 ( .A(x[1297]), .B(y[1297]), .Z(n32725) );
  NANDN U28609 ( .A(x[1298]), .B(y[1298]), .Z(n32730) );
  AND U28610 ( .A(n32725), .B(n32730), .Z(n52307) );
  AND U28611 ( .A(n12436), .B(n52307), .Z(n12437) );
  ANDN U28612 ( .B(x[1298]), .A(y[1298]), .Z(n32727) );
  ANDN U28613 ( .B(x[1299]), .A(y[1299]), .Z(n32737) );
  OR U28614 ( .A(n32727), .B(n32737), .Z(n53351) );
  OR U28615 ( .A(n12437), .B(n53351), .Z(n12438) );
  NAND U28616 ( .A(n53352), .B(n12438), .Z(n12439) );
  NANDN U28617 ( .A(n52306), .B(n12439), .Z(n12440) );
  NANDN U28618 ( .A(n53353), .B(n12440), .Z(n12441) );
  AND U28619 ( .A(n53354), .B(n12441), .Z(n12443) );
  ANDN U28620 ( .B(y[1303]), .A(x[1303]), .Z(n32749) );
  IV U28621 ( .A(n32749), .Z(n53355) );
  ANDN U28622 ( .B(y[1304]), .A(x[1304]), .Z(n27942) );
  ANDN U28623 ( .B(n53355), .A(n27942), .Z(n12442) );
  NANDN U28624 ( .A(n12443), .B(n12442), .Z(n12444) );
  NAND U28625 ( .A(n32755), .B(n12444), .Z(n12445) );
  NANDN U28626 ( .A(y[1304]), .B(x[1304]), .Z(n53356) );
  NANDN U28627 ( .A(n12445), .B(n53356), .Z(n12446) );
  AND U28628 ( .A(n32757), .B(n12446), .Z(n12449) );
  NANDN U28629 ( .A(x[1305]), .B(y[1305]), .Z(n27943) );
  OR U28630 ( .A(n27943), .B(n12447), .Z(n12448) );
  NAND U28631 ( .A(n12449), .B(n12448), .Z(n12450) );
  NAND U28632 ( .A(n52304), .B(n12450), .Z(n12451) );
  NAND U28633 ( .A(n53360), .B(n12451), .Z(n12452) );
  NANDN U28634 ( .A(n53362), .B(n12452), .Z(n12455) );
  NANDN U28635 ( .A(x[1312]), .B(y[1312]), .Z(n12454) );
  NANDN U28636 ( .A(x[1311]), .B(y[1311]), .Z(n12453) );
  NAND U28637 ( .A(n12454), .B(n12453), .Z(n53364) );
  ANDN U28638 ( .B(n12455), .A(n53364), .Z(n12456) );
  OR U28639 ( .A(n53366), .B(n12456), .Z(n12457) );
  NAND U28640 ( .A(n53368), .B(n12457), .Z(n12458) );
  NANDN U28641 ( .A(n53370), .B(n12458), .Z(n12459) );
  NAND U28642 ( .A(n53372), .B(n12459), .Z(n12460) );
  NANDN U28643 ( .A(n53374), .B(n12460), .Z(n12461) );
  AND U28644 ( .A(n53376), .B(n12461), .Z(n12462) );
  OR U28645 ( .A(n53378), .B(n12462), .Z(n12463) );
  NAND U28646 ( .A(n53380), .B(n12463), .Z(n12464) );
  NANDN U28647 ( .A(n53382), .B(n12464), .Z(n12465) );
  NAND U28648 ( .A(n53384), .B(n12465), .Z(n12466) );
  NANDN U28649 ( .A(n53386), .B(n12466), .Z(n12467) );
  AND U28650 ( .A(n53388), .B(n12467), .Z(n12468) );
  OR U28651 ( .A(n53390), .B(n12468), .Z(n12469) );
  NAND U28652 ( .A(n53392), .B(n12469), .Z(n12470) );
  NANDN U28653 ( .A(n53394), .B(n12470), .Z(n12471) );
  NAND U28654 ( .A(n53396), .B(n12471), .Z(n12472) );
  NANDN U28655 ( .A(n53398), .B(n12472), .Z(n12473) );
  AND U28656 ( .A(n53400), .B(n12473), .Z(n12474) );
  OR U28657 ( .A(n53402), .B(n12474), .Z(n12475) );
  NAND U28658 ( .A(n53404), .B(n12475), .Z(n12476) );
  NANDN U28659 ( .A(n53405), .B(n12476), .Z(n12477) );
  NAND U28660 ( .A(n53406), .B(n12477), .Z(n12478) );
  NAND U28661 ( .A(n53407), .B(n12478), .Z(n12479) );
  NANDN U28662 ( .A(n52303), .B(n12479), .Z(n12480) );
  NANDN U28663 ( .A(y[1337]), .B(x[1337]), .Z(n32847) );
  AND U28664 ( .A(n12480), .B(n32847), .Z(n12481) );
  NANDN U28665 ( .A(n53408), .B(n12481), .Z(n12482) );
  NANDN U28666 ( .A(n53409), .B(n12482), .Z(n12484) );
  NANDN U28667 ( .A(y[1338]), .B(x[1338]), .Z(n32846) );
  ANDN U28668 ( .B(x[1339]), .A(y[1339]), .Z(n53410) );
  ANDN U28669 ( .B(n32846), .A(n53410), .Z(n12483) );
  NAND U28670 ( .A(n12484), .B(n12483), .Z(n12485) );
  AND U28671 ( .A(n53413), .B(n12485), .Z(n12486) );
  ANDN U28672 ( .B(x[1340]), .A(y[1340]), .Z(n32852) );
  NANDN U28673 ( .A(y[1341]), .B(x[1341]), .Z(n32856) );
  NANDN U28674 ( .A(n32852), .B(n32856), .Z(n52302) );
  OR U28675 ( .A(n12486), .B(n52302), .Z(n12487) );
  NAND U28676 ( .A(n53414), .B(n12487), .Z(n12488) );
  NANDN U28677 ( .A(n53415), .B(n12488), .Z(n12489) );
  NAND U28678 ( .A(n53416), .B(n12489), .Z(n12490) );
  NANDN U28679 ( .A(n53417), .B(n12490), .Z(n12491) );
  AND U28680 ( .A(n53419), .B(n12491), .Z(n12492) );
  OR U28681 ( .A(n53420), .B(n12492), .Z(n12493) );
  NAND U28682 ( .A(n53421), .B(n12493), .Z(n12494) );
  NANDN U28683 ( .A(n53422), .B(n12494), .Z(n12495) );
  ANDN U28684 ( .B(y[1349]), .A(x[1349]), .Z(n53423) );
  ANDN U28685 ( .B(n12495), .A(n53423), .Z(n12496) );
  ANDN U28686 ( .B(x[1350]), .A(y[1350]), .Z(n27913) );
  OR U28687 ( .A(n12496), .B(n27913), .Z(n12497) );
  NANDN U28688 ( .A(n32888), .B(n12497), .Z(n12498) );
  NAND U28689 ( .A(n52300), .B(n12498), .Z(n12499) );
  NANDN U28690 ( .A(n53425), .B(n12499), .Z(n12500) );
  NANDN U28691 ( .A(n53427), .B(n12500), .Z(n12501) );
  AND U28692 ( .A(n53428), .B(n12501), .Z(n12502) );
  NANDN U28693 ( .A(y[1354]), .B(x[1354]), .Z(n27911) );
  NANDN U28694 ( .A(y[1355]), .B(x[1355]), .Z(n27909) );
  NAND U28695 ( .A(n27911), .B(n27909), .Z(n52299) );
  OR U28696 ( .A(n12502), .B(n52299), .Z(n12503) );
  NAND U28697 ( .A(n53429), .B(n12503), .Z(n12504) );
  NANDN U28698 ( .A(n52298), .B(n12504), .Z(n12505) );
  NAND U28699 ( .A(n52297), .B(n12505), .Z(n12506) );
  NANDN U28700 ( .A(n53430), .B(n12506), .Z(n12507) );
  NANDN U28701 ( .A(x[1359]), .B(y[1359]), .Z(n32909) );
  NANDN U28702 ( .A(x[1360]), .B(y[1360]), .Z(n32916) );
  AND U28703 ( .A(n32909), .B(n32916), .Z(n53433) );
  AND U28704 ( .A(n12507), .B(n53433), .Z(n12508) );
  NANDN U28705 ( .A(y[1360]), .B(x[1360]), .Z(n27905) );
  NANDN U28706 ( .A(y[1361]), .B(x[1361]), .Z(n27904) );
  NAND U28707 ( .A(n27905), .B(n27904), .Z(n52296) );
  OR U28708 ( .A(n12508), .B(n52296), .Z(n12509) );
  NAND U28709 ( .A(n52295), .B(n12509), .Z(n12510) );
  NANDN U28710 ( .A(n52294), .B(n12510), .Z(n12511) );
  NAND U28711 ( .A(n52293), .B(n12511), .Z(n12512) );
  ANDN U28712 ( .B(x[1366]), .A(y[1366]), .Z(n32932) );
  NANDN U28713 ( .A(y[1367]), .B(x[1367]), .Z(n27899) );
  NANDN U28714 ( .A(n32932), .B(n27899), .Z(n52292) );
  NANDN U28715 ( .A(x[1371]), .B(y[1371]), .Z(n32946) );
  XNOR U28716 ( .A(y[1372]), .B(x[1372]), .Z(n12513) );
  AND U28717 ( .A(n32946), .B(n12513), .Z(n53440) );
  ANDN U28718 ( .B(x[1372]), .A(y[1372]), .Z(n32950) );
  ANDN U28719 ( .B(x[1373]), .A(y[1373]), .Z(n32958) );
  OR U28720 ( .A(n32950), .B(n32958), .Z(n52288) );
  NANDN U28721 ( .A(y[1379]), .B(x[1379]), .Z(n27890) );
  NANDN U28722 ( .A(y[1383]), .B(x[1383]), .Z(n12515) );
  NANDN U28723 ( .A(y[1382]), .B(x[1382]), .Z(n12514) );
  AND U28724 ( .A(n12515), .B(n12514), .Z(n53448) );
  AND U28725 ( .A(n12516), .B(n53448), .Z(n12519) );
  NANDN U28726 ( .A(x[1384]), .B(y[1384]), .Z(n12518) );
  NANDN U28727 ( .A(x[1383]), .B(y[1383]), .Z(n12517) );
  NAND U28728 ( .A(n12518), .B(n12517), .Z(n53449) );
  OR U28729 ( .A(n12519), .B(n53449), .Z(n12520) );
  NANDN U28730 ( .A(y[1384]), .B(x[1384]), .Z(n53452) );
  AND U28731 ( .A(n12520), .B(n53452), .Z(n12521) );
  NANDN U28732 ( .A(y[1385]), .B(x[1385]), .Z(n27887) );
  NAND U28733 ( .A(n12521), .B(n27887), .Z(n12522) );
  ANDN U28734 ( .B(y[1386]), .A(x[1386]), .Z(n27883) );
  ANDN U28735 ( .B(n12522), .A(n27883), .Z(n12523) );
  NANDN U28736 ( .A(n52285), .B(n12523), .Z(n12524) );
  NANDN U28737 ( .A(y[1386]), .B(x[1386]), .Z(n27886) );
  AND U28738 ( .A(n12524), .B(n27886), .Z(n12525) );
  NAND U28739 ( .A(n27882), .B(n12525), .Z(n12526) );
  NANDN U28740 ( .A(n27884), .B(n12526), .Z(n12527) );
  ANDN U28741 ( .B(y[1388]), .A(x[1388]), .Z(n27879) );
  OR U28742 ( .A(n12527), .B(n27879), .Z(n12528) );
  NANDN U28743 ( .A(y[1389]), .B(x[1389]), .Z(n53456) );
  AND U28744 ( .A(n12528), .B(n53456), .Z(n12529) );
  NANDN U28745 ( .A(n27881), .B(n12529), .Z(n12530) );
  AND U28746 ( .A(n27880), .B(n12530), .Z(n12531) );
  NANDN U28747 ( .A(x[1390]), .B(y[1390]), .Z(n53457) );
  NAND U28748 ( .A(n12531), .B(n53457), .Z(n12532) );
  NANDN U28749 ( .A(n53458), .B(n12532), .Z(n12533) );
  AND U28750 ( .A(n53459), .B(n12533), .Z(n12534) );
  OR U28751 ( .A(n53460), .B(n12534), .Z(n12535) );
  NAND U28752 ( .A(n53461), .B(n12535), .Z(n12536) );
  NANDN U28753 ( .A(n53462), .B(n12536), .Z(n12537) );
  NANDN U28754 ( .A(n52283), .B(n12537), .Z(n12538) );
  AND U28755 ( .A(n53464), .B(n12538), .Z(n12540) );
  NANDN U28756 ( .A(x[1398]), .B(y[1398]), .Z(n27870) );
  ANDN U28757 ( .B(y[1397]), .A(x[1397]), .Z(n33007) );
  ANDN U28758 ( .B(n27870), .A(n33007), .Z(n12539) );
  NANDN U28759 ( .A(n12540), .B(n12539), .Z(n12541) );
  NANDN U28760 ( .A(y[1398]), .B(x[1398]), .Z(n33013) );
  AND U28761 ( .A(n12541), .B(n33013), .Z(n12542) );
  NANDN U28762 ( .A(y[1399]), .B(x[1399]), .Z(n27869) );
  NAND U28763 ( .A(n12542), .B(n27869), .Z(n12543) );
  NAND U28764 ( .A(n27871), .B(n12543), .Z(n12544) );
  ANDN U28765 ( .B(y[1400]), .A(x[1400]), .Z(n27866) );
  OR U28766 ( .A(n12544), .B(n27866), .Z(n12545) );
  NAND U28767 ( .A(n12546), .B(n12545), .Z(n12547) );
  NANDN U28768 ( .A(n12548), .B(n12547), .Z(n12549) );
  NAND U28769 ( .A(n53472), .B(n12549), .Z(n12550) );
  NANDN U28770 ( .A(n53473), .B(n12550), .Z(n12551) );
  NANDN U28771 ( .A(y[1404]), .B(x[1404]), .Z(n27864) );
  NANDN U28772 ( .A(y[1405]), .B(x[1405]), .Z(n33032) );
  AND U28773 ( .A(n27864), .B(n33032), .Z(n53474) );
  AND U28774 ( .A(n12551), .B(n53474), .Z(n12552) );
  NANDN U28775 ( .A(x[1405]), .B(y[1405]), .Z(n33027) );
  NANDN U28776 ( .A(x[1406]), .B(y[1406]), .Z(n27863) );
  NAND U28777 ( .A(n33027), .B(n27863), .Z(n52282) );
  OR U28778 ( .A(n12552), .B(n52282), .Z(n12553) );
  NAND U28779 ( .A(n53475), .B(n12553), .Z(n12554) );
  NANDN U28780 ( .A(n27862), .B(n12554), .Z(n12555) );
  NAND U28781 ( .A(n53477), .B(n12555), .Z(n12556) );
  NAND U28782 ( .A(n53478), .B(n12556), .Z(n12557) );
  NANDN U28783 ( .A(n53479), .B(n12557), .Z(n12558) );
  NANDN U28784 ( .A(n53480), .B(n12558), .Z(n12559) );
  NANDN U28785 ( .A(y[1412]), .B(x[1412]), .Z(n27856) );
  NANDN U28786 ( .A(y[1413]), .B(x[1413]), .Z(n33055) );
  AND U28787 ( .A(n27856), .B(n33055), .Z(n53483) );
  AND U28788 ( .A(n12559), .B(n53483), .Z(n12560) );
  ANDN U28789 ( .B(y[1413]), .A(x[1413]), .Z(n33051) );
  NANDN U28790 ( .A(x[1414]), .B(y[1414]), .Z(n27854) );
  NANDN U28791 ( .A(n33051), .B(n27854), .Z(n52281) );
  OR U28792 ( .A(n12560), .B(n52281), .Z(n12561) );
  AND U28793 ( .A(n12562), .B(n12561), .Z(n12564) );
  NANDN U28794 ( .A(x[1415]), .B(y[1415]), .Z(n53486) );
  NANDN U28795 ( .A(x[1416]), .B(y[1416]), .Z(n53488) );
  NAND U28796 ( .A(n53486), .B(n53488), .Z(n12563) );
  OR U28797 ( .A(n12564), .B(n12563), .Z(n12565) );
  AND U28798 ( .A(n27852), .B(n12565), .Z(n12566) );
  NAND U28799 ( .A(n33064), .B(n12566), .Z(n12567) );
  NANDN U28800 ( .A(n53490), .B(n12567), .Z(n12568) );
  AND U28801 ( .A(n53491), .B(n12568), .Z(n12569) );
  ANDN U28802 ( .B(y[1419]), .A(x[1419]), .Z(n27850) );
  ANDN U28803 ( .B(y[1420]), .A(x[1420]), .Z(n33072) );
  OR U28804 ( .A(n27850), .B(n33072), .Z(n53492) );
  OR U28805 ( .A(n12569), .B(n53492), .Z(n12570) );
  NANDN U28806 ( .A(y[1420]), .B(x[1420]), .Z(n53493) );
  AND U28807 ( .A(n12570), .B(n53493), .Z(n12571) );
  NANDN U28808 ( .A(y[1421]), .B(x[1421]), .Z(n27848) );
  NAND U28809 ( .A(n12571), .B(n27848), .Z(n12572) );
  ANDN U28810 ( .B(y[1421]), .A(x[1421]), .Z(n52280) );
  ANDN U28811 ( .B(n12572), .A(n52280), .Z(n12573) );
  NANDN U28812 ( .A(n27846), .B(n12573), .Z(n12575) );
  NANDN U28813 ( .A(y[1422]), .B(x[1422]), .Z(n12574) );
  AND U28814 ( .A(n12575), .B(n12574), .Z(n12576) );
  NAND U28815 ( .A(n27845), .B(n12576), .Z(n12577) );
  NANDN U28816 ( .A(n33075), .B(n12577), .Z(n12578) );
  ANDN U28817 ( .B(y[1424]), .A(x[1424]), .Z(n27842) );
  OR U28818 ( .A(n12578), .B(n27842), .Z(n12579) );
  NAND U28819 ( .A(n12580), .B(n12579), .Z(n12581) );
  NANDN U28820 ( .A(n27843), .B(n12581), .Z(n12582) );
  ANDN U28821 ( .B(y[1426]), .A(x[1426]), .Z(n52278) );
  OR U28822 ( .A(n12582), .B(n52278), .Z(n12583) );
  NAND U28823 ( .A(n53499), .B(n12583), .Z(n12584) );
  NANDN U28824 ( .A(n53500), .B(n12584), .Z(n12585) );
  NAND U28825 ( .A(n53501), .B(n12585), .Z(n12586) );
  ANDN U28826 ( .B(y[1430]), .A(x[1430]), .Z(n27839) );
  ANDN U28827 ( .B(n12586), .A(n27839), .Z(n12587) );
  NAND U28828 ( .A(n53502), .B(n12587), .Z(n12588) );
  ANDN U28829 ( .B(x[1430]), .A(y[1430]), .Z(n53503) );
  ANDN U28830 ( .B(n12588), .A(n53503), .Z(n12589) );
  NAND U28831 ( .A(n27838), .B(n12589), .Z(n12590) );
  NAND U28832 ( .A(n27841), .B(n12590), .Z(n12591) );
  ANDN U28833 ( .B(y[1432]), .A(x[1432]), .Z(n27834) );
  OR U28834 ( .A(n12591), .B(n27834), .Z(n12592) );
  NAND U28835 ( .A(n12593), .B(n12592), .Z(n12594) );
  NANDN U28836 ( .A(x[1434]), .B(y[1434]), .Z(n53508) );
  AND U28837 ( .A(n12594), .B(n53508), .Z(n12595) );
  NAND U28838 ( .A(n27836), .B(n12595), .Z(n12596) );
  NANDN U28839 ( .A(n52277), .B(n12596), .Z(n12597) );
  ANDN U28840 ( .B(x[1434]), .A(y[1434]), .Z(n33097) );
  OR U28841 ( .A(n12597), .B(n33097), .Z(n12598) );
  NANDN U28842 ( .A(x[1435]), .B(y[1435]), .Z(n33101) );
  NANDN U28843 ( .A(x[1436]), .B(y[1436]), .Z(n33106) );
  AND U28844 ( .A(n33101), .B(n33106), .Z(n52276) );
  AND U28845 ( .A(n12598), .B(n52276), .Z(n12599) );
  OR U28846 ( .A(n53510), .B(n12599), .Z(n12600) );
  NAND U28847 ( .A(n53511), .B(n12600), .Z(n12601) );
  NANDN U28848 ( .A(n53512), .B(n12601), .Z(n12602) );
  NANDN U28849 ( .A(y[1439]), .B(x[1439]), .Z(n27833) );
  NANDN U28850 ( .A(n12602), .B(n27833), .Z(n12603) );
  AND U28851 ( .A(n33118), .B(n12603), .Z(n12604) );
  NANDN U28852 ( .A(n53513), .B(n12604), .Z(n12605) );
  ANDN U28853 ( .B(x[1440]), .A(y[1440]), .Z(n27832) );
  ANDN U28854 ( .B(n12605), .A(n27832), .Z(n12606) );
  NANDN U28855 ( .A(n27830), .B(n12606), .Z(n12609) );
  NANDN U28856 ( .A(x[1442]), .B(y[1442]), .Z(n12607) );
  NAND U28857 ( .A(n12608), .B(n12607), .Z(n53516) );
  ANDN U28858 ( .B(n12609), .A(n53516), .Z(n12610) );
  NAND U28859 ( .A(n33117), .B(n12610), .Z(n12611) );
  NANDN U28860 ( .A(n52274), .B(n12611), .Z(n12612) );
  NAND U28861 ( .A(n33125), .B(n12612), .Z(n12613) );
  NANDN U28862 ( .A(n53518), .B(n12613), .Z(n12614) );
  AND U28863 ( .A(n53519), .B(n12614), .Z(n12615) );
  NANDN U28864 ( .A(y[1448]), .B(x[1448]), .Z(n33132) );
  NANDN U28865 ( .A(y[1449]), .B(x[1449]), .Z(n33141) );
  NAND U28866 ( .A(n33132), .B(n33141), .Z(n52273) );
  OR U28867 ( .A(n12615), .B(n52273), .Z(n12616) );
  NAND U28868 ( .A(n53520), .B(n12616), .Z(n12617) );
  NANDN U28869 ( .A(n52272), .B(n12617), .Z(n12618) );
  NAND U28870 ( .A(n53522), .B(n12618), .Z(n12619) );
  NANDN U28871 ( .A(n53523), .B(n12619), .Z(n12620) );
  NANDN U28872 ( .A(x[1453]), .B(y[1453]), .Z(n27822) );
  NANDN U28873 ( .A(x[1454]), .B(y[1454]), .Z(n27819) );
  AND U28874 ( .A(n27822), .B(n27819), .Z(n53524) );
  AND U28875 ( .A(n12620), .B(n53524), .Z(n12621) );
  NANDN U28876 ( .A(y[1454]), .B(x[1454]), .Z(n27820) );
  NANDN U28877 ( .A(y[1455]), .B(x[1455]), .Z(n33155) );
  NAND U28878 ( .A(n27820), .B(n33155), .Z(n52271) );
  OR U28879 ( .A(n12621), .B(n52271), .Z(n12622) );
  NAND U28880 ( .A(n52270), .B(n12622), .Z(n12623) );
  NANDN U28881 ( .A(n52269), .B(n12623), .Z(n12624) );
  NAND U28882 ( .A(n53525), .B(n12624), .Z(n12625) );
  NANDN U28883 ( .A(n53526), .B(n12625), .Z(n12626) );
  AND U28884 ( .A(n53527), .B(n12626), .Z(n12627) );
  NANDN U28885 ( .A(y[1460]), .B(x[1460]), .Z(n33170) );
  NANDN U28886 ( .A(y[1461]), .B(x[1461]), .Z(n33178) );
  NAND U28887 ( .A(n33170), .B(n33178), .Z(n52268) );
  OR U28888 ( .A(n12627), .B(n52268), .Z(n12628) );
  NAND U28889 ( .A(n53528), .B(n12628), .Z(n12629) );
  NANDN U28890 ( .A(n33177), .B(n12629), .Z(n12630) );
  NANDN U28891 ( .A(y[1463]), .B(x[1463]), .Z(n27814) );
  NANDN U28892 ( .A(n12630), .B(n27814), .Z(n12631) );
  AND U28893 ( .A(n12632), .B(n12631), .Z(n12634) );
  NANDN U28894 ( .A(y[1465]), .B(x[1465]), .Z(n53534) );
  ANDN U28895 ( .B(x[1464]), .A(y[1464]), .Z(n27813) );
  ANDN U28896 ( .B(n53534), .A(n27813), .Z(n12633) );
  NANDN U28897 ( .A(n12634), .B(n12633), .Z(n12635) );
  NANDN U28898 ( .A(n52267), .B(n12635), .Z(n12636) );
  NANDN U28899 ( .A(n53535), .B(n12636), .Z(n12637) );
  AND U28900 ( .A(n53536), .B(n12637), .Z(n12638) );
  NANDN U28901 ( .A(y[1468]), .B(x[1468]), .Z(n27811) );
  NANDN U28902 ( .A(n12638), .B(n27811), .Z(n12639) );
  ANDN U28903 ( .B(x[1469]), .A(y[1469]), .Z(n27805) );
  OR U28904 ( .A(n12639), .B(n27805), .Z(n12640) );
  NAND U28905 ( .A(n53538), .B(n12640), .Z(n12641) );
  NANDN U28906 ( .A(n27809), .B(n12641), .Z(n12644) );
  ANDN U28907 ( .B(x[1470]), .A(y[1470]), .Z(n27804) );
  NAND U28908 ( .A(n27804), .B(n12642), .Z(n12643) );
  NANDN U28909 ( .A(n12644), .B(n12643), .Z(n12645) );
  AND U28910 ( .A(n53540), .B(n12645), .Z(n12646) );
  OR U28911 ( .A(n53541), .B(n12646), .Z(n12647) );
  NAND U28912 ( .A(n53542), .B(n12647), .Z(n12648) );
  NANDN U28913 ( .A(n53543), .B(n12648), .Z(n12649) );
  NAND U28914 ( .A(n53544), .B(n12649), .Z(n12650) );
  NANDN U28915 ( .A(n53545), .B(n12650), .Z(n12651) );
  AND U28916 ( .A(n53546), .B(n12651), .Z(n12652) );
  OR U28917 ( .A(n53547), .B(n12652), .Z(n12653) );
  NAND U28918 ( .A(n53549), .B(n12653), .Z(n12654) );
  NAND U28919 ( .A(n53550), .B(n12654), .Z(n12656) );
  NANDN U28920 ( .A(x[1482]), .B(y[1482]), .Z(n33231) );
  ANDN U28921 ( .B(y[1481]), .A(x[1481]), .Z(n53551) );
  ANDN U28922 ( .B(n33231), .A(n53551), .Z(n12655) );
  NAND U28923 ( .A(n12656), .B(n12655), .Z(n12657) );
  AND U28924 ( .A(n12658), .B(n12657), .Z(n12660) );
  NANDN U28925 ( .A(x[1483]), .B(y[1483]), .Z(n33230) );
  ANDN U28926 ( .B(y[1484]), .A(x[1484]), .Z(n52265) );
  ANDN U28927 ( .B(n33230), .A(n52265), .Z(n12659) );
  NANDN U28928 ( .A(n12660), .B(n12659), .Z(n12661) );
  AND U28929 ( .A(n53554), .B(n12661), .Z(n12662) );
  ANDN U28930 ( .B(y[1485]), .A(x[1485]), .Z(n33236) );
  NANDN U28931 ( .A(x[1486]), .B(y[1486]), .Z(n33240) );
  NANDN U28932 ( .A(n33236), .B(n33240), .Z(n53555) );
  OR U28933 ( .A(n12662), .B(n53555), .Z(n12663) );
  NAND U28934 ( .A(n53556), .B(n12663), .Z(n12664) );
  NANDN U28935 ( .A(n52264), .B(n12664), .Z(n12665) );
  NAND U28936 ( .A(n53557), .B(n12665), .Z(n12666) );
  NAND U28937 ( .A(n53558), .B(n12666), .Z(n12667) );
  NANDN U28938 ( .A(n53559), .B(n12667), .Z(n12668) );
  NAND U28939 ( .A(n53560), .B(n12668), .Z(n12669) );
  NANDN U28940 ( .A(n53562), .B(n12669), .Z(n12670) );
  AND U28941 ( .A(n53563), .B(n12670), .Z(n12671) );
  OR U28942 ( .A(n53564), .B(n12671), .Z(n12672) );
  NAND U28943 ( .A(n53565), .B(n12672), .Z(n12673) );
  NANDN U28944 ( .A(n52263), .B(n12673), .Z(n12674) );
  NANDN U28945 ( .A(n53566), .B(n12674), .Z(n12675) );
  AND U28946 ( .A(n27788), .B(n12675), .Z(n12676) );
  NANDN U28947 ( .A(n52262), .B(n12676), .Z(n12677) );
  NAND U28948 ( .A(n12678), .B(n12677), .Z(n12679) );
  NAND U28949 ( .A(n53570), .B(n12679), .Z(n12680) );
  ANDN U28950 ( .B(x[1500]), .A(y[1500]), .Z(n27787) );
  OR U28951 ( .A(n12680), .B(n27787), .Z(n12681) );
  NAND U28952 ( .A(n53571), .B(n12681), .Z(n12682) );
  NANDN U28953 ( .A(n53572), .B(n12682), .Z(n12683) );
  NAND U28954 ( .A(n53573), .B(n12683), .Z(n12684) );
  AND U28955 ( .A(n12685), .B(n12684), .Z(n12687) );
  NANDN U28956 ( .A(x[1505]), .B(y[1505]), .Z(n53575) );
  ANDN U28957 ( .B(y[1506]), .A(x[1506]), .Z(n27780) );
  ANDN U28958 ( .B(n53575), .A(n27780), .Z(n12686) );
  NANDN U28959 ( .A(n12687), .B(n12686), .Z(n12688) );
  NANDN U28960 ( .A(y[1507]), .B(x[1507]), .Z(n33300) );
  AND U28961 ( .A(n12688), .B(n33300), .Z(n12689) );
  NANDN U28962 ( .A(y[1506]), .B(x[1506]), .Z(n27783) );
  NAND U28963 ( .A(n12689), .B(n27783), .Z(n12690) );
  NANDN U28964 ( .A(n53580), .B(n12690), .Z(n12691) );
  AND U28965 ( .A(n53581), .B(n12691), .Z(n12692) );
  NANDN U28966 ( .A(x[1509]), .B(y[1509]), .Z(n27779) );
  NANDN U28967 ( .A(x[1510]), .B(y[1510]), .Z(n27774) );
  NAND U28968 ( .A(n27779), .B(n27774), .Z(n52261) );
  OR U28969 ( .A(n12692), .B(n52261), .Z(n12693) );
  NAND U28970 ( .A(n52260), .B(n12693), .Z(n12694) );
  NANDN U28971 ( .A(n53582), .B(n12694), .Z(n12695) );
  NAND U28972 ( .A(n53583), .B(n12695), .Z(n12696) );
  NANDN U28973 ( .A(x[1514]), .B(y[1514]), .Z(n27773) );
  AND U28974 ( .A(n12696), .B(n27773), .Z(n12697) );
  NANDN U28975 ( .A(n53584), .B(n12697), .Z(n12698) );
  ANDN U28976 ( .B(x[1514]), .A(y[1514]), .Z(n53585) );
  ANDN U28977 ( .B(n12698), .A(n53585), .Z(n12699) );
  NAND U28978 ( .A(n33319), .B(n12699), .Z(n12700) );
  NANDN U28979 ( .A(n27772), .B(n12700), .Z(n12701) );
  NANDN U28980 ( .A(x[1516]), .B(y[1516]), .Z(n27771) );
  NANDN U28981 ( .A(n12701), .B(n27771), .Z(n12702) );
  NAND U28982 ( .A(n12703), .B(n12702), .Z(n12704) );
  NANDN U28983 ( .A(n27770), .B(n12704), .Z(n12705) );
  NANDN U28984 ( .A(x[1518]), .B(y[1518]), .Z(n53589) );
  NANDN U28985 ( .A(n12705), .B(n53589), .Z(n12706) );
  AND U28986 ( .A(n12707), .B(n12706), .Z(n12708) );
  OR U28987 ( .A(n53592), .B(n12708), .Z(n12709) );
  NAND U28988 ( .A(n53593), .B(n12709), .Z(n12710) );
  NANDN U28989 ( .A(n53594), .B(n12710), .Z(n12711) );
  NANDN U28990 ( .A(y[1522]), .B(x[1522]), .Z(n53595) );
  AND U28991 ( .A(n12711), .B(n53595), .Z(n12712) );
  NAND U28992 ( .A(n33338), .B(n12712), .Z(n12713) );
  NANDN U28993 ( .A(n52258), .B(n12713), .Z(n12714) );
  ANDN U28994 ( .B(y[1524]), .A(x[1524]), .Z(n27764) );
  OR U28995 ( .A(n12714), .B(n27764), .Z(n12715) );
  AND U28996 ( .A(n12716), .B(n12715), .Z(n12718) );
  NANDN U28997 ( .A(x[1525]), .B(y[1525]), .Z(n27765) );
  ANDN U28998 ( .B(y[1526]), .A(x[1526]), .Z(n53598) );
  ANDN U28999 ( .B(n27765), .A(n53598), .Z(n12717) );
  NANDN U29000 ( .A(n12718), .B(n12717), .Z(n12719) );
  ANDN U29001 ( .B(x[1527]), .A(y[1527]), .Z(n53599) );
  ANDN U29002 ( .B(n12719), .A(n53599), .Z(n12720) );
  NANDN U29003 ( .A(y[1526]), .B(x[1526]), .Z(n27763) );
  NAND U29004 ( .A(n12720), .B(n27763), .Z(n12721) );
  NANDN U29005 ( .A(n53600), .B(n12721), .Z(n12722) );
  AND U29006 ( .A(n53601), .B(n12722), .Z(n12723) );
  OR U29007 ( .A(n53602), .B(n12723), .Z(n12724) );
  NAND U29008 ( .A(n53603), .B(n12724), .Z(n12725) );
  NANDN U29009 ( .A(n53604), .B(n12725), .Z(n12726) );
  NAND U29010 ( .A(n53605), .B(n12726), .Z(n12727) );
  NAND U29011 ( .A(n53607), .B(n12727), .Z(n12730) );
  NANDN U29012 ( .A(y[1535]), .B(x[1535]), .Z(n12729) );
  NANDN U29013 ( .A(y[1534]), .B(x[1534]), .Z(n12728) );
  NAND U29014 ( .A(n12729), .B(n12728), .Z(n53608) );
  ANDN U29015 ( .B(n12730), .A(n53608), .Z(n12731) );
  OR U29016 ( .A(n53609), .B(n12731), .Z(n12732) );
  NAND U29017 ( .A(n53610), .B(n12732), .Z(n12733) );
  NANDN U29018 ( .A(n53611), .B(n12733), .Z(n12734) );
  NAND U29019 ( .A(n53612), .B(n12734), .Z(n12735) );
  NANDN U29020 ( .A(n53613), .B(n12735), .Z(n12736) );
  AND U29021 ( .A(n53614), .B(n12736), .Z(n12737) );
  OR U29022 ( .A(n53615), .B(n12737), .Z(n12738) );
  NAND U29023 ( .A(n53616), .B(n12738), .Z(n12739) );
  NANDN U29024 ( .A(n53617), .B(n12739), .Z(n12740) );
  NANDN U29025 ( .A(n52256), .B(n12740), .Z(n12741) );
  AND U29026 ( .A(n53618), .B(n12741), .Z(n12743) );
  NANDN U29027 ( .A(y[1547]), .B(x[1547]), .Z(n53622) );
  ANDN U29028 ( .B(x[1546]), .A(y[1546]), .Z(n52255) );
  ANDN U29029 ( .B(n53622), .A(n52255), .Z(n12742) );
  NANDN U29030 ( .A(n12743), .B(n12742), .Z(n12744) );
  NANDN U29031 ( .A(n53619), .B(n12744), .Z(n12745) );
  NAND U29032 ( .A(n53620), .B(n12745), .Z(n12746) );
  NANDN U29033 ( .A(n53624), .B(n12746), .Z(n12747) );
  NANDN U29034 ( .A(y[1550]), .B(x[1550]), .Z(n27742) );
  NANDN U29035 ( .A(y[1551]), .B(x[1551]), .Z(n33410) );
  AND U29036 ( .A(n27742), .B(n33410), .Z(n52254) );
  AND U29037 ( .A(n12747), .B(n52254), .Z(n12748) );
  ANDN U29038 ( .B(y[1552]), .A(x[1552]), .Z(n33414) );
  NANDN U29039 ( .A(x[1551]), .B(y[1551]), .Z(n27740) );
  NANDN U29040 ( .A(n33414), .B(n27740), .Z(n53625) );
  OR U29041 ( .A(n12748), .B(n53625), .Z(n12749) );
  NANDN U29042 ( .A(y[1552]), .B(x[1552]), .Z(n53626) );
  AND U29043 ( .A(n12749), .B(n53626), .Z(n12750) );
  NANDN U29044 ( .A(y[1553]), .B(x[1553]), .Z(n33417) );
  NAND U29045 ( .A(n12750), .B(n33417), .Z(n12751) );
  ANDN U29046 ( .B(y[1554]), .A(x[1554]), .Z(n33419) );
  ANDN U29047 ( .B(n12751), .A(n33419), .Z(n12752) );
  NANDN U29048 ( .A(n52253), .B(n12752), .Z(n12753) );
  NANDN U29049 ( .A(y[1554]), .B(x[1554]), .Z(n33416) );
  AND U29050 ( .A(n12753), .B(n33416), .Z(n12754) );
  NAND U29051 ( .A(n27739), .B(n12754), .Z(n12755) );
  NANDN U29052 ( .A(n33420), .B(n12755), .Z(n12756) );
  ANDN U29053 ( .B(y[1556]), .A(x[1556]), .Z(n27736) );
  OR U29054 ( .A(n12756), .B(n27736), .Z(n12757) );
  ANDN U29055 ( .B(x[1558]), .A(y[1558]), .Z(n12760) );
  IV U29056 ( .A(n12760), .Z(n52251) );
  ANDN U29057 ( .B(x[1557]), .A(y[1557]), .Z(n53630) );
  ANDN U29058 ( .B(n52251), .A(n53630), .Z(n33425) );
  AND U29059 ( .A(n12757), .B(n33425), .Z(n12758) );
  NANDN U29060 ( .A(n27738), .B(n12758), .Z(n12759) );
  AND U29061 ( .A(n33427), .B(n12759), .Z(n12762) );
  NANDN U29062 ( .A(x[1557]), .B(y[1557]), .Z(n27737) );
  OR U29063 ( .A(n27737), .B(n12760), .Z(n12761) );
  NAND U29064 ( .A(n12762), .B(n12761), .Z(n12763) );
  NAND U29065 ( .A(n52250), .B(n12763), .Z(n12764) );
  NANDN U29066 ( .A(n53633), .B(n12764), .Z(n12765) );
  NANDN U29067 ( .A(n53635), .B(n12765), .Z(n12766) );
  AND U29068 ( .A(n53637), .B(n12766), .Z(n12767) );
  OR U29069 ( .A(n53639), .B(n12767), .Z(n12768) );
  NAND U29070 ( .A(n53641), .B(n12768), .Z(n12769) );
  NANDN U29071 ( .A(n53642), .B(n12769), .Z(n12770) );
  NANDN U29072 ( .A(x[1565]), .B(y[1565]), .Z(n53645) );
  AND U29073 ( .A(n12770), .B(n53645), .Z(n12771) );
  NAND U29074 ( .A(n27731), .B(n12771), .Z(n12772) );
  NAND U29075 ( .A(n53650), .B(n12772), .Z(n12773) );
  ANDN U29076 ( .B(x[1566]), .A(y[1566]), .Z(n53647) );
  OR U29077 ( .A(n12773), .B(n53647), .Z(n12774) );
  AND U29078 ( .A(n12775), .B(n12774), .Z(n12776) );
  OR U29079 ( .A(n53655), .B(n12776), .Z(n12777) );
  NAND U29080 ( .A(n53657), .B(n12777), .Z(n12778) );
  NANDN U29081 ( .A(n53659), .B(n12778), .Z(n12779) );
  NAND U29082 ( .A(n53661), .B(n12779), .Z(n12780) );
  NANDN U29083 ( .A(n53663), .B(n12780), .Z(n12781) );
  AND U29084 ( .A(n53665), .B(n12781), .Z(n12782) );
  OR U29085 ( .A(n53667), .B(n12782), .Z(n12783) );
  NAND U29086 ( .A(n53669), .B(n12783), .Z(n12784) );
  NANDN U29087 ( .A(n53671), .B(n12784), .Z(n12785) );
  NAND U29088 ( .A(n53673), .B(n12785), .Z(n12786) );
  NANDN U29089 ( .A(n53675), .B(n12786), .Z(n12787) );
  AND U29090 ( .A(n53676), .B(n12787), .Z(n12788) );
  OR U29091 ( .A(n53677), .B(n12788), .Z(n12789) );
  NAND U29092 ( .A(n53678), .B(n12789), .Z(n12790) );
  NAND U29093 ( .A(n33489), .B(n12790), .Z(n12791) );
  NANDN U29094 ( .A(n27711), .B(n12791), .Z(n12792) );
  NAND U29095 ( .A(n53681), .B(n12792), .Z(n12793) );
  NANDN U29096 ( .A(n53684), .B(n12793), .Z(n12794) );
  NANDN U29097 ( .A(n52249), .B(n12794), .Z(n12795) );
  AND U29098 ( .A(n53685), .B(n12795), .Z(n12797) );
  ANDN U29099 ( .B(x[1588]), .A(y[1588]), .Z(n33504) );
  IV U29100 ( .A(n33504), .Z(n53686) );
  ANDN U29101 ( .B(x[1589]), .A(y[1589]), .Z(n52247) );
  ANDN U29102 ( .B(n53686), .A(n52247), .Z(n12796) );
  NANDN U29103 ( .A(n12797), .B(n12796), .Z(n12798) );
  NAND U29104 ( .A(n33509), .B(n12798), .Z(n12799) );
  NANDN U29105 ( .A(n33510), .B(n12799), .Z(n12800) );
  NAND U29106 ( .A(n53691), .B(n12800), .Z(n12801) );
  NANDN U29107 ( .A(n33513), .B(n12801), .Z(n12804) );
  NANDN U29108 ( .A(x[1594]), .B(y[1594]), .Z(n12803) );
  NANDN U29109 ( .A(x[1593]), .B(y[1593]), .Z(n12802) );
  NAND U29110 ( .A(n12803), .B(n12802), .Z(n53694) );
  ANDN U29111 ( .B(n12804), .A(n53694), .Z(n12805) );
  OR U29112 ( .A(n53695), .B(n12805), .Z(n12806) );
  NAND U29113 ( .A(n53696), .B(n12806), .Z(n12807) );
  NANDN U29114 ( .A(n53697), .B(n12807), .Z(n12808) );
  ANDN U29115 ( .B(y[1597]), .A(x[1597]), .Z(n53698) );
  ANDN U29116 ( .B(n12808), .A(n53698), .Z(n12809) );
  NAND U29117 ( .A(n33527), .B(n12809), .Z(n12810) );
  NAND U29118 ( .A(n53699), .B(n12810), .Z(n12811) );
  ANDN U29119 ( .B(x[1599]), .A(y[1599]), .Z(n27704) );
  OR U29120 ( .A(n12811), .B(n27704), .Z(n12812) );
  AND U29121 ( .A(n33528), .B(n12812), .Z(n12813) );
  NANDN U29122 ( .A(n27702), .B(n12813), .Z(n12814) );
  NAND U29123 ( .A(n12815), .B(n12814), .Z(n12816) );
  ANDN U29124 ( .B(y[1602]), .A(x[1602]), .Z(n53703) );
  ANDN U29125 ( .B(n12816), .A(n53703), .Z(n12817) );
  NAND U29126 ( .A(n27703), .B(n12817), .Z(n12818) );
  NAND U29127 ( .A(n53704), .B(n12818), .Z(n12819) );
  ANDN U29128 ( .B(x[1602]), .A(y[1602]), .Z(n27700) );
  OR U29129 ( .A(n12819), .B(n27700), .Z(n12820) );
  AND U29130 ( .A(n53705), .B(n12820), .Z(n12821) );
  OR U29131 ( .A(n53706), .B(n12821), .Z(n12822) );
  NAND U29132 ( .A(n53707), .B(n12822), .Z(n12823) );
  NAND U29133 ( .A(n53708), .B(n12823), .Z(n12824) );
  ANDN U29134 ( .B(x[1607]), .A(y[1607]), .Z(n27698) );
  OR U29135 ( .A(n12824), .B(n27698), .Z(n12825) );
  AND U29136 ( .A(n27699), .B(n12825), .Z(n12826) );
  NANDN U29137 ( .A(n53710), .B(n12826), .Z(n12828) );
  ANDN U29138 ( .B(x[1608]), .A(y[1608]), .Z(n12827) );
  ANDN U29139 ( .B(n12828), .A(n12827), .Z(n12829) );
  NAND U29140 ( .A(n53713), .B(n12829), .Z(n12830) );
  NANDN U29141 ( .A(x[1609]), .B(y[1609]), .Z(n33550) );
  AND U29142 ( .A(n12830), .B(n33550), .Z(n12831) );
  NANDN U29143 ( .A(n53714), .B(n12831), .Z(n12832) );
  NANDN U29144 ( .A(n53715), .B(n12832), .Z(n12833) );
  NAND U29145 ( .A(n53716), .B(n12833), .Z(n12834) );
  NANDN U29146 ( .A(n53717), .B(n12834), .Z(n12835) );
  AND U29147 ( .A(n53718), .B(n12835), .Z(n12836) );
  OR U29148 ( .A(n53719), .B(n12836), .Z(n12837) );
  NAND U29149 ( .A(n53720), .B(n12837), .Z(n12838) );
  NANDN U29150 ( .A(n53721), .B(n12838), .Z(n12839) );
  NAND U29151 ( .A(n53722), .B(n12839), .Z(n12840) );
  NANDN U29152 ( .A(n53723), .B(n12840), .Z(n12841) );
  AND U29153 ( .A(n53724), .B(n12841), .Z(n12842) );
  OR U29154 ( .A(n53725), .B(n12842), .Z(n12843) );
  NAND U29155 ( .A(n53726), .B(n12843), .Z(n12844) );
  NANDN U29156 ( .A(n53727), .B(n12844), .Z(n12845) );
  NAND U29157 ( .A(n53728), .B(n12845), .Z(n12846) );
  NANDN U29158 ( .A(n53730), .B(n12846), .Z(n12847) );
  AND U29159 ( .A(n53731), .B(n12847), .Z(n12848) );
  OR U29160 ( .A(n53732), .B(n12848), .Z(n12849) );
  NAND U29161 ( .A(n53733), .B(n12849), .Z(n12850) );
  NANDN U29162 ( .A(n53734), .B(n12850), .Z(n12851) );
  NAND U29163 ( .A(n53735), .B(n12851), .Z(n12852) );
  AND U29164 ( .A(n12853), .B(n12852), .Z(n12854) );
  ANDN U29165 ( .B(y[1631]), .A(x[1631]), .Z(n33629) );
  NANDN U29166 ( .A(x[1632]), .B(y[1632]), .Z(n27689) );
  IV U29167 ( .A(n27689), .Z(n53739) );
  OR U29168 ( .A(n33629), .B(n53739), .Z(n53737) );
  OR U29169 ( .A(n12854), .B(n53737), .Z(n12855) );
  AND U29170 ( .A(n53738), .B(n12855), .Z(n12856) );
  NANDN U29171 ( .A(n27690), .B(n12856), .Z(n12857) );
  NAND U29172 ( .A(n53741), .B(n12857), .Z(n12858) );
  NANDN U29173 ( .A(n52245), .B(n12858), .Z(n12859) );
  NAND U29174 ( .A(n53742), .B(n12859), .Z(n12860) );
  ANDN U29175 ( .B(x[1637]), .A(y[1637]), .Z(n33648) );
  ANDN U29176 ( .B(n12860), .A(n33648), .Z(n12861) );
  NANDN U29177 ( .A(n52244), .B(n12861), .Z(n12862) );
  NANDN U29178 ( .A(x[1637]), .B(y[1637]), .Z(n52243) );
  AND U29179 ( .A(n12862), .B(n52243), .Z(n12863) );
  NAND U29180 ( .A(n27685), .B(n12863), .Z(n12864) );
  NANDN U29181 ( .A(n33647), .B(n12864), .Z(n12865) );
  ANDN U29182 ( .B(x[1639]), .A(y[1639]), .Z(n27684) );
  OR U29183 ( .A(n12865), .B(n27684), .Z(n12866) );
  AND U29184 ( .A(n27686), .B(n12866), .Z(n12867) );
  NANDN U29185 ( .A(x[1640]), .B(y[1640]), .Z(n27682) );
  NAND U29186 ( .A(n12867), .B(n27682), .Z(n12868) );
  ANDN U29187 ( .B(x[1641]), .A(y[1641]), .Z(n27679) );
  ANDN U29188 ( .B(n12868), .A(n27679), .Z(n12869) );
  NANDN U29189 ( .A(n27683), .B(n12869), .Z(n12870) );
  NANDN U29190 ( .A(x[1641]), .B(y[1641]), .Z(n27681) );
  AND U29191 ( .A(n12870), .B(n27681), .Z(n12871) );
  NAND U29192 ( .A(n52241), .B(n12871), .Z(n12872) );
  NANDN U29193 ( .A(n53748), .B(n12872), .Z(n12873) );
  NAND U29194 ( .A(n53749), .B(n12873), .Z(n12874) );
  NANDN U29195 ( .A(n52240), .B(n12874), .Z(n12875) );
  NANDN U29196 ( .A(x[1645]), .B(y[1645]), .Z(n27674) );
  NANDN U29197 ( .A(x[1646]), .B(y[1646]), .Z(n33666) );
  AND U29198 ( .A(n27674), .B(n33666), .Z(n52239) );
  AND U29199 ( .A(n12875), .B(n52239), .Z(n12878) );
  NANDN U29200 ( .A(y[1648]), .B(x[1648]), .Z(n12882) );
  NANDN U29201 ( .A(y[1647]), .B(x[1647]), .Z(n12876) );
  AND U29202 ( .A(n12882), .B(n12876), .Z(n33668) );
  NANDN U29203 ( .A(y[1646]), .B(x[1646]), .Z(n12877) );
  NAND U29204 ( .A(n33668), .B(n12877), .Z(n52238) );
  OR U29205 ( .A(n12878), .B(n52238), .Z(n12885) );
  XNOR U29206 ( .A(y[1648]), .B(x[1648]), .Z(n12880) );
  NANDN U29207 ( .A(x[1647]), .B(y[1647]), .Z(n12879) );
  NAND U29208 ( .A(n12880), .B(n12879), .Z(n12881) );
  NAND U29209 ( .A(n12882), .B(n12881), .Z(n12884) );
  NANDN U29210 ( .A(x[1649]), .B(y[1649]), .Z(n12883) );
  NAND U29211 ( .A(n12884), .B(n12883), .Z(n53750) );
  ANDN U29212 ( .B(n12885), .A(n53750), .Z(n12886) );
  OR U29213 ( .A(n53752), .B(n12886), .Z(n12887) );
  NAND U29214 ( .A(n53754), .B(n12887), .Z(n12888) );
  NANDN U29215 ( .A(n53756), .B(n12888), .Z(n12889) );
  NAND U29216 ( .A(n53758), .B(n12889), .Z(n12890) );
  NANDN U29217 ( .A(n53760), .B(n12890), .Z(n12891) );
  AND U29218 ( .A(n53762), .B(n12891), .Z(n12892) );
  OR U29219 ( .A(n53764), .B(n12892), .Z(n12893) );
  NAND U29220 ( .A(n53766), .B(n12893), .Z(n12894) );
  NANDN U29221 ( .A(n53768), .B(n12894), .Z(n12895) );
  NAND U29222 ( .A(n53770), .B(n12895), .Z(n12896) );
  NANDN U29223 ( .A(n53772), .B(n12896), .Z(n12897) );
  AND U29224 ( .A(n53774), .B(n12897), .Z(n12898) );
  NANDN U29225 ( .A(y[1660]), .B(x[1660]), .Z(n33694) );
  NANDN U29226 ( .A(y[1661]), .B(x[1661]), .Z(n27658) );
  NAND U29227 ( .A(n33694), .B(n27658), .Z(n53776) );
  OR U29228 ( .A(n12898), .B(n53776), .Z(n12899) );
  ANDN U29229 ( .B(y[1661]), .A(x[1661]), .Z(n52236) );
  ANDN U29230 ( .B(n12899), .A(n52236), .Z(n12900) );
  NANDN U29231 ( .A(y[1662]), .B(x[1662]), .Z(n53780) );
  NANDN U29232 ( .A(n12900), .B(n53780), .Z(n12901) );
  NANDN U29233 ( .A(x[1662]), .B(y[1662]), .Z(n52237) );
  NANDN U29234 ( .A(x[1663]), .B(y[1663]), .Z(n53785) );
  NAND U29235 ( .A(n52237), .B(n53785), .Z(n33703) );
  ANDN U29236 ( .B(n12901), .A(n33703), .Z(n12902) );
  NANDN U29237 ( .A(y[1663]), .B(x[1663]), .Z(n53779) );
  NANDN U29238 ( .A(n12902), .B(n53779), .Z(n12903) );
  NANDN U29239 ( .A(n53783), .B(n12903), .Z(n12904) );
  NANDN U29240 ( .A(n53788), .B(n12904), .Z(n12905) );
  NAND U29241 ( .A(n53790), .B(n12905), .Z(n12906) );
  NANDN U29242 ( .A(n53791), .B(n12906), .Z(n12907) );
  AND U29243 ( .A(n53792), .B(n12907), .Z(n12908) );
  OR U29244 ( .A(n53793), .B(n12908), .Z(n12909) );
  NAND U29245 ( .A(n53794), .B(n12909), .Z(n12910) );
  NANDN U29246 ( .A(n53795), .B(n12910), .Z(n12911) );
  NAND U29247 ( .A(n53796), .B(n12911), .Z(n12912) );
  NANDN U29248 ( .A(y[1673]), .B(x[1673]), .Z(n27648) );
  AND U29249 ( .A(n12912), .B(n27648), .Z(n12913) );
  NAND U29250 ( .A(n53797), .B(n12913), .Z(n12914) );
  ANDN U29251 ( .B(y[1673]), .A(x[1673]), .Z(n53798) );
  ANDN U29252 ( .B(n12914), .A(n53798), .Z(n12915) );
  NAND U29253 ( .A(n33732), .B(n12915), .Z(n12916) );
  NAND U29254 ( .A(n53800), .B(n12916), .Z(n12917) );
  ANDN U29255 ( .B(x[1674]), .A(y[1674]), .Z(n27647) );
  OR U29256 ( .A(n12917), .B(n27647), .Z(n12918) );
  AND U29257 ( .A(n12919), .B(n12918), .Z(n12920) );
  OR U29258 ( .A(n53802), .B(n12920), .Z(n12921) );
  NAND U29259 ( .A(n53803), .B(n12921), .Z(n12922) );
  NANDN U29260 ( .A(n53804), .B(n12922), .Z(n12923) );
  NAND U29261 ( .A(n53805), .B(n12923), .Z(n12924) );
  NANDN U29262 ( .A(n53806), .B(n12924), .Z(n12925) );
  AND U29263 ( .A(n53808), .B(n12925), .Z(n12926) );
  OR U29264 ( .A(n53809), .B(n12926), .Z(n12927) );
  NAND U29265 ( .A(n53810), .B(n12927), .Z(n12928) );
  NANDN U29266 ( .A(n53811), .B(n12928), .Z(n12929) );
  ANDN U29267 ( .B(x[1685]), .A(y[1685]), .Z(n27638) );
  OR U29268 ( .A(n12929), .B(n27638), .Z(n12930) );
  AND U29269 ( .A(n53814), .B(n12930), .Z(n12931) );
  NANDN U29270 ( .A(n27641), .B(n12931), .Z(n12932) );
  AND U29271 ( .A(n12933), .B(n12932), .Z(n12934) );
  NANDN U29272 ( .A(x[1687]), .B(y[1687]), .Z(n27637) );
  NANDN U29273 ( .A(x[1688]), .B(y[1688]), .Z(n27636) );
  NAND U29274 ( .A(n27637), .B(n27636), .Z(n52233) );
  OR U29275 ( .A(n12934), .B(n52233), .Z(n12935) );
  NANDN U29276 ( .A(y[1688]), .B(x[1688]), .Z(n52232) );
  AND U29277 ( .A(n12935), .B(n52232), .Z(n12936) );
  NANDN U29278 ( .A(n27635), .B(n12936), .Z(n12937) );
  AND U29279 ( .A(n27632), .B(n12937), .Z(n12938) );
  NANDN U29280 ( .A(x[1689]), .B(y[1689]), .Z(n52234) );
  NAND U29281 ( .A(n12938), .B(n52234), .Z(n12939) );
  ANDN U29282 ( .B(x[1691]), .A(y[1691]), .Z(n27630) );
  ANDN U29283 ( .B(n12939), .A(n27630), .Z(n12940) );
  NANDN U29284 ( .A(n27634), .B(n12940), .Z(n12941) );
  NANDN U29285 ( .A(x[1692]), .B(y[1692]), .Z(n53819) );
  AND U29286 ( .A(n12941), .B(n53819), .Z(n12942) );
  NAND U29287 ( .A(n27633), .B(n12942), .Z(n12943) );
  NAND U29288 ( .A(n53820), .B(n12943), .Z(n12944) );
  NANDN U29289 ( .A(y[1692]), .B(x[1692]), .Z(n27631) );
  NANDN U29290 ( .A(n12944), .B(n27631), .Z(n12945) );
  AND U29291 ( .A(n53821), .B(n12945), .Z(n12946) );
  NANDN U29292 ( .A(y[1694]), .B(x[1694]), .Z(n33778) );
  NANDN U29293 ( .A(y[1695]), .B(x[1695]), .Z(n33784) );
  AND U29294 ( .A(n33778), .B(n33784), .Z(n53822) );
  NANDN U29295 ( .A(n12946), .B(n53822), .Z(n12947) );
  NANDN U29296 ( .A(n52231), .B(n12947), .Z(n12948) );
  NANDN U29297 ( .A(y[1696]), .B(x[1696]), .Z(n33783) );
  NANDN U29298 ( .A(y[1697]), .B(x[1697]), .Z(n33790) );
  AND U29299 ( .A(n33783), .B(n33790), .Z(n52230) );
  AND U29300 ( .A(n12948), .B(n52230), .Z(n12949) );
  NANDN U29301 ( .A(x[1697]), .B(y[1697]), .Z(n27625) );
  NANDN U29302 ( .A(x[1698]), .B(y[1698]), .Z(n27624) );
  NAND U29303 ( .A(n27625), .B(n27624), .Z(n52229) );
  OR U29304 ( .A(n12949), .B(n52229), .Z(n12950) );
  NAND U29305 ( .A(n52228), .B(n12950), .Z(n12951) );
  NANDN U29306 ( .A(n53825), .B(n12951), .Z(n12952) );
  NAND U29307 ( .A(n53826), .B(n12952), .Z(n12953) );
  NANDN U29308 ( .A(n52227), .B(n12953), .Z(n12954) );
  NANDN U29309 ( .A(y[1702]), .B(x[1702]), .Z(n33801) );
  NANDN U29310 ( .A(y[1703]), .B(x[1703]), .Z(n33808) );
  AND U29311 ( .A(n33801), .B(n33808), .Z(n52226) );
  AND U29312 ( .A(n12954), .B(n52226), .Z(n12955) );
  NANDN U29313 ( .A(x[1703]), .B(y[1703]), .Z(n27619) );
  NANDN U29314 ( .A(x[1704]), .B(y[1704]), .Z(n27618) );
  NAND U29315 ( .A(n27619), .B(n27618), .Z(n52225) );
  OR U29316 ( .A(n12955), .B(n52225), .Z(n12956) );
  NAND U29317 ( .A(n53827), .B(n12956), .Z(n12957) );
  NANDN U29318 ( .A(n53828), .B(n12957), .Z(n12958) );
  NAND U29319 ( .A(n53829), .B(n12958), .Z(n12959) );
  NANDN U29320 ( .A(n52224), .B(n12959), .Z(n12960) );
  AND U29321 ( .A(n53832), .B(n12960), .Z(n12961) );
  ANDN U29322 ( .B(y[1709]), .A(x[1709]), .Z(n33824) );
  NANDN U29323 ( .A(x[1710]), .B(y[1710]), .Z(n27613) );
  NANDN U29324 ( .A(n33824), .B(n27613), .Z(n52223) );
  OR U29325 ( .A(n12961), .B(n52223), .Z(n12962) );
  NAND U29326 ( .A(n53833), .B(n12962), .Z(n12963) );
  NANDN U29327 ( .A(n53834), .B(n12963), .Z(n12964) );
  NANDN U29328 ( .A(n52222), .B(n12964), .Z(n12965) );
  AND U29329 ( .A(n53835), .B(n12965), .Z(n12967) );
  NANDN U29330 ( .A(y[1714]), .B(x[1714]), .Z(n53836) );
  ANDN U29331 ( .B(x[1715]), .A(y[1715]), .Z(n27608) );
  ANDN U29332 ( .B(n53836), .A(n27608), .Z(n12966) );
  NANDN U29333 ( .A(n12967), .B(n12966), .Z(n12968) );
  NANDN U29334 ( .A(n12969), .B(n12968), .Z(n12971) );
  NANDN U29335 ( .A(y[1716]), .B(x[1716]), .Z(n27609) );
  NANDN U29336 ( .A(y[1717]), .B(x[1717]), .Z(n52220) );
  AND U29337 ( .A(n27609), .B(n52220), .Z(n12970) );
  NAND U29338 ( .A(n12971), .B(n12970), .Z(n12972) );
  AND U29339 ( .A(n53839), .B(n12972), .Z(n12973) );
  OR U29340 ( .A(n53840), .B(n12973), .Z(n12974) );
  NAND U29341 ( .A(n53842), .B(n12974), .Z(n12975) );
  NANDN U29342 ( .A(n27605), .B(n12975), .Z(n12976) );
  ANDN U29343 ( .B(x[1721]), .A(y[1721]), .Z(n27600) );
  OR U29344 ( .A(n12976), .B(n27600), .Z(n12977) );
  NAND U29345 ( .A(n27604), .B(n12977), .Z(n12978) );
  NANDN U29346 ( .A(n27603), .B(n12978), .Z(n12981) );
  NANDN U29347 ( .A(y[1722]), .B(x[1722]), .Z(n27601) );
  NANDN U29348 ( .A(n27601), .B(n12979), .Z(n12980) );
  NANDN U29349 ( .A(n12981), .B(n12980), .Z(n12984) );
  NANDN U29350 ( .A(x[1724]), .B(y[1724]), .Z(n12983) );
  NANDN U29351 ( .A(x[1725]), .B(y[1725]), .Z(n12982) );
  NAND U29352 ( .A(n12983), .B(n12982), .Z(n53846) );
  ANDN U29353 ( .B(n12984), .A(n53846), .Z(n12985) );
  NANDN U29354 ( .A(y[1725]), .B(x[1725]), .Z(n53847) );
  NANDN U29355 ( .A(n12985), .B(n53847), .Z(n12986) );
  NANDN U29356 ( .A(n53848), .B(n12986), .Z(n12987) );
  NANDN U29357 ( .A(n53849), .B(n12987), .Z(n12988) );
  XOR U29358 ( .A(x[1728]), .B(y[1728]), .Z(n27598) );
  ANDN U29359 ( .B(n12988), .A(n27598), .Z(n12989) );
  NANDN U29360 ( .A(n53850), .B(n12989), .Z(n12990) );
  NANDN U29361 ( .A(n53852), .B(n12990), .Z(n12991) );
  NAND U29362 ( .A(n53853), .B(n12991), .Z(n12992) );
  NANDN U29363 ( .A(n53854), .B(n12992), .Z(n12993) );
  AND U29364 ( .A(n53855), .B(n12993), .Z(n12994) );
  ANDN U29365 ( .B(x[1732]), .A(y[1732]), .Z(n33879) );
  NANDN U29366 ( .A(y[1733]), .B(x[1733]), .Z(n27593) );
  NANDN U29367 ( .A(n33879), .B(n27593), .Z(n53856) );
  OR U29368 ( .A(n12994), .B(n53856), .Z(n12995) );
  NANDN U29369 ( .A(x[1733]), .B(y[1733]), .Z(n27594) );
  AND U29370 ( .A(n12995), .B(n27594), .Z(n12996) );
  NANDN U29371 ( .A(x[1734]), .B(y[1734]), .Z(n27591) );
  NAND U29372 ( .A(n12996), .B(n27591), .Z(n12997) );
  NANDN U29373 ( .A(y[1735]), .B(x[1735]), .Z(n27589) );
  AND U29374 ( .A(n12997), .B(n27589), .Z(n12998) );
  NANDN U29375 ( .A(n27592), .B(n12998), .Z(n12999) );
  NANDN U29376 ( .A(x[1735]), .B(y[1735]), .Z(n27590) );
  AND U29377 ( .A(n12999), .B(n27590), .Z(n13000) );
  NAND U29378 ( .A(n33889), .B(n13000), .Z(n13001) );
  NAND U29379 ( .A(n53863), .B(n13001), .Z(n13002) );
  ANDN U29380 ( .B(x[1736]), .A(y[1736]), .Z(n27588) );
  OR U29381 ( .A(n13002), .B(n27588), .Z(n13003) );
  AND U29382 ( .A(n33888), .B(n13003), .Z(n13004) );
  NANDN U29383 ( .A(n52219), .B(n13004), .Z(n13005) );
  NANDN U29384 ( .A(y[1739]), .B(x[1739]), .Z(n33894) );
  NANDN U29385 ( .A(y[1738]), .B(x[1738]), .Z(n27587) );
  AND U29386 ( .A(n33894), .B(n27587), .Z(n52218) );
  AND U29387 ( .A(n13005), .B(n52218), .Z(n13008) );
  NANDN U29388 ( .A(x[1739]), .B(y[1739]), .Z(n13007) );
  NANDN U29389 ( .A(x[1740]), .B(y[1740]), .Z(n13006) );
  NAND U29390 ( .A(n13007), .B(n13006), .Z(n52217) );
  OR U29391 ( .A(n13008), .B(n52217), .Z(n13011) );
  NANDN U29392 ( .A(y[1741]), .B(x[1741]), .Z(n13010) );
  NANDN U29393 ( .A(y[1740]), .B(x[1740]), .Z(n13009) );
  AND U29394 ( .A(n13010), .B(n13009), .Z(n52216) );
  AND U29395 ( .A(n13011), .B(n52216), .Z(n13014) );
  NANDN U29396 ( .A(x[1741]), .B(y[1741]), .Z(n13013) );
  NANDN U29397 ( .A(x[1742]), .B(y[1742]), .Z(n13012) );
  NAND U29398 ( .A(n13013), .B(n13012), .Z(n53864) );
  OR U29399 ( .A(n13014), .B(n53864), .Z(n13015) );
  NAND U29400 ( .A(n53865), .B(n13015), .Z(n13016) );
  NANDN U29401 ( .A(n52215), .B(n13016), .Z(n13017) );
  NAND U29402 ( .A(n52214), .B(n13017), .Z(n13018) );
  NAND U29403 ( .A(n53868), .B(n13018), .Z(n13019) );
  NANDN U29404 ( .A(n53869), .B(n13019), .Z(n13020) );
  NANDN U29405 ( .A(n53871), .B(n13020), .Z(n13021) );
  AND U29406 ( .A(n53872), .B(n13021), .Z(n13026) );
  NANDN U29407 ( .A(x[1748]), .B(y[1748]), .Z(n53870) );
  OR U29408 ( .A(n13022), .B(n53870), .Z(n13025) );
  NANDN U29409 ( .A(x[1750]), .B(y[1750]), .Z(n13024) );
  NANDN U29410 ( .A(x[1749]), .B(y[1749]), .Z(n13023) );
  AND U29411 ( .A(n13024), .B(n13023), .Z(n53873) );
  AND U29412 ( .A(n13025), .B(n53873), .Z(n33913) );
  NANDN U29413 ( .A(n13026), .B(n33913), .Z(n13027) );
  NANDN U29414 ( .A(n33914), .B(n13027), .Z(n13032) );
  XNOR U29415 ( .A(y[1752]), .B(x[1752]), .Z(n13029) );
  NANDN U29416 ( .A(x[1751]), .B(y[1751]), .Z(n13028) );
  NAND U29417 ( .A(n13029), .B(n13028), .Z(n13030) );
  NAND U29418 ( .A(n13031), .B(n13030), .Z(n52213) );
  AND U29419 ( .A(n13032), .B(n52213), .Z(n13033) );
  ANDN U29420 ( .B(x[1753]), .A(y[1753]), .Z(n27584) );
  OR U29421 ( .A(n13033), .B(n27584), .Z(n13034) );
  NAND U29422 ( .A(n53876), .B(n13034), .Z(n13035) );
  NANDN U29423 ( .A(n53877), .B(n13035), .Z(n13036) );
  NAND U29424 ( .A(n53878), .B(n13036), .Z(n13037) );
  ANDN U29425 ( .B(x[1757]), .A(y[1757]), .Z(n27578) );
  ANDN U29426 ( .B(n13037), .A(n27578), .Z(n13038) );
  NANDN U29427 ( .A(n53879), .B(n13038), .Z(n13040) );
  NANDN U29428 ( .A(x[1757]), .B(y[1757]), .Z(n53880) );
  NANDN U29429 ( .A(x[1758]), .B(y[1758]), .Z(n53883) );
  AND U29430 ( .A(n53880), .B(n53883), .Z(n13039) );
  NAND U29431 ( .A(n13040), .B(n13039), .Z(n13041) );
  NANDN U29432 ( .A(y[1759]), .B(x[1759]), .Z(n33932) );
  AND U29433 ( .A(n13041), .B(n33932), .Z(n13042) );
  NANDN U29434 ( .A(y[1758]), .B(x[1758]), .Z(n27579) );
  NAND U29435 ( .A(n13042), .B(n27579), .Z(n13043) );
  NANDN U29436 ( .A(n53885), .B(n13043), .Z(n13044) );
  AND U29437 ( .A(n53886), .B(n13044), .Z(n13045) );
  OR U29438 ( .A(n53887), .B(n13045), .Z(n13046) );
  NAND U29439 ( .A(n53888), .B(n13046), .Z(n13047) );
  NANDN U29440 ( .A(n53889), .B(n13047), .Z(n13048) );
  NAND U29441 ( .A(n53890), .B(n13048), .Z(n13049) );
  NAND U29442 ( .A(n52212), .B(n13049), .Z(n13050) );
  NANDN U29443 ( .A(n53891), .B(n13050), .Z(n13051) );
  AND U29444 ( .A(n33949), .B(n13051), .Z(n13052) );
  OR U29445 ( .A(n53893), .B(n13052), .Z(n13053) );
  NAND U29446 ( .A(n33952), .B(n13053), .Z(n13054) );
  NANDN U29447 ( .A(n33954), .B(n13054), .Z(n13055) );
  NANDN U29448 ( .A(x[1770]), .B(y[1770]), .Z(n53895) );
  AND U29449 ( .A(n13055), .B(n53895), .Z(n13056) );
  NAND U29450 ( .A(n33951), .B(n13056), .Z(n13057) );
  NANDN U29451 ( .A(n52209), .B(n13057), .Z(n13058) );
  ANDN U29452 ( .B(x[1770]), .A(y[1770]), .Z(n33955) );
  OR U29453 ( .A(n13058), .B(n33955), .Z(n13059) );
  NAND U29454 ( .A(n53897), .B(n13059), .Z(n13060) );
  NANDN U29455 ( .A(n53898), .B(n13060), .Z(n13061) );
  AND U29456 ( .A(n53899), .B(n13061), .Z(n13063) );
  NANDN U29457 ( .A(y[1774]), .B(x[1774]), .Z(n53900) );
  ANDN U29458 ( .B(x[1775]), .A(y[1775]), .Z(n27564) );
  ANDN U29459 ( .B(n53900), .A(n27564), .Z(n13062) );
  NANDN U29460 ( .A(n13063), .B(n13062), .Z(n13064) );
  NANDN U29461 ( .A(n13065), .B(n13064), .Z(n13066) );
  NANDN U29462 ( .A(y[1776]), .B(x[1776]), .Z(n27565) );
  AND U29463 ( .A(n13066), .B(n27565), .Z(n13067) );
  NAND U29464 ( .A(n27562), .B(n13067), .Z(n13068) );
  NANDN U29465 ( .A(n53905), .B(n13068), .Z(n13069) );
  NAND U29466 ( .A(n53906), .B(n13069), .Z(n13070) );
  NANDN U29467 ( .A(n53907), .B(n13070), .Z(n13071) );
  AND U29468 ( .A(n53908), .B(n13071), .Z(n13072) );
  OR U29469 ( .A(n53909), .B(n13072), .Z(n13073) );
  NAND U29470 ( .A(n53910), .B(n13073), .Z(n13074) );
  NANDN U29471 ( .A(n53911), .B(n13074), .Z(n13075) );
  NAND U29472 ( .A(n52208), .B(n13075), .Z(n13076) );
  NANDN U29473 ( .A(n53912), .B(n13076), .Z(n13079) );
  NANDN U29474 ( .A(y[1787]), .B(x[1787]), .Z(n13078) );
  NANDN U29475 ( .A(y[1786]), .B(x[1786]), .Z(n13077) );
  AND U29476 ( .A(n13078), .B(n13077), .Z(n53913) );
  AND U29477 ( .A(n13079), .B(n53913), .Z(n13082) );
  NANDN U29478 ( .A(x[1787]), .B(y[1787]), .Z(n13081) );
  NANDN U29479 ( .A(x[1788]), .B(y[1788]), .Z(n13080) );
  NAND U29480 ( .A(n13081), .B(n13080), .Z(n53916) );
  OR U29481 ( .A(n13082), .B(n53916), .Z(n13083) );
  NAND U29482 ( .A(n53918), .B(n13083), .Z(n13084) );
  NANDN U29483 ( .A(n52207), .B(n13084), .Z(n13085) );
  NAND U29484 ( .A(n52206), .B(n13085), .Z(n13086) );
  NAND U29485 ( .A(n53919), .B(n13086), .Z(n13087) );
  NANDN U29486 ( .A(n52205), .B(n13087), .Z(n13088) );
  NAND U29487 ( .A(n52204), .B(n13088), .Z(n13089) );
  NANDN U29488 ( .A(n53920), .B(n13089), .Z(n13090) );
  AND U29489 ( .A(n53921), .B(n13090), .Z(n13092) );
  NANDN U29490 ( .A(y[1796]), .B(x[1796]), .Z(n13091) );
  ANDN U29491 ( .B(x[1797]), .A(y[1797]), .Z(n27551) );
  ANDN U29492 ( .B(n13091), .A(n27551), .Z(n53922) );
  NANDN U29493 ( .A(n13092), .B(n53922), .Z(n13093) );
  NAND U29494 ( .A(n53923), .B(n13093), .Z(n13094) );
  NANDN U29495 ( .A(n34005), .B(n13094), .Z(n13095) );
  NAND U29496 ( .A(n34007), .B(n13095), .Z(n13096) );
  NAND U29497 ( .A(n34008), .B(n13096), .Z(n13097) );
  NANDN U29498 ( .A(n34010), .B(n13097), .Z(n13098) );
  NAND U29499 ( .A(n53931), .B(n13098), .Z(n13099) );
  NANDN U29500 ( .A(n53932), .B(n13099), .Z(n13100) );
  NANDN U29501 ( .A(y[1804]), .B(x[1804]), .Z(n34018) );
  AND U29502 ( .A(n13100), .B(n34018), .Z(n13101) );
  NANDN U29503 ( .A(y[1805]), .B(x[1805]), .Z(n27546) );
  NAND U29504 ( .A(n13101), .B(n27546), .Z(n13102) );
  ANDN U29505 ( .B(y[1805]), .A(x[1805]), .Z(n27548) );
  ANDN U29506 ( .B(n13102), .A(n27548), .Z(n13103) );
  NANDN U29507 ( .A(n27545), .B(n13103), .Z(n13105) );
  NANDN U29508 ( .A(y[1806]), .B(x[1806]), .Z(n13104) );
  AND U29509 ( .A(n13105), .B(n13104), .Z(n13106) );
  NAND U29510 ( .A(n27541), .B(n13106), .Z(n13107) );
  NANDN U29511 ( .A(n27542), .B(n13107), .Z(n13108) );
  ANDN U29512 ( .B(y[1808]), .A(x[1808]), .Z(n27539) );
  OR U29513 ( .A(n13108), .B(n27539), .Z(n13109) );
  NANDN U29514 ( .A(y[1809]), .B(x[1809]), .Z(n53939) );
  AND U29515 ( .A(n13109), .B(n53939), .Z(n13110) );
  NANDN U29516 ( .A(n13111), .B(n13110), .Z(n13112) );
  AND U29517 ( .A(n27540), .B(n13112), .Z(n13113) );
  NANDN U29518 ( .A(x[1810]), .B(y[1810]), .Z(n53940) );
  NAND U29519 ( .A(n13113), .B(n53940), .Z(n13114) );
  NANDN U29520 ( .A(n53941), .B(n13114), .Z(n13115) );
  AND U29521 ( .A(n53942), .B(n13115), .Z(n13116) );
  OR U29522 ( .A(n53944), .B(n13116), .Z(n13117) );
  NAND U29523 ( .A(n53945), .B(n13117), .Z(n13118) );
  NANDN U29524 ( .A(n53946), .B(n13118), .Z(n13119) );
  NANDN U29525 ( .A(n52202), .B(n13119), .Z(n13120) );
  NANDN U29526 ( .A(y[1816]), .B(x[1816]), .Z(n34043) );
  NANDN U29527 ( .A(y[1817]), .B(x[1817]), .Z(n27532) );
  AND U29528 ( .A(n34043), .B(n27532), .Z(n52201) );
  AND U29529 ( .A(n13120), .B(n52201), .Z(n13122) );
  NANDN U29530 ( .A(x[1818]), .B(y[1818]), .Z(n34051) );
  ANDN U29531 ( .B(y[1817]), .A(x[1817]), .Z(n52200) );
  ANDN U29532 ( .B(n34051), .A(n52200), .Z(n13121) );
  NANDN U29533 ( .A(n13122), .B(n13121), .Z(n13123) );
  NAND U29534 ( .A(n53947), .B(n13123), .Z(n13124) );
  ANDN U29535 ( .B(x[1819]), .A(y[1819]), .Z(n27529) );
  OR U29536 ( .A(n13124), .B(n27529), .Z(n13125) );
  NAND U29537 ( .A(n13126), .B(n13125), .Z(n13127) );
  NANDN U29538 ( .A(y[1820]), .B(x[1820]), .Z(n27530) );
  AND U29539 ( .A(n13127), .B(n27530), .Z(n13128) );
  NAND U29540 ( .A(n27525), .B(n13128), .Z(n13129) );
  NANDN U29541 ( .A(n27526), .B(n13129), .Z(n13130) );
  ANDN U29542 ( .B(y[1822]), .A(x[1822]), .Z(n27522) );
  OR U29543 ( .A(n13130), .B(n27522), .Z(n13131) );
  NANDN U29544 ( .A(y[1823]), .B(x[1823]), .Z(n52199) );
  AND U29545 ( .A(n13131), .B(n52199), .Z(n13132) );
  NANDN U29546 ( .A(n27524), .B(n13132), .Z(n13133) );
  AND U29547 ( .A(n13134), .B(n13133), .Z(n13135) );
  OR U29548 ( .A(n53954), .B(n13135), .Z(n13136) );
  NAND U29549 ( .A(n53955), .B(n13136), .Z(n13137) );
  NANDN U29550 ( .A(n53957), .B(n13137), .Z(n13138) );
  NAND U29551 ( .A(n53958), .B(n13138), .Z(n13139) );
  NANDN U29552 ( .A(n53959), .B(n13139), .Z(n13140) );
  AND U29553 ( .A(n53960), .B(n13140), .Z(n13141) );
  OR U29554 ( .A(n53961), .B(n13141), .Z(n13142) );
  NAND U29555 ( .A(n53962), .B(n13142), .Z(n13143) );
  NANDN U29556 ( .A(n53963), .B(n13143), .Z(n13144) );
  NAND U29557 ( .A(n53964), .B(n13144), .Z(n13145) );
  NANDN U29558 ( .A(y[1835]), .B(x[1835]), .Z(n27516) );
  AND U29559 ( .A(n13145), .B(n27516), .Z(n13146) );
  NAND U29560 ( .A(n53965), .B(n13146), .Z(n13148) );
  NANDN U29561 ( .A(x[1835]), .B(y[1835]), .Z(n53966) );
  ANDN U29562 ( .B(y[1836]), .A(x[1836]), .Z(n53968) );
  ANDN U29563 ( .B(n53966), .A(n53968), .Z(n13147) );
  NAND U29564 ( .A(n13148), .B(n13147), .Z(n13149) );
  NANDN U29565 ( .A(y[1837]), .B(x[1837]), .Z(n53969) );
  AND U29566 ( .A(n13149), .B(n53969), .Z(n13150) );
  NANDN U29567 ( .A(n27515), .B(n13150), .Z(n13151) );
  AND U29568 ( .A(n53970), .B(n13151), .Z(n13152) );
  NANDN U29569 ( .A(y[1838]), .B(x[1838]), .Z(n34102) );
  NANDN U29570 ( .A(y[1839]), .B(x[1839]), .Z(n34109) );
  NAND U29571 ( .A(n34102), .B(n34109), .Z(n53971) );
  OR U29572 ( .A(n13152), .B(n53971), .Z(n13153) );
  AND U29573 ( .A(n53972), .B(n13153), .Z(n13155) );
  NANDN U29574 ( .A(y[1841]), .B(x[1841]), .Z(n27513) );
  ANDN U29575 ( .B(x[1840]), .A(y[1840]), .Z(n34108) );
  ANDN U29576 ( .B(n27513), .A(n34108), .Z(n13154) );
  NANDN U29577 ( .A(n13155), .B(n13154), .Z(n13156) );
  NANDN U29578 ( .A(n53974), .B(n13156), .Z(n13157) );
  XNOR U29579 ( .A(x[1842]), .B(y[1842]), .Z(n27514) );
  NANDN U29580 ( .A(n13157), .B(n27514), .Z(n13158) );
  AND U29581 ( .A(n13159), .B(n13158), .Z(n13160) );
  OR U29582 ( .A(n53979), .B(n13160), .Z(n13161) );
  NAND U29583 ( .A(n53980), .B(n13161), .Z(n13162) );
  NANDN U29584 ( .A(n53981), .B(n13162), .Z(n13163) );
  NAND U29585 ( .A(n53982), .B(n13163), .Z(n13164) );
  NANDN U29586 ( .A(n53983), .B(n13164), .Z(n13165) );
  AND U29587 ( .A(n53984), .B(n13165), .Z(n13167) );
  ANDN U29588 ( .B(y[1850]), .A(x[1850]), .Z(n27507) );
  ANDN U29589 ( .B(y[1849]), .A(x[1849]), .Z(n53985) );
  NOR U29590 ( .A(n27507), .B(n53985), .Z(n13166) );
  NANDN U29591 ( .A(n13167), .B(n13166), .Z(n13168) );
  ANDN U29592 ( .B(x[1850]), .A(y[1850]), .Z(n53986) );
  ANDN U29593 ( .B(n13168), .A(n53986), .Z(n13169) );
  NAND U29594 ( .A(n13170), .B(n13169), .Z(n13171) );
  NAND U29595 ( .A(n27508), .B(n13171), .Z(n13172) );
  AND U29596 ( .A(n34142), .B(n13172), .Z(n13175) );
  NANDN U29597 ( .A(x[1852]), .B(y[1852]), .Z(n13174) );
  NANDN U29598 ( .A(x[1853]), .B(y[1853]), .Z(n13173) );
  NAND U29599 ( .A(n13174), .B(n13173), .Z(n34144) );
  OR U29600 ( .A(n13175), .B(n34144), .Z(n13178) );
  NANDN U29601 ( .A(y[1854]), .B(x[1854]), .Z(n13177) );
  NANDN U29602 ( .A(y[1853]), .B(x[1853]), .Z(n13176) );
  AND U29603 ( .A(n13177), .B(n13176), .Z(n34146) );
  AND U29604 ( .A(n13178), .B(n34146), .Z(n13183) );
  NANDN U29605 ( .A(x[1855]), .B(y[1855]), .Z(n13180) );
  NANDN U29606 ( .A(x[1854]), .B(y[1854]), .Z(n13179) );
  AND U29607 ( .A(n13180), .B(n13179), .Z(n13182) );
  NANDN U29608 ( .A(x[1856]), .B(y[1856]), .Z(n13181) );
  AND U29609 ( .A(n13182), .B(n13181), .Z(n53990) );
  NANDN U29610 ( .A(n13183), .B(n53990), .Z(n13184) );
  NAND U29611 ( .A(n13185), .B(n13184), .Z(n13186) );
  NANDN U29612 ( .A(x[1857]), .B(y[1857]), .Z(n53992) );
  AND U29613 ( .A(n13186), .B(n53992), .Z(n13187) );
  NAND U29614 ( .A(n27504), .B(n13187), .Z(n13188) );
  NAND U29615 ( .A(n27506), .B(n13188), .Z(n13189) );
  ANDN U29616 ( .B(x[1859]), .A(y[1859]), .Z(n27501) );
  OR U29617 ( .A(n13189), .B(n27501), .Z(n13190) );
  NAND U29618 ( .A(n13191), .B(n13190), .Z(n13192) );
  NANDN U29619 ( .A(n13193), .B(n13192), .Z(n13194) );
  ANDN U29620 ( .B(x[1861]), .A(y[1861]), .Z(n53997) );
  OR U29621 ( .A(n13194), .B(n53997), .Z(n13195) );
  AND U29622 ( .A(n13196), .B(n13195), .Z(n13197) );
  OR U29623 ( .A(n53999), .B(n13197), .Z(n13198) );
  NAND U29624 ( .A(n54000), .B(n13198), .Z(n13199) );
  NANDN U29625 ( .A(n54001), .B(n13199), .Z(n13200) );
  NAND U29626 ( .A(n54002), .B(n13200), .Z(n13201) );
  NAND U29627 ( .A(n52196), .B(n13201), .Z(n13202) );
  NANDN U29628 ( .A(n54003), .B(n13202), .Z(n13203) );
  NANDN U29629 ( .A(y[1868]), .B(x[1868]), .Z(n27488) );
  NANDN U29630 ( .A(y[1869]), .B(x[1869]), .Z(n34175) );
  AND U29631 ( .A(n27488), .B(n34175), .Z(n54004) );
  AND U29632 ( .A(n13203), .B(n54004), .Z(n13204) );
  NANDN U29633 ( .A(x[1869]), .B(y[1869]), .Z(n27486) );
  NANDN U29634 ( .A(x[1870]), .B(y[1870]), .Z(n34177) );
  AND U29635 ( .A(n27486), .B(n34177), .Z(n54005) );
  NANDN U29636 ( .A(n13204), .B(n54005), .Z(n13205) );
  NANDN U29637 ( .A(n54006), .B(n13205), .Z(n13206) );
  AND U29638 ( .A(n54007), .B(n13206), .Z(n13207) );
  OR U29639 ( .A(n54009), .B(n13207), .Z(n13208) );
  NAND U29640 ( .A(n54010), .B(n13208), .Z(n13209) );
  NANDN U29641 ( .A(n54011), .B(n13209), .Z(n13210) );
  NANDN U29642 ( .A(n52195), .B(n13210), .Z(n13211) );
  NANDN U29643 ( .A(y[1876]), .B(x[1876]), .Z(n34192) );
  NANDN U29644 ( .A(y[1877]), .B(x[1877]), .Z(n34201) );
  AND U29645 ( .A(n34192), .B(n34201), .Z(n52194) );
  AND U29646 ( .A(n13211), .B(n52194), .Z(n13212) );
  ANDN U29647 ( .B(y[1878]), .A(x[1878]), .Z(n34204) );
  NANDN U29648 ( .A(x[1877]), .B(y[1877]), .Z(n27480) );
  NANDN U29649 ( .A(n34204), .B(n27480), .Z(n52193) );
  OR U29650 ( .A(n13212), .B(n52193), .Z(n13213) );
  NAND U29651 ( .A(n54012), .B(n13213), .Z(n13214) );
  NANDN U29652 ( .A(n54013), .B(n13214), .Z(n13215) );
  NANDN U29653 ( .A(n52192), .B(n13215), .Z(n13216) );
  AND U29654 ( .A(n54014), .B(n13216), .Z(n13218) );
  NANDN U29655 ( .A(y[1883]), .B(x[1883]), .Z(n27473) );
  ANDN U29656 ( .B(x[1882]), .A(y[1882]), .Z(n27476) );
  ANDN U29657 ( .B(n27473), .A(n27476), .Z(n13217) );
  NANDN U29658 ( .A(n13218), .B(n13217), .Z(n13219) );
  NANDN U29659 ( .A(n54018), .B(n13219), .Z(n13220) );
  NANDN U29660 ( .A(x[1883]), .B(y[1883]), .Z(n54016) );
  NANDN U29661 ( .A(n13220), .B(n54016), .Z(n13221) );
  AND U29662 ( .A(n13222), .B(n13221), .Z(n13223) );
  OR U29663 ( .A(n54020), .B(n13223), .Z(n13224) );
  NAND U29664 ( .A(n52191), .B(n13224), .Z(n13225) );
  NANDN U29665 ( .A(n54022), .B(n13225), .Z(n13227) );
  NANDN U29666 ( .A(y[1889]), .B(x[1889]), .Z(n27467) );
  NANDN U29667 ( .A(y[1888]), .B(x[1888]), .Z(n54023) );
  AND U29668 ( .A(n27467), .B(n54023), .Z(n13226) );
  NAND U29669 ( .A(n13227), .B(n13226), .Z(n13228) );
  AND U29670 ( .A(n54024), .B(n13228), .Z(n13229) );
  NANDN U29671 ( .A(x[1890]), .B(y[1890]), .Z(n27465) );
  NAND U29672 ( .A(n13229), .B(n27465), .Z(n13230) );
  ANDN U29673 ( .B(x[1891]), .A(y[1891]), .Z(n27462) );
  ANDN U29674 ( .B(n13230), .A(n27462), .Z(n13231) );
  NANDN U29675 ( .A(n27466), .B(n13231), .Z(n13232) );
  AND U29676 ( .A(n27464), .B(n13232), .Z(n13233) );
  NAND U29677 ( .A(n27463), .B(n13233), .Z(n13234) );
  NANDN U29678 ( .A(y[1893]), .B(x[1893]), .Z(n54029) );
  AND U29679 ( .A(n13234), .B(n54029), .Z(n13235) );
  NANDN U29680 ( .A(n13236), .B(n13235), .Z(n13237) );
  AND U29681 ( .A(n27459), .B(n13237), .Z(n13238) );
  NANDN U29682 ( .A(x[1893]), .B(y[1893]), .Z(n27460) );
  NAND U29683 ( .A(n13238), .B(n27460), .Z(n13239) );
  NANDN U29684 ( .A(n54031), .B(n13239), .Z(n13240) );
  AND U29685 ( .A(n54032), .B(n13240), .Z(n13241) );
  OR U29686 ( .A(n54033), .B(n13241), .Z(n13242) );
  NAND U29687 ( .A(n54034), .B(n13242), .Z(n13243) );
  NANDN U29688 ( .A(n54035), .B(n13243), .Z(n13244) );
  NANDN U29689 ( .A(n52190), .B(n13244), .Z(n13245) );
  NANDN U29690 ( .A(y[1901]), .B(x[1901]), .Z(n34257) );
  NANDN U29691 ( .A(y[1900]), .B(x[1900]), .Z(n27456) );
  AND U29692 ( .A(n34257), .B(n27456), .Z(n52189) );
  AND U29693 ( .A(n13245), .B(n52189), .Z(n13248) );
  NANDN U29694 ( .A(x[1901]), .B(y[1901]), .Z(n13247) );
  NANDN U29695 ( .A(x[1902]), .B(y[1902]), .Z(n13246) );
  NAND U29696 ( .A(n13247), .B(n13246), .Z(n52188) );
  OR U29697 ( .A(n13248), .B(n52188), .Z(n13251) );
  NANDN U29698 ( .A(y[1903]), .B(x[1903]), .Z(n13250) );
  NANDN U29699 ( .A(y[1902]), .B(x[1902]), .Z(n13249) );
  AND U29700 ( .A(n13250), .B(n13249), .Z(n52187) );
  AND U29701 ( .A(n13251), .B(n52187), .Z(n13254) );
  NANDN U29702 ( .A(x[1903]), .B(y[1903]), .Z(n13253) );
  NANDN U29703 ( .A(x[1904]), .B(y[1904]), .Z(n13252) );
  NAND U29704 ( .A(n13253), .B(n13252), .Z(n54037) );
  OR U29705 ( .A(n13254), .B(n54037), .Z(n13255) );
  NAND U29706 ( .A(n54038), .B(n13255), .Z(n13256) );
  NANDN U29707 ( .A(n54039), .B(n13256), .Z(n13257) );
  NANDN U29708 ( .A(y[1906]), .B(x[1906]), .Z(n54040) );
  AND U29709 ( .A(n13257), .B(n54040), .Z(n13258) );
  NAND U29710 ( .A(n27454), .B(n13258), .Z(n13259) );
  NANDN U29711 ( .A(n52186), .B(n13259), .Z(n13260) );
  ANDN U29712 ( .B(y[1908]), .A(x[1908]), .Z(n27451) );
  OR U29713 ( .A(n13260), .B(n27451), .Z(n13261) );
  NANDN U29714 ( .A(y[1909]), .B(x[1909]), .Z(n52185) );
  AND U29715 ( .A(n13261), .B(n52185), .Z(n13262) );
  NANDN U29716 ( .A(n27453), .B(n13262), .Z(n13263) );
  AND U29717 ( .A(n13264), .B(n13263), .Z(n13265) );
  OR U29718 ( .A(n54045), .B(n13265), .Z(n13266) );
  NAND U29719 ( .A(n54046), .B(n13266), .Z(n13267) );
  NANDN U29720 ( .A(n54047), .B(n13267), .Z(n13268) );
  NANDN U29721 ( .A(n52184), .B(n13268), .Z(n13269) );
  AND U29722 ( .A(n54048), .B(n13269), .Z(n13270) );
  OR U29723 ( .A(n54049), .B(n13270), .Z(n13271) );
  NAND U29724 ( .A(n54050), .B(n13271), .Z(n13272) );
  NANDN U29725 ( .A(n54051), .B(n13272), .Z(n13273) );
  ANDN U29726 ( .B(x[1918]), .A(y[1918]), .Z(n54052) );
  ANDN U29727 ( .B(n13273), .A(n54052), .Z(n13274) );
  NAND U29728 ( .A(n34302), .B(n13274), .Z(n13275) );
  NAND U29729 ( .A(n54053), .B(n13275), .Z(n13278) );
  ANDN U29730 ( .B(x[1920]), .A(y[1920]), .Z(n34303) );
  NANDN U29731 ( .A(n13276), .B(n34303), .Z(n13277) );
  AND U29732 ( .A(n13278), .B(n13277), .Z(n13279) );
  NANDN U29733 ( .A(n34301), .B(n13279), .Z(n13280) );
  AND U29734 ( .A(n54056), .B(n13280), .Z(n13281) );
  ANDN U29735 ( .B(x[1923]), .A(y[1923]), .Z(n52182) );
  OR U29736 ( .A(n13281), .B(n52182), .Z(n13282) );
  NANDN U29737 ( .A(x[1923]), .B(y[1923]), .Z(n27447) );
  NANDN U29738 ( .A(x[1924]), .B(y[1924]), .Z(n27446) );
  AND U29739 ( .A(n27447), .B(n27446), .Z(n54057) );
  AND U29740 ( .A(n13282), .B(n54057), .Z(n13283) );
  ANDN U29741 ( .B(x[1924]), .A(y[1924]), .Z(n34310) );
  ANDN U29742 ( .B(x[1925]), .A(y[1925]), .Z(n34316) );
  OR U29743 ( .A(n34310), .B(n34316), .Z(n52181) );
  OR U29744 ( .A(n13283), .B(n52181), .Z(n13284) );
  NAND U29745 ( .A(n52180), .B(n13284), .Z(n13285) );
  NANDN U29746 ( .A(n54059), .B(n13285), .Z(n13286) );
  AND U29747 ( .A(n54060), .B(n13286), .Z(n13288) );
  ANDN U29748 ( .B(x[1929]), .A(y[1929]), .Z(n27440) );
  NANDN U29749 ( .A(y[1928]), .B(x[1928]), .Z(n13287) );
  NANDN U29750 ( .A(n27440), .B(n13287), .Z(n27442) );
  OR U29751 ( .A(n13288), .B(n27442), .Z(n13289) );
  NAND U29752 ( .A(n54062), .B(n13289), .Z(n13290) );
  NANDN U29753 ( .A(n54063), .B(n13290), .Z(n13291) );
  NANDN U29754 ( .A(n54064), .B(n13291), .Z(n13292) );
  AND U29755 ( .A(n54065), .B(n13292), .Z(n13294) );
  NANDN U29756 ( .A(x[1934]), .B(y[1934]), .Z(n27435) );
  ANDN U29757 ( .B(y[1933]), .A(x[1933]), .Z(n54066) );
  ANDN U29758 ( .B(n27435), .A(n54066), .Z(n13293) );
  NANDN U29759 ( .A(n13294), .B(n13293), .Z(n13295) );
  NAND U29760 ( .A(n54067), .B(n13295), .Z(n13296) );
  ANDN U29761 ( .B(x[1935]), .A(y[1935]), .Z(n27432) );
  OR U29762 ( .A(n13296), .B(n27432), .Z(n13297) );
  AND U29763 ( .A(n27436), .B(n13297), .Z(n13298) );
  NANDN U29764 ( .A(x[1936]), .B(y[1936]), .Z(n34337) );
  AND U29765 ( .A(n13298), .B(n34337), .Z(n13299) );
  NANDN U29766 ( .A(y[1936]), .B(x[1936]), .Z(n27434) );
  NANDN U29767 ( .A(n13299), .B(n27434), .Z(n13300) );
  ANDN U29768 ( .B(x[1937]), .A(y[1937]), .Z(n27430) );
  OR U29769 ( .A(n13300), .B(n27430), .Z(n13301) );
  ANDN U29770 ( .B(y[1938]), .A(x[1938]), .Z(n54072) );
  ANDN U29771 ( .B(n13301), .A(n54072), .Z(n13302) );
  NANDN U29772 ( .A(n34336), .B(n13302), .Z(n13303) );
  AND U29773 ( .A(n13304), .B(n13303), .Z(n13305) );
  ANDN U29774 ( .B(y[1939]), .A(x[1939]), .Z(n34341) );
  NANDN U29775 ( .A(x[1940]), .B(y[1940]), .Z(n27428) );
  NANDN U29776 ( .A(n34341), .B(n27428), .Z(n54075) );
  OR U29777 ( .A(n13305), .B(n54075), .Z(n13306) );
  NAND U29778 ( .A(n54076), .B(n13306), .Z(n13307) );
  NANDN U29779 ( .A(n52179), .B(n13307), .Z(n13308) );
  NANDN U29780 ( .A(y[1942]), .B(x[1942]), .Z(n34348) );
  NANDN U29781 ( .A(y[1943]), .B(x[1943]), .Z(n27426) );
  AND U29782 ( .A(n34348), .B(n27426), .Z(n52178) );
  AND U29783 ( .A(n13308), .B(n52178), .Z(n13309) );
  OR U29784 ( .A(n54077), .B(n13309), .Z(n13310) );
  NAND U29785 ( .A(n54078), .B(n13310), .Z(n13311) );
  NANDN U29786 ( .A(n54079), .B(n13311), .Z(n13312) );
  NAND U29787 ( .A(n54080), .B(n13312), .Z(n13313) );
  NANDN U29788 ( .A(n54081), .B(n13313), .Z(n13314) );
  NANDN U29789 ( .A(y[1948]), .B(x[1948]), .Z(n27421) );
  NANDN U29790 ( .A(y[1949]), .B(x[1949]), .Z(n27420) );
  AND U29791 ( .A(n27421), .B(n27420), .Z(n52177) );
  AND U29792 ( .A(n13314), .B(n52177), .Z(n13315) );
  NANDN U29793 ( .A(x[1949]), .B(y[1949]), .Z(n34370) );
  NANDN U29794 ( .A(x[1950]), .B(y[1950]), .Z(n34377) );
  NAND U29795 ( .A(n34370), .B(n34377), .Z(n54082) );
  OR U29796 ( .A(n13315), .B(n54082), .Z(n13316) );
  NAND U29797 ( .A(n54083), .B(n13316), .Z(n13317) );
  NANDN U29798 ( .A(n52176), .B(n13317), .Z(n13318) );
  NANDN U29799 ( .A(n54086), .B(n13318), .Z(n13319) );
  NANDN U29800 ( .A(x[1953]), .B(y[1953]), .Z(n34382) );
  NANDN U29801 ( .A(x[1954]), .B(y[1954]), .Z(n27414) );
  AND U29802 ( .A(n34382), .B(n27414), .Z(n52175) );
  AND U29803 ( .A(n13319), .B(n52175), .Z(n13320) );
  NANDN U29804 ( .A(y[1954]), .B(x[1954]), .Z(n27415) );
  NANDN U29805 ( .A(y[1955]), .B(x[1955]), .Z(n27411) );
  NAND U29806 ( .A(n27415), .B(n27411), .Z(n54087) );
  OR U29807 ( .A(n13320), .B(n54087), .Z(n13321) );
  NAND U29808 ( .A(n54088), .B(n13321), .Z(n13322) );
  NANDN U29809 ( .A(n52174), .B(n13322), .Z(n13323) );
  NANDN U29810 ( .A(n54089), .B(n13323), .Z(n13324) );
  AND U29811 ( .A(n54090), .B(n13324), .Z(n13325) );
  NANDN U29812 ( .A(x[1959]), .B(y[1959]), .Z(n27409) );
  NANDN U29813 ( .A(x[1960]), .B(y[1960]), .Z(n34408) );
  NAND U29814 ( .A(n27409), .B(n34408), .Z(n54091) );
  OR U29815 ( .A(n13325), .B(n54091), .Z(n13326) );
  NAND U29816 ( .A(n54092), .B(n13326), .Z(n13327) );
  NANDN U29817 ( .A(n52173), .B(n13327), .Z(n13328) );
  NANDN U29818 ( .A(n54093), .B(n13328), .Z(n13329) );
  NANDN U29819 ( .A(x[1963]), .B(y[1963]), .Z(n34414) );
  NANDN U29820 ( .A(x[1964]), .B(y[1964]), .Z(n27408) );
  AND U29821 ( .A(n34414), .B(n27408), .Z(n52172) );
  AND U29822 ( .A(n13329), .B(n52172), .Z(n13330) );
  ANDN U29823 ( .B(x[1964]), .A(y[1964]), .Z(n34415) );
  ANDN U29824 ( .B(x[1965]), .A(y[1965]), .Z(n34417) );
  OR U29825 ( .A(n34415), .B(n34417), .Z(n54094) );
  OR U29826 ( .A(n13330), .B(n54094), .Z(n13331) );
  NAND U29827 ( .A(n54097), .B(n13331), .Z(n13332) );
  NANDN U29828 ( .A(n54099), .B(n13332), .Z(n13333) );
  NANDN U29829 ( .A(y[1967]), .B(x[1967]), .Z(n27406) );
  NANDN U29830 ( .A(n13333), .B(n27406), .Z(n13334) );
  NAND U29831 ( .A(n54100), .B(n13334), .Z(n13335) );
  NANDN U29832 ( .A(n52171), .B(n13335), .Z(n13336) );
  ANDN U29833 ( .B(x[1968]), .A(y[1968]), .Z(n27405) );
  OR U29834 ( .A(n13336), .B(n27405), .Z(n13337) );
  AND U29835 ( .A(n54101), .B(n13337), .Z(n13339) );
  NANDN U29836 ( .A(y[1970]), .B(x[1970]), .Z(n13338) );
  NANDN U29837 ( .A(y[1971]), .B(x[1971]), .Z(n27400) );
  NAND U29838 ( .A(n13338), .B(n27400), .Z(n52168) );
  OR U29839 ( .A(n13339), .B(n52168), .Z(n13340) );
  XNOR U29840 ( .A(y[1972]), .B(x[1972]), .Z(n27401) );
  NANDN U29841 ( .A(x[1971]), .B(y[1971]), .Z(n27402) );
  AND U29842 ( .A(n27401), .B(n27402), .Z(n52167) );
  AND U29843 ( .A(n13340), .B(n52167), .Z(n13342) );
  NANDN U29844 ( .A(y[1972]), .B(x[1972]), .Z(n13341) );
  NANDN U29845 ( .A(y[1973]), .B(x[1973]), .Z(n27398) );
  NAND U29846 ( .A(n13341), .B(n27398), .Z(n52166) );
  OR U29847 ( .A(n13342), .B(n52166), .Z(n13343) );
  NANDN U29848 ( .A(x[1973]), .B(y[1973]), .Z(n54102) );
  AND U29849 ( .A(n13343), .B(n54102), .Z(n13344) );
  ANDN U29850 ( .B(x[1974]), .A(y[1974]), .Z(n27397) );
  OR U29851 ( .A(n13344), .B(n27397), .Z(n13345) );
  NANDN U29852 ( .A(x[1975]), .B(y[1975]), .Z(n54105) );
  NANDN U29853 ( .A(x[1974]), .B(y[1974]), .Z(n52165) );
  AND U29854 ( .A(n54105), .B(n52165), .Z(n34430) );
  AND U29855 ( .A(n13345), .B(n34430), .Z(n13346) );
  NANDN U29856 ( .A(y[1975]), .B(x[1975]), .Z(n27396) );
  NANDN U29857 ( .A(n13346), .B(n27396), .Z(n13349) );
  NANDN U29858 ( .A(x[1976]), .B(y[1976]), .Z(n13347) );
  NANDN U29859 ( .A(n13348), .B(n13347), .Z(n34433) );
  IV U29860 ( .A(n34433), .Z(n54107) );
  AND U29861 ( .A(n13349), .B(n54107), .Z(n13350) );
  ANDN U29862 ( .B(n13351), .A(n13350), .Z(n13352) );
  OR U29863 ( .A(n54109), .B(n13352), .Z(n13353) );
  NANDN U29864 ( .A(y[1978]), .B(x[1978]), .Z(n27395) );
  NANDN U29865 ( .A(y[1979]), .B(x[1979]), .Z(n27393) );
  AND U29866 ( .A(n27395), .B(n27393), .Z(n52164) );
  AND U29867 ( .A(n13353), .B(n52164), .Z(n13354) );
  ANDN U29868 ( .B(y[1979]), .A(x[1979]), .Z(n34438) );
  NANDN U29869 ( .A(x[1980]), .B(y[1980]), .Z(n34443) );
  NANDN U29870 ( .A(n34438), .B(n34443), .Z(n54110) );
  OR U29871 ( .A(n13354), .B(n54110), .Z(n13355) );
  NAND U29872 ( .A(n54111), .B(n13355), .Z(n13356) );
  NANDN U29873 ( .A(n52163), .B(n13356), .Z(n13357) );
  NANDN U29874 ( .A(n54112), .B(n13357), .Z(n13358) );
  NANDN U29875 ( .A(x[1983]), .B(y[1983]), .Z(n27389) );
  NANDN U29876 ( .A(x[1984]), .B(y[1984]), .Z(n34452) );
  AND U29877 ( .A(n27389), .B(n34452), .Z(n52162) );
  AND U29878 ( .A(n13358), .B(n52162), .Z(n13359) );
  ANDN U29879 ( .B(x[1985]), .A(y[1985]), .Z(n34456) );
  NANDN U29880 ( .A(y[1984]), .B(x[1984]), .Z(n27388) );
  NANDN U29881 ( .A(n34456), .B(n27388), .Z(n54113) );
  OR U29882 ( .A(n13359), .B(n54113), .Z(n13360) );
  NANDN U29883 ( .A(x[1985]), .B(y[1985]), .Z(n54114) );
  AND U29884 ( .A(n13360), .B(n54114), .Z(n13361) );
  NANDN U29885 ( .A(x[1986]), .B(y[1986]), .Z(n27385) );
  NAND U29886 ( .A(n13361), .B(n27385), .Z(n13362) );
  NANDN U29887 ( .A(y[1987]), .B(x[1987]), .Z(n54119) );
  AND U29888 ( .A(n13362), .B(n54119), .Z(n13363) );
  NANDN U29889 ( .A(n54117), .B(n13363), .Z(n13364) );
  AND U29890 ( .A(n54120), .B(n13364), .Z(n13365) );
  NANDN U29891 ( .A(x[1987]), .B(y[1987]), .Z(n27386) );
  AND U29892 ( .A(n13365), .B(n27386), .Z(n13366) );
  NANDN U29893 ( .A(y[1988]), .B(x[1988]), .Z(n27384) );
  ANDN U29894 ( .B(x[1989]), .A(y[1989]), .Z(n34466) );
  ANDN U29895 ( .B(n27384), .A(n34466), .Z(n54121) );
  NANDN U29896 ( .A(n13366), .B(n54121), .Z(n13367) );
  NANDN U29897 ( .A(n52161), .B(n13367), .Z(n13368) );
  AND U29898 ( .A(n54122), .B(n13368), .Z(n13369) );
  OR U29899 ( .A(n54123), .B(n13369), .Z(n13370) );
  NAND U29900 ( .A(n54124), .B(n13370), .Z(n13371) );
  NANDN U29901 ( .A(n54125), .B(n13371), .Z(n13372) );
  NANDN U29902 ( .A(n52160), .B(n13372), .Z(n13373) );
  NANDN U29903 ( .A(x[1995]), .B(y[1995]), .Z(n27376) );
  NANDN U29904 ( .A(x[1996]), .B(y[1996]), .Z(n27373) );
  AND U29905 ( .A(n27376), .B(n27373), .Z(n52159) );
  AND U29906 ( .A(n13373), .B(n52159), .Z(n13374) );
  OR U29907 ( .A(n54126), .B(n13374), .Z(n13375) );
  NAND U29908 ( .A(n54127), .B(n13375), .Z(n13376) );
  NANDN U29909 ( .A(n54128), .B(n13376), .Z(n13377) );
  NANDN U29910 ( .A(n52158), .B(n13377), .Z(n13378) );
  AND U29911 ( .A(n54131), .B(n13378), .Z(n13379) );
  ANDN U29912 ( .B(y[2002]), .A(x[2002]), .Z(n34502) );
  NANDN U29913 ( .A(x[2001]), .B(y[2001]), .Z(n27368) );
  NANDN U29914 ( .A(n34502), .B(n27368), .Z(n54132) );
  OR U29915 ( .A(n13379), .B(n54132), .Z(n13380) );
  NAND U29916 ( .A(n13381), .B(n13380), .Z(n13382) );
  NANDN U29917 ( .A(n52157), .B(n13382), .Z(n13383) );
  NANDN U29918 ( .A(y[2005]), .B(x[2005]), .Z(n52156) );
  AND U29919 ( .A(n13383), .B(n52156), .Z(n13384) );
  NANDN U29920 ( .A(y[2004]), .B(x[2004]), .Z(n27365) );
  NAND U29921 ( .A(n13384), .B(n27365), .Z(n13385) );
  NANDN U29922 ( .A(n54136), .B(n13385), .Z(n13386) );
  AND U29923 ( .A(n54137), .B(n13386), .Z(n13387) );
  ANDN U29924 ( .B(y[2007]), .A(x[2007]), .Z(n34510) );
  ANDN U29925 ( .B(y[2008]), .A(x[2008]), .Z(n34516) );
  OR U29926 ( .A(n34510), .B(n34516), .Z(n54138) );
  OR U29927 ( .A(n13387), .B(n54138), .Z(n13388) );
  AND U29928 ( .A(n54139), .B(n13388), .Z(n13389) );
  NANDN U29929 ( .A(y[2009]), .B(x[2009]), .Z(n27362) );
  AND U29930 ( .A(n13389), .B(n27362), .Z(n13390) );
  NANDN U29931 ( .A(x[2009]), .B(y[2009]), .Z(n27363) );
  NANDN U29932 ( .A(n13390), .B(n27363), .Z(n13391) );
  XOR U29933 ( .A(x[2010]), .B(y[2010]), .Z(n27361) );
  OR U29934 ( .A(n13391), .B(n27361), .Z(n13392) );
  AND U29935 ( .A(n54143), .B(n13392), .Z(n13393) );
  NANDN U29936 ( .A(n13394), .B(n13393), .Z(n13395) );
  AND U29937 ( .A(n13396), .B(n13395), .Z(n13397) );
  NANDN U29938 ( .A(y[2012]), .B(x[2012]), .Z(n34524) );
  NANDN U29939 ( .A(y[2013]), .B(x[2013]), .Z(n34529) );
  NAND U29940 ( .A(n34524), .B(n34529), .Z(n54146) );
  OR U29941 ( .A(n13397), .B(n54146), .Z(n13398) );
  NAND U29942 ( .A(n54147), .B(n13398), .Z(n13399) );
  NANDN U29943 ( .A(n52155), .B(n13399), .Z(n13400) );
  NANDN U29944 ( .A(n54148), .B(n13400), .Z(n13401) );
  AND U29945 ( .A(n54149), .B(n13401), .Z(n13403) );
  ANDN U29946 ( .B(y[2018]), .A(x[2018]), .Z(n27353) );
  ANDN U29947 ( .B(y[2017]), .A(x[2017]), .Z(n54150) );
  NOR U29948 ( .A(n27353), .B(n54150), .Z(n13402) );
  NANDN U29949 ( .A(n13403), .B(n13402), .Z(n13404) );
  NANDN U29950 ( .A(n27356), .B(n13404), .Z(n13405) );
  ANDN U29951 ( .B(x[2019]), .A(y[2019]), .Z(n27350) );
  OR U29952 ( .A(n13405), .B(n27350), .Z(n13406) );
  AND U29953 ( .A(n27354), .B(n13406), .Z(n13407) );
  NANDN U29954 ( .A(x[2020]), .B(y[2020]), .Z(n27349) );
  AND U29955 ( .A(n13407), .B(n27349), .Z(n13408) );
  NANDN U29956 ( .A(y[2020]), .B(x[2020]), .Z(n27352) );
  NANDN U29957 ( .A(n13408), .B(n27352), .Z(n13409) );
  ANDN U29958 ( .B(x[2021]), .A(y[2021]), .Z(n27346) );
  OR U29959 ( .A(n13409), .B(n27346), .Z(n13410) );
  NANDN U29960 ( .A(x[2022]), .B(y[2022]), .Z(n34548) );
  AND U29961 ( .A(n13410), .B(n34548), .Z(n13411) );
  NANDN U29962 ( .A(n27348), .B(n13411), .Z(n13412) );
  AND U29963 ( .A(n13413), .B(n13412), .Z(n13414) );
  OR U29964 ( .A(n54158), .B(n13414), .Z(n13415) );
  NAND U29965 ( .A(n54159), .B(n13415), .Z(n13416) );
  NANDN U29966 ( .A(n54160), .B(n13416), .Z(n13417) );
  NANDN U29967 ( .A(y[2027]), .B(x[2027]), .Z(n27344) );
  AND U29968 ( .A(n13417), .B(n27344), .Z(n13418) );
  NAND U29969 ( .A(n54161), .B(n13418), .Z(n13419) );
  NANDN U29970 ( .A(n54163), .B(n13419), .Z(n13420) );
  AND U29971 ( .A(n54164), .B(n13420), .Z(n13421) );
  NANDN U29972 ( .A(y[2028]), .B(x[2028]), .Z(n27343) );
  NAND U29973 ( .A(n13421), .B(n27343), .Z(n13422) );
  NANDN U29974 ( .A(n54167), .B(n13422), .Z(n13423) );
  AND U29975 ( .A(n54168), .B(n13423), .Z(n13424) );
  OR U29976 ( .A(n54169), .B(n13424), .Z(n13425) );
  NAND U29977 ( .A(n52154), .B(n13425), .Z(n13426) );
  NANDN U29978 ( .A(n54170), .B(n13426), .Z(n13427) );
  NANDN U29979 ( .A(n54171), .B(n13427), .Z(n13428) );
  AND U29980 ( .A(n54172), .B(n13428), .Z(n13429) );
  OR U29981 ( .A(n54173), .B(n13429), .Z(n13430) );
  NAND U29982 ( .A(n52153), .B(n13430), .Z(n13431) );
  NANDN U29983 ( .A(n54174), .B(n13431), .Z(n13432) );
  AND U29984 ( .A(n54175), .B(n13432), .Z(n13433) );
  OR U29985 ( .A(n54176), .B(n13433), .Z(n13434) );
  NAND U29986 ( .A(n54178), .B(n13434), .Z(n13435) );
  NANDN U29987 ( .A(n54179), .B(n13435), .Z(n13436) );
  NAND U29988 ( .A(n54180), .B(n13436), .Z(n13437) );
  NANDN U29989 ( .A(n54181), .B(n13437), .Z(n13438) );
  AND U29990 ( .A(n54182), .B(n13438), .Z(n13439) );
  OR U29991 ( .A(n54183), .B(n13439), .Z(n13440) );
  NAND U29992 ( .A(n54184), .B(n13440), .Z(n13441) );
  NANDN U29993 ( .A(n54185), .B(n13441), .Z(n13442) );
  NANDN U29994 ( .A(n54186), .B(n13442), .Z(n13443) );
  AND U29995 ( .A(n27324), .B(n13443), .Z(n13444) );
  NANDN U29996 ( .A(n54187), .B(n13444), .Z(n13445) );
  NANDN U29997 ( .A(x[2052]), .B(y[2052]), .Z(n54190) );
  AND U29998 ( .A(n13445), .B(n54190), .Z(n13446) );
  NAND U29999 ( .A(n54188), .B(n13446), .Z(n13447) );
  ANDN U30000 ( .B(x[2053]), .A(y[2053]), .Z(n54191) );
  ANDN U30001 ( .B(n13447), .A(n54191), .Z(n13448) );
  NANDN U30002 ( .A(y[2052]), .B(x[2052]), .Z(n27325) );
  NAND U30003 ( .A(n13448), .B(n27325), .Z(n13449) );
  NANDN U30004 ( .A(n54192), .B(n13449), .Z(n13450) );
  AND U30005 ( .A(n54193), .B(n13450), .Z(n13451) );
  NANDN U30006 ( .A(x[2055]), .B(y[2055]), .Z(n27322) );
  NANDN U30007 ( .A(x[2056]), .B(y[2056]), .Z(n27321) );
  NAND U30008 ( .A(n27322), .B(n27321), .Z(n54194) );
  OR U30009 ( .A(n13451), .B(n54194), .Z(n13452) );
  ANDN U30010 ( .B(x[2056]), .A(y[2056]), .Z(n54195) );
  ANDN U30011 ( .B(n13452), .A(n54195), .Z(n13453) );
  NANDN U30012 ( .A(n34652), .B(n13453), .Z(n13456) );
  NANDN U30013 ( .A(x[2059]), .B(y[2059]), .Z(n13458) );
  NANDN U30014 ( .A(x[2058]), .B(y[2058]), .Z(n13454) );
  AND U30015 ( .A(n13458), .B(n13454), .Z(n34654) );
  NANDN U30016 ( .A(x[2057]), .B(y[2057]), .Z(n13455) );
  AND U30017 ( .A(n34654), .B(n13455), .Z(n54196) );
  AND U30018 ( .A(n13456), .B(n54196), .Z(n13460) );
  ANDN U30019 ( .B(x[2058]), .A(y[2058]), .Z(n34651) );
  ANDN U30020 ( .B(x[2059]), .A(y[2059]), .Z(n34656) );
  OR U30021 ( .A(n34651), .B(n34656), .Z(n13457) );
  AND U30022 ( .A(n13458), .B(n13457), .Z(n13459) );
  OR U30023 ( .A(n13460), .B(n13459), .Z(n13461) );
  AND U30024 ( .A(n54200), .B(n13461), .Z(n13462) );
  ANDN U30025 ( .B(n13463), .A(n13462), .Z(n13464) );
  ANDN U30026 ( .B(y[2062]), .A(x[2062]), .Z(n27319) );
  OR U30027 ( .A(n13464), .B(n27319), .Z(n13465) );
  AND U30028 ( .A(n54203), .B(n13465), .Z(n13466) );
  ANDN U30029 ( .B(y[2064]), .A(x[2064]), .Z(n27317) );
  NANDN U30030 ( .A(x[2063]), .B(y[2063]), .Z(n27320) );
  NANDN U30031 ( .A(n27317), .B(n27320), .Z(n52152) );
  OR U30032 ( .A(n13466), .B(n52152), .Z(n13467) );
  NAND U30033 ( .A(n54204), .B(n13467), .Z(n13468) );
  NANDN U30034 ( .A(n54205), .B(n13468), .Z(n13469) );
  NANDN U30035 ( .A(n54206), .B(n13469), .Z(n13470) );
  AND U30036 ( .A(n54207), .B(n13470), .Z(n13472) );
  NANDN U30037 ( .A(y[2068]), .B(x[2068]), .Z(n13471) );
  NANDN U30038 ( .A(y[2069]), .B(x[2069]), .Z(n27313) );
  NAND U30039 ( .A(n13471), .B(n27313), .Z(n52151) );
  OR U30040 ( .A(n13472), .B(n52151), .Z(n13473) );
  NAND U30041 ( .A(n54208), .B(n13473), .Z(n13474) );
  NANDN U30042 ( .A(n54209), .B(n13474), .Z(n13475) );
  NANDN U30043 ( .A(n54210), .B(n13475), .Z(n13476) );
  AND U30044 ( .A(n54211), .B(n13476), .Z(n13477) );
  OR U30045 ( .A(n54214), .B(n13477), .Z(n13478) );
  NAND U30046 ( .A(n54216), .B(n13478), .Z(n13479) );
  NANDN U30047 ( .A(n54217), .B(n13479), .Z(n13480) );
  NAND U30048 ( .A(n54220), .B(n13480), .Z(n13481) );
  NANDN U30049 ( .A(n52149), .B(n13481), .Z(n13482) );
  NANDN U30050 ( .A(n27303), .B(n13482), .Z(n13483) );
  NANDN U30051 ( .A(n34711), .B(n13483), .Z(n13484) );
  NAND U30052 ( .A(n54227), .B(n13484), .Z(n13485) );
  AND U30053 ( .A(n54230), .B(n13485), .Z(n13486) );
  NANDN U30054 ( .A(y[2082]), .B(x[2082]), .Z(n34715) );
  NANDN U30055 ( .A(y[2083]), .B(x[2083]), .Z(n34721) );
  NAND U30056 ( .A(n34715), .B(n34721), .Z(n54232) );
  OR U30057 ( .A(n13486), .B(n54232), .Z(n13487) );
  NANDN U30058 ( .A(x[2084]), .B(y[2084]), .Z(n27299) );
  AND U30059 ( .A(n13487), .B(n27299), .Z(n13488) );
  NANDN U30060 ( .A(n54233), .B(n13488), .Z(n13489) );
  NANDN U30061 ( .A(n34720), .B(n13489), .Z(n13493) );
  ANDN U30062 ( .B(y[2086]), .A(x[2086]), .Z(n27302) );
  ANDN U30063 ( .B(y[2085]), .A(x[2085]), .Z(n27300) );
  OR U30064 ( .A(n27302), .B(n27300), .Z(n13490) );
  AND U30065 ( .A(n13491), .B(n13490), .Z(n13492) );
  ANDN U30066 ( .B(n13493), .A(n13492), .Z(n13494) );
  ANDN U30067 ( .B(x[2087]), .A(y[2087]), .Z(n27298) );
  OR U30068 ( .A(n13494), .B(n27298), .Z(n13495) );
  NAND U30069 ( .A(n54241), .B(n13495), .Z(n13496) );
  AND U30070 ( .A(n54244), .B(n13496), .Z(n13497) );
  NANDN U30071 ( .A(y[2089]), .B(x[2089]), .Z(n27296) );
  NAND U30072 ( .A(n13497), .B(n27296), .Z(n13498) );
  NANDN U30073 ( .A(x[2090]), .B(y[2090]), .Z(n27294) );
  AND U30074 ( .A(n13498), .B(n27294), .Z(n13499) );
  NAND U30075 ( .A(n54245), .B(n13499), .Z(n13500) );
  NANDN U30076 ( .A(y[2090]), .B(x[2090]), .Z(n27295) );
  AND U30077 ( .A(n13500), .B(n27295), .Z(n13501) );
  NAND U30078 ( .A(n27292), .B(n13501), .Z(n13502) );
  NANDN U30079 ( .A(n34734), .B(n13502), .Z(n13503) );
  ANDN U30080 ( .B(y[2091]), .A(x[2091]), .Z(n27293) );
  OR U30081 ( .A(n13503), .B(n27293), .Z(n13504) );
  AND U30082 ( .A(n54253), .B(n13504), .Z(n13505) );
  NANDN U30083 ( .A(n13506), .B(n13505), .Z(n13507) );
  AND U30084 ( .A(n13508), .B(n13507), .Z(n13509) );
  NANDN U30085 ( .A(y[2094]), .B(x[2094]), .Z(n34738) );
  NANDN U30086 ( .A(y[2095]), .B(x[2095]), .Z(n34743) );
  NAND U30087 ( .A(n34738), .B(n34743), .Z(n54255) );
  OR U30088 ( .A(n13509), .B(n54255), .Z(n13510) );
  NAND U30089 ( .A(n54256), .B(n13510), .Z(n13511) );
  NANDN U30090 ( .A(n52148), .B(n13511), .Z(n13512) );
  AND U30091 ( .A(n54257), .B(n13512), .Z(n13513) );
  OR U30092 ( .A(n54258), .B(n13513), .Z(n13514) );
  NAND U30093 ( .A(n54259), .B(n13514), .Z(n13515) );
  NANDN U30094 ( .A(n54260), .B(n13515), .Z(n13516) );
  NAND U30095 ( .A(n54261), .B(n13516), .Z(n13517) );
  NANDN U30096 ( .A(n54262), .B(n13517), .Z(n13518) );
  AND U30097 ( .A(n54263), .B(n13518), .Z(n13519) );
  NANDN U30098 ( .A(y[2104]), .B(x[2104]), .Z(n27286) );
  NANDN U30099 ( .A(y[2105]), .B(x[2105]), .Z(n34781) );
  NAND U30100 ( .A(n27286), .B(n34781), .Z(n54264) );
  OR U30101 ( .A(n13519), .B(n54264), .Z(n13520) );
  NAND U30102 ( .A(n54265), .B(n13520), .Z(n13521) );
  NANDN U30103 ( .A(n52147), .B(n13521), .Z(n13522) );
  AND U30104 ( .A(n54267), .B(n13522), .Z(n13524) );
  NANDN U30105 ( .A(y[2108]), .B(x[2108]), .Z(n34788) );
  NANDN U30106 ( .A(y[2109]), .B(x[2109]), .Z(n13523) );
  NAND U30107 ( .A(n34788), .B(n13523), .Z(n52146) );
  OR U30108 ( .A(n13524), .B(n52146), .Z(n13525) );
  NAND U30109 ( .A(n54268), .B(n13525), .Z(n13526) );
  NANDN U30110 ( .A(n34799), .B(n13526), .Z(n13529) );
  NANDN U30111 ( .A(x[2112]), .B(y[2112]), .Z(n13528) );
  NANDN U30112 ( .A(x[2111]), .B(y[2111]), .Z(n13527) );
  AND U30113 ( .A(n13528), .B(n13527), .Z(n34801) );
  AND U30114 ( .A(n13529), .B(n34801), .Z(n13532) );
  NANDN U30115 ( .A(y[2112]), .B(x[2112]), .Z(n13531) );
  NANDN U30116 ( .A(y[2113]), .B(x[2113]), .Z(n13530) );
  NAND U30117 ( .A(n13531), .B(n13530), .Z(n27285) );
  OR U30118 ( .A(n13532), .B(n27285), .Z(n13533) );
  NAND U30119 ( .A(n27284), .B(n13533), .Z(n13534) );
  NANDN U30120 ( .A(n27283), .B(n13534), .Z(n13535) );
  NANDN U30121 ( .A(n54274), .B(n13535), .Z(n13536) );
  AND U30122 ( .A(n54275), .B(n13536), .Z(n13537) );
  OR U30123 ( .A(n54276), .B(n13537), .Z(n13538) );
  NAND U30124 ( .A(n54277), .B(n13538), .Z(n13539) );
  NANDN U30125 ( .A(n54278), .B(n13539), .Z(n13540) );
  NANDN U30126 ( .A(n54279), .B(n13540), .Z(n13541) );
  AND U30127 ( .A(n54280), .B(n13541), .Z(n13543) );
  NANDN U30128 ( .A(y[2122]), .B(x[2122]), .Z(n13542) );
  NANDN U30129 ( .A(y[2123]), .B(x[2123]), .Z(n27280) );
  NAND U30130 ( .A(n13542), .B(n27280), .Z(n54281) );
  OR U30131 ( .A(n13543), .B(n54281), .Z(n13544) );
  NAND U30132 ( .A(n54283), .B(n13544), .Z(n13545) );
  NANDN U30133 ( .A(n54284), .B(n13545), .Z(n13546) );
  NANDN U30134 ( .A(n54285), .B(n13546), .Z(n13547) );
  AND U30135 ( .A(n54286), .B(n13547), .Z(n13550) );
  NANDN U30136 ( .A(x[2127]), .B(y[2127]), .Z(n13549) );
  NANDN U30137 ( .A(x[2128]), .B(y[2128]), .Z(n13548) );
  AND U30138 ( .A(n13549), .B(n13548), .Z(n54287) );
  NANDN U30139 ( .A(n13550), .B(n54287), .Z(n13551) );
  AND U30140 ( .A(n54288), .B(n13551), .Z(n13552) );
  OR U30141 ( .A(n54289), .B(n13552), .Z(n13553) );
  NAND U30142 ( .A(n54290), .B(n13553), .Z(n13554) );
  NANDN U30143 ( .A(n54291), .B(n13554), .Z(n13555) );
  NANDN U30144 ( .A(n54292), .B(n13555), .Z(n13556) );
  AND U30145 ( .A(n54293), .B(n13556), .Z(n13557) );
  OR U30146 ( .A(n54294), .B(n13557), .Z(n13558) );
  NAND U30147 ( .A(n54295), .B(n13558), .Z(n13559) );
  NANDN U30148 ( .A(n54296), .B(n13559), .Z(n13560) );
  NANDN U30149 ( .A(n54297), .B(n13560), .Z(n13561) );
  AND U30150 ( .A(n54298), .B(n13561), .Z(n13562) );
  OR U30151 ( .A(n54299), .B(n13562), .Z(n13563) );
  NAND U30152 ( .A(n54300), .B(n13563), .Z(n13564) );
  NANDN U30153 ( .A(n54301), .B(n13564), .Z(n13565) );
  NANDN U30154 ( .A(n54302), .B(n13565), .Z(n13567) );
  NANDN U30155 ( .A(x[2143]), .B(y[2143]), .Z(n34896) );
  XNOR U30156 ( .A(y[2144]), .B(x[2144]), .Z(n13566) );
  AND U30157 ( .A(n34896), .B(n13566), .Z(n54305) );
  AND U30158 ( .A(n13567), .B(n54305), .Z(n13568) );
  ANDN U30159 ( .B(x[2145]), .A(y[2145]), .Z(n34907) );
  NANDN U30160 ( .A(y[2144]), .B(x[2144]), .Z(n27269) );
  NANDN U30161 ( .A(n34907), .B(n27269), .Z(n52145) );
  OR U30162 ( .A(n13568), .B(n52145), .Z(n13569) );
  NAND U30163 ( .A(n52144), .B(n13569), .Z(n13570) );
  NANDN U30164 ( .A(n54306), .B(n13570), .Z(n13571) );
  ANDN U30165 ( .B(x[2147]), .A(y[2147]), .Z(n27265) );
  OR U30166 ( .A(n13571), .B(n27265), .Z(n13572) );
  NANDN U30167 ( .A(n13573), .B(n13572), .Z(n13574) );
  AND U30168 ( .A(n13575), .B(n13574), .Z(n13576) );
  ANDN U30169 ( .B(y[2149]), .A(x[2149]), .Z(n27264) );
  OR U30170 ( .A(n13576), .B(n27264), .Z(n13577) );
  AND U30171 ( .A(n34914), .B(n13577), .Z(n13580) );
  NANDN U30172 ( .A(x[2150]), .B(y[2150]), .Z(n13578) );
  AND U30173 ( .A(n13579), .B(n13578), .Z(n54311) );
  NANDN U30174 ( .A(n13580), .B(n54311), .Z(n13581) );
  NANDN U30175 ( .A(n13582), .B(n13581), .Z(n13583) );
  ANDN U30176 ( .B(y[2152]), .A(x[2152]), .Z(n54313) );
  ANDN U30177 ( .B(n13583), .A(n54313), .Z(n13584) );
  OR U30178 ( .A(n54314), .B(n13584), .Z(n13585) );
  NAND U30179 ( .A(n54315), .B(n13585), .Z(n13586) );
  NANDN U30180 ( .A(n54316), .B(n13586), .Z(n13587) );
  NANDN U30181 ( .A(n54318), .B(n13587), .Z(n13588) );
  AND U30182 ( .A(n54319), .B(n13588), .Z(n13589) );
  OR U30183 ( .A(n54320), .B(n13589), .Z(n13590) );
  NAND U30184 ( .A(n54321), .B(n13590), .Z(n13591) );
  NAND U30185 ( .A(n54322), .B(n13591), .Z(n13594) );
  NANDN U30186 ( .A(y[2160]), .B(x[2160]), .Z(n13593) );
  NANDN U30187 ( .A(y[2159]), .B(x[2159]), .Z(n13592) );
  NAND U30188 ( .A(n13593), .B(n13592), .Z(n54323) );
  ANDN U30189 ( .B(n13594), .A(n54323), .Z(n13597) );
  NANDN U30190 ( .A(x[2160]), .B(y[2160]), .Z(n13596) );
  NANDN U30191 ( .A(x[2161]), .B(y[2161]), .Z(n13595) );
  AND U30192 ( .A(n13596), .B(n13595), .Z(n54324) );
  NANDN U30193 ( .A(n13597), .B(n54324), .Z(n13598) );
  NANDN U30194 ( .A(n54325), .B(n13598), .Z(n13599) );
  NANDN U30195 ( .A(n27263), .B(n13599), .Z(n13600) );
  NANDN U30196 ( .A(y[2163]), .B(x[2163]), .Z(n34948) );
  AND U30197 ( .A(n13600), .B(n34948), .Z(n13601) );
  ANDN U30198 ( .B(y[2164]), .A(x[2164]), .Z(n27261) );
  OR U30199 ( .A(n13601), .B(n27261), .Z(n13602) );
  NANDN U30200 ( .A(n54329), .B(n13602), .Z(n13603) );
  AND U30201 ( .A(n54330), .B(n13603), .Z(n13604) );
  OR U30202 ( .A(n54331), .B(n13604), .Z(n13605) );
  NAND U30203 ( .A(n54332), .B(n13605), .Z(n13606) );
  NANDN U30204 ( .A(n54333), .B(n13606), .Z(n13607) );
  NANDN U30205 ( .A(x[2170]), .B(y[2170]), .Z(n27258) );
  AND U30206 ( .A(n13607), .B(n27258), .Z(n13608) );
  NAND U30207 ( .A(n54334), .B(n13608), .Z(n13609) );
  NANDN U30208 ( .A(n54336), .B(n13609), .Z(n13610) );
  ANDN U30209 ( .B(y[2172]), .A(x[2172]), .Z(n54337) );
  ANDN U30210 ( .B(n13610), .A(n54337), .Z(n13611) );
  NANDN U30211 ( .A(x[2171]), .B(y[2171]), .Z(n27257) );
  NAND U30212 ( .A(n13611), .B(n27257), .Z(n13612) );
  NANDN U30213 ( .A(n54340), .B(n13612), .Z(n13613) );
  AND U30214 ( .A(n54341), .B(n13613), .Z(n13614) );
  OR U30215 ( .A(n54342), .B(n13614), .Z(n13615) );
  NAND U30216 ( .A(n54343), .B(n13615), .Z(n13616) );
  NANDN U30217 ( .A(n54344), .B(n13616), .Z(n13617) );
  NAND U30218 ( .A(n52143), .B(n13617), .Z(n13618) );
  NANDN U30219 ( .A(n54345), .B(n13618), .Z(n13619) );
  NAND U30220 ( .A(n34991), .B(n13619), .Z(n13620) );
  AND U30221 ( .A(n54346), .B(n13620), .Z(n13621) );
  ANDN U30222 ( .B(y[2180]), .A(x[2180]), .Z(n34994) );
  OR U30223 ( .A(n13621), .B(n34994), .Z(n13622) );
  NANDN U30224 ( .A(n54348), .B(n13622), .Z(n13623) );
  NANDN U30225 ( .A(x[2181]), .B(y[2181]), .Z(n34995) );
  NANDN U30226 ( .A(x[2182]), .B(y[2182]), .Z(n27251) );
  AND U30227 ( .A(n34995), .B(n27251), .Z(n54349) );
  AND U30228 ( .A(n13623), .B(n54349), .Z(n13624) );
  ANDN U30229 ( .B(x[2182]), .A(y[2182]), .Z(n34999) );
  ANDN U30230 ( .B(x[2183]), .A(y[2183]), .Z(n35007) );
  OR U30231 ( .A(n34999), .B(n35007), .Z(n52140) );
  OR U30232 ( .A(n13624), .B(n52140), .Z(n13625) );
  NAND U30233 ( .A(n52139), .B(n13625), .Z(n13626) );
  NANDN U30234 ( .A(n54352), .B(n13626), .Z(n13627) );
  NANDN U30235 ( .A(n54353), .B(n13627), .Z(n13628) );
  AND U30236 ( .A(n54354), .B(n13628), .Z(n13629) );
  XOR U30237 ( .A(y[2188]), .B(x[2188]), .Z(n35021) );
  NANDN U30238 ( .A(x[2187]), .B(y[2187]), .Z(n35017) );
  NANDN U30239 ( .A(n35021), .B(n35017), .Z(n52138) );
  OR U30240 ( .A(n13629), .B(n52138), .Z(n13630) );
  NAND U30241 ( .A(n52137), .B(n13630), .Z(n13631) );
  NANDN U30242 ( .A(n52136), .B(n13631), .Z(n13632) );
  NANDN U30243 ( .A(y[2190]), .B(x[2190]), .Z(n52135) );
  AND U30244 ( .A(n13632), .B(n52135), .Z(n13633) );
  NAND U30245 ( .A(n27248), .B(n13633), .Z(n13634) );
  NANDN U30246 ( .A(n35032), .B(n13634), .Z(n13635) );
  NAND U30247 ( .A(n27249), .B(n13635), .Z(n13636) );
  NAND U30248 ( .A(n54357), .B(n13636), .Z(n13637) );
  NANDN U30249 ( .A(n54358), .B(n13637), .Z(n13638) );
  AND U30250 ( .A(n54360), .B(n13638), .Z(n13639) );
  OR U30251 ( .A(n54361), .B(n13639), .Z(n13640) );
  NAND U30252 ( .A(n54362), .B(n13640), .Z(n13641) );
  NANDN U30253 ( .A(n54363), .B(n13641), .Z(n13642) );
  NAND U30254 ( .A(n52134), .B(n13642), .Z(n13643) );
  NANDN U30255 ( .A(n54364), .B(n13643), .Z(n13644) );
  NANDN U30256 ( .A(x[2200]), .B(y[2200]), .Z(n54365) );
  AND U30257 ( .A(n13644), .B(n54365), .Z(n13645) );
  ANDN U30258 ( .B(x[2200]), .A(y[2200]), .Z(n35046) );
  ANDN U30259 ( .B(x[2201]), .A(y[2201]), .Z(n35053) );
  OR U30260 ( .A(n35046), .B(n35053), .Z(n54366) );
  OR U30261 ( .A(n13645), .B(n54366), .Z(n13646) );
  NAND U30262 ( .A(n54367), .B(n13646), .Z(n13647) );
  NANDN U30263 ( .A(n52133), .B(n13647), .Z(n13648) );
  NANDN U30264 ( .A(n54368), .B(n13648), .Z(n13649) );
  NANDN U30265 ( .A(y[2204]), .B(x[2204]), .Z(n35059) );
  NANDN U30266 ( .A(y[2205]), .B(x[2205]), .Z(n35065) );
  AND U30267 ( .A(n35059), .B(n35065), .Z(n52132) );
  AND U30268 ( .A(n13649), .B(n52132), .Z(n13650) );
  NANDN U30269 ( .A(x[2205]), .B(y[2205]), .Z(n27247) );
  NANDN U30270 ( .A(x[2206]), .B(y[2206]), .Z(n27245) );
  NAND U30271 ( .A(n27247), .B(n27245), .Z(n54369) );
  OR U30272 ( .A(n13650), .B(n54369), .Z(n13651) );
  NAND U30273 ( .A(n54372), .B(n13651), .Z(n13652) );
  NANDN U30274 ( .A(n52131), .B(n13652), .Z(n13653) );
  NAND U30275 ( .A(n54374), .B(n13653), .Z(n13654) );
  ANDN U30276 ( .B(y[2210]), .A(x[2210]), .Z(n27240) );
  ANDN U30277 ( .B(n13654), .A(n27240), .Z(n13655) );
  NANDN U30278 ( .A(n52130), .B(n13655), .Z(n13656) );
  AND U30279 ( .A(n54375), .B(n13656), .Z(n13662) );
  NANDN U30280 ( .A(x[2212]), .B(y[2212]), .Z(n13658) );
  NANDN U30281 ( .A(x[2213]), .B(y[2213]), .Z(n13657) );
  AND U30282 ( .A(n13658), .B(n13657), .Z(n27243) );
  NANDN U30283 ( .A(x[2211]), .B(y[2211]), .Z(n27241) );
  OR U30284 ( .A(n27241), .B(n13659), .Z(n13660) );
  AND U30285 ( .A(n27243), .B(n13660), .Z(n13661) );
  NANDN U30286 ( .A(n13662), .B(n13661), .Z(n13663) );
  NANDN U30287 ( .A(n54376), .B(n13663), .Z(n13664) );
  NANDN U30288 ( .A(n35082), .B(n13664), .Z(n13665) );
  NAND U30289 ( .A(n35084), .B(n13665), .Z(n13666) );
  NANDN U30290 ( .A(n27239), .B(n13666), .Z(n13667) );
  NANDN U30291 ( .A(y[2217]), .B(x[2217]), .Z(n35089) );
  AND U30292 ( .A(n13667), .B(n35089), .Z(n13668) );
  ANDN U30293 ( .B(y[2218]), .A(x[2218]), .Z(n54381) );
  OR U30294 ( .A(n13668), .B(n54381), .Z(n13669) );
  AND U30295 ( .A(n54382), .B(n13669), .Z(n13672) );
  NANDN U30296 ( .A(x[2219]), .B(y[2219]), .Z(n13671) );
  NANDN U30297 ( .A(x[2220]), .B(y[2220]), .Z(n13670) );
  NAND U30298 ( .A(n13671), .B(n13670), .Z(n35094) );
  OR U30299 ( .A(n13672), .B(n35094), .Z(n13675) );
  NANDN U30300 ( .A(y[2221]), .B(x[2221]), .Z(n13674) );
  NANDN U30301 ( .A(y[2220]), .B(x[2220]), .Z(n13673) );
  AND U30302 ( .A(n13674), .B(n13673), .Z(n27238) );
  AND U30303 ( .A(n13675), .B(n27238), .Z(n13676) );
  NANDN U30304 ( .A(x[2221]), .B(y[2221]), .Z(n35098) );
  NANDN U30305 ( .A(x[2222]), .B(y[2222]), .Z(n27237) );
  NAND U30306 ( .A(n35098), .B(n27237), .Z(n52128) );
  OR U30307 ( .A(n13676), .B(n52128), .Z(n13677) );
  NAND U30308 ( .A(n54386), .B(n13677), .Z(n13678) );
  NANDN U30309 ( .A(n54387), .B(n13678), .Z(n13679) );
  NANDN U30310 ( .A(n54388), .B(n13679), .Z(n13680) );
  XNOR U30311 ( .A(y[2226]), .B(x[2226]), .Z(n27233) );
  NANDN U30312 ( .A(x[2225]), .B(y[2225]), .Z(n27235) );
  AND U30313 ( .A(n27233), .B(n27235), .Z(n54389) );
  AND U30314 ( .A(n13680), .B(n54389), .Z(n13682) );
  NANDN U30315 ( .A(y[2227]), .B(x[2227]), .Z(n35114) );
  NANDN U30316 ( .A(y[2226]), .B(x[2226]), .Z(n13681) );
  NAND U30317 ( .A(n35114), .B(n13681), .Z(n52127) );
  OR U30318 ( .A(n13682), .B(n52127), .Z(n13683) );
  NAND U30319 ( .A(n54390), .B(n13683), .Z(n13684) );
  NANDN U30320 ( .A(n27229), .B(n13684), .Z(n13685) );
  NAND U30321 ( .A(n27228), .B(n13685), .Z(n13686) );
  NANDN U30322 ( .A(n27227), .B(n13686), .Z(n13687) );
  NANDN U30323 ( .A(x[2231]), .B(y[2231]), .Z(n35121) );
  NANDN U30324 ( .A(x[2232]), .B(y[2232]), .Z(n35127) );
  AND U30325 ( .A(n35121), .B(n35127), .Z(n54394) );
  AND U30326 ( .A(n13687), .B(n54394), .Z(n13688) );
  ANDN U30327 ( .B(x[2232]), .A(y[2232]), .Z(n35123) );
  NANDN U30328 ( .A(y[2233]), .B(x[2233]), .Z(n27226) );
  NANDN U30329 ( .A(n35123), .B(n27226), .Z(n52126) );
  OR U30330 ( .A(n13688), .B(n52126), .Z(n13689) );
  NAND U30331 ( .A(n52125), .B(n13689), .Z(n13690) );
  NANDN U30332 ( .A(n54396), .B(n13690), .Z(n13691) );
  NANDN U30333 ( .A(n54397), .B(n13691), .Z(n13692) );
  AND U30334 ( .A(n54399), .B(n13692), .Z(n13693) );
  NANDN U30335 ( .A(x[2237]), .B(y[2237]), .Z(n35139) );
  NANDN U30336 ( .A(x[2238]), .B(y[2238]), .Z(n35147) );
  NAND U30337 ( .A(n35139), .B(n35147), .Z(n52124) );
  OR U30338 ( .A(n13693), .B(n52124), .Z(n13694) );
  AND U30339 ( .A(n54400), .B(n13694), .Z(n13695) );
  ANDN U30340 ( .B(y[2239]), .A(x[2239]), .Z(n35146) );
  OR U30341 ( .A(n13695), .B(n35146), .Z(n13696) );
  NANDN U30342 ( .A(y[2240]), .B(x[2240]), .Z(n27224) );
  AND U30343 ( .A(n13696), .B(n27224), .Z(n13697) );
  NANDN U30344 ( .A(x[2240]), .B(y[2240]), .Z(n54401) );
  NANDN U30345 ( .A(x[2241]), .B(y[2241]), .Z(n52122) );
  AND U30346 ( .A(n54401), .B(n52122), .Z(n35154) );
  NANDN U30347 ( .A(n13697), .B(n35154), .Z(n13698) );
  NAND U30348 ( .A(n35155), .B(n13698), .Z(n13699) );
  NANDN U30349 ( .A(n35158), .B(n13699), .Z(n13700) );
  NAND U30350 ( .A(n35160), .B(n13700), .Z(n13701) );
  NANDN U30351 ( .A(x[2244]), .B(y[2244]), .Z(n52120) );
  NANDN U30352 ( .A(x[2245]), .B(y[2245]), .Z(n54409) );
  AND U30353 ( .A(n52120), .B(n54409), .Z(n35161) );
  AND U30354 ( .A(n13701), .B(n35161), .Z(n13702) );
  ANDN U30355 ( .B(x[2245]), .A(y[2245]), .Z(n54406) );
  OR U30356 ( .A(n13702), .B(n54406), .Z(n13703) );
  NANDN U30357 ( .A(x[2246]), .B(y[2246]), .Z(n52118) );
  AND U30358 ( .A(n13703), .B(n52118), .Z(n13704) );
  NANDN U30359 ( .A(y[2246]), .B(x[2246]), .Z(n35164) );
  NANDN U30360 ( .A(y[2247]), .B(x[2247]), .Z(n27222) );
  NAND U30361 ( .A(n35164), .B(n27222), .Z(n54410) );
  OR U30362 ( .A(n13704), .B(n54410), .Z(n13705) );
  NANDN U30363 ( .A(x[2247]), .B(y[2247]), .Z(n27223) );
  NANDN U30364 ( .A(x[2248]), .B(y[2248]), .Z(n27219) );
  AND U30365 ( .A(n27223), .B(n27219), .Z(n54411) );
  AND U30366 ( .A(n13705), .B(n54411), .Z(n13706) );
  NANDN U30367 ( .A(y[2248]), .B(x[2248]), .Z(n27221) );
  NANDN U30368 ( .A(y[2249]), .B(x[2249]), .Z(n35173) );
  NAND U30369 ( .A(n27221), .B(n35173), .Z(n52117) );
  OR U30370 ( .A(n13706), .B(n52117), .Z(n13707) );
  NAND U30371 ( .A(n54412), .B(n13707), .Z(n13708) );
  NANDN U30372 ( .A(n35172), .B(n13708), .Z(n13709) );
  NANDN U30373 ( .A(y[2251]), .B(x[2251]), .Z(n27218) );
  NANDN U30374 ( .A(n13709), .B(n27218), .Z(n13710) );
  NANDN U30375 ( .A(x[2251]), .B(y[2251]), .Z(n35178) );
  AND U30376 ( .A(n13710), .B(n35178), .Z(n13711) );
  NANDN U30377 ( .A(x[2252]), .B(y[2252]), .Z(n35181) );
  NAND U30378 ( .A(n13711), .B(n35181), .Z(n13712) );
  NANDN U30379 ( .A(y[2253]), .B(x[2253]), .Z(n27216) );
  AND U30380 ( .A(n13712), .B(n27216), .Z(n13713) );
  NANDN U30381 ( .A(n27217), .B(n13713), .Z(n13714) );
  NANDN U30382 ( .A(x[2253]), .B(y[2253]), .Z(n35182) );
  AND U30383 ( .A(n13714), .B(n35182), .Z(n13715) );
  NAND U30384 ( .A(n27214), .B(n13715), .Z(n13716) );
  NANDN U30385 ( .A(n27211), .B(n13716), .Z(n13717) );
  ANDN U30386 ( .B(x[2254]), .A(y[2254]), .Z(n27215) );
  OR U30387 ( .A(n13717), .B(n27215), .Z(n13718) );
  AND U30388 ( .A(n13719), .B(n13718), .Z(n13720) );
  ANDN U30389 ( .B(x[2257]), .A(y[2257]), .Z(n35195) );
  NANDN U30390 ( .A(y[2256]), .B(x[2256]), .Z(n27212) );
  NANDN U30391 ( .A(n35195), .B(n27212), .Z(n54421) );
  OR U30392 ( .A(n13720), .B(n54421), .Z(n13721) );
  NAND U30393 ( .A(n54424), .B(n13721), .Z(n13722) );
  NANDN U30394 ( .A(n52116), .B(n13722), .Z(n13723) );
  NANDN U30395 ( .A(n54425), .B(n13723), .Z(n13724) );
  AND U30396 ( .A(n54426), .B(n13724), .Z(n13725) );
  XNOR U30397 ( .A(y[2262]), .B(x[2262]), .Z(n35208) );
  NANDN U30398 ( .A(x[2261]), .B(y[2261]), .Z(n27209) );
  NAND U30399 ( .A(n35208), .B(n27209), .Z(n54427) );
  OR U30400 ( .A(n13725), .B(n54427), .Z(n13726) );
  NAND U30401 ( .A(n54428), .B(n13726), .Z(n13727) );
  NANDN U30402 ( .A(n52115), .B(n13727), .Z(n13728) );
  NANDN U30403 ( .A(n54429), .B(n13728), .Z(n13729) );
  AND U30404 ( .A(n54430), .B(n13729), .Z(n13730) );
  ANDN U30405 ( .B(x[2267]), .A(y[2267]), .Z(n35231) );
  NANDN U30406 ( .A(y[2266]), .B(x[2266]), .Z(n27207) );
  NANDN U30407 ( .A(n35231), .B(n27207), .Z(n54431) );
  OR U30408 ( .A(n13730), .B(n54431), .Z(n13731) );
  NAND U30409 ( .A(n54432), .B(n13731), .Z(n13732) );
  NANDN U30410 ( .A(n35228), .B(n13732), .Z(n13733) );
  ANDN U30411 ( .B(x[2269]), .A(y[2269]), .Z(n27203) );
  OR U30412 ( .A(n13733), .B(n27203), .Z(n13734) );
  NAND U30413 ( .A(n13735), .B(n13734), .Z(n13737) );
  NANDN U30414 ( .A(y[2270]), .B(x[2270]), .Z(n13736) );
  AND U30415 ( .A(n13737), .B(n13736), .Z(n13738) );
  NAND U30416 ( .A(n27201), .B(n13738), .Z(n13739) );
  NANDN U30417 ( .A(n27202), .B(n13739), .Z(n13740) );
  ANDN U30418 ( .B(y[2272]), .A(x[2272]), .Z(n27197) );
  OR U30419 ( .A(n13740), .B(n27197), .Z(n13741) );
  AND U30420 ( .A(n54440), .B(n13741), .Z(n13742) );
  NANDN U30421 ( .A(n27200), .B(n13742), .Z(n13743) );
  AND U30422 ( .A(n13744), .B(n13743), .Z(n13745) );
  NANDN U30423 ( .A(y[2274]), .B(x[2274]), .Z(n35239) );
  NANDN U30424 ( .A(y[2275]), .B(x[2275]), .Z(n27195) );
  NAND U30425 ( .A(n35239), .B(n27195), .Z(n54442) );
  OR U30426 ( .A(n13745), .B(n54442), .Z(n13746) );
  NAND U30427 ( .A(n54443), .B(n13746), .Z(n13747) );
  NANDN U30428 ( .A(n52114), .B(n13747), .Z(n13748) );
  NANDN U30429 ( .A(x[2277]), .B(y[2277]), .Z(n27193) );
  NANDN U30430 ( .A(x[2278]), .B(y[2278]), .Z(n35252) );
  AND U30431 ( .A(n27193), .B(n35252), .Z(n52113) );
  AND U30432 ( .A(n13748), .B(n52113), .Z(n13749) );
  OR U30433 ( .A(n54444), .B(n13749), .Z(n13750) );
  NAND U30434 ( .A(n54445), .B(n13750), .Z(n13751) );
  NANDN U30435 ( .A(n54446), .B(n13751), .Z(n13752) );
  ANDN U30436 ( .B(x[2281]), .A(y[2281]), .Z(n27188) );
  OR U30437 ( .A(n13752), .B(n27188), .Z(n13753) );
  NAND U30438 ( .A(n13754), .B(n13753), .Z(n13755) );
  NANDN U30439 ( .A(n13756), .B(n13755), .Z(n13757) );
  ANDN U30440 ( .B(x[2283]), .A(y[2283]), .Z(n27185) );
  OR U30441 ( .A(n13757), .B(n27185), .Z(n13758) );
  NAND U30442 ( .A(n13759), .B(n13758), .Z(n13760) );
  NANDN U30443 ( .A(n13761), .B(n13760), .Z(n13762) );
  AND U30444 ( .A(n54452), .B(n13762), .Z(n13763) );
  NANDN U30445 ( .A(x[2285]), .B(y[2285]), .Z(n27183) );
  NAND U30446 ( .A(n13763), .B(n27183), .Z(n13764) );
  NANDN U30447 ( .A(n54453), .B(n13764), .Z(n13765) );
  AND U30448 ( .A(n54454), .B(n13765), .Z(n13766) );
  OR U30449 ( .A(n54455), .B(n13766), .Z(n13767) );
  NAND U30450 ( .A(n54456), .B(n13767), .Z(n13768) );
  NANDN U30451 ( .A(n54457), .B(n13768), .Z(n13769) );
  NANDN U30452 ( .A(x[2291]), .B(y[2291]), .Z(n27177) );
  AND U30453 ( .A(n13769), .B(n27177), .Z(n13770) );
  NAND U30454 ( .A(n27173), .B(n13770), .Z(n13771) );
  NANDN U30455 ( .A(n27171), .B(n13771), .Z(n13772) );
  ANDN U30456 ( .B(x[2292]), .A(y[2292]), .Z(n27175) );
  OR U30457 ( .A(n13772), .B(n27175), .Z(n13773) );
  AND U30458 ( .A(n13774), .B(n13773), .Z(n13775) );
  OR U30459 ( .A(n54463), .B(n13775), .Z(n13776) );
  NAND U30460 ( .A(n54464), .B(n13776), .Z(n13777) );
  NANDN U30461 ( .A(n54465), .B(n13777), .Z(n13778) );
  NANDN U30462 ( .A(n52110), .B(n13778), .Z(n13779) );
  AND U30463 ( .A(n54467), .B(n13779), .Z(n13781) );
  NANDN U30464 ( .A(x[2300]), .B(y[2300]), .Z(n27168) );
  NANDN U30465 ( .A(x[2299]), .B(y[2299]), .Z(n54468) );
  AND U30466 ( .A(n27168), .B(n54468), .Z(n13780) );
  NANDN U30467 ( .A(n13781), .B(n13780), .Z(n13782) );
  NANDN U30468 ( .A(n54471), .B(n13782), .Z(n13783) );
  NANDN U30469 ( .A(x[2301]), .B(y[2301]), .Z(n27167) );
  NANDN U30470 ( .A(x[2302]), .B(y[2302]), .Z(n27166) );
  AND U30471 ( .A(n27167), .B(n27166), .Z(n54472) );
  AND U30472 ( .A(n13783), .B(n54472), .Z(n13784) );
  ANDN U30473 ( .B(x[2303]), .A(y[2303]), .Z(n35317) );
  NANDN U30474 ( .A(y[2302]), .B(x[2302]), .Z(n35311) );
  NANDN U30475 ( .A(n35317), .B(n35311), .Z(n52109) );
  OR U30476 ( .A(n13784), .B(n52109), .Z(n13785) );
  NAND U30477 ( .A(n52108), .B(n13785), .Z(n13786) );
  NANDN U30478 ( .A(n52107), .B(n13786), .Z(n13787) );
  AND U30479 ( .A(n35325), .B(n13787), .Z(n13788) );
  NANDN U30480 ( .A(x[2305]), .B(y[2305]), .Z(n52106) );
  NAND U30481 ( .A(n13788), .B(n52106), .Z(n13789) );
  NANDN U30482 ( .A(n54473), .B(n13789), .Z(n13790) );
  AND U30483 ( .A(n54474), .B(n13790), .Z(n13791) );
  OR U30484 ( .A(n54475), .B(n13791), .Z(n13792) );
  NAND U30485 ( .A(n54476), .B(n13792), .Z(n13793) );
  NANDN U30486 ( .A(n54477), .B(n13793), .Z(n13794) );
  NAND U30487 ( .A(n54479), .B(n13794), .Z(n13795) );
  NANDN U30488 ( .A(y[2313]), .B(x[2313]), .Z(n27160) );
  AND U30489 ( .A(n13795), .B(n27160), .Z(n13796) );
  NANDN U30490 ( .A(n54480), .B(n13796), .Z(n13797) );
  AND U30491 ( .A(n54481), .B(n13797), .Z(n13799) );
  NANDN U30492 ( .A(y[2315]), .B(x[2315]), .Z(n27157) );
  ANDN U30493 ( .B(x[2314]), .A(y[2314]), .Z(n27159) );
  ANDN U30494 ( .B(n27157), .A(n27159), .Z(n13798) );
  NANDN U30495 ( .A(n13799), .B(n13798), .Z(n13800) );
  NANDN U30496 ( .A(n54487), .B(n13800), .Z(n13801) );
  NANDN U30497 ( .A(y[2316]), .B(x[2316]), .Z(n54486) );
  AND U30498 ( .A(n13801), .B(n54486), .Z(n13802) );
  NANDN U30499 ( .A(n27151), .B(n13802), .Z(n13803) );
  NAND U30500 ( .A(n54485), .B(n13803), .Z(n13804) );
  NANDN U30501 ( .A(n27156), .B(n13804), .Z(n13805) );
  ANDN U30502 ( .B(n13806), .A(n13805), .Z(n13809) );
  NANDN U30503 ( .A(x[2320]), .B(y[2320]), .Z(n13808) );
  NANDN U30504 ( .A(x[2321]), .B(y[2321]), .Z(n13807) );
  NAND U30505 ( .A(n13808), .B(n13807), .Z(n35358) );
  OR U30506 ( .A(n13809), .B(n35358), .Z(n13810) );
  NANDN U30507 ( .A(y[2321]), .B(x[2321]), .Z(n52104) );
  AND U30508 ( .A(n13810), .B(n52104), .Z(n13811) );
  ANDN U30509 ( .B(y[2322]), .A(x[2322]), .Z(n54490) );
  OR U30510 ( .A(n13811), .B(n54490), .Z(n13812) );
  AND U30511 ( .A(n54491), .B(n13812), .Z(n13813) );
  ANDN U30512 ( .B(y[2323]), .A(x[2323]), .Z(n35364) );
  NANDN U30513 ( .A(x[2324]), .B(y[2324]), .Z(n27149) );
  NANDN U30514 ( .A(n35364), .B(n27149), .Z(n52103) );
  OR U30515 ( .A(n13813), .B(n52103), .Z(n13814) );
  NAND U30516 ( .A(n52102), .B(n13814), .Z(n13815) );
  NANDN U30517 ( .A(n54494), .B(n13815), .Z(n13816) );
  NANDN U30518 ( .A(n54495), .B(n13816), .Z(n13817) );
  NANDN U30519 ( .A(x[2327]), .B(y[2327]), .Z(n27147) );
  NANDN U30520 ( .A(x[2328]), .B(y[2328]), .Z(n27146) );
  AND U30521 ( .A(n27147), .B(n27146), .Z(n54496) );
  AND U30522 ( .A(n13817), .B(n54496), .Z(n13818) );
  NANDN U30523 ( .A(y[2328]), .B(x[2328]), .Z(n35378) );
  NANDN U30524 ( .A(y[2329]), .B(x[2329]), .Z(n35387) );
  NAND U30525 ( .A(n35378), .B(n35387), .Z(n52101) );
  OR U30526 ( .A(n13818), .B(n52101), .Z(n13819) );
  NAND U30527 ( .A(n54497), .B(n13819), .Z(n13820) );
  NANDN U30528 ( .A(n52100), .B(n13820), .Z(n13821) );
  NANDN U30529 ( .A(x[2331]), .B(y[2331]), .Z(n27144) );
  AND U30530 ( .A(n13821), .B(n27144), .Z(n13822) );
  NAND U30531 ( .A(n35394), .B(n13822), .Z(n13823) );
  NANDN U30532 ( .A(n54499), .B(n13823), .Z(n13824) );
  NAND U30533 ( .A(n13825), .B(n13824), .Z(n13826) );
  NAND U30534 ( .A(n35398), .B(n13826), .Z(n13827) );
  NANDN U30535 ( .A(x[2334]), .B(y[2334]), .Z(n27142) );
  NAND U30536 ( .A(n13827), .B(n27142), .Z(n13828) );
  ANDN U30537 ( .B(x[2335]), .A(y[2335]), .Z(n27140) );
  ANDN U30538 ( .B(n13828), .A(n27140), .Z(n13829) );
  NANDN U30539 ( .A(n35397), .B(n13829), .Z(n13830) );
  NANDN U30540 ( .A(x[2335]), .B(y[2335]), .Z(n27143) );
  AND U30541 ( .A(n13830), .B(n27143), .Z(n13831) );
  NAND U30542 ( .A(n27139), .B(n13831), .Z(n13832) );
  NANDN U30543 ( .A(n54505), .B(n13832), .Z(n13833) );
  NANDN U30544 ( .A(y[2336]), .B(x[2336]), .Z(n27141) );
  NANDN U30545 ( .A(n13833), .B(n27141), .Z(n13834) );
  AND U30546 ( .A(n13835), .B(n13834), .Z(n13836) );
  OR U30547 ( .A(n54507), .B(n13836), .Z(n13837) );
  NAND U30548 ( .A(n54508), .B(n13837), .Z(n13838) );
  NANDN U30549 ( .A(n54509), .B(n13838), .Z(n13839) );
  NANDN U30550 ( .A(n52098), .B(n13839), .Z(n13840) );
  NANDN U30551 ( .A(y[2342]), .B(x[2342]), .Z(n27136) );
  NANDN U30552 ( .A(y[2343]), .B(x[2343]), .Z(n35425) );
  AND U30553 ( .A(n27136), .B(n35425), .Z(n52097) );
  AND U30554 ( .A(n13840), .B(n52097), .Z(n13841) );
  OR U30555 ( .A(n54510), .B(n13841), .Z(n13842) );
  NAND U30556 ( .A(n54511), .B(n13842), .Z(n13843) );
  NANDN U30557 ( .A(n54512), .B(n13843), .Z(n13844) );
  NANDN U30558 ( .A(n52096), .B(n13844), .Z(n13845) );
  NANDN U30559 ( .A(x[2347]), .B(y[2347]), .Z(n27130) );
  NANDN U30560 ( .A(x[2348]), .B(y[2348]), .Z(n27127) );
  AND U30561 ( .A(n27130), .B(n27127), .Z(n52095) );
  AND U30562 ( .A(n13845), .B(n52095), .Z(n13846) );
  OR U30563 ( .A(n54513), .B(n13846), .Z(n13847) );
  NAND U30564 ( .A(n54514), .B(n13847), .Z(n13848) );
  NANDN U30565 ( .A(n54515), .B(n13848), .Z(n13849) );
  NANDN U30566 ( .A(n52094), .B(n13849), .Z(n13850) );
  NANDN U30567 ( .A(y[2352]), .B(x[2352]), .Z(n35443) );
  NANDN U30568 ( .A(y[2353]), .B(x[2353]), .Z(n27123) );
  AND U30569 ( .A(n35443), .B(n27123), .Z(n52093) );
  AND U30570 ( .A(n13850), .B(n52093), .Z(n13851) );
  OR U30571 ( .A(n54517), .B(n13851), .Z(n13852) );
  NAND U30572 ( .A(n54518), .B(n13852), .Z(n13853) );
  NANDN U30573 ( .A(n54519), .B(n13853), .Z(n13854) );
  AND U30574 ( .A(n54520), .B(n13854), .Z(n13855) );
  OR U30575 ( .A(n54521), .B(n13855), .Z(n13856) );
  NAND U30576 ( .A(n54522), .B(n13856), .Z(n13857) );
  NAND U30577 ( .A(n54523), .B(n13857), .Z(n13858) );
  NANDN U30578 ( .A(n54524), .B(n13858), .Z(n13859) );
  NAND U30579 ( .A(n54525), .B(n13859), .Z(n13862) );
  NANDN U30580 ( .A(y[2363]), .B(x[2363]), .Z(n13861) );
  NANDN U30581 ( .A(y[2362]), .B(x[2362]), .Z(n13860) );
  NAND U30582 ( .A(n13861), .B(n13860), .Z(n54526) );
  ANDN U30583 ( .B(n13862), .A(n54526), .Z(n13865) );
  NANDN U30584 ( .A(x[2363]), .B(y[2363]), .Z(n13864) );
  NANDN U30585 ( .A(x[2364]), .B(y[2364]), .Z(n13863) );
  NAND U30586 ( .A(n13864), .B(n13863), .Z(n27113) );
  OR U30587 ( .A(n13865), .B(n27113), .Z(n13868) );
  NANDN U30588 ( .A(y[2365]), .B(x[2365]), .Z(n13867) );
  NANDN U30589 ( .A(y[2364]), .B(x[2364]), .Z(n13866) );
  NAND U30590 ( .A(n13867), .B(n13866), .Z(n54528) );
  ANDN U30591 ( .B(n13868), .A(n54528), .Z(n13871) );
  NANDN U30592 ( .A(x[2365]), .B(y[2365]), .Z(n13870) );
  NANDN U30593 ( .A(x[2366]), .B(y[2366]), .Z(n13869) );
  AND U30594 ( .A(n13870), .B(n13869), .Z(n54529) );
  NANDN U30595 ( .A(n13871), .B(n54529), .Z(n13872) );
  AND U30596 ( .A(n54530), .B(n13872), .Z(n13873) );
  OR U30597 ( .A(n54531), .B(n13873), .Z(n13874) );
  NAND U30598 ( .A(n54532), .B(n13874), .Z(n13875) );
  NANDN U30599 ( .A(n54534), .B(n13875), .Z(n13876) );
  NANDN U30600 ( .A(n54535), .B(n13876), .Z(n13877) );
  AND U30601 ( .A(n54536), .B(n13877), .Z(n13878) );
  OR U30602 ( .A(n54537), .B(n13878), .Z(n13879) );
  NAND U30603 ( .A(n54538), .B(n13879), .Z(n13880) );
  NANDN U30604 ( .A(n54539), .B(n13880), .Z(n13881) );
  NANDN U30605 ( .A(n54540), .B(n13881), .Z(n13882) );
  AND U30606 ( .A(n54541), .B(n13882), .Z(n13883) );
  OR U30607 ( .A(n54542), .B(n13883), .Z(n13884) );
  NAND U30608 ( .A(n54543), .B(n13884), .Z(n13885) );
  NANDN U30609 ( .A(n54544), .B(n13885), .Z(n13886) );
  NANDN U30610 ( .A(n54545), .B(n13886), .Z(n13887) );
  AND U30611 ( .A(n54546), .B(n13887), .Z(n13888) );
  ANDN U30612 ( .B(x[2383]), .A(y[2383]), .Z(n35527) );
  NANDN U30613 ( .A(y[2382]), .B(x[2382]), .Z(n35520) );
  NANDN U30614 ( .A(n35527), .B(n35520), .Z(n52092) );
  OR U30615 ( .A(n13888), .B(n52092), .Z(n13889) );
  NAND U30616 ( .A(n52091), .B(n13889), .Z(n13890) );
  NANDN U30617 ( .A(n54547), .B(n13890), .Z(n13891) );
  NANDN U30618 ( .A(y[2385]), .B(x[2385]), .Z(n35533) );
  NANDN U30619 ( .A(n13891), .B(n35533), .Z(n13892) );
  NANDN U30620 ( .A(x[2385]), .B(y[2385]), .Z(n54548) );
  AND U30621 ( .A(n13892), .B(n54548), .Z(n13893) );
  NAND U30622 ( .A(n27098), .B(n13893), .Z(n13894) );
  NANDN U30623 ( .A(n35532), .B(n13894), .Z(n13895) );
  ANDN U30624 ( .B(x[2387]), .A(y[2387]), .Z(n27095) );
  OR U30625 ( .A(n13895), .B(n27095), .Z(n13896) );
  NAND U30626 ( .A(n13897), .B(n13896), .Z(n13898) );
  NAND U30627 ( .A(n27097), .B(n13898), .Z(n13900) );
  NANDN U30628 ( .A(y[2389]), .B(n13900), .Z(n13899) );
  ANDN U30629 ( .B(x[2390]), .A(y[2390]), .Z(n27092) );
  ANDN U30630 ( .B(n13899), .A(n27092), .Z(n13903) );
  XNOR U30631 ( .A(n13900), .B(y[2389]), .Z(n13901) );
  NAND U30632 ( .A(n13901), .B(x[2389]), .Z(n13902) );
  NAND U30633 ( .A(n13903), .B(n13902), .Z(n13906) );
  NANDN U30634 ( .A(x[2391]), .B(y[2391]), .Z(n13905) );
  NANDN U30635 ( .A(x[2390]), .B(y[2390]), .Z(n13904) );
  NAND U30636 ( .A(n13905), .B(n13904), .Z(n54555) );
  ANDN U30637 ( .B(n13906), .A(n54555), .Z(n13909) );
  NANDN U30638 ( .A(y[2391]), .B(x[2391]), .Z(n13908) );
  NANDN U30639 ( .A(y[2392]), .B(x[2392]), .Z(n13907) );
  NAND U30640 ( .A(n13908), .B(n13907), .Z(n35542) );
  OR U30641 ( .A(n13909), .B(n35542), .Z(n13910) );
  NAND U30642 ( .A(n35544), .B(n13910), .Z(n13911) );
  NAND U30643 ( .A(n27091), .B(n13911), .Z(n13912) );
  NANDN U30644 ( .A(x[2394]), .B(y[2394]), .Z(n35547) );
  NAND U30645 ( .A(n13912), .B(n35547), .Z(n13913) );
  NANDN U30646 ( .A(y[2395]), .B(x[2395]), .Z(n54560) );
  AND U30647 ( .A(n13913), .B(n54560), .Z(n13914) );
  NANDN U30648 ( .A(n27090), .B(n13914), .Z(n13915) );
  ANDN U30649 ( .B(y[2396]), .A(x[2396]), .Z(n54561) );
  ANDN U30650 ( .B(n13915), .A(n54561), .Z(n13916) );
  NANDN U30651 ( .A(x[2395]), .B(y[2395]), .Z(n35548) );
  NAND U30652 ( .A(n13916), .B(n35548), .Z(n13917) );
  NANDN U30653 ( .A(n54562), .B(n13917), .Z(n13918) );
  AND U30654 ( .A(n54563), .B(n13918), .Z(n13919) );
  OR U30655 ( .A(n54564), .B(n13919), .Z(n13920) );
  NAND U30656 ( .A(n54565), .B(n13920), .Z(n13921) );
  NANDN U30657 ( .A(n54566), .B(n13921), .Z(n13922) );
  NANDN U30658 ( .A(x[2401]), .B(y[2401]), .Z(n35569) );
  AND U30659 ( .A(n13922), .B(n35569), .Z(n13923) );
  NAND U30660 ( .A(n35575), .B(n13923), .Z(n13924) );
  NANDN U30661 ( .A(n54570), .B(n13924), .Z(n13925) );
  ANDN U30662 ( .B(x[2403]), .A(y[2403]), .Z(n35578) );
  OR U30663 ( .A(n13925), .B(n35578), .Z(n13926) );
  AND U30664 ( .A(n13927), .B(n13926), .Z(n13929) );
  NANDN U30665 ( .A(y[2405]), .B(x[2405]), .Z(n27086) );
  ANDN U30666 ( .B(x[2404]), .A(y[2404]), .Z(n35577) );
  ANDN U30667 ( .B(n27086), .A(n35577), .Z(n13928) );
  NANDN U30668 ( .A(n13929), .B(n13928), .Z(n13930) );
  AND U30669 ( .A(n27088), .B(n13930), .Z(n13931) );
  NANDN U30670 ( .A(n27083), .B(n13931), .Z(n13932) );
  ANDN U30671 ( .B(x[2407]), .A(y[2407]), .Z(n54576) );
  ANDN U30672 ( .B(n13932), .A(n54576), .Z(n13933) );
  NANDN U30673 ( .A(n27085), .B(n13933), .Z(n13934) );
  AND U30674 ( .A(n13935), .B(n13934), .Z(n13936) );
  ANDN U30675 ( .B(x[2408]), .A(y[2408]), .Z(n35585) );
  ANDN U30676 ( .B(x[2409]), .A(y[2409]), .Z(n35591) );
  OR U30677 ( .A(n35585), .B(n35591), .Z(n54577) );
  OR U30678 ( .A(n13936), .B(n54577), .Z(n13937) );
  NAND U30679 ( .A(n54578), .B(n13937), .Z(n13938) );
  NANDN U30680 ( .A(n52088), .B(n13938), .Z(n13939) );
  NANDN U30681 ( .A(n54580), .B(n13939), .Z(n13940) );
  AND U30682 ( .A(n54581), .B(n13940), .Z(n13941) );
  NANDN U30683 ( .A(x[2413]), .B(y[2413]), .Z(n27079) );
  NANDN U30684 ( .A(n13941), .B(n27079), .Z(n13942) );
  ANDN U30685 ( .B(y[2414]), .A(x[2414]), .Z(n35604) );
  OR U30686 ( .A(n13942), .B(n35604), .Z(n13943) );
  NAND U30687 ( .A(n54583), .B(n13943), .Z(n13944) );
  NANDN U30688 ( .A(n35605), .B(n13944), .Z(n13945) );
  NAND U30689 ( .A(n54585), .B(n13945), .Z(n13946) );
  NANDN U30690 ( .A(n54586), .B(n13946), .Z(n13947) );
  AND U30691 ( .A(n54587), .B(n13947), .Z(n13950) );
  NANDN U30692 ( .A(x[2419]), .B(y[2419]), .Z(n13949) );
  NANDN U30693 ( .A(x[2420]), .B(y[2420]), .Z(n13948) );
  AND U30694 ( .A(n13949), .B(n13948), .Z(n54588) );
  NANDN U30695 ( .A(n13950), .B(n54588), .Z(n13953) );
  NANDN U30696 ( .A(y[2421]), .B(x[2421]), .Z(n13952) );
  NANDN U30697 ( .A(y[2420]), .B(x[2420]), .Z(n13951) );
  NAND U30698 ( .A(n13952), .B(n13951), .Z(n54589) );
  ANDN U30699 ( .B(n13953), .A(n54589), .Z(n13956) );
  NANDN U30700 ( .A(x[2421]), .B(y[2421]), .Z(n13955) );
  NANDN U30701 ( .A(x[2422]), .B(y[2422]), .Z(n13954) );
  NAND U30702 ( .A(n13955), .B(n13954), .Z(n35612) );
  OR U30703 ( .A(n13956), .B(n35612), .Z(n13959) );
  NANDN U30704 ( .A(y[2423]), .B(x[2423]), .Z(n13958) );
  NANDN U30705 ( .A(y[2422]), .B(x[2422]), .Z(n13957) );
  AND U30706 ( .A(n13958), .B(n13957), .Z(n35614) );
  AND U30707 ( .A(n13959), .B(n35614), .Z(n13960) );
  NANDN U30708 ( .A(x[2423]), .B(y[2423]), .Z(n35617) );
  NANDN U30709 ( .A(x[2424]), .B(y[2424]), .Z(n35623) );
  NAND U30710 ( .A(n35617), .B(n35623), .Z(n54592) );
  OR U30711 ( .A(n13960), .B(n54592), .Z(n13961) );
  NAND U30712 ( .A(n54593), .B(n13961), .Z(n13962) );
  NANDN U30713 ( .A(n52087), .B(n13962), .Z(n13963) );
  NAND U30714 ( .A(n54594), .B(n13963), .Z(n13964) );
  AND U30715 ( .A(n13965), .B(n13964), .Z(n13967) );
  ANDN U30716 ( .B(x[2429]), .A(y[2429]), .Z(n35639) );
  NANDN U30717 ( .A(y[2428]), .B(x[2428]), .Z(n13966) );
  NANDN U30718 ( .A(n35639), .B(n13966), .Z(n54597) );
  OR U30719 ( .A(n13967), .B(n54597), .Z(n13968) );
  NAND U30720 ( .A(n54600), .B(n13968), .Z(n13969) );
  NANDN U30721 ( .A(n52086), .B(n13969), .Z(n13970) );
  NANDN U30722 ( .A(n54602), .B(n13970), .Z(n13971) );
  AND U30723 ( .A(n54603), .B(n13971), .Z(n13972) );
  NANDN U30724 ( .A(x[2433]), .B(y[2433]), .Z(n35649) );
  NANDN U30725 ( .A(x[2434]), .B(y[2434]), .Z(n35656) );
  NAND U30726 ( .A(n35649), .B(n35656), .Z(n54604) );
  OR U30727 ( .A(n13972), .B(n54604), .Z(n13973) );
  NANDN U30728 ( .A(y[2434]), .B(x[2434]), .Z(n27075) );
  AND U30729 ( .A(n13973), .B(n27075), .Z(n13974) );
  NANDN U30730 ( .A(y[2435]), .B(x[2435]), .Z(n27073) );
  NAND U30731 ( .A(n13974), .B(n27073), .Z(n13975) );
  NANDN U30732 ( .A(n54606), .B(n13975), .Z(n13976) );
  XNOR U30733 ( .A(y[2436]), .B(x[2436]), .Z(n27074) );
  NAND U30734 ( .A(n13976), .B(n27074), .Z(n13977) );
  NANDN U30735 ( .A(n54608), .B(n13977), .Z(n13978) );
  AND U30736 ( .A(n54609), .B(n13978), .Z(n13979) );
  OR U30737 ( .A(n54610), .B(n13979), .Z(n13980) );
  NAND U30738 ( .A(n54611), .B(n13980), .Z(n13981) );
  NANDN U30739 ( .A(n54612), .B(n13981), .Z(n13982) );
  NAND U30740 ( .A(n54613), .B(n13982), .Z(n13983) );
  NANDN U30741 ( .A(n54614), .B(n13983), .Z(n13986) );
  NANDN U30742 ( .A(y[2442]), .B(x[2442]), .Z(n35673) );
  NANDN U30743 ( .A(y[2443]), .B(x[2443]), .Z(n27069) );
  NAND U30744 ( .A(n35673), .B(n27069), .Z(n13984) );
  NAND U30745 ( .A(n13985), .B(n13984), .Z(n52085) );
  AND U30746 ( .A(n13986), .B(n52085), .Z(n13987) );
  ANDN U30747 ( .B(y[2444]), .A(x[2444]), .Z(n27066) );
  OR U30748 ( .A(n13987), .B(n27066), .Z(n13988) );
  NANDN U30749 ( .A(y[2444]), .B(x[2444]), .Z(n27068) );
  NANDN U30750 ( .A(y[2445]), .B(x[2445]), .Z(n27065) );
  AND U30751 ( .A(n27068), .B(n27065), .Z(n54617) );
  AND U30752 ( .A(n13988), .B(n54617), .Z(n13989) );
  XNOR U30753 ( .A(y[2446]), .B(x[2446]), .Z(n27064) );
  NANDN U30754 ( .A(x[2445]), .B(y[2445]), .Z(n27067) );
  NAND U30755 ( .A(n27064), .B(n27067), .Z(n52084) );
  OR U30756 ( .A(n13989), .B(n52084), .Z(n13990) );
  NAND U30757 ( .A(n54619), .B(n13990), .Z(n13991) );
  NANDN U30758 ( .A(n35683), .B(n13991), .Z(n13992) );
  ANDN U30759 ( .B(n13993), .A(n13992), .Z(n13995) );
  ANDN U30760 ( .B(x[2449]), .A(y[2449]), .Z(n35694) );
  NANDN U30761 ( .A(y[2448]), .B(x[2448]), .Z(n13994) );
  NANDN U30762 ( .A(n35694), .B(n13994), .Z(n54622) );
  OR U30763 ( .A(n13995), .B(n54622), .Z(n13996) );
  NAND U30764 ( .A(n54623), .B(n13996), .Z(n13997) );
  NANDN U30765 ( .A(n52083), .B(n13997), .Z(n13998) );
  NANDN U30766 ( .A(x[2451]), .B(y[2451]), .Z(n35699) );
  NANDN U30767 ( .A(x[2452]), .B(y[2452]), .Z(n35704) );
  AND U30768 ( .A(n35699), .B(n35704), .Z(n52082) );
  AND U30769 ( .A(n13998), .B(n52082), .Z(n13999) );
  NANDN U30770 ( .A(y[2452]), .B(x[2452]), .Z(n27062) );
  ANDN U30771 ( .B(x[2453]), .A(y[2453]), .Z(n35708) );
  ANDN U30772 ( .B(n27062), .A(n35708), .Z(n54624) );
  NANDN U30773 ( .A(n13999), .B(n54624), .Z(n14000) );
  NAND U30774 ( .A(n14001), .B(n14000), .Z(n14002) );
  ANDN U30775 ( .B(x[2454]), .A(y[2454]), .Z(n54626) );
  ANDN U30776 ( .B(n14002), .A(n54626), .Z(n14003) );
  NAND U30777 ( .A(n35712), .B(n14003), .Z(n14004) );
  NAND U30778 ( .A(n27061), .B(n14004), .Z(n14005) );
  ANDN U30779 ( .B(y[2456]), .A(x[2456]), .Z(n27057) );
  OR U30780 ( .A(n14005), .B(n27057), .Z(n14006) );
  AND U30781 ( .A(n35711), .B(n14006), .Z(n14007) );
  NANDN U30782 ( .A(y[2457]), .B(x[2457]), .Z(n27055) );
  NAND U30783 ( .A(n14007), .B(n27055), .Z(n14008) );
  NANDN U30784 ( .A(x[2458]), .B(y[2458]), .Z(n27054) );
  AND U30785 ( .A(n14008), .B(n27054), .Z(n14009) );
  NAND U30786 ( .A(n27058), .B(n14009), .Z(n14010) );
  NANDN U30787 ( .A(y[2459]), .B(x[2459]), .Z(n54632) );
  AND U30788 ( .A(n14010), .B(n54632), .Z(n14011) );
  NANDN U30789 ( .A(y[2458]), .B(x[2458]), .Z(n27056) );
  NAND U30790 ( .A(n14011), .B(n27056), .Z(n14012) );
  ANDN U30791 ( .B(y[2459]), .A(x[2459]), .Z(n27053) );
  ANDN U30792 ( .B(n14012), .A(n27053), .Z(n14013) );
  NANDN U30793 ( .A(n27050), .B(n14013), .Z(n14014) );
  NANDN U30794 ( .A(n54634), .B(n14014), .Z(n14015) );
  AND U30795 ( .A(n54635), .B(n14015), .Z(n14016) );
  ANDN U30796 ( .B(x[2463]), .A(y[2463]), .Z(n35726) );
  NANDN U30797 ( .A(y[2462]), .B(x[2462]), .Z(n27048) );
  NANDN U30798 ( .A(n35726), .B(n27048), .Z(n54636) );
  OR U30799 ( .A(n14016), .B(n54636), .Z(n14017) );
  NAND U30800 ( .A(n52080), .B(n14017), .Z(n14018) );
  NANDN U30801 ( .A(n54637), .B(n14018), .Z(n14019) );
  NANDN U30802 ( .A(n54638), .B(n14019), .Z(n14020) );
  AND U30803 ( .A(n54639), .B(n14020), .Z(n14021) );
  NANDN U30804 ( .A(x[2467]), .B(y[2467]), .Z(n35738) );
  NANDN U30805 ( .A(x[2468]), .B(y[2468]), .Z(n27045) );
  NAND U30806 ( .A(n35738), .B(n27045), .Z(n54640) );
  OR U30807 ( .A(n14021), .B(n54640), .Z(n14022) );
  NAND U30808 ( .A(n52079), .B(n14022), .Z(n14023) );
  NANDN U30809 ( .A(n54641), .B(n14023), .Z(n14024) );
  NANDN U30810 ( .A(n54644), .B(n14024), .Z(n14025) );
  AND U30811 ( .A(n54645), .B(n14025), .Z(n14026) );
  OR U30812 ( .A(n54646), .B(n14026), .Z(n14027) );
  NAND U30813 ( .A(n54647), .B(n14027), .Z(n14028) );
  NANDN U30814 ( .A(n54648), .B(n14028), .Z(n14029) );
  NAND U30815 ( .A(n54650), .B(n14029), .Z(n14030) );
  NAND U30816 ( .A(n27037), .B(n14030), .Z(n14031) );
  NAND U30817 ( .A(n35768), .B(n14031), .Z(n14032) );
  NANDN U30818 ( .A(y[2477]), .B(x[2477]), .Z(n52078) );
  AND U30819 ( .A(n14032), .B(n52078), .Z(n14033) );
  ANDN U30820 ( .B(y[2478]), .A(x[2478]), .Z(n35771) );
  OR U30821 ( .A(n14033), .B(n35771), .Z(n14034) );
  NANDN U30822 ( .A(n54652), .B(n14034), .Z(n14035) );
  AND U30823 ( .A(n54653), .B(n14035), .Z(n14036) );
  OR U30824 ( .A(n54654), .B(n14036), .Z(n14037) );
  NAND U30825 ( .A(n54655), .B(n14037), .Z(n14038) );
  NANDN U30826 ( .A(n54656), .B(n14038), .Z(n14039) );
  NANDN U30827 ( .A(n52075), .B(n14039), .Z(n14041) );
  NANDN U30828 ( .A(y[2484]), .B(x[2484]), .Z(n14040) );
  NANDN U30829 ( .A(y[2485]), .B(x[2485]), .Z(n27029) );
  AND U30830 ( .A(n14040), .B(n27029), .Z(n52074) );
  AND U30831 ( .A(n14041), .B(n52074), .Z(n14042) );
  ANDN U30832 ( .B(y[2485]), .A(x[2485]), .Z(n35791) );
  NANDN U30833 ( .A(x[2486]), .B(y[2486]), .Z(n27026) );
  NANDN U30834 ( .A(n35791), .B(n27026), .Z(n52073) );
  OR U30835 ( .A(n14042), .B(n52073), .Z(n14043) );
  NAND U30836 ( .A(n52072), .B(n14043), .Z(n14044) );
  NANDN U30837 ( .A(n54659), .B(n14044), .Z(n14045) );
  NANDN U30838 ( .A(n54660), .B(n14045), .Z(n14046) );
  AND U30839 ( .A(n54661), .B(n14046), .Z(n14047) );
  OR U30840 ( .A(n54662), .B(n14047), .Z(n14048) );
  NAND U30841 ( .A(n54663), .B(n14048), .Z(n14049) );
  NANDN U30842 ( .A(n54664), .B(n14049), .Z(n14050) );
  NANDN U30843 ( .A(n54665), .B(n14050), .Z(n14051) );
  AND U30844 ( .A(n54666), .B(n14051), .Z(n14052) );
  OR U30845 ( .A(n54667), .B(n14052), .Z(n14053) );
  NAND U30846 ( .A(n54668), .B(n14053), .Z(n14054) );
  NANDN U30847 ( .A(n27020), .B(n14054), .Z(n14055) );
  XNOR U30848 ( .A(x[2498]), .B(y[2498]), .Z(n35832) );
  NANDN U30849 ( .A(n14055), .B(n35832), .Z(n14056) );
  NANDN U30850 ( .A(n54669), .B(n14056), .Z(n14057) );
  AND U30851 ( .A(n54671), .B(n14057), .Z(n14058) );
  OR U30852 ( .A(n54672), .B(n14058), .Z(n14059) );
  NAND U30853 ( .A(n54673), .B(n14059), .Z(n14060) );
  NANDN U30854 ( .A(n54674), .B(n14060), .Z(n14061) );
  AND U30855 ( .A(n54675), .B(n14061), .Z(n14062) );
  NANDN U30856 ( .A(y[2504]), .B(x[2504]), .Z(n27015) );
  ANDN U30857 ( .B(x[2505]), .A(y[2505]), .Z(n27013) );
  ANDN U30858 ( .B(n27015), .A(n27013), .Z(n54676) );
  NANDN U30859 ( .A(n14062), .B(n54676), .Z(n14063) );
  NANDN U30860 ( .A(n54677), .B(n14063), .Z(n14064) );
  AND U30861 ( .A(n54678), .B(n14064), .Z(n14065) );
  OR U30862 ( .A(n54679), .B(n14065), .Z(n14066) );
  NAND U30863 ( .A(n54680), .B(n14066), .Z(n14067) );
  NANDN U30864 ( .A(n54681), .B(n14067), .Z(n14068) );
  NAND U30865 ( .A(n54682), .B(n14068), .Z(n14069) );
  ANDN U30866 ( .B(y[2512]), .A(x[2512]), .Z(n27006) );
  ANDN U30867 ( .B(n14069), .A(n27006), .Z(n14070) );
  NANDN U30868 ( .A(n54683), .B(n14070), .Z(n14071) );
  NAND U30869 ( .A(n54684), .B(n14071), .Z(n14072) );
  ANDN U30870 ( .B(x[2513]), .A(y[2513]), .Z(n27003) );
  OR U30871 ( .A(n14072), .B(n27003), .Z(n14073) );
  NAND U30872 ( .A(n14074), .B(n14073), .Z(n14075) );
  AND U30873 ( .A(n27005), .B(n14075), .Z(n14076) );
  NANDN U30874 ( .A(y[2515]), .B(x[2515]), .Z(n27002) );
  NAND U30875 ( .A(n14076), .B(n27002), .Z(n14077) );
  ANDN U30876 ( .B(y[2516]), .A(x[2516]), .Z(n26998) );
  ANDN U30877 ( .B(n14077), .A(n26998), .Z(n14078) );
  ANDN U30878 ( .B(y[2515]), .A(x[2515]), .Z(n35879) );
  ANDN U30879 ( .B(n14078), .A(n35879), .Z(n14080) );
  NANDN U30880 ( .A(y[2517]), .B(x[2517]), .Z(n54691) );
  ANDN U30881 ( .B(x[2516]), .A(y[2516]), .Z(n27001) );
  ANDN U30882 ( .B(n54691), .A(n27001), .Z(n14079) );
  NANDN U30883 ( .A(n14080), .B(n14079), .Z(n14081) );
  ANDN U30884 ( .B(y[2518]), .A(x[2518]), .Z(n54692) );
  ANDN U30885 ( .B(n14081), .A(n54692), .Z(n14082) );
  NANDN U30886 ( .A(x[2517]), .B(y[2517]), .Z(n27000) );
  AND U30887 ( .A(n14082), .B(n27000), .Z(n14083) );
  OR U30888 ( .A(n54693), .B(n14083), .Z(n14084) );
  NAND U30889 ( .A(n54694), .B(n14084), .Z(n14085) );
  NANDN U30890 ( .A(n54695), .B(n14085), .Z(n14086) );
  NAND U30891 ( .A(n52069), .B(n14086), .Z(n14087) );
  NANDN U30892 ( .A(n54696), .B(n14087), .Z(n14088) );
  NANDN U30893 ( .A(x[2523]), .B(y[2523]), .Z(n35899) );
  NANDN U30894 ( .A(x[2524]), .B(y[2524]), .Z(n35908) );
  AND U30895 ( .A(n35899), .B(n35908), .Z(n54697) );
  AND U30896 ( .A(n14088), .B(n54697), .Z(n14089) );
  ANDN U30897 ( .B(x[2524]), .A(y[2524]), .Z(n35903) );
  ANDN U30898 ( .B(x[2525]), .A(y[2525]), .Z(n35913) );
  OR U30899 ( .A(n35903), .B(n35913), .Z(n54698) );
  OR U30900 ( .A(n14089), .B(n54698), .Z(n14090) );
  NAND U30901 ( .A(n54699), .B(n14090), .Z(n14091) );
  NANDN U30902 ( .A(n52068), .B(n14091), .Z(n14092) );
  NANDN U30903 ( .A(x[2527]), .B(y[2527]), .Z(n52067) );
  AND U30904 ( .A(n14092), .B(n52067), .Z(n14093) );
  NAND U30905 ( .A(n26993), .B(n14093), .Z(n14094) );
  NANDN U30906 ( .A(n26990), .B(n14094), .Z(n14095) );
  ANDN U30907 ( .B(x[2528]), .A(y[2528]), .Z(n52066) );
  OR U30908 ( .A(n14095), .B(n52066), .Z(n14096) );
  AND U30909 ( .A(n14097), .B(n14096), .Z(n14098) );
  ANDN U30910 ( .B(x[2531]), .A(y[2531]), .Z(n35928) );
  NANDN U30911 ( .A(y[2530]), .B(x[2530]), .Z(n26991) );
  NANDN U30912 ( .A(n35928), .B(n26991), .Z(n54703) );
  OR U30913 ( .A(n14098), .B(n54703), .Z(n14099) );
  NAND U30914 ( .A(n54704), .B(n14099), .Z(n14100) );
  NANDN U30915 ( .A(n52064), .B(n14100), .Z(n14101) );
  NANDN U30916 ( .A(n54705), .B(n14101), .Z(n14102) );
  AND U30917 ( .A(n54706), .B(n14102), .Z(n14103) );
  ANDN U30918 ( .B(n14104), .A(n14103), .Z(n14105) );
  NANDN U30919 ( .A(y[2536]), .B(x[2536]), .Z(n26985) );
  NANDN U30920 ( .A(y[2537]), .B(x[2537]), .Z(n26982) );
  AND U30921 ( .A(n26985), .B(n26982), .Z(n54708) );
  NANDN U30922 ( .A(n14105), .B(n54708), .Z(n14106) );
  NAND U30923 ( .A(n52063), .B(n14106), .Z(n14107) );
  ANDN U30924 ( .B(y[2537]), .A(x[2537]), .Z(n26983) );
  OR U30925 ( .A(n14107), .B(n26983), .Z(n14109) );
  NANDN U30926 ( .A(y[2538]), .B(x[2538]), .Z(n14108) );
  NANDN U30927 ( .A(y[2539]), .B(x[2539]), .Z(n35945) );
  AND U30928 ( .A(n14108), .B(n35945), .Z(n54710) );
  AND U30929 ( .A(n14109), .B(n54710), .Z(n14111) );
  ANDN U30930 ( .B(y[2539]), .A(x[2539]), .Z(n26981) );
  XNOR U30931 ( .A(x[2540]), .B(y[2540]), .Z(n14110) );
  NANDN U30932 ( .A(n26981), .B(n14110), .Z(n54711) );
  OR U30933 ( .A(n14111), .B(n54711), .Z(n14112) );
  NAND U30934 ( .A(n54712), .B(n14112), .Z(n14113) );
  NANDN U30935 ( .A(n52060), .B(n14113), .Z(n14114) );
  NANDN U30936 ( .A(n54713), .B(n14114), .Z(n14115) );
  AND U30937 ( .A(n54714), .B(n14115), .Z(n14116) );
  ANDN U30938 ( .B(x[2544]), .A(y[2544]), .Z(n26977) );
  ANDN U30939 ( .B(x[2545]), .A(y[2545]), .Z(n35968) );
  OR U30940 ( .A(n26977), .B(n35968), .Z(n54715) );
  OR U30941 ( .A(n14116), .B(n54715), .Z(n14117) );
  NAND U30942 ( .A(n54716), .B(n14117), .Z(n14118) );
  NANDN U30943 ( .A(n54717), .B(n14118), .Z(n14119) );
  NANDN U30944 ( .A(n54718), .B(n14119), .Z(n14120) );
  AND U30945 ( .A(n54719), .B(n14120), .Z(n14122) );
  NANDN U30946 ( .A(x[2549]), .B(y[2549]), .Z(n52058) );
  XOR U30947 ( .A(x[2550]), .B(y[2550]), .Z(n35983) );
  ANDN U30948 ( .B(n52058), .A(n35983), .Z(n14121) );
  NANDN U30949 ( .A(n14122), .B(n14121), .Z(n14123) );
  NANDN U30950 ( .A(n54721), .B(n14123), .Z(n14124) );
  AND U30951 ( .A(n54722), .B(n14124), .Z(n14125) );
  OR U30952 ( .A(n54723), .B(n14125), .Z(n14126) );
  NAND U30953 ( .A(n54724), .B(n14126), .Z(n14127) );
  NANDN U30954 ( .A(n54725), .B(n14127), .Z(n14128) );
  NAND U30955 ( .A(n54726), .B(n14128), .Z(n14129) );
  ANDN U30956 ( .B(x[2557]), .A(y[2557]), .Z(n36005) );
  ANDN U30957 ( .B(n14129), .A(n36005), .Z(n14130) );
  NANDN U30958 ( .A(n54727), .B(n14130), .Z(n14132) );
  NANDN U30959 ( .A(x[2557]), .B(y[2557]), .Z(n54728) );
  NANDN U30960 ( .A(x[2558]), .B(y[2558]), .Z(n54730) );
  AND U30961 ( .A(n54728), .B(n54730), .Z(n14131) );
  NAND U30962 ( .A(n14132), .B(n14131), .Z(n14133) );
  ANDN U30963 ( .B(x[2559]), .A(y[2559]), .Z(n54731) );
  ANDN U30964 ( .B(n14133), .A(n54731), .Z(n14134) );
  NANDN U30965 ( .A(y[2558]), .B(x[2558]), .Z(n36006) );
  NAND U30966 ( .A(n14134), .B(n36006), .Z(n14135) );
  NANDN U30967 ( .A(n54732), .B(n14135), .Z(n14136) );
  AND U30968 ( .A(n54734), .B(n14136), .Z(n14137) );
  NANDN U30969 ( .A(x[2561]), .B(y[2561]), .Z(n36014) );
  NANDN U30970 ( .A(x[2562]), .B(y[2562]), .Z(n36021) );
  NAND U30971 ( .A(n36014), .B(n36021), .Z(n54735) );
  OR U30972 ( .A(n14137), .B(n54735), .Z(n14138) );
  NAND U30973 ( .A(n54736), .B(n14138), .Z(n14139) );
  NANDN U30974 ( .A(x[2563]), .B(y[2563]), .Z(n52057) );
  AND U30975 ( .A(n14139), .B(n52057), .Z(n14140) );
  NAND U30976 ( .A(n26969), .B(n14140), .Z(n14141) );
  NAND U30977 ( .A(n14142), .B(n14141), .Z(n14143) );
  NAND U30978 ( .A(n54740), .B(n14143), .Z(n14144) );
  ANDN U30979 ( .B(y[2565]), .A(x[2565]), .Z(n26968) );
  OR U30980 ( .A(n14144), .B(n26968), .Z(n14145) );
  AND U30981 ( .A(n54741), .B(n14145), .Z(n14146) );
  OR U30982 ( .A(n54742), .B(n14146), .Z(n14147) );
  NAND U30983 ( .A(n54743), .B(n14147), .Z(n14148) );
  NANDN U30984 ( .A(n54744), .B(n14148), .Z(n14149) );
  NANDN U30985 ( .A(n52056), .B(n14149), .Z(n14150) );
  NANDN U30986 ( .A(x[2571]), .B(y[2571]), .Z(n26964) );
  NANDN U30987 ( .A(x[2572]), .B(y[2572]), .Z(n26959) );
  AND U30988 ( .A(n26964), .B(n26959), .Z(n52055) );
  AND U30989 ( .A(n14150), .B(n52055), .Z(n14151) );
  OR U30990 ( .A(n54745), .B(n14151), .Z(n14152) );
  NAND U30991 ( .A(n54746), .B(n14152), .Z(n14153) );
  NANDN U30992 ( .A(n54747), .B(n14153), .Z(n14154) );
  ANDN U30993 ( .B(y[2575]), .A(x[2575]), .Z(n54748) );
  ANDN U30994 ( .B(n14154), .A(n54748), .Z(n14155) );
  NAND U30995 ( .A(n26957), .B(n14155), .Z(n14156) );
  NANDN U30996 ( .A(n54750), .B(n14156), .Z(n14157) );
  NANDN U30997 ( .A(y[2577]), .B(x[2577]), .Z(n26955) );
  NANDN U30998 ( .A(n14157), .B(n26955), .Z(n14158) );
  AND U30999 ( .A(n14159), .B(n14158), .Z(n14161) );
  NANDN U31000 ( .A(y[2579]), .B(x[2579]), .Z(n26951) );
  ANDN U31001 ( .B(x[2578]), .A(y[2578]), .Z(n26954) );
  ANDN U31002 ( .B(n26951), .A(n26954), .Z(n14160) );
  NANDN U31003 ( .A(n14161), .B(n14160), .Z(n14162) );
  NANDN U31004 ( .A(n26952), .B(n14162), .Z(n14163) );
  ANDN U31005 ( .B(y[2580]), .A(x[2580]), .Z(n26948) );
  OR U31006 ( .A(n14163), .B(n26948), .Z(n14164) );
  NANDN U31007 ( .A(y[2581]), .B(x[2581]), .Z(n36064) );
  AND U31008 ( .A(n14164), .B(n36064), .Z(n14165) );
  NAND U31009 ( .A(n26950), .B(n14165), .Z(n14166) );
  AND U31010 ( .A(n14167), .B(n14166), .Z(n14168) );
  OR U31011 ( .A(n54758), .B(n14168), .Z(n14169) );
  NAND U31012 ( .A(n54759), .B(n14169), .Z(n14170) );
  NANDN U31013 ( .A(n54760), .B(n14170), .Z(n14171) );
  NANDN U31014 ( .A(n54761), .B(n14171), .Z(n14172) );
  AND U31015 ( .A(n54762), .B(n14172), .Z(n14174) );
  NANDN U31016 ( .A(x[2587]), .B(y[2587]), .Z(n36084) );
  XNOR U31017 ( .A(y[2588]), .B(x[2588]), .Z(n14173) );
  AND U31018 ( .A(n36084), .B(n14173), .Z(n54763) );
  NANDN U31019 ( .A(n14174), .B(n54763), .Z(n14175) );
  NANDN U31020 ( .A(n52054), .B(n14175), .Z(n14176) );
  XNOR U31021 ( .A(y[2590]), .B(x[2590]), .Z(n36095) );
  NANDN U31022 ( .A(x[2589]), .B(y[2589]), .Z(n26946) );
  AND U31023 ( .A(n36095), .B(n26946), .Z(n52053) );
  AND U31024 ( .A(n14176), .B(n52053), .Z(n14178) );
  NANDN U31025 ( .A(y[2590]), .B(x[2590]), .Z(n14177) );
  NANDN U31026 ( .A(y[2591]), .B(x[2591]), .Z(n26942) );
  NAND U31027 ( .A(n14177), .B(n26942), .Z(n54765) );
  OR U31028 ( .A(n14178), .B(n54765), .Z(n14179) );
  AND U31029 ( .A(n54766), .B(n14179), .Z(n14181) );
  NANDN U31030 ( .A(y[2592]), .B(x[2592]), .Z(n14180) );
  ANDN U31031 ( .B(x[2593]), .A(y[2593]), .Z(n36106) );
  ANDN U31032 ( .B(n14180), .A(n36106), .Z(n54767) );
  NANDN U31033 ( .A(n14181), .B(n54767), .Z(n14182) );
  NANDN U31034 ( .A(n52052), .B(n14182), .Z(n14183) );
  AND U31035 ( .A(n54768), .B(n14183), .Z(n14185) );
  NANDN U31036 ( .A(x[2595]), .B(y[2595]), .Z(n26940) );
  NANDN U31037 ( .A(x[2596]), .B(y[2596]), .Z(n14184) );
  NAND U31038 ( .A(n26940), .B(n14184), .Z(n54769) );
  OR U31039 ( .A(n14185), .B(n54769), .Z(n14186) );
  AND U31040 ( .A(n54770), .B(n14186), .Z(n14187) );
  OR U31041 ( .A(n54771), .B(n14187), .Z(n14188) );
  NAND U31042 ( .A(n54772), .B(n14188), .Z(n14189) );
  NANDN U31043 ( .A(n54773), .B(n14189), .Z(n14190) );
  NANDN U31044 ( .A(n54774), .B(n14190), .Z(n14191) );
  AND U31045 ( .A(n54775), .B(n14191), .Z(n14192) );
  OR U31046 ( .A(n54776), .B(n14192), .Z(n14193) );
  NAND U31047 ( .A(n54777), .B(n14193), .Z(n14194) );
  NANDN U31048 ( .A(n54778), .B(n14194), .Z(n14195) );
  NANDN U31049 ( .A(n54779), .B(n14195), .Z(n14196) );
  AND U31050 ( .A(n54780), .B(n14196), .Z(n14197) );
  OR U31051 ( .A(n54781), .B(n14197), .Z(n14198) );
  NAND U31052 ( .A(n54782), .B(n14198), .Z(n14199) );
  NANDN U31053 ( .A(n54784), .B(n14199), .Z(n14200) );
  AND U31054 ( .A(n54785), .B(n14200), .Z(n14202) );
  NANDN U31055 ( .A(x[2611]), .B(y[2611]), .Z(n26928) );
  XNOR U31056 ( .A(y[2612]), .B(x[2612]), .Z(n14201) );
  AND U31057 ( .A(n26928), .B(n14201), .Z(n54786) );
  NANDN U31058 ( .A(n14202), .B(n54786), .Z(n14203) );
  NANDN U31059 ( .A(n52051), .B(n14203), .Z(n14204) );
  AND U31060 ( .A(n54787), .B(n14204), .Z(n14206) );
  ANDN U31061 ( .B(x[2615]), .A(y[2615]), .Z(n36178) );
  NANDN U31062 ( .A(y[2614]), .B(x[2614]), .Z(n14205) );
  NANDN U31063 ( .A(n36178), .B(n14205), .Z(n54788) );
  OR U31064 ( .A(n14206), .B(n54788), .Z(n14207) );
  NANDN U31065 ( .A(x[2615]), .B(y[2615]), .Z(n54790) );
  AND U31066 ( .A(n14207), .B(n54790), .Z(n14208) );
  XNOR U31067 ( .A(x[2616]), .B(y[2616]), .Z(n36177) );
  NAND U31068 ( .A(n14208), .B(n36177), .Z(n14209) );
  NANDN U31069 ( .A(n54791), .B(n14209), .Z(n14210) );
  AND U31070 ( .A(n36183), .B(n14210), .Z(n14211) );
  NANDN U31071 ( .A(x[2617]), .B(y[2617]), .Z(n54792) );
  NAND U31072 ( .A(n14211), .B(n54792), .Z(n14212) );
  NANDN U31073 ( .A(n54793), .B(n14212), .Z(n14213) );
  AND U31074 ( .A(n54794), .B(n14213), .Z(n14214) );
  OR U31075 ( .A(n54795), .B(n14214), .Z(n14215) );
  NAND U31076 ( .A(n54796), .B(n14215), .Z(n14216) );
  NANDN U31077 ( .A(n54798), .B(n14216), .Z(n14217) );
  NANDN U31078 ( .A(n54799), .B(n14217), .Z(n14218) );
  AND U31079 ( .A(n54800), .B(n14218), .Z(n14219) );
  OR U31080 ( .A(n54801), .B(n14219), .Z(n14220) );
  NAND U31081 ( .A(n54802), .B(n14220), .Z(n14221) );
  NANDN U31082 ( .A(n54803), .B(n14221), .Z(n14222) );
  AND U31083 ( .A(n54804), .B(n14222), .Z(n14223) );
  ANDN U31084 ( .B(n14224), .A(n14223), .Z(n14225) );
  ANDN U31085 ( .B(y[2629]), .A(x[2629]), .Z(n52048) );
  ANDN U31086 ( .B(n14225), .A(n52048), .Z(n14226) );
  OR U31087 ( .A(n54805), .B(n14226), .Z(n14227) );
  AND U31088 ( .A(n14228), .B(n14227), .Z(n14230) );
  ANDN U31089 ( .B(x[2633]), .A(y[2633]), .Z(n36230) );
  NANDN U31090 ( .A(y[2632]), .B(x[2632]), .Z(n14229) );
  NANDN U31091 ( .A(n36230), .B(n14229), .Z(n54807) );
  OR U31092 ( .A(n14230), .B(n54807), .Z(n14231) );
  NAND U31093 ( .A(n54808), .B(n14231), .Z(n14232) );
  NANDN U31094 ( .A(n52046), .B(n14232), .Z(n14233) );
  NANDN U31095 ( .A(n54809), .B(n14233), .Z(n14234) );
  NANDN U31096 ( .A(y[2636]), .B(x[2636]), .Z(n26908) );
  NANDN U31097 ( .A(y[2637]), .B(x[2637]), .Z(n36240) );
  AND U31098 ( .A(n26908), .B(n36240), .Z(n52045) );
  AND U31099 ( .A(n14234), .B(n52045), .Z(n14235) );
  XNOR U31100 ( .A(y[2638]), .B(x[2638]), .Z(n36238) );
  NANDN U31101 ( .A(x[2637]), .B(y[2637]), .Z(n26906) );
  NAND U31102 ( .A(n36238), .B(n26906), .Z(n54811) );
  OR U31103 ( .A(n14235), .B(n54811), .Z(n14236) );
  NAND U31104 ( .A(n54812), .B(n14236), .Z(n14237) );
  NANDN U31105 ( .A(n52044), .B(n14237), .Z(n14238) );
  NANDN U31106 ( .A(n54813), .B(n14238), .Z(n14239) );
  NANDN U31107 ( .A(x[2641]), .B(y[2641]), .Z(n26904) );
  NANDN U31108 ( .A(x[2642]), .B(y[2642]), .Z(n36255) );
  AND U31109 ( .A(n26904), .B(n36255), .Z(n52043) );
  AND U31110 ( .A(n14239), .B(n52043), .Z(n14240) );
  NANDN U31111 ( .A(y[2642]), .B(x[2642]), .Z(n26902) );
  NANDN U31112 ( .A(y[2643]), .B(x[2643]), .Z(n26900) );
  NAND U31113 ( .A(n26902), .B(n26900), .Z(n54814) );
  OR U31114 ( .A(n14240), .B(n54814), .Z(n14241) );
  NAND U31115 ( .A(n54815), .B(n14241), .Z(n14242) );
  NANDN U31116 ( .A(n52042), .B(n14242), .Z(n14243) );
  NANDN U31117 ( .A(n54816), .B(n14243), .Z(n14245) );
  NANDN U31118 ( .A(y[2646]), .B(x[2646]), .Z(n14244) );
  NANDN U31119 ( .A(y[2647]), .B(x[2647]), .Z(n26897) );
  AND U31120 ( .A(n14244), .B(n26897), .Z(n52041) );
  AND U31121 ( .A(n14245), .B(n52041), .Z(n14246) );
  ANDN U31122 ( .B(y[2647]), .A(x[2647]), .Z(n36266) );
  NANDN U31123 ( .A(x[2648]), .B(y[2648]), .Z(n26895) );
  NANDN U31124 ( .A(n36266), .B(n26895), .Z(n54817) );
  OR U31125 ( .A(n14246), .B(n54817), .Z(n14247) );
  NAND U31126 ( .A(n54820), .B(n14247), .Z(n14248) );
  NANDN U31127 ( .A(n52040), .B(n14248), .Z(n14249) );
  NANDN U31128 ( .A(n54822), .B(n14249), .Z(n14251) );
  NANDN U31129 ( .A(x[2651]), .B(y[2651]), .Z(n26892) );
  XNOR U31130 ( .A(y[2652]), .B(x[2652]), .Z(n14250) );
  AND U31131 ( .A(n26892), .B(n14250), .Z(n52039) );
  AND U31132 ( .A(n14251), .B(n52039), .Z(n14252) );
  NANDN U31133 ( .A(y[2652]), .B(x[2652]), .Z(n26890) );
  NANDN U31134 ( .A(y[2653]), .B(x[2653]), .Z(n26887) );
  NAND U31135 ( .A(n26890), .B(n26887), .Z(n54823) );
  OR U31136 ( .A(n14252), .B(n54823), .Z(n14253) );
  NANDN U31137 ( .A(x[2653]), .B(y[2653]), .Z(n26889) );
  NANDN U31138 ( .A(x[2654]), .B(y[2654]), .Z(n26885) );
  AND U31139 ( .A(n26889), .B(n26885), .Z(n54824) );
  AND U31140 ( .A(n14253), .B(n54824), .Z(n14254) );
  NANDN U31141 ( .A(y[2654]), .B(x[2654]), .Z(n26886) );
  NANDN U31142 ( .A(y[2655]), .B(x[2655]), .Z(n26883) );
  NAND U31143 ( .A(n26886), .B(n26883), .Z(n52038) );
  OR U31144 ( .A(n14254), .B(n52038), .Z(n14255) );
  NAND U31145 ( .A(n52037), .B(n14255), .Z(n14256) );
  NANDN U31146 ( .A(n54825), .B(n14256), .Z(n14257) );
  NANDN U31147 ( .A(n54826), .B(n14257), .Z(n14258) );
  NANDN U31148 ( .A(y[2658]), .B(x[2658]), .Z(n36293) );
  NANDN U31149 ( .A(y[2659]), .B(x[2659]), .Z(n36300) );
  AND U31150 ( .A(n36293), .B(n36300), .Z(n54827) );
  AND U31151 ( .A(n14258), .B(n54827), .Z(n14259) );
  NANDN U31152 ( .A(x[2659]), .B(y[2659]), .Z(n26880) );
  NANDN U31153 ( .A(x[2660]), .B(y[2660]), .Z(n26879) );
  NAND U31154 ( .A(n26880), .B(n26879), .Z(n52036) );
  OR U31155 ( .A(n14259), .B(n52036), .Z(n14260) );
  NAND U31156 ( .A(n52035), .B(n14260), .Z(n14261) );
  NANDN U31157 ( .A(n54830), .B(n14261), .Z(n14262) );
  NANDN U31158 ( .A(n54831), .B(n14262), .Z(n14263) );
  NANDN U31159 ( .A(x[2663]), .B(y[2663]), .Z(n26876) );
  NANDN U31160 ( .A(x[2664]), .B(y[2664]), .Z(n26875) );
  AND U31161 ( .A(n26876), .B(n26875), .Z(n54832) );
  AND U31162 ( .A(n14263), .B(n54832), .Z(n14264) );
  NANDN U31163 ( .A(y[2664]), .B(x[2664]), .Z(n36311) );
  NANDN U31164 ( .A(y[2665]), .B(x[2665]), .Z(n36318) );
  NAND U31165 ( .A(n36311), .B(n36318), .Z(n52034) );
  OR U31166 ( .A(n14264), .B(n52034), .Z(n14265) );
  NAND U31167 ( .A(n52033), .B(n14265), .Z(n14266) );
  NANDN U31168 ( .A(n52032), .B(n14266), .Z(n14267) );
  AND U31169 ( .A(n36324), .B(n14267), .Z(n14268) );
  NANDN U31170 ( .A(n26872), .B(n14268), .Z(n14269) );
  NAND U31171 ( .A(n54833), .B(n14269), .Z(n14270) );
  NANDN U31172 ( .A(n52029), .B(n14270), .Z(n14271) );
  NAND U31173 ( .A(n52028), .B(n14271), .Z(n14272) );
  NAND U31174 ( .A(n36337), .B(n14272), .Z(n14273) );
  ANDN U31175 ( .B(y[2671]), .A(x[2671]), .Z(n54836) );
  OR U31176 ( .A(n14273), .B(n54836), .Z(n14274) );
  AND U31177 ( .A(n54839), .B(n14274), .Z(n14275) );
  OR U31178 ( .A(n54840), .B(n14275), .Z(n14276) );
  NAND U31179 ( .A(n54841), .B(n14276), .Z(n14277) );
  NANDN U31180 ( .A(n54842), .B(n14277), .Z(n14278) );
  NANDN U31181 ( .A(n54843), .B(n14278), .Z(n14279) );
  AND U31182 ( .A(n54844), .B(n14279), .Z(n14280) );
  OR U31183 ( .A(n54845), .B(n14280), .Z(n14281) );
  NAND U31184 ( .A(n54846), .B(n14281), .Z(n14282) );
  NANDN U31185 ( .A(n54847), .B(n14282), .Z(n14283) );
  NANDN U31186 ( .A(n54848), .B(n14283), .Z(n14284) );
  NANDN U31187 ( .A(y[2682]), .B(x[2682]), .Z(n26862) );
  NANDN U31188 ( .A(y[2683]), .B(x[2683]), .Z(n26861) );
  AND U31189 ( .A(n26862), .B(n26861), .Z(n54849) );
  AND U31190 ( .A(n14284), .B(n54849), .Z(n14285) );
  NANDN U31191 ( .A(x[2683]), .B(y[2683]), .Z(n36370) );
  NANDN U31192 ( .A(x[2684]), .B(y[2684]), .Z(n36377) );
  NAND U31193 ( .A(n36370), .B(n36377), .Z(n52027) );
  OR U31194 ( .A(n14285), .B(n52027), .Z(n14286) );
  NAND U31195 ( .A(n52026), .B(n14286), .Z(n14287) );
  NANDN U31196 ( .A(n52025), .B(n14287), .Z(n14288) );
  NANDN U31197 ( .A(n54851), .B(n14288), .Z(n14289) );
  AND U31198 ( .A(n54852), .B(n14289), .Z(n14290) );
  NANDN U31199 ( .A(y[2688]), .B(x[2688]), .Z(n26856) );
  NANDN U31200 ( .A(y[2689]), .B(x[2689]), .Z(n26855) );
  NAND U31201 ( .A(n26856), .B(n26855), .Z(n54853) );
  OR U31202 ( .A(n14290), .B(n54853), .Z(n14291) );
  AND U31203 ( .A(n54854), .B(n14291), .Z(n14292) );
  OR U31204 ( .A(n54855), .B(n14292), .Z(n14293) );
  NAND U31205 ( .A(n54856), .B(n14293), .Z(n14294) );
  NANDN U31206 ( .A(n54857), .B(n14294), .Z(n14295) );
  NANDN U31207 ( .A(n54858), .B(n14295), .Z(n14296) );
  AND U31208 ( .A(n54859), .B(n14296), .Z(n14297) );
  OR U31209 ( .A(n54860), .B(n14297), .Z(n14298) );
  NAND U31210 ( .A(n54861), .B(n14298), .Z(n14299) );
  NANDN U31211 ( .A(n54862), .B(n14299), .Z(n14300) );
  NANDN U31212 ( .A(n54863), .B(n14300), .Z(n14301) );
  NANDN U31213 ( .A(x[2699]), .B(y[2699]), .Z(n36414) );
  NANDN U31214 ( .A(x[2700]), .B(y[2700]), .Z(n36420) );
  AND U31215 ( .A(n36414), .B(n36420), .Z(n54864) );
  AND U31216 ( .A(n14301), .B(n54864), .Z(n14302) );
  NANDN U31217 ( .A(y[2700]), .B(x[2700]), .Z(n26840) );
  NANDN U31218 ( .A(y[2701]), .B(x[2701]), .Z(n26838) );
  AND U31219 ( .A(n26840), .B(n26838), .Z(n54865) );
  NANDN U31220 ( .A(n14302), .B(n54865), .Z(n14303) );
  NAND U31221 ( .A(n26839), .B(n14303), .Z(n14304) );
  NANDN U31222 ( .A(x[2701]), .B(y[2701]), .Z(n54867) );
  NANDN U31223 ( .A(n14304), .B(n54867), .Z(n14305) );
  AND U31224 ( .A(n54870), .B(n14305), .Z(n14306) );
  OR U31225 ( .A(n54871), .B(n14306), .Z(n14307) );
  NAND U31226 ( .A(n54872), .B(n14307), .Z(n14308) );
  NANDN U31227 ( .A(n54873), .B(n14308), .Z(n14309) );
  NANDN U31228 ( .A(n54874), .B(n14309), .Z(n14310) );
  AND U31229 ( .A(n54875), .B(n14310), .Z(n14311) );
  NANDN U31230 ( .A(y[2708]), .B(x[2708]), .Z(n26832) );
  NANDN U31231 ( .A(y[2709]), .B(x[2709]), .Z(n36447) );
  NAND U31232 ( .A(n26832), .B(n36447), .Z(n54876) );
  OR U31233 ( .A(n14311), .B(n54876), .Z(n14312) );
  AND U31234 ( .A(n52024), .B(n14312), .Z(n14313) );
  XNOR U31235 ( .A(x[2710]), .B(y[2710]), .Z(n36446) );
  NAND U31236 ( .A(n14313), .B(n36446), .Z(n14314) );
  NANDN U31237 ( .A(n54877), .B(n14314), .Z(n14315) );
  AND U31238 ( .A(n54878), .B(n14315), .Z(n14316) );
  NANDN U31239 ( .A(y[2712]), .B(x[2712]), .Z(n26830) );
  NANDN U31240 ( .A(y[2713]), .B(x[2713]), .Z(n26826) );
  AND U31241 ( .A(n26830), .B(n26826), .Z(n54879) );
  NANDN U31242 ( .A(n14316), .B(n54879), .Z(n14317) );
  NAND U31243 ( .A(n14318), .B(n14317), .Z(n14319) );
  NAND U31244 ( .A(n54882), .B(n14319), .Z(n14320) );
  NAND U31245 ( .A(n36461), .B(n14320), .Z(n14321) );
  OR U31246 ( .A(n54883), .B(n14321), .Z(n14322) );
  AND U31247 ( .A(n54888), .B(n14322), .Z(n14323) );
  OR U31248 ( .A(n54890), .B(n14323), .Z(n14324) );
  NAND U31249 ( .A(n54892), .B(n14324), .Z(n14325) );
  NANDN U31250 ( .A(n54894), .B(n14325), .Z(n14326) );
  NANDN U31251 ( .A(n54896), .B(n14326), .Z(n14327) );
  AND U31252 ( .A(n54898), .B(n14327), .Z(n14328) );
  OR U31253 ( .A(n54900), .B(n14328), .Z(n14329) );
  NAND U31254 ( .A(n54902), .B(n14329), .Z(n14330) );
  NANDN U31255 ( .A(n54904), .B(n14330), .Z(n14331) );
  NANDN U31256 ( .A(n54906), .B(n14331), .Z(n14332) );
  AND U31257 ( .A(n54908), .B(n14332), .Z(n14333) );
  OR U31258 ( .A(n54910), .B(n14333), .Z(n14334) );
  NAND U31259 ( .A(n54912), .B(n14334), .Z(n14335) );
  NANDN U31260 ( .A(n54914), .B(n14335), .Z(n14336) );
  NANDN U31261 ( .A(n54916), .B(n14336), .Z(n14337) );
  AND U31262 ( .A(n54918), .B(n14337), .Z(n14338) );
  OR U31263 ( .A(n54920), .B(n14338), .Z(n14339) );
  NAND U31264 ( .A(n54922), .B(n14339), .Z(n14340) );
  NANDN U31265 ( .A(n54924), .B(n14340), .Z(n14341) );
  NANDN U31266 ( .A(x[2735]), .B(y[2735]), .Z(n52022) );
  AND U31267 ( .A(n14341), .B(n52022), .Z(n14342) );
  NAND U31268 ( .A(n26805), .B(n14342), .Z(n14343) );
  NANDN U31269 ( .A(n26803), .B(n14343), .Z(n14344) );
  ANDN U31270 ( .B(x[2736]), .A(y[2736]), .Z(n26807) );
  OR U31271 ( .A(n14344), .B(n26807), .Z(n14345) );
  AND U31272 ( .A(n14346), .B(n14345), .Z(n14347) );
  NANDN U31273 ( .A(y[2738]), .B(x[2738]), .Z(n26804) );
  NANDN U31274 ( .A(y[2739]), .B(x[2739]), .Z(n26802) );
  NAND U31275 ( .A(n26804), .B(n26802), .Z(n52021) );
  OR U31276 ( .A(n14347), .B(n52021), .Z(n14348) );
  NAND U31277 ( .A(n54931), .B(n14348), .Z(n14349) );
  NANDN U31278 ( .A(n54932), .B(n14349), .Z(n14350) );
  AND U31279 ( .A(n54933), .B(n14350), .Z(n14353) );
  NANDN U31280 ( .A(y[2743]), .B(x[2743]), .Z(n14352) );
  NANDN U31281 ( .A(y[2742]), .B(x[2742]), .Z(n14351) );
  AND U31282 ( .A(n14352), .B(n14351), .Z(n54934) );
  NANDN U31283 ( .A(n14353), .B(n54934), .Z(n14354) );
  NANDN U31284 ( .A(n54935), .B(n14354), .Z(n14355) );
  AND U31285 ( .A(n54936), .B(n14355), .Z(n14356) );
  OR U31286 ( .A(n54937), .B(n14356), .Z(n14357) );
  NAND U31287 ( .A(n54938), .B(n14357), .Z(n14358) );
  NANDN U31288 ( .A(n54939), .B(n14358), .Z(n14359) );
  NAND U31289 ( .A(n54940), .B(n14359), .Z(n14360) );
  AND U31290 ( .A(n14361), .B(n14360), .Z(n14362) );
  OR U31291 ( .A(n54942), .B(n14362), .Z(n14363) );
  NAND U31292 ( .A(n54943), .B(n14363), .Z(n14364) );
  NANDN U31293 ( .A(n54944), .B(n14364), .Z(n14365) );
  NANDN U31294 ( .A(n54945), .B(n14365), .Z(n14366) );
  AND U31295 ( .A(n54946), .B(n14366), .Z(n14367) );
  OR U31296 ( .A(n54947), .B(n14367), .Z(n14368) );
  NAND U31297 ( .A(n54948), .B(n14368), .Z(n14369) );
  NANDN U31298 ( .A(n54949), .B(n14369), .Z(n14370) );
  NANDN U31299 ( .A(n54950), .B(n14370), .Z(n14371) );
  AND U31300 ( .A(n54951), .B(n14371), .Z(n14373) );
  NANDN U31301 ( .A(y[2760]), .B(x[2760]), .Z(n14372) );
  NANDN U31302 ( .A(y[2761]), .B(x[2761]), .Z(n36593) );
  NAND U31303 ( .A(n14372), .B(n36593), .Z(n54952) );
  OR U31304 ( .A(n14373), .B(n54952), .Z(n14374) );
  NAND U31305 ( .A(n52018), .B(n14374), .Z(n14375) );
  NANDN U31306 ( .A(n54953), .B(n14375), .Z(n14376) );
  NANDN U31307 ( .A(n54954), .B(n14376), .Z(n14377) );
  AND U31308 ( .A(n54955), .B(n14377), .Z(n14378) );
  OR U31309 ( .A(n54956), .B(n14378), .Z(n14379) );
  NAND U31310 ( .A(n54957), .B(n14379), .Z(n14380) );
  NAND U31311 ( .A(n54959), .B(n14380), .Z(n14381) );
  XNOR U31312 ( .A(x[2768]), .B(y[2768]), .Z(n36613) );
  NANDN U31313 ( .A(n14381), .B(n36613), .Z(n14382) );
  NANDN U31314 ( .A(n54964), .B(n14382), .Z(n14383) );
  AND U31315 ( .A(n54966), .B(n14383), .Z(n14384) );
  OR U31316 ( .A(n54968), .B(n14384), .Z(n14385) );
  NAND U31317 ( .A(n54970), .B(n14385), .Z(n14386) );
  NANDN U31318 ( .A(n54972), .B(n14386), .Z(n14387) );
  NANDN U31319 ( .A(n54974), .B(n14387), .Z(n14388) );
  AND U31320 ( .A(n54976), .B(n14388), .Z(n14390) );
  XNOR U31321 ( .A(x[2776]), .B(y[2776]), .Z(n26773) );
  NANDN U31322 ( .A(x[2775]), .B(y[2775]), .Z(n54978) );
  AND U31323 ( .A(n26773), .B(n54978), .Z(n14389) );
  NANDN U31324 ( .A(n14390), .B(n14389), .Z(n14391) );
  NAND U31325 ( .A(n54982), .B(n14391), .Z(n14392) );
  NAND U31326 ( .A(n26771), .B(n14392), .Z(n14393) );
  OR U31327 ( .A(n54984), .B(n14393), .Z(n14394) );
  AND U31328 ( .A(n54988), .B(n14394), .Z(n14395) );
  OR U31329 ( .A(n54990), .B(n14395), .Z(n14396) );
  NAND U31330 ( .A(n54992), .B(n14396), .Z(n14397) );
  NANDN U31331 ( .A(n54994), .B(n14397), .Z(n14398) );
  NANDN U31332 ( .A(n54996), .B(n14398), .Z(n14399) );
  AND U31333 ( .A(n54998), .B(n14399), .Z(n14400) );
  OR U31334 ( .A(n54999), .B(n14400), .Z(n14401) );
  NAND U31335 ( .A(n55001), .B(n14401), .Z(n14402) );
  NANDN U31336 ( .A(n55002), .B(n14402), .Z(n14403) );
  NANDN U31337 ( .A(n52017), .B(n14403), .Z(n14404) );
  NANDN U31338 ( .A(y[2788]), .B(x[2788]), .Z(n36671) );
  NANDN U31339 ( .A(y[2789]), .B(x[2789]), .Z(n36677) );
  AND U31340 ( .A(n36671), .B(n36677), .Z(n52016) );
  AND U31341 ( .A(n14404), .B(n52016), .Z(n14405) );
  NOR U31342 ( .A(n26762), .B(n14405), .Z(n14406) );
  XNOR U31343 ( .A(x[2790]), .B(y[2790]), .Z(n36678) );
  NAND U31344 ( .A(n14406), .B(n36678), .Z(n14407) );
  NANDN U31345 ( .A(n55004), .B(n14407), .Z(n14408) );
  AND U31346 ( .A(n55005), .B(n14408), .Z(n14409) );
  OR U31347 ( .A(n55006), .B(n14409), .Z(n14410) );
  NAND U31348 ( .A(n55007), .B(n14410), .Z(n14411) );
  NANDN U31349 ( .A(n55008), .B(n14411), .Z(n14412) );
  NANDN U31350 ( .A(n55009), .B(n14412), .Z(n14415) );
  NANDN U31351 ( .A(y[2797]), .B(x[2797]), .Z(n14414) );
  NANDN U31352 ( .A(y[2796]), .B(x[2796]), .Z(n14413) );
  NAND U31353 ( .A(n14414), .B(n14413), .Z(n55010) );
  ANDN U31354 ( .B(n14415), .A(n55010), .Z(n14416) );
  OR U31355 ( .A(n55011), .B(n14416), .Z(n14417) );
  NAND U31356 ( .A(n55012), .B(n14417), .Z(n14418) );
  NANDN U31357 ( .A(n55013), .B(n14418), .Z(n14419) );
  NANDN U31358 ( .A(n55015), .B(n14419), .Z(n14420) );
  AND U31359 ( .A(n55016), .B(n14420), .Z(n14421) );
  NANDN U31360 ( .A(y[2802]), .B(x[2802]), .Z(n26751) );
  NANDN U31361 ( .A(y[2803]), .B(x[2803]), .Z(n26750) );
  NAND U31362 ( .A(n26751), .B(n26750), .Z(n55017) );
  OR U31363 ( .A(n14421), .B(n55017), .Z(n14422) );
  NAND U31364 ( .A(n52014), .B(n14422), .Z(n14423) );
  NANDN U31365 ( .A(n55018), .B(n14423), .Z(n14424) );
  NANDN U31366 ( .A(n55019), .B(n14424), .Z(n14425) );
  AND U31367 ( .A(n55020), .B(n14425), .Z(n14426) );
  OR U31368 ( .A(n55021), .B(n14426), .Z(n14427) );
  NAND U31369 ( .A(n55022), .B(n14427), .Z(n14428) );
  NANDN U31370 ( .A(n55023), .B(n14428), .Z(n14429) );
  NANDN U31371 ( .A(n55024), .B(n14429), .Z(n14430) );
  AND U31372 ( .A(n55025), .B(n14430), .Z(n14431) );
  OR U31373 ( .A(n55026), .B(n14431), .Z(n14432) );
  NAND U31374 ( .A(n55027), .B(n14432), .Z(n14433) );
  NANDN U31375 ( .A(n55028), .B(n14433), .Z(n14434) );
  AND U31376 ( .A(n36755), .B(n14434), .Z(n14435) );
  NAND U31377 ( .A(n55030), .B(n14435), .Z(n14436) );
  NANDN U31378 ( .A(n55032), .B(n14436), .Z(n14437) );
  AND U31379 ( .A(n26738), .B(n14437), .Z(n14438) );
  NANDN U31380 ( .A(n26739), .B(n14438), .Z(n14439) );
  NAND U31381 ( .A(n52013), .B(n14439), .Z(n14440) );
  NANDN U31382 ( .A(n55035), .B(n14440), .Z(n14441) );
  NAND U31383 ( .A(n55036), .B(n14441), .Z(n14442) );
  NAND U31384 ( .A(n36769), .B(n14442), .Z(n14443) );
  ANDN U31385 ( .B(y[2821]), .A(x[2821]), .Z(n26732) );
  OR U31386 ( .A(n14443), .B(n26732), .Z(n14444) );
  AND U31387 ( .A(n55038), .B(n14444), .Z(n14445) );
  OR U31388 ( .A(n55039), .B(n14445), .Z(n14446) );
  NAND U31389 ( .A(n55040), .B(n14446), .Z(n14447) );
  NANDN U31390 ( .A(n55041), .B(n14447), .Z(n14448) );
  NANDN U31391 ( .A(n55042), .B(n14448), .Z(n14449) );
  AND U31392 ( .A(n55043), .B(n14449), .Z(n14450) );
  OR U31393 ( .A(n55044), .B(n14450), .Z(n14451) );
  NAND U31394 ( .A(n55045), .B(n14451), .Z(n14452) );
  NANDN U31395 ( .A(n55047), .B(n14452), .Z(n14453) );
  NANDN U31396 ( .A(n55048), .B(n14453), .Z(n14454) );
  AND U31397 ( .A(n55049), .B(n14454), .Z(n14455) );
  OR U31398 ( .A(n55050), .B(n14455), .Z(n14456) );
  NAND U31399 ( .A(n55051), .B(n14456), .Z(n14457) );
  NAND U31400 ( .A(n55052), .B(n14457), .Z(n14458) );
  XNOR U31401 ( .A(x[2836]), .B(y[2836]), .Z(n26720) );
  NANDN U31402 ( .A(n14458), .B(n26720), .Z(n14459) );
  NAND U31403 ( .A(n52011), .B(n14459), .Z(n14460) );
  NANDN U31404 ( .A(n55054), .B(n14460), .Z(n14462) );
  NANDN U31405 ( .A(y[2838]), .B(x[2838]), .Z(n14461) );
  NANDN U31406 ( .A(y[2839]), .B(x[2839]), .Z(n26715) );
  AND U31407 ( .A(n14461), .B(n26715), .Z(n55055) );
  AND U31408 ( .A(n14462), .B(n55055), .Z(n14463) );
  NANDN U31409 ( .A(x[2839]), .B(y[2839]), .Z(n36818) );
  NANDN U31410 ( .A(x[2840]), .B(y[2840]), .Z(n26713) );
  NAND U31411 ( .A(n36818), .B(n26713), .Z(n52010) );
  OR U31412 ( .A(n14463), .B(n52010), .Z(n14464) );
  NAND U31413 ( .A(n52009), .B(n14464), .Z(n14465) );
  NANDN U31414 ( .A(n55056), .B(n14465), .Z(n14466) );
  AND U31415 ( .A(n55057), .B(n14466), .Z(n14468) );
  XNOR U31416 ( .A(x[2844]), .B(y[2844]), .Z(n14467) );
  ANDN U31417 ( .B(y[2843]), .A(x[2843]), .Z(n36828) );
  ANDN U31418 ( .B(n14467), .A(n36828), .Z(n55058) );
  NANDN U31419 ( .A(n14468), .B(n55058), .Z(n14469) );
  NANDN U31420 ( .A(n55060), .B(n14469), .Z(n14470) );
  AND U31421 ( .A(n55061), .B(n14470), .Z(n14471) );
  NANDN U31422 ( .A(y[2846]), .B(x[2846]), .Z(n26706) );
  NANDN U31423 ( .A(y[2847]), .B(x[2847]), .Z(n36844) );
  NAND U31424 ( .A(n26706), .B(n36844), .Z(n52008) );
  OR U31425 ( .A(n14471), .B(n52008), .Z(n14472) );
  NAND U31426 ( .A(n52007), .B(n14472), .Z(n14473) );
  NANDN U31427 ( .A(n55062), .B(n14473), .Z(n14474) );
  NANDN U31428 ( .A(n55063), .B(n14474), .Z(n14475) );
  NANDN U31429 ( .A(y[2850]), .B(x[2850]), .Z(n36849) );
  NANDN U31430 ( .A(y[2851]), .B(x[2851]), .Z(n36856) );
  AND U31431 ( .A(n36849), .B(n36856), .Z(n55064) );
  AND U31432 ( .A(n14475), .B(n55064), .Z(n14476) );
  NANDN U31433 ( .A(x[2851]), .B(y[2851]), .Z(n26702) );
  NANDN U31434 ( .A(x[2852]), .B(y[2852]), .Z(n26701) );
  AND U31435 ( .A(n26702), .B(n26701), .Z(n55065) );
  NANDN U31436 ( .A(n14476), .B(n55065), .Z(n14477) );
  NANDN U31437 ( .A(n55066), .B(n14477), .Z(n14478) );
  NANDN U31438 ( .A(x[2853]), .B(y[2853]), .Z(n26700) );
  NANDN U31439 ( .A(x[2854]), .B(y[2854]), .Z(n26699) );
  AND U31440 ( .A(n26700), .B(n26699), .Z(n52006) );
  AND U31441 ( .A(n14478), .B(n52006), .Z(n14479) );
  NANDN U31442 ( .A(y[2854]), .B(x[2854]), .Z(n36861) );
  NANDN U31443 ( .A(y[2855]), .B(x[2855]), .Z(n36870) );
  NAND U31444 ( .A(n36861), .B(n36870), .Z(n55067) );
  OR U31445 ( .A(n14479), .B(n55067), .Z(n14480) );
  AND U31446 ( .A(n55068), .B(n14480), .Z(n14481) );
  NANDN U31447 ( .A(y[2856]), .B(x[2856]), .Z(n36868) );
  NANDN U31448 ( .A(y[2857]), .B(x[2857]), .Z(n36877) );
  NAND U31449 ( .A(n36868), .B(n36877), .Z(n52005) );
  OR U31450 ( .A(n14481), .B(n52005), .Z(n14482) );
  NAND U31451 ( .A(n55071), .B(n14482), .Z(n14483) );
  NANDN U31452 ( .A(n55072), .B(n14483), .Z(n14484) );
  NANDN U31453 ( .A(n55073), .B(n14484), .Z(n14485) );
  NANDN U31454 ( .A(y[2860]), .B(x[2860]), .Z(n36882) );
  NANDN U31455 ( .A(y[2861]), .B(x[2861]), .Z(n36889) );
  AND U31456 ( .A(n36882), .B(n36889), .Z(n55074) );
  AND U31457 ( .A(n14485), .B(n55074), .Z(n14486) );
  NANDN U31458 ( .A(x[2861]), .B(y[2861]), .Z(n26694) );
  NANDN U31459 ( .A(x[2862]), .B(y[2862]), .Z(n36892) );
  NAND U31460 ( .A(n26694), .B(n36892), .Z(n52004) );
  OR U31461 ( .A(n14486), .B(n52004), .Z(n14487) );
  NAND U31462 ( .A(n52003), .B(n14487), .Z(n14488) );
  NANDN U31463 ( .A(n55075), .B(n14488), .Z(n14489) );
  NANDN U31464 ( .A(n55076), .B(n14489), .Z(n14490) );
  NANDN U31465 ( .A(x[2865]), .B(y[2865]), .Z(n36897) );
  NANDN U31466 ( .A(x[2866]), .B(y[2866]), .Z(n36904) );
  AND U31467 ( .A(n36897), .B(n36904), .Z(n55077) );
  AND U31468 ( .A(n14490), .B(n55077), .Z(n14491) );
  NANDN U31469 ( .A(y[2866]), .B(x[2866]), .Z(n26690) );
  NANDN U31470 ( .A(y[2867]), .B(x[2867]), .Z(n26689) );
  NAND U31471 ( .A(n26690), .B(n26689), .Z(n52002) );
  OR U31472 ( .A(n14491), .B(n52002), .Z(n14492) );
  NAND U31473 ( .A(n52001), .B(n14492), .Z(n14493) );
  NANDN U31474 ( .A(n55079), .B(n14493), .Z(n14494) );
  NANDN U31475 ( .A(n55080), .B(n14494), .Z(n14495) );
  NANDN U31476 ( .A(y[2870]), .B(x[2870]), .Z(n26686) );
  NANDN U31477 ( .A(y[2871]), .B(x[2871]), .Z(n26685) );
  AND U31478 ( .A(n26686), .B(n26685), .Z(n55082) );
  AND U31479 ( .A(n14495), .B(n55082), .Z(n14496) );
  NANDN U31480 ( .A(x[2871]), .B(y[2871]), .Z(n36915) );
  NANDN U31481 ( .A(x[2872]), .B(y[2872]), .Z(n26683) );
  NAND U31482 ( .A(n36915), .B(n26683), .Z(n52000) );
  OR U31483 ( .A(n14496), .B(n52000), .Z(n14497) );
  NAND U31484 ( .A(n51999), .B(n14497), .Z(n14498) );
  NANDN U31485 ( .A(n55083), .B(n14498), .Z(n14499) );
  NANDN U31486 ( .A(n55084), .B(n14499), .Z(n14500) );
  NANDN U31487 ( .A(x[2875]), .B(y[2875]), .Z(n36926) );
  NANDN U31488 ( .A(x[2876]), .B(y[2876]), .Z(n26677) );
  AND U31489 ( .A(n36926), .B(n26677), .Z(n55085) );
  AND U31490 ( .A(n14500), .B(n55085), .Z(n14501) );
  NANDN U31491 ( .A(y[2876]), .B(x[2876]), .Z(n26678) );
  NANDN U31492 ( .A(y[2877]), .B(x[2877]), .Z(n26675) );
  NAND U31493 ( .A(n26678), .B(n26675), .Z(n51998) );
  OR U31494 ( .A(n14501), .B(n51998), .Z(n14502) );
  NAND U31495 ( .A(n51997), .B(n14502), .Z(n14503) );
  NANDN U31496 ( .A(n55086), .B(n14503), .Z(n14504) );
  AND U31497 ( .A(n55087), .B(n14504), .Z(n14505) );
  OR U31498 ( .A(n55088), .B(n14505), .Z(n14506) );
  NAND U31499 ( .A(n55090), .B(n14506), .Z(n14507) );
  NANDN U31500 ( .A(n55091), .B(n14507), .Z(n14508) );
  NAND U31501 ( .A(n51996), .B(n14508), .Z(n14509) );
  NANDN U31502 ( .A(n55092), .B(n14509), .Z(n14510) );
  NANDN U31503 ( .A(x[2885]), .B(y[2885]), .Z(n36954) );
  NANDN U31504 ( .A(x[2886]), .B(y[2886]), .Z(n26665) );
  AND U31505 ( .A(n36954), .B(n26665), .Z(n55093) );
  AND U31506 ( .A(n14510), .B(n55093), .Z(n14511) );
  NANDN U31507 ( .A(y[2886]), .B(x[2886]), .Z(n26666) );
  NANDN U31508 ( .A(y[2887]), .B(x[2887]), .Z(n26664) );
  NAND U31509 ( .A(n26666), .B(n26664), .Z(n51995) );
  OR U31510 ( .A(n14511), .B(n51995), .Z(n14512) );
  NANDN U31511 ( .A(x[2887]), .B(y[2887]), .Z(n51994) );
  AND U31512 ( .A(n14512), .B(n51994), .Z(n14515) );
  NANDN U31513 ( .A(x[2888]), .B(y[2888]), .Z(n14513) );
  AND U31514 ( .A(n14514), .B(n14513), .Z(n51993) );
  AND U31515 ( .A(n14515), .B(n51993), .Z(n14516) );
  OR U31516 ( .A(n14517), .B(n14516), .Z(n14518) );
  NANDN U31517 ( .A(x[2890]), .B(y[2890]), .Z(n55096) );
  AND U31518 ( .A(n14518), .B(n55096), .Z(n14519) );
  ANDN U31519 ( .B(x[2890]), .A(y[2890]), .Z(n36965) );
  NANDN U31520 ( .A(y[2891]), .B(x[2891]), .Z(n26662) );
  NANDN U31521 ( .A(n36965), .B(n26662), .Z(n55097) );
  OR U31522 ( .A(n14519), .B(n55097), .Z(n14520) );
  NAND U31523 ( .A(n55098), .B(n14520), .Z(n14521) );
  NANDN U31524 ( .A(n55101), .B(n14521), .Z(n14522) );
  NANDN U31525 ( .A(n55102), .B(n14522), .Z(n14523) );
  AND U31526 ( .A(n55103), .B(n14523), .Z(n14524) );
  OR U31527 ( .A(n55104), .B(n14524), .Z(n14525) );
  NAND U31528 ( .A(n51992), .B(n14525), .Z(n14526) );
  NANDN U31529 ( .A(n55105), .B(n14526), .Z(n14527) );
  NANDN U31530 ( .A(n55106), .B(n14527), .Z(n14528) );
  AND U31531 ( .A(n55107), .B(n14528), .Z(n14529) );
  OR U31532 ( .A(n55108), .B(n14529), .Z(n14530) );
  NAND U31533 ( .A(n51991), .B(n14530), .Z(n14531) );
  NANDN U31534 ( .A(n55109), .B(n14531), .Z(n14532) );
  NANDN U31535 ( .A(n55110), .B(n14532), .Z(n14533) );
  AND U31536 ( .A(n55111), .B(n14533), .Z(n14534) );
  OR U31537 ( .A(n55112), .B(n14534), .Z(n14535) );
  NAND U31538 ( .A(n51990), .B(n14535), .Z(n14536) );
  NANDN U31539 ( .A(n55114), .B(n14536), .Z(n14537) );
  NANDN U31540 ( .A(n55115), .B(n14537), .Z(n14538) );
  AND U31541 ( .A(n55116), .B(n14538), .Z(n14539) );
  OR U31542 ( .A(n55117), .B(n14539), .Z(n14540) );
  NAND U31543 ( .A(n55118), .B(n14540), .Z(n14541) );
  NANDN U31544 ( .A(n55119), .B(n14541), .Z(n14542) );
  NANDN U31545 ( .A(n55120), .B(n14542), .Z(n14543) );
  AND U31546 ( .A(n55121), .B(n14543), .Z(n14544) );
  OR U31547 ( .A(n55122), .B(n14544), .Z(n14545) );
  NAND U31548 ( .A(n55123), .B(n14545), .Z(n14546) );
  NANDN U31549 ( .A(n55124), .B(n14546), .Z(n14547) );
  NANDN U31550 ( .A(n55125), .B(n14547), .Z(n14548) );
  AND U31551 ( .A(n55126), .B(n14548), .Z(n14549) );
  OR U31552 ( .A(n55127), .B(n14549), .Z(n14550) );
  NAND U31553 ( .A(n55128), .B(n14550), .Z(n14551) );
  NANDN U31554 ( .A(n55129), .B(n14551), .Z(n14552) );
  NANDN U31555 ( .A(n55131), .B(n14552), .Z(n14553) );
  AND U31556 ( .A(n55132), .B(n14553), .Z(n14554) );
  OR U31557 ( .A(n55133), .B(n14554), .Z(n14555) );
  NAND U31558 ( .A(n55134), .B(n14555), .Z(n14556) );
  NANDN U31559 ( .A(n55135), .B(n14556), .Z(n14557) );
  NANDN U31560 ( .A(n55136), .B(n14557), .Z(n14558) );
  AND U31561 ( .A(n55137), .B(n14558), .Z(n14559) );
  OR U31562 ( .A(n55138), .B(n14559), .Z(n14560) );
  NAND U31563 ( .A(n55139), .B(n14560), .Z(n14561) );
  NANDN U31564 ( .A(n55140), .B(n14561), .Z(n14562) );
  NANDN U31565 ( .A(n55141), .B(n14562), .Z(n14563) );
  AND U31566 ( .A(n55142), .B(n14563), .Z(n14564) );
  OR U31567 ( .A(n55143), .B(n14564), .Z(n14565) );
  NAND U31568 ( .A(n55144), .B(n14565), .Z(n14566) );
  NAND U31569 ( .A(n55145), .B(n14566), .Z(n14567) );
  XNOR U31570 ( .A(x[2938]), .B(y[2938]), .Z(n37102) );
  NANDN U31571 ( .A(n14567), .B(n37102), .Z(n14568) );
  NANDN U31572 ( .A(n55147), .B(n14568), .Z(n14569) );
  AND U31573 ( .A(n55148), .B(n14569), .Z(n14570) );
  OR U31574 ( .A(n55149), .B(n14570), .Z(n14571) );
  NAND U31575 ( .A(n55151), .B(n14571), .Z(n14572) );
  NANDN U31576 ( .A(n55152), .B(n14572), .Z(n14573) );
  NANDN U31577 ( .A(n55153), .B(n14573), .Z(n14574) );
  AND U31578 ( .A(n55154), .B(n14574), .Z(n14575) );
  NANDN U31579 ( .A(x[2945]), .B(y[2945]), .Z(n26603) );
  NANDN U31580 ( .A(x[2946]), .B(y[2946]), .Z(n26602) );
  AND U31581 ( .A(n26603), .B(n26602), .Z(n55155) );
  NANDN U31582 ( .A(n14575), .B(n55155), .Z(n14576) );
  NANDN U31583 ( .A(n51989), .B(n14576), .Z(n14577) );
  XNOR U31584 ( .A(y[2948]), .B(x[2948]), .Z(n37130) );
  NANDN U31585 ( .A(x[2947]), .B(y[2947]), .Z(n26601) );
  AND U31586 ( .A(n37130), .B(n26601), .Z(n51988) );
  AND U31587 ( .A(n14577), .B(n51988), .Z(n14579) );
  NANDN U31588 ( .A(y[2948]), .B(x[2948]), .Z(n14578) );
  NANDN U31589 ( .A(y[2949]), .B(x[2949]), .Z(n37137) );
  NAND U31590 ( .A(n14578), .B(n37137), .Z(n55156) );
  OR U31591 ( .A(n14579), .B(n55156), .Z(n14580) );
  AND U31592 ( .A(n55157), .B(n14580), .Z(n14581) );
  NANDN U31593 ( .A(y[2950]), .B(x[2950]), .Z(n37136) );
  NANDN U31594 ( .A(y[2951]), .B(x[2951]), .Z(n26595) );
  AND U31595 ( .A(n37136), .B(n26595), .Z(n55158) );
  NANDN U31596 ( .A(n14581), .B(n55158), .Z(n14582) );
  NANDN U31597 ( .A(n55159), .B(n14582), .Z(n14583) );
  AND U31598 ( .A(n55160), .B(n14583), .Z(n14584) );
  NANDN U31599 ( .A(x[2954]), .B(y[2954]), .Z(n55161) );
  NANDN U31600 ( .A(n14584), .B(n55161), .Z(n14585) );
  AND U31601 ( .A(n55162), .B(n14585), .Z(n14586) );
  OR U31602 ( .A(n55163), .B(n14586), .Z(n14587) );
  NAND U31603 ( .A(n55164), .B(n14587), .Z(n14588) );
  NANDN U31604 ( .A(n55165), .B(n14588), .Z(n14589) );
  NANDN U31605 ( .A(n55166), .B(n14589), .Z(n14590) );
  NANDN U31606 ( .A(x[2959]), .B(y[2959]), .Z(n37156) );
  NANDN U31607 ( .A(x[2960]), .B(y[2960]), .Z(n37163) );
  AND U31608 ( .A(n37156), .B(n37163), .Z(n55169) );
  AND U31609 ( .A(n14590), .B(n55169), .Z(n14591) );
  NANDN U31610 ( .A(y[2960]), .B(x[2960]), .Z(n26584) );
  NANDN U31611 ( .A(y[2961]), .B(x[2961]), .Z(n26583) );
  NAND U31612 ( .A(n26584), .B(n26583), .Z(n51987) );
  OR U31613 ( .A(n14591), .B(n51987), .Z(n14592) );
  NAND U31614 ( .A(n51986), .B(n14592), .Z(n14593) );
  NANDN U31615 ( .A(n51985), .B(n14593), .Z(n14595) );
  XNOR U31616 ( .A(x[2964]), .B(y[2964]), .Z(n37171) );
  NANDN U31617 ( .A(x[2963]), .B(y[2963]), .Z(n55171) );
  AND U31618 ( .A(n37171), .B(n55171), .Z(n14594) );
  NAND U31619 ( .A(n14595), .B(n14594), .Z(n14597) );
  NANDN U31620 ( .A(y[2964]), .B(x[2964]), .Z(n14596) );
  NANDN U31621 ( .A(y[2965]), .B(x[2965]), .Z(n37177) );
  AND U31622 ( .A(n14596), .B(n37177), .Z(n51984) );
  AND U31623 ( .A(n14597), .B(n51984), .Z(n14598) );
  NANDN U31624 ( .A(x[2965]), .B(y[2965]), .Z(n26581) );
  NANDN U31625 ( .A(x[2966]), .B(y[2966]), .Z(n26580) );
  NAND U31626 ( .A(n26581), .B(n26580), .Z(n55173) );
  OR U31627 ( .A(n14598), .B(n55173), .Z(n14599) );
  NAND U31628 ( .A(n55174), .B(n14599), .Z(n14600) );
  NANDN U31629 ( .A(n51983), .B(n14600), .Z(n14601) );
  NANDN U31630 ( .A(y[2968]), .B(x[2968]), .Z(n37182) );
  NANDN U31631 ( .A(y[2969]), .B(x[2969]), .Z(n37188) );
  AND U31632 ( .A(n37182), .B(n37188), .Z(n51982) );
  AND U31633 ( .A(n14601), .B(n51982), .Z(n14602) );
  XNOR U31634 ( .A(x[2970]), .B(y[2970]), .Z(n37189) );
  NANDN U31635 ( .A(n14602), .B(n37189), .Z(n14603) );
  ANDN U31636 ( .B(y[2969]), .A(x[2969]), .Z(n26577) );
  OR U31637 ( .A(n14603), .B(n26577), .Z(n14604) );
  AND U31638 ( .A(n55179), .B(n14604), .Z(n14605) );
  OR U31639 ( .A(n55180), .B(n14605), .Z(n14606) );
  NAND U31640 ( .A(n55181), .B(n14606), .Z(n14607) );
  NANDN U31641 ( .A(n55182), .B(n14607), .Z(n14608) );
  NANDN U31642 ( .A(n55183), .B(n14608), .Z(n14609) );
  AND U31643 ( .A(n55184), .B(n14609), .Z(n14610) );
  OR U31644 ( .A(n55185), .B(n14610), .Z(n14611) );
  NAND U31645 ( .A(n55186), .B(n14611), .Z(n14612) );
  NANDN U31646 ( .A(n55187), .B(n14612), .Z(n14613) );
  NANDN U31647 ( .A(n55188), .B(n14613), .Z(n14614) );
  AND U31648 ( .A(n55189), .B(n14614), .Z(n14615) );
  NANDN U31649 ( .A(x[2981]), .B(y[2981]), .Z(n26562) );
  NANDN U31650 ( .A(x[2982]), .B(y[2982]), .Z(n26558) );
  NAND U31651 ( .A(n26562), .B(n26558), .Z(n55190) );
  OR U31652 ( .A(n14615), .B(n55190), .Z(n14616) );
  NAND U31653 ( .A(n51981), .B(n14616), .Z(n14617) );
  NANDN U31654 ( .A(n55191), .B(n14617), .Z(n14618) );
  NANDN U31655 ( .A(n55192), .B(n14618), .Z(n14619) );
  AND U31656 ( .A(n55193), .B(n14619), .Z(n14620) );
  OR U31657 ( .A(n55195), .B(n14620), .Z(n14621) );
  NAND U31658 ( .A(n55196), .B(n14621), .Z(n14622) );
  NANDN U31659 ( .A(n55197), .B(n14622), .Z(n14623) );
  NANDN U31660 ( .A(n55198), .B(n14623), .Z(n14624) );
  AND U31661 ( .A(n55199), .B(n14624), .Z(n14625) );
  NANDN U31662 ( .A(x[2991]), .B(y[2991]), .Z(n26548) );
  NANDN U31663 ( .A(x[2992]), .B(y[2992]), .Z(n26547) );
  AND U31664 ( .A(n26548), .B(n26547), .Z(n55200) );
  NANDN U31665 ( .A(n14625), .B(n55200), .Z(n14626) );
  NANDN U31666 ( .A(n51980), .B(n14626), .Z(n14627) );
  XNOR U31667 ( .A(y[2994]), .B(x[2994]), .Z(n37253) );
  NANDN U31668 ( .A(x[2993]), .B(y[2993]), .Z(n26546) );
  AND U31669 ( .A(n37253), .B(n26546), .Z(n51979) );
  AND U31670 ( .A(n14627), .B(n51979), .Z(n14629) );
  NANDN U31671 ( .A(y[2994]), .B(x[2994]), .Z(n14628) );
  NANDN U31672 ( .A(y[2995]), .B(x[2995]), .Z(n37259) );
  NAND U31673 ( .A(n14628), .B(n37259), .Z(n55201) );
  OR U31674 ( .A(n14629), .B(n55201), .Z(n14630) );
  AND U31675 ( .A(n55202), .B(n14630), .Z(n14631) );
  OR U31676 ( .A(n55203), .B(n14631), .Z(n14632) );
  NAND U31677 ( .A(n55204), .B(n14632), .Z(n14633) );
  NANDN U31678 ( .A(n55205), .B(n14633), .Z(n14634) );
  NANDN U31679 ( .A(n55206), .B(n14634), .Z(n14635) );
  AND U31680 ( .A(n55207), .B(n14635), .Z(n14636) );
  OR U31681 ( .A(n55208), .B(n14636), .Z(n14637) );
  NAND U31682 ( .A(n55209), .B(n14637), .Z(n14638) );
  NANDN U31683 ( .A(n55211), .B(n14638), .Z(n14639) );
  NANDN U31684 ( .A(n55212), .B(n14639), .Z(n14640) );
  NANDN U31685 ( .A(x[3005]), .B(y[3005]), .Z(n26534) );
  NANDN U31686 ( .A(x[3006]), .B(y[3006]), .Z(n26533) );
  AND U31687 ( .A(n26534), .B(n26533), .Z(n55214) );
  AND U31688 ( .A(n14640), .B(n55214), .Z(n14641) );
  NANDN U31689 ( .A(y[3006]), .B(x[3006]), .Z(n37288) );
  NANDN U31690 ( .A(y[3007]), .B(x[3007]), .Z(n37294) );
  AND U31691 ( .A(n37288), .B(n37294), .Z(n55215) );
  NANDN U31692 ( .A(n14641), .B(n55215), .Z(n14642) );
  NAND U31693 ( .A(n37295), .B(n14642), .Z(n14643) );
  NANDN U31694 ( .A(x[3007]), .B(y[3007]), .Z(n55216) );
  NANDN U31695 ( .A(n14643), .B(n55216), .Z(n14644) );
  AND U31696 ( .A(n55218), .B(n14644), .Z(n14645) );
  OR U31697 ( .A(n55219), .B(n14645), .Z(n14646) );
  NAND U31698 ( .A(n55220), .B(n14646), .Z(n14647) );
  NANDN U31699 ( .A(n55221), .B(n14647), .Z(n14648) );
  NAND U31700 ( .A(n55222), .B(n14648), .Z(n14649) );
  AND U31701 ( .A(n14650), .B(n14649), .Z(n14651) );
  OR U31702 ( .A(n55223), .B(n14651), .Z(n14652) );
  NAND U31703 ( .A(n55224), .B(n14652), .Z(n14653) );
  NANDN U31704 ( .A(n55225), .B(n14653), .Z(n14654) );
  NANDN U31705 ( .A(n55226), .B(n14654), .Z(n14655) );
  AND U31706 ( .A(n55227), .B(n14655), .Z(n14656) );
  OR U31707 ( .A(n55229), .B(n14656), .Z(n14657) );
  NAND U31708 ( .A(n55231), .B(n14657), .Z(n14658) );
  NANDN U31709 ( .A(n55233), .B(n14658), .Z(n14659) );
  NANDN U31710 ( .A(n55235), .B(n14659), .Z(n14660) );
  AND U31711 ( .A(n55237), .B(n14660), .Z(n14661) );
  OR U31712 ( .A(n55239), .B(n14661), .Z(n14662) );
  NAND U31713 ( .A(n55241), .B(n14662), .Z(n14663) );
  NANDN U31714 ( .A(n55243), .B(n14663), .Z(n14664) );
  NANDN U31715 ( .A(n55245), .B(n14664), .Z(n14665) );
  AND U31716 ( .A(n55247), .B(n14665), .Z(n14666) );
  OR U31717 ( .A(n55249), .B(n14666), .Z(n14667) );
  NAND U31718 ( .A(n55251), .B(n14667), .Z(n14668) );
  NANDN U31719 ( .A(n55253), .B(n14668), .Z(n14669) );
  NANDN U31720 ( .A(n55255), .B(n14669), .Z(n14670) );
  AND U31721 ( .A(n55257), .B(n14670), .Z(n14671) );
  OR U31722 ( .A(n55259), .B(n14671), .Z(n14672) );
  NAND U31723 ( .A(n55261), .B(n14672), .Z(n14673) );
  NANDN U31724 ( .A(n55263), .B(n14673), .Z(n14674) );
  NANDN U31725 ( .A(n55265), .B(n14674), .Z(n14675) );
  AND U31726 ( .A(n55267), .B(n14675), .Z(n14677) );
  NANDN U31727 ( .A(x[3040]), .B(y[3040]), .Z(n55273) );
  NANDN U31728 ( .A(x[3039]), .B(y[3039]), .Z(n55268) );
  AND U31729 ( .A(n55273), .B(n55268), .Z(n14676) );
  NANDN U31730 ( .A(n14677), .B(n14676), .Z(n14678) );
  NAND U31731 ( .A(n55271), .B(n14678), .Z(n14679) );
  AND U31732 ( .A(n55274), .B(n14679), .Z(n14680) );
  ANDN U31733 ( .B(x[3043]), .A(y[3043]), .Z(n37407) );
  NANDN U31734 ( .A(y[3042]), .B(x[3042]), .Z(n26509) );
  NANDN U31735 ( .A(n37407), .B(n26509), .Z(n55276) );
  OR U31736 ( .A(n14680), .B(n55276), .Z(n14683) );
  NANDN U31737 ( .A(x[3044]), .B(y[3044]), .Z(n14682) );
  NANDN U31738 ( .A(x[3043]), .B(y[3043]), .Z(n14681) );
  AND U31739 ( .A(n14682), .B(n14681), .Z(n55277) );
  AND U31740 ( .A(n14683), .B(n55277), .Z(n14684) );
  ANDN U31741 ( .B(x[3044]), .A(y[3044]), .Z(n37410) );
  ANDN U31742 ( .B(x[3045]), .A(y[3045]), .Z(n37415) );
  OR U31743 ( .A(n37410), .B(n37415), .Z(n55278) );
  OR U31744 ( .A(n14684), .B(n55278), .Z(n14685) );
  AND U31745 ( .A(n55279), .B(n14685), .Z(n14687) );
  XNOR U31746 ( .A(x[3046]), .B(y[3046]), .Z(n14686) );
  NAND U31747 ( .A(n14687), .B(n14686), .Z(n14688) );
  NANDN U31748 ( .A(n55281), .B(n14688), .Z(n14689) );
  AND U31749 ( .A(n55282), .B(n14689), .Z(n14690) );
  OR U31750 ( .A(n55283), .B(n14690), .Z(n14691) );
  AND U31751 ( .A(n14692), .B(n14691), .Z(n14694) );
  NANDN U31752 ( .A(y[3050]), .B(x[3050]), .Z(n14693) );
  NANDN U31753 ( .A(y[3051]), .B(x[3051]), .Z(n26503) );
  NAND U31754 ( .A(n14693), .B(n26503), .Z(n55286) );
  OR U31755 ( .A(n14694), .B(n55286), .Z(n14695) );
  NAND U31756 ( .A(n55287), .B(n14695), .Z(n14696) );
  NANDN U31757 ( .A(n51976), .B(n14696), .Z(n14697) );
  NANDN U31758 ( .A(n55290), .B(n14697), .Z(n14698) );
  NANDN U31759 ( .A(y[3054]), .B(x[3054]), .Z(n26500) );
  NANDN U31760 ( .A(y[3055]), .B(x[3055]), .Z(n37439) );
  AND U31761 ( .A(n26500), .B(n37439), .Z(n51975) );
  AND U31762 ( .A(n14698), .B(n51975), .Z(n14699) );
  NANDN U31763 ( .A(x[3055]), .B(y[3055]), .Z(n26498) );
  NANDN U31764 ( .A(x[3056]), .B(y[3056]), .Z(n26497) );
  NAND U31765 ( .A(n26498), .B(n26497), .Z(n55291) );
  OR U31766 ( .A(n14699), .B(n55291), .Z(n14700) );
  NAND U31767 ( .A(n55292), .B(n14700), .Z(n14701) );
  NANDN U31768 ( .A(n51974), .B(n14701), .Z(n14702) );
  NANDN U31769 ( .A(n55293), .B(n14702), .Z(n14703) );
  XNOR U31770 ( .A(y[3060]), .B(x[3060]), .Z(n37451) );
  NANDN U31771 ( .A(x[3059]), .B(y[3059]), .Z(n26494) );
  AND U31772 ( .A(n37451), .B(n26494), .Z(n51973) );
  AND U31773 ( .A(n14703), .B(n51973), .Z(n14705) );
  NANDN U31774 ( .A(y[3060]), .B(x[3060]), .Z(n14704) );
  NANDN U31775 ( .A(y[3061]), .B(x[3061]), .Z(n37456) );
  NAND U31776 ( .A(n14704), .B(n37456), .Z(n55294) );
  OR U31777 ( .A(n14705), .B(n55294), .Z(n14706) );
  NAND U31778 ( .A(n55295), .B(n14706), .Z(n14707) );
  NANDN U31779 ( .A(n51972), .B(n14707), .Z(n14708) );
  NANDN U31780 ( .A(n55296), .B(n14708), .Z(n14709) );
  AND U31781 ( .A(n55298), .B(n14709), .Z(n14711) );
  NANDN U31782 ( .A(x[3065]), .B(y[3065]), .Z(n26488) );
  XNOR U31783 ( .A(x[3066]), .B(y[3066]), .Z(n14710) );
  NAND U31784 ( .A(n26488), .B(n14710), .Z(n55299) );
  OR U31785 ( .A(n14711), .B(n55299), .Z(n14712) );
  NAND U31786 ( .A(n51971), .B(n14712), .Z(n14713) );
  NANDN U31787 ( .A(n55300), .B(n14713), .Z(n14714) );
  NANDN U31788 ( .A(n55301), .B(n14714), .Z(n14715) );
  AND U31789 ( .A(n55302), .B(n14715), .Z(n14716) );
  NANDN U31790 ( .A(y[3070]), .B(x[3070]), .Z(n37477) );
  NANDN U31791 ( .A(y[3071]), .B(x[3071]), .Z(n37484) );
  NAND U31792 ( .A(n37477), .B(n37484), .Z(n55303) );
  OR U31793 ( .A(n14716), .B(n55303), .Z(n14717) );
  NANDN U31794 ( .A(x[3071]), .B(y[3071]), .Z(n26478) );
  NANDN U31795 ( .A(x[3072]), .B(y[3072]), .Z(n26477) );
  AND U31796 ( .A(n26478), .B(n26477), .Z(n51970) );
  AND U31797 ( .A(n14717), .B(n51970), .Z(n14718) );
  NANDN U31798 ( .A(y[3072]), .B(x[3072]), .Z(n37483) );
  NANDN U31799 ( .A(y[3073]), .B(x[3073]), .Z(n37490) );
  NAND U31800 ( .A(n37483), .B(n37490), .Z(n55304) );
  OR U31801 ( .A(n14718), .B(n55304), .Z(n14719) );
  NAND U31802 ( .A(n55305), .B(n14719), .Z(n14720) );
  NANDN U31803 ( .A(n51969), .B(n14720), .Z(n14721) );
  AND U31804 ( .A(n37496), .B(n14721), .Z(n14722) );
  NAND U31805 ( .A(n55306), .B(n14722), .Z(n14723) );
  NAND U31806 ( .A(n51968), .B(n14723), .Z(n14724) );
  NANDN U31807 ( .A(n55309), .B(n14724), .Z(n14725) );
  NAND U31808 ( .A(n55310), .B(n14725), .Z(n14726) );
  NAND U31809 ( .A(n26472), .B(n14726), .Z(n14727) );
  ANDN U31810 ( .B(y[3079]), .A(x[3079]), .Z(n55311) );
  OR U31811 ( .A(n14727), .B(n55311), .Z(n14728) );
  AND U31812 ( .A(n55312), .B(n14728), .Z(n14729) );
  OR U31813 ( .A(n55313), .B(n14729), .Z(n14730) );
  NAND U31814 ( .A(n55314), .B(n14730), .Z(n14731) );
  NANDN U31815 ( .A(n55315), .B(n14731), .Z(n14732) );
  AND U31816 ( .A(n55316), .B(n14732), .Z(n14733) );
  OR U31817 ( .A(n55317), .B(n14733), .Z(n14734) );
  NAND U31818 ( .A(n55318), .B(n14734), .Z(n14735) );
  NAND U31819 ( .A(n37529), .B(n14735), .Z(n14736) );
  NANDN U31820 ( .A(x[3087]), .B(y[3087]), .Z(n55319) );
  NANDN U31821 ( .A(n14736), .B(n55319), .Z(n14737) );
  AND U31822 ( .A(n55322), .B(n14737), .Z(n14738) );
  OR U31823 ( .A(n55324), .B(n14738), .Z(n14739) );
  NAND U31824 ( .A(n55326), .B(n14739), .Z(n14740) );
  NANDN U31825 ( .A(n55328), .B(n14740), .Z(n14741) );
  NANDN U31826 ( .A(n55330), .B(n14741), .Z(n14742) );
  AND U31827 ( .A(n55332), .B(n14742), .Z(n14743) );
  OR U31828 ( .A(n55334), .B(n14743), .Z(n14744) );
  NAND U31829 ( .A(n55336), .B(n14744), .Z(n14745) );
  NANDN U31830 ( .A(n55338), .B(n14745), .Z(n14746) );
  NANDN U31831 ( .A(n55340), .B(n14746), .Z(n14747) );
  AND U31832 ( .A(n55342), .B(n14747), .Z(n14748) );
  OR U31833 ( .A(n55344), .B(n14748), .Z(n14749) );
  NAND U31834 ( .A(n55346), .B(n14749), .Z(n14750) );
  NANDN U31835 ( .A(n55348), .B(n14750), .Z(n14751) );
  NANDN U31836 ( .A(n55350), .B(n14751), .Z(n14752) );
  AND U31837 ( .A(n55352), .B(n14752), .Z(n14753) );
  OR U31838 ( .A(n55354), .B(n14753), .Z(n14754) );
  NAND U31839 ( .A(n55356), .B(n14754), .Z(n14755) );
  NANDN U31840 ( .A(n55358), .B(n14755), .Z(n14756) );
  NANDN U31841 ( .A(n55360), .B(n14756), .Z(n14757) );
  AND U31842 ( .A(n55362), .B(n14757), .Z(n14758) );
  OR U31843 ( .A(n55363), .B(n14758), .Z(n14759) );
  NAND U31844 ( .A(n55364), .B(n14759), .Z(n14760) );
  NANDN U31845 ( .A(n55365), .B(n14760), .Z(n14761) );
  NANDN U31846 ( .A(n55366), .B(n14761), .Z(n14762) );
  AND U31847 ( .A(n55367), .B(n14762), .Z(n14763) );
  OR U31848 ( .A(n55368), .B(n14763), .Z(n14764) );
  NAND U31849 ( .A(n55369), .B(n14764), .Z(n14765) );
  NAND U31850 ( .A(n55370), .B(n14765), .Z(n14768) );
  NANDN U31851 ( .A(x[3118]), .B(y[3118]), .Z(n14767) );
  NANDN U31852 ( .A(x[3117]), .B(y[3117]), .Z(n14766) );
  NAND U31853 ( .A(n14767), .B(n14766), .Z(n55371) );
  ANDN U31854 ( .B(n14768), .A(n55371), .Z(n14769) );
  NANDN U31855 ( .A(y[3118]), .B(x[3118]), .Z(n37615) );
  NANDN U31856 ( .A(y[3119]), .B(x[3119]), .Z(n26431) );
  AND U31857 ( .A(n37615), .B(n26431), .Z(n55372) );
  NANDN U31858 ( .A(n14769), .B(n55372), .Z(n14770) );
  NANDN U31859 ( .A(n55373), .B(n14770), .Z(n14771) );
  AND U31860 ( .A(n55374), .B(n14771), .Z(n14772) );
  OR U31861 ( .A(n55375), .B(n14772), .Z(n14773) );
  NAND U31862 ( .A(n55376), .B(n14773), .Z(n14774) );
  NANDN U31863 ( .A(n55377), .B(n14774), .Z(n14775) );
  NANDN U31864 ( .A(n55378), .B(n14775), .Z(n14776) );
  AND U31865 ( .A(n55379), .B(n14776), .Z(n14777) );
  NANDN U31866 ( .A(y[3126]), .B(x[3126]), .Z(n26420) );
  NANDN U31867 ( .A(y[3127]), .B(x[3127]), .Z(n26419) );
  NAND U31868 ( .A(n26420), .B(n26419), .Z(n55380) );
  OR U31869 ( .A(n14777), .B(n55380), .Z(n14778) );
  NAND U31870 ( .A(n51966), .B(n14778), .Z(n14779) );
  NANDN U31871 ( .A(n55383), .B(n14779), .Z(n14780) );
  NANDN U31872 ( .A(n55385), .B(n14780), .Z(n14781) );
  AND U31873 ( .A(n55386), .B(n14781), .Z(n14782) );
  NANDN U31874 ( .A(x[3131]), .B(y[3131]), .Z(n26416) );
  NANDN U31875 ( .A(x[3132]), .B(y[3132]), .Z(n26415) );
  AND U31876 ( .A(n26416), .B(n26415), .Z(n55387) );
  NANDN U31877 ( .A(n14782), .B(n55387), .Z(n14783) );
  NANDN U31878 ( .A(n51965), .B(n14783), .Z(n14785) );
  NANDN U31879 ( .A(x[3133]), .B(y[3133]), .Z(n26414) );
  XNOR U31880 ( .A(x[3134]), .B(y[3134]), .Z(n14784) );
  AND U31881 ( .A(n26414), .B(n14784), .Z(n51964) );
  AND U31882 ( .A(n14785), .B(n51964), .Z(n14786) );
  NANDN U31883 ( .A(y[3134]), .B(x[3134]), .Z(n37656) );
  NANDN U31884 ( .A(y[3135]), .B(x[3135]), .Z(n37662) );
  NAND U31885 ( .A(n37656), .B(n37662), .Z(n55388) );
  OR U31886 ( .A(n14786), .B(n55388), .Z(n14787) );
  AND U31887 ( .A(n55389), .B(n14787), .Z(n14788) );
  OR U31888 ( .A(n55390), .B(n14788), .Z(n14789) );
  NAND U31889 ( .A(n55391), .B(n14789), .Z(n14790) );
  NANDN U31890 ( .A(n55392), .B(n14790), .Z(n14792) );
  XNOR U31891 ( .A(x[3140]), .B(y[3140]), .Z(n26408) );
  NANDN U31892 ( .A(x[3139]), .B(y[3139]), .Z(n55393) );
  AND U31893 ( .A(n26408), .B(n55393), .Z(n14791) );
  NAND U31894 ( .A(n14792), .B(n14791), .Z(n14793) );
  AND U31895 ( .A(n55395), .B(n14793), .Z(n14794) );
  OR U31896 ( .A(n55396), .B(n14794), .Z(n14795) );
  NAND U31897 ( .A(n55397), .B(n14795), .Z(n14796) );
  NANDN U31898 ( .A(n55399), .B(n14796), .Z(n14797) );
  NANDN U31899 ( .A(n55400), .B(n14797), .Z(n14798) );
  AND U31900 ( .A(n55401), .B(n14798), .Z(n14799) );
  OR U31901 ( .A(n55402), .B(n14799), .Z(n14800) );
  NAND U31902 ( .A(n55403), .B(n14800), .Z(n14801) );
  NANDN U31903 ( .A(n55404), .B(n14801), .Z(n14802) );
  NANDN U31904 ( .A(n55405), .B(n14802), .Z(n14803) );
  AND U31905 ( .A(n55406), .B(n14803), .Z(n14804) );
  OR U31906 ( .A(n55407), .B(n14804), .Z(n14805) );
  NAND U31907 ( .A(n55408), .B(n14805), .Z(n14806) );
  NANDN U31908 ( .A(n55409), .B(n14806), .Z(n14807) );
  NANDN U31909 ( .A(n55410), .B(n14807), .Z(n14808) );
  AND U31910 ( .A(n55411), .B(n14808), .Z(n14809) );
  NANDN U31911 ( .A(y[3156]), .B(x[3156]), .Z(n37720) );
  NANDN U31912 ( .A(y[3157]), .B(x[3157]), .Z(n37726) );
  NAND U31913 ( .A(n37720), .B(n37726), .Z(n55412) );
  OR U31914 ( .A(n14809), .B(n55412), .Z(n14810) );
  AND U31915 ( .A(n51962), .B(n14810), .Z(n14811) );
  XNOR U31916 ( .A(x[3158]), .B(y[3158]), .Z(n37727) );
  NAND U31917 ( .A(n14811), .B(n37727), .Z(n14812) );
  NANDN U31918 ( .A(n55413), .B(n14812), .Z(n14813) );
  AND U31919 ( .A(n55414), .B(n14813), .Z(n14814) );
  NANDN U31920 ( .A(y[3160]), .B(x[3160]), .Z(n37732) );
  NANDN U31921 ( .A(y[3161]), .B(x[3161]), .Z(n26386) );
  AND U31922 ( .A(n37732), .B(n26386), .Z(n55415) );
  NANDN U31923 ( .A(n14814), .B(n55415), .Z(n14815) );
  NAND U31924 ( .A(n14816), .B(n14815), .Z(n14817) );
  NAND U31925 ( .A(n55418), .B(n14817), .Z(n14818) );
  NAND U31926 ( .A(n26385), .B(n14818), .Z(n14819) );
  NANDN U31927 ( .A(x[3163]), .B(y[3163]), .Z(n55419) );
  NANDN U31928 ( .A(n14819), .B(n55419), .Z(n14820) );
  AND U31929 ( .A(n55421), .B(n14820), .Z(n14821) );
  OR U31930 ( .A(n55422), .B(n14821), .Z(n14822) );
  NAND U31931 ( .A(n55423), .B(n14822), .Z(n14823) );
  NANDN U31932 ( .A(n55424), .B(n14823), .Z(n14824) );
  NANDN U31933 ( .A(n55425), .B(n14824), .Z(n14825) );
  AND U31934 ( .A(n55426), .B(n14825), .Z(n14826) );
  OR U31935 ( .A(n55427), .B(n14826), .Z(n14827) );
  NAND U31936 ( .A(n55428), .B(n14827), .Z(n14828) );
  NANDN U31937 ( .A(n55429), .B(n14828), .Z(n14829) );
  NANDN U31938 ( .A(n55430), .B(n14829), .Z(n14830) );
  AND U31939 ( .A(n55431), .B(n14830), .Z(n14831) );
  OR U31940 ( .A(n55432), .B(n14831), .Z(n14832) );
  NAND U31941 ( .A(n55433), .B(n14832), .Z(n14833) );
  NANDN U31942 ( .A(n55434), .B(n14833), .Z(n14834) );
  NANDN U31943 ( .A(n55436), .B(n14834), .Z(n14835) );
  AND U31944 ( .A(n55437), .B(n14835), .Z(n14836) );
  OR U31945 ( .A(n55438), .B(n14836), .Z(n14837) );
  NAND U31946 ( .A(n55439), .B(n14837), .Z(n14838) );
  NANDN U31947 ( .A(n55440), .B(n14838), .Z(n14839) );
  NANDN U31948 ( .A(n55441), .B(n14839), .Z(n14840) );
  AND U31949 ( .A(n55442), .B(n14840), .Z(n14841) );
  NANDN U31950 ( .A(x[3185]), .B(y[3185]), .Z(n37801) );
  NANDN U31951 ( .A(x[3186]), .B(y[3186]), .Z(n37808) );
  AND U31952 ( .A(n37801), .B(n37808), .Z(n55443) );
  NANDN U31953 ( .A(n14841), .B(n55443), .Z(n14842) );
  NANDN U31954 ( .A(n51960), .B(n14842), .Z(n14843) );
  NANDN U31955 ( .A(x[3187]), .B(y[3187]), .Z(n37807) );
  NANDN U31956 ( .A(x[3188]), .B(y[3188]), .Z(n26357) );
  AND U31957 ( .A(n37807), .B(n26357), .Z(n51959) );
  AND U31958 ( .A(n14843), .B(n51959), .Z(n14844) );
  NANDN U31959 ( .A(y[3188]), .B(x[3188]), .Z(n26358) );
  NANDN U31960 ( .A(y[3189]), .B(x[3189]), .Z(n26355) );
  NAND U31961 ( .A(n26358), .B(n26355), .Z(n51958) );
  OR U31962 ( .A(n14844), .B(n51958), .Z(n14845) );
  AND U31963 ( .A(n26354), .B(n14845), .Z(n14846) );
  NANDN U31964 ( .A(n26356), .B(n14846), .Z(n14848) );
  NANDN U31965 ( .A(y[3190]), .B(x[3190]), .Z(n14847) );
  NANDN U31966 ( .A(y[3191]), .B(x[3191]), .Z(n26353) );
  AND U31967 ( .A(n14847), .B(n26353), .Z(n55444) );
  AND U31968 ( .A(n14848), .B(n55444), .Z(n14850) );
  NANDN U31969 ( .A(x[3192]), .B(y[3192]), .Z(n26351) );
  ANDN U31970 ( .B(y[3191]), .A(x[3191]), .Z(n37817) );
  ANDN U31971 ( .B(n26351), .A(n37817), .Z(n14849) );
  NANDN U31972 ( .A(n14850), .B(n14849), .Z(n14851) );
  AND U31973 ( .A(n14852), .B(n14851), .Z(n14853) );
  OR U31974 ( .A(n55448), .B(n14853), .Z(n14854) );
  NAND U31975 ( .A(n55449), .B(n14854), .Z(n14855) );
  NANDN U31976 ( .A(n55450), .B(n14855), .Z(n14856) );
  NANDN U31977 ( .A(n51953), .B(n14856), .Z(n14857) );
  NANDN U31978 ( .A(x[3197]), .B(y[3197]), .Z(n37834) );
  NANDN U31979 ( .A(x[3198]), .B(y[3198]), .Z(n26346) );
  AND U31980 ( .A(n37834), .B(n26346), .Z(n51952) );
  AND U31981 ( .A(n14857), .B(n51952), .Z(n14858) );
  NANDN U31982 ( .A(y[3198]), .B(x[3198]), .Z(n26347) );
  NANDN U31983 ( .A(y[3199]), .B(x[3199]), .Z(n37841) );
  AND U31984 ( .A(n26347), .B(n37841), .Z(n55451) );
  NANDN U31985 ( .A(n14858), .B(n55451), .Z(n14859) );
  NAND U31986 ( .A(n37842), .B(n14859), .Z(n14860) );
  ANDN U31987 ( .B(y[3199]), .A(x[3199]), .Z(n26345) );
  OR U31988 ( .A(n14860), .B(n26345), .Z(n14862) );
  NANDN U31989 ( .A(y[3200]), .B(x[3200]), .Z(n14861) );
  NANDN U31990 ( .A(y[3201]), .B(x[3201]), .Z(n37848) );
  AND U31991 ( .A(n14861), .B(n37848), .Z(n55452) );
  AND U31992 ( .A(n14862), .B(n55452), .Z(n14863) );
  NANDN U31993 ( .A(x[3201]), .B(y[3201]), .Z(n26344) );
  NANDN U31994 ( .A(x[3202]), .B(y[3202]), .Z(n26343) );
  NAND U31995 ( .A(n26344), .B(n26343), .Z(n51949) );
  OR U31996 ( .A(n14863), .B(n51949), .Z(n14864) );
  NAND U31997 ( .A(n51948), .B(n14864), .Z(n14865) );
  NANDN U31998 ( .A(n55454), .B(n14865), .Z(n14866) );
  AND U31999 ( .A(n55455), .B(n14866), .Z(n14867) );
  OR U32000 ( .A(n55456), .B(n14867), .Z(n14868) );
  NAND U32001 ( .A(n55457), .B(n14868), .Z(n14869) );
  NANDN U32002 ( .A(n55458), .B(n14869), .Z(n14870) );
  NAND U32003 ( .A(n51947), .B(n14870), .Z(n14871) );
  NANDN U32004 ( .A(n55459), .B(n14871), .Z(n14872) );
  NANDN U32005 ( .A(y[3210]), .B(x[3210]), .Z(n37871) );
  NANDN U32006 ( .A(y[3211]), .B(x[3211]), .Z(n37877) );
  AND U32007 ( .A(n37871), .B(n37877), .Z(n55460) );
  AND U32008 ( .A(n14872), .B(n55460), .Z(n14873) );
  XNOR U32009 ( .A(y[3212]), .B(x[3212]), .Z(n37878) );
  NANDN U32010 ( .A(x[3211]), .B(y[3211]), .Z(n26334) );
  NAND U32011 ( .A(n37878), .B(n26334), .Z(n51946) );
  OR U32012 ( .A(n14873), .B(n51946), .Z(n14874) );
  NAND U32013 ( .A(n51945), .B(n14874), .Z(n14875) );
  NANDN U32014 ( .A(n55461), .B(n14875), .Z(n14876) );
  NANDN U32015 ( .A(n55462), .B(n14876), .Z(n14877) );
  XNOR U32016 ( .A(y[3216]), .B(x[3216]), .Z(n37890) );
  NANDN U32017 ( .A(x[3215]), .B(y[3215]), .Z(n26330) );
  AND U32018 ( .A(n37890), .B(n26330), .Z(n55463) );
  AND U32019 ( .A(n14877), .B(n55463), .Z(n14879) );
  NANDN U32020 ( .A(y[3216]), .B(x[3216]), .Z(n14878) );
  NANDN U32021 ( .A(y[3217]), .B(x[3217]), .Z(n37896) );
  NAND U32022 ( .A(n14878), .B(n37896), .Z(n51944) );
  OR U32023 ( .A(n14879), .B(n51944), .Z(n14880) );
  NAND U32024 ( .A(n51943), .B(n14880), .Z(n14881) );
  NANDN U32025 ( .A(n55465), .B(n14881), .Z(n14882) );
  NANDN U32026 ( .A(n55466), .B(n14882), .Z(n14884) );
  NANDN U32027 ( .A(y[3220]), .B(x[3220]), .Z(n14883) );
  NANDN U32028 ( .A(y[3221]), .B(x[3221]), .Z(n37908) );
  AND U32029 ( .A(n14883), .B(n37908), .Z(n55467) );
  AND U32030 ( .A(n14884), .B(n55467), .Z(n14885) );
  ANDN U32031 ( .B(y[3221]), .A(x[3221]), .Z(n26324) );
  NANDN U32032 ( .A(x[3222]), .B(y[3222]), .Z(n26323) );
  NANDN U32033 ( .A(n26324), .B(n26323), .Z(n51942) );
  OR U32034 ( .A(n14885), .B(n51942), .Z(n14886) );
  NAND U32035 ( .A(n51941), .B(n14886), .Z(n14887) );
  NANDN U32036 ( .A(n55468), .B(n14887), .Z(n14888) );
  AND U32037 ( .A(n55469), .B(n14888), .Z(n14889) );
  OR U32038 ( .A(n55470), .B(n14889), .Z(n14890) );
  NAND U32039 ( .A(n55471), .B(n14890), .Z(n14891) );
  NAND U32040 ( .A(n55472), .B(n14891), .Z(n14892) );
  XNOR U32041 ( .A(x[3228]), .B(y[3228]), .Z(n37926) );
  NANDN U32042 ( .A(n14892), .B(n37926), .Z(n14893) );
  NAND U32043 ( .A(n51940), .B(n14893), .Z(n14894) );
  NANDN U32044 ( .A(n55476), .B(n14894), .Z(n14895) );
  NAND U32045 ( .A(n55478), .B(n14895), .Z(n14896) );
  AND U32046 ( .A(n14897), .B(n14896), .Z(n14899) );
  NANDN U32047 ( .A(y[3232]), .B(x[3232]), .Z(n14898) );
  NANDN U32048 ( .A(y[3233]), .B(x[3233]), .Z(n37942) );
  NAND U32049 ( .A(n14898), .B(n37942), .Z(n55481) );
  OR U32050 ( .A(n14899), .B(n55481), .Z(n14900) );
  NAND U32051 ( .A(n55482), .B(n14900), .Z(n14901) );
  NANDN U32052 ( .A(n51939), .B(n14901), .Z(n14902) );
  NANDN U32053 ( .A(n55483), .B(n14902), .Z(n14903) );
  AND U32054 ( .A(n55484), .B(n14903), .Z(n14904) );
  OR U32055 ( .A(n55485), .B(n14904), .Z(n14905) );
  NAND U32056 ( .A(n55486), .B(n14905), .Z(n14906) );
  NANDN U32057 ( .A(n55487), .B(n14906), .Z(n14907) );
  NANDN U32058 ( .A(n51938), .B(n14907), .Z(n14908) );
  NANDN U32059 ( .A(x[3241]), .B(y[3241]), .Z(n37962) );
  NANDN U32060 ( .A(x[3242]), .B(y[3242]), .Z(n37969) );
  AND U32061 ( .A(n37962), .B(n37969), .Z(n51937) );
  AND U32062 ( .A(n14908), .B(n51937), .Z(n14909) );
  NANDN U32063 ( .A(y[3242]), .B(x[3242]), .Z(n26305) );
  NANDN U32064 ( .A(y[3243]), .B(x[3243]), .Z(n26304) );
  NAND U32065 ( .A(n26305), .B(n26304), .Z(n55488) );
  OR U32066 ( .A(n14909), .B(n55488), .Z(n14910) );
  NAND U32067 ( .A(n55491), .B(n14910), .Z(n14911) );
  NANDN U32068 ( .A(n51936), .B(n14911), .Z(n14912) );
  NANDN U32069 ( .A(n55492), .B(n14912), .Z(n14913) );
  NANDN U32070 ( .A(y[3246]), .B(x[3246]), .Z(n26301) );
  NANDN U32071 ( .A(y[3247]), .B(x[3247]), .Z(n26298) );
  AND U32072 ( .A(n26301), .B(n26298), .Z(n51935) );
  AND U32073 ( .A(n14913), .B(n51935), .Z(n14914) );
  NANDN U32074 ( .A(x[3247]), .B(y[3247]), .Z(n26299) );
  NANDN U32075 ( .A(x[3248]), .B(y[3248]), .Z(n37986) );
  NAND U32076 ( .A(n26299), .B(n37986), .Z(n55493) );
  OR U32077 ( .A(n14914), .B(n55493), .Z(n14915) );
  NAND U32078 ( .A(n55494), .B(n14915), .Z(n14916) );
  NANDN U32079 ( .A(n51934), .B(n14916), .Z(n14917) );
  NANDN U32080 ( .A(n55495), .B(n14917), .Z(n14919) );
  NANDN U32081 ( .A(x[3251]), .B(y[3251]), .Z(n37991) );
  XNOR U32082 ( .A(x[3252]), .B(y[3252]), .Z(n14918) );
  AND U32083 ( .A(n37991), .B(n14918), .Z(n51933) );
  AND U32084 ( .A(n14919), .B(n51933), .Z(n14920) );
  NANDN U32085 ( .A(y[3252]), .B(x[3252]), .Z(n26293) );
  NANDN U32086 ( .A(y[3253]), .B(x[3253]), .Z(n38000) );
  NAND U32087 ( .A(n26293), .B(n38000), .Z(n55496) );
  OR U32088 ( .A(n14920), .B(n55496), .Z(n14921) );
  NAND U32089 ( .A(n55497), .B(n14921), .Z(n14922) );
  NANDN U32090 ( .A(n51932), .B(n14922), .Z(n14923) );
  NANDN U32091 ( .A(n55499), .B(n14923), .Z(n14924) );
  NANDN U32092 ( .A(y[3256]), .B(x[3256]), .Z(n38006) );
  NANDN U32093 ( .A(y[3257]), .B(x[3257]), .Z(n38013) );
  AND U32094 ( .A(n38006), .B(n38013), .Z(n51931) );
  AND U32095 ( .A(n14924), .B(n51931), .Z(n14925) );
  NANDN U32096 ( .A(x[3257]), .B(y[3257]), .Z(n26289) );
  NANDN U32097 ( .A(x[3258]), .B(y[3258]), .Z(n26288) );
  NAND U32098 ( .A(n26289), .B(n26288), .Z(n55500) );
  OR U32099 ( .A(n14925), .B(n55500), .Z(n14926) );
  NAND U32100 ( .A(n55501), .B(n14926), .Z(n14927) );
  NANDN U32101 ( .A(n55502), .B(n14927), .Z(n14928) );
  NANDN U32102 ( .A(n55503), .B(n14928), .Z(n14929) );
  NANDN U32103 ( .A(x[3261]), .B(y[3261]), .Z(n26285) );
  NANDN U32104 ( .A(x[3262]), .B(y[3262]), .Z(n26284) );
  AND U32105 ( .A(n26285), .B(n26284), .Z(n55504) );
  AND U32106 ( .A(n14929), .B(n55504), .Z(n14930) );
  NANDN U32107 ( .A(y[3262]), .B(x[3262]), .Z(n38024) );
  NANDN U32108 ( .A(y[3263]), .B(x[3263]), .Z(n38031) );
  NAND U32109 ( .A(n38024), .B(n38031), .Z(n55505) );
  OR U32110 ( .A(n14930), .B(n55505), .Z(n14931) );
  NAND U32111 ( .A(n55506), .B(n14931), .Z(n14932) );
  NANDN U32112 ( .A(n51930), .B(n14932), .Z(n14933) );
  NANDN U32113 ( .A(n55507), .B(n14933), .Z(n14934) );
  AND U32114 ( .A(n55509), .B(n14934), .Z(n14936) );
  XNOR U32115 ( .A(x[3268]), .B(y[3268]), .Z(n26279) );
  NANDN U32116 ( .A(x[3267]), .B(y[3267]), .Z(n51928) );
  AND U32117 ( .A(n26279), .B(n51928), .Z(n14935) );
  NANDN U32118 ( .A(n14936), .B(n14935), .Z(n14937) );
  NANDN U32119 ( .A(n55510), .B(n14937), .Z(n14938) );
  AND U32120 ( .A(n55511), .B(n14938), .Z(n14939) );
  OR U32121 ( .A(n55512), .B(n14939), .Z(n14940) );
  NAND U32122 ( .A(n51927), .B(n14940), .Z(n14941) );
  NANDN U32123 ( .A(n55513), .B(n14941), .Z(n14942) );
  NANDN U32124 ( .A(n55514), .B(n14942), .Z(n14943) );
  AND U32125 ( .A(n55515), .B(n14943), .Z(n14944) );
  OR U32126 ( .A(n55516), .B(n14944), .Z(n14945) );
  NAND U32127 ( .A(n51926), .B(n14945), .Z(n14946) );
  NANDN U32128 ( .A(n55517), .B(n14946), .Z(n14947) );
  NANDN U32129 ( .A(n55518), .B(n14947), .Z(n14948) );
  AND U32130 ( .A(n55519), .B(n14948), .Z(n14949) );
  OR U32131 ( .A(n55520), .B(n14949), .Z(n14950) );
  NAND U32132 ( .A(n51925), .B(n14950), .Z(n14951) );
  NANDN U32133 ( .A(n55522), .B(n14951), .Z(n14952) );
  NANDN U32134 ( .A(n55523), .B(n14952), .Z(n14953) );
  AND U32135 ( .A(n55524), .B(n14953), .Z(n14954) );
  OR U32136 ( .A(n55525), .B(n14954), .Z(n14955) );
  NAND U32137 ( .A(n51924), .B(n14955), .Z(n14956) );
  NANDN U32138 ( .A(n55526), .B(n14956), .Z(n14957) );
  NANDN U32139 ( .A(n55527), .B(n14957), .Z(n14958) );
  AND U32140 ( .A(n55528), .B(n14958), .Z(n14959) );
  OR U32141 ( .A(n55529), .B(n14959), .Z(n14960) );
  NAND U32142 ( .A(n51923), .B(n14960), .Z(n14961) );
  NANDN U32143 ( .A(n55530), .B(n14961), .Z(n14962) );
  NANDN U32144 ( .A(n55531), .B(n14962), .Z(n14963) );
  AND U32145 ( .A(n55532), .B(n14963), .Z(n14964) );
  OR U32146 ( .A(n55534), .B(n14964), .Z(n14965) );
  NAND U32147 ( .A(n51922), .B(n14965), .Z(n14966) );
  NANDN U32148 ( .A(n55535), .B(n14966), .Z(n14967) );
  NANDN U32149 ( .A(n55536), .B(n14967), .Z(n14968) );
  AND U32150 ( .A(n55537), .B(n14968), .Z(n14969) );
  OR U32151 ( .A(n55538), .B(n14969), .Z(n14970) );
  NAND U32152 ( .A(n51921), .B(n14970), .Z(n14971) );
  NANDN U32153 ( .A(n55539), .B(n14971), .Z(n14973) );
  XNOR U32154 ( .A(x[3304]), .B(y[3304]), .Z(n38147) );
  NANDN U32155 ( .A(x[3303]), .B(y[3303]), .Z(n55540) );
  AND U32156 ( .A(n38147), .B(n55540), .Z(n14972) );
  NAND U32157 ( .A(n14973), .B(n14972), .Z(n14975) );
  NANDN U32158 ( .A(y[3304]), .B(x[3304]), .Z(n14974) );
  NANDN U32159 ( .A(y[3305]), .B(x[3305]), .Z(n38153) );
  AND U32160 ( .A(n14974), .B(n38153), .Z(n51920) );
  AND U32161 ( .A(n14975), .B(n51920), .Z(n14976) );
  NANDN U32162 ( .A(x[3305]), .B(y[3305]), .Z(n26241) );
  NANDN U32163 ( .A(x[3306]), .B(y[3306]), .Z(n26240) );
  NAND U32164 ( .A(n26241), .B(n26240), .Z(n55542) );
  OR U32165 ( .A(n14976), .B(n55542), .Z(n14977) );
  NAND U32166 ( .A(n55543), .B(n14977), .Z(n14978) );
  NANDN U32167 ( .A(n51919), .B(n14978), .Z(n14979) );
  NANDN U32168 ( .A(n55546), .B(n14979), .Z(n14980) );
  NANDN U32169 ( .A(x[3309]), .B(y[3309]), .Z(n26237) );
  NANDN U32170 ( .A(x[3310]), .B(y[3310]), .Z(n26236) );
  AND U32171 ( .A(n26237), .B(n26236), .Z(n51918) );
  AND U32172 ( .A(n14980), .B(n51918), .Z(n14981) );
  NANDN U32173 ( .A(y[3310]), .B(x[3310]), .Z(n38164) );
  NANDN U32174 ( .A(y[3311]), .B(x[3311]), .Z(n38171) );
  NAND U32175 ( .A(n38164), .B(n38171), .Z(n55547) );
  OR U32176 ( .A(n14981), .B(n55547), .Z(n14982) );
  NAND U32177 ( .A(n55548), .B(n14982), .Z(n14983) );
  NANDN U32178 ( .A(n51917), .B(n14983), .Z(n14984) );
  NANDN U32179 ( .A(n55549), .B(n14984), .Z(n14985) );
  NANDN U32180 ( .A(y[3314]), .B(x[3314]), .Z(n38176) );
  NANDN U32181 ( .A(y[3315]), .B(x[3315]), .Z(n38183) );
  AND U32182 ( .A(n38176), .B(n38183), .Z(n51916) );
  AND U32183 ( .A(n14985), .B(n51916), .Z(n14986) );
  NANDN U32184 ( .A(x[3315]), .B(y[3315]), .Z(n26231) );
  NANDN U32185 ( .A(x[3316]), .B(y[3316]), .Z(n26230) );
  NAND U32186 ( .A(n26231), .B(n26230), .Z(n55550) );
  OR U32187 ( .A(n14986), .B(n55550), .Z(n14987) );
  NAND U32188 ( .A(n55551), .B(n14987), .Z(n14988) );
  NANDN U32189 ( .A(n51915), .B(n14988), .Z(n14989) );
  NANDN U32190 ( .A(n55552), .B(n14989), .Z(n14990) );
  NANDN U32191 ( .A(x[3319]), .B(y[3319]), .Z(n26227) );
  NANDN U32192 ( .A(x[3320]), .B(y[3320]), .Z(n26226) );
  AND U32193 ( .A(n26227), .B(n26226), .Z(n51914) );
  AND U32194 ( .A(n14990), .B(n51914), .Z(n14991) );
  NANDN U32195 ( .A(y[3320]), .B(x[3320]), .Z(n38194) );
  NANDN U32196 ( .A(y[3321]), .B(x[3321]), .Z(n38201) );
  NAND U32197 ( .A(n38194), .B(n38201), .Z(n55554) );
  OR U32198 ( .A(n14991), .B(n55554), .Z(n14992) );
  NAND U32199 ( .A(n55555), .B(n14992), .Z(n14993) );
  NANDN U32200 ( .A(n51913), .B(n14993), .Z(n14994) );
  NANDN U32201 ( .A(n55556), .B(n14994), .Z(n14995) );
  AND U32202 ( .A(n55557), .B(n14995), .Z(n14996) );
  NANDN U32203 ( .A(x[3325]), .B(y[3325]), .Z(n26221) );
  NANDN U32204 ( .A(x[3326]), .B(y[3326]), .Z(n38217) );
  NAND U32205 ( .A(n26221), .B(n38217), .Z(n55558) );
  OR U32206 ( .A(n14996), .B(n55558), .Z(n14997) );
  NAND U32207 ( .A(n55559), .B(n14997), .Z(n14998) );
  NANDN U32208 ( .A(n51912), .B(n14998), .Z(n14999) );
  NANDN U32209 ( .A(n55560), .B(n14999), .Z(n15000) );
  AND U32210 ( .A(n55561), .B(n15000), .Z(n15001) );
  OR U32211 ( .A(n55562), .B(n15001), .Z(n15002) );
  NAND U32212 ( .A(n55563), .B(n15002), .Z(n15003) );
  NANDN U32213 ( .A(n55565), .B(n15003), .Z(n15004) );
  NANDN U32214 ( .A(n51911), .B(n15004), .Z(n15005) );
  NANDN U32215 ( .A(y[3334]), .B(x[3334]), .Z(n38238) );
  NANDN U32216 ( .A(y[3335]), .B(x[3335]), .Z(n38245) );
  AND U32217 ( .A(n38238), .B(n38245), .Z(n51910) );
  AND U32218 ( .A(n15005), .B(n51910), .Z(n15006) );
  NANDN U32219 ( .A(x[3335]), .B(y[3335]), .Z(n26213) );
  NANDN U32220 ( .A(x[3336]), .B(y[3336]), .Z(n26212) );
  NAND U32221 ( .A(n26213), .B(n26212), .Z(n55566) );
  OR U32222 ( .A(n15006), .B(n55566), .Z(n15007) );
  NAND U32223 ( .A(n55567), .B(n15007), .Z(n15008) );
  NANDN U32224 ( .A(n51909), .B(n15008), .Z(n15009) );
  NANDN U32225 ( .A(n55568), .B(n15009), .Z(n15011) );
  NANDN U32226 ( .A(x[3339]), .B(y[3339]), .Z(n26209) );
  XNOR U32227 ( .A(x[3340]), .B(y[3340]), .Z(n15010) );
  AND U32228 ( .A(n26209), .B(n15010), .Z(n51908) );
  AND U32229 ( .A(n15011), .B(n51908), .Z(n15012) );
  NANDN U32230 ( .A(y[3340]), .B(x[3340]), .Z(n26207) );
  NANDN U32231 ( .A(y[3341]), .B(x[3341]), .Z(n26204) );
  NAND U32232 ( .A(n26207), .B(n26204), .Z(n55569) );
  OR U32233 ( .A(n15012), .B(n55569), .Z(n15013) );
  NAND U32234 ( .A(n55570), .B(n15013), .Z(n15014) );
  NANDN U32235 ( .A(n51907), .B(n15014), .Z(n15016) );
  NANDN U32236 ( .A(x[3343]), .B(y[3343]), .Z(n51906) );
  NANDN U32237 ( .A(x[3344]), .B(y[3344]), .Z(n51905) );
  AND U32238 ( .A(n51906), .B(n51905), .Z(n15015) );
  NAND U32239 ( .A(n15016), .B(n15015), .Z(n15017) );
  AND U32240 ( .A(n15018), .B(n15017), .Z(n15019) );
  OR U32241 ( .A(n55575), .B(n15019), .Z(n15020) );
  NAND U32242 ( .A(n55576), .B(n15020), .Z(n15021) );
  NANDN U32243 ( .A(n55577), .B(n15021), .Z(n15022) );
  NANDN U32244 ( .A(n55578), .B(n15022), .Z(n15023) );
  NANDN U32245 ( .A(x[3349]), .B(y[3349]), .Z(n38277) );
  NANDN U32246 ( .A(x[3350]), .B(y[3350]), .Z(n26194) );
  AND U32247 ( .A(n38277), .B(n26194), .Z(n55579) );
  AND U32248 ( .A(n15023), .B(n55579), .Z(n15024) );
  NANDN U32249 ( .A(y[3350]), .B(x[3350]), .Z(n26195) );
  NANDN U32250 ( .A(y[3351]), .B(x[3351]), .Z(n26192) );
  NAND U32251 ( .A(n26195), .B(n26192), .Z(n51904) );
  OR U32252 ( .A(n15024), .B(n51904), .Z(n15025) );
  NAND U32253 ( .A(n51903), .B(n15025), .Z(n15026) );
  NANDN U32254 ( .A(n51902), .B(n15026), .Z(n15028) );
  XNOR U32255 ( .A(x[3354]), .B(y[3354]), .Z(n26190) );
  NANDN U32256 ( .A(x[3353]), .B(y[3353]), .Z(n51900) );
  AND U32257 ( .A(n26190), .B(n51900), .Z(n15027) );
  NAND U32258 ( .A(n15028), .B(n15027), .Z(n15030) );
  NANDN U32259 ( .A(y[3354]), .B(x[3354]), .Z(n15029) );
  NANDN U32260 ( .A(y[3355]), .B(x[3355]), .Z(n26188) );
  AND U32261 ( .A(n15029), .B(n26188), .Z(n55580) );
  AND U32262 ( .A(n15030), .B(n55580), .Z(n15031) );
  NANDN U32263 ( .A(x[3355]), .B(y[3355]), .Z(n38292) );
  NANDN U32264 ( .A(x[3356]), .B(y[3356]), .Z(n26186) );
  NAND U32265 ( .A(n38292), .B(n26186), .Z(n51899) );
  OR U32266 ( .A(n15031), .B(n51899), .Z(n15032) );
  NAND U32267 ( .A(n51898), .B(n15032), .Z(n15033) );
  NANDN U32268 ( .A(n55583), .B(n15033), .Z(n15034) );
  NANDN U32269 ( .A(n55584), .B(n15034), .Z(n15035) );
  AND U32270 ( .A(n55585), .B(n15035), .Z(n15036) );
  OR U32271 ( .A(n55586), .B(n15036), .Z(n15037) );
  NAND U32272 ( .A(n55587), .B(n15037), .Z(n15038) );
  NANDN U32273 ( .A(n55588), .B(n15038), .Z(n15039) );
  NANDN U32274 ( .A(n55589), .B(n15039), .Z(n15040) );
  NANDN U32275 ( .A(y[3364]), .B(x[3364]), .Z(n38316) );
  NANDN U32276 ( .A(y[3365]), .B(x[3365]), .Z(n38323) );
  AND U32277 ( .A(n38316), .B(n38323), .Z(n55590) );
  AND U32278 ( .A(n15040), .B(n55590), .Z(n15041) );
  NANDN U32279 ( .A(x[3365]), .B(y[3365]), .Z(n26177) );
  NANDN U32280 ( .A(x[3366]), .B(y[3366]), .Z(n26176) );
  NAND U32281 ( .A(n26177), .B(n26176), .Z(n51897) );
  OR U32282 ( .A(n15041), .B(n51897), .Z(n15042) );
  NAND U32283 ( .A(n51896), .B(n15042), .Z(n15043) );
  NANDN U32284 ( .A(n55592), .B(n15043), .Z(n15044) );
  NANDN U32285 ( .A(n55593), .B(n15044), .Z(n15045) );
  NANDN U32286 ( .A(x[3369]), .B(y[3369]), .Z(n26173) );
  NANDN U32287 ( .A(x[3370]), .B(y[3370]), .Z(n26172) );
  AND U32288 ( .A(n26173), .B(n26172), .Z(n55594) );
  AND U32289 ( .A(n15045), .B(n55594), .Z(n15046) );
  NANDN U32290 ( .A(y[3370]), .B(x[3370]), .Z(n38334) );
  NANDN U32291 ( .A(y[3371]), .B(x[3371]), .Z(n38341) );
  NAND U32292 ( .A(n38334), .B(n38341), .Z(n51895) );
  OR U32293 ( .A(n15046), .B(n51895), .Z(n15047) );
  NAND U32294 ( .A(n51894), .B(n15047), .Z(n15048) );
  NANDN U32295 ( .A(n55595), .B(n15048), .Z(n15049) );
  NANDN U32296 ( .A(n55596), .B(n15049), .Z(n15050) );
  AND U32297 ( .A(n55597), .B(n15050), .Z(n15051) );
  NANDN U32298 ( .A(x[3375]), .B(y[3375]), .Z(n26167) );
  NANDN U32299 ( .A(x[3376]), .B(y[3376]), .Z(n38357) );
  NAND U32300 ( .A(n26167), .B(n38357), .Z(n51893) );
  OR U32301 ( .A(n15051), .B(n51893), .Z(n15052) );
  NAND U32302 ( .A(n51892), .B(n15052), .Z(n15053) );
  NANDN U32303 ( .A(n55598), .B(n15053), .Z(n15054) );
  NANDN U32304 ( .A(n55599), .B(n15054), .Z(n15055) );
  NANDN U32305 ( .A(x[3379]), .B(y[3379]), .Z(n26165) );
  NANDN U32306 ( .A(x[3380]), .B(y[3380]), .Z(n26164) );
  AND U32307 ( .A(n26165), .B(n26164), .Z(n55600) );
  AND U32308 ( .A(n15055), .B(n55600), .Z(n15056) );
  NANDN U32309 ( .A(y[3380]), .B(x[3380]), .Z(n38366) );
  NANDN U32310 ( .A(y[3381]), .B(x[3381]), .Z(n38375) );
  AND U32311 ( .A(n38366), .B(n38375), .Z(n55603) );
  NANDN U32312 ( .A(n15056), .B(n55603), .Z(n15057) );
  NAND U32313 ( .A(n38373), .B(n15057), .Z(n15058) );
  NANDN U32314 ( .A(x[3381]), .B(y[3381]), .Z(n55604) );
  NANDN U32315 ( .A(n15058), .B(n55604), .Z(n15060) );
  NANDN U32316 ( .A(y[3382]), .B(x[3382]), .Z(n15059) );
  NANDN U32317 ( .A(y[3383]), .B(x[3383]), .Z(n38381) );
  AND U32318 ( .A(n15059), .B(n38381), .Z(n51891) );
  AND U32319 ( .A(n15060), .B(n51891), .Z(n15061) );
  ANDN U32320 ( .B(y[3383]), .A(x[3383]), .Z(n38377) );
  NANDN U32321 ( .A(x[3384]), .B(y[3384]), .Z(n26163) );
  NANDN U32322 ( .A(n38377), .B(n26163), .Z(n55606) );
  OR U32323 ( .A(n15061), .B(n55606), .Z(n15062) );
  NAND U32324 ( .A(n55607), .B(n15062), .Z(n15063) );
  NANDN U32325 ( .A(n51890), .B(n15063), .Z(n15064) );
  NANDN U32326 ( .A(n55608), .B(n15064), .Z(n15065) );
  NANDN U32327 ( .A(x[3387]), .B(y[3387]), .Z(n26160) );
  NANDN U32328 ( .A(x[3388]), .B(y[3388]), .Z(n26157) );
  AND U32329 ( .A(n26160), .B(n26157), .Z(n51889) );
  AND U32330 ( .A(n15065), .B(n51889), .Z(n15066) );
  NANDN U32331 ( .A(y[3388]), .B(x[3388]), .Z(n26158) );
  NANDN U32332 ( .A(y[3389]), .B(x[3389]), .Z(n26155) );
  AND U32333 ( .A(n26158), .B(n26155), .Z(n55609) );
  NANDN U32334 ( .A(n15066), .B(n55609), .Z(n15067) );
  NAND U32335 ( .A(n26154), .B(n15067), .Z(n15068) );
  ANDN U32336 ( .B(y[3389]), .A(x[3389]), .Z(n26156) );
  OR U32337 ( .A(n15068), .B(n26156), .Z(n15070) );
  NANDN U32338 ( .A(y[3390]), .B(x[3390]), .Z(n15069) );
  NANDN U32339 ( .A(y[3391]), .B(x[3391]), .Z(n26153) );
  AND U32340 ( .A(n15069), .B(n26153), .Z(n51888) );
  AND U32341 ( .A(n15070), .B(n51888), .Z(n15071) );
  NANDN U32342 ( .A(x[3391]), .B(y[3391]), .Z(n38397) );
  NANDN U32343 ( .A(x[3392]), .B(y[3392]), .Z(n26151) );
  NAND U32344 ( .A(n38397), .B(n26151), .Z(n55612) );
  OR U32345 ( .A(n15071), .B(n55612), .Z(n15072) );
  NAND U32346 ( .A(n55615), .B(n15072), .Z(n15073) );
  NANDN U32347 ( .A(n51887), .B(n15073), .Z(n15074) );
  NAND U32348 ( .A(n51886), .B(n15074), .Z(n15075) );
  AND U32349 ( .A(n15076), .B(n15075), .Z(n15078) );
  NANDN U32350 ( .A(y[3396]), .B(x[3396]), .Z(n15077) );
  NANDN U32351 ( .A(y[3397]), .B(x[3397]), .Z(n38413) );
  NAND U32352 ( .A(n15077), .B(n38413), .Z(n55619) );
  OR U32353 ( .A(n15078), .B(n55619), .Z(n15079) );
  AND U32354 ( .A(n38414), .B(n15079), .Z(n15080) );
  NANDN U32355 ( .A(x[3397]), .B(y[3397]), .Z(n55620) );
  AND U32356 ( .A(n15080), .B(n55620), .Z(n15081) );
  OR U32357 ( .A(n55622), .B(n15081), .Z(n15082) );
  NAND U32358 ( .A(n55623), .B(n15082), .Z(n15083) );
  NANDN U32359 ( .A(n55624), .B(n15083), .Z(n15084) );
  NAND U32360 ( .A(n55625), .B(n15084), .Z(n15085) );
  NANDN U32361 ( .A(n55626), .B(n15085), .Z(n15086) );
  NANDN U32362 ( .A(x[3403]), .B(y[3403]), .Z(n26141) );
  NANDN U32363 ( .A(x[3404]), .B(y[3404]), .Z(n26140) );
  AND U32364 ( .A(n26141), .B(n26140), .Z(n51885) );
  AND U32365 ( .A(n15086), .B(n51885), .Z(n15087) );
  NANDN U32366 ( .A(y[3404]), .B(x[3404]), .Z(n38431) );
  NANDN U32367 ( .A(y[3405]), .B(x[3405]), .Z(n38438) );
  NAND U32368 ( .A(n38431), .B(n38438), .Z(n55627) );
  OR U32369 ( .A(n15087), .B(n55627), .Z(n15088) );
  NAND U32370 ( .A(n55628), .B(n15088), .Z(n15089) );
  NANDN U32371 ( .A(n51884), .B(n15089), .Z(n15090) );
  AND U32372 ( .A(n38444), .B(n15090), .Z(n15091) );
  NAND U32373 ( .A(n51883), .B(n15091), .Z(n15092) );
  NANDN U32374 ( .A(n55632), .B(n15092), .Z(n15093) );
  AND U32375 ( .A(n55633), .B(n15093), .Z(n15094) );
  OR U32376 ( .A(n55634), .B(n15094), .Z(n15095) );
  NAND U32377 ( .A(n55635), .B(n15095), .Z(n15096) );
  NANDN U32378 ( .A(n55636), .B(n15096), .Z(n15097) );
  NANDN U32379 ( .A(n55637), .B(n15097), .Z(n15098) );
  AND U32380 ( .A(n55638), .B(n15098), .Z(n15099) );
  OR U32381 ( .A(n55639), .B(n15099), .Z(n15100) );
  NAND U32382 ( .A(n55640), .B(n15100), .Z(n15101) );
  NAND U32383 ( .A(n55641), .B(n15101), .Z(n15102) );
  XNOR U32384 ( .A(x[3418]), .B(y[3418]), .Z(n26127) );
  NANDN U32385 ( .A(n15102), .B(n26127), .Z(n15103) );
  NANDN U32386 ( .A(n55643), .B(n15103), .Z(n15104) );
  AND U32387 ( .A(n55644), .B(n15104), .Z(n15105) );
  OR U32388 ( .A(n55646), .B(n15105), .Z(n15106) );
  NAND U32389 ( .A(n55647), .B(n15106), .Z(n15107) );
  NANDN U32390 ( .A(n55648), .B(n15107), .Z(n15109) );
  XNOR U32391 ( .A(x[3424]), .B(y[3424]), .Z(n38489) );
  NANDN U32392 ( .A(x[3423]), .B(y[3423]), .Z(n55649) );
  AND U32393 ( .A(n38489), .B(n55649), .Z(n15108) );
  NAND U32394 ( .A(n15109), .B(n15108), .Z(n15110) );
  AND U32395 ( .A(n55651), .B(n15110), .Z(n15111) );
  OR U32396 ( .A(n55652), .B(n15111), .Z(n15112) );
  NAND U32397 ( .A(n55653), .B(n15112), .Z(n15113) );
  NANDN U32398 ( .A(n55654), .B(n15113), .Z(n15114) );
  NANDN U32399 ( .A(n55655), .B(n15114), .Z(n15115) );
  NANDN U32400 ( .A(x[3429]), .B(y[3429]), .Z(n26119) );
  NANDN U32401 ( .A(x[3430]), .B(y[3430]), .Z(n26116) );
  AND U32402 ( .A(n26119), .B(n26116), .Z(n55656) );
  AND U32403 ( .A(n15115), .B(n55656), .Z(n15116) );
  NANDN U32404 ( .A(y[3430]), .B(x[3430]), .Z(n26118) );
  ANDN U32405 ( .B(x[3431]), .A(y[3431]), .Z(n38512) );
  ANDN U32406 ( .B(n26118), .A(n38512), .Z(n55657) );
  NANDN U32407 ( .A(n15116), .B(n55657), .Z(n15117) );
  NAND U32408 ( .A(n38513), .B(n15117), .Z(n15118) );
  NANDN U32409 ( .A(x[3431]), .B(y[3431]), .Z(n55658) );
  NANDN U32410 ( .A(n15118), .B(n55658), .Z(n15119) );
  AND U32411 ( .A(n55660), .B(n15119), .Z(n15120) );
  OR U32412 ( .A(n55661), .B(n15120), .Z(n15121) );
  NAND U32413 ( .A(n55662), .B(n15121), .Z(n15122) );
  NANDN U32414 ( .A(n55664), .B(n15122), .Z(n15123) );
  NANDN U32415 ( .A(n55666), .B(n15123), .Z(n15124) );
  AND U32416 ( .A(n55668), .B(n15124), .Z(n15125) );
  OR U32417 ( .A(n55670), .B(n15125), .Z(n15126) );
  NAND U32418 ( .A(n55672), .B(n15126), .Z(n15127) );
  NANDN U32419 ( .A(n55674), .B(n15127), .Z(n15128) );
  NANDN U32420 ( .A(n55676), .B(n15128), .Z(n15129) );
  AND U32421 ( .A(n55678), .B(n15129), .Z(n15130) );
  OR U32422 ( .A(n55680), .B(n15130), .Z(n15131) );
  NAND U32423 ( .A(n55682), .B(n15131), .Z(n15132) );
  NANDN U32424 ( .A(n55684), .B(n15132), .Z(n15133) );
  NANDN U32425 ( .A(n55686), .B(n15133), .Z(n15134) );
  AND U32426 ( .A(n55688), .B(n15134), .Z(n15135) );
  OR U32427 ( .A(n55690), .B(n15135), .Z(n15136) );
  NAND U32428 ( .A(n55692), .B(n15136), .Z(n15137) );
  NANDN U32429 ( .A(n55694), .B(n15137), .Z(n15138) );
  NANDN U32430 ( .A(n55696), .B(n15138), .Z(n15139) );
  AND U32431 ( .A(n55698), .B(n15139), .Z(n15140) );
  OR U32432 ( .A(n55700), .B(n15140), .Z(n15141) );
  NAND U32433 ( .A(n55702), .B(n15141), .Z(n15142) );
  NANDN U32434 ( .A(n55704), .B(n15142), .Z(n15143) );
  NANDN U32435 ( .A(n55706), .B(n15143), .Z(n15144) );
  AND U32436 ( .A(n55708), .B(n15144), .Z(n15145) );
  OR U32437 ( .A(n55710), .B(n15145), .Z(n15146) );
  NAND U32438 ( .A(n55712), .B(n15146), .Z(n15147) );
  NANDN U32439 ( .A(n55714), .B(n15147), .Z(n15149) );
  XNOR U32440 ( .A(x[3462]), .B(y[3462]), .Z(n38591) );
  NANDN U32441 ( .A(x[3461]), .B(y[3461]), .Z(n55715) );
  AND U32442 ( .A(n38591), .B(n55715), .Z(n15148) );
  NAND U32443 ( .A(n15149), .B(n15148), .Z(n15150) );
  AND U32444 ( .A(n55720), .B(n15150), .Z(n15151) );
  OR U32445 ( .A(n55722), .B(n15151), .Z(n15152) );
  NAND U32446 ( .A(n55724), .B(n15152), .Z(n15153) );
  NANDN U32447 ( .A(n55726), .B(n15153), .Z(n15154) );
  NANDN U32448 ( .A(n55728), .B(n15154), .Z(n15155) );
  AND U32449 ( .A(n55730), .B(n15155), .Z(n15156) );
  OR U32450 ( .A(n55732), .B(n15156), .Z(n15157) );
  NAND U32451 ( .A(n55734), .B(n15157), .Z(n15158) );
  NANDN U32452 ( .A(n55736), .B(n15158), .Z(n15159) );
  NANDN U32453 ( .A(n55738), .B(n15159), .Z(n15160) );
  AND U32454 ( .A(n55740), .B(n15160), .Z(n15161) );
  OR U32455 ( .A(n55742), .B(n15161), .Z(n15162) );
  NAND U32456 ( .A(n55744), .B(n15162), .Z(n15163) );
  NANDN U32457 ( .A(n55745), .B(n15163), .Z(n15164) );
  NAND U32458 ( .A(n55746), .B(n15164), .Z(n15165) );
  AND U32459 ( .A(n15166), .B(n15165), .Z(n15167) );
  OR U32460 ( .A(n55747), .B(n15167), .Z(n15168) );
  NAND U32461 ( .A(n55748), .B(n15168), .Z(n15169) );
  NANDN U32462 ( .A(n55749), .B(n15169), .Z(n15170) );
  NANDN U32463 ( .A(n55750), .B(n15170), .Z(n15171) );
  AND U32464 ( .A(n55751), .B(n15171), .Z(n15172) );
  OR U32465 ( .A(n55752), .B(n15172), .Z(n15173) );
  NAND U32466 ( .A(n55753), .B(n15173), .Z(n15174) );
  NANDN U32467 ( .A(n55754), .B(n15174), .Z(n15175) );
  NANDN U32468 ( .A(n55755), .B(n15175), .Z(n15176) );
  AND U32469 ( .A(n55756), .B(n15176), .Z(n15177) );
  OR U32470 ( .A(n55757), .B(n15177), .Z(n15178) );
  NAND U32471 ( .A(n55758), .B(n15178), .Z(n15179) );
  NANDN U32472 ( .A(n55759), .B(n15179), .Z(n15180) );
  NANDN U32473 ( .A(n51880), .B(n15180), .Z(n15181) );
  NANDN U32474 ( .A(y[3492]), .B(x[3492]), .Z(n38677) );
  NANDN U32475 ( .A(y[3493]), .B(x[3493]), .Z(n26044) );
  AND U32476 ( .A(n38677), .B(n26044), .Z(n51879) );
  AND U32477 ( .A(n15181), .B(n51879), .Z(n15182) );
  OR U32478 ( .A(n55762), .B(n15182), .Z(n15183) );
  NAND U32479 ( .A(n55763), .B(n15183), .Z(n15184) );
  NAND U32480 ( .A(n55764), .B(n15184), .Z(n15185) );
  XNOR U32481 ( .A(y[3496]), .B(x[3496]), .Z(n26041) );
  NANDN U32482 ( .A(n15185), .B(n26041), .Z(n15186) );
  NAND U32483 ( .A(n55765), .B(n15186), .Z(n15187) );
  NAND U32484 ( .A(n55766), .B(n15187), .Z(n15188) );
  ANDN U32485 ( .B(y[3497]), .A(x[3497]), .Z(n26039) );
  OR U32486 ( .A(n15188), .B(n26039), .Z(n15189) );
  AND U32487 ( .A(n55767), .B(n15189), .Z(n15190) );
  NANDN U32488 ( .A(x[3499]), .B(y[3499]), .Z(n26037) );
  NANDN U32489 ( .A(x[3500]), .B(y[3500]), .Z(n26034) );
  NAND U32490 ( .A(n26037), .B(n26034), .Z(n55768) );
  OR U32491 ( .A(n15190), .B(n55768), .Z(n15191) );
  AND U32492 ( .A(n55769), .B(n15191), .Z(n15192) );
  OR U32493 ( .A(n55770), .B(n15192), .Z(n15193) );
  NAND U32494 ( .A(n55771), .B(n15193), .Z(n15194) );
  NANDN U32495 ( .A(n55772), .B(n15194), .Z(n15195) );
  AND U32496 ( .A(n55773), .B(n15195), .Z(n15196) );
  XNOR U32497 ( .A(x[3506]), .B(y[3506]), .Z(n38711) );
  NANDN U32498 ( .A(n15196), .B(n38711), .Z(n15197) );
  NANDN U32499 ( .A(x[3505]), .B(y[3505]), .Z(n55774) );
  NANDN U32500 ( .A(n15197), .B(n55774), .Z(n15198) );
  AND U32501 ( .A(n55776), .B(n15198), .Z(n15199) );
  OR U32502 ( .A(n55777), .B(n15199), .Z(n15200) );
  NAND U32503 ( .A(n55779), .B(n15200), .Z(n15201) );
  NANDN U32504 ( .A(n55780), .B(n15201), .Z(n15202) );
  NANDN U32505 ( .A(n55781), .B(n15202), .Z(n15203) );
  NANDN U32506 ( .A(x[3511]), .B(y[3511]), .Z(n38724) );
  NANDN U32507 ( .A(x[3512]), .B(y[3512]), .Z(n38731) );
  AND U32508 ( .A(n38724), .B(n38731), .Z(n55782) );
  AND U32509 ( .A(n15203), .B(n55782), .Z(n15204) );
  NANDN U32510 ( .A(y[3512]), .B(x[3512]), .Z(n26022) );
  NANDN U32511 ( .A(y[3513]), .B(x[3513]), .Z(n26021) );
  NAND U32512 ( .A(n26022), .B(n26021), .Z(n51876) );
  OR U32513 ( .A(n15204), .B(n51876), .Z(n15205) );
  NAND U32514 ( .A(n51875), .B(n15205), .Z(n15206) );
  NANDN U32515 ( .A(n51874), .B(n15206), .Z(n15207) );
  NANDN U32516 ( .A(n55783), .B(n15207), .Z(n15208) );
  AND U32517 ( .A(n55784), .B(n15208), .Z(n15209) );
  OR U32518 ( .A(n55785), .B(n15209), .Z(n15210) );
  NAND U32519 ( .A(n55786), .B(n15210), .Z(n15211) );
  NANDN U32520 ( .A(n55787), .B(n15211), .Z(n15212) );
  NANDN U32521 ( .A(n55788), .B(n15212), .Z(n15213) );
  AND U32522 ( .A(n55789), .B(n15213), .Z(n15214) );
  OR U32523 ( .A(n55790), .B(n15214), .Z(n15215) );
  NAND U32524 ( .A(n55792), .B(n15215), .Z(n15216) );
  NANDN U32525 ( .A(n55793), .B(n15216), .Z(n15217) );
  AND U32526 ( .A(n26010), .B(n15217), .Z(n15218) );
  NANDN U32527 ( .A(x[3525]), .B(y[3525]), .Z(n55795) );
  NAND U32528 ( .A(n15218), .B(n55795), .Z(n15219) );
  NANDN U32529 ( .A(n55796), .B(n15219), .Z(n15220) );
  AND U32530 ( .A(n55797), .B(n15220), .Z(n15221) );
  NANDN U32531 ( .A(y[3528]), .B(x[3528]), .Z(n38775) );
  NANDN U32532 ( .A(y[3529]), .B(x[3529]), .Z(n38782) );
  NAND U32533 ( .A(n38775), .B(n38782), .Z(n51873) );
  OR U32534 ( .A(n15221), .B(n51873), .Z(n15222) );
  NAND U32535 ( .A(n51872), .B(n15222), .Z(n15223) );
  NANDN U32536 ( .A(n51871), .B(n15223), .Z(n15224) );
  NAND U32537 ( .A(n38787), .B(n15224), .Z(n15225) );
  ANDN U32538 ( .B(y[3531]), .A(x[3531]), .Z(n26005) );
  OR U32539 ( .A(n15225), .B(n26005), .Z(n15226) );
  NAND U32540 ( .A(n55798), .B(n15226), .Z(n15227) );
  NANDN U32541 ( .A(n51868), .B(n15227), .Z(n15228) );
  NANDN U32542 ( .A(y[3534]), .B(x[3534]), .Z(n26003) );
  NANDN U32543 ( .A(y[3535]), .B(x[3535]), .Z(n25999) );
  AND U32544 ( .A(n26003), .B(n25999), .Z(n51867) );
  AND U32545 ( .A(n15228), .B(n51867), .Z(n15230) );
  XNOR U32546 ( .A(x[3536]), .B(y[3536]), .Z(n26000) );
  ANDN U32547 ( .B(y[3535]), .A(x[3535]), .Z(n26001) );
  ANDN U32548 ( .B(n26000), .A(n26001), .Z(n15229) );
  NANDN U32549 ( .A(n15230), .B(n15229), .Z(n15231) );
  AND U32550 ( .A(n55802), .B(n15231), .Z(n15232) );
  OR U32551 ( .A(n55803), .B(n15232), .Z(n15233) );
  NAND U32552 ( .A(n55804), .B(n15233), .Z(n15234) );
  NANDN U32553 ( .A(n55805), .B(n15234), .Z(n15235) );
  AND U32554 ( .A(n55806), .B(n15235), .Z(n15237) );
  XNOR U32555 ( .A(x[3542]), .B(y[3542]), .Z(n38813) );
  NANDN U32556 ( .A(x[3541]), .B(y[3541]), .Z(n51865) );
  NAND U32557 ( .A(n38813), .B(n51865), .Z(n15236) );
  OR U32558 ( .A(n15237), .B(n15236), .Z(n15239) );
  NANDN U32559 ( .A(y[3542]), .B(x[3542]), .Z(n15238) );
  NANDN U32560 ( .A(y[3543]), .B(x[3543]), .Z(n38819) );
  AND U32561 ( .A(n15238), .B(n38819), .Z(n55807) );
  AND U32562 ( .A(n15239), .B(n55807), .Z(n15240) );
  NANDN U32563 ( .A(x[3543]), .B(y[3543]), .Z(n25993) );
  NANDN U32564 ( .A(x[3544]), .B(y[3544]), .Z(n25992) );
  NAND U32565 ( .A(n25993), .B(n25992), .Z(n51864) );
  OR U32566 ( .A(n15240), .B(n51864), .Z(n15241) );
  NAND U32567 ( .A(n55808), .B(n15241), .Z(n15242) );
  NANDN U32568 ( .A(n55809), .B(n15242), .Z(n15243) );
  AND U32569 ( .A(n55810), .B(n15243), .Z(n15244) );
  OR U32570 ( .A(n55811), .B(n15244), .Z(n15245) );
  NAND U32571 ( .A(n55812), .B(n15245), .Z(n15246) );
  NAND U32572 ( .A(n55814), .B(n15246), .Z(n15248) );
  XOR U32573 ( .A(x[3550]), .B(y[3550]), .Z(n15247) );
  OR U32574 ( .A(n15248), .B(n15247), .Z(n15249) );
  NAND U32575 ( .A(n55817), .B(n15249), .Z(n15250) );
  NANDN U32576 ( .A(n55818), .B(n15250), .Z(n15251) );
  AND U32577 ( .A(n55819), .B(n15251), .Z(n15252) );
  NANDN U32578 ( .A(x[3553]), .B(y[3553]), .Z(n25984) );
  NANDN U32579 ( .A(x[3554]), .B(y[3554]), .Z(n38852) );
  NAND U32580 ( .A(n25984), .B(n38852), .Z(n51863) );
  OR U32581 ( .A(n15252), .B(n51863), .Z(n15253) );
  NANDN U32582 ( .A(y[3554]), .B(x[3554]), .Z(n25982) );
  NANDN U32583 ( .A(y[3555]), .B(x[3555]), .Z(n38854) );
  AND U32584 ( .A(n25982), .B(n38854), .Z(n51862) );
  AND U32585 ( .A(n15253), .B(n51862), .Z(n15254) );
  OR U32586 ( .A(n55820), .B(n15254), .Z(n15255) );
  NAND U32587 ( .A(n55821), .B(n15255), .Z(n15256) );
  NANDN U32588 ( .A(n55822), .B(n15256), .Z(n15257) );
  AND U32589 ( .A(n55823), .B(n15257), .Z(n15258) );
  NANDN U32590 ( .A(x[3559]), .B(y[3559]), .Z(n38863) );
  NANDN U32591 ( .A(x[3560]), .B(y[3560]), .Z(n38870) );
  AND U32592 ( .A(n38863), .B(n38870), .Z(n51861) );
  NANDN U32593 ( .A(n15258), .B(n51861), .Z(n15259) );
  NANDN U32594 ( .A(n55824), .B(n15259), .Z(n15260) );
  AND U32595 ( .A(n55825), .B(n15260), .Z(n15261) );
  OR U32596 ( .A(n55826), .B(n15261), .Z(n15262) );
  NAND U32597 ( .A(n55827), .B(n15262), .Z(n15263) );
  NANDN U32598 ( .A(n55829), .B(n15263), .Z(n15264) );
  NANDN U32599 ( .A(x[3565]), .B(y[3565]), .Z(n25972) );
  NANDN U32600 ( .A(x[3566]), .B(y[3566]), .Z(n25969) );
  AND U32601 ( .A(n25972), .B(n25969), .Z(n51860) );
  AND U32602 ( .A(n15264), .B(n51860), .Z(n15265) );
  ANDN U32603 ( .B(x[3567]), .A(y[3567]), .Z(n38888) );
  NANDN U32604 ( .A(y[3566]), .B(x[3566]), .Z(n25971) );
  NANDN U32605 ( .A(n38888), .B(n25971), .Z(n55830) );
  OR U32606 ( .A(n15265), .B(n55830), .Z(n15266) );
  AND U32607 ( .A(n15267), .B(n15266), .Z(n15268) );
  OR U32608 ( .A(n55833), .B(n15268), .Z(n15269) );
  NAND U32609 ( .A(n55834), .B(n15269), .Z(n15270) );
  NANDN U32610 ( .A(n55835), .B(n15270), .Z(n15271) );
  AND U32611 ( .A(n25964), .B(n15271), .Z(n15272) );
  NANDN U32612 ( .A(n25965), .B(n15272), .Z(n15273) );
  NAND U32613 ( .A(n55838), .B(n15273), .Z(n15274) );
  NANDN U32614 ( .A(n55839), .B(n15274), .Z(n15275) );
  AND U32615 ( .A(n55840), .B(n15275), .Z(n15276) );
  NANDN U32616 ( .A(x[3575]), .B(y[3575]), .Z(n38905) );
  NANDN U32617 ( .A(x[3576]), .B(y[3576]), .Z(n38912) );
  NAND U32618 ( .A(n38905), .B(n38912), .Z(n55841) );
  OR U32619 ( .A(n15276), .B(n55841), .Z(n15277) );
  NANDN U32620 ( .A(y[3576]), .B(x[3576]), .Z(n25959) );
  NANDN U32621 ( .A(y[3577]), .B(x[3577]), .Z(n25958) );
  AND U32622 ( .A(n25959), .B(n25958), .Z(n51859) );
  AND U32623 ( .A(n15277), .B(n51859), .Z(n15278) );
  NANDN U32624 ( .A(x[3577]), .B(y[3577]), .Z(n38911) );
  NANDN U32625 ( .A(x[3578]), .B(y[3578]), .Z(n38920) );
  NAND U32626 ( .A(n38911), .B(n38920), .Z(n55842) );
  OR U32627 ( .A(n15278), .B(n55842), .Z(n15279) );
  NAND U32628 ( .A(n55843), .B(n15279), .Z(n15280) );
  NANDN U32629 ( .A(n51858), .B(n15280), .Z(n15281) );
  AND U32630 ( .A(n55845), .B(n15281), .Z(n15282) );
  OR U32631 ( .A(n55846), .B(n15282), .Z(n15283) );
  NAND U32632 ( .A(n55847), .B(n15283), .Z(n15284) );
  AND U32633 ( .A(n38934), .B(n15284), .Z(n15285) );
  NANDN U32634 ( .A(x[3583]), .B(y[3583]), .Z(n55848) );
  AND U32635 ( .A(n15285), .B(n55848), .Z(n15287) );
  NANDN U32636 ( .A(y[3584]), .B(x[3584]), .Z(n15286) );
  NANDN U32637 ( .A(y[3585]), .B(x[3585]), .Z(n38939) );
  NAND U32638 ( .A(n15286), .B(n38939), .Z(n55850) );
  OR U32639 ( .A(n15287), .B(n55850), .Z(n15288) );
  AND U32640 ( .A(n55851), .B(n15288), .Z(n15289) );
  OR U32641 ( .A(n55852), .B(n15289), .Z(n15290) );
  NAND U32642 ( .A(n55853), .B(n15290), .Z(n15291) );
  NANDN U32643 ( .A(n55854), .B(n15291), .Z(n15292) );
  AND U32644 ( .A(n55855), .B(n15292), .Z(n15293) );
  NANDN U32645 ( .A(y[3590]), .B(x[3590]), .Z(n25949) );
  NANDN U32646 ( .A(y[3591]), .B(x[3591]), .Z(n38960) );
  AND U32647 ( .A(n25949), .B(n38960), .Z(n55856) );
  NANDN U32648 ( .A(n15293), .B(n55856), .Z(n15294) );
  NANDN U32649 ( .A(n55857), .B(n15294), .Z(n15295) );
  AND U32650 ( .A(n55858), .B(n15295), .Z(n15296) );
  OR U32651 ( .A(n55859), .B(n15296), .Z(n15297) );
  NAND U32652 ( .A(n51857), .B(n15297), .Z(n15298) );
  NANDN U32653 ( .A(n55860), .B(n15298), .Z(n15299) );
  NANDN U32654 ( .A(y[3596]), .B(x[3596]), .Z(n25943) );
  NANDN U32655 ( .A(y[3597]), .B(x[3597]), .Z(n38979) );
  AND U32656 ( .A(n25943), .B(n38979), .Z(n55863) );
  AND U32657 ( .A(n15299), .B(n55863), .Z(n15300) );
  XNOR U32658 ( .A(y[3598]), .B(x[3598]), .Z(n38978) );
  NANDN U32659 ( .A(x[3597]), .B(y[3597]), .Z(n38973) );
  NAND U32660 ( .A(n38978), .B(n38973), .Z(n51856) );
  OR U32661 ( .A(n15300), .B(n51856), .Z(n15302) );
  NANDN U32662 ( .A(y[3598]), .B(x[3598]), .Z(n15301) );
  NANDN U32663 ( .A(y[3599]), .B(x[3599]), .Z(n38985) );
  AND U32664 ( .A(n15301), .B(n38985), .Z(n51855) );
  AND U32665 ( .A(n15302), .B(n51855), .Z(n15303) );
  OR U32666 ( .A(n55864), .B(n15303), .Z(n15304) );
  NAND U32667 ( .A(n55865), .B(n15304), .Z(n15305) );
  NANDN U32668 ( .A(n55866), .B(n15305), .Z(n15306) );
  AND U32669 ( .A(n55867), .B(n15306), .Z(n15307) );
  NANDN U32670 ( .A(x[3603]), .B(y[3603]), .Z(n25937) );
  NANDN U32671 ( .A(x[3604]), .B(y[3604]), .Z(n39000) );
  AND U32672 ( .A(n25937), .B(n39000), .Z(n51854) );
  NANDN U32673 ( .A(n15307), .B(n51854), .Z(n15308) );
  NANDN U32674 ( .A(n55868), .B(n15308), .Z(n15309) );
  AND U32675 ( .A(n55869), .B(n15309), .Z(n15310) );
  OR U32676 ( .A(n55870), .B(n15310), .Z(n15311) );
  NAND U32677 ( .A(n55871), .B(n15311), .Z(n15312) );
  NANDN U32678 ( .A(n55872), .B(n15312), .Z(n15313) );
  AND U32679 ( .A(n55873), .B(n15313), .Z(n15314) );
  NANDN U32680 ( .A(y[3610]), .B(x[3610]), .Z(n25931) );
  NANDN U32681 ( .A(y[3611]), .B(x[3611]), .Z(n25930) );
  NAND U32682 ( .A(n25931), .B(n25930), .Z(n55874) );
  OR U32683 ( .A(n15314), .B(n55874), .Z(n15315) );
  AND U32684 ( .A(n55876), .B(n15315), .Z(n15316) );
  NANDN U32685 ( .A(y[3612]), .B(x[3612]), .Z(n25929) );
  NANDN U32686 ( .A(y[3613]), .B(x[3613]), .Z(n25927) );
  AND U32687 ( .A(n25929), .B(n25927), .Z(n55877) );
  NANDN U32688 ( .A(n15316), .B(n55877), .Z(n15317) );
  NANDN U32689 ( .A(n15318), .B(n15317), .Z(n15320) );
  NANDN U32690 ( .A(y[3614]), .B(x[3614]), .Z(n15319) );
  NANDN U32691 ( .A(y[3615]), .B(x[3615]), .Z(n25926) );
  AND U32692 ( .A(n15319), .B(n25926), .Z(n55879) );
  AND U32693 ( .A(n15320), .B(n55879), .Z(n15321) );
  NANDN U32694 ( .A(x[3615]), .B(y[3615]), .Z(n39029) );
  NANDN U32695 ( .A(x[3616]), .B(y[3616]), .Z(n25924) );
  NAND U32696 ( .A(n39029), .B(n25924), .Z(n51851) );
  OR U32697 ( .A(n15321), .B(n51851), .Z(n15322) );
  NAND U32698 ( .A(n51850), .B(n15322), .Z(n15323) );
  NANDN U32699 ( .A(n55880), .B(n15323), .Z(n15324) );
  NANDN U32700 ( .A(y[3618]), .B(x[3618]), .Z(n39035) );
  NANDN U32701 ( .A(y[3619]), .B(x[3619]), .Z(n25922) );
  AND U32702 ( .A(n39035), .B(n25922), .Z(n55881) );
  AND U32703 ( .A(n15324), .B(n55881), .Z(n15325) );
  NANDN U32704 ( .A(x[3619]), .B(y[3619]), .Z(n39039) );
  NANDN U32705 ( .A(x[3620]), .B(y[3620]), .Z(n39046) );
  NAND U32706 ( .A(n39039), .B(n39046), .Z(n55882) );
  OR U32707 ( .A(n15325), .B(n55882), .Z(n15326) );
  NANDN U32708 ( .A(y[3620]), .B(x[3620]), .Z(n25921) );
  NANDN U32709 ( .A(y[3621]), .B(x[3621]), .Z(n25920) );
  AND U32710 ( .A(n25921), .B(n25920), .Z(n55883) );
  AND U32711 ( .A(n15326), .B(n55883), .Z(n15327) );
  NANDN U32712 ( .A(x[3621]), .B(y[3621]), .Z(n39045) );
  NANDN U32713 ( .A(x[3622]), .B(y[3622]), .Z(n39052) );
  NAND U32714 ( .A(n39045), .B(n39052), .Z(n51849) );
  OR U32715 ( .A(n15327), .B(n51849), .Z(n15328) );
  NAND U32716 ( .A(n51848), .B(n15328), .Z(n15329) );
  NANDN U32717 ( .A(n55885), .B(n15329), .Z(n15330) );
  NANDN U32718 ( .A(y[3624]), .B(x[3624]), .Z(n25917) );
  NANDN U32719 ( .A(y[3625]), .B(x[3625]), .Z(n25916) );
  AND U32720 ( .A(n25917), .B(n25916), .Z(n55886) );
  AND U32721 ( .A(n15330), .B(n55886), .Z(n15331) );
  NANDN U32722 ( .A(x[3625]), .B(y[3625]), .Z(n39058) );
  NANDN U32723 ( .A(x[3626]), .B(y[3626]), .Z(n39065) );
  NAND U32724 ( .A(n39058), .B(n39065), .Z(n51847) );
  OR U32725 ( .A(n15331), .B(n51847), .Z(n15332) );
  NAND U32726 ( .A(n51846), .B(n15332), .Z(n15333) );
  NANDN U32727 ( .A(n55887), .B(n15333), .Z(n15334) );
  NANDN U32728 ( .A(y[3628]), .B(x[3628]), .Z(n25913) );
  NANDN U32729 ( .A(y[3629]), .B(x[3629]), .Z(n39073) );
  AND U32730 ( .A(n25913), .B(n39073), .Z(n55888) );
  AND U32731 ( .A(n15334), .B(n55888), .Z(n15336) );
  XNOR U32732 ( .A(x[3630]), .B(y[3630]), .Z(n39074) );
  ANDN U32733 ( .B(y[3629]), .A(x[3629]), .Z(n39069) );
  ANDN U32734 ( .B(n39074), .A(n39069), .Z(n15335) );
  NANDN U32735 ( .A(n15336), .B(n15335), .Z(n15338) );
  NANDN U32736 ( .A(y[3630]), .B(x[3630]), .Z(n15337) );
  NANDN U32737 ( .A(y[3631]), .B(x[3631]), .Z(n39080) );
  AND U32738 ( .A(n15337), .B(n39080), .Z(n55889) );
  AND U32739 ( .A(n15338), .B(n55889), .Z(n15339) );
  NANDN U32740 ( .A(x[3631]), .B(y[3631]), .Z(n25912) );
  NANDN U32741 ( .A(x[3632]), .B(y[3632]), .Z(n25911) );
  NAND U32742 ( .A(n25912), .B(n25911), .Z(n51843) );
  OR U32743 ( .A(n15339), .B(n51843), .Z(n15340) );
  NAND U32744 ( .A(n51842), .B(n15340), .Z(n15341) );
  NANDN U32745 ( .A(n55892), .B(n15341), .Z(n15342) );
  NANDN U32746 ( .A(y[3634]), .B(x[3634]), .Z(n39085) );
  NANDN U32747 ( .A(y[3635]), .B(x[3635]), .Z(n39091) );
  AND U32748 ( .A(n39085), .B(n39091), .Z(n55894) );
  AND U32749 ( .A(n15342), .B(n55894), .Z(n15343) );
  XNOR U32750 ( .A(y[3636]), .B(x[3636]), .Z(n39092) );
  NANDN U32751 ( .A(x[3635]), .B(y[3635]), .Z(n25908) );
  NAND U32752 ( .A(n39092), .B(n25908), .Z(n55895) );
  OR U32753 ( .A(n15343), .B(n55895), .Z(n15345) );
  NANDN U32754 ( .A(y[3636]), .B(x[3636]), .Z(n15344) );
  NANDN U32755 ( .A(y[3637]), .B(x[3637]), .Z(n39098) );
  AND U32756 ( .A(n15344), .B(n39098), .Z(n55896) );
  AND U32757 ( .A(n15345), .B(n55896), .Z(n15346) );
  NANDN U32758 ( .A(x[3637]), .B(y[3637]), .Z(n25906) );
  NANDN U32759 ( .A(x[3638]), .B(y[3638]), .Z(n25905) );
  NAND U32760 ( .A(n25906), .B(n25905), .Z(n51841) );
  OR U32761 ( .A(n15346), .B(n51841), .Z(n15347) );
  NAND U32762 ( .A(n51840), .B(n15347), .Z(n15348) );
  NANDN U32763 ( .A(n55897), .B(n15348), .Z(n15349) );
  NANDN U32764 ( .A(y[3640]), .B(x[3640]), .Z(n39104) );
  NANDN U32765 ( .A(y[3641]), .B(x[3641]), .Z(n39113) );
  AND U32766 ( .A(n39104), .B(n39113), .Z(n55898) );
  AND U32767 ( .A(n15349), .B(n55898), .Z(n15350) );
  ANDN U32768 ( .B(y[3641]), .A(x[3641]), .Z(n39108) );
  NANDN U32769 ( .A(x[3642]), .B(y[3642]), .Z(n25903) );
  NANDN U32770 ( .A(n39108), .B(n25903), .Z(n51839) );
  OR U32771 ( .A(n15350), .B(n51839), .Z(n15351) );
  NAND U32772 ( .A(n51838), .B(n15351), .Z(n15352) );
  NANDN U32773 ( .A(n55899), .B(n15352), .Z(n15353) );
  AND U32774 ( .A(n55902), .B(n15353), .Z(n15354) );
  ANDN U32775 ( .B(n51837), .A(n15354), .Z(n15355) );
  NAND U32776 ( .A(n39124), .B(n15355), .Z(n15356) );
  NANDN U32777 ( .A(n55903), .B(n15356), .Z(n15357) );
  NANDN U32778 ( .A(x[3648]), .B(y[3648]), .Z(n55906) );
  AND U32779 ( .A(n15357), .B(n55906), .Z(n15358) );
  NAND U32780 ( .A(n55904), .B(n15358), .Z(n15359) );
  NANDN U32781 ( .A(n55905), .B(n15359), .Z(n15360) );
  AND U32782 ( .A(n55908), .B(n15360), .Z(n15362) );
  NANDN U32783 ( .A(y[3650]), .B(x[3650]), .Z(n15361) );
  NANDN U32784 ( .A(y[3651]), .B(x[3651]), .Z(n25895) );
  NAND U32785 ( .A(n15361), .B(n25895), .Z(n55909) );
  OR U32786 ( .A(n15362), .B(n55909), .Z(n15363) );
  NAND U32787 ( .A(n55910), .B(n15363), .Z(n15364) );
  NANDN U32788 ( .A(n51835), .B(n15364), .Z(n15365) );
  AND U32789 ( .A(n55912), .B(n15365), .Z(n15366) );
  NANDN U32790 ( .A(y[3654]), .B(x[3654]), .Z(n25893) );
  NANDN U32791 ( .A(y[3655]), .B(x[3655]), .Z(n25890) );
  NAND U32792 ( .A(n25893), .B(n25890), .Z(n55913) );
  OR U32793 ( .A(n15366), .B(n55913), .Z(n15367) );
  AND U32794 ( .A(n15368), .B(n15367), .Z(n15370) );
  NANDN U32795 ( .A(y[3656]), .B(x[3656]), .Z(n15369) );
  NANDN U32796 ( .A(y[3657]), .B(x[3657]), .Z(n25888) );
  NAND U32797 ( .A(n15369), .B(n25888), .Z(n55916) );
  OR U32798 ( .A(n15370), .B(n55916), .Z(n15371) );
  NAND U32799 ( .A(n55917), .B(n15371), .Z(n15372) );
  NANDN U32800 ( .A(n51834), .B(n15372), .Z(n15373) );
  NANDN U32801 ( .A(x[3659]), .B(y[3659]), .Z(n25885) );
  NANDN U32802 ( .A(x[3660]), .B(y[3660]), .Z(n25882) );
  AND U32803 ( .A(n25885), .B(n25882), .Z(n51833) );
  AND U32804 ( .A(n15373), .B(n51833), .Z(n15374) );
  NANDN U32805 ( .A(y[3660]), .B(x[3660]), .Z(n25883) );
  NANDN U32806 ( .A(y[3661]), .B(x[3661]), .Z(n25880) );
  NAND U32807 ( .A(n25883), .B(n25880), .Z(n55918) );
  OR U32808 ( .A(n15374), .B(n55918), .Z(n15375) );
  AND U32809 ( .A(n15376), .B(n15375), .Z(n15378) );
  NANDN U32810 ( .A(y[3662]), .B(x[3662]), .Z(n15377) );
  NANDN U32811 ( .A(y[3663]), .B(x[3663]), .Z(n25879) );
  NAND U32812 ( .A(n15377), .B(n25879), .Z(n55921) );
  OR U32813 ( .A(n15378), .B(n55921), .Z(n15379) );
  NAND U32814 ( .A(n55922), .B(n15379), .Z(n15380) );
  NANDN U32815 ( .A(n51832), .B(n15380), .Z(n15381) );
  NANDN U32816 ( .A(x[3665]), .B(y[3665]), .Z(n25876) );
  NANDN U32817 ( .A(x[3666]), .B(y[3666]), .Z(n25875) );
  AND U32818 ( .A(n25876), .B(n25875), .Z(n51831) );
  AND U32819 ( .A(n15381), .B(n51831), .Z(n15382) );
  NANDN U32820 ( .A(y[3666]), .B(x[3666]), .Z(n39171) );
  NANDN U32821 ( .A(y[3667]), .B(x[3667]), .Z(n39178) );
  NAND U32822 ( .A(n39171), .B(n39178), .Z(n55924) );
  OR U32823 ( .A(n15382), .B(n55924), .Z(n15383) );
  NANDN U32824 ( .A(x[3667]), .B(y[3667]), .Z(n25874) );
  NANDN U32825 ( .A(x[3668]), .B(y[3668]), .Z(n25873) );
  AND U32826 ( .A(n25874), .B(n25873), .Z(n55925) );
  AND U32827 ( .A(n15383), .B(n55925), .Z(n15384) );
  NANDN U32828 ( .A(y[3668]), .B(x[3668]), .Z(n39177) );
  NANDN U32829 ( .A(y[3669]), .B(x[3669]), .Z(n39184) );
  NAND U32830 ( .A(n39177), .B(n39184), .Z(n55926) );
  OR U32831 ( .A(n15384), .B(n55926), .Z(n15385) );
  NAND U32832 ( .A(n55927), .B(n15385), .Z(n15386) );
  NANDN U32833 ( .A(n51830), .B(n15386), .Z(n15387) );
  NANDN U32834 ( .A(x[3671]), .B(y[3671]), .Z(n39187) );
  NANDN U32835 ( .A(x[3672]), .B(y[3672]), .Z(n25869) );
  AND U32836 ( .A(n39187), .B(n25869), .Z(n51829) );
  AND U32837 ( .A(n15387), .B(n51829), .Z(n15388) );
  NANDN U32838 ( .A(y[3672]), .B(x[3672]), .Z(n25870) );
  NANDN U32839 ( .A(y[3673]), .B(x[3673]), .Z(n25867) );
  AND U32840 ( .A(n25870), .B(n25867), .Z(n55928) );
  NANDN U32841 ( .A(n15388), .B(n55928), .Z(n15389) );
  NANDN U32842 ( .A(n51828), .B(n15389), .Z(n15390) );
  NANDN U32843 ( .A(y[3674]), .B(x[3674]), .Z(n25866) );
  NANDN U32844 ( .A(y[3675]), .B(x[3675]), .Z(n25862) );
  AND U32845 ( .A(n25866), .B(n25862), .Z(n51827) );
  AND U32846 ( .A(n15390), .B(n51827), .Z(n15391) );
  NANDN U32847 ( .A(x[3675]), .B(y[3675]), .Z(n25864) );
  NANDN U32848 ( .A(x[3676]), .B(y[3676]), .Z(n39203) );
  NAND U32849 ( .A(n25864), .B(n39203), .Z(n55931) );
  OR U32850 ( .A(n15391), .B(n55931), .Z(n15392) );
  NAND U32851 ( .A(n55933), .B(n15392), .Z(n15393) );
  NANDN U32852 ( .A(n51826), .B(n15393), .Z(n15394) );
  NANDN U32853 ( .A(y[3678]), .B(x[3678]), .Z(n25860) );
  NANDN U32854 ( .A(y[3679]), .B(x[3679]), .Z(n25857) );
  AND U32855 ( .A(n25860), .B(n25857), .Z(n51825) );
  AND U32856 ( .A(n15394), .B(n51825), .Z(n15395) );
  NANDN U32857 ( .A(x[3679]), .B(y[3679]), .Z(n25858) );
  NANDN U32858 ( .A(x[3680]), .B(y[3680]), .Z(n25855) );
  NAND U32859 ( .A(n25858), .B(n25855), .Z(n55934) );
  OR U32860 ( .A(n15395), .B(n55934), .Z(n15396) );
  NANDN U32861 ( .A(y[3680]), .B(x[3680]), .Z(n25856) );
  NANDN U32862 ( .A(y[3681]), .B(x[3681]), .Z(n39213) );
  AND U32863 ( .A(n25856), .B(n39213), .Z(n55935) );
  AND U32864 ( .A(n15396), .B(n55935), .Z(n15397) );
  NANDN U32865 ( .A(x[3681]), .B(y[3681]), .Z(n25854) );
  NANDN U32866 ( .A(x[3682]), .B(y[3682]), .Z(n39217) );
  AND U32867 ( .A(n25854), .B(n39217), .Z(n55936) );
  NANDN U32868 ( .A(n15397), .B(n55936), .Z(n15398) );
  NANDN U32869 ( .A(y[3682]), .B(x[3682]), .Z(n39212) );
  NANDN U32870 ( .A(y[3683]), .B(x[3683]), .Z(n25853) );
  AND U32871 ( .A(n39212), .B(n25853), .Z(n55937) );
  AND U32872 ( .A(n15398), .B(n55937), .Z(n15399) );
  ANDN U32873 ( .B(n55938), .A(n15399), .Z(n15400) );
  OR U32874 ( .A(n55939), .B(n15400), .Z(n15401) );
  NAND U32875 ( .A(n55940), .B(n15401), .Z(n15402) );
  NANDN U32876 ( .A(n55941), .B(n15402), .Z(n15403) );
  NANDN U32877 ( .A(x[3687]), .B(y[3687]), .Z(n39228) );
  NANDN U32878 ( .A(x[3688]), .B(y[3688]), .Z(n39235) );
  AND U32879 ( .A(n39228), .B(n39235), .Z(n51824) );
  AND U32880 ( .A(n15403), .B(n51824), .Z(n15404) );
  NANDN U32881 ( .A(y[3688]), .B(x[3688]), .Z(n25848) );
  NANDN U32882 ( .A(y[3689]), .B(x[3689]), .Z(n25847) );
  NAND U32883 ( .A(n25848), .B(n25847), .Z(n55943) );
  OR U32884 ( .A(n15404), .B(n55943), .Z(n15405) );
  NANDN U32885 ( .A(x[3689]), .B(y[3689]), .Z(n39234) );
  NANDN U32886 ( .A(x[3690]), .B(y[3690]), .Z(n25845) );
  AND U32887 ( .A(n39234), .B(n25845), .Z(n55944) );
  AND U32888 ( .A(n15405), .B(n55944), .Z(n15406) );
  NANDN U32889 ( .A(y[3690]), .B(x[3690]), .Z(n25846) );
  NANDN U32890 ( .A(y[3691]), .B(x[3691]), .Z(n25842) );
  NAND U32891 ( .A(n25846), .B(n25842), .Z(n51823) );
  OR U32892 ( .A(n15406), .B(n51823), .Z(n15407) );
  NAND U32893 ( .A(n51822), .B(n15407), .Z(n15408) );
  NANDN U32894 ( .A(n55945), .B(n15408), .Z(n15409) );
  AND U32895 ( .A(n39248), .B(n15409), .Z(n15410) );
  NANDN U32896 ( .A(x[3693]), .B(y[3693]), .Z(n55946) );
  AND U32897 ( .A(n15410), .B(n55946), .Z(n15412) );
  NANDN U32898 ( .A(y[3694]), .B(x[3694]), .Z(n15411) );
  NANDN U32899 ( .A(y[3695]), .B(x[3695]), .Z(n25840) );
  NAND U32900 ( .A(n15411), .B(n25840), .Z(n55948) );
  OR U32901 ( .A(n15412), .B(n55948), .Z(n15413) );
  NANDN U32902 ( .A(x[3695]), .B(y[3695]), .Z(n39250) );
  NANDN U32903 ( .A(x[3696]), .B(y[3696]), .Z(n25838) );
  AND U32904 ( .A(n39250), .B(n25838), .Z(n55949) );
  AND U32905 ( .A(n15413), .B(n55949), .Z(n15414) );
  NANDN U32906 ( .A(y[3696]), .B(x[3696]), .Z(n25839) );
  NANDN U32907 ( .A(y[3697]), .B(x[3697]), .Z(n25836) );
  NAND U32908 ( .A(n25839), .B(n25836), .Z(n51821) );
  OR U32909 ( .A(n15414), .B(n51821), .Z(n15415) );
  NAND U32910 ( .A(n51820), .B(n15415), .Z(n15416) );
  NANDN U32911 ( .A(n55951), .B(n15416), .Z(n15417) );
  AND U32912 ( .A(n55952), .B(n15417), .Z(n15418) );
  NANDN U32913 ( .A(y[3700]), .B(x[3700]), .Z(n25833) );
  NANDN U32914 ( .A(y[3701]), .B(x[3701]), .Z(n25832) );
  NAND U32915 ( .A(n25833), .B(n25832), .Z(n55953) );
  OR U32916 ( .A(n15418), .B(n55953), .Z(n15419) );
  NAND U32917 ( .A(n55954), .B(n15419), .Z(n15420) );
  NANDN U32918 ( .A(n51819), .B(n15420), .Z(n15421) );
  NANDN U32919 ( .A(x[3703]), .B(y[3703]), .Z(n25829) );
  NANDN U32920 ( .A(x[3704]), .B(y[3704]), .Z(n25826) );
  AND U32921 ( .A(n25829), .B(n25826), .Z(n51818) );
  AND U32922 ( .A(n15421), .B(n51818), .Z(n15422) );
  NANDN U32923 ( .A(y[3704]), .B(x[3704]), .Z(n25827) );
  NANDN U32924 ( .A(y[3705]), .B(x[3705]), .Z(n25824) );
  AND U32925 ( .A(n25827), .B(n25824), .Z(n55955) );
  NANDN U32926 ( .A(n15422), .B(n55955), .Z(n15423) );
  AND U32927 ( .A(n15424), .B(n15423), .Z(n15425) );
  OR U32928 ( .A(n55958), .B(n15425), .Z(n15426) );
  NAND U32929 ( .A(n55959), .B(n15426), .Z(n15427) );
  NANDN U32930 ( .A(n55960), .B(n15427), .Z(n15428) );
  AND U32931 ( .A(n55961), .B(n15428), .Z(n15429) );
  NANDN U32932 ( .A(y[3710]), .B(x[3710]), .Z(n39289) );
  NANDN U32933 ( .A(y[3711]), .B(x[3711]), .Z(n39296) );
  NAND U32934 ( .A(n39289), .B(n39296), .Z(n55963) );
  OR U32935 ( .A(n15429), .B(n55963), .Z(n15430) );
  AND U32936 ( .A(n55964), .B(n15430), .Z(n15431) );
  OR U32937 ( .A(n55965), .B(n15431), .Z(n15432) );
  NAND U32938 ( .A(n55966), .B(n15432), .Z(n15433) );
  NANDN U32939 ( .A(n55967), .B(n15433), .Z(n15434) );
  NANDN U32940 ( .A(x[3715]), .B(y[3715]), .Z(n39304) );
  NANDN U32941 ( .A(x[3716]), .B(y[3716]), .Z(n39311) );
  AND U32942 ( .A(n39304), .B(n39311), .Z(n51817) );
  AND U32943 ( .A(n15434), .B(n51817), .Z(n15435) );
  NANDN U32944 ( .A(y[3716]), .B(x[3716]), .Z(n25816) );
  NANDN U32945 ( .A(y[3717]), .B(x[3717]), .Z(n25815) );
  NAND U32946 ( .A(n25816), .B(n25815), .Z(n55968) );
  OR U32947 ( .A(n15435), .B(n55968), .Z(n15436) );
  NAND U32948 ( .A(n55969), .B(n15436), .Z(n15437) );
  NANDN U32949 ( .A(n51816), .B(n15437), .Z(n15438) );
  NAND U32950 ( .A(n51815), .B(n15438), .Z(n15439) );
  NAND U32951 ( .A(n55970), .B(n15439), .Z(n15440) );
  ANDN U32952 ( .B(y[3721]), .A(x[3721]), .Z(n25810) );
  ANDN U32953 ( .B(n15440), .A(n25810), .Z(n15441) );
  NAND U32954 ( .A(n25809), .B(n15441), .Z(n15442) );
  NAND U32955 ( .A(n55973), .B(n15442), .Z(n15443) );
  XOR U32956 ( .A(x[3724]), .B(y[3724]), .Z(n39329) );
  ANDN U32957 ( .B(n15443), .A(n39329), .Z(n15444) );
  NANDN U32958 ( .A(x[3723]), .B(y[3723]), .Z(n55974) );
  AND U32959 ( .A(n15444), .B(n55974), .Z(n15445) );
  OR U32960 ( .A(n55978), .B(n15445), .Z(n15446) );
  NAND U32961 ( .A(n55979), .B(n15446), .Z(n15447) );
  NANDN U32962 ( .A(n55980), .B(n15447), .Z(n15448) );
  AND U32963 ( .A(n55981), .B(n15448), .Z(n15449) );
  OR U32964 ( .A(n55982), .B(n15449), .Z(n15450) );
  NAND U32965 ( .A(n15451), .B(n15450), .Z(n15453) );
  NANDN U32966 ( .A(y[3730]), .B(x[3730]), .Z(n15452) );
  NANDN U32967 ( .A(y[3731]), .B(x[3731]), .Z(n39351) );
  AND U32968 ( .A(n15452), .B(n39351), .Z(n55985) );
  AND U32969 ( .A(n15453), .B(n55985), .Z(n15455) );
  XNOR U32970 ( .A(x[3732]), .B(y[3732]), .Z(n39352) );
  ANDN U32971 ( .B(y[3731]), .A(x[3731]), .Z(n25802) );
  ANDN U32972 ( .B(n39352), .A(n25802), .Z(n15454) );
  NANDN U32973 ( .A(n15455), .B(n15454), .Z(n15457) );
  NANDN U32974 ( .A(y[3732]), .B(x[3732]), .Z(n15456) );
  NANDN U32975 ( .A(y[3733]), .B(x[3733]), .Z(n39358) );
  AND U32976 ( .A(n15456), .B(n39358), .Z(n55986) );
  AND U32977 ( .A(n15457), .B(n55986), .Z(n15458) );
  NANDN U32978 ( .A(x[3733]), .B(y[3733]), .Z(n25801) );
  NANDN U32979 ( .A(x[3734]), .B(y[3734]), .Z(n25800) );
  NAND U32980 ( .A(n25801), .B(n25800), .Z(n51812) );
  OR U32981 ( .A(n15458), .B(n51812), .Z(n15459) );
  NAND U32982 ( .A(n51811), .B(n15459), .Z(n15460) );
  NANDN U32983 ( .A(n55987), .B(n15460), .Z(n15461) );
  AND U32984 ( .A(n55988), .B(n15461), .Z(n15462) );
  NANDN U32985 ( .A(x[3737]), .B(y[3737]), .Z(n25797) );
  NANDN U32986 ( .A(x[3738]), .B(y[3738]), .Z(n25796) );
  NAND U32987 ( .A(n25797), .B(n25796), .Z(n55990) );
  OR U32988 ( .A(n15462), .B(n55990), .Z(n15463) );
  NANDN U32989 ( .A(y[3738]), .B(x[3738]), .Z(n39372) );
  NANDN U32990 ( .A(y[3739]), .B(x[3739]), .Z(n25794) );
  AND U32991 ( .A(n39372), .B(n25794), .Z(n55991) );
  AND U32992 ( .A(n15463), .B(n55991), .Z(n15464) );
  NANDN U32993 ( .A(x[3739]), .B(y[3739]), .Z(n25795) );
  NANDN U32994 ( .A(x[3740]), .B(y[3740]), .Z(n25792) );
  NAND U32995 ( .A(n25795), .B(n25792), .Z(n51810) );
  OR U32996 ( .A(n15464), .B(n51810), .Z(n15465) );
  NAND U32997 ( .A(n51809), .B(n15465), .Z(n15466) );
  NANDN U32998 ( .A(n55992), .B(n15466), .Z(n15467) );
  AND U32999 ( .A(n55993), .B(n15467), .Z(n15468) );
  NANDN U33000 ( .A(x[3743]), .B(y[3743]), .Z(n25789) );
  NANDN U33001 ( .A(x[3744]), .B(y[3744]), .Z(n25788) );
  AND U33002 ( .A(n25789), .B(n25788), .Z(n51808) );
  NANDN U33003 ( .A(n15468), .B(n51808), .Z(n15469) );
  NANDN U33004 ( .A(n55994), .B(n15469), .Z(n15470) );
  NANDN U33005 ( .A(x[3745]), .B(y[3745]), .Z(n25787) );
  NANDN U33006 ( .A(x[3746]), .B(y[3746]), .Z(n25786) );
  AND U33007 ( .A(n25787), .B(n25786), .Z(n55995) );
  AND U33008 ( .A(n15470), .B(n55995), .Z(n15471) );
  NANDN U33009 ( .A(y[3746]), .B(x[3746]), .Z(n39392) );
  NANDN U33010 ( .A(y[3747]), .B(x[3747]), .Z(n25783) );
  NAND U33011 ( .A(n39392), .B(n25783), .Z(n51807) );
  OR U33012 ( .A(n15471), .B(n51807), .Z(n15472) );
  NAND U33013 ( .A(n51806), .B(n15472), .Z(n15473) );
  NANDN U33014 ( .A(n51805), .B(n15473), .Z(n15474) );
  AND U33015 ( .A(n55997), .B(n15474), .Z(n15476) );
  NANDN U33016 ( .A(y[3750]), .B(x[3750]), .Z(n15475) );
  NANDN U33017 ( .A(y[3751]), .B(x[3751]), .Z(n25780) );
  NAND U33018 ( .A(n15475), .B(n25780), .Z(n55998) );
  OR U33019 ( .A(n15476), .B(n55998), .Z(n15477) );
  AND U33020 ( .A(n55999), .B(n15477), .Z(n15478) );
  NANDN U33021 ( .A(y[3752]), .B(x[3752]), .Z(n25779) );
  NANDN U33022 ( .A(y[3753]), .B(x[3753]), .Z(n25775) );
  NAND U33023 ( .A(n25779), .B(n25775), .Z(n56000) );
  OR U33024 ( .A(n15478), .B(n56000), .Z(n15479) );
  NAND U33025 ( .A(n51804), .B(n15479), .Z(n15480) );
  NANDN U33026 ( .A(n56001), .B(n15480), .Z(n15481) );
  AND U33027 ( .A(n56002), .B(n15481), .Z(n15483) );
  NANDN U33028 ( .A(y[3756]), .B(x[3756]), .Z(n15482) );
  NANDN U33029 ( .A(y[3757]), .B(x[3757]), .Z(n25772) );
  AND U33030 ( .A(n15482), .B(n25772), .Z(n56003) );
  NANDN U33031 ( .A(n15483), .B(n56003), .Z(n15484) );
  NANDN U33032 ( .A(n56004), .B(n15484), .Z(n15485) );
  AND U33033 ( .A(n56005), .B(n15485), .Z(n15486) );
  OR U33034 ( .A(n56006), .B(n15486), .Z(n15487) );
  NAND U33035 ( .A(n56007), .B(n15487), .Z(n15488) );
  NANDN U33036 ( .A(n56008), .B(n15488), .Z(n15489) );
  AND U33037 ( .A(n56010), .B(n15489), .Z(n15490) );
  NANDN U33038 ( .A(x[3763]), .B(y[3763]), .Z(n25767) );
  NANDN U33039 ( .A(x[3764]), .B(y[3764]), .Z(n25766) );
  NAND U33040 ( .A(n25767), .B(n25766), .Z(n56011) );
  OR U33041 ( .A(n15490), .B(n56011), .Z(n15491) );
  AND U33042 ( .A(n56012), .B(n15491), .Z(n15492) );
  NANDN U33043 ( .A(x[3765]), .B(y[3765]), .Z(n25765) );
  NANDN U33044 ( .A(x[3766]), .B(y[3766]), .Z(n25764) );
  NAND U33045 ( .A(n25765), .B(n25764), .Z(n56013) );
  OR U33046 ( .A(n15492), .B(n56013), .Z(n15493) );
  NAND U33047 ( .A(n51803), .B(n15493), .Z(n15494) );
  NANDN U33048 ( .A(n56014), .B(n15494), .Z(n15495) );
  NANDN U33049 ( .A(y[3768]), .B(x[3768]), .Z(n25761) );
  NANDN U33050 ( .A(y[3769]), .B(x[3769]), .Z(n25758) );
  AND U33051 ( .A(n25761), .B(n25758), .Z(n56015) );
  AND U33052 ( .A(n15495), .B(n56015), .Z(n15496) );
  NANDN U33053 ( .A(x[3769]), .B(y[3769]), .Z(n25759) );
  NANDN U33054 ( .A(x[3770]), .B(y[3770]), .Z(n39461) );
  NAND U33055 ( .A(n25759), .B(n39461), .Z(n51802) );
  OR U33056 ( .A(n15496), .B(n51802), .Z(n15497) );
  NAND U33057 ( .A(n51801), .B(n15497), .Z(n15498) );
  AND U33058 ( .A(n39465), .B(n15498), .Z(n15499) );
  NANDN U33059 ( .A(x[3771]), .B(y[3771]), .Z(n56016) );
  AND U33060 ( .A(n15499), .B(n56016), .Z(n15501) );
  NANDN U33061 ( .A(y[3772]), .B(x[3772]), .Z(n15500) );
  NANDN U33062 ( .A(y[3773]), .B(x[3773]), .Z(n39471) );
  NAND U33063 ( .A(n15500), .B(n39471), .Z(n51800) );
  OR U33064 ( .A(n15501), .B(n51800), .Z(n15502) );
  NANDN U33065 ( .A(x[3773]), .B(y[3773]), .Z(n25756) );
  NANDN U33066 ( .A(x[3774]), .B(y[3774]), .Z(n25755) );
  AND U33067 ( .A(n25756), .B(n25755), .Z(n51799) );
  AND U33068 ( .A(n15502), .B(n51799), .Z(n15503) );
  NANDN U33069 ( .A(y[3774]), .B(x[3774]), .Z(n39470) );
  NANDN U33070 ( .A(y[3775]), .B(x[3775]), .Z(n25753) );
  NAND U33071 ( .A(n39470), .B(n25753), .Z(n56019) );
  OR U33072 ( .A(n15503), .B(n56019), .Z(n15504) );
  NAND U33073 ( .A(n15505), .B(n15504), .Z(n15506) );
  NANDN U33074 ( .A(n56022), .B(n15506), .Z(n15507) );
  AND U33075 ( .A(n25752), .B(n15507), .Z(n15508) );
  NANDN U33076 ( .A(x[3777]), .B(y[3777]), .Z(n56023) );
  AND U33077 ( .A(n15508), .B(n56023), .Z(n15510) );
  NANDN U33078 ( .A(y[3778]), .B(x[3778]), .Z(n15509) );
  NANDN U33079 ( .A(y[3779]), .B(x[3779]), .Z(n39486) );
  NAND U33080 ( .A(n15509), .B(n39486), .Z(n56025) );
  OR U33081 ( .A(n15510), .B(n56025), .Z(n15511) );
  AND U33082 ( .A(n39485), .B(n15511), .Z(n15512) );
  ANDN U33083 ( .B(y[3779]), .A(x[3779]), .Z(n56026) );
  ANDN U33084 ( .B(n15512), .A(n56026), .Z(n15514) );
  NANDN U33085 ( .A(y[3780]), .B(x[3780]), .Z(n15513) );
  NANDN U33086 ( .A(y[3781]), .B(x[3781]), .Z(n39492) );
  NAND U33087 ( .A(n15513), .B(n39492), .Z(n56028) );
  OR U33088 ( .A(n15514), .B(n56028), .Z(n15515) );
  AND U33089 ( .A(n56029), .B(n15515), .Z(n15516) );
  OR U33090 ( .A(n56030), .B(n15516), .Z(n15517) );
  NAND U33091 ( .A(n56031), .B(n15517), .Z(n15518) );
  NANDN U33092 ( .A(n56032), .B(n15518), .Z(n15519) );
  AND U33093 ( .A(n56033), .B(n15519), .Z(n15520) );
  NANDN U33094 ( .A(y[3786]), .B(x[3786]), .Z(n25746) );
  NANDN U33095 ( .A(y[3787]), .B(x[3787]), .Z(n25742) );
  AND U33096 ( .A(n25746), .B(n25742), .Z(n56034) );
  NANDN U33097 ( .A(n15520), .B(n56034), .Z(n15521) );
  NANDN U33098 ( .A(n56036), .B(n15521), .Z(n15522) );
  AND U33099 ( .A(n56037), .B(n15522), .Z(n15523) );
  OR U33100 ( .A(n56038), .B(n15523), .Z(n15524) );
  NAND U33101 ( .A(n56039), .B(n15524), .Z(n15525) );
  NANDN U33102 ( .A(n56040), .B(n15525), .Z(n15526) );
  AND U33103 ( .A(n56041), .B(n15526), .Z(n15527) );
  NANDN U33104 ( .A(x[3793]), .B(y[3793]), .Z(n25736) );
  NANDN U33105 ( .A(x[3794]), .B(y[3794]), .Z(n39528) );
  NAND U33106 ( .A(n25736), .B(n39528), .Z(n56042) );
  OR U33107 ( .A(n15527), .B(n56042), .Z(n15528) );
  NAND U33108 ( .A(n56043), .B(n15528), .Z(n15529) );
  AND U33109 ( .A(n56044), .B(n15529), .Z(n15530) );
  NANDN U33110 ( .A(y[3796]), .B(x[3796]), .Z(n25732) );
  NANDN U33111 ( .A(y[3797]), .B(x[3797]), .Z(n25730) );
  AND U33112 ( .A(n25732), .B(n25730), .Z(n56045) );
  NANDN U33113 ( .A(n15530), .B(n56045), .Z(n15531) );
  NAND U33114 ( .A(n15532), .B(n15531), .Z(n15533) );
  AND U33115 ( .A(n56046), .B(n15533), .Z(n15535) );
  NANDN U33116 ( .A(x[3799]), .B(y[3799]), .Z(n56047) );
  ANDN U33117 ( .B(y[3800]), .A(x[3800]), .Z(n25726) );
  ANDN U33118 ( .B(n56047), .A(n25726), .Z(n15534) );
  NANDN U33119 ( .A(n15535), .B(n15534), .Z(n15536) );
  NANDN U33120 ( .A(n56048), .B(n15536), .Z(n15537) );
  AND U33121 ( .A(n56049), .B(n15537), .Z(n15538) );
  NANDN U33122 ( .A(x[3801]), .B(y[3801]), .Z(n25727) );
  NAND U33123 ( .A(n15538), .B(n25727), .Z(n15539) );
  NANDN U33124 ( .A(n56053), .B(n15539), .Z(n15540) );
  AND U33125 ( .A(n56054), .B(n15540), .Z(n15541) );
  NANDN U33126 ( .A(y[3804]), .B(x[3804]), .Z(n25723) );
  NANDN U33127 ( .A(y[3805]), .B(x[3805]), .Z(n39554) );
  NAND U33128 ( .A(n25723), .B(n39554), .Z(n56055) );
  OR U33129 ( .A(n15541), .B(n56055), .Z(n15542) );
  NAND U33130 ( .A(n51796), .B(n15542), .Z(n15543) );
  NANDN U33131 ( .A(n56056), .B(n15543), .Z(n15544) );
  NANDN U33132 ( .A(x[3807]), .B(y[3807]), .Z(n39557) );
  NANDN U33133 ( .A(x[3808]), .B(y[3808]), .Z(n39564) );
  AND U33134 ( .A(n39557), .B(n39564), .Z(n56057) );
  AND U33135 ( .A(n15544), .B(n56057), .Z(n15545) );
  NANDN U33136 ( .A(y[3808]), .B(x[3808]), .Z(n25721) );
  NANDN U33137 ( .A(y[3809]), .B(x[3809]), .Z(n25720) );
  NAND U33138 ( .A(n25721), .B(n25720), .Z(n51795) );
  OR U33139 ( .A(n15545), .B(n51795), .Z(n15546) );
  NANDN U33140 ( .A(x[3809]), .B(y[3809]), .Z(n39563) );
  NANDN U33141 ( .A(x[3810]), .B(y[3810]), .Z(n39570) );
  AND U33142 ( .A(n39563), .B(n39570), .Z(n51794) );
  AND U33143 ( .A(n15546), .B(n51794), .Z(n15547) );
  NANDN U33144 ( .A(y[3810]), .B(x[3810]), .Z(n25719) );
  NANDN U33145 ( .A(y[3811]), .B(x[3811]), .Z(n25718) );
  NAND U33146 ( .A(n25719), .B(n25718), .Z(n56058) );
  OR U33147 ( .A(n15547), .B(n56058), .Z(n15548) );
  NAND U33148 ( .A(n56059), .B(n15548), .Z(n15549) );
  NANDN U33149 ( .A(n56060), .B(n15549), .Z(n15550) );
  NANDN U33150 ( .A(x[3813]), .B(y[3813]), .Z(n39575) );
  NANDN U33151 ( .A(x[3814]), .B(y[3814]), .Z(n39584) );
  AND U33152 ( .A(n39575), .B(n39584), .Z(n56061) );
  AND U33153 ( .A(n15550), .B(n56061), .Z(n15551) );
  NANDN U33154 ( .A(y[3814]), .B(x[3814]), .Z(n25715) );
  ANDN U33155 ( .B(x[3815]), .A(y[3815]), .Z(n39588) );
  ANDN U33156 ( .B(n25715), .A(n39588), .Z(n56064) );
  NANDN U33157 ( .A(n15551), .B(n56064), .Z(n15552) );
  NANDN U33158 ( .A(n56065), .B(n15552), .Z(n15553) );
  AND U33159 ( .A(n56066), .B(n15553), .Z(n15554) );
  XNOR U33160 ( .A(y[3818]), .B(x[3818]), .Z(n25714) );
  NANDN U33161 ( .A(x[3817]), .B(y[3817]), .Z(n39590) );
  NAND U33162 ( .A(n25714), .B(n39590), .Z(n56067) );
  OR U33163 ( .A(n15554), .B(n56067), .Z(n15555) );
  NAND U33164 ( .A(n51793), .B(n15555), .Z(n15556) );
  NANDN U33165 ( .A(n56068), .B(n15556), .Z(n15558) );
  NANDN U33166 ( .A(y[3820]), .B(x[3820]), .Z(n15557) );
  NANDN U33167 ( .A(y[3821]), .B(x[3821]), .Z(n39603) );
  AND U33168 ( .A(n15557), .B(n39603), .Z(n56069) );
  AND U33169 ( .A(n15558), .B(n56069), .Z(n15559) );
  XNOR U33170 ( .A(y[3822]), .B(x[3822]), .Z(n39604) );
  NANDN U33171 ( .A(x[3821]), .B(y[3821]), .Z(n25709) );
  NAND U33172 ( .A(n39604), .B(n25709), .Z(n51792) );
  OR U33173 ( .A(n15559), .B(n51792), .Z(n15561) );
  NANDN U33174 ( .A(y[3822]), .B(x[3822]), .Z(n15560) );
  NANDN U33175 ( .A(y[3823]), .B(x[3823]), .Z(n39609) );
  AND U33176 ( .A(n15560), .B(n39609), .Z(n51791) );
  AND U33177 ( .A(n15561), .B(n51791), .Z(n15562) );
  XNOR U33178 ( .A(y[3824]), .B(x[3824]), .Z(n39610) );
  NANDN U33179 ( .A(x[3823]), .B(y[3823]), .Z(n25707) );
  NAND U33180 ( .A(n39610), .B(n25707), .Z(n56070) );
  OR U33181 ( .A(n15562), .B(n56070), .Z(n15563) );
  NAND U33182 ( .A(n56071), .B(n15563), .Z(n15564) );
  NANDN U33183 ( .A(n56072), .B(n15564), .Z(n15566) );
  NANDN U33184 ( .A(y[3826]), .B(x[3826]), .Z(n15565) );
  NANDN U33185 ( .A(y[3827]), .B(x[3827]), .Z(n39621) );
  AND U33186 ( .A(n15565), .B(n39621), .Z(n56075) );
  AND U33187 ( .A(n15566), .B(n56075), .Z(n15567) );
  XNOR U33188 ( .A(y[3828]), .B(x[3828]), .Z(n39622) );
  NANDN U33189 ( .A(x[3827]), .B(y[3827]), .Z(n25703) );
  NAND U33190 ( .A(n39622), .B(n25703), .Z(n51790) );
  OR U33191 ( .A(n15567), .B(n51790), .Z(n15568) );
  NAND U33192 ( .A(n51789), .B(n15568), .Z(n15569) );
  NANDN U33193 ( .A(n56076), .B(n15569), .Z(n15570) );
  NANDN U33194 ( .A(y[3830]), .B(x[3830]), .Z(n39627) );
  NANDN U33195 ( .A(y[3831]), .B(x[3831]), .Z(n25698) );
  AND U33196 ( .A(n39627), .B(n25698), .Z(n56077) );
  AND U33197 ( .A(n15570), .B(n56077), .Z(n15571) );
  ANDN U33198 ( .B(n15572), .A(n15571), .Z(n15574) );
  NANDN U33199 ( .A(y[3832]), .B(x[3832]), .Z(n15573) );
  NANDN U33200 ( .A(y[3833]), .B(x[3833]), .Z(n25696) );
  AND U33201 ( .A(n15573), .B(n25696), .Z(n56078) );
  NANDN U33202 ( .A(n15574), .B(n56078), .Z(n15575) );
  AND U33203 ( .A(n25697), .B(n15575), .Z(n15576) );
  NAND U33204 ( .A(n51786), .B(n15576), .Z(n15577) );
  NANDN U33205 ( .A(n56079), .B(n15577), .Z(n15578) );
  AND U33206 ( .A(n39642), .B(n15578), .Z(n15579) );
  NAND U33207 ( .A(n56080), .B(n15579), .Z(n15580) );
  NAND U33208 ( .A(n56084), .B(n15580), .Z(n15581) );
  NANDN U33209 ( .A(n56085), .B(n15581), .Z(n15582) );
  NAND U33210 ( .A(n56086), .B(n15582), .Z(n15583) );
  AND U33211 ( .A(n39654), .B(n15583), .Z(n15584) );
  NAND U33212 ( .A(n56088), .B(n15584), .Z(n15585) );
  NANDN U33213 ( .A(n56089), .B(n15585), .Z(n15586) );
  AND U33214 ( .A(n39660), .B(n15586), .Z(n15587) );
  NANDN U33215 ( .A(x[3841]), .B(y[3841]), .Z(n56090) );
  AND U33216 ( .A(n15587), .B(n56090), .Z(n15588) );
  ANDN U33217 ( .B(n51784), .A(n15588), .Z(n15589) );
  NANDN U33218 ( .A(x[3843]), .B(y[3843]), .Z(n39663) );
  NANDN U33219 ( .A(x[3844]), .B(y[3844]), .Z(n25691) );
  NAND U33220 ( .A(n39663), .B(n25691), .Z(n56092) );
  OR U33221 ( .A(n15589), .B(n56092), .Z(n15590) );
  NAND U33222 ( .A(n56093), .B(n15590), .Z(n15591) );
  NANDN U33223 ( .A(n51783), .B(n15591), .Z(n15592) );
  NANDN U33224 ( .A(y[3846]), .B(x[3846]), .Z(n25688) );
  NANDN U33225 ( .A(y[3847]), .B(x[3847]), .Z(n25687) );
  AND U33226 ( .A(n25688), .B(n25687), .Z(n51782) );
  AND U33227 ( .A(n15592), .B(n51782), .Z(n15593) );
  ANDN U33228 ( .B(y[3848]), .A(x[3848]), .Z(n39681) );
  NANDN U33229 ( .A(x[3847]), .B(y[3847]), .Z(n39673) );
  NANDN U33230 ( .A(n39681), .B(n39673), .Z(n56094) );
  OR U33231 ( .A(n15593), .B(n56094), .Z(n15594) );
  AND U33232 ( .A(n56097), .B(n15594), .Z(n15595) );
  NANDN U33233 ( .A(x[3849]), .B(y[3849]), .Z(n39679) );
  NANDN U33234 ( .A(x[3850]), .B(y[3850]), .Z(n25684) );
  NAND U33235 ( .A(n39679), .B(n25684), .Z(n56098) );
  OR U33236 ( .A(n15595), .B(n56098), .Z(n15596) );
  NAND U33237 ( .A(n56099), .B(n15596), .Z(n15597) );
  NANDN U33238 ( .A(n51781), .B(n15597), .Z(n15598) );
  NAND U33239 ( .A(n56100), .B(n15598), .Z(n15599) );
  AND U33240 ( .A(n25679), .B(n15599), .Z(n15600) );
  NANDN U33241 ( .A(n25680), .B(n15600), .Z(n15602) );
  NANDN U33242 ( .A(y[3854]), .B(x[3854]), .Z(n15601) );
  NANDN U33243 ( .A(y[3855]), .B(x[3855]), .Z(n39699) );
  AND U33244 ( .A(n15601), .B(n39699), .Z(n56103) );
  AND U33245 ( .A(n15602), .B(n56103), .Z(n15603) );
  ANDN U33246 ( .B(y[3855]), .A(x[3855]), .Z(n39696) );
  NANDN U33247 ( .A(x[3856]), .B(y[3856]), .Z(n25677) );
  NANDN U33248 ( .A(n39696), .B(n25677), .Z(n56104) );
  OR U33249 ( .A(n15603), .B(n56104), .Z(n15604) );
  NAND U33250 ( .A(n56105), .B(n15604), .Z(n15605) );
  NANDN U33251 ( .A(n51780), .B(n15605), .Z(n15606) );
  NANDN U33252 ( .A(y[3858]), .B(x[3858]), .Z(n39704) );
  NANDN U33253 ( .A(y[3859]), .B(x[3859]), .Z(n39711) );
  AND U33254 ( .A(n39704), .B(n39711), .Z(n51779) );
  AND U33255 ( .A(n15606), .B(n51779), .Z(n15607) );
  NANDN U33256 ( .A(x[3859]), .B(y[3859]), .Z(n25674) );
  NANDN U33257 ( .A(x[3860]), .B(y[3860]), .Z(n25673) );
  NAND U33258 ( .A(n25674), .B(n25673), .Z(n56107) );
  OR U33259 ( .A(n15607), .B(n56107), .Z(n15608) );
  AND U33260 ( .A(n56108), .B(n15608), .Z(n15609) );
  OR U33261 ( .A(n56109), .B(n15609), .Z(n15610) );
  NAND U33262 ( .A(n56110), .B(n15610), .Z(n15611) );
  NANDN U33263 ( .A(n56111), .B(n15611), .Z(n15612) );
  AND U33264 ( .A(n56112), .B(n15612), .Z(n15613) );
  NANDN U33265 ( .A(x[3865]), .B(y[3865]), .Z(n25668) );
  NANDN U33266 ( .A(x[3866]), .B(y[3866]), .Z(n39731) );
  AND U33267 ( .A(n25668), .B(n39731), .Z(n51778) );
  NANDN U33268 ( .A(n15613), .B(n51778), .Z(n15614) );
  NANDN U33269 ( .A(n56113), .B(n15614), .Z(n15615) );
  AND U33270 ( .A(n56114), .B(n15615), .Z(n15616) );
  NANDN U33271 ( .A(y[3868]), .B(x[3868]), .Z(n25664) );
  NANDN U33272 ( .A(y[3869]), .B(x[3869]), .Z(n25663) );
  NAND U33273 ( .A(n25664), .B(n25663), .Z(n56115) );
  OR U33274 ( .A(n15616), .B(n56115), .Z(n15617) );
  NAND U33275 ( .A(n56116), .B(n15617), .Z(n15618) );
  NANDN U33276 ( .A(n51777), .B(n15618), .Z(n15619) );
  NANDN U33277 ( .A(x[3871]), .B(y[3871]), .Z(n25660) );
  NANDN U33278 ( .A(x[3872]), .B(y[3872]), .Z(n39747) );
  AND U33279 ( .A(n25660), .B(n39747), .Z(n51776) );
  AND U33280 ( .A(n15619), .B(n51776), .Z(n15620) );
  NANDN U33281 ( .A(y[3872]), .B(x[3872]), .Z(n39744) );
  NANDN U33282 ( .A(y[3873]), .B(x[3873]), .Z(n39750) );
  AND U33283 ( .A(n39744), .B(n39750), .Z(n56119) );
  NANDN U33284 ( .A(n15620), .B(n56119), .Z(n15621) );
  AND U33285 ( .A(n39751), .B(n15621), .Z(n15622) );
  NANDN U33286 ( .A(x[3873]), .B(y[3873]), .Z(n56121) );
  AND U33287 ( .A(n15622), .B(n56121), .Z(n15623) );
  OR U33288 ( .A(n56122), .B(n15623), .Z(n15624) );
  NAND U33289 ( .A(n56123), .B(n15624), .Z(n15625) );
  NANDN U33290 ( .A(n56124), .B(n15625), .Z(n15626) );
  AND U33291 ( .A(n25654), .B(n15626), .Z(n15627) );
  NANDN U33292 ( .A(n25655), .B(n15627), .Z(n15628) );
  NAND U33293 ( .A(n56125), .B(n15628), .Z(n15629) );
  NAND U33294 ( .A(n39765), .B(n15629), .Z(n15630) );
  ANDN U33295 ( .B(y[3879]), .A(x[3879]), .Z(n56127) );
  OR U33296 ( .A(n15630), .B(n56127), .Z(n15631) );
  NAND U33297 ( .A(n51773), .B(n15631), .Z(n15633) );
  XNOR U33298 ( .A(x[3882]), .B(y[3882]), .Z(n39771) );
  NANDN U33299 ( .A(x[3881]), .B(y[3881]), .Z(n56128) );
  NAND U33300 ( .A(n39771), .B(n56128), .Z(n15632) );
  ANDN U33301 ( .B(n15633), .A(n15632), .Z(n15634) );
  OR U33302 ( .A(n56130), .B(n15634), .Z(n15635) );
  NAND U33303 ( .A(n56131), .B(n15635), .Z(n15636) );
  NANDN U33304 ( .A(n56132), .B(n15636), .Z(n15637) );
  AND U33305 ( .A(n56134), .B(n15637), .Z(n15638) );
  NANDN U33306 ( .A(y[3886]), .B(x[3886]), .Z(n25647) );
  NANDN U33307 ( .A(y[3887]), .B(x[3887]), .Z(n39784) );
  NAND U33308 ( .A(n25647), .B(n39784), .Z(n56135) );
  OR U33309 ( .A(n15638), .B(n56135), .Z(n15639) );
  AND U33310 ( .A(n15640), .B(n15639), .Z(n15641) );
  OR U33311 ( .A(n56138), .B(n15641), .Z(n15642) );
  NAND U33312 ( .A(n56139), .B(n15642), .Z(n15643) );
  NANDN U33313 ( .A(n56140), .B(n15643), .Z(n15644) );
  AND U33314 ( .A(n56141), .B(n15644), .Z(n15645) );
  NANDN U33315 ( .A(y[3892]), .B(x[3892]), .Z(n25639) );
  NANDN U33316 ( .A(y[3893]), .B(x[3893]), .Z(n25638) );
  AND U33317 ( .A(n25639), .B(n25638), .Z(n51772) );
  NANDN U33318 ( .A(n15645), .B(n51772), .Z(n15646) );
  NANDN U33319 ( .A(n56142), .B(n15646), .Z(n15647) );
  NANDN U33320 ( .A(y[3894]), .B(x[3894]), .Z(n25637) );
  NANDN U33321 ( .A(y[3895]), .B(x[3895]), .Z(n25636) );
  AND U33322 ( .A(n25637), .B(n25636), .Z(n56143) );
  AND U33323 ( .A(n15647), .B(n56143), .Z(n15648) );
  ANDN U33324 ( .B(y[3895]), .A(x[3895]), .Z(n39803) );
  ANDN U33325 ( .B(y[3896]), .A(x[3896]), .Z(n39812) );
  OR U33326 ( .A(n39803), .B(n39812), .Z(n56144) );
  OR U33327 ( .A(n15648), .B(n56144), .Z(n15649) );
  NAND U33328 ( .A(n56145), .B(n15649), .Z(n15650) );
  NANDN U33329 ( .A(n51771), .B(n15650), .Z(n15651) );
  NANDN U33330 ( .A(y[3898]), .B(x[3898]), .Z(n25633) );
  NANDN U33331 ( .A(y[3899]), .B(x[3899]), .Z(n39820) );
  AND U33332 ( .A(n25633), .B(n39820), .Z(n51770) );
  AND U33333 ( .A(n15651), .B(n51770), .Z(n15652) );
  NANDN U33334 ( .A(x[3899]), .B(y[3899]), .Z(n25631) );
  NANDN U33335 ( .A(x[3900]), .B(y[3900]), .Z(n39822) );
  NAND U33336 ( .A(n25631), .B(n39822), .Z(n56147) );
  OR U33337 ( .A(n15652), .B(n56147), .Z(n15653) );
  AND U33338 ( .A(n56148), .B(n15653), .Z(n15654) );
  OR U33339 ( .A(n56149), .B(n15654), .Z(n15655) );
  NAND U33340 ( .A(n56150), .B(n15655), .Z(n15656) );
  NANDN U33341 ( .A(n56151), .B(n15656), .Z(n15657) );
  AND U33342 ( .A(n56152), .B(n15657), .Z(n15658) );
  OR U33343 ( .A(n56153), .B(n15658), .Z(n15659) );
  NAND U33344 ( .A(n56154), .B(n15659), .Z(n15660) );
  NANDN U33345 ( .A(n51769), .B(n15660), .Z(n15661) );
  NANDN U33346 ( .A(y[3908]), .B(x[3908]), .Z(n39843) );
  NANDN U33347 ( .A(y[3909]), .B(x[3909]), .Z(n39850) );
  AND U33348 ( .A(n39843), .B(n39850), .Z(n51768) );
  AND U33349 ( .A(n15661), .B(n51768), .Z(n15663) );
  NANDN U33350 ( .A(x[3909]), .B(y[3909]), .Z(n25623) );
  XNOR U33351 ( .A(y[3910]), .B(x[3910]), .Z(n15662) );
  NAND U33352 ( .A(n25623), .B(n15662), .Z(n56155) );
  OR U33353 ( .A(n15663), .B(n56155), .Z(n15664) );
  AND U33354 ( .A(n56156), .B(n15664), .Z(n15665) );
  NANDN U33355 ( .A(x[3911]), .B(y[3911]), .Z(n25621) );
  NANDN U33356 ( .A(x[3912]), .B(y[3912]), .Z(n25620) );
  NAND U33357 ( .A(n25621), .B(n25620), .Z(n51767) );
  OR U33358 ( .A(n15665), .B(n51767), .Z(n15666) );
  NAND U33359 ( .A(n51766), .B(n15666), .Z(n15667) );
  NANDN U33360 ( .A(n56159), .B(n15667), .Z(n15668) );
  NANDN U33361 ( .A(y[3914]), .B(x[3914]), .Z(n25617) );
  NANDN U33362 ( .A(y[3915]), .B(x[3915]), .Z(n39867) );
  AND U33363 ( .A(n25617), .B(n39867), .Z(n56160) );
  AND U33364 ( .A(n15668), .B(n56160), .Z(n15669) );
  NANDN U33365 ( .A(x[3915]), .B(y[3915]), .Z(n25615) );
  NANDN U33366 ( .A(x[3916]), .B(y[3916]), .Z(n25614) );
  AND U33367 ( .A(n25615), .B(n25614), .Z(n56161) );
  NANDN U33368 ( .A(n15669), .B(n56161), .Z(n15670) );
  NANDN U33369 ( .A(n56162), .B(n15670), .Z(n15671) );
  AND U33370 ( .A(n56163), .B(n15671), .Z(n15672) );
  OR U33371 ( .A(n56164), .B(n15672), .Z(n15673) );
  NAND U33372 ( .A(n56165), .B(n15673), .Z(n15674) );
  NANDN U33373 ( .A(n56166), .B(n15674), .Z(n15675) );
  NANDN U33374 ( .A(x[3921]), .B(y[3921]), .Z(n39881) );
  NANDN U33375 ( .A(x[3922]), .B(y[3922]), .Z(n39888) );
  AND U33376 ( .A(n39881), .B(n39888), .Z(n51765) );
  AND U33377 ( .A(n15675), .B(n51765), .Z(n15676) );
  NANDN U33378 ( .A(y[3922]), .B(x[3922]), .Z(n25609) );
  NANDN U33379 ( .A(y[3923]), .B(x[3923]), .Z(n25608) );
  NAND U33380 ( .A(n25609), .B(n25608), .Z(n56167) );
  OR U33381 ( .A(n15676), .B(n56167), .Z(n15677) );
  NANDN U33382 ( .A(x[3923]), .B(y[3923]), .Z(n39887) );
  NANDN U33383 ( .A(x[3924]), .B(y[3924]), .Z(n39894) );
  AND U33384 ( .A(n39887), .B(n39894), .Z(n56168) );
  AND U33385 ( .A(n15677), .B(n56168), .Z(n15678) );
  NANDN U33386 ( .A(y[3924]), .B(x[3924]), .Z(n25607) );
  NANDN U33387 ( .A(y[3925]), .B(x[3925]), .Z(n25606) );
  NAND U33388 ( .A(n25607), .B(n25606), .Z(n51764) );
  OR U33389 ( .A(n15678), .B(n51764), .Z(n15679) );
  NAND U33390 ( .A(n51763), .B(n15679), .Z(n15680) );
  NANDN U33391 ( .A(n56171), .B(n15680), .Z(n15681) );
  NANDN U33392 ( .A(x[3927]), .B(y[3927]), .Z(n39899) );
  NANDN U33393 ( .A(x[3928]), .B(y[3928]), .Z(n25602) );
  AND U33394 ( .A(n39899), .B(n25602), .Z(n56173) );
  AND U33395 ( .A(n15681), .B(n56173), .Z(n15682) );
  NANDN U33396 ( .A(y[3928]), .B(x[3928]), .Z(n25603) );
  NANDN U33397 ( .A(y[3929]), .B(x[3929]), .Z(n25599) );
  AND U33398 ( .A(n25603), .B(n25599), .Z(n56174) );
  NANDN U33399 ( .A(n15682), .B(n56174), .Z(n15683) );
  NAND U33400 ( .A(n56175), .B(n15683), .Z(n15684) );
  NANDN U33401 ( .A(n56176), .B(n15684), .Z(n15685) );
  AND U33402 ( .A(n39913), .B(n15685), .Z(n15686) );
  NAND U33403 ( .A(n51761), .B(n15686), .Z(n15687) );
  NANDN U33404 ( .A(n56177), .B(n15687), .Z(n15688) );
  AND U33405 ( .A(n39918), .B(n15688), .Z(n15689) );
  NANDN U33406 ( .A(x[3933]), .B(y[3933]), .Z(n56178) );
  AND U33407 ( .A(n15689), .B(n56178), .Z(n15691) );
  NANDN U33408 ( .A(y[3934]), .B(x[3934]), .Z(n15690) );
  NANDN U33409 ( .A(y[3935]), .B(x[3935]), .Z(n25597) );
  NAND U33410 ( .A(n15690), .B(n25597), .Z(n56180) );
  OR U33411 ( .A(n15691), .B(n56180), .Z(n15692) );
  NANDN U33412 ( .A(x[3935]), .B(y[3935]), .Z(n39921) );
  NANDN U33413 ( .A(x[3936]), .B(y[3936]), .Z(n25595) );
  AND U33414 ( .A(n39921), .B(n25595), .Z(n56181) );
  AND U33415 ( .A(n15692), .B(n56181), .Z(n15693) );
  NANDN U33416 ( .A(y[3936]), .B(x[3936]), .Z(n25596) );
  NANDN U33417 ( .A(y[3937]), .B(x[3937]), .Z(n25593) );
  NAND U33418 ( .A(n25596), .B(n25593), .Z(n51760) );
  OR U33419 ( .A(n15693), .B(n51760), .Z(n15694) );
  NAND U33420 ( .A(n51759), .B(n15694), .Z(n15695) );
  NANDN U33421 ( .A(n56184), .B(n15695), .Z(n15696) );
  NANDN U33422 ( .A(x[3939]), .B(y[3939]), .Z(n39931) );
  NANDN U33423 ( .A(x[3940]), .B(y[3940]), .Z(n39938) );
  AND U33424 ( .A(n39931), .B(n39938), .Z(n56185) );
  AND U33425 ( .A(n15696), .B(n56185), .Z(n15697) );
  NANDN U33426 ( .A(y[3940]), .B(x[3940]), .Z(n25590) );
  NANDN U33427 ( .A(y[3941]), .B(x[3941]), .Z(n25589) );
  AND U33428 ( .A(n25590), .B(n25589), .Z(n56186) );
  NANDN U33429 ( .A(n15697), .B(n56186), .Z(n15698) );
  NANDN U33430 ( .A(n56187), .B(n15698), .Z(n15699) );
  AND U33431 ( .A(n56188), .B(n15699), .Z(n15700) );
  OR U33432 ( .A(n56189), .B(n15700), .Z(n15701) );
  NAND U33433 ( .A(n56190), .B(n15701), .Z(n15702) );
  NANDN U33434 ( .A(n51758), .B(n15702), .Z(n15703) );
  NANDN U33435 ( .A(y[3946]), .B(x[3946]), .Z(n25582) );
  NANDN U33436 ( .A(y[3947]), .B(x[3947]), .Z(n25581) );
  AND U33437 ( .A(n25582), .B(n25581), .Z(n51757) );
  AND U33438 ( .A(n15703), .B(n51757), .Z(n15705) );
  ANDN U33439 ( .B(y[3947]), .A(x[3947]), .Z(n39953) );
  XNOR U33440 ( .A(y[3948]), .B(x[3948]), .Z(n15704) );
  NANDN U33441 ( .A(n39953), .B(n15704), .Z(n56191) );
  OR U33442 ( .A(n15705), .B(n56191), .Z(n15706) );
  NAND U33443 ( .A(n56192), .B(n15706), .Z(n15707) );
  NANDN U33444 ( .A(n51756), .B(n15707), .Z(n15708) );
  NANDN U33445 ( .A(y[3950]), .B(x[3950]), .Z(n25576) );
  NANDN U33446 ( .A(y[3951]), .B(x[3951]), .Z(n25572) );
  AND U33447 ( .A(n25576), .B(n25572), .Z(n51755) );
  AND U33448 ( .A(n15708), .B(n51755), .Z(n15709) );
  NOR U33449 ( .A(n25574), .B(n15709), .Z(n15710) );
  NAND U33450 ( .A(n15711), .B(n15710), .Z(n15712) );
  AND U33451 ( .A(n56195), .B(n15712), .Z(n15714) );
  NANDN U33452 ( .A(x[3954]), .B(y[3954]), .Z(n51754) );
  ANDN U33453 ( .B(y[3953]), .A(x[3953]), .Z(n25571) );
  ANDN U33454 ( .B(n51754), .A(n25571), .Z(n15713) );
  NANDN U33455 ( .A(n15714), .B(n15713), .Z(n15715) );
  NANDN U33456 ( .A(n56196), .B(n15715), .Z(n15716) );
  AND U33457 ( .A(n56197), .B(n15716), .Z(n15717) );
  OR U33458 ( .A(n56198), .B(n15717), .Z(n15718) );
  AND U33459 ( .A(n15719), .B(n15718), .Z(n15720) );
  OR U33460 ( .A(n56201), .B(n15720), .Z(n15721) );
  NAND U33461 ( .A(n56202), .B(n15721), .Z(n15722) );
  NANDN U33462 ( .A(n56203), .B(n15722), .Z(n15723) );
  AND U33463 ( .A(n56204), .B(n15723), .Z(n15724) );
  OR U33464 ( .A(n56205), .B(n15724), .Z(n15725) );
  AND U33465 ( .A(n15726), .B(n15725), .Z(n15727) );
  OR U33466 ( .A(n56210), .B(n15727), .Z(n15728) );
  NAND U33467 ( .A(n56211), .B(n15728), .Z(n15729) );
  NANDN U33468 ( .A(n56212), .B(n15729), .Z(n15730) );
  AND U33469 ( .A(n56213), .B(n15730), .Z(n15731) );
  NANDN U33470 ( .A(y[3968]), .B(x[3968]), .Z(n40004) );
  NANDN U33471 ( .A(y[3969]), .B(x[3969]), .Z(n40011) );
  NAND U33472 ( .A(n40004), .B(n40011), .Z(n56214) );
  OR U33473 ( .A(n15731), .B(n56214), .Z(n15732) );
  NAND U33474 ( .A(n56215), .B(n15732), .Z(n15734) );
  NANDN U33475 ( .A(y[3970]), .B(x[3970]), .Z(n15733) );
  NANDN U33476 ( .A(y[3971]), .B(x[3971]), .Z(n25554) );
  AND U33477 ( .A(n15733), .B(n25554), .Z(n56216) );
  AND U33478 ( .A(n15734), .B(n56216), .Z(n15736) );
  NANDN U33479 ( .A(x[3971]), .B(y[3971]), .Z(n25555) );
  XNOR U33480 ( .A(x[3972]), .B(y[3972]), .Z(n15735) );
  NAND U33481 ( .A(n25555), .B(n15735), .Z(n56217) );
  OR U33482 ( .A(n15736), .B(n56217), .Z(n15737) );
  NANDN U33483 ( .A(y[3972]), .B(x[3972]), .Z(n25553) );
  NANDN U33484 ( .A(y[3973]), .B(x[3973]), .Z(n25549) );
  AND U33485 ( .A(n25553), .B(n25549), .Z(n56218) );
  AND U33486 ( .A(n15737), .B(n56218), .Z(n15738) );
  XNOR U33487 ( .A(y[3974]), .B(x[3974]), .Z(n25550) );
  NANDN U33488 ( .A(x[3973]), .B(y[3973]), .Z(n25552) );
  NAND U33489 ( .A(n25550), .B(n25552), .Z(n51751) );
  OR U33490 ( .A(n15738), .B(n51751), .Z(n15739) );
  NAND U33491 ( .A(n51750), .B(n15739), .Z(n15740) );
  NANDN U33492 ( .A(n56219), .B(n15740), .Z(n15741) );
  AND U33493 ( .A(n56220), .B(n15741), .Z(n15742) );
  NANDN U33494 ( .A(x[3977]), .B(y[3977]), .Z(n25547) );
  NANDN U33495 ( .A(x[3978]), .B(y[3978]), .Z(n25546) );
  AND U33496 ( .A(n25547), .B(n25546), .Z(n51749) );
  NANDN U33497 ( .A(n15742), .B(n51749), .Z(n15743) );
  NANDN U33498 ( .A(n56223), .B(n15743), .Z(n15744) );
  XNOR U33499 ( .A(y[3980]), .B(x[3980]), .Z(n40040) );
  NANDN U33500 ( .A(x[3979]), .B(y[3979]), .Z(n25545) );
  AND U33501 ( .A(n40040), .B(n25545), .Z(n56224) );
  AND U33502 ( .A(n15744), .B(n56224), .Z(n15746) );
  NANDN U33503 ( .A(y[3980]), .B(x[3980]), .Z(n15745) );
  NANDN U33504 ( .A(y[3981]), .B(x[3981]), .Z(n40047) );
  NAND U33505 ( .A(n15745), .B(n40047), .Z(n51748) );
  OR U33506 ( .A(n15746), .B(n51748), .Z(n15747) );
  NAND U33507 ( .A(n51747), .B(n15747), .Z(n15748) );
  NANDN U33508 ( .A(n56225), .B(n15748), .Z(n15749) );
  AND U33509 ( .A(n25541), .B(n15749), .Z(n15750) );
  NANDN U33510 ( .A(x[3983]), .B(y[3983]), .Z(n56227) );
  AND U33511 ( .A(n15750), .B(n56227), .Z(n15752) );
  NANDN U33512 ( .A(y[3984]), .B(x[3984]), .Z(n15751) );
  NANDN U33513 ( .A(y[3985]), .B(x[3985]), .Z(n25539) );
  NAND U33514 ( .A(n15751), .B(n25539), .Z(n56228) );
  OR U33515 ( .A(n15752), .B(n56228), .Z(n15753) );
  AND U33516 ( .A(n56229), .B(n15753), .Z(n15754) );
  NANDN U33517 ( .A(y[3986]), .B(x[3986]), .Z(n25538) );
  NANDN U33518 ( .A(y[3987]), .B(x[3987]), .Z(n25536) );
  AND U33519 ( .A(n25538), .B(n25536), .Z(n56230) );
  NANDN U33520 ( .A(n15754), .B(n56230), .Z(n15755) );
  AND U33521 ( .A(n25537), .B(n15755), .Z(n15756) );
  NANDN U33522 ( .A(x[3987]), .B(y[3987]), .Z(n51745) );
  AND U33523 ( .A(n15756), .B(n51745), .Z(n15757) );
  OR U33524 ( .A(n56232), .B(n15757), .Z(n15758) );
  NAND U33525 ( .A(n56233), .B(n15758), .Z(n15759) );
  NANDN U33526 ( .A(n56234), .B(n15759), .Z(n15760) );
  AND U33527 ( .A(n25532), .B(n15760), .Z(n15761) );
  NANDN U33528 ( .A(x[3991]), .B(y[3991]), .Z(n56235) );
  AND U33529 ( .A(n15761), .B(n56235), .Z(n15762) );
  OR U33530 ( .A(n56237), .B(n15762), .Z(n15763) );
  AND U33531 ( .A(n15764), .B(n15763), .Z(n15765) );
  OR U33532 ( .A(n56238), .B(n15765), .Z(n15766) );
  NAND U33533 ( .A(n56239), .B(n15766), .Z(n15767) );
  NANDN U33534 ( .A(n56240), .B(n15767), .Z(n15768) );
  AND U33535 ( .A(n25526), .B(n15768), .Z(n15769) );
  NANDN U33536 ( .A(x[3997]), .B(y[3997]), .Z(n56241) );
  AND U33537 ( .A(n15769), .B(n56241), .Z(n15771) );
  ANDN U33538 ( .B(x[3999]), .A(y[3999]), .Z(n40090) );
  NANDN U33539 ( .A(y[3998]), .B(x[3998]), .Z(n15770) );
  NANDN U33540 ( .A(n40090), .B(n15770), .Z(n56243) );
  OR U33541 ( .A(n15771), .B(n56243), .Z(n15772) );
  XOR U33542 ( .A(x[4000]), .B(y[4000]), .Z(n40089) );
  ANDN U33543 ( .B(n15772), .A(n40089), .Z(n15773) );
  NANDN U33544 ( .A(x[3999]), .B(y[3999]), .Z(n51741) );
  AND U33545 ( .A(n15773), .B(n51741), .Z(n15775) );
  NANDN U33546 ( .A(y[4000]), .B(x[4000]), .Z(n15774) );
  NANDN U33547 ( .A(y[4001]), .B(x[4001]), .Z(n25523) );
  NAND U33548 ( .A(n15774), .B(n25523), .Z(n56244) );
  OR U33549 ( .A(n15775), .B(n56244), .Z(n15776) );
  AND U33550 ( .A(n15777), .B(n15776), .Z(n15779) );
  NANDN U33551 ( .A(y[4002]), .B(x[4002]), .Z(n15778) );
  NANDN U33552 ( .A(y[4003]), .B(x[4003]), .Z(n25522) );
  NAND U33553 ( .A(n15778), .B(n25522), .Z(n56249) );
  OR U33554 ( .A(n15779), .B(n56249), .Z(n15780) );
  NAND U33555 ( .A(n56251), .B(n15780), .Z(n15781) );
  NANDN U33556 ( .A(n51740), .B(n15781), .Z(n15782) );
  NANDN U33557 ( .A(x[4005]), .B(y[4005]), .Z(n25519) );
  NANDN U33558 ( .A(x[4006]), .B(y[4006]), .Z(n40107) );
  AND U33559 ( .A(n25519), .B(n40107), .Z(n51739) );
  AND U33560 ( .A(n15782), .B(n51739), .Z(n15783) );
  NANDN U33561 ( .A(y[4006]), .B(x[4006]), .Z(n25517) );
  NANDN U33562 ( .A(y[4007]), .B(x[4007]), .Z(n25516) );
  NAND U33563 ( .A(n25517), .B(n25516), .Z(n56252) );
  OR U33564 ( .A(n15783), .B(n56252), .Z(n15785) );
  NANDN U33565 ( .A(x[4007]), .B(y[4007]), .Z(n40106) );
  XNOR U33566 ( .A(x[4008]), .B(y[4008]), .Z(n15784) );
  AND U33567 ( .A(n40106), .B(n15784), .Z(n56253) );
  AND U33568 ( .A(n15785), .B(n56253), .Z(n15786) );
  NANDN U33569 ( .A(y[4008]), .B(x[4008]), .Z(n25515) );
  NANDN U33570 ( .A(y[4009]), .B(x[4009]), .Z(n25514) );
  NAND U33571 ( .A(n25515), .B(n25514), .Z(n56254) );
  OR U33572 ( .A(n15786), .B(n56254), .Z(n15787) );
  NAND U33573 ( .A(n56255), .B(n15787), .Z(n15788) );
  NANDN U33574 ( .A(n56256), .B(n15788), .Z(n15789) );
  AND U33575 ( .A(n56257), .B(n15789), .Z(n15790) );
  NANDN U33576 ( .A(y[4012]), .B(x[4012]), .Z(n25511) );
  NANDN U33577 ( .A(y[4013]), .B(x[4013]), .Z(n40127) );
  NAND U33578 ( .A(n25511), .B(n40127), .Z(n56258) );
  OR U33579 ( .A(n15790), .B(n56258), .Z(n15791) );
  NAND U33580 ( .A(n56259), .B(n15791), .Z(n15792) );
  NANDN U33581 ( .A(n51738), .B(n15792), .Z(n15793) );
  NAND U33582 ( .A(n51737), .B(n15793), .Z(n15794) );
  NAND U33583 ( .A(n56262), .B(n15794), .Z(n15795) );
  NANDN U33584 ( .A(n56263), .B(n15795), .Z(n15796) );
  AND U33585 ( .A(n56264), .B(n15796), .Z(n15797) );
  NANDN U33586 ( .A(x[4019]), .B(y[4019]), .Z(n25505) );
  NANDN U33587 ( .A(x[4020]), .B(y[4020]), .Z(n25504) );
  AND U33588 ( .A(n25505), .B(n25504), .Z(n56265) );
  NANDN U33589 ( .A(n15797), .B(n56265), .Z(n15798) );
  NANDN U33590 ( .A(n51736), .B(n15798), .Z(n15799) );
  NANDN U33591 ( .A(x[4021]), .B(y[4021]), .Z(n25503) );
  NANDN U33592 ( .A(x[4022]), .B(y[4022]), .Z(n25502) );
  AND U33593 ( .A(n25503), .B(n25502), .Z(n51735) );
  AND U33594 ( .A(n15799), .B(n51735), .Z(n15800) );
  NANDN U33595 ( .A(y[4022]), .B(x[4022]), .Z(n40151) );
  NANDN U33596 ( .A(y[4023]), .B(x[4023]), .Z(n40158) );
  NAND U33597 ( .A(n40151), .B(n40158), .Z(n56266) );
  OR U33598 ( .A(n15800), .B(n56266), .Z(n15801) );
  NAND U33599 ( .A(n56267), .B(n15801), .Z(n15802) );
  NANDN U33600 ( .A(n51734), .B(n15802), .Z(n15803) );
  NAND U33601 ( .A(n51733), .B(n15803), .Z(n15804) );
  NAND U33602 ( .A(n56270), .B(n15804), .Z(n15805) );
  NAND U33603 ( .A(n56273), .B(n15805), .Z(n15806) );
  ANDN U33604 ( .B(n25497), .A(n15806), .Z(n15807) );
  OR U33605 ( .A(n56274), .B(n15807), .Z(n15808) );
  NAND U33606 ( .A(n56275), .B(n15808), .Z(n15809) );
  NANDN U33607 ( .A(n51732), .B(n15809), .Z(n15810) );
  AND U33608 ( .A(n40178), .B(n15810), .Z(n15811) );
  NANDN U33609 ( .A(x[4031]), .B(y[4031]), .Z(n51731) );
  AND U33610 ( .A(n15811), .B(n51731), .Z(n15813) );
  NANDN U33611 ( .A(y[4032]), .B(x[4032]), .Z(n15812) );
  NANDN U33612 ( .A(y[4033]), .B(x[4033]), .Z(n40183) );
  NAND U33613 ( .A(n15812), .B(n40183), .Z(n56277) );
  OR U33614 ( .A(n15813), .B(n56277), .Z(n15814) );
  AND U33615 ( .A(n15815), .B(n15814), .Z(n15817) );
  NANDN U33616 ( .A(y[4034]), .B(x[4034]), .Z(n15816) );
  NANDN U33617 ( .A(y[4035]), .B(x[4035]), .Z(n40190) );
  NAND U33618 ( .A(n15816), .B(n40190), .Z(n56280) );
  OR U33619 ( .A(n15817), .B(n56280), .Z(n15818) );
  NAND U33620 ( .A(n56281), .B(n15818), .Z(n15819) );
  NANDN U33621 ( .A(n51730), .B(n15819), .Z(n15820) );
  NANDN U33622 ( .A(x[4037]), .B(y[4037]), .Z(n25489) );
  NANDN U33623 ( .A(x[4038]), .B(y[4038]), .Z(n25488) );
  AND U33624 ( .A(n25489), .B(n25488), .Z(n51729) );
  AND U33625 ( .A(n15820), .B(n51729), .Z(n15821) );
  NANDN U33626 ( .A(y[4038]), .B(x[4038]), .Z(n40198) );
  NANDN U33627 ( .A(y[4039]), .B(x[4039]), .Z(n25486) );
  NAND U33628 ( .A(n40198), .B(n25486), .Z(n51728) );
  OR U33629 ( .A(n15821), .B(n51728), .Z(n15822) );
  AND U33630 ( .A(n56283), .B(n15822), .Z(n15823) );
  NANDN U33631 ( .A(y[4040]), .B(x[4040]), .Z(n25485) );
  NANDN U33632 ( .A(y[4041]), .B(x[4041]), .Z(n40207) );
  NAND U33633 ( .A(n25485), .B(n40207), .Z(n51727) );
  OR U33634 ( .A(n15823), .B(n51727), .Z(n15824) );
  NAND U33635 ( .A(n56284), .B(n15824), .Z(n15825) );
  NANDN U33636 ( .A(n51726), .B(n15825), .Z(n15826) );
  NANDN U33637 ( .A(x[4043]), .B(y[4043]), .Z(n25481) );
  NANDN U33638 ( .A(x[4044]), .B(y[4044]), .Z(n25480) );
  AND U33639 ( .A(n25481), .B(n25480), .Z(n51725) );
  AND U33640 ( .A(n15826), .B(n51725), .Z(n15827) );
  NANDN U33641 ( .A(y[4044]), .B(x[4044]), .Z(n40212) );
  NANDN U33642 ( .A(y[4045]), .B(x[4045]), .Z(n40219) );
  AND U33643 ( .A(n40212), .B(n40219), .Z(n56285) );
  NANDN U33644 ( .A(n15827), .B(n56285), .Z(n15828) );
  NANDN U33645 ( .A(n56286), .B(n15828), .Z(n15829) );
  AND U33646 ( .A(n56287), .B(n15829), .Z(n15830) );
  OR U33647 ( .A(n56288), .B(n15830), .Z(n15831) );
  NAND U33648 ( .A(n56289), .B(n15831), .Z(n15832) );
  NANDN U33649 ( .A(n56291), .B(n15832), .Z(n15833) );
  AND U33650 ( .A(n56292), .B(n15833), .Z(n15835) );
  NANDN U33651 ( .A(x[4051]), .B(y[4051]), .Z(n40232) );
  XNOR U33652 ( .A(y[4052]), .B(x[4052]), .Z(n15834) );
  NAND U33653 ( .A(n40232), .B(n15834), .Z(n56293) );
  OR U33654 ( .A(n15835), .B(n56293), .Z(n15836) );
  NANDN U33655 ( .A(y[4052]), .B(x[4052]), .Z(n25471) );
  NANDN U33656 ( .A(y[4053]), .B(x[4053]), .Z(n25470) );
  AND U33657 ( .A(n25471), .B(n25470), .Z(n51724) );
  AND U33658 ( .A(n15836), .B(n51724), .Z(n15837) );
  NANDN U33659 ( .A(x[4053]), .B(y[4053]), .Z(n40238) );
  NANDN U33660 ( .A(x[4054]), .B(y[4054]), .Z(n40245) );
  NAND U33661 ( .A(n40238), .B(n40245), .Z(n56294) );
  OR U33662 ( .A(n15837), .B(n56294), .Z(n15838) );
  NAND U33663 ( .A(n56295), .B(n15838), .Z(n15839) );
  NANDN U33664 ( .A(n51723), .B(n15839), .Z(n15840) );
  NANDN U33665 ( .A(y[4056]), .B(x[4056]), .Z(n40247) );
  NANDN U33666 ( .A(y[4057]), .B(x[4057]), .Z(n40254) );
  AND U33667 ( .A(n40247), .B(n40254), .Z(n51722) );
  AND U33668 ( .A(n15840), .B(n51722), .Z(n15841) );
  NANDN U33669 ( .A(x[4057]), .B(y[4057]), .Z(n25467) );
  NANDN U33670 ( .A(x[4058]), .B(y[4058]), .Z(n40259) );
  AND U33671 ( .A(n25467), .B(n40259), .Z(n56296) );
  NANDN U33672 ( .A(n15841), .B(n56296), .Z(n15842) );
  NANDN U33673 ( .A(n56297), .B(n15842), .Z(n15843) );
  AND U33674 ( .A(n56298), .B(n15843), .Z(n15844) );
  OR U33675 ( .A(n56299), .B(n15844), .Z(n15845) );
  NAND U33676 ( .A(n56300), .B(n15845), .Z(n15846) );
  NANDN U33677 ( .A(n56301), .B(n15846), .Z(n15847) );
  AND U33678 ( .A(n56303), .B(n15847), .Z(n15848) );
  NANDN U33679 ( .A(y[4064]), .B(x[4064]), .Z(n40276) );
  NANDN U33680 ( .A(y[4065]), .B(x[4065]), .Z(n25460) );
  NAND U33681 ( .A(n40276), .B(n25460), .Z(n56304) );
  OR U33682 ( .A(n15848), .B(n56304), .Z(n15849) );
  NANDN U33683 ( .A(x[4065]), .B(y[4065]), .Z(n25461) );
  NANDN U33684 ( .A(x[4066]), .B(y[4066]), .Z(n25458) );
  AND U33685 ( .A(n25461), .B(n25458), .Z(n51721) );
  AND U33686 ( .A(n15849), .B(n51721), .Z(n15850) );
  NANDN U33687 ( .A(y[4066]), .B(x[4066]), .Z(n25459) );
  NANDN U33688 ( .A(y[4067]), .B(x[4067]), .Z(n40285) );
  NAND U33689 ( .A(n25459), .B(n40285), .Z(n56306) );
  OR U33690 ( .A(n15850), .B(n56306), .Z(n15851) );
  NAND U33691 ( .A(n56307), .B(n15851), .Z(n15852) );
  NANDN U33692 ( .A(n51720), .B(n15852), .Z(n15853) );
  NANDN U33693 ( .A(x[4069]), .B(y[4069]), .Z(n25455) );
  NANDN U33694 ( .A(x[4070]), .B(y[4070]), .Z(n25454) );
  AND U33695 ( .A(n25455), .B(n25454), .Z(n51719) );
  AND U33696 ( .A(n15853), .B(n51719), .Z(n15854) );
  NANDN U33697 ( .A(y[4070]), .B(x[4070]), .Z(n40290) );
  NANDN U33698 ( .A(y[4071]), .B(x[4071]), .Z(n40297) );
  AND U33699 ( .A(n40290), .B(n40297), .Z(n56308) );
  NANDN U33700 ( .A(n15854), .B(n56308), .Z(n15855) );
  NANDN U33701 ( .A(n56309), .B(n15855), .Z(n15856) );
  AND U33702 ( .A(n56310), .B(n15856), .Z(n15857) );
  OR U33703 ( .A(n56311), .B(n15857), .Z(n15858) );
  NAND U33704 ( .A(n56312), .B(n15858), .Z(n15859) );
  NANDN U33705 ( .A(n56313), .B(n15859), .Z(n15860) );
  AND U33706 ( .A(n56314), .B(n15860), .Z(n15861) );
  NANDN U33707 ( .A(x[4077]), .B(y[4077]), .Z(n25447) );
  NANDN U33708 ( .A(x[4078]), .B(y[4078]), .Z(n25444) );
  NAND U33709 ( .A(n25447), .B(n25444), .Z(n56315) );
  OR U33710 ( .A(n15861), .B(n56315), .Z(n15862) );
  NAND U33711 ( .A(n56317), .B(n15862), .Z(n15863) );
  XNOR U33712 ( .A(y[4080]), .B(x[4080]), .Z(n40319) );
  NANDN U33713 ( .A(x[4079]), .B(y[4079]), .Z(n25443) );
  AND U33714 ( .A(n40319), .B(n25443), .Z(n51718) );
  AND U33715 ( .A(n15863), .B(n51718), .Z(n15865) );
  NANDN U33716 ( .A(y[4080]), .B(x[4080]), .Z(n15864) );
  NANDN U33717 ( .A(y[4081]), .B(x[4081]), .Z(n25441) );
  AND U33718 ( .A(n15864), .B(n25441), .Z(n56318) );
  NANDN U33719 ( .A(n15865), .B(n56318), .Z(n15866) );
  NAND U33720 ( .A(n15867), .B(n15866), .Z(n15869) );
  NANDN U33721 ( .A(y[4082]), .B(x[4082]), .Z(n15868) );
  NANDN U33722 ( .A(y[4083]), .B(x[4083]), .Z(n25439) );
  AND U33723 ( .A(n15868), .B(n25439), .Z(n51717) );
  AND U33724 ( .A(n15869), .B(n51717), .Z(n15871) );
  XNOR U33725 ( .A(x[4084]), .B(y[4084]), .Z(n25440) );
  ANDN U33726 ( .B(y[4083]), .A(x[4083]), .Z(n56321) );
  ANDN U33727 ( .B(n25440), .A(n56321), .Z(n15870) );
  NANDN U33728 ( .A(n15871), .B(n15870), .Z(n15873) );
  NANDN U33729 ( .A(y[4084]), .B(x[4084]), .Z(n15872) );
  NANDN U33730 ( .A(y[4085]), .B(x[4085]), .Z(n25438) );
  AND U33731 ( .A(n15872), .B(n25438), .Z(n51715) );
  AND U33732 ( .A(n15873), .B(n51715), .Z(n15874) );
  ANDN U33733 ( .B(y[4085]), .A(x[4085]), .Z(n40331) );
  NANDN U33734 ( .A(x[4086]), .B(y[4086]), .Z(n40338) );
  NANDN U33735 ( .A(n40331), .B(n40338), .Z(n56322) );
  OR U33736 ( .A(n15874), .B(n56322), .Z(n15875) );
  NAND U33737 ( .A(n56323), .B(n15875), .Z(n15876) );
  NANDN U33738 ( .A(n51714), .B(n15876), .Z(n15878) );
  NANDN U33739 ( .A(y[4088]), .B(x[4088]), .Z(n15877) );
  NANDN U33740 ( .A(y[4089]), .B(x[4089]), .Z(n40346) );
  AND U33741 ( .A(n15877), .B(n40346), .Z(n51713) );
  AND U33742 ( .A(n15878), .B(n51713), .Z(n15879) );
  NANDN U33743 ( .A(x[4089]), .B(y[4089]), .Z(n25435) );
  NANDN U33744 ( .A(x[4090]), .B(y[4090]), .Z(n25434) );
  AND U33745 ( .A(n25435), .B(n25434), .Z(n56325) );
  NANDN U33746 ( .A(n15879), .B(n56325), .Z(n15880) );
  NANDN U33747 ( .A(n56326), .B(n15880), .Z(n15881) );
  AND U33748 ( .A(n25433), .B(n15881), .Z(n15882) );
  NANDN U33749 ( .A(x[4091]), .B(y[4091]), .Z(n51711) );
  AND U33750 ( .A(n15882), .B(n51711), .Z(n15884) );
  NANDN U33751 ( .A(y[4092]), .B(x[4092]), .Z(n15883) );
  NANDN U33752 ( .A(y[4093]), .B(x[4093]), .Z(n25430) );
  NAND U33753 ( .A(n15883), .B(n25430), .Z(n56327) );
  OR U33754 ( .A(n15884), .B(n56327), .Z(n15885) );
  AND U33755 ( .A(n56328), .B(n15885), .Z(n15886) );
  NANDN U33756 ( .A(y[4094]), .B(x[4094]), .Z(n25429) );
  NANDN U33757 ( .A(y[4095]), .B(x[4095]), .Z(n40361) );
  AND U33758 ( .A(n25429), .B(n40361), .Z(n51710) );
  NANDN U33759 ( .A(n15886), .B(n51710), .Z(n15887) );
  NANDN U33760 ( .A(n15888), .B(n15887), .Z(n15890) );
  NANDN U33761 ( .A(y[4096]), .B(x[4096]), .Z(n15889) );
  NANDN U33762 ( .A(y[4097]), .B(x[4097]), .Z(n40367) );
  AND U33763 ( .A(n15889), .B(n40367), .Z(n56331) );
  AND U33764 ( .A(n15890), .B(n56331), .Z(n15891) );
  NANDN U33765 ( .A(x[4097]), .B(y[4097]), .Z(n25427) );
  NANDN U33766 ( .A(x[4098]), .B(y[4098]), .Z(n25426) );
  NAND U33767 ( .A(n25427), .B(n25426), .Z(n56332) );
  OR U33768 ( .A(n15891), .B(n56332), .Z(n15892) );
  NAND U33769 ( .A(n56333), .B(n15892), .Z(n15893) );
  NANDN U33770 ( .A(n51709), .B(n15893), .Z(n15894) );
  NANDN U33771 ( .A(y[4100]), .B(x[4100]), .Z(n40372) );
  NANDN U33772 ( .A(y[4101]), .B(x[4101]), .Z(n25424) );
  AND U33773 ( .A(n40372), .B(n25424), .Z(n51708) );
  AND U33774 ( .A(n15894), .B(n51708), .Z(n15895) );
  NANDN U33775 ( .A(x[4101]), .B(y[4101]), .Z(n40375) );
  NANDN U33776 ( .A(x[4102]), .B(y[4102]), .Z(n40382) );
  NAND U33777 ( .A(n40375), .B(n40382), .Z(n56336) );
  OR U33778 ( .A(n15895), .B(n56336), .Z(n15896) );
  NANDN U33779 ( .A(y[4102]), .B(x[4102]), .Z(n25423) );
  NANDN U33780 ( .A(y[4103]), .B(x[4103]), .Z(n25422) );
  AND U33781 ( .A(n25423), .B(n25422), .Z(n56337) );
  AND U33782 ( .A(n15896), .B(n56337), .Z(n15897) );
  NANDN U33783 ( .A(x[4103]), .B(y[4103]), .Z(n40381) );
  NANDN U33784 ( .A(x[4104]), .B(y[4104]), .Z(n40388) );
  NAND U33785 ( .A(n40381), .B(n40388), .Z(n56338) );
  OR U33786 ( .A(n15897), .B(n56338), .Z(n15898) );
  NAND U33787 ( .A(n56339), .B(n15898), .Z(n15899) );
  NANDN U33788 ( .A(n51707), .B(n15899), .Z(n15900) );
  NANDN U33789 ( .A(y[4106]), .B(x[4106]), .Z(n25419) );
  NANDN U33790 ( .A(y[4107]), .B(x[4107]), .Z(n25418) );
  AND U33791 ( .A(n25419), .B(n25418), .Z(n51706) );
  AND U33792 ( .A(n15900), .B(n51706), .Z(n15902) );
  NANDN U33793 ( .A(x[4107]), .B(y[4107]), .Z(n40393) );
  XNOR U33794 ( .A(x[4108]), .B(y[4108]), .Z(n15901) );
  NAND U33795 ( .A(n40393), .B(n15901), .Z(n56340) );
  OR U33796 ( .A(n15902), .B(n56340), .Z(n15903) );
  NAND U33797 ( .A(n56341), .B(n15903), .Z(n15904) );
  NANDN U33798 ( .A(n56342), .B(n15904), .Z(n15905) );
  AND U33799 ( .A(n56343), .B(n15905), .Z(n15906) );
  NANDN U33800 ( .A(x[4111]), .B(y[4111]), .Z(n40405) );
  NANDN U33801 ( .A(x[4112]), .B(y[4112]), .Z(n40412) );
  NAND U33802 ( .A(n40405), .B(n40412), .Z(n56344) );
  OR U33803 ( .A(n15906), .B(n56344), .Z(n15907) );
  AND U33804 ( .A(n56345), .B(n15907), .Z(n15908) );
  OR U33805 ( .A(n56347), .B(n15908), .Z(n15909) );
  NAND U33806 ( .A(n56348), .B(n15909), .Z(n15910) );
  NANDN U33807 ( .A(n56349), .B(n15910), .Z(n15911) );
  AND U33808 ( .A(n56350), .B(n15911), .Z(n15912) );
  NANDN U33809 ( .A(x[4117]), .B(y[4117]), .Z(n40424) );
  NANDN U33810 ( .A(x[4118]), .B(y[4118]), .Z(n40433) );
  AND U33811 ( .A(n40424), .B(n40433), .Z(n56351) );
  NANDN U33812 ( .A(n15912), .B(n56351), .Z(n15913) );
  NANDN U33813 ( .A(n51705), .B(n15913), .Z(n15914) );
  NANDN U33814 ( .A(x[4119]), .B(y[4119]), .Z(n40432) );
  NANDN U33815 ( .A(x[4120]), .B(y[4120]), .Z(n40439) );
  AND U33816 ( .A(n40432), .B(n40439), .Z(n51704) );
  AND U33817 ( .A(n15914), .B(n51704), .Z(n15915) );
  NANDN U33818 ( .A(y[4120]), .B(x[4120]), .Z(n25407) );
  NANDN U33819 ( .A(y[4121]), .B(x[4121]), .Z(n25406) );
  NAND U33820 ( .A(n25407), .B(n25406), .Z(n56352) );
  OR U33821 ( .A(n15915), .B(n56352), .Z(n15916) );
  NAND U33822 ( .A(n56353), .B(n15916), .Z(n15917) );
  NANDN U33823 ( .A(n56354), .B(n15917), .Z(n15918) );
  AND U33824 ( .A(n56355), .B(n15918), .Z(n15919) );
  NANDN U33825 ( .A(y[4124]), .B(x[4124]), .Z(n25403) );
  NANDN U33826 ( .A(y[4125]), .B(x[4125]), .Z(n25402) );
  NAND U33827 ( .A(n25403), .B(n25402), .Z(n56356) );
  OR U33828 ( .A(n15919), .B(n56356), .Z(n15920) );
  AND U33829 ( .A(n56357), .B(n15920), .Z(n15921) );
  NANDN U33830 ( .A(y[4126]), .B(x[4126]), .Z(n25401) );
  NANDN U33831 ( .A(y[4127]), .B(x[4127]), .Z(n40457) );
  AND U33832 ( .A(n25401), .B(n40457), .Z(n51703) );
  NANDN U33833 ( .A(n15921), .B(n51703), .Z(n15922) );
  NANDN U33834 ( .A(n15923), .B(n15922), .Z(n15925) );
  NANDN U33835 ( .A(y[4128]), .B(x[4128]), .Z(n15924) );
  NANDN U33836 ( .A(y[4129]), .B(x[4129]), .Z(n40464) );
  AND U33837 ( .A(n15924), .B(n40464), .Z(n56361) );
  AND U33838 ( .A(n15925), .B(n56361), .Z(n15926) );
  NANDN U33839 ( .A(x[4129]), .B(y[4129]), .Z(n25399) );
  NANDN U33840 ( .A(x[4130]), .B(y[4130]), .Z(n40469) );
  NAND U33841 ( .A(n25399), .B(n40469), .Z(n56362) );
  OR U33842 ( .A(n15926), .B(n56362), .Z(n15927) );
  NAND U33843 ( .A(n56363), .B(n15927), .Z(n15928) );
  NANDN U33844 ( .A(n51702), .B(n15928), .Z(n15929) );
  NANDN U33845 ( .A(y[4132]), .B(x[4132]), .Z(n40471) );
  NANDN U33846 ( .A(y[4133]), .B(x[4133]), .Z(n40477) );
  AND U33847 ( .A(n40471), .B(n40477), .Z(n51701) );
  AND U33848 ( .A(n15929), .B(n51701), .Z(n15931) );
  XNOR U33849 ( .A(x[4134]), .B(y[4134]), .Z(n40478) );
  NANDN U33850 ( .A(x[4133]), .B(y[4133]), .Z(n56364) );
  NAND U33851 ( .A(n40478), .B(n56364), .Z(n15930) );
  OR U33852 ( .A(n15931), .B(n15930), .Z(n15933) );
  NANDN U33853 ( .A(y[4134]), .B(x[4134]), .Z(n15932) );
  NANDN U33854 ( .A(y[4135]), .B(x[4135]), .Z(n25396) );
  AND U33855 ( .A(n15932), .B(n25396), .Z(n56366) );
  AND U33856 ( .A(n15933), .B(n56366), .Z(n15934) );
  ANDN U33857 ( .B(y[4135]), .A(x[4135]), .Z(n25397) );
  NANDN U33858 ( .A(x[4136]), .B(y[4136]), .Z(n25394) );
  NANDN U33859 ( .A(n25397), .B(n25394), .Z(n56367) );
  OR U33860 ( .A(n15934), .B(n56367), .Z(n15935) );
  NAND U33861 ( .A(n56368), .B(n15935), .Z(n15936) );
  NANDN U33862 ( .A(n51700), .B(n15936), .Z(n15937) );
  NANDN U33863 ( .A(y[4138]), .B(x[4138]), .Z(n40488) );
  NANDN U33864 ( .A(y[4139]), .B(x[4139]), .Z(n40495) );
  AND U33865 ( .A(n40488), .B(n40495), .Z(n51699) );
  AND U33866 ( .A(n15937), .B(n51699), .Z(n15938) );
  NANDN U33867 ( .A(x[4139]), .B(y[4139]), .Z(n25391) );
  NANDN U33868 ( .A(x[4140]), .B(y[4140]), .Z(n25390) );
  NAND U33869 ( .A(n25391), .B(n25390), .Z(n56370) );
  OR U33870 ( .A(n15938), .B(n56370), .Z(n15939) );
  NANDN U33871 ( .A(y[4140]), .B(x[4140]), .Z(n40494) );
  NANDN U33872 ( .A(y[4141]), .B(x[4141]), .Z(n40501) );
  AND U33873 ( .A(n40494), .B(n40501), .Z(n56371) );
  AND U33874 ( .A(n15939), .B(n56371), .Z(n15940) );
  NANDN U33875 ( .A(x[4141]), .B(y[4141]), .Z(n25389) );
  NANDN U33876 ( .A(x[4142]), .B(y[4142]), .Z(n40504) );
  NAND U33877 ( .A(n25389), .B(n40504), .Z(n56372) );
  OR U33878 ( .A(n15940), .B(n56372), .Z(n15941) );
  NAND U33879 ( .A(n56373), .B(n15941), .Z(n15942) );
  NANDN U33880 ( .A(n51698), .B(n15942), .Z(n15943) );
  NANDN U33881 ( .A(y[4144]), .B(x[4144]), .Z(n25387) );
  NANDN U33882 ( .A(y[4145]), .B(x[4145]), .Z(n25386) );
  AND U33883 ( .A(n25387), .B(n25386), .Z(n51697) );
  AND U33884 ( .A(n15943), .B(n51697), .Z(n15944) );
  ANDN U33885 ( .B(y[4146]), .A(x[4146]), .Z(n40516) );
  NANDN U33886 ( .A(x[4145]), .B(y[4145]), .Z(n40509) );
  NANDN U33887 ( .A(n40516), .B(n40509), .Z(n56374) );
  OR U33888 ( .A(n15944), .B(n56374), .Z(n15945) );
  NAND U33889 ( .A(n56375), .B(n15945), .Z(n15946) );
  AND U33890 ( .A(n25384), .B(n15946), .Z(n15947) );
  NANDN U33891 ( .A(x[4147]), .B(y[4147]), .Z(n51695) );
  AND U33892 ( .A(n15947), .B(n51695), .Z(n15949) );
  NANDN U33893 ( .A(y[4148]), .B(x[4148]), .Z(n15948) );
  NANDN U33894 ( .A(y[4149]), .B(x[4149]), .Z(n25382) );
  NAND U33895 ( .A(n15948), .B(n25382), .Z(n56378) );
  OR U33896 ( .A(n15949), .B(n56378), .Z(n15950) );
  NAND U33897 ( .A(n56379), .B(n15950), .Z(n15951) );
  NANDN U33898 ( .A(y[4150]), .B(x[4150]), .Z(n25381) );
  NANDN U33899 ( .A(y[4151]), .B(x[4151]), .Z(n25379) );
  AND U33900 ( .A(n25381), .B(n25379), .Z(n51694) );
  AND U33901 ( .A(n15951), .B(n51694), .Z(n15952) );
  NOR U33902 ( .A(n40525), .B(n15952), .Z(n15953) );
  NAND U33903 ( .A(n25380), .B(n15953), .Z(n15954) );
  NANDN U33904 ( .A(n56382), .B(n15954), .Z(n15955) );
  AND U33905 ( .A(n40534), .B(n15955), .Z(n15956) );
  NANDN U33906 ( .A(x[4153]), .B(y[4153]), .Z(n51692) );
  AND U33907 ( .A(n15956), .B(n51692), .Z(n15957) );
  ANDN U33908 ( .B(n56383), .A(n15957), .Z(n15958) );
  XNOR U33909 ( .A(y[4156]), .B(x[4156]), .Z(n40540) );
  NANDN U33910 ( .A(x[4155]), .B(y[4155]), .Z(n25378) );
  NAND U33911 ( .A(n40540), .B(n25378), .Z(n51691) );
  OR U33912 ( .A(n15958), .B(n51691), .Z(n15959) );
  NAND U33913 ( .A(n51690), .B(n15959), .Z(n15960) );
  NANDN U33914 ( .A(n56384), .B(n15960), .Z(n15961) );
  AND U33915 ( .A(n56385), .B(n15961), .Z(n15963) );
  NANDN U33916 ( .A(x[4159]), .B(y[4159]), .Z(n25374) );
  XNOR U33917 ( .A(y[4160]), .B(x[4160]), .Z(n15962) );
  AND U33918 ( .A(n25374), .B(n15962), .Z(n51689) );
  NANDN U33919 ( .A(n15963), .B(n51689), .Z(n15964) );
  NANDN U33920 ( .A(n56388), .B(n15964), .Z(n15965) );
  NANDN U33921 ( .A(x[4161]), .B(y[4161]), .Z(n25372) );
  NANDN U33922 ( .A(x[4162]), .B(y[4162]), .Z(n25371) );
  AND U33923 ( .A(n25372), .B(n25371), .Z(n56389) );
  AND U33924 ( .A(n15965), .B(n56389), .Z(n15966) );
  NANDN U33925 ( .A(y[4162]), .B(x[4162]), .Z(n40557) );
  NANDN U33926 ( .A(y[4163]), .B(x[4163]), .Z(n25369) );
  NAND U33927 ( .A(n40557), .B(n25369), .Z(n51688) );
  OR U33928 ( .A(n15966), .B(n51688), .Z(n15967) );
  NAND U33929 ( .A(n51687), .B(n15967), .Z(n15968) );
  NANDN U33930 ( .A(n51686), .B(n15968), .Z(n15969) );
  AND U33931 ( .A(n56390), .B(n15969), .Z(n15971) );
  NANDN U33932 ( .A(y[4166]), .B(x[4166]), .Z(n15970) );
  NANDN U33933 ( .A(y[4167]), .B(x[4167]), .Z(n40574) );
  NAND U33934 ( .A(n15970), .B(n40574), .Z(n51685) );
  OR U33935 ( .A(n15971), .B(n51685), .Z(n15972) );
  AND U33936 ( .A(n56391), .B(n15972), .Z(n15973) );
  NANDN U33937 ( .A(y[4168]), .B(x[4168]), .Z(n40573) );
  NANDN U33938 ( .A(y[4169]), .B(x[4169]), .Z(n40580) );
  NAND U33939 ( .A(n40573), .B(n40580), .Z(n51684) );
  OR U33940 ( .A(n15973), .B(n51684), .Z(n15974) );
  NAND U33941 ( .A(n56392), .B(n15974), .Z(n15975) );
  AND U33942 ( .A(n56393), .B(n15975), .Z(n15976) );
  OR U33943 ( .A(n56394), .B(n15976), .Z(n15977) );
  NAND U33944 ( .A(n56396), .B(n15977), .Z(n15978) );
  NANDN U33945 ( .A(n56397), .B(n15978), .Z(n15979) );
  AND U33946 ( .A(n56398), .B(n15979), .Z(n15980) );
  ANDN U33947 ( .B(y[4175]), .A(x[4175]), .Z(n40596) );
  NANDN U33948 ( .A(x[4176]), .B(y[4176]), .Z(n25357) );
  NANDN U33949 ( .A(n40596), .B(n25357), .Z(n56399) );
  OR U33950 ( .A(n15980), .B(n56399), .Z(n15981) );
  AND U33951 ( .A(n56400), .B(n15981), .Z(n15982) );
  NANDN U33952 ( .A(x[4177]), .B(y[4177]), .Z(n25356) );
  NANDN U33953 ( .A(x[4178]), .B(y[4178]), .Z(n25355) );
  NAND U33954 ( .A(n25356), .B(n25355), .Z(n56401) );
  OR U33955 ( .A(n15982), .B(n56401), .Z(n15983) );
  NAND U33956 ( .A(n51683), .B(n15983), .Z(n15984) );
  NANDN U33957 ( .A(n56402), .B(n15984), .Z(n15985) );
  NANDN U33958 ( .A(y[4180]), .B(x[4180]), .Z(n40612) );
  NANDN U33959 ( .A(y[4181]), .B(x[4181]), .Z(n25353) );
  AND U33960 ( .A(n40612), .B(n25353), .Z(n56403) );
  AND U33961 ( .A(n15985), .B(n56403), .Z(n15986) );
  NANDN U33962 ( .A(x[4181]), .B(y[4181]), .Z(n40615) );
  NANDN U33963 ( .A(x[4182]), .B(y[4182]), .Z(n40622) );
  AND U33964 ( .A(n40615), .B(n40622), .Z(n56404) );
  NANDN U33965 ( .A(n15986), .B(n56404), .Z(n15987) );
  NANDN U33966 ( .A(n56405), .B(n15987), .Z(n15988) );
  AND U33967 ( .A(n56406), .B(n15988), .Z(n15989) );
  OR U33968 ( .A(n56407), .B(n15989), .Z(n15990) );
  NAND U33969 ( .A(n56408), .B(n15990), .Z(n15991) );
  NANDN U33970 ( .A(n56409), .B(n15991), .Z(n15992) );
  AND U33971 ( .A(n56410), .B(n15992), .Z(n15993) );
  ANDN U33972 ( .B(x[4189]), .A(y[4189]), .Z(n40646) );
  NANDN U33973 ( .A(y[4188]), .B(x[4188]), .Z(n25346) );
  NANDN U33974 ( .A(n40646), .B(n25346), .Z(n56412) );
  OR U33975 ( .A(n15993), .B(n56412), .Z(n15994) );
  AND U33976 ( .A(n56413), .B(n15994), .Z(n15995) );
  ANDN U33977 ( .B(x[4190]), .A(y[4190]), .Z(n40644) );
  NANDN U33978 ( .A(y[4191]), .B(x[4191]), .Z(n25344) );
  NANDN U33979 ( .A(n40644), .B(n25344), .Z(n56414) );
  OR U33980 ( .A(n15995), .B(n56414), .Z(n15996) );
  NAND U33981 ( .A(n51682), .B(n15996), .Z(n15997) );
  NANDN U33982 ( .A(n56415), .B(n15997), .Z(n15998) );
  XNOR U33983 ( .A(y[4194]), .B(x[4194]), .Z(n40658) );
  NANDN U33984 ( .A(x[4193]), .B(y[4193]), .Z(n40654) );
  AND U33985 ( .A(n40658), .B(n40654), .Z(n56416) );
  AND U33986 ( .A(n15998), .B(n56416), .Z(n16000) );
  NANDN U33987 ( .A(y[4194]), .B(x[4194]), .Z(n15999) );
  NANDN U33988 ( .A(y[4195]), .B(x[4195]), .Z(n25343) );
  AND U33989 ( .A(n15999), .B(n25343), .Z(n56417) );
  NANDN U33990 ( .A(n16000), .B(n56417), .Z(n16001) );
  NANDN U33991 ( .A(n56418), .B(n16001), .Z(n16002) );
  AND U33992 ( .A(n56419), .B(n16002), .Z(n16003) );
  OR U33993 ( .A(n56420), .B(n16003), .Z(n16004) );
  NAND U33994 ( .A(n56421), .B(n16004), .Z(n16005) );
  NANDN U33995 ( .A(n56422), .B(n16005), .Z(n16006) );
  NAND U33996 ( .A(n56423), .B(n16006), .Z(n16007) );
  AND U33997 ( .A(n40683), .B(n16007), .Z(n16008) );
  NAND U33998 ( .A(n25337), .B(n16008), .Z(n16009) );
  NANDN U33999 ( .A(n56424), .B(n16009), .Z(n16010) );
  AND U34000 ( .A(n40689), .B(n16010), .Z(n16011) );
  NANDN U34001 ( .A(x[4203]), .B(y[4203]), .Z(n56427) );
  AND U34002 ( .A(n16011), .B(n56427), .Z(n16012) );
  ANDN U34003 ( .B(n56430), .A(n16012), .Z(n16013) );
  OR U34004 ( .A(n56431), .B(n16013), .Z(n16014) );
  NAND U34005 ( .A(n56432), .B(n16014), .Z(n16015) );
  NANDN U34006 ( .A(n56433), .B(n16015), .Z(n16016) );
  AND U34007 ( .A(n56434), .B(n16016), .Z(n16017) );
  NANDN U34008 ( .A(x[4209]), .B(y[4209]), .Z(n25332) );
  NANDN U34009 ( .A(x[4210]), .B(y[4210]), .Z(n25331) );
  NAND U34010 ( .A(n25332), .B(n25331), .Z(n56435) );
  OR U34011 ( .A(n16017), .B(n56435), .Z(n16018) );
  NAND U34012 ( .A(n56436), .B(n16018), .Z(n16019) );
  AND U34013 ( .A(n56437), .B(n16019), .Z(n16020) );
  OR U34014 ( .A(n56438), .B(n16020), .Z(n16021) );
  AND U34015 ( .A(n16022), .B(n16021), .Z(n16023) );
  OR U34016 ( .A(n56439), .B(n16023), .Z(n16024) );
  NAND U34017 ( .A(n56440), .B(n16024), .Z(n16025) );
  NANDN U34018 ( .A(n56441), .B(n16025), .Z(n16026) );
  AND U34019 ( .A(n56442), .B(n16026), .Z(n16027) );
  ANDN U34020 ( .B(x[4219]), .A(y[4219]), .Z(n40736) );
  NANDN U34021 ( .A(y[4218]), .B(x[4218]), .Z(n40728) );
  NANDN U34022 ( .A(n40736), .B(n40728), .Z(n56443) );
  OR U34023 ( .A(n16027), .B(n56443), .Z(n16028) );
  AND U34024 ( .A(n56444), .B(n16028), .Z(n16029) );
  OR U34025 ( .A(n56446), .B(n16029), .Z(n16030) );
  NAND U34026 ( .A(n56448), .B(n16030), .Z(n16031) );
  NANDN U34027 ( .A(n56450), .B(n16031), .Z(n16032) );
  NAND U34028 ( .A(n56452), .B(n16032), .Z(n16033) );
  NAND U34029 ( .A(n56453), .B(n16033), .Z(n16034) );
  NANDN U34030 ( .A(n56456), .B(n16034), .Z(n16035) );
  AND U34031 ( .A(n56458), .B(n16035), .Z(n16036) );
  OR U34032 ( .A(n56460), .B(n16036), .Z(n16037) );
  NAND U34033 ( .A(n56462), .B(n16037), .Z(n16038) );
  NANDN U34034 ( .A(n56464), .B(n16038), .Z(n16039) );
  NAND U34035 ( .A(n56466), .B(n16039), .Z(n16040) );
  AND U34036 ( .A(n25311), .B(n16040), .Z(n16041) );
  NAND U34037 ( .A(n56470), .B(n16041), .Z(n16042) );
  NANDN U34038 ( .A(n56472), .B(n16042), .Z(n16043) );
  AND U34039 ( .A(n56474), .B(n16043), .Z(n16044) );
  OR U34040 ( .A(n56476), .B(n16044), .Z(n16045) );
  AND U34041 ( .A(n16046), .B(n16045), .Z(n16047) );
  OR U34042 ( .A(n56480), .B(n16047), .Z(n16048) );
  NAND U34043 ( .A(n56482), .B(n16048), .Z(n16049) );
  NANDN U34044 ( .A(n56484), .B(n16049), .Z(n16050) );
  AND U34045 ( .A(n56485), .B(n16050), .Z(n16051) );
  NANDN U34046 ( .A(y[4240]), .B(x[4240]), .Z(n25301) );
  NANDN U34047 ( .A(y[4241]), .B(x[4241]), .Z(n40798) );
  NAND U34048 ( .A(n25301), .B(n40798), .Z(n56486) );
  OR U34049 ( .A(n16051), .B(n56486), .Z(n16052) );
  AND U34050 ( .A(n56487), .B(n16052), .Z(n16053) );
  OR U34051 ( .A(n56488), .B(n16053), .Z(n16054) );
  NAND U34052 ( .A(n56489), .B(n16054), .Z(n16055) );
  NANDN U34053 ( .A(n56490), .B(n16055), .Z(n16056) );
  AND U34054 ( .A(n56491), .B(n16056), .Z(n16058) );
  ANDN U34055 ( .B(x[4247]), .A(y[4247]), .Z(n40815) );
  NANDN U34056 ( .A(y[4246]), .B(x[4246]), .Z(n16057) );
  NANDN U34057 ( .A(n40815), .B(n16057), .Z(n56492) );
  OR U34058 ( .A(n16058), .B(n56492), .Z(n16059) );
  AND U34059 ( .A(n16060), .B(n16059), .Z(n16062) );
  NANDN U34060 ( .A(y[4248]), .B(x[4248]), .Z(n16061) );
  NANDN U34061 ( .A(y[4249]), .B(x[4249]), .Z(n25294) );
  NAND U34062 ( .A(n16061), .B(n25294), .Z(n56493) );
  OR U34063 ( .A(n16062), .B(n56493), .Z(n16063) );
  NAND U34064 ( .A(n56494), .B(n16063), .Z(n16064) );
  NANDN U34065 ( .A(n56495), .B(n16064), .Z(n16065) );
  NANDN U34066 ( .A(x[4251]), .B(y[4251]), .Z(n25291) );
  NANDN U34067 ( .A(x[4252]), .B(y[4252]), .Z(n40830) );
  AND U34068 ( .A(n25291), .B(n40830), .Z(n56496) );
  AND U34069 ( .A(n16065), .B(n56496), .Z(n16066) );
  NANDN U34070 ( .A(y[4252]), .B(x[4252]), .Z(n40825) );
  NANDN U34071 ( .A(y[4253]), .B(x[4253]), .Z(n25290) );
  NAND U34072 ( .A(n40825), .B(n25290), .Z(n51673) );
  OR U34073 ( .A(n16066), .B(n51673), .Z(n16067) );
  NAND U34074 ( .A(n51672), .B(n16067), .Z(n16068) );
  NANDN U34075 ( .A(n56499), .B(n16068), .Z(n16069) );
  AND U34076 ( .A(n56500), .B(n16069), .Z(n16070) );
  ANDN U34077 ( .B(x[4257]), .A(y[4257]), .Z(n40845) );
  NANDN U34078 ( .A(y[4256]), .B(x[4256]), .Z(n25287) );
  NANDN U34079 ( .A(n40845), .B(n25287), .Z(n56501) );
  OR U34080 ( .A(n16070), .B(n56501), .Z(n16071) );
  XOR U34081 ( .A(x[4258]), .B(y[4258]), .Z(n40846) );
  ANDN U34082 ( .B(n16071), .A(n40846), .Z(n16072) );
  NANDN U34083 ( .A(x[4257]), .B(y[4257]), .Z(n56502) );
  AND U34084 ( .A(n16072), .B(n56502), .Z(n16074) );
  NANDN U34085 ( .A(y[4258]), .B(x[4258]), .Z(n16073) );
  NANDN U34086 ( .A(y[4259]), .B(x[4259]), .Z(n40852) );
  NAND U34087 ( .A(n16073), .B(n40852), .Z(n56504) );
  OR U34088 ( .A(n16074), .B(n56504), .Z(n16075) );
  NAND U34089 ( .A(n56505), .B(n16075), .Z(n16076) );
  NANDN U34090 ( .A(y[4260]), .B(x[4260]), .Z(n40851) );
  NANDN U34091 ( .A(y[4261]), .B(x[4261]), .Z(n25286) );
  AND U34092 ( .A(n40851), .B(n25286), .Z(n56506) );
  AND U34093 ( .A(n16076), .B(n56506), .Z(n16078) );
  NANDN U34094 ( .A(x[4261]), .B(y[4261]), .Z(n40856) );
  XNOR U34095 ( .A(y[4262]), .B(x[4262]), .Z(n16077) );
  NAND U34096 ( .A(n40856), .B(n16077), .Z(n51671) );
  OR U34097 ( .A(n16078), .B(n51671), .Z(n16079) );
  NANDN U34098 ( .A(y[4262]), .B(x[4262]), .Z(n25285) );
  NANDN U34099 ( .A(y[4263]), .B(x[4263]), .Z(n25281) );
  AND U34100 ( .A(n25285), .B(n25281), .Z(n51670) );
  AND U34101 ( .A(n16079), .B(n51670), .Z(n16080) );
  XNOR U34102 ( .A(y[4264]), .B(x[4264]), .Z(n25282) );
  NANDN U34103 ( .A(x[4263]), .B(y[4263]), .Z(n25283) );
  NAND U34104 ( .A(n25282), .B(n25283), .Z(n56507) );
  OR U34105 ( .A(n16080), .B(n56507), .Z(n16081) );
  NAND U34106 ( .A(n56508), .B(n16081), .Z(n16082) );
  AND U34107 ( .A(n56509), .B(n16082), .Z(n16083) );
  OR U34108 ( .A(n56510), .B(n16083), .Z(n16084) );
  NAND U34109 ( .A(n56512), .B(n16084), .Z(n16085) );
  NANDN U34110 ( .A(n56513), .B(n16085), .Z(n16086) );
  NAND U34111 ( .A(n25274), .B(n16086), .Z(n16087) );
  ANDN U34112 ( .B(y[4269]), .A(x[4269]), .Z(n25275) );
  OR U34113 ( .A(n16087), .B(n25275), .Z(n16088) );
  NAND U34114 ( .A(n56514), .B(n16088), .Z(n16089) );
  NANDN U34115 ( .A(n56515), .B(n16089), .Z(n16090) );
  AND U34116 ( .A(n56516), .B(n16090), .Z(n16091) );
  NOR U34117 ( .A(n25268), .B(n16091), .Z(n16092) );
  XNOR U34118 ( .A(x[4274]), .B(y[4274]), .Z(n40888) );
  AND U34119 ( .A(n16092), .B(n40888), .Z(n16093) );
  OR U34120 ( .A(n56519), .B(n16093), .Z(n16094) );
  NAND U34121 ( .A(n56520), .B(n16094), .Z(n16095) );
  NANDN U34122 ( .A(n56521), .B(n16095), .Z(n16096) );
  AND U34123 ( .A(n56522), .B(n16096), .Z(n16097) );
  NANDN U34124 ( .A(y[4278]), .B(x[4278]), .Z(n40900) );
  ANDN U34125 ( .B(x[4279]), .A(y[4279]), .Z(n40906) );
  ANDN U34126 ( .B(n40900), .A(n40906), .Z(n56523) );
  NANDN U34127 ( .A(n16097), .B(n56523), .Z(n16098) );
  NANDN U34128 ( .A(n56524), .B(n16098), .Z(n16100) );
  NANDN U34129 ( .A(y[4280]), .B(x[4280]), .Z(n16099) );
  NANDN U34130 ( .A(y[4281]), .B(x[4281]), .Z(n25262) );
  AND U34131 ( .A(n16099), .B(n25262), .Z(n56525) );
  AND U34132 ( .A(n16100), .B(n56525), .Z(n16102) );
  NANDN U34133 ( .A(x[4281]), .B(y[4281]), .Z(n40910) );
  XNOR U34134 ( .A(x[4282]), .B(y[4282]), .Z(n16101) );
  NAND U34135 ( .A(n40910), .B(n16101), .Z(n56526) );
  OR U34136 ( .A(n16102), .B(n56526), .Z(n16103) );
  NAND U34137 ( .A(n56529), .B(n16103), .Z(n16104) );
  NANDN U34138 ( .A(n51667), .B(n16104), .Z(n16105) );
  NANDN U34139 ( .A(y[4284]), .B(x[4284]), .Z(n25257) );
  NANDN U34140 ( .A(y[4285]), .B(x[4285]), .Z(n25256) );
  AND U34141 ( .A(n25257), .B(n25256), .Z(n51666) );
  AND U34142 ( .A(n16105), .B(n51666), .Z(n16106) );
  ANDN U34143 ( .B(y[4286]), .A(x[4286]), .Z(n40928) );
  NANDN U34144 ( .A(x[4285]), .B(y[4285]), .Z(n40920) );
  NANDN U34145 ( .A(n40928), .B(n40920), .Z(n51665) );
  OR U34146 ( .A(n16106), .B(n51665), .Z(n16107) );
  AND U34147 ( .A(n56530), .B(n16107), .Z(n16108) );
  OR U34148 ( .A(n56531), .B(n16108), .Z(n16109) );
  NAND U34149 ( .A(n56532), .B(n16109), .Z(n16110) );
  NANDN U34150 ( .A(n56533), .B(n16110), .Z(n16111) );
  AND U34151 ( .A(n56534), .B(n16111), .Z(n16112) );
  NANDN U34152 ( .A(x[4291]), .B(y[4291]), .Z(n40937) );
  NANDN U34153 ( .A(x[4292]), .B(y[4292]), .Z(n25250) );
  AND U34154 ( .A(n40937), .B(n25250), .Z(n51664) );
  NANDN U34155 ( .A(n16112), .B(n51664), .Z(n16113) );
  NANDN U34156 ( .A(n56535), .B(n16113), .Z(n16114) );
  XNOR U34157 ( .A(y[4294]), .B(x[4294]), .Z(n40948) );
  NANDN U34158 ( .A(x[4293]), .B(y[4293]), .Z(n25249) );
  AND U34159 ( .A(n40948), .B(n25249), .Z(n56536) );
  AND U34160 ( .A(n16114), .B(n56536), .Z(n16116) );
  NANDN U34161 ( .A(y[4294]), .B(x[4294]), .Z(n16115) );
  NANDN U34162 ( .A(y[4295]), .B(x[4295]), .Z(n25246) );
  NAND U34163 ( .A(n16115), .B(n25246), .Z(n56537) );
  OR U34164 ( .A(n16116), .B(n56537), .Z(n16117) );
  NAND U34165 ( .A(n56540), .B(n16117), .Z(n16118) );
  NANDN U34166 ( .A(n51663), .B(n16118), .Z(n16119) );
  AND U34167 ( .A(n56541), .B(n16119), .Z(n16121) );
  ANDN U34168 ( .B(x[4299]), .A(y[4299]), .Z(n40965) );
  NANDN U34169 ( .A(y[4298]), .B(x[4298]), .Z(n16120) );
  NANDN U34170 ( .A(n40965), .B(n16120), .Z(n56542) );
  OR U34171 ( .A(n16121), .B(n56542), .Z(n16122) );
  NAND U34172 ( .A(n56543), .B(n16122), .Z(n16123) );
  AND U34173 ( .A(n56544), .B(n16123), .Z(n16124) );
  ANDN U34174 ( .B(n56545), .A(n16124), .Z(n16125) );
  NAND U34175 ( .A(n25239), .B(n16125), .Z(n16126) );
  NANDN U34176 ( .A(n56547), .B(n16126), .Z(n16127) );
  AND U34177 ( .A(n40975), .B(n16127), .Z(n16128) );
  NANDN U34178 ( .A(x[4303]), .B(y[4303]), .Z(n51661) );
  NAND U34179 ( .A(n16128), .B(n51661), .Z(n16129) );
  NANDN U34180 ( .A(n56548), .B(n16129), .Z(n16130) );
  AND U34181 ( .A(n56549), .B(n16130), .Z(n16131) );
  OR U34182 ( .A(n56550), .B(n16131), .Z(n16132) );
  NAND U34183 ( .A(n56551), .B(n16132), .Z(n16133) );
  NANDN U34184 ( .A(n51660), .B(n16133), .Z(n16134) );
  NANDN U34185 ( .A(x[4309]), .B(y[4309]), .Z(n40988) );
  NANDN U34186 ( .A(x[4310]), .B(y[4310]), .Z(n40995) );
  AND U34187 ( .A(n40988), .B(n40995), .Z(n51659) );
  AND U34188 ( .A(n16134), .B(n51659), .Z(n16135) );
  NANDN U34189 ( .A(y[4310]), .B(x[4310]), .Z(n25232) );
  NANDN U34190 ( .A(y[4311]), .B(x[4311]), .Z(n25231) );
  NAND U34191 ( .A(n25232), .B(n25231), .Z(n56553) );
  OR U34192 ( .A(n16135), .B(n56553), .Z(n16136) );
  AND U34193 ( .A(n56554), .B(n16136), .Z(n16137) );
  OR U34194 ( .A(n56555), .B(n16137), .Z(n16138) );
  NAND U34195 ( .A(n56556), .B(n16138), .Z(n16139) );
  NANDN U34196 ( .A(n56557), .B(n16139), .Z(n16140) );
  AND U34197 ( .A(n56558), .B(n16140), .Z(n16141) );
  OR U34198 ( .A(n56559), .B(n16141), .Z(n16142) );
  NAND U34199 ( .A(n56560), .B(n16142), .Z(n16143) );
  NANDN U34200 ( .A(n56561), .B(n16143), .Z(n16144) );
  AND U34201 ( .A(n56562), .B(n16144), .Z(n16145) );
  OR U34202 ( .A(n56563), .B(n16145), .Z(n16146) );
  AND U34203 ( .A(n16147), .B(n16146), .Z(n16148) );
  OR U34204 ( .A(n56566), .B(n16148), .Z(n16149) );
  NAND U34205 ( .A(n56567), .B(n16149), .Z(n16150) );
  NANDN U34206 ( .A(n56568), .B(n16150), .Z(n16151) );
  AND U34207 ( .A(n56569), .B(n16151), .Z(n16153) );
  NANDN U34208 ( .A(y[4326]), .B(x[4326]), .Z(n16152) );
  NANDN U34209 ( .A(y[4327]), .B(x[4327]), .Z(n25223) );
  NAND U34210 ( .A(n16152), .B(n25223), .Z(n56571) );
  OR U34211 ( .A(n16153), .B(n56571), .Z(n16154) );
  AND U34212 ( .A(n56572), .B(n16154), .Z(n16155) );
  OR U34213 ( .A(n56573), .B(n16155), .Z(n16156) );
  NAND U34214 ( .A(n56574), .B(n16156), .Z(n16157) );
  NANDN U34215 ( .A(n56575), .B(n16157), .Z(n16158) );
  AND U34216 ( .A(n56576), .B(n16158), .Z(n16159) );
  OR U34217 ( .A(n56577), .B(n16159), .Z(n16160) );
  NAND U34218 ( .A(n56578), .B(n16160), .Z(n16161) );
  NANDN U34219 ( .A(n51658), .B(n16161), .Z(n16162) );
  AND U34220 ( .A(n41074), .B(n16162), .Z(n16163) );
  NAND U34221 ( .A(n51657), .B(n16163), .Z(n16164) );
  NANDN U34222 ( .A(n56580), .B(n16164), .Z(n16165) );
  NANDN U34223 ( .A(x[4337]), .B(y[4337]), .Z(n25213) );
  NANDN U34224 ( .A(x[4338]), .B(y[4338]), .Z(n25212) );
  AND U34225 ( .A(n25213), .B(n25212), .Z(n56581) );
  AND U34226 ( .A(n16165), .B(n56581), .Z(n16166) );
  NANDN U34227 ( .A(y[4338]), .B(x[4338]), .Z(n41079) );
  NANDN U34228 ( .A(y[4339]), .B(x[4339]), .Z(n41086) );
  NAND U34229 ( .A(n41079), .B(n41086), .Z(n51656) );
  OR U34230 ( .A(n16166), .B(n51656), .Z(n16167) );
  NAND U34231 ( .A(n51655), .B(n16167), .Z(n16168) );
  NANDN U34232 ( .A(n56584), .B(n16168), .Z(n16169) );
  NANDN U34233 ( .A(x[4341]), .B(y[4341]), .Z(n25209) );
  NANDN U34234 ( .A(x[4342]), .B(y[4342]), .Z(n25208) );
  AND U34235 ( .A(n25209), .B(n25208), .Z(n56586) );
  AND U34236 ( .A(n16169), .B(n56586), .Z(n16170) );
  NANDN U34237 ( .A(y[4342]), .B(x[4342]), .Z(n41091) );
  NANDN U34238 ( .A(y[4343]), .B(x[4343]), .Z(n41098) );
  NAND U34239 ( .A(n41091), .B(n41098), .Z(n56587) );
  OR U34240 ( .A(n16170), .B(n56587), .Z(n16171) );
  NANDN U34241 ( .A(x[4343]), .B(y[4343]), .Z(n25207) );
  NANDN U34242 ( .A(x[4344]), .B(y[4344]), .Z(n25206) );
  AND U34243 ( .A(n25207), .B(n25206), .Z(n56588) );
  AND U34244 ( .A(n16171), .B(n56588), .Z(n16172) );
  NANDN U34245 ( .A(y[4344]), .B(x[4344]), .Z(n41097) );
  NANDN U34246 ( .A(y[4345]), .B(x[4345]), .Z(n41104) );
  NAND U34247 ( .A(n41097), .B(n41104), .Z(n51654) );
  OR U34248 ( .A(n16172), .B(n51654), .Z(n16173) );
  NAND U34249 ( .A(n51653), .B(n16173), .Z(n16174) );
  NANDN U34250 ( .A(n56589), .B(n16174), .Z(n16175) );
  NANDN U34251 ( .A(x[4347]), .B(y[4347]), .Z(n25203) );
  NANDN U34252 ( .A(x[4348]), .B(y[4348]), .Z(n25202) );
  AND U34253 ( .A(n25203), .B(n25202), .Z(n56590) );
  AND U34254 ( .A(n16175), .B(n56590), .Z(n16176) );
  NANDN U34255 ( .A(y[4348]), .B(x[4348]), .Z(n41109) );
  NANDN U34256 ( .A(y[4349]), .B(x[4349]), .Z(n25200) );
  NAND U34257 ( .A(n41109), .B(n25200), .Z(n51652) );
  OR U34258 ( .A(n16176), .B(n51652), .Z(n16177) );
  NAND U34259 ( .A(n51651), .B(n16177), .Z(n16178) );
  NANDN U34260 ( .A(n56591), .B(n16178), .Z(n16181) );
  NANDN U34261 ( .A(x[4352]), .B(y[4352]), .Z(n16180) );
  NANDN U34262 ( .A(x[4351]), .B(y[4351]), .Z(n16179) );
  AND U34263 ( .A(n16180), .B(n16179), .Z(n56594) );
  AND U34264 ( .A(n16181), .B(n56594), .Z(n16184) );
  NANDN U34265 ( .A(y[4352]), .B(x[4352]), .Z(n16183) );
  NANDN U34266 ( .A(y[4353]), .B(x[4353]), .Z(n16182) );
  NAND U34267 ( .A(n16183), .B(n16182), .Z(n56596) );
  OR U34268 ( .A(n16184), .B(n56596), .Z(n16185) );
  NANDN U34269 ( .A(x[4353]), .B(y[4353]), .Z(n41124) );
  NANDN U34270 ( .A(x[4354]), .B(y[4354]), .Z(n25198) );
  AND U34271 ( .A(n41124), .B(n25198), .Z(n56597) );
  AND U34272 ( .A(n16185), .B(n56597), .Z(n16186) );
  ANDN U34273 ( .B(x[4354]), .A(y[4354]), .Z(n41126) );
  NANDN U34274 ( .A(y[4355]), .B(x[4355]), .Z(n41130) );
  NANDN U34275 ( .A(n41126), .B(n41130), .Z(n51650) );
  OR U34276 ( .A(n16186), .B(n51650), .Z(n16187) );
  NAND U34277 ( .A(n51649), .B(n16187), .Z(n16188) );
  NANDN U34278 ( .A(n56598), .B(n16188), .Z(n16189) );
  XNOR U34279 ( .A(y[4358]), .B(x[4358]), .Z(n25196) );
  NANDN U34280 ( .A(x[4357]), .B(y[4357]), .Z(n41134) );
  AND U34281 ( .A(n25196), .B(n41134), .Z(n56599) );
  AND U34282 ( .A(n16189), .B(n56599), .Z(n16191) );
  NANDN U34283 ( .A(y[4358]), .B(x[4358]), .Z(n16190) );
  NANDN U34284 ( .A(y[4359]), .B(x[4359]), .Z(n25193) );
  NAND U34285 ( .A(n16190), .B(n25193), .Z(n51648) );
  OR U34286 ( .A(n16191), .B(n51648), .Z(n16192) );
  AND U34287 ( .A(n16193), .B(n16192), .Z(n16194) );
  OR U34288 ( .A(n56602), .B(n16194), .Z(n16195) );
  NAND U34289 ( .A(n56604), .B(n16195), .Z(n16196) );
  NANDN U34290 ( .A(n56605), .B(n16196), .Z(n16197) );
  AND U34291 ( .A(n25190), .B(n16197), .Z(n16198) );
  NANDN U34292 ( .A(x[4363]), .B(y[4363]), .Z(n56606) );
  AND U34293 ( .A(n16198), .B(n56606), .Z(n16200) );
  NANDN U34294 ( .A(y[4364]), .B(x[4364]), .Z(n16199) );
  NANDN U34295 ( .A(y[4365]), .B(x[4365]), .Z(n25186) );
  AND U34296 ( .A(n16199), .B(n25186), .Z(n51647) );
  NANDN U34297 ( .A(n16200), .B(n51647), .Z(n16201) );
  NAND U34298 ( .A(n16202), .B(n16201), .Z(n16203) );
  AND U34299 ( .A(n56610), .B(n16203), .Z(n16205) );
  NANDN U34300 ( .A(x[4367]), .B(y[4367]), .Z(n41160) );
  XNOR U34301 ( .A(x[4368]), .B(y[4368]), .Z(n16204) );
  NAND U34302 ( .A(n41160), .B(n16204), .Z(n56611) );
  OR U34303 ( .A(n16205), .B(n56611), .Z(n16206) );
  AND U34304 ( .A(n56612), .B(n16206), .Z(n16207) );
  NANDN U34305 ( .A(x[4369]), .B(y[4369]), .Z(n25184) );
  NANDN U34306 ( .A(x[4370]), .B(y[4370]), .Z(n25183) );
  NAND U34307 ( .A(n25184), .B(n25183), .Z(n51645) );
  OR U34308 ( .A(n16207), .B(n51645), .Z(n16208) );
  NAND U34309 ( .A(n56613), .B(n16208), .Z(n16209) );
  NANDN U34310 ( .A(n56614), .B(n16209), .Z(n16210) );
  AND U34311 ( .A(n56615), .B(n16210), .Z(n16212) );
  XNOR U34312 ( .A(x[4374]), .B(y[4374]), .Z(n41179) );
  NANDN U34313 ( .A(x[4373]), .B(y[4373]), .Z(n51643) );
  NAND U34314 ( .A(n41179), .B(n51643), .Z(n16211) );
  OR U34315 ( .A(n16212), .B(n16211), .Z(n16214) );
  NANDN U34316 ( .A(y[4374]), .B(x[4374]), .Z(n16213) );
  NANDN U34317 ( .A(y[4375]), .B(x[4375]), .Z(n25178) );
  AND U34318 ( .A(n16213), .B(n25178), .Z(n56618) );
  AND U34319 ( .A(n16214), .B(n56618), .Z(n16215) );
  NANDN U34320 ( .A(x[4375]), .B(y[4375]), .Z(n41181) );
  NANDN U34321 ( .A(x[4376]), .B(y[4376]), .Z(n25176) );
  NAND U34322 ( .A(n41181), .B(n25176), .Z(n51642) );
  OR U34323 ( .A(n16215), .B(n51642), .Z(n16216) );
  NAND U34324 ( .A(n51641), .B(n16216), .Z(n16217) );
  NANDN U34325 ( .A(n56620), .B(n16217), .Z(n16218) );
  NANDN U34326 ( .A(y[4378]), .B(x[4378]), .Z(n25173) );
  NANDN U34327 ( .A(y[4379]), .B(x[4379]), .Z(n25172) );
  AND U34328 ( .A(n25173), .B(n25172), .Z(n56621) );
  AND U34329 ( .A(n16218), .B(n56621), .Z(n16219) );
  ANDN U34330 ( .B(y[4380]), .A(x[4380]), .Z(n41199) );
  NANDN U34331 ( .A(x[4379]), .B(y[4379]), .Z(n41191) );
  NANDN U34332 ( .A(n41199), .B(n41191), .Z(n56622) );
  OR U34333 ( .A(n16219), .B(n56622), .Z(n16220) );
  NANDN U34334 ( .A(y[4380]), .B(x[4380]), .Z(n25171) );
  NANDN U34335 ( .A(y[4381]), .B(x[4381]), .Z(n41201) );
  AND U34336 ( .A(n25171), .B(n41201), .Z(n56623) );
  AND U34337 ( .A(n16220), .B(n56623), .Z(n16221) );
  XNOR U34338 ( .A(y[4382]), .B(x[4382]), .Z(n41203) );
  NANDN U34339 ( .A(x[4381]), .B(y[4381]), .Z(n41197) );
  NAND U34340 ( .A(n41203), .B(n41197), .Z(n51640) );
  OR U34341 ( .A(n16221), .B(n51640), .Z(n16222) );
  NAND U34342 ( .A(n51639), .B(n16222), .Z(n16223) );
  NANDN U34343 ( .A(n56624), .B(n16223), .Z(n16224) );
  AND U34344 ( .A(n56625), .B(n16224), .Z(n16225) );
  XNOR U34345 ( .A(y[4386]), .B(x[4386]), .Z(n41215) );
  ANDN U34346 ( .B(y[4385]), .A(x[4385]), .Z(n41213) );
  ANDN U34347 ( .B(n41215), .A(n41213), .Z(n56627) );
  NANDN U34348 ( .A(n16225), .B(n56627), .Z(n16226) );
  NANDN U34349 ( .A(n56628), .B(n16226), .Z(n16227) );
  XNOR U34350 ( .A(y[4388]), .B(x[4388]), .Z(n41221) );
  NANDN U34351 ( .A(x[4387]), .B(y[4387]), .Z(n25167) );
  AND U34352 ( .A(n41221), .B(n25167), .Z(n56629) );
  AND U34353 ( .A(n16227), .B(n56629), .Z(n16229) );
  NANDN U34354 ( .A(y[4388]), .B(x[4388]), .Z(n16228) );
  NANDN U34355 ( .A(y[4389]), .B(x[4389]), .Z(n41227) );
  NAND U34356 ( .A(n16228), .B(n41227), .Z(n51638) );
  OR U34357 ( .A(n16229), .B(n51638), .Z(n16230) );
  NAND U34358 ( .A(n51637), .B(n16230), .Z(n16231) );
  NANDN U34359 ( .A(n56630), .B(n16231), .Z(n16232) );
  AND U34360 ( .A(n56631), .B(n16232), .Z(n16233) );
  NANDN U34361 ( .A(y[4392]), .B(x[4392]), .Z(n25163) );
  NANDN U34362 ( .A(y[4393]), .B(x[4393]), .Z(n25161) );
  NAND U34363 ( .A(n25163), .B(n25161), .Z(n56632) );
  OR U34364 ( .A(n16233), .B(n56632), .Z(n16234) );
  AND U34365 ( .A(n16235), .B(n16234), .Z(n16237) );
  NANDN U34366 ( .A(y[4394]), .B(x[4394]), .Z(n16236) );
  NANDN U34367 ( .A(y[4395]), .B(x[4395]), .Z(n25159) );
  NAND U34368 ( .A(n16236), .B(n25159), .Z(n56635) );
  OR U34369 ( .A(n16237), .B(n56635), .Z(n16238) );
  NAND U34370 ( .A(n56636), .B(n16238), .Z(n16239) );
  NANDN U34371 ( .A(n56637), .B(n16239), .Z(n16240) );
  AND U34372 ( .A(n56639), .B(n16240), .Z(n16242) );
  NANDN U34373 ( .A(y[4398]), .B(x[4398]), .Z(n16241) );
  NANDN U34374 ( .A(y[4399]), .B(x[4399]), .Z(n41257) );
  NAND U34375 ( .A(n16241), .B(n41257), .Z(n56640) );
  OR U34376 ( .A(n16242), .B(n56640), .Z(n16243) );
  AND U34377 ( .A(n56641), .B(n16243), .Z(n16244) );
  OR U34378 ( .A(n56642), .B(n16244), .Z(n16245) );
  NAND U34379 ( .A(n56643), .B(n16245), .Z(n16246) );
  NANDN U34380 ( .A(n56644), .B(n16246), .Z(n16247) );
  NAND U34381 ( .A(n56645), .B(n16247), .Z(n16248) );
  NAND U34382 ( .A(n51636), .B(n16248), .Z(n16249) );
  NAND U34383 ( .A(n25148), .B(n16249), .Z(n16250) );
  ANDN U34384 ( .B(y[4405]), .A(x[4405]), .Z(n25149) );
  OR U34385 ( .A(n16250), .B(n25149), .Z(n16252) );
  NANDN U34386 ( .A(y[4406]), .B(x[4406]), .Z(n16251) );
  NANDN U34387 ( .A(y[4407]), .B(x[4407]), .Z(n41278) );
  AND U34388 ( .A(n16251), .B(n41278), .Z(n56648) );
  AND U34389 ( .A(n16252), .B(n56648), .Z(n16253) );
  OR U34390 ( .A(n16254), .B(n16253), .Z(n16255) );
  NAND U34391 ( .A(n56649), .B(n16255), .Z(n16256) );
  NANDN U34392 ( .A(n51633), .B(n16256), .Z(n16257) );
  NANDN U34393 ( .A(y[4410]), .B(x[4410]), .Z(n41283) );
  NANDN U34394 ( .A(y[4411]), .B(x[4411]), .Z(n41290) );
  AND U34395 ( .A(n41283), .B(n41290), .Z(n51632) );
  AND U34396 ( .A(n16257), .B(n51632), .Z(n16258) );
  XNOR U34397 ( .A(x[4414]), .B(y[4414]), .Z(n41295) );
  NANDN U34398 ( .A(x[4413]), .B(y[4413]), .Z(n56655) );
  NANDN U34399 ( .A(y[4414]), .B(x[4414]), .Z(n16259) );
  NANDN U34400 ( .A(y[4415]), .B(x[4415]), .Z(n25143) );
  AND U34401 ( .A(n16259), .B(n25143), .Z(n56657) );
  NANDN U34402 ( .A(x[4415]), .B(y[4415]), .Z(n41298) );
  NANDN U34403 ( .A(x[4416]), .B(y[4416]), .Z(n25141) );
  NAND U34404 ( .A(n41298), .B(n25141), .Z(n51631) );
  NANDN U34405 ( .A(y[4418]), .B(x[4418]), .Z(n25138) );
  NANDN U34406 ( .A(y[4419]), .B(x[4419]), .Z(n25137) );
  AND U34407 ( .A(n25138), .B(n25137), .Z(n56659) );
  NANDN U34408 ( .A(x[4419]), .B(y[4419]), .Z(n41308) );
  NANDN U34409 ( .A(x[4420]), .B(y[4420]), .Z(n41315) );
  NAND U34410 ( .A(n41308), .B(n41315), .Z(n56660) );
  NANDN U34411 ( .A(y[4420]), .B(x[4420]), .Z(n25136) );
  NANDN U34412 ( .A(y[4421]), .B(x[4421]), .Z(n25134) );
  AND U34413 ( .A(n25136), .B(n25134), .Z(n56661) );
  XNOR U34414 ( .A(y[4422]), .B(x[4422]), .Z(n25135) );
  NANDN U34415 ( .A(x[4421]), .B(y[4421]), .Z(n41314) );
  NAND U34416 ( .A(n25135), .B(n41314), .Z(n51629) );
  NANDN U34417 ( .A(y[4424]), .B(x[4424]), .Z(n16260) );
  NANDN U34418 ( .A(y[4425]), .B(x[4425]), .Z(n25128) );
  AND U34419 ( .A(n16260), .B(n25128), .Z(n56664) );
  XNOR U34420 ( .A(y[4426]), .B(x[4426]), .Z(n25129) );
  NANDN U34421 ( .A(x[4425]), .B(y[4425]), .Z(n25130) );
  NAND U34422 ( .A(n25129), .B(n25130), .Z(n51627) );
  NAND U34423 ( .A(n25125), .B(n16261), .Z(n16262) );
  ANDN U34424 ( .B(y[4427]), .A(x[4427]), .Z(n25126) );
  OR U34425 ( .A(n16262), .B(n25126), .Z(n16263) );
  NAND U34426 ( .A(n56667), .B(n16263), .Z(n16265) );
  ANDN U34427 ( .B(y[4429]), .A(x[4429]), .Z(n56668) );
  XNOR U34428 ( .A(x[4430]), .B(y[4430]), .Z(n41336) );
  NANDN U34429 ( .A(n56668), .B(n41336), .Z(n16264) );
  ANDN U34430 ( .B(n16265), .A(n16264), .Z(n16266) );
  OR U34431 ( .A(n56670), .B(n16266), .Z(n16267) );
  NAND U34432 ( .A(n56672), .B(n16267), .Z(n16268) );
  NANDN U34433 ( .A(n56673), .B(n16268), .Z(n16269) );
  AND U34434 ( .A(n56674), .B(n16269), .Z(n16271) );
  ANDN U34435 ( .B(x[4435]), .A(y[4435]), .Z(n41356) );
  NANDN U34436 ( .A(y[4434]), .B(x[4434]), .Z(n16270) );
  NANDN U34437 ( .A(n41356), .B(n16270), .Z(n56675) );
  OR U34438 ( .A(n16271), .B(n56675), .Z(n16272) );
  AND U34439 ( .A(n56676), .B(n16272), .Z(n16274) );
  ANDN U34440 ( .B(x[4437]), .A(y[4437]), .Z(n41364) );
  NANDN U34441 ( .A(y[4436]), .B(x[4436]), .Z(n16273) );
  NANDN U34442 ( .A(n41364), .B(n16273), .Z(n56677) );
  OR U34443 ( .A(n16274), .B(n56677), .Z(n16275) );
  NAND U34444 ( .A(n51625), .B(n16275), .Z(n16276) );
  NANDN U34445 ( .A(n56678), .B(n16276), .Z(n16277) );
  XNOR U34446 ( .A(y[4440]), .B(x[4440]), .Z(n41373) );
  NANDN U34447 ( .A(x[4439]), .B(y[4439]), .Z(n41367) );
  AND U34448 ( .A(n41373), .B(n41367), .Z(n56679) );
  AND U34449 ( .A(n16277), .B(n56679), .Z(n16279) );
  NANDN U34450 ( .A(y[4440]), .B(x[4440]), .Z(n16278) );
  NANDN U34451 ( .A(y[4441]), .B(x[4441]), .Z(n41379) );
  AND U34452 ( .A(n16278), .B(n41379), .Z(n56680) );
  NANDN U34453 ( .A(n16279), .B(n56680), .Z(n16280) );
  NANDN U34454 ( .A(n56681), .B(n16280), .Z(n16281) );
  AND U34455 ( .A(n56682), .B(n16281), .Z(n16282) );
  OR U34456 ( .A(n56683), .B(n16282), .Z(n16283) );
  NAND U34457 ( .A(n56684), .B(n16283), .Z(n16284) );
  NANDN U34458 ( .A(n56685), .B(n16284), .Z(n16285) );
  AND U34459 ( .A(n56686), .B(n16285), .Z(n16286) );
  XNOR U34460 ( .A(y[4448]), .B(x[4448]), .Z(n41403) );
  NANDN U34461 ( .A(x[4447]), .B(y[4447]), .Z(n41397) );
  AND U34462 ( .A(n41403), .B(n41397), .Z(n51624) );
  NANDN U34463 ( .A(n16286), .B(n51624), .Z(n16287) );
  NANDN U34464 ( .A(n51623), .B(n16287), .Z(n16288) );
  AND U34465 ( .A(n25117), .B(n16288), .Z(n16289) );
  NANDN U34466 ( .A(x[4449]), .B(y[4449]), .Z(n56688) );
  AND U34467 ( .A(n16289), .B(n56688), .Z(n16291) );
  NANDN U34468 ( .A(y[4450]), .B(x[4450]), .Z(n16290) );
  NANDN U34469 ( .A(y[4451]), .B(x[4451]), .Z(n41413) );
  NAND U34470 ( .A(n16290), .B(n41413), .Z(n51622) );
  OR U34471 ( .A(n16291), .B(n51622), .Z(n16292) );
  XNOR U34472 ( .A(y[4452]), .B(x[4452]), .Z(n41414) );
  NANDN U34473 ( .A(x[4451]), .B(y[4451]), .Z(n41410) );
  AND U34474 ( .A(n41414), .B(n41410), .Z(n56690) );
  AND U34475 ( .A(n16292), .B(n56690), .Z(n16294) );
  NANDN U34476 ( .A(y[4452]), .B(x[4452]), .Z(n16293) );
  NANDN U34477 ( .A(y[4453]), .B(x[4453]), .Z(n25116) );
  NAND U34478 ( .A(n16293), .B(n25116), .Z(n51621) );
  OR U34479 ( .A(n16294), .B(n51621), .Z(n16295) );
  NAND U34480 ( .A(n51620), .B(n16295), .Z(n16296) );
  NANDN U34481 ( .A(n56691), .B(n16296), .Z(n16297) );
  XNOR U34482 ( .A(y[4456]), .B(x[4456]), .Z(n41426) );
  NANDN U34483 ( .A(x[4455]), .B(y[4455]), .Z(n25113) );
  AND U34484 ( .A(n41426), .B(n25113), .Z(n56692) );
  AND U34485 ( .A(n16297), .B(n56692), .Z(n16299) );
  NANDN U34486 ( .A(y[4456]), .B(x[4456]), .Z(n16298) );
  NANDN U34487 ( .A(y[4457]), .B(x[4457]), .Z(n25111) );
  AND U34488 ( .A(n16298), .B(n25111), .Z(n56693) );
  NANDN U34489 ( .A(n16299), .B(n56693), .Z(n16300) );
  NAND U34490 ( .A(n56694), .B(n16300), .Z(n16301) );
  NANDN U34491 ( .A(n56695), .B(n16301), .Z(n16302) );
  AND U34492 ( .A(n25109), .B(n16302), .Z(n16303) );
  NANDN U34493 ( .A(x[4459]), .B(y[4459]), .Z(n51617) );
  AND U34494 ( .A(n16303), .B(n51617), .Z(n16305) );
  NANDN U34495 ( .A(y[4460]), .B(x[4460]), .Z(n16304) );
  NANDN U34496 ( .A(y[4461]), .B(x[4461]), .Z(n41441) );
  NAND U34497 ( .A(n16304), .B(n41441), .Z(n56698) );
  OR U34498 ( .A(n16305), .B(n56698), .Z(n16306) );
  AND U34499 ( .A(n41442), .B(n16306), .Z(n16307) );
  NANDN U34500 ( .A(x[4461]), .B(y[4461]), .Z(n56699) );
  AND U34501 ( .A(n16307), .B(n56699), .Z(n16309) );
  NANDN U34502 ( .A(y[4462]), .B(x[4462]), .Z(n16308) );
  NANDN U34503 ( .A(y[4463]), .B(x[4463]), .Z(n25106) );
  NAND U34504 ( .A(n16308), .B(n25106), .Z(n56701) );
  OR U34505 ( .A(n16309), .B(n56701), .Z(n16310) );
  AND U34506 ( .A(n56702), .B(n16310), .Z(n16312) );
  NANDN U34507 ( .A(y[4464]), .B(x[4464]), .Z(n16311) );
  NANDN U34508 ( .A(y[4465]), .B(x[4465]), .Z(n25104) );
  NAND U34509 ( .A(n16311), .B(n25104), .Z(n51616) );
  OR U34510 ( .A(n16312), .B(n51616), .Z(n16313) );
  NAND U34511 ( .A(n56703), .B(n16313), .Z(n16314) );
  NANDN U34512 ( .A(n56704), .B(n16314), .Z(n16315) );
  XNOR U34513 ( .A(y[4468]), .B(x[4468]), .Z(n41459) );
  NANDN U34514 ( .A(x[4467]), .B(y[4467]), .Z(n25102) );
  AND U34515 ( .A(n41459), .B(n25102), .Z(n56705) );
  AND U34516 ( .A(n16315), .B(n56705), .Z(n16317) );
  NANDN U34517 ( .A(y[4468]), .B(x[4468]), .Z(n16316) );
  NANDN U34518 ( .A(y[4469]), .B(x[4469]), .Z(n41464) );
  AND U34519 ( .A(n16316), .B(n41464), .Z(n56706) );
  NANDN U34520 ( .A(n16317), .B(n56706), .Z(n16318) );
  NANDN U34521 ( .A(n56707), .B(n16318), .Z(n16319) );
  AND U34522 ( .A(n56709), .B(n16319), .Z(n16320) );
  XNOR U34523 ( .A(y[4472]), .B(x[4472]), .Z(n41471) );
  NANDN U34524 ( .A(x[4471]), .B(y[4471]), .Z(n25098) );
  NAND U34525 ( .A(n41471), .B(n25098), .Z(n56710) );
  OR U34526 ( .A(n16320), .B(n56710), .Z(n16321) );
  NAND U34527 ( .A(n56712), .B(n16321), .Z(n16322) );
  NANDN U34528 ( .A(n51615), .B(n16322), .Z(n16324) );
  NANDN U34529 ( .A(y[4474]), .B(x[4474]), .Z(n16323) );
  NANDN U34530 ( .A(y[4475]), .B(x[4475]), .Z(n41486) );
  AND U34531 ( .A(n16323), .B(n41486), .Z(n51614) );
  AND U34532 ( .A(n16324), .B(n51614), .Z(n16325) );
  XNOR U34533 ( .A(y[4476]), .B(x[4476]), .Z(n41485) );
  NANDN U34534 ( .A(x[4475]), .B(y[4475]), .Z(n25096) );
  AND U34535 ( .A(n41485), .B(n25096), .Z(n56713) );
  NANDN U34536 ( .A(n16325), .B(n56713), .Z(n16326) );
  NANDN U34537 ( .A(n56714), .B(n16326), .Z(n16327) );
  AND U34538 ( .A(n51612), .B(n16327), .Z(n16328) );
  NAND U34539 ( .A(n41491), .B(n16328), .Z(n16329) );
  NANDN U34540 ( .A(n56715), .B(n16329), .Z(n16330) );
  AND U34541 ( .A(n56716), .B(n16330), .Z(n16331) );
  OR U34542 ( .A(n56717), .B(n16331), .Z(n16332) );
  NAND U34543 ( .A(n56718), .B(n16332), .Z(n16333) );
  NANDN U34544 ( .A(n56719), .B(n16333), .Z(n16334) );
  AND U34545 ( .A(n56720), .B(n16334), .Z(n16336) );
  NANDN U34546 ( .A(y[4484]), .B(x[4484]), .Z(n16335) );
  NANDN U34547 ( .A(y[4485]), .B(x[4485]), .Z(n25085) );
  NAND U34548 ( .A(n16335), .B(n25085), .Z(n56721) );
  OR U34549 ( .A(n16336), .B(n56721), .Z(n16337) );
  NAND U34550 ( .A(n16338), .B(n16337), .Z(n16340) );
  NANDN U34551 ( .A(y[4486]), .B(x[4486]), .Z(n16339) );
  NANDN U34552 ( .A(y[4487]), .B(x[4487]), .Z(n25084) );
  AND U34553 ( .A(n16339), .B(n25084), .Z(n51611) );
  AND U34554 ( .A(n16340), .B(n51611), .Z(n16341) );
  NANDN U34555 ( .A(x[4488]), .B(y[4488]), .Z(n25083) );
  ANDN U34556 ( .B(y[4487]), .A(x[4487]), .Z(n41515) );
  ANDN U34557 ( .B(n25083), .A(n41515), .Z(n56726) );
  NANDN U34558 ( .A(n16341), .B(n56726), .Z(n16342) );
  NAND U34559 ( .A(n16343), .B(n16342), .Z(n16344) );
  AND U34560 ( .A(n56728), .B(n16344), .Z(n16345) );
  NANDN U34561 ( .A(x[4490]), .B(y[4490]), .Z(n25079) );
  NAND U34562 ( .A(n16345), .B(n25079), .Z(n16346) );
  NANDN U34563 ( .A(y[4491]), .B(x[4491]), .Z(n56731) );
  AND U34564 ( .A(n16346), .B(n56731), .Z(n16347) );
  NANDN U34565 ( .A(n25081), .B(n16347), .Z(n16349) );
  NANDN U34566 ( .A(x[4492]), .B(y[4492]), .Z(n25077) );
  NANDN U34567 ( .A(x[4493]), .B(y[4493]), .Z(n25076) );
  NANDN U34568 ( .A(x[4494]), .B(y[4494]), .Z(n25073) );
  NAND U34569 ( .A(n25076), .B(n25073), .Z(n16351) );
  ANDN U34570 ( .B(n25077), .A(n16351), .Z(n56732) );
  NANDN U34571 ( .A(x[4491]), .B(y[4491]), .Z(n25080) );
  AND U34572 ( .A(n56732), .B(n25080), .Z(n16348) );
  NAND U34573 ( .A(n16349), .B(n16348), .Z(n16354) );
  NANDN U34574 ( .A(y[4493]), .B(x[4493]), .Z(n25074) );
  NANDN U34575 ( .A(y[4492]), .B(x[4492]), .Z(n25078) );
  NAND U34576 ( .A(n25074), .B(n25078), .Z(n16350) );
  NANDN U34577 ( .A(n16351), .B(n16350), .Z(n16352) );
  ANDN U34578 ( .B(x[4495]), .A(y[4495]), .Z(n41532) );
  ANDN U34579 ( .B(n16352), .A(n41532), .Z(n16353) );
  NANDN U34580 ( .A(y[4494]), .B(x[4494]), .Z(n25075) );
  AND U34581 ( .A(n16353), .B(n25075), .Z(n56733) );
  AND U34582 ( .A(n16354), .B(n56733), .Z(n16355) );
  XNOR U34583 ( .A(y[4496]), .B(x[4496]), .Z(n41533) );
  NANDN U34584 ( .A(x[4495]), .B(y[4495]), .Z(n25072) );
  NAND U34585 ( .A(n41533), .B(n25072), .Z(n56734) );
  OR U34586 ( .A(n16355), .B(n56734), .Z(n16356) );
  NAND U34587 ( .A(n56735), .B(n16356), .Z(n16357) );
  NANDN U34588 ( .A(n51610), .B(n16357), .Z(n16358) );
  AND U34589 ( .A(n56736), .B(n16358), .Z(n16359) );
  XNOR U34590 ( .A(y[4500]), .B(x[4500]), .Z(n41549) );
  NANDN U34591 ( .A(x[4499]), .B(y[4499]), .Z(n41543) );
  AND U34592 ( .A(n41549), .B(n41543), .Z(n56738) );
  NANDN U34593 ( .A(n16359), .B(n56738), .Z(n16360) );
  AND U34594 ( .A(n56739), .B(n16360), .Z(n16361) );
  OR U34595 ( .A(n56740), .B(n16361), .Z(n16362) );
  NAND U34596 ( .A(n56741), .B(n16362), .Z(n16363) );
  NANDN U34597 ( .A(n56742), .B(n16363), .Z(n16364) );
  AND U34598 ( .A(n56743), .B(n16364), .Z(n16365) );
  NANDN U34599 ( .A(x[4505]), .B(y[4505]), .Z(n25068) );
  NANDN U34600 ( .A(x[4506]), .B(y[4506]), .Z(n41571) );
  NAND U34601 ( .A(n25068), .B(n41571), .Z(n56744) );
  OR U34602 ( .A(n16365), .B(n56744), .Z(n16366) );
  AND U34603 ( .A(n56745), .B(n16366), .Z(n16367) );
  OR U34604 ( .A(n56746), .B(n16367), .Z(n16368) );
  NAND U34605 ( .A(n56747), .B(n16368), .Z(n16369) );
  NANDN U34606 ( .A(n56748), .B(n16369), .Z(n16370) );
  AND U34607 ( .A(n56749), .B(n16370), .Z(n16371) );
  XNOR U34608 ( .A(y[4512]), .B(x[4512]), .Z(n41586) );
  NANDN U34609 ( .A(x[4511]), .B(y[4511]), .Z(n41582) );
  AND U34610 ( .A(n41586), .B(n41582), .Z(n51609) );
  NANDN U34611 ( .A(n16371), .B(n51609), .Z(n16372) );
  NANDN U34612 ( .A(n56750), .B(n16372), .Z(n16373) );
  XNOR U34613 ( .A(y[4514]), .B(x[4514]), .Z(n41592) );
  NANDN U34614 ( .A(x[4513]), .B(y[4513]), .Z(n25060) );
  AND U34615 ( .A(n41592), .B(n25060), .Z(n56751) );
  AND U34616 ( .A(n16373), .B(n56751), .Z(n16375) );
  NANDN U34617 ( .A(y[4514]), .B(x[4514]), .Z(n16374) );
  NANDN U34618 ( .A(y[4515]), .B(x[4515]), .Z(n25056) );
  NAND U34619 ( .A(n16374), .B(n25056), .Z(n51608) );
  OR U34620 ( .A(n16375), .B(n51608), .Z(n16376) );
  NAND U34621 ( .A(n51607), .B(n16376), .Z(n16377) );
  NANDN U34622 ( .A(n56754), .B(n16377), .Z(n16378) );
  AND U34623 ( .A(n25054), .B(n16378), .Z(n16379) );
  NANDN U34624 ( .A(x[4517]), .B(y[4517]), .Z(n56755) );
  AND U34625 ( .A(n16379), .B(n56755), .Z(n16381) );
  NANDN U34626 ( .A(y[4518]), .B(x[4518]), .Z(n16380) );
  NANDN U34627 ( .A(y[4519]), .B(x[4519]), .Z(n41606) );
  NAND U34628 ( .A(n16380), .B(n41606), .Z(n56757) );
  OR U34629 ( .A(n16381), .B(n56757), .Z(n16382) );
  AND U34630 ( .A(n56758), .B(n16382), .Z(n16384) );
  NANDN U34631 ( .A(y[4520]), .B(x[4520]), .Z(n16383) );
  NANDN U34632 ( .A(y[4521]), .B(x[4521]), .Z(n41613) );
  NAND U34633 ( .A(n16383), .B(n41613), .Z(n51606) );
  OR U34634 ( .A(n16384), .B(n51606), .Z(n16385) );
  NAND U34635 ( .A(n51605), .B(n16385), .Z(n16386) );
  NANDN U34636 ( .A(n56759), .B(n16386), .Z(n16387) );
  NAND U34637 ( .A(n56760), .B(n16387), .Z(n16388) );
  NAND U34638 ( .A(n56761), .B(n16388), .Z(n16389) );
  NANDN U34639 ( .A(n56762), .B(n16389), .Z(n16390) );
  AND U34640 ( .A(n56763), .B(n16390), .Z(n16391) );
  OR U34641 ( .A(n56764), .B(n16391), .Z(n16392) );
  NAND U34642 ( .A(n56766), .B(n16392), .Z(n16393) );
  NAND U34643 ( .A(n41639), .B(n16393), .Z(n16394) );
  ANDN U34644 ( .B(y[4529]), .A(x[4529]), .Z(n25045) );
  OR U34645 ( .A(n16394), .B(n25045), .Z(n16395) );
  NAND U34646 ( .A(n56772), .B(n16395), .Z(n16397) );
  XNOR U34647 ( .A(x[4532]), .B(y[4532]), .Z(n41646) );
  NANDN U34648 ( .A(x[4531]), .B(y[4531]), .Z(n56774) );
  NAND U34649 ( .A(n41646), .B(n56774), .Z(n16396) );
  ANDN U34650 ( .B(n16397), .A(n16396), .Z(n16398) );
  OR U34651 ( .A(n56777), .B(n16398), .Z(n16399) );
  NAND U34652 ( .A(n56780), .B(n16399), .Z(n16400) );
  NANDN U34653 ( .A(n56782), .B(n16400), .Z(n16401) );
  AND U34654 ( .A(n56784), .B(n16401), .Z(n16403) );
  NANDN U34655 ( .A(y[4536]), .B(x[4536]), .Z(n16402) );
  NANDN U34656 ( .A(y[4537]), .B(x[4537]), .Z(n25039) );
  NAND U34657 ( .A(n16402), .B(n25039), .Z(n56786) );
  OR U34658 ( .A(n16403), .B(n56786), .Z(n16404) );
  AND U34659 ( .A(n16405), .B(n16404), .Z(n16406) );
  OR U34660 ( .A(n56791), .B(n16406), .Z(n16407) );
  NAND U34661 ( .A(n56794), .B(n16407), .Z(n16408) );
  NANDN U34662 ( .A(n56796), .B(n16408), .Z(n16409) );
  AND U34663 ( .A(n56798), .B(n16409), .Z(n16410) );
  NANDN U34664 ( .A(y[4542]), .B(x[4542]), .Z(n41672) );
  NANDN U34665 ( .A(y[4543]), .B(x[4543]), .Z(n41678) );
  NAND U34666 ( .A(n41672), .B(n41678), .Z(n56800) );
  OR U34667 ( .A(n16410), .B(n56800), .Z(n16411) );
  AND U34668 ( .A(n56802), .B(n16411), .Z(n16412) );
  OR U34669 ( .A(n56804), .B(n16412), .Z(n16413) );
  NAND U34670 ( .A(n56806), .B(n16413), .Z(n16414) );
  NANDN U34671 ( .A(n56807), .B(n16414), .Z(n16415) );
  AND U34672 ( .A(n25030), .B(n16415), .Z(n16416) );
  NANDN U34673 ( .A(x[4547]), .B(y[4547]), .Z(n56808) );
  AND U34674 ( .A(n16416), .B(n56808), .Z(n16418) );
  NANDN U34675 ( .A(y[4548]), .B(x[4548]), .Z(n16417) );
  NANDN U34676 ( .A(y[4549]), .B(x[4549]), .Z(n25027) );
  NAND U34677 ( .A(n16417), .B(n25027), .Z(n56810) );
  OR U34678 ( .A(n16418), .B(n56810), .Z(n16419) );
  AND U34679 ( .A(n16420), .B(n16419), .Z(n16422) );
  NANDN U34680 ( .A(y[4550]), .B(x[4550]), .Z(n16421) );
  NANDN U34681 ( .A(y[4551]), .B(x[4551]), .Z(n41700) );
  AND U34682 ( .A(n16421), .B(n41700), .Z(n56813) );
  NANDN U34683 ( .A(n16422), .B(n56813), .Z(n16423) );
  AND U34684 ( .A(n41699), .B(n16423), .Z(n16424) );
  ANDN U34685 ( .B(y[4551]), .A(x[4551]), .Z(n51603) );
  ANDN U34686 ( .B(n16424), .A(n51603), .Z(n16425) );
  OR U34687 ( .A(n56814), .B(n16425), .Z(n16426) );
  NAND U34688 ( .A(n56815), .B(n16426), .Z(n16427) );
  NANDN U34689 ( .A(n56816), .B(n16427), .Z(n16428) );
  AND U34690 ( .A(n56817), .B(n16428), .Z(n16430) );
  NANDN U34691 ( .A(y[4556]), .B(x[4556]), .Z(n16429) );
  NANDN U34692 ( .A(y[4557]), .B(x[4557]), .Z(n25022) );
  NAND U34693 ( .A(n16429), .B(n25022), .Z(n56818) );
  OR U34694 ( .A(n16430), .B(n56818), .Z(n16431) );
  AND U34695 ( .A(n56819), .B(n16431), .Z(n16432) );
  OR U34696 ( .A(n56820), .B(n16432), .Z(n16433) );
  NAND U34697 ( .A(n56822), .B(n16433), .Z(n16434) );
  NANDN U34698 ( .A(n56823), .B(n16434), .Z(n16435) );
  AND U34699 ( .A(n56824), .B(n16435), .Z(n16437) );
  NANDN U34700 ( .A(y[4562]), .B(x[4562]), .Z(n16436) );
  NANDN U34701 ( .A(y[4563]), .B(x[4563]), .Z(n25016) );
  NAND U34702 ( .A(n16436), .B(n25016), .Z(n56825) );
  OR U34703 ( .A(n16437), .B(n56825), .Z(n16438) );
  NAND U34704 ( .A(n16439), .B(n16438), .Z(n16440) );
  AND U34705 ( .A(n56826), .B(n16440), .Z(n16441) );
  ANDN U34706 ( .B(n56828), .A(n16441), .Z(n16442) );
  NAND U34707 ( .A(n25015), .B(n16442), .Z(n16443) );
  NANDN U34708 ( .A(n56829), .B(n16443), .Z(n16444) );
  AND U34709 ( .A(n25013), .B(n16444), .Z(n16445) );
  NANDN U34710 ( .A(x[4567]), .B(y[4567]), .Z(n56830) );
  AND U34711 ( .A(n16445), .B(n56830), .Z(n16446) );
  OR U34712 ( .A(n56832), .B(n16446), .Z(n16447) );
  AND U34713 ( .A(n41748), .B(n16447), .Z(n16448) );
  ANDN U34714 ( .B(y[4569]), .A(x[4569]), .Z(n56833) );
  ANDN U34715 ( .B(n16448), .A(n56833), .Z(n16450) );
  NANDN U34716 ( .A(y[4570]), .B(x[4570]), .Z(n16449) );
  NANDN U34717 ( .A(y[4571]), .B(x[4571]), .Z(n41755) );
  NAND U34718 ( .A(n16449), .B(n41755), .Z(n56835) );
  OR U34719 ( .A(n16450), .B(n56835), .Z(n16451) );
  AND U34720 ( .A(n56836), .B(n16451), .Z(n16452) );
  NANDN U34721 ( .A(y[4572]), .B(x[4572]), .Z(n41754) );
  NANDN U34722 ( .A(y[4573]), .B(x[4573]), .Z(n41761) );
  AND U34723 ( .A(n41754), .B(n41761), .Z(n56837) );
  NANDN U34724 ( .A(n16452), .B(n56837), .Z(n16453) );
  NANDN U34725 ( .A(n16454), .B(n16453), .Z(n16455) );
  AND U34726 ( .A(n56842), .B(n16455), .Z(n16456) );
  OR U34727 ( .A(n56843), .B(n16456), .Z(n16457) );
  NAND U34728 ( .A(n56844), .B(n16457), .Z(n16458) );
  NANDN U34729 ( .A(n56845), .B(n16458), .Z(n16459) );
  NAND U34730 ( .A(n56846), .B(n16459), .Z(n16460) );
  XNOR U34731 ( .A(y[4580]), .B(x[4580]), .Z(n41784) );
  NANDN U34732 ( .A(x[4579]), .B(y[4579]), .Z(n41778) );
  AND U34733 ( .A(n41784), .B(n41778), .Z(n56847) );
  AND U34734 ( .A(n16460), .B(n56847), .Z(n16461) );
  ANDN U34735 ( .B(n56848), .A(n16461), .Z(n16462) );
  OR U34736 ( .A(n56849), .B(n16462), .Z(n16463) );
  NAND U34737 ( .A(n56850), .B(n16463), .Z(n16464) );
  NANDN U34738 ( .A(n56851), .B(n16464), .Z(n16465) );
  AND U34739 ( .A(n56852), .B(n16465), .Z(n16466) );
  ANDN U34740 ( .B(n56854), .A(n16466), .Z(n16468) );
  NAND U34741 ( .A(n16468), .B(n16467), .Z(n16469) );
  NANDN U34742 ( .A(n56855), .B(n16469), .Z(n16470) );
  AND U34743 ( .A(n25007), .B(n16470), .Z(n16471) );
  NANDN U34744 ( .A(n56856), .B(n16471), .Z(n16472) );
  NANDN U34745 ( .A(n56858), .B(n16472), .Z(n16473) );
  AND U34746 ( .A(n56860), .B(n16473), .Z(n16474) );
  OR U34747 ( .A(n56861), .B(n16474), .Z(n16475) );
  NAND U34748 ( .A(n56862), .B(n16475), .Z(n16476) );
  NANDN U34749 ( .A(n56863), .B(n16476), .Z(n16477) );
  AND U34750 ( .A(n56864), .B(n16477), .Z(n16479) );
  NANDN U34751 ( .A(y[4594]), .B(x[4594]), .Z(n16478) );
  NANDN U34752 ( .A(y[4595]), .B(x[4595]), .Z(n24998) );
  AND U34753 ( .A(n16478), .B(n24998), .Z(n56865) );
  NANDN U34754 ( .A(n16479), .B(n56865), .Z(n16480) );
  XNOR U34755 ( .A(y[4596]), .B(x[4596]), .Z(n24999) );
  NANDN U34756 ( .A(x[4595]), .B(y[4595]), .Z(n25000) );
  AND U34757 ( .A(n24999), .B(n25000), .Z(n51600) );
  AND U34758 ( .A(n16480), .B(n51600), .Z(n16482) );
  NANDN U34759 ( .A(y[4596]), .B(x[4596]), .Z(n16481) );
  NANDN U34760 ( .A(y[4597]), .B(x[4597]), .Z(n24994) );
  NAND U34761 ( .A(n16481), .B(n24994), .Z(n56866) );
  OR U34762 ( .A(n16482), .B(n56866), .Z(n16483) );
  NAND U34763 ( .A(n56867), .B(n16483), .Z(n16484) );
  NANDN U34764 ( .A(n51599), .B(n16484), .Z(n16485) );
  XNOR U34765 ( .A(y[4600]), .B(x[4600]), .Z(n24993) );
  NANDN U34766 ( .A(x[4599]), .B(y[4599]), .Z(n41838) );
  AND U34767 ( .A(n24993), .B(n41838), .Z(n51598) );
  AND U34768 ( .A(n16485), .B(n51598), .Z(n16487) );
  NANDN U34769 ( .A(y[4600]), .B(x[4600]), .Z(n16486) );
  NANDN U34770 ( .A(y[4601]), .B(x[4601]), .Z(n41848) );
  NAND U34771 ( .A(n16486), .B(n41848), .Z(n56868) );
  OR U34772 ( .A(n16487), .B(n56868), .Z(n16488) );
  XNOR U34773 ( .A(y[4602]), .B(x[4602]), .Z(n41849) );
  NANDN U34774 ( .A(x[4601]), .B(y[4601]), .Z(n41845) );
  AND U34775 ( .A(n41849), .B(n41845), .Z(n56869) );
  AND U34776 ( .A(n16488), .B(n56869), .Z(n16490) );
  NANDN U34777 ( .A(y[4602]), .B(x[4602]), .Z(n16489) );
  NANDN U34778 ( .A(y[4603]), .B(x[4603]), .Z(n41854) );
  NAND U34779 ( .A(n16489), .B(n41854), .Z(n56870) );
  OR U34780 ( .A(n16490), .B(n56870), .Z(n16491) );
  NAND U34781 ( .A(n56873), .B(n16491), .Z(n16492) );
  NANDN U34782 ( .A(n51597), .B(n16492), .Z(n16493) );
  XNOR U34783 ( .A(y[4606]), .B(x[4606]), .Z(n41861) );
  NANDN U34784 ( .A(x[4605]), .B(y[4605]), .Z(n24988) );
  AND U34785 ( .A(n41861), .B(n24988), .Z(n51596) );
  AND U34786 ( .A(n16493), .B(n51596), .Z(n16495) );
  NANDN U34787 ( .A(y[4606]), .B(x[4606]), .Z(n16494) );
  NANDN U34788 ( .A(y[4607]), .B(x[4607]), .Z(n41866) );
  AND U34789 ( .A(n16494), .B(n41866), .Z(n56875) );
  NANDN U34790 ( .A(n16495), .B(n56875), .Z(n16496) );
  AND U34791 ( .A(n16497), .B(n16496), .Z(n16498) );
  OR U34792 ( .A(n56878), .B(n16498), .Z(n16499) );
  NAND U34793 ( .A(n56879), .B(n16499), .Z(n16500) );
  NANDN U34794 ( .A(n56880), .B(n16500), .Z(n16501) );
  AND U34795 ( .A(n24982), .B(n16501), .Z(n16502) );
  NANDN U34796 ( .A(x[4611]), .B(y[4611]), .Z(n51594) );
  AND U34797 ( .A(n16502), .B(n51594), .Z(n16504) );
  NANDN U34798 ( .A(y[4612]), .B(x[4612]), .Z(n16503) );
  NANDN U34799 ( .A(y[4613]), .B(x[4613]), .Z(n41883) );
  NAND U34800 ( .A(n16503), .B(n41883), .Z(n56881) );
  OR U34801 ( .A(n16504), .B(n56881), .Z(n16505) );
  AND U34802 ( .A(n56882), .B(n16505), .Z(n16506) );
  NANDN U34803 ( .A(y[4614]), .B(x[4614]), .Z(n41882) );
  ANDN U34804 ( .B(x[4615]), .A(y[4615]), .Z(n41890) );
  ANDN U34805 ( .B(n41882), .A(n41890), .Z(n56883) );
  NANDN U34806 ( .A(n16506), .B(n56883), .Z(n16507) );
  NAND U34807 ( .A(n56885), .B(n16507), .Z(n16508) );
  NANDN U34808 ( .A(n56886), .B(n16508), .Z(n16509) );
  AND U34809 ( .A(n24977), .B(n16509), .Z(n16510) );
  NANDN U34810 ( .A(x[4617]), .B(y[4617]), .Z(n51592) );
  AND U34811 ( .A(n16510), .B(n51592), .Z(n16512) );
  ANDN U34812 ( .B(x[4619]), .A(y[4619]), .Z(n41898) );
  NANDN U34813 ( .A(y[4618]), .B(x[4618]), .Z(n16511) );
  NANDN U34814 ( .A(n41898), .B(n16511), .Z(n56888) );
  OR U34815 ( .A(n16512), .B(n56888), .Z(n16513) );
  AND U34816 ( .A(n16514), .B(n16513), .Z(n16516) );
  NANDN U34817 ( .A(y[4620]), .B(x[4620]), .Z(n16515) );
  NANDN U34818 ( .A(y[4621]), .B(x[4621]), .Z(n41904) );
  NAND U34819 ( .A(n16515), .B(n41904), .Z(n56891) );
  OR U34820 ( .A(n16516), .B(n56891), .Z(n16517) );
  NAND U34821 ( .A(n56892), .B(n16517), .Z(n16518) );
  NANDN U34822 ( .A(n51591), .B(n16518), .Z(n16519) );
  XNOR U34823 ( .A(y[4624]), .B(x[4624]), .Z(n24974) );
  NANDN U34824 ( .A(x[4623]), .B(y[4623]), .Z(n41908) );
  AND U34825 ( .A(n24974), .B(n41908), .Z(n51590) );
  AND U34826 ( .A(n16519), .B(n51590), .Z(n16521) );
  ANDN U34827 ( .B(x[4625]), .A(y[4625]), .Z(n41919) );
  NANDN U34828 ( .A(y[4624]), .B(x[4624]), .Z(n16520) );
  NANDN U34829 ( .A(n41919), .B(n16520), .Z(n56893) );
  OR U34830 ( .A(n16521), .B(n56893), .Z(n16522) );
  XNOR U34831 ( .A(y[4626]), .B(x[4626]), .Z(n41920) );
  NANDN U34832 ( .A(x[4625]), .B(y[4625]), .Z(n41914) );
  AND U34833 ( .A(n41920), .B(n41914), .Z(n56894) );
  AND U34834 ( .A(n16522), .B(n56894), .Z(n16524) );
  ANDN U34835 ( .B(x[4627]), .A(y[4627]), .Z(n41927) );
  NANDN U34836 ( .A(y[4626]), .B(x[4626]), .Z(n16523) );
  NANDN U34837 ( .A(n41927), .B(n16523), .Z(n56897) );
  OR U34838 ( .A(n16524), .B(n56897), .Z(n16525) );
  NAND U34839 ( .A(n56898), .B(n16525), .Z(n16526) );
  NANDN U34840 ( .A(n51589), .B(n16526), .Z(n16527) );
  XNOR U34841 ( .A(y[4630]), .B(x[4630]), .Z(n41936) );
  NANDN U34842 ( .A(x[4629]), .B(y[4629]), .Z(n41930) );
  AND U34843 ( .A(n41936), .B(n41930), .Z(n51588) );
  AND U34844 ( .A(n16527), .B(n51588), .Z(n16529) );
  NANDN U34845 ( .A(y[4630]), .B(x[4630]), .Z(n16528) );
  ANDN U34846 ( .B(x[4631]), .A(y[4631]), .Z(n41943) );
  ANDN U34847 ( .B(n16528), .A(n41943), .Z(n56899) );
  NANDN U34848 ( .A(n16529), .B(n56899), .Z(n16530) );
  NANDN U34849 ( .A(n56900), .B(n16530), .Z(n16531) );
  AND U34850 ( .A(n56901), .B(n16531), .Z(n16532) );
  OR U34851 ( .A(n56902), .B(n16532), .Z(n16533) );
  NAND U34852 ( .A(n56903), .B(n16533), .Z(n16534) );
  NANDN U34853 ( .A(n56904), .B(n16534), .Z(n16535) );
  AND U34854 ( .A(n56905), .B(n16535), .Z(n16536) );
  NANDN U34855 ( .A(x[4637]), .B(y[4637]), .Z(n56906) );
  NANDN U34856 ( .A(n16536), .B(n56906), .Z(n16537) );
  NAND U34857 ( .A(n41963), .B(n16537), .Z(n16538) );
  NAND U34858 ( .A(n56908), .B(n16538), .Z(n16539) );
  NANDN U34859 ( .A(y[4639]), .B(x[4639]), .Z(n51587) );
  AND U34860 ( .A(n16539), .B(n51587), .Z(n16540) );
  NANDN U34861 ( .A(y[4638]), .B(x[4638]), .Z(n41962) );
  AND U34862 ( .A(n16540), .B(n41962), .Z(n16541) );
  XNOR U34863 ( .A(y[4640]), .B(x[4640]), .Z(n24971) );
  NANDN U34864 ( .A(x[4639]), .B(y[4639]), .Z(n41966) );
  NAND U34865 ( .A(n24971), .B(n41966), .Z(n56911) );
  OR U34866 ( .A(n16541), .B(n56911), .Z(n16542) );
  NAND U34867 ( .A(n56912), .B(n16542), .Z(n16543) );
  AND U34868 ( .A(n56913), .B(n16543), .Z(n16545) );
  NANDN U34869 ( .A(y[4642]), .B(x[4642]), .Z(n16544) );
  NANDN U34870 ( .A(y[4643]), .B(x[4643]), .Z(n41978) );
  AND U34871 ( .A(n16544), .B(n41978), .Z(n51586) );
  NANDN U34872 ( .A(n16545), .B(n51586), .Z(n16546) );
  NAND U34873 ( .A(n16547), .B(n16546), .Z(n16548) );
  AND U34874 ( .A(n56916), .B(n16548), .Z(n16549) );
  ANDN U34875 ( .B(n51584), .A(n16549), .Z(n16550) );
  NAND U34876 ( .A(n24967), .B(n16550), .Z(n16551) );
  NANDN U34877 ( .A(n24964), .B(n16551), .Z(n16552) );
  ANDN U34878 ( .B(x[4646]), .A(y[4646]), .Z(n56917) );
  OR U34879 ( .A(n16552), .B(n56917), .Z(n16553) );
  NAND U34880 ( .A(n16554), .B(n16553), .Z(n16555) );
  NANDN U34881 ( .A(n16556), .B(n16555), .Z(n16557) );
  XNOR U34882 ( .A(y[4650]), .B(x[4650]), .Z(n41993) );
  NANDN U34883 ( .A(x[4649]), .B(y[4649]), .Z(n41989) );
  AND U34884 ( .A(n41993), .B(n41989), .Z(n56922) );
  AND U34885 ( .A(n16557), .B(n56922), .Z(n16559) );
  NANDN U34886 ( .A(y[4650]), .B(x[4650]), .Z(n16558) );
  NANDN U34887 ( .A(y[4651]), .B(x[4651]), .Z(n24961) );
  NAND U34888 ( .A(n16558), .B(n24961), .Z(n51582) );
  OR U34889 ( .A(n16559), .B(n51582), .Z(n16560) );
  AND U34890 ( .A(n16561), .B(n16560), .Z(n16562) );
  OR U34891 ( .A(n56926), .B(n16562), .Z(n16563) );
  NAND U34892 ( .A(n56927), .B(n16563), .Z(n16564) );
  NANDN U34893 ( .A(n56928), .B(n16564), .Z(n16565) );
  AND U34894 ( .A(n56929), .B(n16565), .Z(n16567) );
  ANDN U34895 ( .B(x[4657]), .A(y[4657]), .Z(n42019) );
  NANDN U34896 ( .A(y[4656]), .B(x[4656]), .Z(n16566) );
  NANDN U34897 ( .A(n42019), .B(n16566), .Z(n56930) );
  OR U34898 ( .A(n16567), .B(n56930), .Z(n16568) );
  AND U34899 ( .A(n56931), .B(n16568), .Z(n16569) );
  OR U34900 ( .A(n56932), .B(n16569), .Z(n16570) );
  NAND U34901 ( .A(n56933), .B(n16570), .Z(n16571) );
  NANDN U34902 ( .A(n56934), .B(n16571), .Z(n16572) );
  AND U34903 ( .A(n24958), .B(n16572), .Z(n16573) );
  ANDN U34904 ( .B(y[4661]), .A(x[4661]), .Z(n56935) );
  ANDN U34905 ( .B(n16573), .A(n56935), .Z(n16575) );
  NANDN U34906 ( .A(y[4662]), .B(x[4662]), .Z(n16574) );
  NANDN U34907 ( .A(y[4663]), .B(x[4663]), .Z(n24956) );
  NAND U34908 ( .A(n16574), .B(n24956), .Z(n56936) );
  OR U34909 ( .A(n16575), .B(n56936), .Z(n16576) );
  AND U34910 ( .A(n56938), .B(n16576), .Z(n16577) );
  OR U34911 ( .A(n56939), .B(n16577), .Z(n16578) );
  NAND U34912 ( .A(n56940), .B(n16578), .Z(n16579) );
  NANDN U34913 ( .A(n56941), .B(n16579), .Z(n16580) );
  AND U34914 ( .A(n56942), .B(n16580), .Z(n16582) );
  NANDN U34915 ( .A(y[4668]), .B(x[4668]), .Z(n16581) );
  NANDN U34916 ( .A(y[4669]), .B(x[4669]), .Z(n42054) );
  NAND U34917 ( .A(n16581), .B(n42054), .Z(n56943) );
  OR U34918 ( .A(n16582), .B(n56943), .Z(n16583) );
  AND U34919 ( .A(n56944), .B(n16583), .Z(n16584) );
  OR U34920 ( .A(n56945), .B(n16584), .Z(n16585) );
  NAND U34921 ( .A(n56946), .B(n16585), .Z(n16586) );
  NANDN U34922 ( .A(n56947), .B(n16586), .Z(n16587) );
  AND U34923 ( .A(n56948), .B(n16587), .Z(n16589) );
  NANDN U34924 ( .A(y[4674]), .B(x[4674]), .Z(n16588) );
  NANDN U34925 ( .A(y[4675]), .B(x[4675]), .Z(n42072) );
  NAND U34926 ( .A(n16588), .B(n42072), .Z(n56949) );
  OR U34927 ( .A(n16589), .B(n56949), .Z(n16590) );
  AND U34928 ( .A(n16591), .B(n16590), .Z(n16593) );
  NANDN U34929 ( .A(y[4676]), .B(x[4676]), .Z(n16592) );
  NANDN U34930 ( .A(y[4677]), .B(x[4677]), .Z(n42078) );
  NAND U34931 ( .A(n16592), .B(n42078), .Z(n56950) );
  OR U34932 ( .A(n16593), .B(n56950), .Z(n16594) );
  NAND U34933 ( .A(n56951), .B(n16594), .Z(n16595) );
  NANDN U34934 ( .A(n56952), .B(n16595), .Z(n16596) );
  NAND U34935 ( .A(n24943), .B(n16596), .Z(n16597) );
  ANDN U34936 ( .B(y[4679]), .A(x[4679]), .Z(n56953) );
  OR U34937 ( .A(n16597), .B(n56953), .Z(n16598) );
  NAND U34938 ( .A(n56956), .B(n16598), .Z(n16600) );
  XNOR U34939 ( .A(x[4682]), .B(y[4682]), .Z(n42089) );
  NANDN U34940 ( .A(x[4681]), .B(y[4681]), .Z(n51577) );
  NAND U34941 ( .A(n42089), .B(n51577), .Z(n16599) );
  ANDN U34942 ( .B(n16600), .A(n16599), .Z(n16601) );
  OR U34943 ( .A(n56958), .B(n16601), .Z(n16602) );
  NAND U34944 ( .A(n56959), .B(n16602), .Z(n16603) );
  NANDN U34945 ( .A(n56960), .B(n16603), .Z(n16604) );
  AND U34946 ( .A(n56961), .B(n16604), .Z(n16606) );
  NANDN U34947 ( .A(y[4686]), .B(x[4686]), .Z(n16605) );
  NANDN U34948 ( .A(y[4687]), .B(x[4687]), .Z(n24935) );
  AND U34949 ( .A(n16605), .B(n24935), .Z(n56962) );
  NANDN U34950 ( .A(n16606), .B(n56962), .Z(n16607) );
  NAND U34951 ( .A(n16608), .B(n16607), .Z(n16609) );
  AND U34952 ( .A(n56963), .B(n16609), .Z(n16610) );
  ANDN U34953 ( .B(n56965), .A(n16610), .Z(n16611) );
  NAND U34954 ( .A(n42112), .B(n16611), .Z(n16612) );
  NANDN U34955 ( .A(n56966), .B(n16612), .Z(n16613) );
  AND U34956 ( .A(n24934), .B(n16613), .Z(n16614) );
  NANDN U34957 ( .A(n42114), .B(n16614), .Z(n16615) );
  NAND U34958 ( .A(n56969), .B(n16615), .Z(n16616) );
  NANDN U34959 ( .A(n56970), .B(n16616), .Z(n16617) );
  AND U34960 ( .A(n56972), .B(n16617), .Z(n16619) );
  XNOR U34961 ( .A(x[4696]), .B(y[4696]), .Z(n24930) );
  ANDN U34962 ( .B(y[4695]), .A(x[4695]), .Z(n56974) );
  ANDN U34963 ( .B(n24930), .A(n56974), .Z(n16618) );
  NANDN U34964 ( .A(n16619), .B(n16618), .Z(n16620) );
  AND U34965 ( .A(n56976), .B(n16620), .Z(n16621) );
  OR U34966 ( .A(n56977), .B(n16621), .Z(n16622) );
  NAND U34967 ( .A(n56978), .B(n16622), .Z(n16623) );
  NANDN U34968 ( .A(n56979), .B(n16623), .Z(n16624) );
  AND U34969 ( .A(n56980), .B(n16624), .Z(n16625) );
  XNOR U34970 ( .A(y[4702]), .B(x[4702]), .Z(n42144) );
  NANDN U34971 ( .A(x[4701]), .B(y[4701]), .Z(n24924) );
  NAND U34972 ( .A(n42144), .B(n24924), .Z(n56981) );
  OR U34973 ( .A(n16625), .B(n56981), .Z(n16626) );
  AND U34974 ( .A(n56982), .B(n16626), .Z(n16627) );
  OR U34975 ( .A(n56983), .B(n16627), .Z(n16628) );
  NAND U34976 ( .A(n56984), .B(n16628), .Z(n16629) );
  NANDN U34977 ( .A(n56985), .B(n16629), .Z(n16630) );
  AND U34978 ( .A(n56986), .B(n16630), .Z(n16632) );
  XNOR U34979 ( .A(x[4708]), .B(y[4708]), .Z(n24916) );
  NANDN U34980 ( .A(x[4707]), .B(y[4707]), .Z(n56988) );
  NAND U34981 ( .A(n24916), .B(n56988), .Z(n16631) );
  OR U34982 ( .A(n16632), .B(n16631), .Z(n16634) );
  NANDN U34983 ( .A(y[4708]), .B(x[4708]), .Z(n16633) );
  NANDN U34984 ( .A(y[4709]), .B(x[4709]), .Z(n42165) );
  AND U34985 ( .A(n16633), .B(n42165), .Z(n51574) );
  AND U34986 ( .A(n16634), .B(n51574), .Z(n16636) );
  XNOR U34987 ( .A(x[4710]), .B(y[4710]), .Z(n42164) );
  ANDN U34988 ( .B(y[4709]), .A(x[4709]), .Z(n56989) );
  ANDN U34989 ( .B(n42164), .A(n56989), .Z(n16635) );
  NANDN U34990 ( .A(n16636), .B(n16635), .Z(n16637) );
  NANDN U34991 ( .A(n56991), .B(n16637), .Z(n16638) );
  AND U34992 ( .A(n56993), .B(n16638), .Z(n16639) );
  OR U34993 ( .A(n56994), .B(n16639), .Z(n16640) );
  NAND U34994 ( .A(n56995), .B(n16640), .Z(n16641) );
  NANDN U34995 ( .A(n56996), .B(n16641), .Z(n16642) );
  AND U34996 ( .A(n56997), .B(n16642), .Z(n16644) );
  NANDN U34997 ( .A(y[4716]), .B(x[4716]), .Z(n16643) );
  NANDN U34998 ( .A(y[4717]), .B(x[4717]), .Z(n24909) );
  NAND U34999 ( .A(n16643), .B(n24909), .Z(n56998) );
  OR U35000 ( .A(n16644), .B(n56998), .Z(n16645) );
  AND U35001 ( .A(n56999), .B(n16645), .Z(n16646) );
  OR U35002 ( .A(n57000), .B(n16646), .Z(n16647) );
  NAND U35003 ( .A(n57001), .B(n16647), .Z(n16648) );
  NANDN U35004 ( .A(n57002), .B(n16648), .Z(n16649) );
  AND U35005 ( .A(n57003), .B(n16649), .Z(n16650) );
  NANDN U35006 ( .A(y[4722]), .B(x[4722]), .Z(n24902) );
  NANDN U35007 ( .A(y[4723]), .B(x[4723]), .Z(n24900) );
  NAND U35008 ( .A(n24902), .B(n24900), .Z(n57004) );
  OR U35009 ( .A(n16650), .B(n57004), .Z(n16651) );
  NAND U35010 ( .A(n16652), .B(n16651), .Z(n16654) );
  NANDN U35011 ( .A(y[4724]), .B(x[4724]), .Z(n16653) );
  NANDN U35012 ( .A(y[4725]), .B(x[4725]), .Z(n24897) );
  AND U35013 ( .A(n16653), .B(n24897), .Z(n51573) );
  AND U35014 ( .A(n16654), .B(n51573), .Z(n16655) );
  NOR U35015 ( .A(n24899), .B(n16655), .Z(n16656) );
  NAND U35016 ( .A(n24898), .B(n16656), .Z(n16657) );
  NANDN U35017 ( .A(n57009), .B(n16657), .Z(n16658) );
  AND U35018 ( .A(n24895), .B(n16658), .Z(n16659) );
  NANDN U35019 ( .A(n24896), .B(n16659), .Z(n16660) );
  NAND U35020 ( .A(n57012), .B(n16660), .Z(n16661) );
  NANDN U35021 ( .A(n42219), .B(n16661), .Z(n16662) );
  ANDN U35022 ( .B(y[4729]), .A(x[4729]), .Z(n24893) );
  OR U35023 ( .A(n16662), .B(n24893), .Z(n16663) );
  NAND U35024 ( .A(n51570), .B(n16663), .Z(n16665) );
  XNOR U35025 ( .A(x[4732]), .B(y[4732]), .Z(n24892) );
  NANDN U35026 ( .A(x[4731]), .B(y[4731]), .Z(n57015) );
  NAND U35027 ( .A(n24892), .B(n57015), .Z(n16664) );
  ANDN U35028 ( .B(n16665), .A(n16664), .Z(n16666) );
  OR U35029 ( .A(n57017), .B(n16666), .Z(n16667) );
  NAND U35030 ( .A(n57018), .B(n16667), .Z(n16668) );
  NANDN U35031 ( .A(n57019), .B(n16668), .Z(n16669) );
  AND U35032 ( .A(n57020), .B(n16669), .Z(n16671) );
  ANDN U35033 ( .B(x[4737]), .A(y[4737]), .Z(n42244) );
  NANDN U35034 ( .A(y[4736]), .B(x[4736]), .Z(n16670) );
  NANDN U35035 ( .A(n42244), .B(n16670), .Z(n57021) );
  OR U35036 ( .A(n16671), .B(n57021), .Z(n16672) );
  AND U35037 ( .A(n57022), .B(n16672), .Z(n16673) );
  OR U35038 ( .A(n57023), .B(n16673), .Z(n16674) );
  NAND U35039 ( .A(n57024), .B(n16674), .Z(n16675) );
  NANDN U35040 ( .A(n57025), .B(n16675), .Z(n16676) );
  AND U35041 ( .A(n57026), .B(n16676), .Z(n16678) );
  ANDN U35042 ( .B(x[4743]), .A(y[4743]), .Z(n42265) );
  NANDN U35043 ( .A(y[4742]), .B(x[4742]), .Z(n16677) );
  NANDN U35044 ( .A(n42265), .B(n16677), .Z(n57027) );
  OR U35045 ( .A(n16678), .B(n57027), .Z(n16679) );
  AND U35046 ( .A(n16680), .B(n16679), .Z(n16681) );
  OR U35047 ( .A(n57031), .B(n16681), .Z(n16682) );
  NAND U35048 ( .A(n57032), .B(n16682), .Z(n16683) );
  NANDN U35049 ( .A(n57033), .B(n16683), .Z(n16684) );
  AND U35050 ( .A(n24886), .B(n16684), .Z(n16685) );
  NANDN U35051 ( .A(x[4747]), .B(y[4747]), .Z(n57034) );
  AND U35052 ( .A(n16685), .B(n57034), .Z(n16687) );
  NANDN U35053 ( .A(y[4748]), .B(x[4748]), .Z(n16686) );
  NANDN U35054 ( .A(y[4749]), .B(x[4749]), .Z(n24883) );
  NAND U35055 ( .A(n16686), .B(n24883), .Z(n51569) );
  OR U35056 ( .A(n16687), .B(n51569), .Z(n16688) );
  XNOR U35057 ( .A(y[4750]), .B(x[4750]), .Z(n24884) );
  NANDN U35058 ( .A(x[4749]), .B(y[4749]), .Z(n42279) );
  AND U35059 ( .A(n24884), .B(n42279), .Z(n57036) );
  AND U35060 ( .A(n16688), .B(n57036), .Z(n16690) );
  NANDN U35061 ( .A(y[4750]), .B(x[4750]), .Z(n16689) );
  NANDN U35062 ( .A(y[4751]), .B(x[4751]), .Z(n42285) );
  NAND U35063 ( .A(n16689), .B(n42285), .Z(n51568) );
  OR U35064 ( .A(n16690), .B(n51568), .Z(n16691) );
  NAND U35065 ( .A(n51567), .B(n16691), .Z(n16692) );
  NANDN U35066 ( .A(n57037), .B(n16692), .Z(n16693) );
  XNOR U35067 ( .A(y[4754]), .B(x[4754]), .Z(n42292) );
  NANDN U35068 ( .A(x[4753]), .B(y[4753]), .Z(n24879) );
  AND U35069 ( .A(n42292), .B(n24879), .Z(n57038) );
  AND U35070 ( .A(n16693), .B(n57038), .Z(n16695) );
  NANDN U35071 ( .A(y[4754]), .B(x[4754]), .Z(n16694) );
  NANDN U35072 ( .A(y[4755]), .B(x[4755]), .Z(n42297) );
  AND U35073 ( .A(n16694), .B(n42297), .Z(n57039) );
  NANDN U35074 ( .A(n16695), .B(n57039), .Z(n16696) );
  NANDN U35075 ( .A(n57040), .B(n16696), .Z(n16697) );
  AND U35076 ( .A(n57042), .B(n16697), .Z(n16698) );
  OR U35077 ( .A(n57043), .B(n16698), .Z(n16699) );
  NAND U35078 ( .A(n57044), .B(n16699), .Z(n16700) );
  NANDN U35079 ( .A(n57045), .B(n16700), .Z(n16702) );
  NANDN U35080 ( .A(y[4760]), .B(x[4760]), .Z(n16701) );
  NANDN U35081 ( .A(y[4761]), .B(x[4761]), .Z(n42315) );
  AND U35082 ( .A(n16701), .B(n42315), .Z(n51566) );
  AND U35083 ( .A(n16702), .B(n51566), .Z(n16703) );
  XNOR U35084 ( .A(y[4762]), .B(x[4762]), .Z(n42316) );
  NANDN U35085 ( .A(x[4761]), .B(y[4761]), .Z(n24871) );
  NAND U35086 ( .A(n42316), .B(n24871), .Z(n57046) );
  OR U35087 ( .A(n16703), .B(n57046), .Z(n16705) );
  NANDN U35088 ( .A(y[4762]), .B(x[4762]), .Z(n16704) );
  NANDN U35089 ( .A(y[4763]), .B(x[4763]), .Z(n42321) );
  AND U35090 ( .A(n16704), .B(n42321), .Z(n57047) );
  AND U35091 ( .A(n16705), .B(n57047), .Z(n16706) );
  ANDN U35092 ( .B(y[4763]), .A(x[4763]), .Z(n24869) );
  XNOR U35093 ( .A(y[4764]), .B(x[4764]), .Z(n42322) );
  NANDN U35094 ( .A(n24869), .B(n42322), .Z(n51565) );
  OR U35095 ( .A(n16706), .B(n51565), .Z(n16707) );
  NAND U35096 ( .A(n51564), .B(n16707), .Z(n16708) );
  NAND U35097 ( .A(n42328), .B(n16708), .Z(n16709) );
  ANDN U35098 ( .B(n57048), .A(n16709), .Z(n16711) );
  NANDN U35099 ( .A(y[4766]), .B(x[4766]), .Z(n16710) );
  NANDN U35100 ( .A(y[4767]), .B(x[4767]), .Z(n42334) );
  NAND U35101 ( .A(n16710), .B(n42334), .Z(n51562) );
  OR U35102 ( .A(n16711), .B(n51562), .Z(n16712) );
  NAND U35103 ( .A(n51561), .B(n16712), .Z(n16713) );
  NANDN U35104 ( .A(n57051), .B(n16713), .Z(n16714) );
  AND U35105 ( .A(n24866), .B(n16714), .Z(n16715) );
  NANDN U35106 ( .A(x[4769]), .B(y[4769]), .Z(n57055) );
  AND U35107 ( .A(n16715), .B(n57055), .Z(n16717) );
  NANDN U35108 ( .A(y[4770]), .B(x[4770]), .Z(n16716) );
  NANDN U35109 ( .A(y[4771]), .B(x[4771]), .Z(n24862) );
  NAND U35110 ( .A(n16716), .B(n24862), .Z(n57056) );
  OR U35111 ( .A(n16717), .B(n57056), .Z(n16718) );
  AND U35112 ( .A(n57057), .B(n16718), .Z(n16719) );
  OR U35113 ( .A(n57058), .B(n16719), .Z(n16720) );
  NAND U35114 ( .A(n57059), .B(n16720), .Z(n16721) );
  NANDN U35115 ( .A(n57060), .B(n16721), .Z(n16722) );
  AND U35116 ( .A(n42355), .B(n16722), .Z(n16723) );
  NAND U35117 ( .A(n57062), .B(n16723), .Z(n16724) );
  NAND U35118 ( .A(n51560), .B(n16724), .Z(n16725) );
  NAND U35119 ( .A(n24858), .B(n16725), .Z(n16726) );
  ANDN U35120 ( .B(n57063), .A(n16726), .Z(n16727) );
  OR U35121 ( .A(n57065), .B(n16727), .Z(n16728) );
  NAND U35122 ( .A(n57066), .B(n16728), .Z(n16729) );
  NANDN U35123 ( .A(n57067), .B(n16729), .Z(n16730) );
  NAND U35124 ( .A(n57069), .B(n16730), .Z(n16731) );
  NAND U35125 ( .A(n51559), .B(n16731), .Z(n16732) );
  NANDN U35126 ( .A(n57070), .B(n16732), .Z(n16734) );
  NANDN U35127 ( .A(y[4784]), .B(x[4784]), .Z(n16733) );
  NANDN U35128 ( .A(y[4785]), .B(x[4785]), .Z(n42382) );
  AND U35129 ( .A(n16733), .B(n42382), .Z(n57071) );
  AND U35130 ( .A(n16734), .B(n57071), .Z(n16735) );
  XNOR U35131 ( .A(y[4786]), .B(x[4786]), .Z(n42383) );
  NANDN U35132 ( .A(x[4785]), .B(y[4785]), .Z(n24850) );
  AND U35133 ( .A(n42383), .B(n24850), .Z(n57072) );
  NANDN U35134 ( .A(n16735), .B(n57072), .Z(n16736) );
  NANDN U35135 ( .A(n57073), .B(n16736), .Z(n16737) );
  AND U35136 ( .A(n57074), .B(n16737), .Z(n16738) );
  OR U35137 ( .A(n57075), .B(n16738), .Z(n16739) );
  NAND U35138 ( .A(n57076), .B(n16739), .Z(n16740) );
  NANDN U35139 ( .A(n57077), .B(n16740), .Z(n16741) );
  NAND U35140 ( .A(n57078), .B(n16741), .Z(n16742) );
  NAND U35141 ( .A(n51558), .B(n16742), .Z(n16743) );
  NANDN U35142 ( .A(n57079), .B(n16743), .Z(n16744) );
  NANDN U35143 ( .A(y[4795]), .B(x[4795]), .Z(n51556) );
  AND U35144 ( .A(n16744), .B(n51556), .Z(n16745) );
  NANDN U35145 ( .A(y[4794]), .B(x[4794]), .Z(n57080) );
  AND U35146 ( .A(n16745), .B(n57080), .Z(n16746) );
  NANDN U35147 ( .A(x[4795]), .B(y[4795]), .Z(n24840) );
  NANDN U35148 ( .A(x[4796]), .B(y[4796]), .Z(n51557) );
  NAND U35149 ( .A(n24840), .B(n51557), .Z(n57081) );
  OR U35150 ( .A(n16746), .B(n57081), .Z(n16747) );
  AND U35151 ( .A(n57084), .B(n16747), .Z(n16748) );
  OR U35152 ( .A(n57085), .B(n16748), .Z(n16749) );
  NAND U35153 ( .A(n57086), .B(n16749), .Z(n16750) );
  NANDN U35154 ( .A(n57087), .B(n16750), .Z(n16751) );
  AND U35155 ( .A(n57088), .B(n16751), .Z(n16752) );
  OR U35156 ( .A(n57089), .B(n16752), .Z(n16753) );
  NAND U35157 ( .A(n57090), .B(n16753), .Z(n16754) );
  NANDN U35158 ( .A(n57091), .B(n16754), .Z(n16755) );
  AND U35159 ( .A(n57092), .B(n16755), .Z(n16756) );
  NANDN U35160 ( .A(y[4805]), .B(x[4805]), .Z(n24827) );
  NAND U35161 ( .A(n16756), .B(n24827), .Z(n16757) );
  ANDN U35162 ( .B(y[4806]), .A(x[4806]), .Z(n24824) );
  ANDN U35163 ( .B(n16757), .A(n24824), .Z(n16758) );
  NANDN U35164 ( .A(n24828), .B(n16758), .Z(n16759) );
  NANDN U35165 ( .A(y[4807]), .B(x[4807]), .Z(n51555) );
  AND U35166 ( .A(n16759), .B(n51555), .Z(n16760) );
  NANDN U35167 ( .A(y[4806]), .B(x[4806]), .Z(n24826) );
  AND U35168 ( .A(n16760), .B(n24826), .Z(n16761) );
  ANDN U35169 ( .B(n16762), .A(n16761), .Z(n16764) );
  NANDN U35170 ( .A(y[4808]), .B(x[4808]), .Z(n16763) );
  ANDN U35171 ( .B(x[4809]), .A(y[4809]), .Z(n42443) );
  ANDN U35172 ( .B(n16763), .A(n42443), .Z(n57097) );
  NANDN U35173 ( .A(n16764), .B(n57097), .Z(n16765) );
  NANDN U35174 ( .A(n16766), .B(n16765), .Z(n16768) );
  NANDN U35175 ( .A(y[4810]), .B(x[4810]), .Z(n16767) );
  NANDN U35176 ( .A(y[4811]), .B(x[4811]), .Z(n24821) );
  AND U35177 ( .A(n16767), .B(n24821), .Z(n57099) );
  AND U35178 ( .A(n16768), .B(n57099), .Z(n16769) );
  NANDN U35179 ( .A(x[4811]), .B(y[4811]), .Z(n42446) );
  NANDN U35180 ( .A(x[4812]), .B(y[4812]), .Z(n24820) );
  NAND U35181 ( .A(n42446), .B(n24820), .Z(n51551) );
  OR U35182 ( .A(n16769), .B(n51551), .Z(n16770) );
  NAND U35183 ( .A(n51550), .B(n16770), .Z(n16771) );
  NANDN U35184 ( .A(n57100), .B(n16771), .Z(n16772) );
  NANDN U35185 ( .A(y[4814]), .B(x[4814]), .Z(n24817) );
  NANDN U35186 ( .A(y[4815]), .B(x[4815]), .Z(n42459) );
  AND U35187 ( .A(n24817), .B(n42459), .Z(n57101) );
  AND U35188 ( .A(n16772), .B(n57101), .Z(n16774) );
  NANDN U35189 ( .A(x[4815]), .B(y[4815]), .Z(n24815) );
  XNOR U35190 ( .A(x[4816]), .B(y[4816]), .Z(n16773) );
  AND U35191 ( .A(n24815), .B(n16773), .Z(n57102) );
  NANDN U35192 ( .A(n16774), .B(n57102), .Z(n16775) );
  NANDN U35193 ( .A(n57103), .B(n16775), .Z(n16776) );
  AND U35194 ( .A(n57104), .B(n16776), .Z(n16777) );
  OR U35195 ( .A(n57105), .B(n16777), .Z(n16778) );
  NAND U35196 ( .A(n57106), .B(n16778), .Z(n16779) );
  NANDN U35197 ( .A(n57107), .B(n16779), .Z(n16780) );
  AND U35198 ( .A(n24807), .B(n16780), .Z(n16781) );
  NANDN U35199 ( .A(x[4821]), .B(y[4821]), .Z(n51548) );
  NAND U35200 ( .A(n16781), .B(n51548), .Z(n16782) );
  NANDN U35201 ( .A(n57108), .B(n16782), .Z(n16783) );
  NANDN U35202 ( .A(x[4823]), .B(y[4823]), .Z(n42476) );
  NANDN U35203 ( .A(x[4824]), .B(y[4824]), .Z(n24803) );
  AND U35204 ( .A(n42476), .B(n24803), .Z(n57111) );
  AND U35205 ( .A(n16783), .B(n57111), .Z(n16784) );
  NANDN U35206 ( .A(y[4824]), .B(x[4824]), .Z(n24804) );
  NANDN U35207 ( .A(y[4825]), .B(x[4825]), .Z(n24800) );
  AND U35208 ( .A(n24804), .B(n24800), .Z(n57112) );
  NANDN U35209 ( .A(n16784), .B(n57112), .Z(n16785) );
  NAND U35210 ( .A(n57113), .B(n16785), .Z(n16786) );
  NANDN U35211 ( .A(n57114), .B(n16786), .Z(n16787) );
  AND U35212 ( .A(n24798), .B(n16787), .Z(n16788) );
  NANDN U35213 ( .A(x[4827]), .B(y[4827]), .Z(n51546) );
  AND U35214 ( .A(n16788), .B(n51546), .Z(n16790) );
  NANDN U35215 ( .A(y[4828]), .B(x[4828]), .Z(n16789) );
  NANDN U35216 ( .A(y[4829]), .B(x[4829]), .Z(n24795) );
  NAND U35217 ( .A(n16789), .B(n24795), .Z(n57115) );
  OR U35218 ( .A(n16790), .B(n57115), .Z(n16791) );
  AND U35219 ( .A(n57116), .B(n16791), .Z(n16792) );
  OR U35220 ( .A(n57117), .B(n16792), .Z(n16793) );
  NAND U35221 ( .A(n57118), .B(n16793), .Z(n16794) );
  NANDN U35222 ( .A(n57119), .B(n16794), .Z(n16795) );
  AND U35223 ( .A(n57120), .B(n16795), .Z(n16797) );
  NANDN U35224 ( .A(y[4834]), .B(x[4834]), .Z(n16796) );
  NANDN U35225 ( .A(y[4835]), .B(x[4835]), .Z(n24786) );
  NAND U35226 ( .A(n16796), .B(n24786), .Z(n57121) );
  OR U35227 ( .A(n16797), .B(n57121), .Z(n16798) );
  AND U35228 ( .A(n16799), .B(n16798), .Z(n16800) );
  OR U35229 ( .A(n57124), .B(n16800), .Z(n16801) );
  NAND U35230 ( .A(n57126), .B(n16801), .Z(n16802) );
  NANDN U35231 ( .A(n51545), .B(n16802), .Z(n16803) );
  XOR U35232 ( .A(x[4840]), .B(y[4840]), .Z(n42516) );
  ANDN U35233 ( .B(n16803), .A(n42516), .Z(n16804) );
  NANDN U35234 ( .A(x[4839]), .B(y[4839]), .Z(n51544) );
  AND U35235 ( .A(n16804), .B(n51544), .Z(n16806) );
  NANDN U35236 ( .A(y[4840]), .B(x[4840]), .Z(n16805) );
  NANDN U35237 ( .A(y[4841]), .B(x[4841]), .Z(n24781) );
  NAND U35238 ( .A(n16805), .B(n24781), .Z(n57128) );
  OR U35239 ( .A(n16806), .B(n57128), .Z(n16807) );
  AND U35240 ( .A(n24782), .B(n16807), .Z(n16808) );
  NANDN U35241 ( .A(x[4841]), .B(y[4841]), .Z(n57130) );
  AND U35242 ( .A(n16808), .B(n57130), .Z(n16809) );
  OR U35243 ( .A(n57131), .B(n16809), .Z(n16810) );
  NAND U35244 ( .A(n16811), .B(n16810), .Z(n16813) );
  NANDN U35245 ( .A(y[4844]), .B(x[4844]), .Z(n16812) );
  NANDN U35246 ( .A(y[4845]), .B(x[4845]), .Z(n24777) );
  AND U35247 ( .A(n16812), .B(n24777), .Z(n57134) );
  AND U35248 ( .A(n16813), .B(n57134), .Z(n16814) );
  NOR U35249 ( .A(n42526), .B(n16814), .Z(n16815) );
  NAND U35250 ( .A(n24778), .B(n16815), .Z(n16816) );
  NANDN U35251 ( .A(n57137), .B(n16816), .Z(n16817) );
  AND U35252 ( .A(n57138), .B(n16817), .Z(n16818) );
  NANDN U35253 ( .A(y[4848]), .B(x[4848]), .Z(n24775) );
  NANDN U35254 ( .A(y[4849]), .B(x[4849]), .Z(n24772) );
  NAND U35255 ( .A(n24775), .B(n24772), .Z(n57139) );
  OR U35256 ( .A(n16818), .B(n57139), .Z(n16819) );
  AND U35257 ( .A(n16820), .B(n16819), .Z(n16821) );
  OR U35258 ( .A(n57145), .B(n16821), .Z(n16822) );
  NAND U35259 ( .A(n57146), .B(n16822), .Z(n16823) );
  NANDN U35260 ( .A(n57147), .B(n16823), .Z(n16824) );
  AND U35261 ( .A(n24768), .B(n16824), .Z(n16825) );
  NANDN U35262 ( .A(x[4853]), .B(y[4853]), .Z(n51542) );
  AND U35263 ( .A(n16825), .B(n51542), .Z(n16827) );
  NANDN U35264 ( .A(y[4854]), .B(x[4854]), .Z(n16826) );
  NANDN U35265 ( .A(y[4855]), .B(x[4855]), .Z(n24765) );
  NAND U35266 ( .A(n16826), .B(n24765), .Z(n57148) );
  OR U35267 ( .A(n16827), .B(n57148), .Z(n16828) );
  AND U35268 ( .A(n24766), .B(n16828), .Z(n16829) );
  NANDN U35269 ( .A(x[4855]), .B(y[4855]), .Z(n57149) );
  AND U35270 ( .A(n16829), .B(n57149), .Z(n16830) );
  OR U35271 ( .A(n57151), .B(n16830), .Z(n16831) );
  NAND U35272 ( .A(n16832), .B(n16831), .Z(n16834) );
  NANDN U35273 ( .A(y[4858]), .B(x[4858]), .Z(n16833) );
  NANDN U35274 ( .A(y[4859]), .B(x[4859]), .Z(n24761) );
  AND U35275 ( .A(n16833), .B(n24761), .Z(n57154) );
  AND U35276 ( .A(n16834), .B(n57154), .Z(n16835) );
  NOR U35277 ( .A(n42557), .B(n16835), .Z(n16836) );
  NAND U35278 ( .A(n24762), .B(n16836), .Z(n16837) );
  NANDN U35279 ( .A(n57158), .B(n16837), .Z(n16838) );
  AND U35280 ( .A(n24760), .B(n16838), .Z(n16839) );
  NANDN U35281 ( .A(x[4861]), .B(y[4861]), .Z(n51540) );
  NAND U35282 ( .A(n16839), .B(n51540), .Z(n16840) );
  NANDN U35283 ( .A(n57159), .B(n16840), .Z(n16841) );
  AND U35284 ( .A(n24758), .B(n16841), .Z(n16842) );
  NANDN U35285 ( .A(x[4863]), .B(y[4863]), .Z(n57160) );
  AND U35286 ( .A(n16842), .B(n57160), .Z(n16844) );
  NANDN U35287 ( .A(y[4864]), .B(x[4864]), .Z(n16843) );
  NANDN U35288 ( .A(y[4865]), .B(x[4865]), .Z(n24755) );
  AND U35289 ( .A(n16843), .B(n24755), .Z(n51539) );
  NANDN U35290 ( .A(n16844), .B(n51539), .Z(n16845) );
  NAND U35291 ( .A(n16846), .B(n16845), .Z(n16847) );
  AND U35292 ( .A(n57164), .B(n16847), .Z(n16848) );
  NOR U35293 ( .A(n24754), .B(n16848), .Z(n16849) );
  NAND U35294 ( .A(n42579), .B(n16849), .Z(n16850) );
  NANDN U35295 ( .A(n57167), .B(n16850), .Z(n16851) );
  AND U35296 ( .A(n24753), .B(n16851), .Z(n16852) );
  NANDN U35297 ( .A(x[4869]), .B(y[4869]), .Z(n51537) );
  AND U35298 ( .A(n16852), .B(n51537), .Z(n16854) );
  NANDN U35299 ( .A(y[4870]), .B(x[4870]), .Z(n16853) );
  NANDN U35300 ( .A(y[4871]), .B(x[4871]), .Z(n24750) );
  NAND U35301 ( .A(n16853), .B(n24750), .Z(n57168) );
  OR U35302 ( .A(n16854), .B(n57168), .Z(n16855) );
  AND U35303 ( .A(n24751), .B(n16855), .Z(n16856) );
  NANDN U35304 ( .A(x[4871]), .B(y[4871]), .Z(n57171) );
  AND U35305 ( .A(n16856), .B(n57171), .Z(n16857) );
  OR U35306 ( .A(n57174), .B(n16857), .Z(n16858) );
  NAND U35307 ( .A(n16859), .B(n16858), .Z(n16861) );
  NANDN U35308 ( .A(y[4874]), .B(x[4874]), .Z(n16860) );
  NANDN U35309 ( .A(y[4875]), .B(x[4875]), .Z(n24745) );
  AND U35310 ( .A(n16860), .B(n24745), .Z(n57177) );
  AND U35311 ( .A(n16861), .B(n57177), .Z(n16863) );
  XNOR U35312 ( .A(x[4876]), .B(y[4876]), .Z(n24746) );
  ANDN U35313 ( .B(y[4875]), .A(x[4875]), .Z(n24747) );
  ANDN U35314 ( .B(n24746), .A(n24747), .Z(n16862) );
  NANDN U35315 ( .A(n16863), .B(n16862), .Z(n16865) );
  NANDN U35316 ( .A(y[4876]), .B(x[4876]), .Z(n16864) );
  NANDN U35317 ( .A(y[4877]), .B(x[4877]), .Z(n24743) );
  AND U35318 ( .A(n16864), .B(n24743), .Z(n57180) );
  AND U35319 ( .A(n16865), .B(n57180), .Z(n16866) );
  XNOR U35320 ( .A(y[4878]), .B(x[4878]), .Z(n24744) );
  NANDN U35321 ( .A(x[4877]), .B(y[4877]), .Z(n42597) );
  NAND U35322 ( .A(n24744), .B(n42597), .Z(n57181) );
  OR U35323 ( .A(n16866), .B(n57181), .Z(n16867) );
  NAND U35324 ( .A(n57182), .B(n16867), .Z(n16868) );
  NANDN U35325 ( .A(n51536), .B(n16868), .Z(n16869) );
  NAND U35326 ( .A(n51535), .B(n16869), .Z(n16870) );
  AND U35327 ( .A(n57184), .B(n16870), .Z(n16872) );
  NANDN U35328 ( .A(y[4882]), .B(x[4882]), .Z(n16871) );
  NANDN U35329 ( .A(y[4883]), .B(x[4883]), .Z(n24734) );
  AND U35330 ( .A(n16871), .B(n24734), .Z(n57185) );
  NANDN U35331 ( .A(n16872), .B(n57185), .Z(n16873) );
  AND U35332 ( .A(n57187), .B(n16873), .Z(n16874) );
  NANDN U35333 ( .A(y[4884]), .B(x[4884]), .Z(n24733) );
  NANDN U35334 ( .A(y[4885]), .B(x[4885]), .Z(n24730) );
  NAND U35335 ( .A(n24733), .B(n24730), .Z(n57188) );
  OR U35336 ( .A(n16874), .B(n57188), .Z(n16875) );
  AND U35337 ( .A(n24731), .B(n16875), .Z(n16876) );
  NANDN U35338 ( .A(x[4885]), .B(y[4885]), .Z(n57189) );
  AND U35339 ( .A(n16876), .B(n57189), .Z(n16878) );
  NANDN U35340 ( .A(y[4886]), .B(x[4886]), .Z(n16877) );
  NANDN U35341 ( .A(y[4887]), .B(x[4887]), .Z(n24729) );
  NAND U35342 ( .A(n16877), .B(n24729), .Z(n57191) );
  OR U35343 ( .A(n16878), .B(n57191), .Z(n16879) );
  AND U35344 ( .A(n57192), .B(n16879), .Z(n16880) );
  OR U35345 ( .A(n57193), .B(n16880), .Z(n16881) );
  NAND U35346 ( .A(n57194), .B(n16881), .Z(n16882) );
  NANDN U35347 ( .A(n57195), .B(n16882), .Z(n16883) );
  AND U35348 ( .A(n57196), .B(n16883), .Z(n16884) );
  NANDN U35349 ( .A(y[4893]), .B(x[4893]), .Z(n24719) );
  ANDN U35350 ( .B(x[4892]), .A(y[4892]), .Z(n42632) );
  ANDN U35351 ( .B(n24719), .A(n42632), .Z(n57197) );
  NANDN U35352 ( .A(n16884), .B(n57197), .Z(n16885) );
  NANDN U35353 ( .A(n57198), .B(n16885), .Z(n16886) );
  NANDN U35354 ( .A(y[4894]), .B(x[4894]), .Z(n24718) );
  NANDN U35355 ( .A(y[4895]), .B(x[4895]), .Z(n42643) );
  AND U35356 ( .A(n24718), .B(n42643), .Z(n57199) );
  AND U35357 ( .A(n16886), .B(n57199), .Z(n16887) );
  NANDN U35358 ( .A(x[4895]), .B(y[4895]), .Z(n24716) );
  NANDN U35359 ( .A(x[4896]), .B(y[4896]), .Z(n24715) );
  AND U35360 ( .A(n24716), .B(n24715), .Z(n57200) );
  NANDN U35361 ( .A(n16887), .B(n57200), .Z(n16888) );
  NAND U35362 ( .A(n57201), .B(n16888), .Z(n16889) );
  NANDN U35363 ( .A(n57202), .B(n16889), .Z(n16890) );
  AND U35364 ( .A(n57204), .B(n16890), .Z(n16891) );
  NANDN U35365 ( .A(x[4899]), .B(y[4899]), .Z(n24710) );
  NANDN U35366 ( .A(x[4900]), .B(y[4900]), .Z(n24709) );
  NAND U35367 ( .A(n24710), .B(n24709), .Z(n57205) );
  OR U35368 ( .A(n16891), .B(n57205), .Z(n16892) );
  AND U35369 ( .A(n57206), .B(n16892), .Z(n16893) );
  OR U35370 ( .A(n57207), .B(n16893), .Z(n16894) );
  NAND U35371 ( .A(n57208), .B(n16894), .Z(n16895) );
  NANDN U35372 ( .A(n57209), .B(n16895), .Z(n16896) );
  NAND U35373 ( .A(n57210), .B(n16896), .Z(n16897) );
  AND U35374 ( .A(n24701), .B(n16897), .Z(n16898) );
  NANDN U35375 ( .A(n24702), .B(n16898), .Z(n16900) );
  NANDN U35376 ( .A(y[4906]), .B(x[4906]), .Z(n16899) );
  NANDN U35377 ( .A(y[4907]), .B(x[4907]), .Z(n24698) );
  AND U35378 ( .A(n16899), .B(n24698), .Z(n57211) );
  AND U35379 ( .A(n16900), .B(n57211), .Z(n16901) );
  NANDN U35380 ( .A(x[4907]), .B(y[4907]), .Z(n24699) );
  NANDN U35381 ( .A(x[4908]), .B(y[4908]), .Z(n24696) );
  NAND U35382 ( .A(n24699), .B(n24696), .Z(n51532) );
  OR U35383 ( .A(n16901), .B(n51532), .Z(n16902) );
  NAND U35384 ( .A(n51531), .B(n16902), .Z(n16903) );
  NANDN U35385 ( .A(n57212), .B(n16903), .Z(n16904) );
  NANDN U35386 ( .A(y[4910]), .B(x[4910]), .Z(n24693) );
  NANDN U35387 ( .A(y[4911]), .B(x[4911]), .Z(n42681) );
  AND U35388 ( .A(n24693), .B(n42681), .Z(n57213) );
  AND U35389 ( .A(n16904), .B(n57213), .Z(n16905) );
  NANDN U35390 ( .A(x[4911]), .B(y[4911]), .Z(n24691) );
  NANDN U35391 ( .A(x[4912]), .B(y[4912]), .Z(n24690) );
  AND U35392 ( .A(n24691), .B(n24690), .Z(n57215) );
  NANDN U35393 ( .A(n16905), .B(n57215), .Z(n16906) );
  NANDN U35394 ( .A(n57216), .B(n16906), .Z(n16907) );
  AND U35395 ( .A(n24689), .B(n16907), .Z(n16908) );
  NANDN U35396 ( .A(x[4913]), .B(y[4913]), .Z(n57218) );
  AND U35397 ( .A(n16908), .B(n57218), .Z(n16909) );
  OR U35398 ( .A(n57219), .B(n16909), .Z(n16910) );
  NAND U35399 ( .A(n16911), .B(n16910), .Z(n16913) );
  NANDN U35400 ( .A(y[4916]), .B(x[4916]), .Z(n16912) );
  NANDN U35401 ( .A(y[4917]), .B(x[4917]), .Z(n24684) );
  AND U35402 ( .A(n16912), .B(n24684), .Z(n57222) );
  AND U35403 ( .A(n16913), .B(n57222), .Z(n16914) );
  ANDN U35404 ( .B(n16915), .A(n16914), .Z(n16917) );
  NANDN U35405 ( .A(y[4918]), .B(x[4918]), .Z(n16916) );
  NANDN U35406 ( .A(y[4919]), .B(x[4919]), .Z(n24683) );
  NAND U35407 ( .A(n16916), .B(n24683), .Z(n51529) );
  OR U35408 ( .A(n16917), .B(n51529), .Z(n16918) );
  NAND U35409 ( .A(n51528), .B(n16918), .Z(n16919) );
  NANDN U35410 ( .A(n57224), .B(n16919), .Z(n16920) );
  NANDN U35411 ( .A(x[4921]), .B(y[4921]), .Z(n24680) );
  NANDN U35412 ( .A(x[4922]), .B(y[4922]), .Z(n24677) );
  AND U35413 ( .A(n24680), .B(n24677), .Z(n57225) );
  AND U35414 ( .A(n16920), .B(n57225), .Z(n16921) );
  ANDN U35415 ( .B(x[4923]), .A(y[4923]), .Z(n42707) );
  NANDN U35416 ( .A(y[4922]), .B(x[4922]), .Z(n24678) );
  NANDN U35417 ( .A(n42707), .B(n24678), .Z(n51527) );
  OR U35418 ( .A(n16921), .B(n51527), .Z(n16922) );
  NAND U35419 ( .A(n16923), .B(n16922), .Z(n16925) );
  NANDN U35420 ( .A(y[4924]), .B(x[4924]), .Z(n16924) );
  NANDN U35421 ( .A(y[4925]), .B(x[4925]), .Z(n24675) );
  AND U35422 ( .A(n16924), .B(n24675), .Z(n57230) );
  AND U35423 ( .A(n16925), .B(n57230), .Z(n16926) );
  NOR U35424 ( .A(n42710), .B(n16926), .Z(n16927) );
  NAND U35425 ( .A(n24676), .B(n16927), .Z(n16928) );
  NANDN U35426 ( .A(n57231), .B(n16928), .Z(n16929) );
  AND U35427 ( .A(n24674), .B(n16929), .Z(n16930) );
  NANDN U35428 ( .A(x[4927]), .B(y[4927]), .Z(n57232) );
  AND U35429 ( .A(n16930), .B(n57232), .Z(n16931) );
  OR U35430 ( .A(n57234), .B(n16931), .Z(n16932) );
  AND U35431 ( .A(n24672), .B(n16932), .Z(n16933) );
  NANDN U35432 ( .A(x[4929]), .B(y[4929]), .Z(n57235) );
  AND U35433 ( .A(n16933), .B(n57235), .Z(n16935) );
  NANDN U35434 ( .A(y[4930]), .B(x[4930]), .Z(n16934) );
  NANDN U35435 ( .A(y[4931]), .B(x[4931]), .Z(n24669) );
  NAND U35436 ( .A(n16934), .B(n24669), .Z(n51524) );
  OR U35437 ( .A(n16935), .B(n51524), .Z(n16936) );
  AND U35438 ( .A(n57238), .B(n16936), .Z(n16937) );
  NANDN U35439 ( .A(y[4932]), .B(x[4932]), .Z(n24670) );
  NANDN U35440 ( .A(y[4933]), .B(x[4933]), .Z(n24666) );
  NAND U35441 ( .A(n24670), .B(n24666), .Z(n57239) );
  OR U35442 ( .A(n16937), .B(n57239), .Z(n16938) );
  NAND U35443 ( .A(n16939), .B(n16938), .Z(n16940) );
  NANDN U35444 ( .A(n57242), .B(n16940), .Z(n16941) );
  AND U35445 ( .A(n24664), .B(n16941), .Z(n16942) );
  NANDN U35446 ( .A(n24665), .B(n16942), .Z(n16943) );
  NAND U35447 ( .A(n57244), .B(n16943), .Z(n16944) );
  NANDN U35448 ( .A(n57245), .B(n16944), .Z(n16945) );
  AND U35449 ( .A(n57246), .B(n16945), .Z(n16946) );
  ANDN U35450 ( .B(n57248), .A(n16946), .Z(n16947) );
  NANDN U35451 ( .A(n42745), .B(n16947), .Z(n16948) );
  NANDN U35452 ( .A(n57249), .B(n16948), .Z(n16949) );
  AND U35453 ( .A(n24659), .B(n16949), .Z(n16950) );
  NANDN U35454 ( .A(x[4941]), .B(y[4941]), .Z(n57250) );
  AND U35455 ( .A(n16950), .B(n57250), .Z(n16952) );
  NANDN U35456 ( .A(y[4942]), .B(x[4942]), .Z(n16951) );
  NANDN U35457 ( .A(y[4943]), .B(x[4943]), .Z(n42753) );
  NAND U35458 ( .A(n16951), .B(n42753), .Z(n57252) );
  OR U35459 ( .A(n16952), .B(n57252), .Z(n16953) );
  AND U35460 ( .A(n57254), .B(n16953), .Z(n16954) );
  NAND U35461 ( .A(n42754), .B(n16954), .Z(n16955) );
  NAND U35462 ( .A(n57256), .B(n16955), .Z(n16956) );
  NANDN U35463 ( .A(n16957), .B(n16956), .Z(n16958) );
  AND U35464 ( .A(n57257), .B(n16958), .Z(n16959) );
  ANDN U35465 ( .B(n57259), .A(n16959), .Z(n16960) );
  NAND U35466 ( .A(n42764), .B(n16960), .Z(n16961) );
  NANDN U35467 ( .A(y[4954]), .B(x[4954]), .Z(n16962) );
  NANDN U35468 ( .A(y[4955]), .B(x[4955]), .Z(n42782) );
  AND U35469 ( .A(n16962), .B(n42782), .Z(n51519) );
  ANDN U35470 ( .B(y[4957]), .A(x[4957]), .Z(n57272) );
  NANDN U35471 ( .A(x[4959]), .B(y[4959]), .Z(n51517) );
  NANDN U35472 ( .A(y[4960]), .B(x[4960]), .Z(n16963) );
  NANDN U35473 ( .A(y[4961]), .B(x[4961]), .Z(n24642) );
  AND U35474 ( .A(n16963), .B(n24642), .Z(n57275) );
  NAND U35475 ( .A(n16965), .B(n16964), .Z(n16966) );
  AND U35476 ( .A(n57276), .B(n16966), .Z(n16967) );
  NOR U35477 ( .A(n42798), .B(n16967), .Z(n16968) );
  NAND U35478 ( .A(n42802), .B(n16968), .Z(n16969) );
  NANDN U35479 ( .A(n57279), .B(n16969), .Z(n16970) );
  AND U35480 ( .A(n24641), .B(n16970), .Z(n16971) );
  NANDN U35481 ( .A(n57280), .B(n16971), .Z(n16972) );
  NAND U35482 ( .A(n57284), .B(n16972), .Z(n16973) );
  NAND U35483 ( .A(n57285), .B(n16973), .Z(n16974) );
  AND U35484 ( .A(n57286), .B(n16974), .Z(n16976) );
  XNOR U35485 ( .A(x[4970]), .B(y[4970]), .Z(n24636) );
  NANDN U35486 ( .A(x[4969]), .B(y[4969]), .Z(n57288) );
  AND U35487 ( .A(n24636), .B(n57288), .Z(n16975) );
  NANDN U35488 ( .A(n16976), .B(n16975), .Z(n16977) );
  AND U35489 ( .A(n57289), .B(n16977), .Z(n16978) );
  OR U35490 ( .A(n57290), .B(n16978), .Z(n16979) );
  NAND U35491 ( .A(n57291), .B(n16979), .Z(n16980) );
  NANDN U35492 ( .A(n57292), .B(n16980), .Z(n16981) );
  AND U35493 ( .A(n57293), .B(n16981), .Z(n16982) );
  NANDN U35494 ( .A(x[4975]), .B(y[4975]), .Z(n24626) );
  NANDN U35495 ( .A(x[4976]), .B(y[4976]), .Z(n24623) );
  NAND U35496 ( .A(n24626), .B(n24623), .Z(n51514) );
  OR U35497 ( .A(n16982), .B(n51514), .Z(n16983) );
  NANDN U35498 ( .A(y[4976]), .B(x[4976]), .Z(n24624) );
  NANDN U35499 ( .A(y[4977]), .B(x[4977]), .Z(n24620) );
  AND U35500 ( .A(n24624), .B(n24620), .Z(n51513) );
  AND U35501 ( .A(n16983), .B(n51513), .Z(n16984) );
  XNOR U35502 ( .A(y[4978]), .B(x[4978]), .Z(n24621) );
  NANDN U35503 ( .A(x[4977]), .B(y[4977]), .Z(n24622) );
  NAND U35504 ( .A(n24621), .B(n24622), .Z(n57294) );
  OR U35505 ( .A(n16984), .B(n57294), .Z(n16985) );
  NAND U35506 ( .A(n57295), .B(n16985), .Z(n16986) );
  NANDN U35507 ( .A(n16987), .B(n16986), .Z(n16988) );
  AND U35508 ( .A(n57298), .B(n16988), .Z(n16989) );
  NOR U35509 ( .A(n57299), .B(n16989), .Z(n16990) );
  NAND U35510 ( .A(n24619), .B(n16990), .Z(n16991) );
  NANDN U35511 ( .A(n57302), .B(n16991), .Z(n16992) );
  AND U35512 ( .A(n42848), .B(n16992), .Z(n16993) );
  NANDN U35513 ( .A(x[4983]), .B(y[4983]), .Z(n57303) );
  AND U35514 ( .A(n16993), .B(n57303), .Z(n16995) );
  NANDN U35515 ( .A(y[4984]), .B(x[4984]), .Z(n16994) );
  NANDN U35516 ( .A(y[4985]), .B(x[4985]), .Z(n24616) );
  NAND U35517 ( .A(n16994), .B(n24616), .Z(n57305) );
  OR U35518 ( .A(n16995), .B(n57305), .Z(n16996) );
  AND U35519 ( .A(n24617), .B(n16996), .Z(n16997) );
  ANDN U35520 ( .B(y[4985]), .A(x[4985]), .Z(n57306) );
  ANDN U35521 ( .B(n16997), .A(n57306), .Z(n16999) );
  NANDN U35522 ( .A(y[4986]), .B(x[4986]), .Z(n16998) );
  NANDN U35523 ( .A(y[4987]), .B(x[4987]), .Z(n42857) );
  AND U35524 ( .A(n16998), .B(n42857), .Z(n57308) );
  NANDN U35525 ( .A(n16999), .B(n57308), .Z(n17000) );
  NAND U35526 ( .A(n17001), .B(n17000), .Z(n17003) );
  NANDN U35527 ( .A(y[4988]), .B(x[4988]), .Z(n17002) );
  NANDN U35528 ( .A(y[4989]), .B(x[4989]), .Z(n24614) );
  AND U35529 ( .A(n17002), .B(n24614), .Z(n51510) );
  AND U35530 ( .A(n17003), .B(n51510), .Z(n17004) );
  NOR U35531 ( .A(n57311), .B(n17004), .Z(n17005) );
  NAND U35532 ( .A(n24615), .B(n17005), .Z(n17006) );
  NANDN U35533 ( .A(n57313), .B(n17006), .Z(n17007) );
  AND U35534 ( .A(n42869), .B(n17007), .Z(n17008) );
  NANDN U35535 ( .A(n42865), .B(n17008), .Z(n17009) );
  NAND U35536 ( .A(n57317), .B(n17009), .Z(n17010) );
  NANDN U35537 ( .A(n57318), .B(n17010), .Z(n17011) );
  AND U35538 ( .A(n57319), .B(n17011), .Z(n17012) );
  NOR U35539 ( .A(n42876), .B(n17012), .Z(n17013) );
  NAND U35540 ( .A(n42881), .B(n17013), .Z(n17014) );
  NANDN U35541 ( .A(n57322), .B(n17014), .Z(n17015) );
  AND U35542 ( .A(n24610), .B(n17015), .Z(n17016) );
  NANDN U35543 ( .A(x[4997]), .B(y[4997]), .Z(n57323) );
  AND U35544 ( .A(n17016), .B(n57323), .Z(n17018) );
  NANDN U35545 ( .A(y[4998]), .B(x[4998]), .Z(n17017) );
  NANDN U35546 ( .A(y[4999]), .B(x[4999]), .Z(n24608) );
  AND U35547 ( .A(n17017), .B(n24608), .Z(n57325) );
  NANDN U35548 ( .A(n17018), .B(n57325), .Z(n17019) );
  AND U35549 ( .A(n57326), .B(n17019), .Z(n17020) );
  NANDN U35550 ( .A(y[5000]), .B(x[5000]), .Z(n24607) );
  NANDN U35551 ( .A(y[5001]), .B(x[5001]), .Z(n24604) );
  AND U35552 ( .A(n24607), .B(n24604), .Z(n57327) );
  NANDN U35553 ( .A(n17020), .B(n57327), .Z(n17021) );
  NAND U35554 ( .A(n17022), .B(n17021), .Z(n17024) );
  NANDN U35555 ( .A(y[5002]), .B(x[5002]), .Z(n17023) );
  NANDN U35556 ( .A(y[5003]), .B(x[5003]), .Z(n42900) );
  AND U35557 ( .A(n17023), .B(n42900), .Z(n51509) );
  AND U35558 ( .A(n17024), .B(n51509), .Z(n17025) );
  NOR U35559 ( .A(n42897), .B(n17025), .Z(n17026) );
  NAND U35560 ( .A(n42901), .B(n17026), .Z(n17027) );
  NANDN U35561 ( .A(n51508), .B(n17027), .Z(n17028) );
  AND U35562 ( .A(n57333), .B(n17028), .Z(n17029) );
  NANDN U35563 ( .A(y[5006]), .B(x[5006]), .Z(n24601) );
  NANDN U35564 ( .A(y[5007]), .B(x[5007]), .Z(n42910) );
  AND U35565 ( .A(n24601), .B(n42910), .Z(n57334) );
  NANDN U35566 ( .A(n17029), .B(n57334), .Z(n17030) );
  NAND U35567 ( .A(n17031), .B(n17030), .Z(n17033) );
  NANDN U35568 ( .A(y[5008]), .B(x[5008]), .Z(n17032) );
  NANDN U35569 ( .A(y[5009]), .B(x[5009]), .Z(n24598) );
  AND U35570 ( .A(n17032), .B(n24598), .Z(n51507) );
  AND U35571 ( .A(n17033), .B(n51507), .Z(n17035) );
  XNOR U35572 ( .A(x[5010]), .B(y[5010]), .Z(n24599) );
  ANDN U35573 ( .B(y[5009]), .A(x[5009]), .Z(n57337) );
  ANDN U35574 ( .B(n24599), .A(n57337), .Z(n17034) );
  NANDN U35575 ( .A(n17035), .B(n17034), .Z(n17037) );
  NANDN U35576 ( .A(y[5010]), .B(x[5010]), .Z(n17036) );
  NANDN U35577 ( .A(y[5011]), .B(x[5011]), .Z(n24595) );
  AND U35578 ( .A(n17036), .B(n24595), .Z(n57339) );
  AND U35579 ( .A(n17037), .B(n57339), .Z(n17038) );
  NOR U35580 ( .A(n24597), .B(n17038), .Z(n17039) );
  NAND U35581 ( .A(n24596), .B(n17039), .Z(n17040) );
  NANDN U35582 ( .A(n57342), .B(n17040), .Z(n17041) );
  AND U35583 ( .A(n57343), .B(n17041), .Z(n17042) );
  NANDN U35584 ( .A(y[5014]), .B(x[5014]), .Z(n24592) );
  NANDN U35585 ( .A(y[5015]), .B(x[5015]), .Z(n42928) );
  AND U35586 ( .A(n24592), .B(n42928), .Z(n57344) );
  NANDN U35587 ( .A(n17042), .B(n57344), .Z(n17043) );
  NAND U35588 ( .A(n17044), .B(n17043), .Z(n17046) );
  NANDN U35589 ( .A(y[5016]), .B(x[5016]), .Z(n17045) );
  NANDN U35590 ( .A(y[5017]), .B(x[5017]), .Z(n24589) );
  AND U35591 ( .A(n17045), .B(n24589), .Z(n51506) );
  AND U35592 ( .A(n17046), .B(n51506), .Z(n17047) );
  NOR U35593 ( .A(n57349), .B(n17047), .Z(n17048) );
  NAND U35594 ( .A(n24590), .B(n17048), .Z(n17049) );
  NANDN U35595 ( .A(n51505), .B(n17049), .Z(n17050) );
  NANDN U35596 ( .A(x[5019]), .B(y[5019]), .Z(n42936) );
  NANDN U35597 ( .A(x[5020]), .B(y[5020]), .Z(n24586) );
  AND U35598 ( .A(n42936), .B(n24586), .Z(n51504) );
  AND U35599 ( .A(n17050), .B(n51504), .Z(n17051) );
  NANDN U35600 ( .A(y[5020]), .B(x[5020]), .Z(n24587) );
  NANDN U35601 ( .A(y[5021]), .B(x[5021]), .Z(n24584) );
  NAND U35602 ( .A(n24587), .B(n24584), .Z(n57352) );
  OR U35603 ( .A(n17051), .B(n57352), .Z(n17052) );
  AND U35604 ( .A(n24585), .B(n17052), .Z(n17053) );
  NANDN U35605 ( .A(x[5021]), .B(y[5021]), .Z(n57354) );
  AND U35606 ( .A(n17053), .B(n57354), .Z(n17055) );
  NANDN U35607 ( .A(y[5022]), .B(x[5022]), .Z(n17054) );
  NANDN U35608 ( .A(y[5023]), .B(x[5023]), .Z(n24582) );
  NAND U35609 ( .A(n17054), .B(n24582), .Z(n57355) );
  OR U35610 ( .A(n17055), .B(n57355), .Z(n17056) );
  AND U35611 ( .A(n17057), .B(n17056), .Z(n17059) );
  NANDN U35612 ( .A(y[5024]), .B(x[5024]), .Z(n17058) );
  NANDN U35613 ( .A(y[5025]), .B(x[5025]), .Z(n24580) );
  NAND U35614 ( .A(n17058), .B(n24580), .Z(n51503) );
  OR U35615 ( .A(n17059), .B(n51503), .Z(n17060) );
  NAND U35616 ( .A(n57358), .B(n17060), .Z(n17061) );
  NANDN U35617 ( .A(n57359), .B(n17061), .Z(n17062) );
  AND U35618 ( .A(n42958), .B(n17062), .Z(n17063) );
  NANDN U35619 ( .A(x[5027]), .B(y[5027]), .Z(n57360) );
  AND U35620 ( .A(n17063), .B(n57360), .Z(n17064) );
  OR U35621 ( .A(n57364), .B(n17064), .Z(n17065) );
  AND U35622 ( .A(n17066), .B(n17065), .Z(n17067) );
  OR U35623 ( .A(n57367), .B(n17067), .Z(n17068) );
  NAND U35624 ( .A(n57368), .B(n17068), .Z(n17069) );
  NANDN U35625 ( .A(n57369), .B(n17069), .Z(n17070) );
  AND U35626 ( .A(n57370), .B(n17070), .Z(n17071) );
  NANDN U35627 ( .A(y[5034]), .B(x[5034]), .Z(n24571) );
  NANDN U35628 ( .A(y[5035]), .B(x[5035]), .Z(n24568) );
  NAND U35629 ( .A(n24571), .B(n24568), .Z(n57371) );
  OR U35630 ( .A(n17071), .B(n57371), .Z(n17072) );
  AND U35631 ( .A(n57372), .B(n17072), .Z(n17073) );
  OR U35632 ( .A(n57373), .B(n17073), .Z(n17074) );
  NAND U35633 ( .A(n17075), .B(n17074), .Z(n17076) );
  NANDN U35634 ( .A(n57374), .B(n17076), .Z(n17077) );
  AND U35635 ( .A(n57375), .B(n17077), .Z(n17078) );
  OR U35636 ( .A(n57376), .B(n17078), .Z(n17079) );
  AND U35637 ( .A(n17080), .B(n17079), .Z(n17082) );
  NANDN U35638 ( .A(y[5042]), .B(x[5042]), .Z(n17081) );
  NANDN U35639 ( .A(y[5043]), .B(x[5043]), .Z(n24558) );
  NAND U35640 ( .A(n17081), .B(n24558), .Z(n51500) );
  OR U35641 ( .A(n17082), .B(n51500), .Z(n17083) );
  NAND U35642 ( .A(n51499), .B(n17083), .Z(n17084) );
  NANDN U35643 ( .A(n57380), .B(n17084), .Z(n17085) );
  AND U35644 ( .A(n24555), .B(n17085), .Z(n17086) );
  NANDN U35645 ( .A(x[5045]), .B(y[5045]), .Z(n57382) );
  AND U35646 ( .A(n17086), .B(n57382), .Z(n17088) );
  NANDN U35647 ( .A(y[5046]), .B(x[5046]), .Z(n17087) );
  NANDN U35648 ( .A(y[5047]), .B(x[5047]), .Z(n24552) );
  NAND U35649 ( .A(n17087), .B(n24552), .Z(n57383) );
  OR U35650 ( .A(n17088), .B(n57383), .Z(n17089) );
  AND U35651 ( .A(n57384), .B(n17089), .Z(n17090) );
  NANDN U35652 ( .A(y[5048]), .B(x[5048]), .Z(n24551) );
  NANDN U35653 ( .A(y[5049]), .B(x[5049]), .Z(n24548) );
  NAND U35654 ( .A(n24551), .B(n24548), .Z(n57385) );
  OR U35655 ( .A(n17090), .B(n57385), .Z(n17091) );
  NANDN U35656 ( .A(x[5049]), .B(y[5049]), .Z(n51497) );
  AND U35657 ( .A(n17091), .B(n51497), .Z(n17092) );
  XNOR U35658 ( .A(x[5050]), .B(y[5050]), .Z(n24549) );
  NAND U35659 ( .A(n17092), .B(n24549), .Z(n17093) );
  NANDN U35660 ( .A(n57386), .B(n17093), .Z(n17094) );
  AND U35661 ( .A(n43010), .B(n17094), .Z(n17095) );
  NANDN U35662 ( .A(x[5051]), .B(y[5051]), .Z(n57387) );
  AND U35663 ( .A(n17095), .B(n57387), .Z(n17096) );
  OR U35664 ( .A(n57389), .B(n17096), .Z(n17097) );
  AND U35665 ( .A(n24547), .B(n17097), .Z(n17098) );
  ANDN U35666 ( .B(y[5053]), .A(x[5053]), .Z(n57390) );
  ANDN U35667 ( .B(n17098), .A(n57390), .Z(n17100) );
  NANDN U35668 ( .A(y[5054]), .B(x[5054]), .Z(n17099) );
  NANDN U35669 ( .A(y[5055]), .B(x[5055]), .Z(n24544) );
  NAND U35670 ( .A(n17099), .B(n24544), .Z(n57393) );
  OR U35671 ( .A(n17100), .B(n57393), .Z(n17101) );
  AND U35672 ( .A(n57394), .B(n17101), .Z(n17102) );
  OR U35673 ( .A(n57395), .B(n17102), .Z(n17103) );
  NAND U35674 ( .A(n57396), .B(n17103), .Z(n17104) );
  NANDN U35675 ( .A(n57397), .B(n17104), .Z(n17105) );
  AND U35676 ( .A(n43028), .B(n17105), .Z(n17106) );
  NANDN U35677 ( .A(x[5059]), .B(y[5059]), .Z(n57398) );
  AND U35678 ( .A(n17106), .B(n57398), .Z(n17108) );
  NANDN U35679 ( .A(y[5060]), .B(x[5060]), .Z(n17107) );
  NANDN U35680 ( .A(y[5061]), .B(x[5061]), .Z(n24536) );
  AND U35681 ( .A(n17107), .B(n24536), .Z(n57400) );
  NANDN U35682 ( .A(n17108), .B(n57400), .Z(n17109) );
  NAND U35683 ( .A(n17110), .B(n17109), .Z(n17111) );
  AND U35684 ( .A(n57401), .B(n17111), .Z(n17112) );
  ANDN U35685 ( .B(n57403), .A(n17112), .Z(n17113) );
  NAND U35686 ( .A(n43038), .B(n17113), .Z(n17114) );
  NANDN U35687 ( .A(n57404), .B(n17114), .Z(n17115) );
  AND U35688 ( .A(n24535), .B(n17115), .Z(n17116) );
  ANDN U35689 ( .B(y[5065]), .A(x[5065]), .Z(n57405) );
  ANDN U35690 ( .B(n17116), .A(n57405), .Z(n17117) );
  OR U35691 ( .A(n57407), .B(n17117), .Z(n17118) );
  AND U35692 ( .A(n43048), .B(n17118), .Z(n17119) );
  NANDN U35693 ( .A(x[5067]), .B(y[5067]), .Z(n57409) );
  AND U35694 ( .A(n17119), .B(n57409), .Z(n17121) );
  NANDN U35695 ( .A(y[5068]), .B(x[5068]), .Z(n17120) );
  NANDN U35696 ( .A(y[5069]), .B(x[5069]), .Z(n24532) );
  NAND U35697 ( .A(n17120), .B(n24532), .Z(n57411) );
  OR U35698 ( .A(n17121), .B(n57411), .Z(n17122) );
  AND U35699 ( .A(n57412), .B(n17122), .Z(n17123) );
  NANDN U35700 ( .A(y[5070]), .B(x[5070]), .Z(n24531) );
  NANDN U35701 ( .A(y[5071]), .B(x[5071]), .Z(n24528) );
  NAND U35702 ( .A(n24531), .B(n24528), .Z(n57413) );
  OR U35703 ( .A(n17123), .B(n57413), .Z(n17124) );
  NAND U35704 ( .A(n17125), .B(n17124), .Z(n17126) );
  NANDN U35705 ( .A(n57416), .B(n17126), .Z(n17127) );
  AND U35706 ( .A(n57417), .B(n17127), .Z(n17128) );
  OR U35707 ( .A(n57418), .B(n17128), .Z(n17129) );
  AND U35708 ( .A(n17130), .B(n17129), .Z(n17131) );
  OR U35709 ( .A(n57419), .B(n17131), .Z(n17132) );
  NAND U35710 ( .A(n57420), .B(n17132), .Z(n17133) );
  NANDN U35711 ( .A(n57422), .B(n17133), .Z(n17134) );
  AND U35712 ( .A(n43076), .B(n17134), .Z(n17135) );
  NANDN U35713 ( .A(x[5079]), .B(y[5079]), .Z(n57423) );
  AND U35714 ( .A(n17135), .B(n57423), .Z(n17137) );
  NANDN U35715 ( .A(y[5080]), .B(x[5080]), .Z(n17136) );
  NANDN U35716 ( .A(y[5081]), .B(x[5081]), .Z(n24518) );
  AND U35717 ( .A(n17136), .B(n24518), .Z(n57425) );
  NANDN U35718 ( .A(n17137), .B(n57425), .Z(n17138) );
  NAND U35719 ( .A(n17139), .B(n17138), .Z(n17140) );
  AND U35720 ( .A(n57426), .B(n17140), .Z(n17141) );
  ANDN U35721 ( .B(n17142), .A(n17141), .Z(n17143) );
  ANDN U35722 ( .B(n51490), .A(n17143), .Z(n17144) );
  NOR U35723 ( .A(n57429), .B(n17144), .Z(n17145) );
  NAND U35724 ( .A(n24517), .B(n17145), .Z(n17146) );
  NANDN U35725 ( .A(n57431), .B(n17146), .Z(n17147) );
  AND U35726 ( .A(n24515), .B(n17147), .Z(n17148) );
  NANDN U35727 ( .A(x[5087]), .B(y[5087]), .Z(n57432) );
  NAND U35728 ( .A(n17148), .B(n57432), .Z(n17149) );
  NANDN U35729 ( .A(n57434), .B(n17149), .Z(n17150) );
  AND U35730 ( .A(n57437), .B(n17150), .Z(n17151) );
  OR U35731 ( .A(n57438), .B(n17151), .Z(n17152) );
  NAND U35732 ( .A(n57439), .B(n17152), .Z(n17153) );
  NANDN U35733 ( .A(n57440), .B(n17153), .Z(n17154) );
  AND U35734 ( .A(n24505), .B(n17154), .Z(n17155) );
  NANDN U35735 ( .A(x[5093]), .B(y[5093]), .Z(n57441) );
  NAND U35736 ( .A(n17155), .B(n57441), .Z(n17157) );
  NANDN U35737 ( .A(y[5094]), .B(x[5094]), .Z(n17156) );
  NANDN U35738 ( .A(y[5095]), .B(x[5095]), .Z(n43112) );
  AND U35739 ( .A(n17156), .B(n43112), .Z(n57443) );
  AND U35740 ( .A(n17157), .B(n57443), .Z(n17158) );
  NOR U35741 ( .A(n43109), .B(n17158), .Z(n17159) );
  NAND U35742 ( .A(n43113), .B(n17159), .Z(n17160) );
  NANDN U35743 ( .A(n57444), .B(n17160), .Z(n17161) );
  AND U35744 ( .A(n57445), .B(n17161), .Z(n17162) );
  OR U35745 ( .A(n57446), .B(n17162), .Z(n17163) );
  NAND U35746 ( .A(n57447), .B(n17163), .Z(n17164) );
  NANDN U35747 ( .A(n57448), .B(n17164), .Z(n17165) );
  AND U35748 ( .A(n57449), .B(n17165), .Z(n17166) );
  OR U35749 ( .A(n57450), .B(n17166), .Z(n17167) );
  NAND U35750 ( .A(n57451), .B(n17167), .Z(n17168) );
  NANDN U35751 ( .A(n57452), .B(n17168), .Z(n17169) );
  AND U35752 ( .A(n24491), .B(n17169), .Z(n17170) );
  NANDN U35753 ( .A(x[5105]), .B(y[5105]), .Z(n57454) );
  AND U35754 ( .A(n17170), .B(n57454), .Z(n17172) );
  NANDN U35755 ( .A(y[5106]), .B(x[5106]), .Z(n17171) );
  NANDN U35756 ( .A(y[5107]), .B(x[5107]), .Z(n24488) );
  NAND U35757 ( .A(n17171), .B(n24488), .Z(n57456) );
  OR U35758 ( .A(n17172), .B(n57456), .Z(n17173) );
  AND U35759 ( .A(n24489), .B(n17173), .Z(n17174) );
  NANDN U35760 ( .A(x[5107]), .B(y[5107]), .Z(n51486) );
  AND U35761 ( .A(n17174), .B(n51486), .Z(n17176) );
  NANDN U35762 ( .A(y[5108]), .B(x[5108]), .Z(n17175) );
  NANDN U35763 ( .A(y[5109]), .B(x[5109]), .Z(n24486) );
  NAND U35764 ( .A(n17175), .B(n24486), .Z(n57457) );
  OR U35765 ( .A(n17176), .B(n57457), .Z(n17177) );
  NAND U35766 ( .A(n17178), .B(n17177), .Z(n17179) );
  AND U35767 ( .A(n57458), .B(n17179), .Z(n17180) );
  NOR U35768 ( .A(n43148), .B(n17180), .Z(n17181) );
  NAND U35769 ( .A(n43152), .B(n17181), .Z(n17182) );
  NANDN U35770 ( .A(n57461), .B(n17182), .Z(n17183) );
  AND U35771 ( .A(n24485), .B(n17183), .Z(n17184) );
  NANDN U35772 ( .A(n57462), .B(n17184), .Z(n17185) );
  NANDN U35773 ( .A(n57464), .B(n17185), .Z(n17186) );
  AND U35774 ( .A(n24483), .B(n17186), .Z(n17187) );
  NANDN U35775 ( .A(x[5115]), .B(y[5115]), .Z(n51482) );
  AND U35776 ( .A(n17187), .B(n51482), .Z(n17189) );
  NANDN U35777 ( .A(y[5116]), .B(x[5116]), .Z(n17188) );
  NANDN U35778 ( .A(y[5117]), .B(x[5117]), .Z(n24480) );
  AND U35779 ( .A(n17188), .B(n24480), .Z(n57466) );
  NANDN U35780 ( .A(n17189), .B(n57466), .Z(n17190) );
  NAND U35781 ( .A(n17191), .B(n17190), .Z(n17192) );
  AND U35782 ( .A(n57470), .B(n17192), .Z(n17193) );
  NANDN U35783 ( .A(x[5119]), .B(y[5119]), .Z(n24479) );
  NANDN U35784 ( .A(x[5120]), .B(y[5120]), .Z(n24476) );
  NAND U35785 ( .A(n24479), .B(n24476), .Z(n57471) );
  OR U35786 ( .A(n17193), .B(n57471), .Z(n17194) );
  AND U35787 ( .A(n57472), .B(n17194), .Z(n17195) );
  OR U35788 ( .A(n57473), .B(n17195), .Z(n17196) );
  NAND U35789 ( .A(n57474), .B(n17196), .Z(n17197) );
  NANDN U35790 ( .A(n57475), .B(n17197), .Z(n17198) );
  AND U35791 ( .A(n57476), .B(n17198), .Z(n17199) );
  XNOR U35792 ( .A(y[5126]), .B(x[5126]), .Z(n24466) );
  NANDN U35793 ( .A(x[5125]), .B(y[5125]), .Z(n24467) );
  NAND U35794 ( .A(n24466), .B(n24467), .Z(n57477) );
  OR U35795 ( .A(n17199), .B(n57477), .Z(n17200) );
  NAND U35796 ( .A(n57478), .B(n17200), .Z(n17201) );
  AND U35797 ( .A(n43187), .B(n17201), .Z(n17202) );
  NANDN U35798 ( .A(x[5127]), .B(y[5127]), .Z(n51480) );
  AND U35799 ( .A(n17202), .B(n51480), .Z(n17204) );
  NANDN U35800 ( .A(y[5128]), .B(x[5128]), .Z(n17203) );
  NANDN U35801 ( .A(y[5129]), .B(x[5129]), .Z(n24463) );
  AND U35802 ( .A(n17203), .B(n24463), .Z(n57479) );
  NANDN U35803 ( .A(n17204), .B(n57479), .Z(n17205) );
  NAND U35804 ( .A(n17206), .B(n17205), .Z(n17208) );
  NANDN U35805 ( .A(y[5130]), .B(x[5130]), .Z(n17207) );
  NANDN U35806 ( .A(y[5131]), .B(x[5131]), .Z(n43197) );
  AND U35807 ( .A(n17207), .B(n43197), .Z(n51479) );
  AND U35808 ( .A(n17208), .B(n51479), .Z(n17209) );
  NOR U35809 ( .A(n43194), .B(n17209), .Z(n17210) );
  NAND U35810 ( .A(n43198), .B(n17210), .Z(n17211) );
  NANDN U35811 ( .A(n57486), .B(n17211), .Z(n17212) );
  AND U35812 ( .A(n24462), .B(n17212), .Z(n17213) );
  ANDN U35813 ( .B(y[5133]), .A(x[5133]), .Z(n57487) );
  ANDN U35814 ( .B(n17213), .A(n57487), .Z(n17215) );
  NANDN U35815 ( .A(y[5134]), .B(x[5134]), .Z(n17214) );
  NANDN U35816 ( .A(y[5135]), .B(x[5135]), .Z(n43208) );
  AND U35817 ( .A(n17214), .B(n43208), .Z(n57489) );
  NANDN U35818 ( .A(n17215), .B(n57489), .Z(n17216) );
  NAND U35819 ( .A(n43209), .B(n17216), .Z(n17217) );
  ANDN U35820 ( .B(y[5135]), .A(x[5135]), .Z(n43205) );
  OR U35821 ( .A(n17217), .B(n43205), .Z(n17218) );
  NAND U35822 ( .A(n57490), .B(n17218), .Z(n17220) );
  NANDN U35823 ( .A(x[5137]), .B(y[5137]), .Z(n24460) );
  XNOR U35824 ( .A(x[5138]), .B(y[5138]), .Z(n24459) );
  NAND U35825 ( .A(n24460), .B(n24459), .Z(n17219) );
  ANDN U35826 ( .B(n17220), .A(n17219), .Z(n17222) );
  NANDN U35827 ( .A(y[5138]), .B(x[5138]), .Z(n17221) );
  NANDN U35828 ( .A(y[5139]), .B(x[5139]), .Z(n24456) );
  NAND U35829 ( .A(n17221), .B(n24456), .Z(n57493) );
  OR U35830 ( .A(n17222), .B(n57493), .Z(n17223) );
  NAND U35831 ( .A(n57494), .B(n17223), .Z(n17224) );
  NANDN U35832 ( .A(n51476), .B(n17224), .Z(n17225) );
  XNOR U35833 ( .A(y[5142]), .B(x[5142]), .Z(n24452) );
  NANDN U35834 ( .A(x[5141]), .B(y[5141]), .Z(n24453) );
  AND U35835 ( .A(n24452), .B(n24453), .Z(n51475) );
  AND U35836 ( .A(n17225), .B(n51475), .Z(n17227) );
  NANDN U35837 ( .A(y[5142]), .B(x[5142]), .Z(n17226) );
  NANDN U35838 ( .A(y[5143]), .B(x[5143]), .Z(n24448) );
  NAND U35839 ( .A(n17226), .B(n24448), .Z(n57497) );
  OR U35840 ( .A(n17227), .B(n57497), .Z(n17228) );
  AND U35841 ( .A(n57498), .B(n17228), .Z(n17229) );
  NANDN U35842 ( .A(y[5144]), .B(x[5144]), .Z(n24447) );
  NANDN U35843 ( .A(y[5145]), .B(x[5145]), .Z(n24444) );
  NAND U35844 ( .A(n24447), .B(n24444), .Z(n57499) );
  OR U35845 ( .A(n17229), .B(n57499), .Z(n17230) );
  AND U35846 ( .A(n57500), .B(n17230), .Z(n17232) );
  NAND U35847 ( .A(n17232), .B(n17231), .Z(n17233) );
  NANDN U35848 ( .A(n57502), .B(n17233), .Z(n17234) );
  AND U35849 ( .A(n43236), .B(n17234), .Z(n17235) );
  NANDN U35850 ( .A(n43232), .B(n17235), .Z(n17236) );
  NAND U35851 ( .A(n57503), .B(n17236), .Z(n17237) );
  NANDN U35852 ( .A(n51472), .B(n17237), .Z(n17238) );
  AND U35853 ( .A(n57504), .B(n17238), .Z(n17239) );
  ANDN U35854 ( .B(n57505), .A(n17239), .Z(n17240) );
  NAND U35855 ( .A(n43247), .B(n17240), .Z(n17241) );
  NANDN U35856 ( .A(n51471), .B(n17241), .Z(n17242) );
  NANDN U35857 ( .A(x[5153]), .B(y[5153]), .Z(n24440) );
  NANDN U35858 ( .A(x[5154]), .B(y[5154]), .Z(n24437) );
  AND U35859 ( .A(n24440), .B(n24437), .Z(n51470) );
  AND U35860 ( .A(n17242), .B(n51470), .Z(n17243) );
  NANDN U35861 ( .A(y[5154]), .B(x[5154]), .Z(n24438) );
  NANDN U35862 ( .A(y[5155]), .B(x[5155]), .Z(n24435) );
  NAND U35863 ( .A(n24438), .B(n24435), .Z(n57509) );
  OR U35864 ( .A(n17243), .B(n57509), .Z(n17244) );
  AND U35865 ( .A(n24436), .B(n17244), .Z(n17245) );
  NANDN U35866 ( .A(x[5155]), .B(y[5155]), .Z(n57510) );
  AND U35867 ( .A(n17245), .B(n57510), .Z(n17247) );
  NANDN U35868 ( .A(y[5156]), .B(x[5156]), .Z(n17246) );
  NANDN U35869 ( .A(y[5157]), .B(x[5157]), .Z(n24433) );
  NAND U35870 ( .A(n17246), .B(n24433), .Z(n57512) );
  OR U35871 ( .A(n17247), .B(n57512), .Z(n17248) );
  AND U35872 ( .A(n17249), .B(n17248), .Z(n17250) );
  OR U35873 ( .A(n57515), .B(n17250), .Z(n17251) );
  NAND U35874 ( .A(n57516), .B(n17251), .Z(n17252) );
  NANDN U35875 ( .A(n57517), .B(n17252), .Z(n17253) );
  AND U35876 ( .A(n57518), .B(n17253), .Z(n17254) );
  OR U35877 ( .A(n57519), .B(n17254), .Z(n17255) );
  NAND U35878 ( .A(n17256), .B(n17255), .Z(n17258) );
  NANDN U35879 ( .A(y[5164]), .B(x[5164]), .Z(n17257) );
  NANDN U35880 ( .A(y[5165]), .B(x[5165]), .Z(n24423) );
  AND U35881 ( .A(n17257), .B(n24423), .Z(n57522) );
  AND U35882 ( .A(n17258), .B(n57522), .Z(n17259) );
  NOR U35883 ( .A(n24425), .B(n17259), .Z(n17260) );
  NAND U35884 ( .A(n24424), .B(n17260), .Z(n17261) );
  NANDN U35885 ( .A(n57524), .B(n17261), .Z(n17262) );
  AND U35886 ( .A(n57525), .B(n17262), .Z(n17263) );
  NANDN U35887 ( .A(y[5168]), .B(x[5168]), .Z(n24421) );
  NANDN U35888 ( .A(y[5169]), .B(x[5169]), .Z(n24418) );
  NAND U35889 ( .A(n24421), .B(n24418), .Z(n57526) );
  OR U35890 ( .A(n17263), .B(n57526), .Z(n17264) );
  AND U35891 ( .A(n24419), .B(n17264), .Z(n17265) );
  NANDN U35892 ( .A(x[5169]), .B(y[5169]), .Z(n57527) );
  AND U35893 ( .A(n17265), .B(n57527), .Z(n17267) );
  NANDN U35894 ( .A(y[5170]), .B(x[5170]), .Z(n17266) );
  NANDN U35895 ( .A(y[5171]), .B(x[5171]), .Z(n43292) );
  NAND U35896 ( .A(n17266), .B(n43292), .Z(n57529) );
  OR U35897 ( .A(n17267), .B(n57529), .Z(n17268) );
  NAND U35898 ( .A(n17269), .B(n17268), .Z(n17270) );
  AND U35899 ( .A(n57530), .B(n17270), .Z(n17271) );
  NOR U35900 ( .A(n57532), .B(n17271), .Z(n17272) );
  NAND U35901 ( .A(n24417), .B(n17272), .Z(n17273) );
  NANDN U35902 ( .A(n57533), .B(n17273), .Z(n17274) );
  AND U35903 ( .A(n43304), .B(n17274), .Z(n17275) );
  NANDN U35904 ( .A(n43300), .B(n17275), .Z(n17276) );
  NAND U35905 ( .A(n57536), .B(n17276), .Z(n17277) );
  NANDN U35906 ( .A(n57537), .B(n17277), .Z(n17278) );
  AND U35907 ( .A(n57538), .B(n17278), .Z(n17279) );
  ANDN U35908 ( .B(n17280), .A(n17279), .Z(n17281) );
  ANDN U35909 ( .B(n51465), .A(n17281), .Z(n17282) );
  NOR U35910 ( .A(n57543), .B(n17282), .Z(n17283) );
  NAND U35911 ( .A(n24411), .B(n17283), .Z(n17284) );
  NANDN U35912 ( .A(n57545), .B(n17284), .Z(n17285) );
  XOR U35913 ( .A(x[5184]), .B(y[5184]), .Z(n43326) );
  ANDN U35914 ( .B(n17285), .A(n43326), .Z(n17286) );
  NANDN U35915 ( .A(n24409), .B(n17286), .Z(n17287) );
  NAND U35916 ( .A(n57548), .B(n17287), .Z(n17288) );
  NANDN U35917 ( .A(n57549), .B(n17288), .Z(n17289) );
  NANDN U35918 ( .A(y[5186]), .B(x[5186]), .Z(n24406) );
  NANDN U35919 ( .A(y[5187]), .B(x[5187]), .Z(n43333) );
  AND U35920 ( .A(n24406), .B(n43333), .Z(n57550) );
  AND U35921 ( .A(n17289), .B(n57550), .Z(n17290) );
  NOR U35922 ( .A(n24404), .B(n17290), .Z(n17291) );
  NAND U35923 ( .A(n43334), .B(n17291), .Z(n17292) );
  NANDN U35924 ( .A(n51462), .B(n17292), .Z(n17293) );
  AND U35925 ( .A(n57552), .B(n17293), .Z(n17294) );
  NANDN U35926 ( .A(y[5190]), .B(x[5190]), .Z(n24401) );
  NANDN U35927 ( .A(y[5191]), .B(x[5191]), .Z(n24398) );
  NAND U35928 ( .A(n24401), .B(n24398), .Z(n57553) );
  OR U35929 ( .A(n17294), .B(n57553), .Z(n17295) );
  AND U35930 ( .A(n24399), .B(n17295), .Z(n17296) );
  NANDN U35931 ( .A(x[5191]), .B(y[5191]), .Z(n51460) );
  AND U35932 ( .A(n17296), .B(n51460), .Z(n17298) );
  NANDN U35933 ( .A(y[5192]), .B(x[5192]), .Z(n17297) );
  NANDN U35934 ( .A(y[5193]), .B(x[5193]), .Z(n24396) );
  NAND U35935 ( .A(n17297), .B(n24396), .Z(n57555) );
  OR U35936 ( .A(n17298), .B(n57555), .Z(n17299) );
  NAND U35937 ( .A(n17300), .B(n17299), .Z(n17302) );
  NANDN U35938 ( .A(y[5194]), .B(x[5194]), .Z(n17301) );
  NANDN U35939 ( .A(y[5195]), .B(x[5195]), .Z(n43352) );
  AND U35940 ( .A(n17301), .B(n43352), .Z(n51459) );
  AND U35941 ( .A(n17302), .B(n51459), .Z(n17303) );
  NOR U35942 ( .A(n43349), .B(n17303), .Z(n17304) );
  NAND U35943 ( .A(n43353), .B(n17304), .Z(n17305) );
  NANDN U35944 ( .A(n57560), .B(n17305), .Z(n17306) );
  AND U35945 ( .A(n24395), .B(n17306), .Z(n17307) );
  ANDN U35946 ( .B(y[5197]), .A(x[5197]), .Z(n57561) );
  ANDN U35947 ( .B(n17307), .A(n57561), .Z(n17309) );
  NANDN U35948 ( .A(y[5198]), .B(x[5198]), .Z(n17308) );
  NANDN U35949 ( .A(y[5199]), .B(x[5199]), .Z(n43363) );
  AND U35950 ( .A(n17308), .B(n43363), .Z(n57563) );
  NANDN U35951 ( .A(n17309), .B(n57563), .Z(n17310) );
  NAND U35952 ( .A(n43364), .B(n17310), .Z(n17311) );
  ANDN U35953 ( .B(y[5199]), .A(x[5199]), .Z(n43360) );
  OR U35954 ( .A(n17311), .B(n43360), .Z(n17312) );
  NAND U35955 ( .A(n57566), .B(n17312), .Z(n17313) );
  NANDN U35956 ( .A(n51456), .B(n17313), .Z(n17314) );
  ANDN U35957 ( .B(n24393), .A(n17314), .Z(n17316) );
  NANDN U35958 ( .A(y[5202]), .B(x[5202]), .Z(n17315) );
  NANDN U35959 ( .A(y[5203]), .B(x[5203]), .Z(n24390) );
  NAND U35960 ( .A(n17315), .B(n24390), .Z(n57567) );
  OR U35961 ( .A(n17316), .B(n57567), .Z(n17317) );
  NAND U35962 ( .A(n57568), .B(n17317), .Z(n17318) );
  NANDN U35963 ( .A(n51454), .B(n17318), .Z(n17319) );
  NANDN U35964 ( .A(x[5205]), .B(y[5205]), .Z(n24387) );
  NANDN U35965 ( .A(x[5206]), .B(y[5206]), .Z(n24384) );
  AND U35966 ( .A(n24387), .B(n24384), .Z(n51453) );
  AND U35967 ( .A(n17319), .B(n51453), .Z(n17320) );
  NANDN U35968 ( .A(y[5206]), .B(x[5206]), .Z(n24385) );
  NANDN U35969 ( .A(y[5207]), .B(x[5207]), .Z(n43381) );
  NAND U35970 ( .A(n24385), .B(n43381), .Z(n57569) );
  OR U35971 ( .A(n17320), .B(n57569), .Z(n17321) );
  NAND U35972 ( .A(n17322), .B(n17321), .Z(n17324) );
  NANDN U35973 ( .A(y[5208]), .B(x[5208]), .Z(n17323) );
  NANDN U35974 ( .A(y[5209]), .B(x[5209]), .Z(n24382) );
  AND U35975 ( .A(n17323), .B(n24382), .Z(n51452) );
  AND U35976 ( .A(n17324), .B(n51452), .Z(n17325) );
  NOR U35977 ( .A(n57572), .B(n17325), .Z(n17326) );
  NAND U35978 ( .A(n24383), .B(n17326), .Z(n17327) );
  NANDN U35979 ( .A(n57576), .B(n17327), .Z(n17328) );
  AND U35980 ( .A(n43392), .B(n17328), .Z(n17329) );
  NANDN U35981 ( .A(x[5211]), .B(y[5211]), .Z(n51450) );
  AND U35982 ( .A(n17329), .B(n51450), .Z(n17331) );
  NANDN U35983 ( .A(y[5212]), .B(x[5212]), .Z(n17330) );
  NANDN U35984 ( .A(y[5213]), .B(x[5213]), .Z(n24380) );
  NAND U35985 ( .A(n17330), .B(n24380), .Z(n57577) );
  OR U35986 ( .A(n17331), .B(n57577), .Z(n17332) );
  AND U35987 ( .A(n24381), .B(n17332), .Z(n17333) );
  NANDN U35988 ( .A(x[5213]), .B(y[5213]), .Z(n57579) );
  AND U35989 ( .A(n17333), .B(n57579), .Z(n17334) );
  OR U35990 ( .A(n57580), .B(n17334), .Z(n17335) );
  AND U35991 ( .A(n17336), .B(n17335), .Z(n17338) );
  NANDN U35992 ( .A(y[5216]), .B(x[5216]), .Z(n17337) );
  NANDN U35993 ( .A(y[5217]), .B(x[5217]), .Z(n24375) );
  NAND U35994 ( .A(n17337), .B(n24375), .Z(n51448) );
  OR U35995 ( .A(n17338), .B(n51448), .Z(n17339) );
  NAND U35996 ( .A(n51447), .B(n17339), .Z(n17340) );
  NANDN U35997 ( .A(n57582), .B(n17340), .Z(n17341) );
  NAND U35998 ( .A(n43411), .B(n17341), .Z(n17342) );
  NANDN U35999 ( .A(x[5219]), .B(y[5219]), .Z(n57586) );
  NANDN U36000 ( .A(n17342), .B(n57586), .Z(n17343) );
  NAND U36001 ( .A(n51446), .B(n17343), .Z(n17344) );
  NANDN U36002 ( .A(n57587), .B(n17344), .Z(n17345) );
  AND U36003 ( .A(n57588), .B(n17345), .Z(n17347) );
  NANDN U36004 ( .A(x[5223]), .B(y[5223]), .Z(n51444) );
  XNOR U36005 ( .A(x[5224]), .B(y[5224]), .Z(n43422) );
  NAND U36006 ( .A(n51444), .B(n43422), .Z(n17346) );
  OR U36007 ( .A(n17347), .B(n17346), .Z(n17348) );
  AND U36008 ( .A(n57589), .B(n17348), .Z(n17349) );
  XNOR U36009 ( .A(x[5226]), .B(y[5226]), .Z(n24371) );
  NANDN U36010 ( .A(n17349), .B(n24371), .Z(n17350) );
  ANDN U36011 ( .B(y[5225]), .A(x[5225]), .Z(n57591) );
  OR U36012 ( .A(n17350), .B(n57591), .Z(n17351) );
  NAND U36013 ( .A(n51443), .B(n17351), .Z(n17352) );
  NANDN U36014 ( .A(n57592), .B(n17352), .Z(n17353) );
  AND U36015 ( .A(n57593), .B(n17353), .Z(n17354) );
  OR U36016 ( .A(n17355), .B(n17354), .Z(n17356) );
  NAND U36017 ( .A(n57596), .B(n17356), .Z(n17357) );
  NAND U36018 ( .A(n43440), .B(n17357), .Z(n17358) );
  NANDN U36019 ( .A(x[5231]), .B(y[5231]), .Z(n57598) );
  NANDN U36020 ( .A(n17358), .B(n57598), .Z(n17359) );
  NAND U36021 ( .A(n57599), .B(n17359), .Z(n17360) );
  AND U36022 ( .A(n57600), .B(n17360), .Z(n17361) );
  NANDN U36023 ( .A(y[5234]), .B(x[5234]), .Z(n24361) );
  NANDN U36024 ( .A(y[5235]), .B(x[5235]), .Z(n43449) );
  AND U36025 ( .A(n24361), .B(n43449), .Z(n57601) );
  NANDN U36026 ( .A(n17361), .B(n57601), .Z(n17362) );
  NAND U36027 ( .A(n17363), .B(n17362), .Z(n17364) );
  AND U36028 ( .A(n57604), .B(n17364), .Z(n17365) );
  NOR U36029 ( .A(n57606), .B(n17365), .Z(n17366) );
  NAND U36030 ( .A(n24359), .B(n17366), .Z(n17367) );
  NANDN U36031 ( .A(n57607), .B(n17367), .Z(n17368) );
  AND U36032 ( .A(n43460), .B(n17368), .Z(n17369) );
  NANDN U36033 ( .A(x[5239]), .B(y[5239]), .Z(n57608) );
  NAND U36034 ( .A(n17369), .B(n57608), .Z(n17370) );
  NANDN U36035 ( .A(n57610), .B(n17370), .Z(n17371) );
  AND U36036 ( .A(n24357), .B(n17371), .Z(n17372) );
  ANDN U36037 ( .B(y[5241]), .A(x[5241]), .Z(n57611) );
  ANDN U36038 ( .B(n17372), .A(n57611), .Z(n17374) );
  NANDN U36039 ( .A(y[5242]), .B(x[5242]), .Z(n17373) );
  NANDN U36040 ( .A(y[5243]), .B(x[5243]), .Z(n24354) );
  NAND U36041 ( .A(n17373), .B(n24354), .Z(n57613) );
  OR U36042 ( .A(n17374), .B(n57613), .Z(n17375) );
  NAND U36043 ( .A(n57615), .B(n17375), .Z(n17376) );
  AND U36044 ( .A(n57616), .B(n17376), .Z(n17377) );
  ANDN U36045 ( .B(n57618), .A(n17377), .Z(n17378) );
  NAND U36046 ( .A(n24351), .B(n17378), .Z(n17379) );
  NANDN U36047 ( .A(n57619), .B(n17379), .Z(n17380) );
  AND U36048 ( .A(n24349), .B(n17380), .Z(n17381) );
  NANDN U36049 ( .A(n43475), .B(n17381), .Z(n17382) );
  NAND U36050 ( .A(n57621), .B(n17382), .Z(n17383) );
  NANDN U36051 ( .A(n57622), .B(n17383), .Z(n17384) );
  AND U36052 ( .A(n57623), .B(n17384), .Z(n17386) );
  XNOR U36053 ( .A(x[5252]), .B(y[5252]), .Z(n24344) );
  NANDN U36054 ( .A(x[5251]), .B(y[5251]), .Z(n57625) );
  AND U36055 ( .A(n24344), .B(n57625), .Z(n17385) );
  NANDN U36056 ( .A(n17386), .B(n17385), .Z(n17388) );
  NANDN U36057 ( .A(y[5252]), .B(x[5252]), .Z(n17387) );
  NANDN U36058 ( .A(y[5253]), .B(x[5253]), .Z(n24340) );
  AND U36059 ( .A(n17387), .B(n24340), .Z(n51439) );
  AND U36060 ( .A(n17388), .B(n51439), .Z(n17389) );
  NOR U36061 ( .A(n24342), .B(n17389), .Z(n17390) );
  NAND U36062 ( .A(n24341), .B(n17390), .Z(n17391) );
  NANDN U36063 ( .A(n57628), .B(n17391), .Z(n17392) );
  AND U36064 ( .A(n43497), .B(n17392), .Z(n17393) );
  NANDN U36065 ( .A(n43493), .B(n17393), .Z(n17394) );
  NAND U36066 ( .A(n57632), .B(n17394), .Z(n17395) );
  NANDN U36067 ( .A(n57633), .B(n17395), .Z(n17396) );
  NANDN U36068 ( .A(y[5258]), .B(x[5258]), .Z(n24337) );
  NANDN U36069 ( .A(y[5259]), .B(x[5259]), .Z(n43506) );
  AND U36070 ( .A(n24337), .B(n43506), .Z(n57634) );
  AND U36071 ( .A(n17396), .B(n57634), .Z(n17397) );
  NOR U36072 ( .A(n24335), .B(n17397), .Z(n17398) );
  NAND U36073 ( .A(n43507), .B(n17398), .Z(n17399) );
  NANDN U36074 ( .A(n57637), .B(n17399), .Z(n17400) );
  AND U36075 ( .A(n24334), .B(n17400), .Z(n17401) );
  NANDN U36076 ( .A(n57638), .B(n17401), .Z(n17402) );
  NAND U36077 ( .A(n57640), .B(n17402), .Z(n17403) );
  NAND U36078 ( .A(n43518), .B(n17403), .Z(n17404) );
  ANDN U36079 ( .B(y[5263]), .A(x[5263]), .Z(n43514) );
  OR U36080 ( .A(n17404), .B(n43514), .Z(n17405) );
  NAND U36081 ( .A(n57641), .B(n17405), .Z(n17407) );
  NANDN U36082 ( .A(x[5265]), .B(y[5265]), .Z(n24332) );
  XNOR U36083 ( .A(x[5266]), .B(y[5266]), .Z(n24331) );
  NAND U36084 ( .A(n24332), .B(n24331), .Z(n17406) );
  ANDN U36085 ( .B(n17407), .A(n17406), .Z(n17409) );
  NANDN U36086 ( .A(y[5266]), .B(x[5266]), .Z(n17408) );
  NANDN U36087 ( .A(y[5267]), .B(x[5267]), .Z(n24328) );
  NAND U36088 ( .A(n17408), .B(n24328), .Z(n57646) );
  OR U36089 ( .A(n17409), .B(n57646), .Z(n17410) );
  NAND U36090 ( .A(n57648), .B(n17410), .Z(n17411) );
  NANDN U36091 ( .A(n51436), .B(n17411), .Z(n17412) );
  XNOR U36092 ( .A(y[5270]), .B(x[5270]), .Z(n24324) );
  NANDN U36093 ( .A(x[5269]), .B(y[5269]), .Z(n24325) );
  AND U36094 ( .A(n24324), .B(n24325), .Z(n51435) );
  AND U36095 ( .A(n17412), .B(n51435), .Z(n17414) );
  ANDN U36096 ( .B(x[5271]), .A(y[5271]), .Z(n43537) );
  NANDN U36097 ( .A(y[5270]), .B(x[5270]), .Z(n17413) );
  NANDN U36098 ( .A(n43537), .B(n17413), .Z(n57649) );
  OR U36099 ( .A(n17414), .B(n57649), .Z(n17415) );
  AND U36100 ( .A(n17416), .B(n17415), .Z(n17418) );
  NANDN U36101 ( .A(y[5272]), .B(x[5272]), .Z(n17417) );
  NANDN U36102 ( .A(y[5273]), .B(x[5273]), .Z(n24321) );
  NAND U36103 ( .A(n17417), .B(n24321), .Z(n57652) );
  OR U36104 ( .A(n17418), .B(n57652), .Z(n17419) );
  NAND U36105 ( .A(n57653), .B(n17419), .Z(n17420) );
  NANDN U36106 ( .A(n51434), .B(n17420), .Z(n17421) );
  NANDN U36107 ( .A(x[5275]), .B(y[5275]), .Z(n24318) );
  NANDN U36108 ( .A(x[5276]), .B(y[5276]), .Z(n24315) );
  AND U36109 ( .A(n24318), .B(n24315), .Z(n51433) );
  AND U36110 ( .A(n17421), .B(n51433), .Z(n17422) );
  NANDN U36111 ( .A(y[5276]), .B(x[5276]), .Z(n24316) );
  NANDN U36112 ( .A(y[5277]), .B(x[5277]), .Z(n24313) );
  NAND U36113 ( .A(n24316), .B(n24313), .Z(n57654) );
  OR U36114 ( .A(n17422), .B(n57654), .Z(n17423) );
  AND U36115 ( .A(n17424), .B(n17423), .Z(n17426) );
  NANDN U36116 ( .A(y[5278]), .B(x[5278]), .Z(n17425) );
  NANDN U36117 ( .A(y[5279]), .B(x[5279]), .Z(n24312) );
  NAND U36118 ( .A(n17425), .B(n24312), .Z(n57660) );
  OR U36119 ( .A(n17426), .B(n57660), .Z(n17427) );
  NANDN U36120 ( .A(x[5281]), .B(y[5281]), .Z(n24309) );
  NANDN U36121 ( .A(x[5282]), .B(y[5282]), .Z(n24306) );
  AND U36122 ( .A(n24309), .B(n24306), .Z(n51431) );
  NANDN U36123 ( .A(y[5282]), .B(x[5282]), .Z(n24307) );
  NANDN U36124 ( .A(y[5283]), .B(x[5283]), .Z(n43563) );
  NAND U36125 ( .A(n24307), .B(n43563), .Z(n57662) );
  NANDN U36126 ( .A(y[5284]), .B(x[5284]), .Z(n17428) );
  NANDN U36127 ( .A(y[5285]), .B(x[5285]), .Z(n24304) );
  NAND U36128 ( .A(n17428), .B(n24304), .Z(n57665) );
  NANDN U36129 ( .A(x[5287]), .B(y[5287]), .Z(n24301) );
  NANDN U36130 ( .A(x[5288]), .B(y[5288]), .Z(n43577) );
  AND U36131 ( .A(n24301), .B(n43577), .Z(n51429) );
  NANDN U36132 ( .A(y[5288]), .B(x[5288]), .Z(n24299) );
  NANDN U36133 ( .A(y[5289]), .B(x[5289]), .Z(n24298) );
  NAND U36134 ( .A(n24299), .B(n24298), .Z(n57669) );
  NANDN U36135 ( .A(y[5290]), .B(x[5290]), .Z(n24297) );
  NANDN U36136 ( .A(y[5291]), .B(x[5291]), .Z(n24294) );
  NAND U36137 ( .A(n24297), .B(n24294), .Z(n57672) );
  NANDN U36138 ( .A(y[5294]), .B(x[5294]), .Z(n24291) );
  NANDN U36139 ( .A(y[5295]), .B(x[5295]), .Z(n24288) );
  NAND U36140 ( .A(n24291), .B(n24288), .Z(n57677) );
  AND U36141 ( .A(n57678), .B(n17429), .Z(n17430) );
  OR U36142 ( .A(n57679), .B(n17430), .Z(n17431) );
  NAND U36143 ( .A(n57680), .B(n17431), .Z(n17432) );
  NANDN U36144 ( .A(n57681), .B(n17432), .Z(n17433) );
  NAND U36145 ( .A(n43600), .B(n17433), .Z(n17434) );
  ANDN U36146 ( .B(y[5299]), .A(x[5299]), .Z(n24281) );
  OR U36147 ( .A(n17434), .B(n24281), .Z(n17435) );
  NAND U36148 ( .A(n57682), .B(n17435), .Z(n17436) );
  NANDN U36149 ( .A(n57683), .B(n17436), .Z(n17437) );
  NANDN U36150 ( .A(y[5302]), .B(x[5302]), .Z(n24278) );
  NANDN U36151 ( .A(y[5303]), .B(x[5303]), .Z(n43609) );
  AND U36152 ( .A(n24278), .B(n43609), .Z(n51426) );
  AND U36153 ( .A(n17437), .B(n51426), .Z(n17438) );
  NOR U36154 ( .A(n24276), .B(n17438), .Z(n17439) );
  NAND U36155 ( .A(n43610), .B(n17439), .Z(n17440) );
  NANDN U36156 ( .A(n57687), .B(n17440), .Z(n17441) );
  AND U36157 ( .A(n24275), .B(n17441), .Z(n17442) );
  ANDN U36158 ( .B(y[5305]), .A(x[5305]), .Z(n51424) );
  ANDN U36159 ( .B(n17442), .A(n51424), .Z(n17444) );
  NANDN U36160 ( .A(y[5306]), .B(x[5306]), .Z(n17443) );
  NANDN U36161 ( .A(y[5307]), .B(x[5307]), .Z(n24272) );
  NAND U36162 ( .A(n17443), .B(n24272), .Z(n51423) );
  OR U36163 ( .A(n17444), .B(n51423), .Z(n17445) );
  AND U36164 ( .A(n24273), .B(n17445), .Z(n17446) );
  NANDN U36165 ( .A(x[5307]), .B(y[5307]), .Z(n57689) );
  AND U36166 ( .A(n17446), .B(n57689), .Z(n17448) );
  NANDN U36167 ( .A(y[5308]), .B(x[5308]), .Z(n17447) );
  NANDN U36168 ( .A(y[5309]), .B(x[5309]), .Z(n24270) );
  NAND U36169 ( .A(n17447), .B(n24270), .Z(n57690) );
  OR U36170 ( .A(n17448), .B(n57690), .Z(n17449) );
  AND U36171 ( .A(n57691), .B(n17449), .Z(n17450) );
  OR U36172 ( .A(n57692), .B(n17450), .Z(n17451) );
  NANDN U36173 ( .A(y[5314]), .B(x[5314]), .Z(n24265) );
  NANDN U36174 ( .A(y[5315]), .B(x[5315]), .Z(n24261) );
  AND U36175 ( .A(n24265), .B(n24261), .Z(n51420) );
  NANDN U36176 ( .A(y[5316]), .B(x[5316]), .Z(n17452) );
  NANDN U36177 ( .A(y[5317]), .B(x[5317]), .Z(n24258) );
  AND U36178 ( .A(n17452), .B(n24258), .Z(n57698) );
  NANDN U36179 ( .A(y[5320]), .B(x[5320]), .Z(n24256) );
  NANDN U36180 ( .A(y[5321]), .B(x[5321]), .Z(n24253) );
  AND U36181 ( .A(n24256), .B(n24253), .Z(n51417) );
  AND U36182 ( .A(n57704), .B(n17453), .Z(n17454) );
  NOR U36183 ( .A(n57706), .B(n17454), .Z(n17455) );
  NAND U36184 ( .A(n24252), .B(n17455), .Z(n17456) );
  NANDN U36185 ( .A(n57707), .B(n17456), .Z(n17457) );
  AND U36186 ( .A(n43666), .B(n17457), .Z(n17458) );
  NANDN U36187 ( .A(x[5327]), .B(y[5327]), .Z(n57708) );
  AND U36188 ( .A(n17458), .B(n57708), .Z(n17459) );
  OR U36189 ( .A(n57712), .B(n17459), .Z(n17460) );
  AND U36190 ( .A(n24250), .B(n17460), .Z(n17461) );
  NANDN U36191 ( .A(n57713), .B(n17461), .Z(n17463) );
  NANDN U36192 ( .A(y[5330]), .B(x[5330]), .Z(n17462) );
  NANDN U36193 ( .A(y[5331]), .B(x[5331]), .Z(n24248) );
  AND U36194 ( .A(n17462), .B(n24248), .Z(n57715) );
  AND U36195 ( .A(n17463), .B(n57715), .Z(n17464) );
  NANDN U36196 ( .A(x[5331]), .B(y[5331]), .Z(n43673) );
  NANDN U36197 ( .A(x[5332]), .B(y[5332]), .Z(n24246) );
  AND U36198 ( .A(n43673), .B(n24246), .Z(n57716) );
  NANDN U36199 ( .A(n17464), .B(n57716), .Z(n17465) );
  AND U36200 ( .A(n57717), .B(n17465), .Z(n17466) );
  ANDN U36201 ( .B(n17467), .A(n17466), .Z(n17469) );
  NANDN U36202 ( .A(y[5334]), .B(x[5334]), .Z(n17468) );
  NANDN U36203 ( .A(y[5335]), .B(x[5335]), .Z(n24241) );
  AND U36204 ( .A(n17468), .B(n24241), .Z(n51414) );
  NANDN U36205 ( .A(n17469), .B(n51414), .Z(n17470) );
  NAND U36206 ( .A(n17471), .B(n17470), .Z(n17472) );
  NAND U36207 ( .A(n57721), .B(n17472), .Z(n17473) );
  NANDN U36208 ( .A(x[5337]), .B(y[5337]), .Z(n24240) );
  NANDN U36209 ( .A(x[5338]), .B(y[5338]), .Z(n24237) );
  AND U36210 ( .A(n24240), .B(n24237), .Z(n51412) );
  AND U36211 ( .A(n17473), .B(n51412), .Z(n17474) );
  NANDN U36212 ( .A(y[5338]), .B(x[5338]), .Z(n24238) );
  NANDN U36213 ( .A(y[5339]), .B(x[5339]), .Z(n43692) );
  NAND U36214 ( .A(n24238), .B(n43692), .Z(n57722) );
  OR U36215 ( .A(n17474), .B(n57722), .Z(n17475) );
  AND U36216 ( .A(n17476), .B(n17475), .Z(n17478) );
  NANDN U36217 ( .A(y[5340]), .B(x[5340]), .Z(n17477) );
  NANDN U36218 ( .A(y[5341]), .B(x[5341]), .Z(n24234) );
  NAND U36219 ( .A(n17477), .B(n24234), .Z(n57728) );
  OR U36220 ( .A(n17478), .B(n57728), .Z(n17479) );
  NAND U36221 ( .A(n57729), .B(n17479), .Z(n17480) );
  NANDN U36222 ( .A(n51411), .B(n17480), .Z(n17481) );
  XNOR U36223 ( .A(y[5344]), .B(x[5344]), .Z(n24231) );
  NANDN U36224 ( .A(x[5343]), .B(y[5343]), .Z(n24232) );
  AND U36225 ( .A(n24231), .B(n24232), .Z(n51410) );
  AND U36226 ( .A(n17481), .B(n51410), .Z(n17483) );
  NANDN U36227 ( .A(y[5344]), .B(x[5344]), .Z(n17482) );
  NANDN U36228 ( .A(y[5345]), .B(x[5345]), .Z(n24226) );
  NAND U36229 ( .A(n17482), .B(n24226), .Z(n57730) );
  OR U36230 ( .A(n17483), .B(n57730), .Z(n17484) );
  XNOR U36231 ( .A(y[5346]), .B(x[5346]), .Z(n24227) );
  NANDN U36232 ( .A(x[5345]), .B(y[5345]), .Z(n24228) );
  AND U36233 ( .A(n24227), .B(n24228), .Z(n57731) );
  AND U36234 ( .A(n17484), .B(n57731), .Z(n17486) );
  NANDN U36235 ( .A(y[5346]), .B(x[5346]), .Z(n17485) );
  NANDN U36236 ( .A(y[5347]), .B(x[5347]), .Z(n24222) );
  AND U36237 ( .A(n17485), .B(n24222), .Z(n57732) );
  NANDN U36238 ( .A(n17486), .B(n57732), .Z(n17487) );
  NAND U36239 ( .A(n57733), .B(n17487), .Z(n17488) );
  NANDN U36240 ( .A(n51409), .B(n17488), .Z(n17489) );
  AND U36241 ( .A(n24220), .B(n17489), .Z(n17490) );
  NANDN U36242 ( .A(x[5349]), .B(y[5349]), .Z(n51408) );
  AND U36243 ( .A(n17490), .B(n51408), .Z(n17492) );
  NANDN U36244 ( .A(y[5350]), .B(x[5350]), .Z(n17491) );
  NANDN U36245 ( .A(y[5351]), .B(x[5351]), .Z(n43718) );
  NAND U36246 ( .A(n17491), .B(n43718), .Z(n57737) );
  OR U36247 ( .A(n17492), .B(n57737), .Z(n17493) );
  AND U36248 ( .A(n17494), .B(n17493), .Z(n17496) );
  NANDN U36249 ( .A(y[5352]), .B(x[5352]), .Z(n17495) );
  NANDN U36250 ( .A(y[5353]), .B(x[5353]), .Z(n24217) );
  NAND U36251 ( .A(n17495), .B(n24217), .Z(n57740) );
  OR U36252 ( .A(n17496), .B(n57740), .Z(n17497) );
  NAND U36253 ( .A(n57741), .B(n17497), .Z(n17498) );
  NANDN U36254 ( .A(n51407), .B(n17498), .Z(n17499) );
  NANDN U36255 ( .A(x[5355]), .B(y[5355]), .Z(n24214) );
  NANDN U36256 ( .A(x[5356]), .B(y[5356]), .Z(n43731) );
  AND U36257 ( .A(n24214), .B(n43731), .Z(n51406) );
  AND U36258 ( .A(n17499), .B(n51406), .Z(n17500) );
  NANDN U36259 ( .A(y[5356]), .B(x[5356]), .Z(n24212) );
  NANDN U36260 ( .A(y[5357]), .B(x[5357]), .Z(n24210) );
  NAND U36261 ( .A(n24212), .B(n24210), .Z(n51405) );
  OR U36262 ( .A(n17500), .B(n51405), .Z(n17501) );
  NAND U36263 ( .A(n17502), .B(n17501), .Z(n17504) );
  NANDN U36264 ( .A(y[5358]), .B(x[5358]), .Z(n17503) );
  NANDN U36265 ( .A(y[5359]), .B(x[5359]), .Z(n43738) );
  AND U36266 ( .A(n17503), .B(n43738), .Z(n51404) );
  AND U36267 ( .A(n17504), .B(n51404), .Z(n17505) );
  NOR U36268 ( .A(n43735), .B(n17505), .Z(n17506) );
  NAND U36269 ( .A(n43739), .B(n17506), .Z(n17507) );
  NANDN U36270 ( .A(n57747), .B(n17507), .Z(n17508) );
  AND U36271 ( .A(n24208), .B(n17508), .Z(n17509) );
  NANDN U36272 ( .A(x[5361]), .B(y[5361]), .Z(n24209) );
  AND U36273 ( .A(n17509), .B(n24209), .Z(n17511) );
  NANDN U36274 ( .A(y[5362]), .B(x[5362]), .Z(n17510) );
  NANDN U36275 ( .A(y[5363]), .B(x[5363]), .Z(n43748) );
  NAND U36276 ( .A(n17510), .B(n43748), .Z(n57749) );
  OR U36277 ( .A(n17511), .B(n57749), .Z(n17512) );
  AND U36278 ( .A(n43749), .B(n17512), .Z(n17513) );
  NANDN U36279 ( .A(x[5363]), .B(y[5363]), .Z(n57750) );
  AND U36280 ( .A(n17513), .B(n57750), .Z(n17515) );
  NANDN U36281 ( .A(y[5364]), .B(x[5364]), .Z(n17514) );
  NANDN U36282 ( .A(y[5365]), .B(x[5365]), .Z(n24204) );
  NAND U36283 ( .A(n17514), .B(n24204), .Z(n57752) );
  OR U36284 ( .A(n17515), .B(n57752), .Z(n17516) );
  AND U36285 ( .A(n57753), .B(n17516), .Z(n17518) );
  NANDN U36286 ( .A(y[5366]), .B(x[5366]), .Z(n17517) );
  NANDN U36287 ( .A(y[5367]), .B(x[5367]), .Z(n24200) );
  NAND U36288 ( .A(n17517), .B(n24200), .Z(n51401) );
  OR U36289 ( .A(n17518), .B(n51401), .Z(n17519) );
  NAND U36290 ( .A(n51400), .B(n17519), .Z(n17520) );
  NANDN U36291 ( .A(n57754), .B(n17520), .Z(n17521) );
  AND U36292 ( .A(n57755), .B(n17521), .Z(n17522) );
  OR U36293 ( .A(n57756), .B(n17522), .Z(n17523) );
  NAND U36294 ( .A(n17524), .B(n17523), .Z(n17526) );
  NANDN U36295 ( .A(y[5372]), .B(x[5372]), .Z(n17525) );
  NANDN U36296 ( .A(y[5373]), .B(x[5373]), .Z(n24194) );
  AND U36297 ( .A(n17525), .B(n24194), .Z(n57760) );
  AND U36298 ( .A(n17526), .B(n57760), .Z(n17527) );
  NOR U36299 ( .A(n51398), .B(n17527), .Z(n17528) );
  NAND U36300 ( .A(n24195), .B(n17528), .Z(n17529) );
  NANDN U36301 ( .A(n57761), .B(n17529), .Z(n17530) );
  AND U36302 ( .A(n24193), .B(n17530), .Z(n17531) );
  NAND U36303 ( .A(n57763), .B(n17531), .Z(n17532) );
  NAND U36304 ( .A(n51397), .B(n17532), .Z(n17533) );
  NANDN U36305 ( .A(n57764), .B(n17533), .Z(n17534) );
  NAND U36306 ( .A(n57765), .B(n17534), .Z(n17535) );
  AND U36307 ( .A(n43786), .B(n17535), .Z(n17536) );
  NAND U36308 ( .A(n51395), .B(n17536), .Z(n17537) );
  NANDN U36309 ( .A(n57766), .B(n17537), .Z(n17538) );
  AND U36310 ( .A(n24187), .B(n17538), .Z(n17539) );
  NAND U36311 ( .A(n57770), .B(n17539), .Z(n17540) );
  NANDN U36312 ( .A(n57772), .B(n17540), .Z(n17541) );
  AND U36313 ( .A(n43796), .B(n17541), .Z(n17542) );
  NANDN U36314 ( .A(x[5383]), .B(y[5383]), .Z(n57773) );
  AND U36315 ( .A(n17542), .B(n57773), .Z(n17544) );
  NANDN U36316 ( .A(y[5384]), .B(x[5384]), .Z(n17543) );
  NANDN U36317 ( .A(y[5385]), .B(x[5385]), .Z(n24183) );
  NAND U36318 ( .A(n17543), .B(n24183), .Z(n51394) );
  OR U36319 ( .A(n17544), .B(n51394), .Z(n17545) );
  NAND U36320 ( .A(n57775), .B(n17545), .Z(n17546) );
  AND U36321 ( .A(n57776), .B(n17546), .Z(n17547) );
  ANDN U36322 ( .B(n57778), .A(n17547), .Z(n17548) );
  NAND U36323 ( .A(n43807), .B(n17548), .Z(n17549) );
  NANDN U36324 ( .A(n57779), .B(n17549), .Z(n17550) );
  AND U36325 ( .A(n24182), .B(n17550), .Z(n17551) );
  ANDN U36326 ( .B(y[5389]), .A(x[5389]), .Z(n57780) );
  ANDN U36327 ( .B(n17551), .A(n57780), .Z(n17553) );
  NANDN U36328 ( .A(y[5390]), .B(x[5390]), .Z(n17552) );
  NANDN U36329 ( .A(y[5391]), .B(x[5391]), .Z(n43817) );
  AND U36330 ( .A(n17552), .B(n43817), .Z(n57782) );
  NANDN U36331 ( .A(n17553), .B(n57782), .Z(n17554) );
  NAND U36332 ( .A(n43818), .B(n17554), .Z(n17555) );
  ANDN U36333 ( .B(y[5391]), .A(x[5391]), .Z(n43814) );
  OR U36334 ( .A(n17555), .B(n43814), .Z(n17556) );
  NAND U36335 ( .A(n57785), .B(n17556), .Z(n17557) );
  NANDN U36336 ( .A(n51391), .B(n17557), .Z(n17558) );
  XNOR U36337 ( .A(x[5394]), .B(y[5394]), .Z(n24180) );
  NANDN U36338 ( .A(n17558), .B(n24180), .Z(n17559) );
  AND U36339 ( .A(n57787), .B(n17559), .Z(n17560) );
  ANDN U36340 ( .B(n57789), .A(n17560), .Z(n17561) );
  NAND U36341 ( .A(n24178), .B(n17561), .Z(n17562) );
  NANDN U36342 ( .A(n57790), .B(n17562), .Z(n17563) );
  AND U36343 ( .A(n24176), .B(n17563), .Z(n17564) );
  NANDN U36344 ( .A(x[5397]), .B(y[5397]), .Z(n57791) );
  AND U36345 ( .A(n17564), .B(n57791), .Z(n17566) );
  NANDN U36346 ( .A(y[5398]), .B(x[5398]), .Z(n17565) );
  NANDN U36347 ( .A(y[5399]), .B(x[5399]), .Z(n24173) );
  NAND U36348 ( .A(n17565), .B(n24173), .Z(n57793) );
  OR U36349 ( .A(n17566), .B(n57793), .Z(n17567) );
  AND U36350 ( .A(n24174), .B(n17567), .Z(n17568) );
  NANDN U36351 ( .A(x[5399]), .B(y[5399]), .Z(n57794) );
  AND U36352 ( .A(n17568), .B(n57794), .Z(n17570) );
  NANDN U36353 ( .A(y[5400]), .B(x[5400]), .Z(n17569) );
  NANDN U36354 ( .A(y[5401]), .B(x[5401]), .Z(n24171) );
  NAND U36355 ( .A(n17569), .B(n24171), .Z(n57796) );
  OR U36356 ( .A(n17570), .B(n57796), .Z(n17571) );
  AND U36357 ( .A(n57797), .B(n17571), .Z(n17572) );
  NANDN U36358 ( .A(y[5402]), .B(x[5402]), .Z(n24170) );
  NANDN U36359 ( .A(y[5403]), .B(x[5403]), .Z(n43843) );
  NAND U36360 ( .A(n24170), .B(n43843), .Z(n57798) );
  OR U36361 ( .A(n17572), .B(n57798), .Z(n17573) );
  NAND U36362 ( .A(n17574), .B(n17573), .Z(n17575) );
  NANDN U36363 ( .A(n57801), .B(n17575), .Z(n17576) );
  AND U36364 ( .A(n24168), .B(n17576), .Z(n17577) );
  ANDN U36365 ( .B(y[5405]), .A(x[5405]), .Z(n57802) );
  ANDN U36366 ( .B(n17577), .A(n57802), .Z(n17579) );
  NANDN U36367 ( .A(y[5406]), .B(x[5406]), .Z(n17578) );
  NANDN U36368 ( .A(y[5407]), .B(x[5407]), .Z(n43854) );
  AND U36369 ( .A(n17578), .B(n43854), .Z(n57805) );
  NANDN U36370 ( .A(n17579), .B(n57805), .Z(n17580) );
  NAND U36371 ( .A(n43855), .B(n17580), .Z(n17581) );
  ANDN U36372 ( .B(y[5407]), .A(x[5407]), .Z(n43851) );
  OR U36373 ( .A(n17581), .B(n43851), .Z(n17582) );
  NAND U36374 ( .A(n57808), .B(n17582), .Z(n17584) );
  ANDN U36375 ( .B(y[5409]), .A(x[5409]), .Z(n51389) );
  XNOR U36376 ( .A(x[5410]), .B(y[5410]), .Z(n24166) );
  NANDN U36377 ( .A(n51389), .B(n24166), .Z(n17583) );
  ANDN U36378 ( .B(n17584), .A(n17583), .Z(n17586) );
  NANDN U36379 ( .A(y[5410]), .B(x[5410]), .Z(n17585) );
  NANDN U36380 ( .A(y[5411]), .B(x[5411]), .Z(n43864) );
  NAND U36381 ( .A(n17585), .B(n43864), .Z(n57809) );
  OR U36382 ( .A(n17586), .B(n57809), .Z(n17587) );
  NAND U36383 ( .A(n17588), .B(n17587), .Z(n17589) );
  NANDN U36384 ( .A(n57812), .B(n17589), .Z(n17590) );
  AND U36385 ( .A(n24164), .B(n17590), .Z(n17591) );
  NANDN U36386 ( .A(n57813), .B(n17591), .Z(n17592) );
  NANDN U36387 ( .A(n51388), .B(n17592), .Z(n17593) );
  AND U36388 ( .A(n43875), .B(n17593), .Z(n17594) );
  NANDN U36389 ( .A(x[5415]), .B(y[5415]), .Z(n57817) );
  AND U36390 ( .A(n17594), .B(n57817), .Z(n17595) );
  OR U36391 ( .A(n57820), .B(n17595), .Z(n17596) );
  NAND U36392 ( .A(n17597), .B(n17596), .Z(n17598) );
  AND U36393 ( .A(n57821), .B(n17598), .Z(n17599) );
  ANDN U36394 ( .B(n57823), .A(n17599), .Z(n17600) );
  NAND U36395 ( .A(n43885), .B(n17600), .Z(n17601) );
  NANDN U36396 ( .A(n57824), .B(n17601), .Z(n17602) );
  AND U36397 ( .A(n24160), .B(n17602), .Z(n17603) );
  NANDN U36398 ( .A(n57825), .B(n17603), .Z(n17604) );
  NANDN U36399 ( .A(n51385), .B(n17604), .Z(n17605) );
  XOR U36400 ( .A(x[5424]), .B(y[5424]), .Z(n43895) );
  ANDN U36401 ( .B(n17605), .A(n43895), .Z(n17606) );
  NANDN U36402 ( .A(x[5423]), .B(y[5423]), .Z(n57827) );
  AND U36403 ( .A(n17606), .B(n57827), .Z(n17607) );
  OR U36404 ( .A(n57829), .B(n17607), .Z(n17608) );
  NAND U36405 ( .A(n17609), .B(n17608), .Z(n17610) );
  AND U36406 ( .A(n57832), .B(n17610), .Z(n17611) );
  NOR U36407 ( .A(n43902), .B(n17611), .Z(n17612) );
  NAND U36408 ( .A(n24156), .B(n17612), .Z(n17613) );
  NANDN U36409 ( .A(n57835), .B(n17613), .Z(n17614) );
  AND U36410 ( .A(n24154), .B(n17614), .Z(n17615) );
  NANDN U36411 ( .A(x[5429]), .B(y[5429]), .Z(n57836) );
  NAND U36412 ( .A(n17615), .B(n57836), .Z(n17616) );
  NANDN U36413 ( .A(n57838), .B(n17616), .Z(n17617) );
  AND U36414 ( .A(n43914), .B(n17617), .Z(n17618) );
  NANDN U36415 ( .A(x[5431]), .B(y[5431]), .Z(n57839) );
  AND U36416 ( .A(n17618), .B(n57839), .Z(n17619) );
  OR U36417 ( .A(n57841), .B(n17619), .Z(n17620) );
  NAND U36418 ( .A(n17621), .B(n17620), .Z(n17622) );
  AND U36419 ( .A(n57842), .B(n17622), .Z(n17623) );
  ANDN U36420 ( .B(n57844), .A(n17623), .Z(n17624) );
  NAND U36421 ( .A(n43924), .B(n17624), .Z(n17625) );
  NANDN U36422 ( .A(n57845), .B(n17625), .Z(n17626) );
  AND U36423 ( .A(n24150), .B(n17626), .Z(n17627) );
  NANDN U36424 ( .A(n57846), .B(n17627), .Z(n17628) );
  NANDN U36425 ( .A(n57848), .B(n17628), .Z(n17629) );
  AND U36426 ( .A(n43934), .B(n17629), .Z(n17630) );
  NANDN U36427 ( .A(x[5439]), .B(y[5439]), .Z(n57850) );
  AND U36428 ( .A(n17630), .B(n57850), .Z(n17631) );
  OR U36429 ( .A(n57852), .B(n17631), .Z(n17632) );
  NAND U36430 ( .A(n17633), .B(n17632), .Z(n17634) );
  AND U36431 ( .A(n57853), .B(n17634), .Z(n17635) );
  ANDN U36432 ( .B(n57855), .A(n17635), .Z(n17636) );
  NAND U36433 ( .A(n43944), .B(n17636), .Z(n17637) );
  NANDN U36434 ( .A(n57856), .B(n17637), .Z(n17638) );
  AND U36435 ( .A(n24146), .B(n17638), .Z(n17639) );
  NANDN U36436 ( .A(n57857), .B(n17639), .Z(n17640) );
  NANDN U36437 ( .A(n57859), .B(n17640), .Z(n17641) );
  AND U36438 ( .A(n43954), .B(n17641), .Z(n17642) );
  NANDN U36439 ( .A(x[5447]), .B(y[5447]), .Z(n57860) );
  AND U36440 ( .A(n17642), .B(n57860), .Z(n17643) );
  OR U36441 ( .A(n57862), .B(n17643), .Z(n17644) );
  NAND U36442 ( .A(n17645), .B(n17644), .Z(n17646) );
  NAND U36443 ( .A(n57864), .B(n17646), .Z(n17647) );
  AND U36444 ( .A(n24142), .B(n17647), .Z(n17648) );
  NAND U36445 ( .A(n57865), .B(n17648), .Z(n17649) );
  NANDN U36446 ( .A(n57868), .B(n17649), .Z(n17650) );
  AND U36447 ( .A(n24140), .B(n17650), .Z(n17651) );
  NANDN U36448 ( .A(x[5453]), .B(y[5453]), .Z(n57869) );
  NAND U36449 ( .A(n17651), .B(n57869), .Z(n17652) );
  NANDN U36450 ( .A(n57871), .B(n17652), .Z(n17653) );
  AND U36451 ( .A(n43972), .B(n17653), .Z(n17654) );
  NANDN U36452 ( .A(x[5455]), .B(y[5455]), .Z(n57872) );
  AND U36453 ( .A(n17654), .B(n57872), .Z(n17655) );
  OR U36454 ( .A(n57874), .B(n17655), .Z(n17656) );
  NAND U36455 ( .A(n17657), .B(n17656), .Z(n17658) );
  AND U36456 ( .A(n57875), .B(n17658), .Z(n17659) );
  ANDN U36457 ( .B(n57877), .A(n17659), .Z(n17660) );
  NAND U36458 ( .A(n43982), .B(n17660), .Z(n17661) );
  NANDN U36459 ( .A(n57878), .B(n17661), .Z(n17662) );
  AND U36460 ( .A(n57879), .B(n17662), .Z(n17664) );
  NANDN U36461 ( .A(y[5462]), .B(x[5462]), .Z(n17663) );
  NANDN U36462 ( .A(y[5463]), .B(x[5463]), .Z(n24131) );
  NAND U36463 ( .A(n17663), .B(n24131), .Z(n57880) );
  OR U36464 ( .A(n17664), .B(n57880), .Z(n17665) );
  AND U36465 ( .A(n24132), .B(n17665), .Z(n17666) );
  NANDN U36466 ( .A(x[5463]), .B(y[5463]), .Z(n51373) );
  AND U36467 ( .A(n17666), .B(n51373), .Z(n17668) );
  NANDN U36468 ( .A(y[5464]), .B(x[5464]), .Z(n17667) );
  NANDN U36469 ( .A(y[5465]), .B(x[5465]), .Z(n24128) );
  NAND U36470 ( .A(n17667), .B(n24128), .Z(n57882) );
  OR U36471 ( .A(n17668), .B(n57882), .Z(n17669) );
  NAND U36472 ( .A(n57883), .B(n17669), .Z(n17671) );
  NANDN U36473 ( .A(y[5466]), .B(x[5466]), .Z(n17670) );
  NANDN U36474 ( .A(y[5467]), .B(x[5467]), .Z(n44001) );
  AND U36475 ( .A(n17670), .B(n44001), .Z(n51372) );
  AND U36476 ( .A(n17671), .B(n51372), .Z(n17672) );
  NOR U36477 ( .A(n43997), .B(n17672), .Z(n17673) );
  NAND U36478 ( .A(n44002), .B(n17673), .Z(n17674) );
  NANDN U36479 ( .A(n57886), .B(n17674), .Z(n17675) );
  AND U36480 ( .A(n24126), .B(n17675), .Z(n17676) );
  NANDN U36481 ( .A(x[5469]), .B(y[5469]), .Z(n24127) );
  AND U36482 ( .A(n17676), .B(n24127), .Z(n17678) );
  NANDN U36483 ( .A(y[5470]), .B(x[5470]), .Z(n17677) );
  NANDN U36484 ( .A(y[5471]), .B(x[5471]), .Z(n44011) );
  NAND U36485 ( .A(n17677), .B(n44011), .Z(n57887) );
  OR U36486 ( .A(n17678), .B(n57887), .Z(n17679) );
  AND U36487 ( .A(n44012), .B(n17679), .Z(n17680) );
  NANDN U36488 ( .A(x[5471]), .B(y[5471]), .Z(n57888) );
  AND U36489 ( .A(n17680), .B(n57888), .Z(n17682) );
  NANDN U36490 ( .A(y[5472]), .B(x[5472]), .Z(n17681) );
  NANDN U36491 ( .A(y[5473]), .B(x[5473]), .Z(n24123) );
  NAND U36492 ( .A(n17681), .B(n24123), .Z(n57890) );
  OR U36493 ( .A(n17682), .B(n57890), .Z(n17683) );
  AND U36494 ( .A(n57891), .B(n17683), .Z(n17684) );
  NANDN U36495 ( .A(y[5474]), .B(x[5474]), .Z(n24122) );
  NANDN U36496 ( .A(y[5475]), .B(x[5475]), .Z(n24119) );
  NAND U36497 ( .A(n24122), .B(n24119), .Z(n51369) );
  OR U36498 ( .A(n17684), .B(n51369), .Z(n17685) );
  NAND U36499 ( .A(n51368), .B(n17685), .Z(n17686) );
  NANDN U36500 ( .A(n57894), .B(n17686), .Z(n17687) );
  AND U36501 ( .A(n24117), .B(n17687), .Z(n17688) );
  ANDN U36502 ( .B(y[5477]), .A(x[5477]), .Z(n57896) );
  ANDN U36503 ( .B(n17688), .A(n57896), .Z(n17690) );
  NANDN U36504 ( .A(y[5478]), .B(x[5478]), .Z(n17689) );
  NANDN U36505 ( .A(y[5479]), .B(x[5479]), .Z(n24114) );
  NAND U36506 ( .A(n17689), .B(n24114), .Z(n57897) );
  OR U36507 ( .A(n17690), .B(n57897), .Z(n17691) );
  NANDN U36508 ( .A(x[5479]), .B(y[5479]), .Z(n24115) );
  NANDN U36509 ( .A(x[5480]), .B(y[5480]), .Z(n24112) );
  AND U36510 ( .A(n24115), .B(n24112), .Z(n57898) );
  AND U36511 ( .A(n17691), .B(n57898), .Z(n17692) );
  NANDN U36512 ( .A(y[5480]), .B(x[5480]), .Z(n24113) );
  NANDN U36513 ( .A(y[5481]), .B(x[5481]), .Z(n24110) );
  NAND U36514 ( .A(n24113), .B(n24110), .Z(n51367) );
  OR U36515 ( .A(n17692), .B(n51367), .Z(n17693) );
  NAND U36516 ( .A(n51366), .B(n17693), .Z(n17694) );
  NANDN U36517 ( .A(n57899), .B(n17694), .Z(n17695) );
  AND U36518 ( .A(n57900), .B(n17695), .Z(n17696) );
  NANDN U36519 ( .A(y[5484]), .B(x[5484]), .Z(n24106) );
  NANDN U36520 ( .A(y[5485]), .B(x[5485]), .Z(n24102) );
  NAND U36521 ( .A(n24106), .B(n24102), .Z(n57901) );
  OR U36522 ( .A(n17696), .B(n57901), .Z(n17697) );
  AND U36523 ( .A(n17698), .B(n17697), .Z(n17699) );
  OR U36524 ( .A(n57904), .B(n17699), .Z(n17700) );
  NAND U36525 ( .A(n57906), .B(n17700), .Z(n17701) );
  NANDN U36526 ( .A(n57907), .B(n17701), .Z(n17702) );
  AND U36527 ( .A(n24099), .B(n17702), .Z(n17703) );
  NAND U36528 ( .A(n57909), .B(n17703), .Z(n17704) );
  NAND U36529 ( .A(n51365), .B(n17704), .Z(n17705) );
  ANDN U36530 ( .B(y[5491]), .A(x[5491]), .Z(n44054) );
  ANDN U36531 ( .B(n17705), .A(n44054), .Z(n17706) );
  NAND U36532 ( .A(n44058), .B(n17706), .Z(n17708) );
  NANDN U36533 ( .A(y[5492]), .B(x[5492]), .Z(n17707) );
  NANDN U36534 ( .A(y[5493]), .B(x[5493]), .Z(n24096) );
  AND U36535 ( .A(n17707), .B(n24096), .Z(n57912) );
  AND U36536 ( .A(n17708), .B(n57912), .Z(n17709) );
  ANDN U36537 ( .B(n17710), .A(n17709), .Z(n17711) );
  OR U36538 ( .A(n57915), .B(n17711), .Z(n17712) );
  NAND U36539 ( .A(n57916), .B(n17712), .Z(n17713) );
  NANDN U36540 ( .A(n57917), .B(n17713), .Z(n17714) );
  AND U36541 ( .A(n24092), .B(n17714), .Z(n17715) );
  NANDN U36542 ( .A(x[5497]), .B(y[5497]), .Z(n57919) );
  AND U36543 ( .A(n17715), .B(n57919), .Z(n17716) );
  OR U36544 ( .A(n57922), .B(n17716), .Z(n17717) );
  AND U36545 ( .A(n17718), .B(n17717), .Z(n17720) );
  NANDN U36546 ( .A(y[5500]), .B(x[5500]), .Z(n17719) );
  NANDN U36547 ( .A(y[5501]), .B(x[5501]), .Z(n24086) );
  NAND U36548 ( .A(n17719), .B(n24086), .Z(n51363) );
  OR U36549 ( .A(n17720), .B(n51363), .Z(n17721) );
  NAND U36550 ( .A(n51362), .B(n17721), .Z(n17722) );
  NANDN U36551 ( .A(n57924), .B(n17722), .Z(n17723) );
  AND U36552 ( .A(n44086), .B(n17723), .Z(n17724) );
  NAND U36553 ( .A(n57926), .B(n17724), .Z(n17725) );
  NAND U36554 ( .A(n51361), .B(n17725), .Z(n17726) );
  NAND U36555 ( .A(n24085), .B(n17726), .Z(n17727) );
  ANDN U36556 ( .B(y[5505]), .A(x[5505]), .Z(n57927) );
  OR U36557 ( .A(n17727), .B(n57927), .Z(n17728) );
  NAND U36558 ( .A(n57929), .B(n17728), .Z(n17730) );
  XNOR U36559 ( .A(x[5508]), .B(y[5508]), .Z(n44096) );
  NANDN U36560 ( .A(x[5507]), .B(y[5507]), .Z(n57931) );
  NAND U36561 ( .A(n44096), .B(n57931), .Z(n17729) );
  ANDN U36562 ( .B(n17730), .A(n17729), .Z(n17731) );
  OR U36563 ( .A(n57933), .B(n17731), .Z(n17732) );
  NAND U36564 ( .A(n57934), .B(n17732), .Z(n17733) );
  NANDN U36565 ( .A(n57935), .B(n17733), .Z(n17734) );
  NAND U36566 ( .A(n24079), .B(n17734), .Z(n17735) );
  ANDN U36567 ( .B(y[5511]), .A(x[5511]), .Z(n24080) );
  OR U36568 ( .A(n17735), .B(n24080), .Z(n17736) );
  NAND U36569 ( .A(n57936), .B(n17736), .Z(n17738) );
  XNOR U36570 ( .A(x[5514]), .B(y[5514]), .Z(n24077) );
  NANDN U36571 ( .A(x[5513]), .B(y[5513]), .Z(n57937) );
  NAND U36572 ( .A(n24077), .B(n57937), .Z(n17737) );
  ANDN U36573 ( .B(n17738), .A(n17737), .Z(n17740) );
  NANDN U36574 ( .A(y[5514]), .B(x[5514]), .Z(n17739) );
  NANDN U36575 ( .A(y[5515]), .B(x[5515]), .Z(n24075) );
  NAND U36576 ( .A(n17739), .B(n24075), .Z(n51357) );
  OR U36577 ( .A(n17740), .B(n51357), .Z(n17741) );
  NAND U36578 ( .A(n51356), .B(n17741), .Z(n17742) );
  NANDN U36579 ( .A(n57938), .B(n17742), .Z(n17743) );
  NANDN U36580 ( .A(x[5517]), .B(y[5517]), .Z(n57939) );
  AND U36581 ( .A(n17743), .B(n57939), .Z(n17744) );
  NANDN U36582 ( .A(x[5518]), .B(y[5518]), .Z(n24071) );
  AND U36583 ( .A(n17744), .B(n24071), .Z(n17745) );
  NANDN U36584 ( .A(y[5518]), .B(x[5518]), .Z(n24072) );
  NANDN U36585 ( .A(y[5519]), .B(x[5519]), .Z(n57944) );
  AND U36586 ( .A(n24072), .B(n57944), .Z(n57941) );
  NANDN U36587 ( .A(n17745), .B(n57941), .Z(n17746) );
  NANDN U36588 ( .A(x[5520]), .B(y[5520]), .Z(n57942) );
  AND U36589 ( .A(n17746), .B(n57942), .Z(n17747) );
  NANDN U36590 ( .A(x[5519]), .B(y[5519]), .Z(n24070) );
  AND U36591 ( .A(n17747), .B(n24070), .Z(n17748) );
  OR U36592 ( .A(n57947), .B(n17748), .Z(n17749) );
  NAND U36593 ( .A(n17750), .B(n17749), .Z(n17752) );
  NANDN U36594 ( .A(y[5522]), .B(x[5522]), .Z(n17751) );
  NANDN U36595 ( .A(y[5523]), .B(x[5523]), .Z(n44132) );
  AND U36596 ( .A(n17751), .B(n44132), .Z(n57950) );
  AND U36597 ( .A(n17752), .B(n57950), .Z(n17753) );
  NOR U36598 ( .A(n44129), .B(n17753), .Z(n17754) );
  NAND U36599 ( .A(n44133), .B(n17754), .Z(n17755) );
  NANDN U36600 ( .A(n57951), .B(n17755), .Z(n17756) );
  AND U36601 ( .A(n24066), .B(n17756), .Z(n17757) );
  NANDN U36602 ( .A(n57953), .B(n17757), .Z(n17758) );
  NAND U36603 ( .A(n51353), .B(n17758), .Z(n17759) );
  NANDN U36604 ( .A(n57954), .B(n17759), .Z(n17760) );
  AND U36605 ( .A(n57955), .B(n17760), .Z(n17761) );
  ANDN U36606 ( .B(n17762), .A(n17761), .Z(n17763) );
  ANDN U36607 ( .B(n57957), .A(n17763), .Z(n17764) );
  ANDN U36608 ( .B(n57959), .A(n17764), .Z(n17765) );
  NAND U36609 ( .A(n24059), .B(n17765), .Z(n17766) );
  NANDN U36610 ( .A(n57960), .B(n17766), .Z(n17767) );
  AND U36611 ( .A(n24057), .B(n17767), .Z(n17768) );
  NANDN U36612 ( .A(x[5533]), .B(y[5533]), .Z(n57961) );
  AND U36613 ( .A(n17768), .B(n57961), .Z(n17770) );
  NANDN U36614 ( .A(y[5534]), .B(x[5534]), .Z(n17769) );
  NANDN U36615 ( .A(y[5535]), .B(x[5535]), .Z(n44159) );
  NAND U36616 ( .A(n17769), .B(n44159), .Z(n57963) );
  OR U36617 ( .A(n17770), .B(n57963), .Z(n17771) );
  AND U36618 ( .A(n44160), .B(n17771), .Z(n17772) );
  NANDN U36619 ( .A(x[5535]), .B(y[5535]), .Z(n57964) );
  AND U36620 ( .A(n17772), .B(n57964), .Z(n17774) );
  NANDN U36621 ( .A(y[5536]), .B(x[5536]), .Z(n17773) );
  NANDN U36622 ( .A(y[5537]), .B(x[5537]), .Z(n24054) );
  NAND U36623 ( .A(n17773), .B(n24054), .Z(n57966) );
  OR U36624 ( .A(n17774), .B(n57966), .Z(n17775) );
  AND U36625 ( .A(n57967), .B(n17775), .Z(n17776) );
  OR U36626 ( .A(n57968), .B(n17776), .Z(n17777) );
  NAND U36627 ( .A(n57969), .B(n17777), .Z(n17778) );
  NANDN U36628 ( .A(n57971), .B(n17778), .Z(n17779) );
  NAND U36629 ( .A(n24048), .B(n17779), .Z(n17780) );
  ANDN U36630 ( .B(y[5541]), .A(x[5541]), .Z(n57972) );
  OR U36631 ( .A(n17780), .B(n57972), .Z(n17781) );
  NAND U36632 ( .A(n57974), .B(n17781), .Z(n17782) );
  NANDN U36633 ( .A(n57975), .B(n17782), .Z(n17783) );
  AND U36634 ( .A(n57976), .B(n17783), .Z(n17784) );
  ANDN U36635 ( .B(n51350), .A(n17784), .Z(n17785) );
  NAND U36636 ( .A(n24042), .B(n17785), .Z(n17786) );
  NANDN U36637 ( .A(n51348), .B(n17786), .Z(n17787) );
  AND U36638 ( .A(n44188), .B(n17787), .Z(n17788) );
  NANDN U36639 ( .A(n44184), .B(n17788), .Z(n17789) );
  NAND U36640 ( .A(n57979), .B(n17789), .Z(n17790) );
  AND U36641 ( .A(n24040), .B(n17790), .Z(n17791) );
  ANDN U36642 ( .B(y[5549]), .A(x[5549]), .Z(n57980) );
  ANDN U36643 ( .B(n17791), .A(n57980), .Z(n17793) );
  NANDN U36644 ( .A(y[5550]), .B(x[5550]), .Z(n17792) );
  NANDN U36645 ( .A(y[5551]), .B(x[5551]), .Z(n44198) );
  AND U36646 ( .A(n17792), .B(n44198), .Z(n57983) );
  NANDN U36647 ( .A(n17793), .B(n57983), .Z(n17794) );
  NAND U36648 ( .A(n17795), .B(n17794), .Z(n17796) );
  AND U36649 ( .A(n57984), .B(n17796), .Z(n17797) );
  NOR U36650 ( .A(n57986), .B(n17797), .Z(n17798) );
  NAND U36651 ( .A(n24038), .B(n17798), .Z(n17799) );
  NANDN U36652 ( .A(n57987), .B(n17799), .Z(n17800) );
  AND U36653 ( .A(n44209), .B(n17800), .Z(n17801) );
  NANDN U36654 ( .A(x[5555]), .B(y[5555]), .Z(n57988) );
  AND U36655 ( .A(n17801), .B(n57988), .Z(n17803) );
  NANDN U36656 ( .A(y[5556]), .B(x[5556]), .Z(n17802) );
  NANDN U36657 ( .A(y[5557]), .B(x[5557]), .Z(n24035) );
  NAND U36658 ( .A(n17802), .B(n24035), .Z(n57990) );
  OR U36659 ( .A(n17803), .B(n57990), .Z(n17804) );
  AND U36660 ( .A(n24036), .B(n17804), .Z(n17805) );
  ANDN U36661 ( .B(y[5557]), .A(x[5557]), .Z(n57991) );
  ANDN U36662 ( .B(n17805), .A(n57991), .Z(n17807) );
  NANDN U36663 ( .A(y[5558]), .B(x[5558]), .Z(n17806) );
  NANDN U36664 ( .A(y[5559]), .B(x[5559]), .Z(n44219) );
  AND U36665 ( .A(n17806), .B(n44219), .Z(n57993) );
  NANDN U36666 ( .A(n17807), .B(n57993), .Z(n17808) );
  NAND U36667 ( .A(n17809), .B(n17808), .Z(n17810) );
  AND U36668 ( .A(n57995), .B(n17810), .Z(n17811) );
  NOR U36669 ( .A(n57997), .B(n17811), .Z(n17812) );
  NAND U36670 ( .A(n24034), .B(n17812), .Z(n17813) );
  NANDN U36671 ( .A(n57999), .B(n17813), .Z(n17814) );
  AND U36672 ( .A(n44230), .B(n17814), .Z(n17815) );
  NANDN U36673 ( .A(x[5563]), .B(y[5563]), .Z(n58000) );
  AND U36674 ( .A(n17815), .B(n58000), .Z(n17817) );
  NANDN U36675 ( .A(y[5564]), .B(x[5564]), .Z(n17816) );
  NANDN U36676 ( .A(y[5565]), .B(x[5565]), .Z(n24031) );
  NAND U36677 ( .A(n17816), .B(n24031), .Z(n58002) );
  OR U36678 ( .A(n17817), .B(n58002), .Z(n17818) );
  AND U36679 ( .A(n24032), .B(n17818), .Z(n17819) );
  ANDN U36680 ( .B(y[5565]), .A(x[5565]), .Z(n58003) );
  ANDN U36681 ( .B(n17819), .A(n58003), .Z(n17821) );
  NANDN U36682 ( .A(y[5566]), .B(x[5566]), .Z(n17820) );
  NANDN U36683 ( .A(y[5567]), .B(x[5567]), .Z(n24030) );
  NAND U36684 ( .A(n17820), .B(n24030), .Z(n58005) );
  OR U36685 ( .A(n17821), .B(n58005), .Z(n17822) );
  AND U36686 ( .A(n58006), .B(n17822), .Z(n17823) );
  OR U36687 ( .A(n58007), .B(n17823), .Z(n17824) );
  NAND U36688 ( .A(n58008), .B(n17824), .Z(n17825) );
  NANDN U36689 ( .A(n58009), .B(n17825), .Z(n17826) );
  AND U36690 ( .A(n58010), .B(n17826), .Z(n17828) );
  NANDN U36691 ( .A(y[5572]), .B(x[5572]), .Z(n17827) );
  NANDN U36692 ( .A(y[5573]), .B(x[5573]), .Z(n24019) );
  AND U36693 ( .A(n17827), .B(n24019), .Z(n58011) );
  NANDN U36694 ( .A(n17828), .B(n58011), .Z(n17829) );
  NANDN U36695 ( .A(n58012), .B(n17829), .Z(n17830) );
  AND U36696 ( .A(n58013), .B(n17830), .Z(n17831) );
  OR U36697 ( .A(n58015), .B(n17831), .Z(n17832) );
  NAND U36698 ( .A(n58016), .B(n17832), .Z(n17833) );
  NANDN U36699 ( .A(n58017), .B(n17833), .Z(n17834) );
  NAND U36700 ( .A(n58018), .B(n17834), .Z(n17835) );
  AND U36701 ( .A(n44274), .B(n17835), .Z(n17836) );
  NAND U36702 ( .A(n58020), .B(n17836), .Z(n17837) );
  NANDN U36703 ( .A(n58021), .B(n17837), .Z(n17838) );
  AND U36704 ( .A(n58022), .B(n17838), .Z(n17840) );
  NANDN U36705 ( .A(y[5582]), .B(x[5582]), .Z(n17839) );
  NANDN U36706 ( .A(y[5583]), .B(x[5583]), .Z(n24013) );
  AND U36707 ( .A(n17839), .B(n24013), .Z(n58023) );
  NANDN U36708 ( .A(n17840), .B(n58023), .Z(n17841) );
  NAND U36709 ( .A(n17842), .B(n17841), .Z(n17843) );
  AND U36710 ( .A(n58024), .B(n17843), .Z(n17844) );
  ANDN U36711 ( .B(n17845), .A(n17844), .Z(n17847) );
  NANDN U36712 ( .A(y[5586]), .B(x[5586]), .Z(n17846) );
  NANDN U36713 ( .A(y[5587]), .B(x[5587]), .Z(n24009) );
  NAND U36714 ( .A(n17846), .B(n24009), .Z(n58027) );
  OR U36715 ( .A(n17847), .B(n58027), .Z(n17848) );
  AND U36716 ( .A(n58028), .B(n17848), .Z(n17849) );
  NANDN U36717 ( .A(y[5588]), .B(x[5588]), .Z(n24008) );
  NANDN U36718 ( .A(y[5589]), .B(x[5589]), .Z(n24005) );
  AND U36719 ( .A(n24008), .B(n24005), .Z(n58029) );
  NANDN U36720 ( .A(n17849), .B(n58029), .Z(n17850) );
  AND U36721 ( .A(n24006), .B(n17850), .Z(n17851) );
  NANDN U36722 ( .A(x[5589]), .B(y[5589]), .Z(n51340) );
  NAND U36723 ( .A(n17851), .B(n51340), .Z(n17852) );
  NANDN U36724 ( .A(n58031), .B(n17852), .Z(n17853) );
  AND U36725 ( .A(n58032), .B(n17853), .Z(n17854) );
  OR U36726 ( .A(n58033), .B(n17854), .Z(n17855) );
  NAND U36727 ( .A(n58034), .B(n17855), .Z(n17856) );
  NANDN U36728 ( .A(n58035), .B(n17856), .Z(n17857) );
  AND U36729 ( .A(n58036), .B(n17857), .Z(n17859) );
  NANDN U36730 ( .A(y[5596]), .B(x[5596]), .Z(n17858) );
  NANDN U36731 ( .A(y[5597]), .B(x[5597]), .Z(n23993) );
  NAND U36732 ( .A(n17858), .B(n23993), .Z(n58037) );
  OR U36733 ( .A(n17859), .B(n58037), .Z(n17860) );
  AND U36734 ( .A(n17861), .B(n17860), .Z(n17862) );
  OR U36735 ( .A(n58040), .B(n17862), .Z(n17863) );
  NAND U36736 ( .A(n58041), .B(n17863), .Z(n17864) );
  NANDN U36737 ( .A(n58042), .B(n17864), .Z(n17865) );
  AND U36738 ( .A(n23988), .B(n17865), .Z(n17866) );
  NANDN U36739 ( .A(x[5601]), .B(y[5601]), .Z(n51338) );
  AND U36740 ( .A(n17866), .B(n51338), .Z(n17868) );
  NANDN U36741 ( .A(y[5602]), .B(x[5602]), .Z(n17867) );
  NANDN U36742 ( .A(y[5603]), .B(x[5603]), .Z(n23985) );
  AND U36743 ( .A(n17867), .B(n23985), .Z(n58044) );
  NANDN U36744 ( .A(n17868), .B(n58044), .Z(n17869) );
  AND U36745 ( .A(n23986), .B(n17869), .Z(n17870) );
  NANDN U36746 ( .A(x[5603]), .B(y[5603]), .Z(n58045) );
  AND U36747 ( .A(n17870), .B(n58045), .Z(n17872) );
  NANDN U36748 ( .A(y[5604]), .B(x[5604]), .Z(n17871) );
  NANDN U36749 ( .A(y[5605]), .B(x[5605]), .Z(n23984) );
  NAND U36750 ( .A(n17871), .B(n23984), .Z(n58048) );
  OR U36751 ( .A(n17872), .B(n58048), .Z(n17873) );
  AND U36752 ( .A(n58049), .B(n17873), .Z(n17874) );
  OR U36753 ( .A(n58050), .B(n17874), .Z(n17875) );
  NAND U36754 ( .A(n17876), .B(n17875), .Z(n17877) );
  NANDN U36755 ( .A(n58051), .B(n17877), .Z(n17878) );
  AND U36756 ( .A(n58052), .B(n17878), .Z(n17879) );
  NANDN U36757 ( .A(y[5610]), .B(x[5610]), .Z(n23978) );
  ANDN U36758 ( .B(x[5611]), .A(y[5611]), .Z(n44345) );
  ANDN U36759 ( .B(n23978), .A(n44345), .Z(n58053) );
  NANDN U36760 ( .A(n17879), .B(n58053), .Z(n17880) );
  NAND U36761 ( .A(n17881), .B(n17880), .Z(n17883) );
  NANDN U36762 ( .A(y[5612]), .B(x[5612]), .Z(n17882) );
  NANDN U36763 ( .A(y[5613]), .B(x[5613]), .Z(n23974) );
  AND U36764 ( .A(n17882), .B(n23974), .Z(n58056) );
  AND U36765 ( .A(n17883), .B(n58056), .Z(n17885) );
  XNOR U36766 ( .A(x[5614]), .B(y[5614]), .Z(n23975) );
  ANDN U36767 ( .B(y[5613]), .A(x[5613]), .Z(n44348) );
  ANDN U36768 ( .B(n23975), .A(n44348), .Z(n17884) );
  NANDN U36769 ( .A(n17885), .B(n17884), .Z(n17887) );
  NANDN U36770 ( .A(y[5614]), .B(x[5614]), .Z(n17886) );
  NANDN U36771 ( .A(y[5615]), .B(x[5615]), .Z(n23972) );
  AND U36772 ( .A(n17886), .B(n23972), .Z(n58057) );
  AND U36773 ( .A(n17887), .B(n58057), .Z(n17888) );
  XNOR U36774 ( .A(y[5616]), .B(x[5616]), .Z(n23973) );
  NANDN U36775 ( .A(x[5615]), .B(y[5615]), .Z(n44353) );
  NAND U36776 ( .A(n23973), .B(n44353), .Z(n51333) );
  OR U36777 ( .A(n17888), .B(n51333), .Z(n17889) );
  NAND U36778 ( .A(n51332), .B(n17889), .Z(n17890) );
  NANDN U36779 ( .A(n58060), .B(n17890), .Z(n17891) );
  NAND U36780 ( .A(n58061), .B(n17891), .Z(n17892) );
  AND U36781 ( .A(n23968), .B(n17892), .Z(n17893) );
  NAND U36782 ( .A(n51330), .B(n17893), .Z(n17894) );
  NANDN U36783 ( .A(n58062), .B(n17894), .Z(n17895) );
  AND U36784 ( .A(n58063), .B(n17895), .Z(n17896) );
  NANDN U36785 ( .A(y[5622]), .B(x[5622]), .Z(n23965) );
  NANDN U36786 ( .A(y[5623]), .B(x[5623]), .Z(n23962) );
  NAND U36787 ( .A(n23965), .B(n23962), .Z(n58064) );
  OR U36788 ( .A(n17896), .B(n58064), .Z(n17897) );
  AND U36789 ( .A(n23963), .B(n17897), .Z(n17898) );
  NANDN U36790 ( .A(x[5623]), .B(y[5623]), .Z(n58065) );
  AND U36791 ( .A(n17898), .B(n58065), .Z(n17900) );
  NANDN U36792 ( .A(y[5624]), .B(x[5624]), .Z(n17899) );
  NANDN U36793 ( .A(y[5625]), .B(x[5625]), .Z(n23960) );
  NAND U36794 ( .A(n17899), .B(n23960), .Z(n58067) );
  OR U36795 ( .A(n17900), .B(n58067), .Z(n17901) );
  NAND U36796 ( .A(n17902), .B(n17901), .Z(n17903) );
  AND U36797 ( .A(n58068), .B(n17903), .Z(n17904) );
  ANDN U36798 ( .B(n58070), .A(n17904), .Z(n17905) );
  NAND U36799 ( .A(n23959), .B(n17905), .Z(n17906) );
  NANDN U36800 ( .A(n58071), .B(n17906), .Z(n17907) );
  AND U36801 ( .A(n23957), .B(n17907), .Z(n17908) );
  NANDN U36802 ( .A(x[5629]), .B(y[5629]), .Z(n58073) );
  AND U36803 ( .A(n17908), .B(n58073), .Z(n17909) );
  OR U36804 ( .A(n58076), .B(n17909), .Z(n17910) );
  AND U36805 ( .A(n44393), .B(n17910), .Z(n17911) );
  NANDN U36806 ( .A(x[5631]), .B(y[5631]), .Z(n58077) );
  AND U36807 ( .A(n17911), .B(n58077), .Z(n17913) );
  NANDN U36808 ( .A(y[5632]), .B(x[5632]), .Z(n17912) );
  NANDN U36809 ( .A(y[5633]), .B(x[5633]), .Z(n23954) );
  AND U36810 ( .A(n17912), .B(n23954), .Z(n58079) );
  NANDN U36811 ( .A(n17913), .B(n58079), .Z(n17914) );
  NAND U36812 ( .A(n17915), .B(n17914), .Z(n17916) );
  AND U36813 ( .A(n58080), .B(n17916), .Z(n17917) );
  ANDN U36814 ( .B(n58082), .A(n17917), .Z(n17918) );
  NAND U36815 ( .A(n23953), .B(n17918), .Z(n17919) );
  NANDN U36816 ( .A(n58083), .B(n17919), .Z(n17920) );
  AND U36817 ( .A(n23951), .B(n17920), .Z(n17921) );
  NANDN U36818 ( .A(x[5637]), .B(y[5637]), .Z(n58084) );
  AND U36819 ( .A(n17921), .B(n58084), .Z(n17923) );
  NANDN U36820 ( .A(y[5638]), .B(x[5638]), .Z(n17922) );
  NANDN U36821 ( .A(y[5639]), .B(x[5639]), .Z(n23948) );
  NAND U36822 ( .A(n17922), .B(n23948), .Z(n58086) );
  OR U36823 ( .A(n17923), .B(n58086), .Z(n17924) );
  AND U36824 ( .A(n23949), .B(n17924), .Z(n17925) );
  NANDN U36825 ( .A(x[5639]), .B(y[5639]), .Z(n58087) );
  AND U36826 ( .A(n17925), .B(n58087), .Z(n17927) );
  NANDN U36827 ( .A(y[5640]), .B(x[5640]), .Z(n17926) );
  NANDN U36828 ( .A(y[5641]), .B(x[5641]), .Z(n23946) );
  AND U36829 ( .A(n17926), .B(n23946), .Z(n58089) );
  NANDN U36830 ( .A(n17927), .B(n58089), .Z(n17928) );
  NAND U36831 ( .A(n17929), .B(n17928), .Z(n17930) );
  AND U36832 ( .A(n58092), .B(n17930), .Z(n17931) );
  ANDN U36833 ( .B(n58094), .A(n17931), .Z(n17932) );
  NAND U36834 ( .A(n23945), .B(n17932), .Z(n17933) );
  NANDN U36835 ( .A(n58095), .B(n17933), .Z(n17934) );
  AND U36836 ( .A(n23943), .B(n17934), .Z(n17935) );
  NANDN U36837 ( .A(x[5645]), .B(y[5645]), .Z(n58096) );
  AND U36838 ( .A(n17935), .B(n58096), .Z(n17937) );
  NANDN U36839 ( .A(y[5646]), .B(x[5646]), .Z(n17936) );
  NANDN U36840 ( .A(y[5647]), .B(x[5647]), .Z(n23939) );
  AND U36841 ( .A(n17936), .B(n23939), .Z(n58098) );
  NANDN U36842 ( .A(n17937), .B(n58098), .Z(n17938) );
  NAND U36843 ( .A(n23940), .B(n17938), .Z(n17939) );
  ANDN U36844 ( .B(y[5647]), .A(x[5647]), .Z(n23941) );
  OR U36845 ( .A(n17939), .B(n23941), .Z(n17940) );
  NAND U36846 ( .A(n58101), .B(n17940), .Z(n17942) );
  XNOR U36847 ( .A(x[5650]), .B(y[5650]), .Z(n23938) );
  NANDN U36848 ( .A(x[5649]), .B(y[5649]), .Z(n51322) );
  NAND U36849 ( .A(n23938), .B(n51322), .Z(n17941) );
  ANDN U36850 ( .B(n17942), .A(n17941), .Z(n17943) );
  OR U36851 ( .A(n58102), .B(n17943), .Z(n17944) );
  NAND U36852 ( .A(n58103), .B(n17944), .Z(n17945) );
  NANDN U36853 ( .A(n58104), .B(n17945), .Z(n17946) );
  AND U36854 ( .A(n23933), .B(n17946), .Z(n17947) );
  NANDN U36855 ( .A(x[5653]), .B(y[5653]), .Z(n58105) );
  AND U36856 ( .A(n17947), .B(n58105), .Z(n17949) );
  NANDN U36857 ( .A(y[5654]), .B(x[5654]), .Z(n17948) );
  NANDN U36858 ( .A(y[5655]), .B(x[5655]), .Z(n44446) );
  NAND U36859 ( .A(n17948), .B(n44446), .Z(n58107) );
  OR U36860 ( .A(n17949), .B(n58107), .Z(n17950) );
  XOR U36861 ( .A(x[5656]), .B(y[5656]), .Z(n44445) );
  ANDN U36862 ( .B(n17950), .A(n44445), .Z(n17951) );
  NANDN U36863 ( .A(x[5655]), .B(y[5655]), .Z(n51320) );
  AND U36864 ( .A(n17951), .B(n51320), .Z(n17953) );
  NANDN U36865 ( .A(y[5656]), .B(x[5656]), .Z(n17952) );
  NANDN U36866 ( .A(y[5657]), .B(x[5657]), .Z(n23930) );
  NAND U36867 ( .A(n17952), .B(n23930), .Z(n58110) );
  OR U36868 ( .A(n17953), .B(n58110), .Z(n17954) );
  NAND U36869 ( .A(n17955), .B(n17954), .Z(n17957) );
  NANDN U36870 ( .A(y[5658]), .B(x[5658]), .Z(n17956) );
  NANDN U36871 ( .A(y[5659]), .B(x[5659]), .Z(n23927) );
  AND U36872 ( .A(n17956), .B(n23927), .Z(n51319) );
  AND U36873 ( .A(n17957), .B(n51319), .Z(n17958) );
  NOR U36874 ( .A(n23929), .B(n17958), .Z(n17959) );
  NAND U36875 ( .A(n23928), .B(n17959), .Z(n17960) );
  NANDN U36876 ( .A(n58115), .B(n17960), .Z(n17961) );
  AND U36877 ( .A(n23926), .B(n17961), .Z(n17962) );
  NANDN U36878 ( .A(x[5661]), .B(y[5661]), .Z(n58116) );
  NAND U36879 ( .A(n17962), .B(n58116), .Z(n17963) );
  NANDN U36880 ( .A(n58118), .B(n17963), .Z(n17964) );
  AND U36881 ( .A(n23924), .B(n17964), .Z(n17965) );
  NANDN U36882 ( .A(x[5663]), .B(y[5663]), .Z(n51317) );
  AND U36883 ( .A(n17965), .B(n51317), .Z(n17967) );
  NANDN U36884 ( .A(y[5664]), .B(x[5664]), .Z(n17966) );
  NANDN U36885 ( .A(y[5665]), .B(x[5665]), .Z(n23922) );
  NAND U36886 ( .A(n17966), .B(n23922), .Z(n58119) );
  OR U36887 ( .A(n17967), .B(n58119), .Z(n17968) );
  AND U36888 ( .A(n58121), .B(n17968), .Z(n17969) );
  OR U36889 ( .A(n58122), .B(n17969), .Z(n17970) );
  NAND U36890 ( .A(n17971), .B(n17970), .Z(n17972) );
  NAND U36891 ( .A(n58125), .B(n17972), .Z(n17973) );
  AND U36892 ( .A(n23917), .B(n17973), .Z(n17974) );
  NANDN U36893 ( .A(n44473), .B(n17974), .Z(n17975) );
  NAND U36894 ( .A(n58126), .B(n17975), .Z(n17976) );
  NANDN U36895 ( .A(n51314), .B(n17976), .Z(n17977) );
  NANDN U36896 ( .A(y[5672]), .B(x[5672]), .Z(n23914) );
  NANDN U36897 ( .A(y[5673]), .B(x[5673]), .Z(n23911) );
  AND U36898 ( .A(n23914), .B(n23911), .Z(n51313) );
  AND U36899 ( .A(n17977), .B(n51313), .Z(n17979) );
  XNOR U36900 ( .A(x[5674]), .B(y[5674]), .Z(n23912) );
  NANDN U36901 ( .A(x[5673]), .B(y[5673]), .Z(n58127) );
  AND U36902 ( .A(n23912), .B(n58127), .Z(n17978) );
  NANDN U36903 ( .A(n17979), .B(n17978), .Z(n17980) );
  AND U36904 ( .A(n58128), .B(n17980), .Z(n17981) );
  ANDN U36905 ( .B(n58129), .A(n17981), .Z(n17982) );
  NAND U36906 ( .A(n23910), .B(n17982), .Z(n17983) );
  NANDN U36907 ( .A(n58131), .B(n17983), .Z(n17984) );
  AND U36908 ( .A(n23908), .B(n17984), .Z(n17985) );
  NANDN U36909 ( .A(x[5677]), .B(y[5677]), .Z(n58135) );
  AND U36910 ( .A(n17985), .B(n58135), .Z(n17987) );
  NANDN U36911 ( .A(y[5678]), .B(x[5678]), .Z(n17986) );
  NANDN U36912 ( .A(y[5679]), .B(x[5679]), .Z(n23905) );
  NAND U36913 ( .A(n17986), .B(n23905), .Z(n58137) );
  OR U36914 ( .A(n17987), .B(n58137), .Z(n17988) );
  AND U36915 ( .A(n23906), .B(n17988), .Z(n17989) );
  NANDN U36916 ( .A(x[5679]), .B(y[5679]), .Z(n58138) );
  AND U36917 ( .A(n17989), .B(n58138), .Z(n17991) );
  NANDN U36918 ( .A(y[5680]), .B(x[5680]), .Z(n17990) );
  NANDN U36919 ( .A(y[5681]), .B(x[5681]), .Z(n23903) );
  AND U36920 ( .A(n17990), .B(n23903), .Z(n58140) );
  NANDN U36921 ( .A(n17991), .B(n58140), .Z(n17992) );
  NAND U36922 ( .A(n17993), .B(n17992), .Z(n17994) );
  AND U36923 ( .A(n58143), .B(n17994), .Z(n17995) );
  NOR U36924 ( .A(n23902), .B(n17995), .Z(n17996) );
  NAND U36925 ( .A(n44508), .B(n17996), .Z(n17997) );
  NANDN U36926 ( .A(n58144), .B(n17997), .Z(n17998) );
  AND U36927 ( .A(n23901), .B(n17998), .Z(n17999) );
  NANDN U36928 ( .A(x[5685]), .B(y[5685]), .Z(n58146) );
  AND U36929 ( .A(n17999), .B(n58146), .Z(n18001) );
  NANDN U36930 ( .A(y[5686]), .B(x[5686]), .Z(n18000) );
  NANDN U36931 ( .A(y[5687]), .B(x[5687]), .Z(n23897) );
  AND U36932 ( .A(n18000), .B(n23897), .Z(n51309) );
  NANDN U36933 ( .A(n18001), .B(n51309), .Z(n18002) );
  NAND U36934 ( .A(n23898), .B(n18002), .Z(n18003) );
  ANDN U36935 ( .B(y[5687]), .A(x[5687]), .Z(n23899) );
  OR U36936 ( .A(n18003), .B(n23899), .Z(n18004) );
  NAND U36937 ( .A(n58150), .B(n18004), .Z(n18006) );
  XNOR U36938 ( .A(x[5690]), .B(y[5690]), .Z(n23896) );
  NANDN U36939 ( .A(x[5689]), .B(y[5689]), .Z(n58151) );
  NAND U36940 ( .A(n23896), .B(n58151), .Z(n18005) );
  ANDN U36941 ( .B(n18006), .A(n18005), .Z(n18007) );
  OR U36942 ( .A(n58153), .B(n18007), .Z(n18008) );
  NAND U36943 ( .A(n58154), .B(n18008), .Z(n18009) );
  NANDN U36944 ( .A(n58155), .B(n18009), .Z(n18010) );
  AND U36945 ( .A(n23891), .B(n18010), .Z(n18011) );
  NANDN U36946 ( .A(x[5693]), .B(y[5693]), .Z(n51307) );
  AND U36947 ( .A(n18011), .B(n51307), .Z(n18013) );
  NANDN U36948 ( .A(y[5694]), .B(x[5694]), .Z(n18012) );
  NANDN U36949 ( .A(y[5695]), .B(x[5695]), .Z(n23887) );
  AND U36950 ( .A(n18012), .B(n23887), .Z(n51306) );
  NANDN U36951 ( .A(n18013), .B(n51306), .Z(n18014) );
  NAND U36952 ( .A(n23888), .B(n18014), .Z(n18015) );
  ANDN U36953 ( .B(y[5695]), .A(x[5695]), .Z(n23889) );
  OR U36954 ( .A(n18015), .B(n23889), .Z(n18016) );
  NAND U36955 ( .A(n58158), .B(n18016), .Z(n18018) );
  XNOR U36956 ( .A(x[5698]), .B(y[5698]), .Z(n23886) );
  NANDN U36957 ( .A(x[5697]), .B(y[5697]), .Z(n51304) );
  NAND U36958 ( .A(n23886), .B(n51304), .Z(n18017) );
  ANDN U36959 ( .B(n18018), .A(n18017), .Z(n18019) );
  OR U36960 ( .A(n58159), .B(n18019), .Z(n18020) );
  NAND U36961 ( .A(n58161), .B(n18020), .Z(n18021) );
  NANDN U36962 ( .A(n58162), .B(n18021), .Z(n18022) );
  AND U36963 ( .A(n23881), .B(n18022), .Z(n18023) );
  NANDN U36964 ( .A(x[5701]), .B(y[5701]), .Z(n58163) );
  AND U36965 ( .A(n18023), .B(n58163), .Z(n18025) );
  NANDN U36966 ( .A(y[5702]), .B(x[5702]), .Z(n18024) );
  NANDN U36967 ( .A(y[5703]), .B(x[5703]), .Z(n23879) );
  NAND U36968 ( .A(n18024), .B(n23879), .Z(n58165) );
  OR U36969 ( .A(n18025), .B(n58165), .Z(n18026) );
  AND U36970 ( .A(n58166), .B(n18026), .Z(n18027) );
  OR U36971 ( .A(n58167), .B(n18027), .Z(n18028) );
  NAND U36972 ( .A(n58168), .B(n18028), .Z(n18029) );
  NANDN U36973 ( .A(n58169), .B(n18029), .Z(n18030) );
  AND U36974 ( .A(n44561), .B(n18030), .Z(n18031) );
  NANDN U36975 ( .A(x[5707]), .B(y[5707]), .Z(n58170) );
  AND U36976 ( .A(n18031), .B(n58170), .Z(n18033) );
  NANDN U36977 ( .A(y[5708]), .B(x[5708]), .Z(n18032) );
  NANDN U36978 ( .A(y[5709]), .B(x[5709]), .Z(n23871) );
  NAND U36979 ( .A(n18032), .B(n23871), .Z(n58172) );
  OR U36980 ( .A(n18033), .B(n58172), .Z(n18034) );
  AND U36981 ( .A(n23872), .B(n18034), .Z(n18035) );
  NANDN U36982 ( .A(x[5709]), .B(y[5709]), .Z(n51302) );
  AND U36983 ( .A(n18035), .B(n51302), .Z(n18037) );
  ANDN U36984 ( .B(x[5711]), .A(y[5711]), .Z(n44572) );
  NANDN U36985 ( .A(y[5710]), .B(x[5710]), .Z(n18036) );
  NANDN U36986 ( .A(n44572), .B(n18036), .Z(n58173) );
  OR U36987 ( .A(n18037), .B(n58173), .Z(n18038) );
  NAND U36988 ( .A(n18039), .B(n18038), .Z(n18041) );
  NANDN U36989 ( .A(y[5712]), .B(x[5712]), .Z(n18040) );
  NANDN U36990 ( .A(y[5713]), .B(x[5713]), .Z(n23868) );
  AND U36991 ( .A(n18040), .B(n23868), .Z(n51301) );
  AND U36992 ( .A(n18041), .B(n51301), .Z(n18042) );
  NOR U36993 ( .A(n44573), .B(n18042), .Z(n18043) );
  NAND U36994 ( .A(n23869), .B(n18043), .Z(n18044) );
  NANDN U36995 ( .A(n51299), .B(n18044), .Z(n18045) );
  XNOR U36996 ( .A(y[5716]), .B(x[5716]), .Z(n23867) );
  NANDN U36997 ( .A(x[5715]), .B(y[5715]), .Z(n44578) );
  AND U36998 ( .A(n23867), .B(n44578), .Z(n51298) );
  AND U36999 ( .A(n18045), .B(n51298), .Z(n18047) );
  NANDN U37000 ( .A(y[5716]), .B(x[5716]), .Z(n18046) );
  NANDN U37001 ( .A(y[5717]), .B(x[5717]), .Z(n23864) );
  AND U37002 ( .A(n18046), .B(n23864), .Z(n58179) );
  NANDN U37003 ( .A(n18047), .B(n58179), .Z(n18048) );
  NAND U37004 ( .A(n18049), .B(n18048), .Z(n18051) );
  NANDN U37005 ( .A(y[5718]), .B(x[5718]), .Z(n18050) );
  NANDN U37006 ( .A(y[5719]), .B(x[5719]), .Z(n23862) );
  AND U37007 ( .A(n18050), .B(n23862), .Z(n51297) );
  AND U37008 ( .A(n18051), .B(n51297), .Z(n18052) );
  ANDN U37009 ( .B(n18053), .A(n18052), .Z(n18054) );
  ANDN U37010 ( .B(n58184), .A(n18054), .Z(n18055) );
  ANDN U37011 ( .B(n58185), .A(n18055), .Z(n18056) );
  NAND U37012 ( .A(n23861), .B(n18056), .Z(n18057) );
  NANDN U37013 ( .A(n58187), .B(n18057), .Z(n18058) );
  AND U37014 ( .A(n23859), .B(n18058), .Z(n18059) );
  NANDN U37015 ( .A(x[5723]), .B(y[5723]), .Z(n51295) );
  AND U37016 ( .A(n18059), .B(n51295), .Z(n18061) );
  NANDN U37017 ( .A(y[5724]), .B(x[5724]), .Z(n18060) );
  NANDN U37018 ( .A(y[5725]), .B(x[5725]), .Z(n23856) );
  NAND U37019 ( .A(n18060), .B(n23856), .Z(n58189) );
  OR U37020 ( .A(n18061), .B(n58189), .Z(n18062) );
  AND U37021 ( .A(n23857), .B(n18062), .Z(n18063) );
  NANDN U37022 ( .A(x[5725]), .B(y[5725]), .Z(n58190) );
  AND U37023 ( .A(n18063), .B(n58190), .Z(n18065) );
  NANDN U37024 ( .A(y[5726]), .B(x[5726]), .Z(n18064) );
  NANDN U37025 ( .A(y[5727]), .B(x[5727]), .Z(n23854) );
  AND U37026 ( .A(n18064), .B(n23854), .Z(n51294) );
  NANDN U37027 ( .A(n18065), .B(n51294), .Z(n18066) );
  NAND U37028 ( .A(n18067), .B(n18066), .Z(n18068) );
  AND U37029 ( .A(n58194), .B(n18068), .Z(n18069) );
  ANDN U37030 ( .B(n58195), .A(n18069), .Z(n18070) );
  NAND U37031 ( .A(n23853), .B(n18070), .Z(n18071) );
  NANDN U37032 ( .A(n51293), .B(n18071), .Z(n18072) );
  XNOR U37033 ( .A(y[5732]), .B(x[5732]), .Z(n44618) );
  NANDN U37034 ( .A(x[5731]), .B(y[5731]), .Z(n44613) );
  AND U37035 ( .A(n44618), .B(n44613), .Z(n51292) );
  AND U37036 ( .A(n18072), .B(n51292), .Z(n18074) );
  NANDN U37037 ( .A(y[5732]), .B(x[5732]), .Z(n18073) );
  NANDN U37038 ( .A(y[5733]), .B(x[5733]), .Z(n44624) );
  AND U37039 ( .A(n18073), .B(n44624), .Z(n58197) );
  NANDN U37040 ( .A(n18074), .B(n58197), .Z(n18075) );
  NAND U37041 ( .A(n18076), .B(n18075), .Z(n18077) );
  AND U37042 ( .A(n58201), .B(n18077), .Z(n18078) );
  NOR U37043 ( .A(n58202), .B(n18078), .Z(n18079) );
  NAND U37044 ( .A(n44631), .B(n18079), .Z(n18080) );
  NANDN U37045 ( .A(n58204), .B(n18080), .Z(n18081) );
  AND U37046 ( .A(n23851), .B(n18081), .Z(n18082) );
  NANDN U37047 ( .A(x[5737]), .B(y[5737]), .Z(n51290) );
  NAND U37048 ( .A(n18082), .B(n51290), .Z(n18083) );
  NANDN U37049 ( .A(n58205), .B(n18083), .Z(n18084) );
  AND U37050 ( .A(n23849), .B(n18084), .Z(n18085) );
  NANDN U37051 ( .A(x[5739]), .B(y[5739]), .Z(n58206) );
  AND U37052 ( .A(n18085), .B(n58206), .Z(n18086) );
  OR U37053 ( .A(n58208), .B(n18086), .Z(n18087) );
  NAND U37054 ( .A(n18088), .B(n18087), .Z(n18089) );
  AND U37055 ( .A(n58210), .B(n18089), .Z(n18090) );
  ANDN U37056 ( .B(n58211), .A(n18090), .Z(n18091) );
  NAND U37057 ( .A(n23845), .B(n18091), .Z(n18092) );
  NANDN U37058 ( .A(n58214), .B(n18092), .Z(n18093) );
  AND U37059 ( .A(n23843), .B(n18093), .Z(n18094) );
  NANDN U37060 ( .A(x[5745]), .B(y[5745]), .Z(n51287) );
  AND U37061 ( .A(n18094), .B(n51287), .Z(n18096) );
  NANDN U37062 ( .A(y[5746]), .B(x[5746]), .Z(n18095) );
  NANDN U37063 ( .A(y[5747]), .B(x[5747]), .Z(n23841) );
  AND U37064 ( .A(n18095), .B(n23841), .Z(n58215) );
  NANDN U37065 ( .A(n18096), .B(n58215), .Z(n18097) );
  AND U37066 ( .A(n58216), .B(n18097), .Z(n18098) );
  NANDN U37067 ( .A(y[5748]), .B(x[5748]), .Z(n23840) );
  NANDN U37068 ( .A(y[5749]), .B(x[5749]), .Z(n23838) );
  AND U37069 ( .A(n23840), .B(n23838), .Z(n51286) );
  NANDN U37070 ( .A(n18098), .B(n51286), .Z(n18099) );
  NAND U37071 ( .A(n18100), .B(n18099), .Z(n18101) );
  AND U37072 ( .A(n58219), .B(n18101), .Z(n18102) );
  ANDN U37073 ( .B(n51284), .A(n18102), .Z(n18103) );
  NAND U37074 ( .A(n23837), .B(n18103), .Z(n18104) );
  NANDN U37075 ( .A(n58220), .B(n18104), .Z(n18105) );
  AND U37076 ( .A(n23835), .B(n18105), .Z(n18106) );
  NANDN U37077 ( .A(x[5753]), .B(y[5753]), .Z(n58222) );
  AND U37078 ( .A(n18106), .B(n58222), .Z(n18108) );
  NANDN U37079 ( .A(y[5754]), .B(x[5754]), .Z(n18107) );
  NANDN U37080 ( .A(y[5755]), .B(x[5755]), .Z(n23832) );
  NAND U37081 ( .A(n18107), .B(n23832), .Z(n58223) );
  OR U37082 ( .A(n18108), .B(n58223), .Z(n18109) );
  AND U37083 ( .A(n58225), .B(n18109), .Z(n18110) );
  NAND U37084 ( .A(n23833), .B(n18110), .Z(n18111) );
  NAND U37085 ( .A(n58227), .B(n18111), .Z(n18112) );
  ANDN U37086 ( .B(y[5757]), .A(x[5757]), .Z(n44677) );
  ANDN U37087 ( .B(n18112), .A(n44677), .Z(n18113) );
  NAND U37088 ( .A(n23831), .B(n18113), .Z(n18115) );
  NANDN U37089 ( .A(y[5758]), .B(x[5758]), .Z(n18114) );
  NANDN U37090 ( .A(y[5759]), .B(x[5759]), .Z(n23828) );
  AND U37091 ( .A(n18114), .B(n23828), .Z(n58230) );
  AND U37092 ( .A(n18115), .B(n58230), .Z(n18117) );
  XNOR U37093 ( .A(x[5760]), .B(y[5760]), .Z(n23829) );
  ANDN U37094 ( .B(y[5759]), .A(x[5759]), .Z(n44682) );
  ANDN U37095 ( .B(n23829), .A(n44682), .Z(n18116) );
  NANDN U37096 ( .A(n18117), .B(n18116), .Z(n18119) );
  NANDN U37097 ( .A(y[5760]), .B(x[5760]), .Z(n18118) );
  NANDN U37098 ( .A(y[5761]), .B(x[5761]), .Z(n23827) );
  AND U37099 ( .A(n18118), .B(n23827), .Z(n58231) );
  AND U37100 ( .A(n18119), .B(n58231), .Z(n18120) );
  NANDN U37101 ( .A(x[5761]), .B(y[5761]), .Z(n44688) );
  NANDN U37102 ( .A(x[5762]), .B(y[5762]), .Z(n23824) );
  NAND U37103 ( .A(n44688), .B(n23824), .Z(n51281) );
  OR U37104 ( .A(n18120), .B(n51281), .Z(n18121) );
  NAND U37105 ( .A(n51280), .B(n18121), .Z(n18122) );
  NANDN U37106 ( .A(n58232), .B(n18122), .Z(n18123) );
  NANDN U37107 ( .A(y[5764]), .B(x[5764]), .Z(n23822) );
  NANDN U37108 ( .A(y[5765]), .B(x[5765]), .Z(n23819) );
  AND U37109 ( .A(n23822), .B(n23819), .Z(n58233) );
  AND U37110 ( .A(n18123), .B(n58233), .Z(n18124) );
  NANDN U37111 ( .A(x[5765]), .B(y[5765]), .Z(n23820) );
  NANDN U37112 ( .A(x[5766]), .B(y[5766]), .Z(n23817) );
  NAND U37113 ( .A(n23820), .B(n23817), .Z(n58234) );
  OR U37114 ( .A(n18124), .B(n58234), .Z(n18125) );
  NANDN U37115 ( .A(y[5766]), .B(x[5766]), .Z(n23818) );
  NANDN U37116 ( .A(y[5767]), .B(x[5767]), .Z(n44704) );
  AND U37117 ( .A(n23818), .B(n44704), .Z(n58237) );
  AND U37118 ( .A(n18125), .B(n58237), .Z(n18126) );
  NANDN U37119 ( .A(x[5767]), .B(y[5767]), .Z(n23816) );
  NANDN U37120 ( .A(x[5768]), .B(y[5768]), .Z(n23815) );
  NAND U37121 ( .A(n23816), .B(n23815), .Z(n51279) );
  OR U37122 ( .A(n18126), .B(n51279), .Z(n18127) );
  NAND U37123 ( .A(n58239), .B(n18127), .Z(n18128) );
  NANDN U37124 ( .A(n58240), .B(n18128), .Z(n18129) );
  NANDN U37125 ( .A(y[5770]), .B(x[5770]), .Z(n44708) );
  NANDN U37126 ( .A(y[5771]), .B(x[5771]), .Z(n44716) );
  AND U37127 ( .A(n44708), .B(n44716), .Z(n58241) );
  AND U37128 ( .A(n18129), .B(n58241), .Z(n18130) );
  NANDN U37129 ( .A(x[5771]), .B(y[5771]), .Z(n23812) );
  NANDN U37130 ( .A(x[5772]), .B(y[5772]), .Z(n23811) );
  NAND U37131 ( .A(n23812), .B(n23811), .Z(n51278) );
  OR U37132 ( .A(n18130), .B(n51278), .Z(n18131) );
  NAND U37133 ( .A(n51277), .B(n18131), .Z(n18132) );
  AND U37134 ( .A(n23810), .B(n18132), .Z(n18133) );
  NANDN U37135 ( .A(x[5773]), .B(y[5773]), .Z(n58242) );
  AND U37136 ( .A(n18133), .B(n58242), .Z(n18135) );
  NANDN U37137 ( .A(y[5774]), .B(x[5774]), .Z(n18134) );
  NANDN U37138 ( .A(y[5775]), .B(x[5775]), .Z(n23807) );
  NAND U37139 ( .A(n18134), .B(n23807), .Z(n58244) );
  OR U37140 ( .A(n18135), .B(n58244), .Z(n18136) );
  AND U37141 ( .A(n58245), .B(n18136), .Z(n18137) );
  OR U37142 ( .A(n58246), .B(n18137), .Z(n18138) );
  NAND U37143 ( .A(n58247), .B(n18138), .Z(n18139) );
  NANDN U37144 ( .A(n58248), .B(n18139), .Z(n18140) );
  AND U37145 ( .A(n23800), .B(n18140), .Z(n18141) );
  NANDN U37146 ( .A(x[5779]), .B(y[5779]), .Z(n58250) );
  AND U37147 ( .A(n18141), .B(n58250), .Z(n18143) );
  NANDN U37148 ( .A(y[5780]), .B(x[5780]), .Z(n18142) );
  NANDN U37149 ( .A(y[5781]), .B(x[5781]), .Z(n23797) );
  AND U37150 ( .A(n18142), .B(n23797), .Z(n58252) );
  NANDN U37151 ( .A(n18143), .B(n58252), .Z(n18144) );
  NAND U37152 ( .A(n18145), .B(n18144), .Z(n18146) );
  AND U37153 ( .A(n58253), .B(n18146), .Z(n18147) );
  ANDN U37154 ( .B(n58255), .A(n18147), .Z(n18148) );
  NAND U37155 ( .A(n23796), .B(n18148), .Z(n18149) );
  NANDN U37156 ( .A(n58256), .B(n18149), .Z(n18150) );
  AND U37157 ( .A(n23794), .B(n18150), .Z(n18151) );
  NANDN U37158 ( .A(x[5785]), .B(y[5785]), .Z(n58257) );
  AND U37159 ( .A(n18151), .B(n58257), .Z(n18152) );
  OR U37160 ( .A(n58259), .B(n18152), .Z(n18153) );
  AND U37161 ( .A(n23792), .B(n18153), .Z(n18154) );
  NANDN U37162 ( .A(x[5787]), .B(y[5787]), .Z(n58260) );
  AND U37163 ( .A(n18154), .B(n58260), .Z(n18156) );
  NANDN U37164 ( .A(y[5788]), .B(x[5788]), .Z(n18155) );
  NANDN U37165 ( .A(y[5789]), .B(x[5789]), .Z(n44753) );
  AND U37166 ( .A(n18155), .B(n44753), .Z(n58262) );
  NANDN U37167 ( .A(n18156), .B(n58262), .Z(n18157) );
  NAND U37168 ( .A(n18158), .B(n18157), .Z(n18159) );
  AND U37169 ( .A(n58263), .B(n18159), .Z(n18160) );
  ANDN U37170 ( .B(n51271), .A(n18160), .Z(n18161) );
  NAND U37171 ( .A(n44761), .B(n18161), .Z(n18162) );
  NANDN U37172 ( .A(n51270), .B(n18162), .Z(n18163) );
  AND U37173 ( .A(n23790), .B(n18163), .Z(n18164) );
  NANDN U37174 ( .A(x[5793]), .B(y[5793]), .Z(n58266) );
  AND U37175 ( .A(n18164), .B(n58266), .Z(n18166) );
  NANDN U37176 ( .A(y[5794]), .B(x[5794]), .Z(n18165) );
  NANDN U37177 ( .A(y[5795]), .B(x[5795]), .Z(n23787) );
  NAND U37178 ( .A(n18165), .B(n23787), .Z(n58268) );
  OR U37179 ( .A(n18166), .B(n58268), .Z(n18167) );
  AND U37180 ( .A(n23788), .B(n18167), .Z(n18168) );
  NANDN U37181 ( .A(x[5795]), .B(y[5795]), .Z(n58269) );
  AND U37182 ( .A(n18168), .B(n58269), .Z(n18170) );
  NANDN U37183 ( .A(y[5796]), .B(x[5796]), .Z(n18169) );
  NANDN U37184 ( .A(y[5797]), .B(x[5797]), .Z(n23785) );
  AND U37185 ( .A(n18169), .B(n23785), .Z(n58271) );
  NANDN U37186 ( .A(n18170), .B(n58271), .Z(n18171) );
  NAND U37187 ( .A(n18172), .B(n18171), .Z(n18173) );
  AND U37188 ( .A(n58274), .B(n18173), .Z(n18174) );
  ANDN U37189 ( .B(n58276), .A(n18174), .Z(n18175) );
  NANDN U37190 ( .A(n44780), .B(n18175), .Z(n18176) );
  NANDN U37191 ( .A(n58277), .B(n18176), .Z(n18177) );
  AND U37192 ( .A(n23784), .B(n18177), .Z(n18178) );
  NANDN U37193 ( .A(x[5801]), .B(y[5801]), .Z(n58278) );
  AND U37194 ( .A(n18178), .B(n58278), .Z(n18180) );
  NANDN U37195 ( .A(y[5802]), .B(x[5802]), .Z(n18179) );
  NANDN U37196 ( .A(y[5803]), .B(x[5803]), .Z(n23781) );
  NAND U37197 ( .A(n18179), .B(n23781), .Z(n58280) );
  OR U37198 ( .A(n18180), .B(n58280), .Z(n18181) );
  AND U37199 ( .A(n23782), .B(n18181), .Z(n18182) );
  NANDN U37200 ( .A(x[5803]), .B(y[5803]), .Z(n58281) );
  AND U37201 ( .A(n18182), .B(n58281), .Z(n18184) );
  NANDN U37202 ( .A(y[5804]), .B(x[5804]), .Z(n18183) );
  NANDN U37203 ( .A(y[5805]), .B(x[5805]), .Z(n23779) );
  AND U37204 ( .A(n18183), .B(n23779), .Z(n58284) );
  NANDN U37205 ( .A(n18184), .B(n58284), .Z(n18185) );
  NAND U37206 ( .A(n18186), .B(n18185), .Z(n18187) );
  AND U37207 ( .A(n58290), .B(n18187), .Z(n18188) );
  ANDN U37208 ( .B(n58292), .A(n18188), .Z(n18189) );
  NAND U37209 ( .A(n23778), .B(n18189), .Z(n18190) );
  NANDN U37210 ( .A(n58296), .B(n18190), .Z(n18191) );
  AND U37211 ( .A(n23776), .B(n18191), .Z(n18192) );
  NANDN U37212 ( .A(x[5809]), .B(y[5809]), .Z(n58298) );
  AND U37213 ( .A(n18192), .B(n58298), .Z(n18194) );
  NANDN U37214 ( .A(y[5810]), .B(x[5810]), .Z(n18193) );
  NANDN U37215 ( .A(y[5811]), .B(x[5811]), .Z(n23773) );
  NAND U37216 ( .A(n18193), .B(n23773), .Z(n58301) );
  OR U37217 ( .A(n18194), .B(n58301), .Z(n18195) );
  AND U37218 ( .A(n23774), .B(n18195), .Z(n18196) );
  NANDN U37219 ( .A(x[5811]), .B(y[5811]), .Z(n58304) );
  AND U37220 ( .A(n18196), .B(n58304), .Z(n18198) );
  NANDN U37221 ( .A(y[5812]), .B(x[5812]), .Z(n18197) );
  NANDN U37222 ( .A(y[5813]), .B(x[5813]), .Z(n23772) );
  NAND U37223 ( .A(n18197), .B(n23772), .Z(n58307) );
  OR U37224 ( .A(n18198), .B(n58307), .Z(n18199) );
  AND U37225 ( .A(n58310), .B(n18199), .Z(n18200) );
  OR U37226 ( .A(n58312), .B(n18200), .Z(n18201) );
  NAND U37227 ( .A(n18202), .B(n18201), .Z(n18203) );
  NANDN U37228 ( .A(n58316), .B(n18203), .Z(n18204) );
  AND U37229 ( .A(n58318), .B(n18204), .Z(n18206) );
  NANDN U37230 ( .A(y[5818]), .B(x[5818]), .Z(n18205) );
  NANDN U37231 ( .A(y[5819]), .B(x[5819]), .Z(n23764) );
  AND U37232 ( .A(n18205), .B(n23764), .Z(n58319) );
  NANDN U37233 ( .A(n18206), .B(n58319), .Z(n18207) );
  NAND U37234 ( .A(n18208), .B(n18207), .Z(n18209) );
  AND U37235 ( .A(n58321), .B(n18209), .Z(n18210) );
  NOR U37236 ( .A(n44826), .B(n18210), .Z(n18211) );
  NAND U37237 ( .A(n23763), .B(n18211), .Z(n18212) );
  NANDN U37238 ( .A(n58324), .B(n18212), .Z(n18213) );
  AND U37239 ( .A(n58325), .B(n18213), .Z(n18214) );
  NANDN U37240 ( .A(y[5824]), .B(x[5824]), .Z(n23759) );
  NANDN U37241 ( .A(y[5825]), .B(x[5825]), .Z(n23756) );
  AND U37242 ( .A(n23759), .B(n23756), .Z(n58326) );
  NANDN U37243 ( .A(n18214), .B(n58326), .Z(n18215) );
  NANDN U37244 ( .A(y[5828]), .B(x[5828]), .Z(n18216) );
  NANDN U37245 ( .A(y[5829]), .B(x[5829]), .Z(n23754) );
  AND U37246 ( .A(n18216), .B(n23754), .Z(n51260) );
  NANDN U37247 ( .A(y[5836]), .B(x[5836]), .Z(n18217) );
  NANDN U37248 ( .A(y[5837]), .B(x[5837]), .Z(n23744) );
  AND U37249 ( .A(n18217), .B(n23744), .Z(n51259) );
  AND U37250 ( .A(n18218), .B(n51259), .Z(n18219) );
  NOR U37251 ( .A(n44863), .B(n18219), .Z(n18220) );
  NAND U37252 ( .A(n23745), .B(n18220), .Z(n18221) );
  NANDN U37253 ( .A(n58343), .B(n18221), .Z(n18222) );
  AND U37254 ( .A(n23743), .B(n18222), .Z(n18223) );
  NANDN U37255 ( .A(x[5839]), .B(y[5839]), .Z(n58344) );
  AND U37256 ( .A(n18223), .B(n58344), .Z(n18224) );
  OR U37257 ( .A(n58346), .B(n18224), .Z(n18225) );
  AND U37258 ( .A(n23741), .B(n18225), .Z(n18226) );
  NANDN U37259 ( .A(x[5841]), .B(y[5841]), .Z(n51257) );
  AND U37260 ( .A(n18226), .B(n51257), .Z(n18228) );
  NANDN U37261 ( .A(y[5842]), .B(x[5842]), .Z(n18227) );
  NANDN U37262 ( .A(y[5843]), .B(x[5843]), .Z(n23738) );
  AND U37263 ( .A(n18227), .B(n23738), .Z(n58347) );
  NANDN U37264 ( .A(n18228), .B(n58347), .Z(n18229) );
  NAND U37265 ( .A(n18230), .B(n18229), .Z(n18232) );
  NANDN U37266 ( .A(y[5844]), .B(x[5844]), .Z(n18231) );
  NANDN U37267 ( .A(y[5845]), .B(x[5845]), .Z(n23736) );
  AND U37268 ( .A(n18231), .B(n23736), .Z(n51256) );
  AND U37269 ( .A(n18232), .B(n51256), .Z(n18233) );
  NOR U37270 ( .A(n44880), .B(n18233), .Z(n18234) );
  NAND U37271 ( .A(n23737), .B(n18234), .Z(n18235) );
  NANDN U37272 ( .A(n58353), .B(n18235), .Z(n18236) );
  AND U37273 ( .A(n23735), .B(n18236), .Z(n18237) );
  NANDN U37274 ( .A(x[5847]), .B(y[5847]), .Z(n58354) );
  AND U37275 ( .A(n18237), .B(n58354), .Z(n18239) );
  NANDN U37276 ( .A(y[5848]), .B(x[5848]), .Z(n18238) );
  NANDN U37277 ( .A(y[5849]), .B(x[5849]), .Z(n23732) );
  NAND U37278 ( .A(n18238), .B(n23732), .Z(n58356) );
  OR U37279 ( .A(n18239), .B(n58356), .Z(n18240) );
  AND U37280 ( .A(n23733), .B(n18240), .Z(n18241) );
  NANDN U37281 ( .A(x[5849]), .B(y[5849]), .Z(n51254) );
  AND U37282 ( .A(n18241), .B(n51254), .Z(n18243) );
  NANDN U37283 ( .A(y[5850]), .B(x[5850]), .Z(n18242) );
  ANDN U37284 ( .B(x[5851]), .A(y[5851]), .Z(n44898) );
  ANDN U37285 ( .B(n18242), .A(n44898), .Z(n58357) );
  NANDN U37286 ( .A(n18243), .B(n58357), .Z(n18244) );
  NAND U37287 ( .A(n18245), .B(n18244), .Z(n18247) );
  NANDN U37288 ( .A(y[5852]), .B(x[5852]), .Z(n18246) );
  NANDN U37289 ( .A(y[5853]), .B(x[5853]), .Z(n23730) );
  AND U37290 ( .A(n18246), .B(n23730), .Z(n51253) );
  AND U37291 ( .A(n18247), .B(n51253), .Z(n18248) );
  NOR U37292 ( .A(n44899), .B(n18248), .Z(n18249) );
  NAND U37293 ( .A(n23731), .B(n18249), .Z(n18250) );
  NANDN U37294 ( .A(n58362), .B(n18250), .Z(n18251) );
  AND U37295 ( .A(n23729), .B(n18251), .Z(n18252) );
  NANDN U37296 ( .A(x[5855]), .B(y[5855]), .Z(n58363) );
  NAND U37297 ( .A(n18252), .B(n58363), .Z(n18253) );
  NANDN U37298 ( .A(n58365), .B(n18253), .Z(n18254) );
  AND U37299 ( .A(n58367), .B(n18254), .Z(n18255) );
  OR U37300 ( .A(n58368), .B(n18255), .Z(n18256) );
  NAND U37301 ( .A(n58369), .B(n18256), .Z(n18257) );
  NANDN U37302 ( .A(n58370), .B(n18257), .Z(n18258) );
  AND U37303 ( .A(n23720), .B(n18258), .Z(n18259) );
  NANDN U37304 ( .A(x[5861]), .B(y[5861]), .Z(n58371) );
  AND U37305 ( .A(n18259), .B(n58371), .Z(n18261) );
  NANDN U37306 ( .A(y[5862]), .B(x[5862]), .Z(n18260) );
  NANDN U37307 ( .A(y[5863]), .B(x[5863]), .Z(n23717) );
  NAND U37308 ( .A(n18260), .B(n23717), .Z(n51252) );
  OR U37309 ( .A(n18261), .B(n51252), .Z(n18262) );
  AND U37310 ( .A(n23718), .B(n18262), .Z(n18263) );
  NANDN U37311 ( .A(x[5863]), .B(y[5863]), .Z(n58374) );
  AND U37312 ( .A(n18263), .B(n58374), .Z(n18265) );
  NANDN U37313 ( .A(y[5864]), .B(x[5864]), .Z(n18264) );
  NANDN U37314 ( .A(y[5865]), .B(x[5865]), .Z(n23716) );
  NAND U37315 ( .A(n18264), .B(n23716), .Z(n58375) );
  OR U37316 ( .A(n18265), .B(n58375), .Z(n18266) );
  NAND U37317 ( .A(n58376), .B(n18266), .Z(n18267) );
  NANDN U37318 ( .A(y[5866]), .B(x[5866]), .Z(n23715) );
  NANDN U37319 ( .A(y[5867]), .B(x[5867]), .Z(n23711) );
  AND U37320 ( .A(n23715), .B(n23711), .Z(n51251) );
  AND U37321 ( .A(n18267), .B(n51251), .Z(n18268) );
  NOR U37322 ( .A(n23713), .B(n18268), .Z(n18269) );
  NAND U37323 ( .A(n23712), .B(n18269), .Z(n18270) );
  NANDN U37324 ( .A(n58379), .B(n18270), .Z(n18271) );
  AND U37325 ( .A(n23710), .B(n18271), .Z(n18272) );
  NANDN U37326 ( .A(n44934), .B(n18272), .Z(n18273) );
  NAND U37327 ( .A(n58381), .B(n18273), .Z(n18274) );
  NANDN U37328 ( .A(n51248), .B(n18274), .Z(n18275) );
  NANDN U37329 ( .A(y[5872]), .B(x[5872]), .Z(n23707) );
  NANDN U37330 ( .A(y[5873]), .B(x[5873]), .Z(n23703) );
  AND U37331 ( .A(n23707), .B(n23703), .Z(n51247) );
  AND U37332 ( .A(n18275), .B(n51247), .Z(n18276) );
  NOR U37333 ( .A(n23705), .B(n18276), .Z(n18277) );
  NAND U37334 ( .A(n23704), .B(n18277), .Z(n18278) );
  NANDN U37335 ( .A(n58384), .B(n18278), .Z(n18279) );
  AND U37336 ( .A(n23702), .B(n18279), .Z(n18280) );
  NAND U37337 ( .A(n51245), .B(n18280), .Z(n18281) );
  NANDN U37338 ( .A(n58385), .B(n18281), .Z(n18282) );
  AND U37339 ( .A(n44955), .B(n18282), .Z(n18283) );
  NANDN U37340 ( .A(x[5877]), .B(y[5877]), .Z(n58386) );
  AND U37341 ( .A(n18283), .B(n58386), .Z(n18284) );
  OR U37342 ( .A(n58389), .B(n18284), .Z(n18285) );
  NAND U37343 ( .A(n18286), .B(n18285), .Z(n18288) );
  NANDN U37344 ( .A(y[5880]), .B(x[5880]), .Z(n18287) );
  NANDN U37345 ( .A(y[5881]), .B(x[5881]), .Z(n23697) );
  AND U37346 ( .A(n18287), .B(n23697), .Z(n58392) );
  AND U37347 ( .A(n18288), .B(n58392), .Z(n18289) );
  NOR U37348 ( .A(n44962), .B(n18289), .Z(n18290) );
  NAND U37349 ( .A(n23698), .B(n18290), .Z(n18291) );
  NANDN U37350 ( .A(n58395), .B(n18291), .Z(n18292) );
  AND U37351 ( .A(n23696), .B(n18292), .Z(n18293) );
  NANDN U37352 ( .A(x[5883]), .B(y[5883]), .Z(n51243) );
  NAND U37353 ( .A(n18293), .B(n51243), .Z(n18294) );
  NANDN U37354 ( .A(n58396), .B(n18294), .Z(n18295) );
  AND U37355 ( .A(n23694), .B(n18295), .Z(n18296) );
  NANDN U37356 ( .A(x[5885]), .B(y[5885]), .Z(n58398) );
  AND U37357 ( .A(n18296), .B(n58398), .Z(n18297) );
  OR U37358 ( .A(n58399), .B(n18297), .Z(n18298) );
  NAND U37359 ( .A(n18299), .B(n18298), .Z(n18301) );
  NANDN U37360 ( .A(y[5888]), .B(x[5888]), .Z(n18300) );
  NANDN U37361 ( .A(y[5889]), .B(x[5889]), .Z(n23689) );
  AND U37362 ( .A(n18300), .B(n23689), .Z(n58402) );
  AND U37363 ( .A(n18301), .B(n58402), .Z(n18302) );
  NOR U37364 ( .A(n44979), .B(n18302), .Z(n18303) );
  NAND U37365 ( .A(n23690), .B(n18303), .Z(n18304) );
  NANDN U37366 ( .A(n58406), .B(n18304), .Z(n18305) );
  AND U37367 ( .A(n23688), .B(n18305), .Z(n18306) );
  NANDN U37368 ( .A(x[5891]), .B(y[5891]), .Z(n51241) );
  NAND U37369 ( .A(n18306), .B(n51241), .Z(n18307) );
  NANDN U37370 ( .A(n58407), .B(n18307), .Z(n18308) );
  AND U37371 ( .A(n23686), .B(n18308), .Z(n18309) );
  NANDN U37372 ( .A(x[5893]), .B(y[5893]), .Z(n58409) );
  AND U37373 ( .A(n18309), .B(n58409), .Z(n18310) );
  OR U37374 ( .A(n58410), .B(n18310), .Z(n18311) );
  NAND U37375 ( .A(n18312), .B(n18311), .Z(n18314) );
  NANDN U37376 ( .A(y[5896]), .B(x[5896]), .Z(n18313) );
  NANDN U37377 ( .A(y[5897]), .B(x[5897]), .Z(n23681) );
  AND U37378 ( .A(n18313), .B(n23681), .Z(n58413) );
  AND U37379 ( .A(n18314), .B(n58413), .Z(n18315) );
  NOR U37380 ( .A(n44996), .B(n18315), .Z(n18316) );
  NAND U37381 ( .A(n23682), .B(n18316), .Z(n18317) );
  NANDN U37382 ( .A(n58416), .B(n18317), .Z(n18318) );
  AND U37383 ( .A(n23680), .B(n18318), .Z(n18319) );
  NANDN U37384 ( .A(x[5899]), .B(y[5899]), .Z(n51239) );
  NAND U37385 ( .A(n18319), .B(n51239), .Z(n18320) );
  NANDN U37386 ( .A(n58417), .B(n18320), .Z(n18321) );
  AND U37387 ( .A(n23678), .B(n18321), .Z(n18322) );
  NANDN U37388 ( .A(x[5901]), .B(y[5901]), .Z(n58422) );
  AND U37389 ( .A(n18322), .B(n58422), .Z(n18323) );
  OR U37390 ( .A(n58423), .B(n18323), .Z(n18324) );
  NAND U37391 ( .A(n18325), .B(n18324), .Z(n18327) );
  NANDN U37392 ( .A(y[5904]), .B(x[5904]), .Z(n18326) );
  NANDN U37393 ( .A(y[5905]), .B(x[5905]), .Z(n23673) );
  AND U37394 ( .A(n18326), .B(n23673), .Z(n58426) );
  AND U37395 ( .A(n18327), .B(n58426), .Z(n18328) );
  NOR U37396 ( .A(n45013), .B(n18328), .Z(n18329) );
  NAND U37397 ( .A(n23674), .B(n18329), .Z(n18330) );
  NANDN U37398 ( .A(n58429), .B(n18330), .Z(n18331) );
  AND U37399 ( .A(n23672), .B(n18331), .Z(n18332) );
  NANDN U37400 ( .A(x[5907]), .B(y[5907]), .Z(n51237) );
  NAND U37401 ( .A(n18332), .B(n51237), .Z(n18333) );
  NANDN U37402 ( .A(n58430), .B(n18333), .Z(n18334) );
  AND U37403 ( .A(n23670), .B(n18334), .Z(n18335) );
  NANDN U37404 ( .A(x[5909]), .B(y[5909]), .Z(n58432) );
  AND U37405 ( .A(n18335), .B(n58432), .Z(n18336) );
  OR U37406 ( .A(n58433), .B(n18336), .Z(n18337) );
  NAND U37407 ( .A(n18338), .B(n18337), .Z(n18340) );
  NANDN U37408 ( .A(y[5912]), .B(x[5912]), .Z(n18339) );
  NANDN U37409 ( .A(y[5913]), .B(x[5913]), .Z(n23665) );
  AND U37410 ( .A(n18339), .B(n23665), .Z(n58436) );
  AND U37411 ( .A(n18340), .B(n58436), .Z(n18341) );
  NOR U37412 ( .A(n45030), .B(n18341), .Z(n18342) );
  NAND U37413 ( .A(n23666), .B(n18342), .Z(n18343) );
  NANDN U37414 ( .A(n58441), .B(n18343), .Z(n18344) );
  AND U37415 ( .A(n23664), .B(n18344), .Z(n18345) );
  NANDN U37416 ( .A(x[5915]), .B(y[5915]), .Z(n51235) );
  NAND U37417 ( .A(n18345), .B(n51235), .Z(n18346) );
  NANDN U37418 ( .A(n58442), .B(n18346), .Z(n18347) );
  AND U37419 ( .A(n23662), .B(n18347), .Z(n18348) );
  NANDN U37420 ( .A(x[5917]), .B(y[5917]), .Z(n58443) );
  AND U37421 ( .A(n18348), .B(n58443), .Z(n18350) );
  NANDN U37422 ( .A(y[5918]), .B(x[5918]), .Z(n18349) );
  NANDN U37423 ( .A(y[5919]), .B(x[5919]), .Z(n23659) );
  NAND U37424 ( .A(n18349), .B(n23659), .Z(n58445) );
  OR U37425 ( .A(n18350), .B(n58445), .Z(n18351) );
  XNOR U37426 ( .A(y[5920]), .B(x[5920]), .Z(n23660) );
  NANDN U37427 ( .A(x[5919]), .B(y[5919]), .Z(n45043) );
  AND U37428 ( .A(n23660), .B(n45043), .Z(n58446) );
  AND U37429 ( .A(n18351), .B(n58446), .Z(n18353) );
  NANDN U37430 ( .A(y[5920]), .B(x[5920]), .Z(n18352) );
  NANDN U37431 ( .A(y[5921]), .B(x[5921]), .Z(n23658) );
  NAND U37432 ( .A(n18352), .B(n23658), .Z(n51234) );
  OR U37433 ( .A(n18353), .B(n51234), .Z(n18354) );
  NAND U37434 ( .A(n51233), .B(n18354), .Z(n18355) );
  NAND U37435 ( .A(n58447), .B(n18355), .Z(n18356) );
  AND U37436 ( .A(n23654), .B(n18356), .Z(n18357) );
  NANDN U37437 ( .A(x[5923]), .B(y[5923]), .Z(n58450) );
  AND U37438 ( .A(n18357), .B(n58450), .Z(n18358) );
  OR U37439 ( .A(n58451), .B(n18358), .Z(n18359) );
  NAND U37440 ( .A(n18360), .B(n18359), .Z(n18362) );
  NANDN U37441 ( .A(y[5926]), .B(x[5926]), .Z(n18361) );
  NANDN U37442 ( .A(y[5927]), .B(x[5927]), .Z(n23650) );
  AND U37443 ( .A(n18361), .B(n23650), .Z(n58454) );
  AND U37444 ( .A(n18362), .B(n58454), .Z(n18363) );
  ANDN U37445 ( .B(n18364), .A(n18363), .Z(n18365) );
  ANDN U37446 ( .B(n58457), .A(n18365), .Z(n18366) );
  NOR U37447 ( .A(n45066), .B(n18366), .Z(n18367) );
  NAND U37448 ( .A(n23649), .B(n18367), .Z(n18368) );
  NANDN U37449 ( .A(n58458), .B(n18368), .Z(n18369) );
  AND U37450 ( .A(n45074), .B(n18369), .Z(n18370) );
  NANDN U37451 ( .A(x[5931]), .B(y[5931]), .Z(n58459) );
  AND U37452 ( .A(n18370), .B(n58459), .Z(n18372) );
  NANDN U37453 ( .A(y[5932]), .B(x[5932]), .Z(n18371) );
  NANDN U37454 ( .A(y[5933]), .B(x[5933]), .Z(n23646) );
  NAND U37455 ( .A(n18371), .B(n23646), .Z(n58461) );
  OR U37456 ( .A(n18372), .B(n58461), .Z(n18373) );
  AND U37457 ( .A(n23647), .B(n18373), .Z(n18374) );
  NANDN U37458 ( .A(x[5933]), .B(y[5933]), .Z(n58462) );
  AND U37459 ( .A(n18374), .B(n58462), .Z(n18376) );
  NANDN U37460 ( .A(y[5934]), .B(x[5934]), .Z(n18375) );
  NANDN U37461 ( .A(y[5935]), .B(x[5935]), .Z(n23644) );
  NAND U37462 ( .A(n18375), .B(n23644), .Z(n51229) );
  OR U37463 ( .A(n18376), .B(n51229), .Z(n18377) );
  XNOR U37464 ( .A(y[5936]), .B(x[5936]), .Z(n23645) );
  NANDN U37465 ( .A(x[5935]), .B(y[5935]), .Z(n45081) );
  AND U37466 ( .A(n23645), .B(n45081), .Z(n51228) );
  AND U37467 ( .A(n18377), .B(n51228), .Z(n18379) );
  NANDN U37468 ( .A(y[5936]), .B(x[5936]), .Z(n18378) );
  NANDN U37469 ( .A(y[5937]), .B(x[5937]), .Z(n23642) );
  NAND U37470 ( .A(n18378), .B(n23642), .Z(n58464) );
  OR U37471 ( .A(n18379), .B(n58464), .Z(n18380) );
  NAND U37472 ( .A(n18381), .B(n18380), .Z(n18382) );
  NANDN U37473 ( .A(n58467), .B(n18382), .Z(n18383) );
  AND U37474 ( .A(n23641), .B(n18383), .Z(n18384) );
  NANDN U37475 ( .A(x[5939]), .B(y[5939]), .Z(n58468) );
  AND U37476 ( .A(n18384), .B(n58468), .Z(n18386) );
  NANDN U37477 ( .A(y[5940]), .B(x[5940]), .Z(n18385) );
  NANDN U37478 ( .A(y[5941]), .B(x[5941]), .Z(n23638) );
  AND U37479 ( .A(n18385), .B(n23638), .Z(n58470) );
  NANDN U37480 ( .A(n18386), .B(n58470), .Z(n18387) );
  NAND U37481 ( .A(n23639), .B(n18387), .Z(n18388) );
  ANDN U37482 ( .B(y[5941]), .A(x[5941]), .Z(n45095) );
  OR U37483 ( .A(n18388), .B(n45095), .Z(n18389) );
  NAND U37484 ( .A(n58473), .B(n18389), .Z(n18391) );
  XNOR U37485 ( .A(x[5944]), .B(y[5944]), .Z(n23637) );
  NANDN U37486 ( .A(x[5943]), .B(y[5943]), .Z(n51226) );
  NAND U37487 ( .A(n23637), .B(n51226), .Z(n18390) );
  ANDN U37488 ( .B(n18391), .A(n18390), .Z(n18393) );
  NANDN U37489 ( .A(y[5944]), .B(x[5944]), .Z(n18392) );
  NANDN U37490 ( .A(y[5945]), .B(x[5945]), .Z(n23634) );
  NAND U37491 ( .A(n18392), .B(n23634), .Z(n58476) );
  OR U37492 ( .A(n18393), .B(n58476), .Z(n18394) );
  NAND U37493 ( .A(n18395), .B(n18394), .Z(n18396) );
  NANDN U37494 ( .A(n58480), .B(n18396), .Z(n18397) );
  AND U37495 ( .A(n23633), .B(n18397), .Z(n18398) );
  NANDN U37496 ( .A(n45108), .B(n18398), .Z(n18399) );
  NAND U37497 ( .A(n58483), .B(n18399), .Z(n18400) );
  NAND U37498 ( .A(n23631), .B(n18400), .Z(n18401) );
  ANDN U37499 ( .B(y[5949]), .A(x[5949]), .Z(n45113) );
  OR U37500 ( .A(n18401), .B(n45113), .Z(n18402) );
  NAND U37501 ( .A(n58486), .B(n18402), .Z(n18404) );
  XNOR U37502 ( .A(x[5952]), .B(y[5952]), .Z(n45121) );
  NANDN U37503 ( .A(x[5951]), .B(y[5951]), .Z(n51224) );
  NAND U37504 ( .A(n45121), .B(n51224), .Z(n18403) );
  ANDN U37505 ( .B(n18404), .A(n18403), .Z(n18405) );
  OR U37506 ( .A(n58487), .B(n18405), .Z(n18406) );
  NAND U37507 ( .A(n58488), .B(n18406), .Z(n18407) );
  NANDN U37508 ( .A(n58489), .B(n18407), .Z(n18408) );
  AND U37509 ( .A(n45133), .B(n18408), .Z(n18409) );
  NANDN U37510 ( .A(x[5955]), .B(y[5955]), .Z(n58490) );
  AND U37511 ( .A(n18409), .B(n58490), .Z(n18411) );
  NANDN U37512 ( .A(y[5956]), .B(x[5956]), .Z(n18410) );
  NANDN U37513 ( .A(y[5957]), .B(x[5957]), .Z(n23625) );
  NAND U37514 ( .A(n18410), .B(n23625), .Z(n58493) );
  OR U37515 ( .A(n18411), .B(n58493), .Z(n18412) );
  AND U37516 ( .A(n23626), .B(n18412), .Z(n18413) );
  NANDN U37517 ( .A(x[5957]), .B(y[5957]), .Z(n51222) );
  AND U37518 ( .A(n18413), .B(n51222), .Z(n18415) );
  NANDN U37519 ( .A(y[5958]), .B(x[5958]), .Z(n18414) );
  NANDN U37520 ( .A(y[5959]), .B(x[5959]), .Z(n23624) );
  NAND U37521 ( .A(n18414), .B(n23624), .Z(n58494) );
  OR U37522 ( .A(n18415), .B(n58494), .Z(n18416) );
  NAND U37523 ( .A(n58495), .B(n18416), .Z(n18417) );
  NANDN U37524 ( .A(y[5960]), .B(x[5960]), .Z(n23623) );
  NANDN U37525 ( .A(y[5961]), .B(x[5961]), .Z(n23619) );
  AND U37526 ( .A(n23623), .B(n23619), .Z(n51221) );
  AND U37527 ( .A(n18417), .B(n51221), .Z(n18418) );
  NOR U37528 ( .A(n23621), .B(n18418), .Z(n18419) );
  NAND U37529 ( .A(n23620), .B(n18419), .Z(n18420) );
  NANDN U37530 ( .A(n58498), .B(n18420), .Z(n18421) );
  AND U37531 ( .A(n23618), .B(n18421), .Z(n18422) );
  NANDN U37532 ( .A(x[5963]), .B(y[5963]), .Z(n51219) );
  NAND U37533 ( .A(n18422), .B(n51219), .Z(n18423) );
  NANDN U37534 ( .A(n58499), .B(n18423), .Z(n18424) );
  AND U37535 ( .A(n58500), .B(n18424), .Z(n18425) );
  OR U37536 ( .A(n58501), .B(n18425), .Z(n18426) );
  NAND U37537 ( .A(n58502), .B(n18426), .Z(n18427) );
  NANDN U37538 ( .A(n58503), .B(n18427), .Z(n18428) );
  AND U37539 ( .A(n23611), .B(n18428), .Z(n18429) );
  NANDN U37540 ( .A(x[5969]), .B(y[5969]), .Z(n51217) );
  AND U37541 ( .A(n18429), .B(n51217), .Z(n18431) );
  NANDN U37542 ( .A(y[5970]), .B(x[5970]), .Z(n18430) );
  NANDN U37543 ( .A(y[5971]), .B(x[5971]), .Z(n23608) );
  NAND U37544 ( .A(n18430), .B(n23608), .Z(n58504) );
  OR U37545 ( .A(n18431), .B(n58504), .Z(n18432) );
  AND U37546 ( .A(n23609), .B(n18432), .Z(n18433) );
  NANDN U37547 ( .A(x[5971]), .B(y[5971]), .Z(n58507) );
  AND U37548 ( .A(n18433), .B(n58507), .Z(n18434) );
  OR U37549 ( .A(n58510), .B(n18434), .Z(n18435) );
  NAND U37550 ( .A(n18436), .B(n18435), .Z(n18438) );
  NANDN U37551 ( .A(y[5974]), .B(x[5974]), .Z(n18437) );
  NANDN U37552 ( .A(y[5975]), .B(x[5975]), .Z(n23603) );
  AND U37553 ( .A(n18437), .B(n23603), .Z(n58513) );
  AND U37554 ( .A(n18438), .B(n58513), .Z(n18439) );
  NOR U37555 ( .A(n23605), .B(n18439), .Z(n18440) );
  NAND U37556 ( .A(n23604), .B(n18440), .Z(n18441) );
  NANDN U37557 ( .A(n58516), .B(n18441), .Z(n18442) );
  AND U37558 ( .A(n23602), .B(n18442), .Z(n18443) );
  NANDN U37559 ( .A(x[5977]), .B(y[5977]), .Z(n51215) );
  AND U37560 ( .A(n18443), .B(n51215), .Z(n18445) );
  NANDN U37561 ( .A(y[5978]), .B(x[5978]), .Z(n18444) );
  NANDN U37562 ( .A(y[5979]), .B(x[5979]), .Z(n23599) );
  AND U37563 ( .A(n18444), .B(n23599), .Z(n58517) );
  NANDN U37564 ( .A(n18445), .B(n58517), .Z(n18446) );
  NAND U37565 ( .A(n23600), .B(n18446), .Z(n18447) );
  NANDN U37566 ( .A(x[5979]), .B(y[5979]), .Z(n58519) );
  NANDN U37567 ( .A(n18447), .B(n58519), .Z(n18448) );
  NAND U37568 ( .A(n51214), .B(n18448), .Z(n18449) );
  NANDN U37569 ( .A(n45187), .B(n18449), .Z(n18450) );
  XNOR U37570 ( .A(x[5982]), .B(y[5982]), .Z(n23598) );
  NANDN U37571 ( .A(n18450), .B(n23598), .Z(n18452) );
  NANDN U37572 ( .A(y[5982]), .B(x[5982]), .Z(n18451) );
  NANDN U37573 ( .A(y[5983]), .B(x[5983]), .Z(n23595) );
  AND U37574 ( .A(n18451), .B(n23595), .Z(n58522) );
  AND U37575 ( .A(n18452), .B(n58522), .Z(n18453) );
  NOR U37576 ( .A(n58525), .B(n18453), .Z(n18454) );
  NAND U37577 ( .A(n23596), .B(n18454), .Z(n18455) );
  NANDN U37578 ( .A(n58528), .B(n18455), .Z(n18456) );
  AND U37579 ( .A(n23594), .B(n18456), .Z(n18457) );
  ANDN U37580 ( .B(y[5985]), .A(x[5985]), .Z(n51212) );
  ANDN U37581 ( .B(n18457), .A(n51212), .Z(n18459) );
  NANDN U37582 ( .A(y[5986]), .B(x[5986]), .Z(n18458) );
  NANDN U37583 ( .A(y[5987]), .B(x[5987]), .Z(n23591) );
  NAND U37584 ( .A(n18458), .B(n23591), .Z(n58529) );
  OR U37585 ( .A(n18459), .B(n58529), .Z(n18460) );
  AND U37586 ( .A(n23592), .B(n18460), .Z(n18461) );
  NANDN U37587 ( .A(x[5987]), .B(y[5987]), .Z(n58530) );
  AND U37588 ( .A(n18461), .B(n58530), .Z(n18463) );
  NANDN U37589 ( .A(y[5988]), .B(x[5988]), .Z(n18462) );
  NANDN U37590 ( .A(y[5989]), .B(x[5989]), .Z(n23589) );
  AND U37591 ( .A(n18462), .B(n23589), .Z(n51211) );
  NANDN U37592 ( .A(n18463), .B(n51211), .Z(n18464) );
  NAND U37593 ( .A(n18465), .B(n18464), .Z(n18467) );
  NANDN U37594 ( .A(y[5990]), .B(x[5990]), .Z(n18466) );
  NANDN U37595 ( .A(y[5991]), .B(x[5991]), .Z(n23586) );
  AND U37596 ( .A(n18466), .B(n23586), .Z(n58534) );
  AND U37597 ( .A(n18467), .B(n58534), .Z(n18468) );
  NOR U37598 ( .A(n23588), .B(n18468), .Z(n18469) );
  NAND U37599 ( .A(n23587), .B(n18469), .Z(n18470) );
  NANDN U37600 ( .A(n58537), .B(n18470), .Z(n18471) );
  AND U37601 ( .A(n23585), .B(n18471), .Z(n18472) );
  NANDN U37602 ( .A(x[5993]), .B(y[5993]), .Z(n51209) );
  AND U37603 ( .A(n18472), .B(n51209), .Z(n18474) );
  NANDN U37604 ( .A(y[5994]), .B(x[5994]), .Z(n18473) );
  NANDN U37605 ( .A(y[5995]), .B(x[5995]), .Z(n23582) );
  NAND U37606 ( .A(n18473), .B(n23582), .Z(n58539) );
  OR U37607 ( .A(n18474), .B(n58539), .Z(n18475) );
  AND U37608 ( .A(n23583), .B(n18475), .Z(n18476) );
  NAND U37609 ( .A(n58540), .B(n18476), .Z(n18477) );
  NAND U37610 ( .A(n51208), .B(n18477), .Z(n18478) );
  ANDN U37611 ( .B(y[5997]), .A(x[5997]), .Z(n45221) );
  ANDN U37612 ( .B(n18478), .A(n45221), .Z(n18479) );
  NAND U37613 ( .A(n23581), .B(n18479), .Z(n18481) );
  NANDN U37614 ( .A(y[5998]), .B(x[5998]), .Z(n18480) );
  NANDN U37615 ( .A(y[5999]), .B(x[5999]), .Z(n23578) );
  AND U37616 ( .A(n18480), .B(n23578), .Z(n58544) );
  AND U37617 ( .A(n18481), .B(n58544), .Z(n18482) );
  NOR U37618 ( .A(n45226), .B(n18482), .Z(n18483) );
  NAND U37619 ( .A(n23579), .B(n18483), .Z(n18484) );
  NANDN U37620 ( .A(n58547), .B(n18484), .Z(n18485) );
  AND U37621 ( .A(n23577), .B(n18485), .Z(n18486) );
  NANDN U37622 ( .A(x[6001]), .B(y[6001]), .Z(n51206) );
  AND U37623 ( .A(n18486), .B(n51206), .Z(n18488) );
  NANDN U37624 ( .A(y[6002]), .B(x[6002]), .Z(n18487) );
  NANDN U37625 ( .A(y[6003]), .B(x[6003]), .Z(n23574) );
  NAND U37626 ( .A(n18487), .B(n23574), .Z(n58548) );
  OR U37627 ( .A(n18488), .B(n58548), .Z(n18489) );
  AND U37628 ( .A(n23575), .B(n18489), .Z(n18490) );
  NANDN U37629 ( .A(x[6003]), .B(y[6003]), .Z(n58549) );
  AND U37630 ( .A(n18490), .B(n58549), .Z(n18492) );
  NANDN U37631 ( .A(y[6004]), .B(x[6004]), .Z(n18491) );
  NANDN U37632 ( .A(y[6005]), .B(x[6005]), .Z(n23572) );
  AND U37633 ( .A(n18491), .B(n23572), .Z(n51205) );
  NANDN U37634 ( .A(n18492), .B(n51205), .Z(n18493) );
  NAND U37635 ( .A(n18494), .B(n18493), .Z(n18496) );
  NANDN U37636 ( .A(y[6006]), .B(x[6006]), .Z(n18495) );
  NANDN U37637 ( .A(y[6007]), .B(x[6007]), .Z(n23570) );
  AND U37638 ( .A(n18495), .B(n23570), .Z(n58555) );
  AND U37639 ( .A(n18496), .B(n58555), .Z(n18497) );
  NOR U37640 ( .A(n45244), .B(n18497), .Z(n18498) );
  NAND U37641 ( .A(n23571), .B(n18498), .Z(n18499) );
  NANDN U37642 ( .A(n58558), .B(n18499), .Z(n18500) );
  AND U37643 ( .A(n23569), .B(n18500), .Z(n18501) );
  NANDN U37644 ( .A(x[6009]), .B(y[6009]), .Z(n51203) );
  AND U37645 ( .A(n18501), .B(n51203), .Z(n18503) );
  NANDN U37646 ( .A(y[6010]), .B(x[6010]), .Z(n18502) );
  NANDN U37647 ( .A(y[6011]), .B(x[6011]), .Z(n23566) );
  NAND U37648 ( .A(n18502), .B(n23566), .Z(n58559) );
  OR U37649 ( .A(n18503), .B(n58559), .Z(n18504) );
  AND U37650 ( .A(n23567), .B(n18504), .Z(n18505) );
  NANDN U37651 ( .A(x[6011]), .B(y[6011]), .Z(n58560) );
  AND U37652 ( .A(n18505), .B(n58560), .Z(n18507) );
  NANDN U37653 ( .A(y[6012]), .B(x[6012]), .Z(n18506) );
  NANDN U37654 ( .A(y[6013]), .B(x[6013]), .Z(n23564) );
  AND U37655 ( .A(n18506), .B(n23564), .Z(n51202) );
  NANDN U37656 ( .A(n18507), .B(n51202), .Z(n18508) );
  NAND U37657 ( .A(n18509), .B(n18508), .Z(n18511) );
  NANDN U37658 ( .A(y[6014]), .B(x[6014]), .Z(n18510) );
  NANDN U37659 ( .A(y[6015]), .B(x[6015]), .Z(n23562) );
  AND U37660 ( .A(n18510), .B(n23562), .Z(n58565) );
  AND U37661 ( .A(n18511), .B(n58565), .Z(n18512) );
  NOR U37662 ( .A(n45262), .B(n18512), .Z(n18513) );
  NAND U37663 ( .A(n23563), .B(n18513), .Z(n18514) );
  NANDN U37664 ( .A(n58568), .B(n18514), .Z(n18515) );
  AND U37665 ( .A(n23561), .B(n18515), .Z(n18516) );
  NANDN U37666 ( .A(x[6017]), .B(y[6017]), .Z(n51200) );
  AND U37667 ( .A(n18516), .B(n51200), .Z(n18518) );
  ANDN U37668 ( .B(x[6019]), .A(y[6019]), .Z(n45274) );
  NANDN U37669 ( .A(y[6018]), .B(x[6018]), .Z(n18517) );
  NANDN U37670 ( .A(n45274), .B(n18517), .Z(n58569) );
  OR U37671 ( .A(n18518), .B(n58569), .Z(n18519) );
  AND U37672 ( .A(n45275), .B(n18519), .Z(n18520) );
  NANDN U37673 ( .A(x[6019]), .B(y[6019]), .Z(n58571) );
  AND U37674 ( .A(n18520), .B(n58571), .Z(n18522) );
  NANDN U37675 ( .A(y[6020]), .B(x[6020]), .Z(n18521) );
  NANDN U37676 ( .A(y[6021]), .B(x[6021]), .Z(n23558) );
  NAND U37677 ( .A(n18521), .B(n23558), .Z(n58572) );
  OR U37678 ( .A(n18522), .B(n58572), .Z(n18523) );
  AND U37679 ( .A(n58573), .B(n18523), .Z(n18525) );
  NANDN U37680 ( .A(y[6022]), .B(x[6022]), .Z(n18524) );
  NANDN U37681 ( .A(y[6023]), .B(x[6023]), .Z(n23555) );
  NAND U37682 ( .A(n18524), .B(n23555), .Z(n58574) );
  OR U37683 ( .A(n18525), .B(n58574), .Z(n18526) );
  NAND U37684 ( .A(n18527), .B(n18526), .Z(n18528) );
  NANDN U37685 ( .A(n58575), .B(n18528), .Z(n18529) );
  AND U37686 ( .A(n23554), .B(n18529), .Z(n18530) );
  NANDN U37687 ( .A(x[6025]), .B(y[6025]), .Z(n58580) );
  AND U37688 ( .A(n18530), .B(n58580), .Z(n18532) );
  NANDN U37689 ( .A(y[6026]), .B(x[6026]), .Z(n18531) );
  NANDN U37690 ( .A(y[6027]), .B(x[6027]), .Z(n23551) );
  NAND U37691 ( .A(n18531), .B(n23551), .Z(n58581) );
  OR U37692 ( .A(n18532), .B(n58581), .Z(n18533) );
  AND U37693 ( .A(n23552), .B(n18533), .Z(n18534) );
  NANDN U37694 ( .A(x[6027]), .B(y[6027]), .Z(n58582) );
  AND U37695 ( .A(n18534), .B(n58582), .Z(n18536) );
  NANDN U37696 ( .A(y[6028]), .B(x[6028]), .Z(n18535) );
  NANDN U37697 ( .A(y[6029]), .B(x[6029]), .Z(n23549) );
  NAND U37698 ( .A(n18535), .B(n23549), .Z(n58584) );
  OR U37699 ( .A(n18536), .B(n58584), .Z(n18537) );
  AND U37700 ( .A(n18538), .B(n18537), .Z(n18540) );
  NANDN U37701 ( .A(y[6030]), .B(x[6030]), .Z(n18539) );
  ANDN U37702 ( .B(x[6031]), .A(y[6031]), .Z(n45301) );
  ANDN U37703 ( .B(n18539), .A(n45301), .Z(n58587) );
  NANDN U37704 ( .A(n18540), .B(n58587), .Z(n18541) );
  AND U37705 ( .A(n45302), .B(n18541), .Z(n18542) );
  NANDN U37706 ( .A(x[6031]), .B(y[6031]), .Z(n51196) );
  NAND U37707 ( .A(n18542), .B(n51196), .Z(n18543) );
  AND U37708 ( .A(n58588), .B(n18543), .Z(n18544) );
  ANDN U37709 ( .B(n58590), .A(n18544), .Z(n18545) );
  NAND U37710 ( .A(n23548), .B(n18545), .Z(n18546) );
  NANDN U37711 ( .A(n58591), .B(n18546), .Z(n18547) );
  AND U37712 ( .A(n23545), .B(n18547), .Z(n18548) );
  NANDN U37713 ( .A(n23546), .B(n18548), .Z(n18549) );
  NAND U37714 ( .A(n58594), .B(n18549), .Z(n18550) );
  NANDN U37715 ( .A(n58595), .B(n18550), .Z(n18551) );
  AND U37716 ( .A(n58596), .B(n18551), .Z(n18552) );
  ANDN U37717 ( .B(n58598), .A(n18552), .Z(n18553) );
  NAND U37718 ( .A(n45322), .B(n18553), .Z(n18554) );
  NANDN U37719 ( .A(n58599), .B(n18554), .Z(n18555) );
  AND U37720 ( .A(n23542), .B(n18555), .Z(n18556) );
  NANDN U37721 ( .A(x[6041]), .B(y[6041]), .Z(n58600) );
  NAND U37722 ( .A(n18556), .B(n58600), .Z(n18557) );
  NANDN U37723 ( .A(n58602), .B(n18557), .Z(n18558) );
  AND U37724 ( .A(n23540), .B(n18558), .Z(n18559) );
  NANDN U37725 ( .A(x[6043]), .B(y[6043]), .Z(n58603) );
  AND U37726 ( .A(n18559), .B(n58603), .Z(n18560) );
  OR U37727 ( .A(n58605), .B(n18560), .Z(n18561) );
  NAND U37728 ( .A(n18562), .B(n18561), .Z(n18563) );
  AND U37729 ( .A(n58606), .B(n18563), .Z(n18565) );
  XNOR U37730 ( .A(x[6048]), .B(y[6048]), .Z(n23536) );
  NANDN U37731 ( .A(x[6047]), .B(y[6047]), .Z(n58608) );
  AND U37732 ( .A(n23536), .B(n58608), .Z(n18564) );
  NANDN U37733 ( .A(n18565), .B(n18564), .Z(n18566) );
  AND U37734 ( .A(n58609), .B(n18566), .Z(n18567) );
  OR U37735 ( .A(n58610), .B(n18567), .Z(n18568) );
  NAND U37736 ( .A(n58612), .B(n18568), .Z(n18569) );
  NANDN U37737 ( .A(n58613), .B(n18569), .Z(n18570) );
  AND U37738 ( .A(n58614), .B(n18570), .Z(n18571) );
  NANDN U37739 ( .A(x[6053]), .B(y[6053]), .Z(n23527) );
  NANDN U37740 ( .A(x[6054]), .B(y[6054]), .Z(n23524) );
  AND U37741 ( .A(n23527), .B(n23524), .Z(n58615) );
  NANDN U37742 ( .A(n18571), .B(n58615), .Z(n18572) );
  NANDN U37743 ( .A(n58616), .B(n18572), .Z(n18573) );
  AND U37744 ( .A(n58617), .B(n18573), .Z(n18574) );
  NAND U37745 ( .A(n23523), .B(n18574), .Z(n18575) );
  NANDN U37746 ( .A(n58619), .B(n18575), .Z(n18576) );
  AND U37747 ( .A(n18577), .B(n18576), .Z(n18578) );
  OR U37748 ( .A(n58620), .B(n18578), .Z(n18579) );
  NAND U37749 ( .A(n58621), .B(n18579), .Z(n18580) );
  NANDN U37750 ( .A(n58622), .B(n18580), .Z(n18581) );
  AND U37751 ( .A(n58623), .B(n18581), .Z(n18582) );
  NANDN U37752 ( .A(y[6062]), .B(x[6062]), .Z(n23514) );
  NANDN U37753 ( .A(y[6063]), .B(x[6063]), .Z(n23511) );
  NAND U37754 ( .A(n23514), .B(n23511), .Z(n58624) );
  OR U37755 ( .A(n18582), .B(n58624), .Z(n18583) );
  AND U37756 ( .A(n18584), .B(n18583), .Z(n18585) );
  OR U37757 ( .A(n58625), .B(n18585), .Z(n18586) );
  NAND U37758 ( .A(n58627), .B(n18586), .Z(n18587) );
  NANDN U37759 ( .A(n58628), .B(n18587), .Z(n18588) );
  AND U37760 ( .A(n58629), .B(n18588), .Z(n18589) );
  NANDN U37761 ( .A(y[6068]), .B(x[6068]), .Z(n23505) );
  NANDN U37762 ( .A(y[6069]), .B(x[6069]), .Z(n23501) );
  AND U37763 ( .A(n23505), .B(n23501), .Z(n58630) );
  NANDN U37764 ( .A(n18589), .B(n58630), .Z(n18590) );
  NAND U37765 ( .A(n18591), .B(n18590), .Z(n18592) );
  AND U37766 ( .A(n58631), .B(n18592), .Z(n18593) );
  ANDN U37767 ( .B(n58633), .A(n18593), .Z(n18594) );
  NAND U37768 ( .A(n23500), .B(n18594), .Z(n18595) );
  NANDN U37769 ( .A(n58634), .B(n18595), .Z(n18596) );
  AND U37770 ( .A(n23498), .B(n18596), .Z(n18597) );
  NANDN U37771 ( .A(x[6073]), .B(y[6073]), .Z(n58635) );
  AND U37772 ( .A(n18597), .B(n58635), .Z(n18599) );
  NANDN U37773 ( .A(y[6074]), .B(x[6074]), .Z(n18598) );
  NANDN U37774 ( .A(y[6075]), .B(x[6075]), .Z(n23494) );
  AND U37775 ( .A(n18598), .B(n23494), .Z(n58637) );
  NANDN U37776 ( .A(n18599), .B(n58637), .Z(n18600) );
  NAND U37777 ( .A(n23495), .B(n18600), .Z(n18601) );
  ANDN U37778 ( .B(y[6075]), .A(x[6075]), .Z(n23496) );
  OR U37779 ( .A(n18601), .B(n23496), .Z(n18602) );
  NAND U37780 ( .A(n58640), .B(n18602), .Z(n18604) );
  XNOR U37781 ( .A(x[6078]), .B(y[6078]), .Z(n23493) );
  NANDN U37782 ( .A(x[6077]), .B(y[6077]), .Z(n51185) );
  NAND U37783 ( .A(n23493), .B(n51185), .Z(n18603) );
  ANDN U37784 ( .B(n18604), .A(n18603), .Z(n18606) );
  NANDN U37785 ( .A(y[6078]), .B(x[6078]), .Z(n18605) );
  NANDN U37786 ( .A(y[6079]), .B(x[6079]), .Z(n23490) );
  NAND U37787 ( .A(n18605), .B(n23490), .Z(n58643) );
  OR U37788 ( .A(n18606), .B(n58643), .Z(n18607) );
  NAND U37789 ( .A(n18608), .B(n18607), .Z(n18609) );
  NANDN U37790 ( .A(n58647), .B(n18609), .Z(n18610) );
  AND U37791 ( .A(n23489), .B(n18610), .Z(n18611) );
  NANDN U37792 ( .A(x[6081]), .B(y[6081]), .Z(n58648) );
  NAND U37793 ( .A(n18611), .B(n58648), .Z(n18612) );
  NANDN U37794 ( .A(n58650), .B(n18612), .Z(n18613) );
  AND U37795 ( .A(n23487), .B(n18613), .Z(n18614) );
  NANDN U37796 ( .A(x[6083]), .B(y[6083]), .Z(n58651) );
  AND U37797 ( .A(n18614), .B(n58651), .Z(n18615) );
  OR U37798 ( .A(n58653), .B(n18615), .Z(n18616) );
  NAND U37799 ( .A(n18617), .B(n18616), .Z(n18618) );
  AND U37800 ( .A(n58654), .B(n18618), .Z(n18619) );
  ANDN U37801 ( .B(n58656), .A(n18619), .Z(n18620) );
  NAND U37802 ( .A(n23483), .B(n18620), .Z(n18621) );
  NANDN U37803 ( .A(n58657), .B(n18621), .Z(n18622) );
  AND U37804 ( .A(n23481), .B(n18622), .Z(n18623) );
  NANDN U37805 ( .A(x[6089]), .B(y[6089]), .Z(n58658) );
  NAND U37806 ( .A(n18623), .B(n58658), .Z(n18624) );
  NANDN U37807 ( .A(n58660), .B(n18624), .Z(n18625) );
  AND U37808 ( .A(n23479), .B(n18625), .Z(n18626) );
  NANDN U37809 ( .A(x[6091]), .B(y[6091]), .Z(n58662) );
  AND U37810 ( .A(n18626), .B(n58662), .Z(n18627) );
  OR U37811 ( .A(n58664), .B(n18627), .Z(n18628) );
  NAND U37812 ( .A(n18629), .B(n18628), .Z(n18630) );
  AND U37813 ( .A(n58665), .B(n18630), .Z(n18631) );
  ANDN U37814 ( .B(n51179), .A(n18631), .Z(n18632) );
  NAND U37815 ( .A(n45439), .B(n18632), .Z(n18633) );
  NANDN U37816 ( .A(n51178), .B(n18633), .Z(n18634) );
  AND U37817 ( .A(n23475), .B(n18634), .Z(n18635) );
  NANDN U37818 ( .A(x[6097]), .B(y[6097]), .Z(n58666) );
  NAND U37819 ( .A(n18635), .B(n58666), .Z(n18636) );
  NANDN U37820 ( .A(n58668), .B(n18636), .Z(n18637) );
  AND U37821 ( .A(n23473), .B(n18637), .Z(n18638) );
  NANDN U37822 ( .A(x[6099]), .B(y[6099]), .Z(n58669) );
  AND U37823 ( .A(n18638), .B(n58669), .Z(n18639) );
  OR U37824 ( .A(n58671), .B(n18639), .Z(n18640) );
  NAND U37825 ( .A(n18641), .B(n18640), .Z(n18642) );
  AND U37826 ( .A(n58672), .B(n18642), .Z(n18643) );
  ANDN U37827 ( .B(n58674), .A(n18643), .Z(n18644) );
  NAND U37828 ( .A(n23469), .B(n18644), .Z(n18645) );
  NANDN U37829 ( .A(n58677), .B(n18645), .Z(n18646) );
  AND U37830 ( .A(n23467), .B(n18646), .Z(n18647) );
  NANDN U37831 ( .A(x[6105]), .B(y[6105]), .Z(n58678) );
  NAND U37832 ( .A(n18647), .B(n58678), .Z(n18648) );
  NANDN U37833 ( .A(n51175), .B(n18648), .Z(n18649) );
  AND U37834 ( .A(n23465), .B(n18649), .Z(n18650) );
  NANDN U37835 ( .A(x[6107]), .B(y[6107]), .Z(n58680) );
  AND U37836 ( .A(n18650), .B(n58680), .Z(n18652) );
  NANDN U37837 ( .A(y[6108]), .B(x[6108]), .Z(n18651) );
  NANDN U37838 ( .A(y[6109]), .B(x[6109]), .Z(n23462) );
  AND U37839 ( .A(n18651), .B(n23462), .Z(n58682) );
  NANDN U37840 ( .A(n18652), .B(n58682), .Z(n18653) );
  NAND U37841 ( .A(n18654), .B(n18653), .Z(n18655) );
  AND U37842 ( .A(n58683), .B(n18655), .Z(n18656) );
  ANDN U37843 ( .B(n58685), .A(n18656), .Z(n18657) );
  NAND U37844 ( .A(n23461), .B(n18657), .Z(n18658) );
  NANDN U37845 ( .A(n58686), .B(n18658), .Z(n18659) );
  AND U37846 ( .A(n23459), .B(n18659), .Z(n18660) );
  NANDN U37847 ( .A(x[6113]), .B(y[6113]), .Z(n58687) );
  AND U37848 ( .A(n18660), .B(n58687), .Z(n18662) );
  NANDN U37849 ( .A(y[6114]), .B(x[6114]), .Z(n18661) );
  NANDN U37850 ( .A(y[6115]), .B(x[6115]), .Z(n23456) );
  NAND U37851 ( .A(n18661), .B(n23456), .Z(n58689) );
  OR U37852 ( .A(n18662), .B(n58689), .Z(n18663) );
  AND U37853 ( .A(n23457), .B(n18663), .Z(n18664) );
  NANDN U37854 ( .A(x[6115]), .B(y[6115]), .Z(n58691) );
  AND U37855 ( .A(n18664), .B(n58691), .Z(n18665) );
  OR U37856 ( .A(n58693), .B(n18665), .Z(n18666) );
  NAND U37857 ( .A(n18667), .B(n18666), .Z(n18668) );
  AND U37858 ( .A(n58694), .B(n18668), .Z(n18669) );
  ANDN U37859 ( .B(n58696), .A(n18669), .Z(n18670) );
  NAND U37860 ( .A(n23453), .B(n18670), .Z(n18671) );
  NANDN U37861 ( .A(n58697), .B(n18671), .Z(n18672) );
  AND U37862 ( .A(n23451), .B(n18672), .Z(n18673) );
  NANDN U37863 ( .A(x[6121]), .B(y[6121]), .Z(n58698) );
  AND U37864 ( .A(n18673), .B(n58698), .Z(n18675) );
  NANDN U37865 ( .A(y[6122]), .B(x[6122]), .Z(n18674) );
  ANDN U37866 ( .B(x[6123]), .A(y[6123]), .Z(n45499) );
  ANDN U37867 ( .B(n18674), .A(n45499), .Z(n58700) );
  NANDN U37868 ( .A(n18675), .B(n58700), .Z(n18676) );
  AND U37869 ( .A(n58701), .B(n18676), .Z(n18678) );
  NANDN U37870 ( .A(y[6124]), .B(x[6124]), .Z(n18677) );
  NANDN U37871 ( .A(y[6125]), .B(x[6125]), .Z(n23448) );
  AND U37872 ( .A(n18677), .B(n23448), .Z(n58702) );
  NANDN U37873 ( .A(n18678), .B(n58702), .Z(n18679) );
  NAND U37874 ( .A(n18680), .B(n18679), .Z(n18682) );
  NANDN U37875 ( .A(y[6126]), .B(x[6126]), .Z(n18681) );
  NANDN U37876 ( .A(y[6127]), .B(x[6127]), .Z(n23446) );
  AND U37877 ( .A(n18681), .B(n23446), .Z(n51170) );
  AND U37878 ( .A(n18682), .B(n51170), .Z(n18683) );
  NOR U37879 ( .A(n45507), .B(n18683), .Z(n18684) );
  NAND U37880 ( .A(n23447), .B(n18684), .Z(n18685) );
  NANDN U37881 ( .A(n58707), .B(n18685), .Z(n18686) );
  AND U37882 ( .A(n23445), .B(n18686), .Z(n18687) );
  NANDN U37883 ( .A(x[6129]), .B(y[6129]), .Z(n58709) );
  AND U37884 ( .A(n18687), .B(n58709), .Z(n18688) );
  OR U37885 ( .A(n58711), .B(n18688), .Z(n18689) );
  AND U37886 ( .A(n23443), .B(n18689), .Z(n18690) );
  NANDN U37887 ( .A(x[6131]), .B(y[6131]), .Z(n51168) );
  AND U37888 ( .A(n18690), .B(n51168), .Z(n18692) );
  NANDN U37889 ( .A(y[6132]), .B(x[6132]), .Z(n18691) );
  NANDN U37890 ( .A(y[6133]), .B(x[6133]), .Z(n23440) );
  AND U37891 ( .A(n18691), .B(n23440), .Z(n58712) );
  NANDN U37892 ( .A(n18692), .B(n58712), .Z(n18693) );
  NAND U37893 ( .A(n18694), .B(n18693), .Z(n18696) );
  NANDN U37894 ( .A(y[6134]), .B(x[6134]), .Z(n18695) );
  NANDN U37895 ( .A(y[6135]), .B(x[6135]), .Z(n23438) );
  AND U37896 ( .A(n18695), .B(n23438), .Z(n51167) );
  AND U37897 ( .A(n18696), .B(n51167), .Z(n18697) );
  NOR U37898 ( .A(n45524), .B(n18697), .Z(n18698) );
  NAND U37899 ( .A(n23439), .B(n18698), .Z(n18699) );
  NANDN U37900 ( .A(n58717), .B(n18699), .Z(n18700) );
  AND U37901 ( .A(n23437), .B(n18700), .Z(n18701) );
  NANDN U37902 ( .A(n45529), .B(n18701), .Z(n18702) );
  NAND U37903 ( .A(n58720), .B(n18702), .Z(n18703) );
  NAND U37904 ( .A(n58721), .B(n18703), .Z(n18704) );
  AND U37905 ( .A(n58722), .B(n18704), .Z(n18705) );
  NOR U37906 ( .A(n58724), .B(n18705), .Z(n18706) );
  NAND U37907 ( .A(n23432), .B(n18706), .Z(n18707) );
  NANDN U37908 ( .A(n58727), .B(n18707), .Z(n18708) );
  AND U37909 ( .A(n23430), .B(n18708), .Z(n18709) );
  ANDN U37910 ( .B(y[6143]), .A(x[6143]), .Z(n58728) );
  ANDN U37911 ( .B(n18709), .A(n58728), .Z(n18711) );
  NANDN U37912 ( .A(y[6144]), .B(x[6144]), .Z(n18710) );
  NANDN U37913 ( .A(y[6145]), .B(x[6145]), .Z(n23427) );
  AND U37914 ( .A(n18710), .B(n23427), .Z(n58729) );
  NANDN U37915 ( .A(n18711), .B(n58729), .Z(n18712) );
  NANDN U37916 ( .A(x[6145]), .B(y[6145]), .Z(n23428) );
  NANDN U37917 ( .A(x[6146]), .B(y[6146]), .Z(n23425) );
  AND U37918 ( .A(n23428), .B(n23425), .Z(n51165) );
  AND U37919 ( .A(n18712), .B(n51165), .Z(n18713) );
  NANDN U37920 ( .A(y[6146]), .B(x[6146]), .Z(n23426) );
  NANDN U37921 ( .A(y[6147]), .B(x[6147]), .Z(n23423) );
  AND U37922 ( .A(n23426), .B(n23423), .Z(n58730) );
  NANDN U37923 ( .A(n18713), .B(n58730), .Z(n18714) );
  NAND U37924 ( .A(n18715), .B(n18714), .Z(n18717) );
  NANDN U37925 ( .A(y[6148]), .B(x[6148]), .Z(n18716) );
  NANDN U37926 ( .A(y[6149]), .B(x[6149]), .Z(n23421) );
  AND U37927 ( .A(n18716), .B(n23421), .Z(n51164) );
  AND U37928 ( .A(n18717), .B(n51164), .Z(n18718) );
  NOR U37929 ( .A(n58733), .B(n18718), .Z(n18719) );
  NAND U37930 ( .A(n23422), .B(n18719), .Z(n18720) );
  NANDN U37931 ( .A(n58735), .B(n18720), .Z(n18721) );
  AND U37932 ( .A(n45562), .B(n18721), .Z(n18722) );
  NANDN U37933 ( .A(x[6151]), .B(y[6151]), .Z(n58736) );
  AND U37934 ( .A(n18722), .B(n58736), .Z(n18723) );
  OR U37935 ( .A(n58739), .B(n18723), .Z(n18724) );
  AND U37936 ( .A(n23420), .B(n18724), .Z(n18725) );
  ANDN U37937 ( .B(y[6153]), .A(x[6153]), .Z(n51162) );
  ANDN U37938 ( .B(n18725), .A(n51162), .Z(n18727) );
  NANDN U37939 ( .A(y[6154]), .B(x[6154]), .Z(n18726) );
  NANDN U37940 ( .A(y[6155]), .B(x[6155]), .Z(n45571) );
  AND U37941 ( .A(n18726), .B(n45571), .Z(n58740) );
  NANDN U37942 ( .A(n18727), .B(n58740), .Z(n18728) );
  NAND U37943 ( .A(n18729), .B(n18728), .Z(n18731) );
  NANDN U37944 ( .A(y[6156]), .B(x[6156]), .Z(n18730) );
  NANDN U37945 ( .A(y[6157]), .B(x[6157]), .Z(n23417) );
  AND U37946 ( .A(n18730), .B(n23417), .Z(n51161) );
  AND U37947 ( .A(n18731), .B(n51161), .Z(n18732) );
  NOR U37948 ( .A(n58743), .B(n18732), .Z(n18733) );
  NAND U37949 ( .A(n23418), .B(n18733), .Z(n18734) );
  NANDN U37950 ( .A(n58745), .B(n18734), .Z(n18735) );
  AND U37951 ( .A(n45582), .B(n18735), .Z(n18736) );
  NANDN U37952 ( .A(x[6159]), .B(y[6159]), .Z(n58746) );
  AND U37953 ( .A(n18736), .B(n58746), .Z(n18738) );
  NANDN U37954 ( .A(y[6160]), .B(x[6160]), .Z(n18737) );
  NANDN U37955 ( .A(y[6161]), .B(x[6161]), .Z(n23415) );
  NAND U37956 ( .A(n18737), .B(n23415), .Z(n58748) );
  OR U37957 ( .A(n18738), .B(n58748), .Z(n18739) );
  AND U37958 ( .A(n23416), .B(n18739), .Z(n18740) );
  ANDN U37959 ( .B(y[6161]), .A(x[6161]), .Z(n51159) );
  ANDN U37960 ( .B(n18740), .A(n51159), .Z(n18742) );
  NANDN U37961 ( .A(y[6162]), .B(x[6162]), .Z(n18741) );
  NANDN U37962 ( .A(y[6163]), .B(x[6163]), .Z(n23414) );
  NAND U37963 ( .A(n18741), .B(n23414), .Z(n58749) );
  OR U37964 ( .A(n18742), .B(n58749), .Z(n18743) );
  AND U37965 ( .A(n58750), .B(n18743), .Z(n18744) );
  OR U37966 ( .A(n58752), .B(n18744), .Z(n18745) );
  NAND U37967 ( .A(n18746), .B(n18745), .Z(n18747) );
  NANDN U37968 ( .A(n51158), .B(n18747), .Z(n18748) );
  NANDN U37969 ( .A(x[6167]), .B(y[6167]), .Z(n23409) );
  NANDN U37970 ( .A(x[6168]), .B(y[6168]), .Z(n23406) );
  AND U37971 ( .A(n23409), .B(n23406), .Z(n51157) );
  AND U37972 ( .A(n18748), .B(n51157), .Z(n18749) );
  NANDN U37973 ( .A(y[6168]), .B(x[6168]), .Z(n23407) );
  NANDN U37974 ( .A(y[6169]), .B(x[6169]), .Z(n23404) );
  AND U37975 ( .A(n23407), .B(n23404), .Z(n58755) );
  NANDN U37976 ( .A(n18749), .B(n58755), .Z(n18750) );
  NAND U37977 ( .A(n18751), .B(n18750), .Z(n18753) );
  NANDN U37978 ( .A(y[6170]), .B(x[6170]), .Z(n18752) );
  NANDN U37979 ( .A(y[6171]), .B(x[6171]), .Z(n23401) );
  AND U37980 ( .A(n18752), .B(n23401), .Z(n51156) );
  AND U37981 ( .A(n18753), .B(n51156), .Z(n18754) );
  NOR U37982 ( .A(n23403), .B(n18754), .Z(n18755) );
  NAND U37983 ( .A(n23402), .B(n18755), .Z(n18756) );
  NANDN U37984 ( .A(n58760), .B(n18756), .Z(n18757) );
  AND U37985 ( .A(n23400), .B(n18757), .Z(n18758) );
  NANDN U37986 ( .A(x[6173]), .B(y[6173]), .Z(n58761) );
  AND U37987 ( .A(n18758), .B(n58761), .Z(n18760) );
  NANDN U37988 ( .A(y[6174]), .B(x[6174]), .Z(n18759) );
  NANDN U37989 ( .A(y[6175]), .B(x[6175]), .Z(n45616) );
  NAND U37990 ( .A(n18759), .B(n45616), .Z(n58763) );
  OR U37991 ( .A(n18760), .B(n58763), .Z(n18761) );
  AND U37992 ( .A(n51155), .B(n18761), .Z(n18762) );
  NAND U37993 ( .A(n45617), .B(n18762), .Z(n18763) );
  NANDN U37994 ( .A(n58766), .B(n18763), .Z(n18764) );
  AND U37995 ( .A(n23398), .B(n18764), .Z(n18765) );
  NAND U37996 ( .A(n58770), .B(n18765), .Z(n18767) );
  NANDN U37997 ( .A(y[6178]), .B(x[6178]), .Z(n18766) );
  NANDN U37998 ( .A(y[6179]), .B(x[6179]), .Z(n45627) );
  AND U37999 ( .A(n18766), .B(n45627), .Z(n51153) );
  AND U38000 ( .A(n18767), .B(n51153), .Z(n18768) );
  NOR U38001 ( .A(n45624), .B(n18768), .Z(n18769) );
  NAND U38002 ( .A(n45628), .B(n18769), .Z(n18770) );
  NANDN U38003 ( .A(n58773), .B(n18770), .Z(n18771) );
  AND U38004 ( .A(n23396), .B(n18771), .Z(n18772) );
  ANDN U38005 ( .B(y[6181]), .A(x[6181]), .Z(n58774) );
  ANDN U38006 ( .B(n18772), .A(n58774), .Z(n18773) );
  OR U38007 ( .A(n58776), .B(n18773), .Z(n18774) );
  AND U38008 ( .A(n45638), .B(n18774), .Z(n18775) );
  NANDN U38009 ( .A(x[6183]), .B(y[6183]), .Z(n51152) );
  AND U38010 ( .A(n18775), .B(n51152), .Z(n18777) );
  NANDN U38011 ( .A(y[6184]), .B(x[6184]), .Z(n18776) );
  NANDN U38012 ( .A(y[6185]), .B(x[6185]), .Z(n23393) );
  AND U38013 ( .A(n18776), .B(n23393), .Z(n58777) );
  NANDN U38014 ( .A(n18777), .B(n58777), .Z(n18778) );
  NAND U38015 ( .A(n18779), .B(n18778), .Z(n18781) );
  NANDN U38016 ( .A(y[6186]), .B(x[6186]), .Z(n18780) );
  NANDN U38017 ( .A(y[6187]), .B(x[6187]), .Z(n45648) );
  AND U38018 ( .A(n18780), .B(n45648), .Z(n51150) );
  AND U38019 ( .A(n18781), .B(n51150), .Z(n18782) );
  NOR U38020 ( .A(n45645), .B(n18782), .Z(n18783) );
  NAND U38021 ( .A(n45649), .B(n18783), .Z(n18784) );
  NANDN U38022 ( .A(n58783), .B(n18784), .Z(n18785) );
  AND U38023 ( .A(n23392), .B(n18785), .Z(n18786) );
  ANDN U38024 ( .B(y[6189]), .A(x[6189]), .Z(n58784) );
  ANDN U38025 ( .B(n18786), .A(n58784), .Z(n18788) );
  NANDN U38026 ( .A(y[6190]), .B(x[6190]), .Z(n18787) );
  NANDN U38027 ( .A(y[6191]), .B(x[6191]), .Z(n45658) );
  NAND U38028 ( .A(n18787), .B(n45658), .Z(n58786) );
  OR U38029 ( .A(n18788), .B(n58786), .Z(n18789) );
  AND U38030 ( .A(n45659), .B(n18789), .Z(n18790) );
  NANDN U38031 ( .A(x[6191]), .B(y[6191]), .Z(n51149) );
  AND U38032 ( .A(n18790), .B(n51149), .Z(n18792) );
  NANDN U38033 ( .A(y[6192]), .B(x[6192]), .Z(n18791) );
  NANDN U38034 ( .A(y[6193]), .B(x[6193]), .Z(n23389) );
  AND U38035 ( .A(n18791), .B(n23389), .Z(n58787) );
  NANDN U38036 ( .A(n18792), .B(n58787), .Z(n18793) );
  NAND U38037 ( .A(n18794), .B(n18793), .Z(n18796) );
  NANDN U38038 ( .A(y[6194]), .B(x[6194]), .Z(n18795) );
  NANDN U38039 ( .A(y[6195]), .B(x[6195]), .Z(n45669) );
  AND U38040 ( .A(n18795), .B(n45669), .Z(n51147) );
  AND U38041 ( .A(n18796), .B(n51147), .Z(n18797) );
  NOR U38042 ( .A(n45666), .B(n18797), .Z(n18798) );
  NAND U38043 ( .A(n45670), .B(n18798), .Z(n18799) );
  NANDN U38044 ( .A(n51146), .B(n18799), .Z(n18800) );
  AND U38045 ( .A(n23387), .B(n18800), .Z(n18801) );
  NANDN U38046 ( .A(x[6197]), .B(y[6197]), .Z(n23388) );
  AND U38047 ( .A(n18801), .B(n23388), .Z(n18803) );
  NANDN U38048 ( .A(y[6198]), .B(x[6198]), .Z(n18802) );
  NANDN U38049 ( .A(y[6199]), .B(x[6199]), .Z(n45679) );
  NAND U38050 ( .A(n18802), .B(n45679), .Z(n58795) );
  OR U38051 ( .A(n18803), .B(n58795), .Z(n18804) );
  AND U38052 ( .A(n45680), .B(n18804), .Z(n18805) );
  NANDN U38053 ( .A(x[6199]), .B(y[6199]), .Z(n51145) );
  AND U38054 ( .A(n18805), .B(n51145), .Z(n18807) );
  NANDN U38055 ( .A(y[6200]), .B(x[6200]), .Z(n18806) );
  NANDN U38056 ( .A(y[6201]), .B(x[6201]), .Z(n23384) );
  AND U38057 ( .A(n18806), .B(n23384), .Z(n58796) );
  NANDN U38058 ( .A(n18807), .B(n58796), .Z(n18808) );
  NAND U38059 ( .A(n18809), .B(n18808), .Z(n18811) );
  NANDN U38060 ( .A(y[6202]), .B(x[6202]), .Z(n18810) );
  NANDN U38061 ( .A(y[6203]), .B(x[6203]), .Z(n45690) );
  AND U38062 ( .A(n18810), .B(n45690), .Z(n51143) );
  AND U38063 ( .A(n18811), .B(n51143), .Z(n18812) );
  NOR U38064 ( .A(n45687), .B(n18812), .Z(n18813) );
  NAND U38065 ( .A(n45691), .B(n18813), .Z(n18814) );
  NANDN U38066 ( .A(n51142), .B(n18814), .Z(n18815) );
  AND U38067 ( .A(n23382), .B(n18815), .Z(n18816) );
  NANDN U38068 ( .A(x[6205]), .B(y[6205]), .Z(n23383) );
  AND U38069 ( .A(n18816), .B(n23383), .Z(n18818) );
  NANDN U38070 ( .A(y[6206]), .B(x[6206]), .Z(n18817) );
  NANDN U38071 ( .A(y[6207]), .B(x[6207]), .Z(n45700) );
  NAND U38072 ( .A(n18817), .B(n45700), .Z(n58803) );
  OR U38073 ( .A(n18818), .B(n58803), .Z(n18819) );
  AND U38074 ( .A(n45701), .B(n18819), .Z(n18820) );
  NANDN U38075 ( .A(x[6207]), .B(y[6207]), .Z(n51141) );
  AND U38076 ( .A(n18820), .B(n51141), .Z(n18822) );
  NANDN U38077 ( .A(y[6208]), .B(x[6208]), .Z(n18821) );
  NANDN U38078 ( .A(y[6209]), .B(x[6209]), .Z(n23379) );
  AND U38079 ( .A(n18821), .B(n23379), .Z(n58805) );
  NANDN U38080 ( .A(n18822), .B(n58805), .Z(n18823) );
  NAND U38081 ( .A(n18824), .B(n18823), .Z(n18826) );
  NANDN U38082 ( .A(y[6210]), .B(x[6210]), .Z(n18825) );
  NANDN U38083 ( .A(y[6211]), .B(x[6211]), .Z(n45711) );
  AND U38084 ( .A(n18825), .B(n45711), .Z(n51138) );
  AND U38085 ( .A(n18826), .B(n51138), .Z(n18827) );
  NOR U38086 ( .A(n45708), .B(n18827), .Z(n18828) );
  NAND U38087 ( .A(n45712), .B(n18828), .Z(n18829) );
  NANDN U38088 ( .A(n58809), .B(n18829), .Z(n18830) );
  AND U38089 ( .A(n23378), .B(n18830), .Z(n18831) );
  NANDN U38090 ( .A(n58810), .B(n18831), .Z(n18832) );
  NAND U38091 ( .A(n58812), .B(n18832), .Z(n18833) );
  AND U38092 ( .A(n45722), .B(n18833), .Z(n18834) );
  NANDN U38093 ( .A(x[6215]), .B(y[6215]), .Z(n51137) );
  AND U38094 ( .A(n18834), .B(n51137), .Z(n18836) );
  NANDN U38095 ( .A(y[6216]), .B(x[6216]), .Z(n18835) );
  NANDN U38096 ( .A(y[6217]), .B(x[6217]), .Z(n23375) );
  AND U38097 ( .A(n18835), .B(n23375), .Z(n58814) );
  NANDN U38098 ( .A(n18836), .B(n58814), .Z(n18837) );
  NAND U38099 ( .A(n18838), .B(n18837), .Z(n18840) );
  NANDN U38100 ( .A(y[6218]), .B(x[6218]), .Z(n18839) );
  NANDN U38101 ( .A(y[6219]), .B(x[6219]), .Z(n45732) );
  AND U38102 ( .A(n18839), .B(n45732), .Z(n51135) );
  AND U38103 ( .A(n18840), .B(n51135), .Z(n18841) );
  NOR U38104 ( .A(n45729), .B(n18841), .Z(n18842) );
  NAND U38105 ( .A(n45733), .B(n18842), .Z(n18843) );
  NANDN U38106 ( .A(n58820), .B(n18843), .Z(n18844) );
  AND U38107 ( .A(n23374), .B(n18844), .Z(n18845) );
  ANDN U38108 ( .B(y[6221]), .A(x[6221]), .Z(n58821) );
  ANDN U38109 ( .B(n18845), .A(n58821), .Z(n18847) );
  NANDN U38110 ( .A(y[6222]), .B(x[6222]), .Z(n18846) );
  NANDN U38111 ( .A(y[6223]), .B(x[6223]), .Z(n23371) );
  NAND U38112 ( .A(n18846), .B(n23371), .Z(n58823) );
  OR U38113 ( .A(n18847), .B(n58823), .Z(n18848) );
  AND U38114 ( .A(n23372), .B(n18848), .Z(n18849) );
  NANDN U38115 ( .A(x[6223]), .B(y[6223]), .Z(n51133) );
  AND U38116 ( .A(n18849), .B(n51133), .Z(n18851) );
  NANDN U38117 ( .A(y[6224]), .B(x[6224]), .Z(n18850) );
  NANDN U38118 ( .A(y[6225]), .B(x[6225]), .Z(n23368) );
  NAND U38119 ( .A(n18850), .B(n23368), .Z(n58824) );
  OR U38120 ( .A(n18851), .B(n58824), .Z(n18852) );
  AND U38121 ( .A(n58825), .B(n18852), .Z(n18853) );
  OR U38122 ( .A(n58826), .B(n18853), .Z(n18854) );
  NAND U38123 ( .A(n18855), .B(n18854), .Z(n18856) );
  NANDN U38124 ( .A(n58829), .B(n18856), .Z(n18857) );
  AND U38125 ( .A(n23366), .B(n18857), .Z(n18858) );
  NANDN U38126 ( .A(x[6229]), .B(y[6229]), .Z(n23367) );
  AND U38127 ( .A(n18858), .B(n23367), .Z(n18860) );
  NANDN U38128 ( .A(y[6230]), .B(x[6230]), .Z(n18859) );
  NANDN U38129 ( .A(y[6231]), .B(x[6231]), .Z(n45761) );
  AND U38130 ( .A(n18859), .B(n45761), .Z(n58832) );
  NANDN U38131 ( .A(n18860), .B(n58832), .Z(n18861) );
  NAND U38132 ( .A(n45762), .B(n18861), .Z(n18862) );
  NANDN U38133 ( .A(x[6231]), .B(y[6231]), .Z(n58834) );
  NANDN U38134 ( .A(n18862), .B(n58834), .Z(n18863) );
  NAND U38135 ( .A(n51130), .B(n18863), .Z(n18865) );
  ANDN U38136 ( .B(y[6233]), .A(x[6233]), .Z(n58835) );
  XNOR U38137 ( .A(x[6234]), .B(y[6234]), .Z(n23364) );
  NANDN U38138 ( .A(n58835), .B(n23364), .Z(n18864) );
  ANDN U38139 ( .B(n18865), .A(n18864), .Z(n18866) );
  OR U38140 ( .A(n58837), .B(n18866), .Z(n18867) );
  NAND U38141 ( .A(n18868), .B(n18867), .Z(n18869) );
  NANDN U38142 ( .A(n58840), .B(n18869), .Z(n18870) );
  AND U38143 ( .A(n23362), .B(n18870), .Z(n18871) );
  NANDN U38144 ( .A(n51128), .B(n18871), .Z(n18872) );
  NANDN U38145 ( .A(n58841), .B(n18872), .Z(n18873) );
  AND U38146 ( .A(n23360), .B(n18873), .Z(n18874) );
  NANDN U38147 ( .A(x[6239]), .B(y[6239]), .Z(n58842) );
  AND U38148 ( .A(n18874), .B(n58842), .Z(n18876) );
  NANDN U38149 ( .A(y[6240]), .B(x[6240]), .Z(n18875) );
  NANDN U38150 ( .A(y[6241]), .B(x[6241]), .Z(n23357) );
  AND U38151 ( .A(n18875), .B(n23357), .Z(n58845) );
  NANDN U38152 ( .A(n18876), .B(n58845), .Z(n18877) );
  NANDN U38153 ( .A(x[6241]), .B(y[6241]), .Z(n23358) );
  NANDN U38154 ( .A(x[6242]), .B(y[6242]), .Z(n23355) );
  AND U38155 ( .A(n23358), .B(n23355), .Z(n58846) );
  AND U38156 ( .A(n18877), .B(n58846), .Z(n18878) );
  NANDN U38157 ( .A(y[6242]), .B(x[6242]), .Z(n23356) );
  NANDN U38158 ( .A(y[6243]), .B(x[6243]), .Z(n23353) );
  NAND U38159 ( .A(n23356), .B(n23353), .Z(n51127) );
  OR U38160 ( .A(n18878), .B(n51127), .Z(n18879) );
  NAND U38161 ( .A(n51126), .B(n18879), .Z(n18880) );
  NANDN U38162 ( .A(n58847), .B(n18880), .Z(n18881) );
  AND U38163 ( .A(n23350), .B(n18881), .Z(n18882) );
  NANDN U38164 ( .A(x[6245]), .B(y[6245]), .Z(n58848) );
  AND U38165 ( .A(n18882), .B(n58848), .Z(n18884) );
  NANDN U38166 ( .A(y[6246]), .B(x[6246]), .Z(n18883) );
  NANDN U38167 ( .A(y[6247]), .B(x[6247]), .Z(n23347) );
  AND U38168 ( .A(n18883), .B(n23347), .Z(n58850) );
  NANDN U38169 ( .A(n18884), .B(n58850), .Z(n18885) );
  NAND U38170 ( .A(n18886), .B(n18885), .Z(n18887) );
  AND U38171 ( .A(n58851), .B(n18887), .Z(n18889) );
  XNOR U38172 ( .A(x[6250]), .B(y[6250]), .Z(n23346) );
  NANDN U38173 ( .A(x[6249]), .B(y[6249]), .Z(n58852) );
  AND U38174 ( .A(n23346), .B(n58852), .Z(n18888) );
  NANDN U38175 ( .A(n18889), .B(n18888), .Z(n18891) );
  NANDN U38176 ( .A(y[6250]), .B(x[6250]), .Z(n18890) );
  NANDN U38177 ( .A(y[6251]), .B(x[6251]), .Z(n23342) );
  AND U38178 ( .A(n18890), .B(n23342), .Z(n58854) );
  AND U38179 ( .A(n18891), .B(n58854), .Z(n18892) );
  NOR U38180 ( .A(n23344), .B(n18892), .Z(n18893) );
  NAND U38181 ( .A(n23343), .B(n18893), .Z(n18894) );
  NANDN U38182 ( .A(n58856), .B(n18894), .Z(n18895) );
  AND U38183 ( .A(n23341), .B(n18895), .Z(n18896) );
  NANDN U38184 ( .A(x[6253]), .B(y[6253]), .Z(n58858) );
  AND U38185 ( .A(n18896), .B(n58858), .Z(n18898) );
  NANDN U38186 ( .A(y[6254]), .B(x[6254]), .Z(n18897) );
  NANDN U38187 ( .A(y[6255]), .B(x[6255]), .Z(n45814) );
  NAND U38188 ( .A(n18897), .B(n45814), .Z(n58859) );
  OR U38189 ( .A(n18898), .B(n58859), .Z(n18899) );
  AND U38190 ( .A(n45815), .B(n18899), .Z(n18900) );
  NANDN U38191 ( .A(x[6255]), .B(y[6255]), .Z(n58860) );
  NANDN U38192 ( .A(y[6256]), .B(x[6256]), .Z(n18901) );
  NANDN U38193 ( .A(y[6257]), .B(x[6257]), .Z(n23338) );
  AND U38194 ( .A(n18901), .B(n23338), .Z(n58862) );
  NANDN U38195 ( .A(y[6258]), .B(x[6258]), .Z(n18902) );
  NANDN U38196 ( .A(y[6259]), .B(x[6259]), .Z(n23336) );
  AND U38197 ( .A(n18902), .B(n23336), .Z(n58865) );
  NANDN U38198 ( .A(x[6261]), .B(y[6261]), .Z(n58870) );
  NANDN U38199 ( .A(y[6262]), .B(x[6262]), .Z(n18903) );
  NANDN U38200 ( .A(y[6263]), .B(x[6263]), .Z(n23332) );
  NAND U38201 ( .A(n18903), .B(n23332), .Z(n58872) );
  NANDN U38202 ( .A(x[6263]), .B(y[6263]), .Z(n58873) );
  NANDN U38203 ( .A(y[6264]), .B(x[6264]), .Z(n18904) );
  NANDN U38204 ( .A(y[6265]), .B(x[6265]), .Z(n23330) );
  NAND U38205 ( .A(n18904), .B(n23330), .Z(n51118) );
  NANDN U38206 ( .A(x[6265]), .B(y[6265]), .Z(n23331) );
  NANDN U38207 ( .A(x[6266]), .B(y[6266]), .Z(n23328) );
  AND U38208 ( .A(n23331), .B(n23328), .Z(n51117) );
  NANDN U38209 ( .A(y[6266]), .B(x[6266]), .Z(n23329) );
  NANDN U38210 ( .A(y[6267]), .B(x[6267]), .Z(n45841) );
  NAND U38211 ( .A(n23329), .B(n45841), .Z(n58874) );
  NANDN U38212 ( .A(x[6267]), .B(y[6267]), .Z(n58875) );
  NANDN U38213 ( .A(n58877), .B(n18905), .Z(n18906) );
  AND U38214 ( .A(n23327), .B(n18906), .Z(n18907) );
  ANDN U38215 ( .B(y[6269]), .A(x[6269]), .Z(n58878) );
  ANDN U38216 ( .B(n18907), .A(n58878), .Z(n18909) );
  NANDN U38217 ( .A(y[6270]), .B(x[6270]), .Z(n18908) );
  NANDN U38218 ( .A(y[6271]), .B(x[6271]), .Z(n45851) );
  NAND U38219 ( .A(n18908), .B(n45851), .Z(n58880) );
  OR U38220 ( .A(n18909), .B(n58880), .Z(n18910) );
  AND U38221 ( .A(n45852), .B(n18910), .Z(n18911) );
  NANDN U38222 ( .A(x[6271]), .B(y[6271]), .Z(n58881) );
  AND U38223 ( .A(n18911), .B(n58881), .Z(n18913) );
  NANDN U38224 ( .A(y[6272]), .B(x[6272]), .Z(n18912) );
  NANDN U38225 ( .A(y[6273]), .B(x[6273]), .Z(n23324) );
  AND U38226 ( .A(n18912), .B(n23324), .Z(n58884) );
  NANDN U38227 ( .A(n18913), .B(n58884), .Z(n18914) );
  NAND U38228 ( .A(n18915), .B(n18914), .Z(n18916) );
  AND U38229 ( .A(n58885), .B(n18916), .Z(n18917) );
  ANDN U38230 ( .B(n58887), .A(n18917), .Z(n18918) );
  NAND U38231 ( .A(n45862), .B(n18918), .Z(n18919) );
  NANDN U38232 ( .A(n58888), .B(n18919), .Z(n18920) );
  AND U38233 ( .A(n23323), .B(n18920), .Z(n18921) );
  NANDN U38234 ( .A(n58889), .B(n18921), .Z(n18922) );
  NAND U38235 ( .A(n58891), .B(n18922), .Z(n18924) );
  XOR U38236 ( .A(x[6280]), .B(y[6280]), .Z(n18923) );
  ANDN U38237 ( .B(n18924), .A(n18923), .Z(n18925) );
  NANDN U38238 ( .A(x[6279]), .B(y[6279]), .Z(n58892) );
  AND U38239 ( .A(n18925), .B(n58892), .Z(n18927) );
  NANDN U38240 ( .A(y[6280]), .B(x[6280]), .Z(n18926) );
  NANDN U38241 ( .A(y[6281]), .B(x[6281]), .Z(n23319) );
  AND U38242 ( .A(n18926), .B(n23319), .Z(n58894) );
  NANDN U38243 ( .A(n18927), .B(n58894), .Z(n18928) );
  NAND U38244 ( .A(n18929), .B(n18928), .Z(n18930) );
  AND U38245 ( .A(n58896), .B(n18930), .Z(n18931) );
  ANDN U38246 ( .B(n58898), .A(n18931), .Z(n18932) );
  NAND U38247 ( .A(n45882), .B(n18932), .Z(n18933) );
  NANDN U38248 ( .A(n58899), .B(n18933), .Z(n18934) );
  AND U38249 ( .A(n23318), .B(n18934), .Z(n18935) );
  ANDN U38250 ( .B(y[6285]), .A(x[6285]), .Z(n58900) );
  ANDN U38251 ( .B(n18935), .A(n58900), .Z(n18937) );
  NANDN U38252 ( .A(y[6286]), .B(x[6286]), .Z(n18936) );
  NANDN U38253 ( .A(y[6287]), .B(x[6287]), .Z(n23315) );
  NAND U38254 ( .A(n18936), .B(n23315), .Z(n58902) );
  OR U38255 ( .A(n18937), .B(n58902), .Z(n18938) );
  AND U38256 ( .A(n23316), .B(n18938), .Z(n18939) );
  NANDN U38257 ( .A(x[6287]), .B(y[6287]), .Z(n58903) );
  AND U38258 ( .A(n18939), .B(n58903), .Z(n18941) );
  NANDN U38259 ( .A(y[6288]), .B(x[6288]), .Z(n18940) );
  NANDN U38260 ( .A(y[6289]), .B(x[6289]), .Z(n23312) );
  AND U38261 ( .A(n18940), .B(n23312), .Z(n58905) );
  NANDN U38262 ( .A(n18941), .B(n58905), .Z(n18942) );
  NAND U38263 ( .A(n18943), .B(n18942), .Z(n18944) );
  AND U38264 ( .A(n58906), .B(n18944), .Z(n18945) );
  ANDN U38265 ( .B(n58908), .A(n18945), .Z(n18946) );
  NAND U38266 ( .A(n23311), .B(n18946), .Z(n18947) );
  NANDN U38267 ( .A(n58909), .B(n18947), .Z(n18948) );
  AND U38268 ( .A(n23309), .B(n18948), .Z(n18949) );
  NANDN U38269 ( .A(x[6293]), .B(y[6293]), .Z(n58910) );
  AND U38270 ( .A(n18949), .B(n58910), .Z(n18951) );
  NANDN U38271 ( .A(y[6294]), .B(x[6294]), .Z(n18950) );
  NANDN U38272 ( .A(y[6295]), .B(x[6295]), .Z(n45907) );
  NAND U38273 ( .A(n18950), .B(n45907), .Z(n58912) );
  OR U38274 ( .A(n18951), .B(n58912), .Z(n18952) );
  AND U38275 ( .A(n45908), .B(n18952), .Z(n18953) );
  NANDN U38276 ( .A(x[6295]), .B(y[6295]), .Z(n58914) );
  AND U38277 ( .A(n18953), .B(n58914), .Z(n18955) );
  NANDN U38278 ( .A(y[6296]), .B(x[6296]), .Z(n18954) );
  NANDN U38279 ( .A(y[6297]), .B(x[6297]), .Z(n23306) );
  AND U38280 ( .A(n18954), .B(n23306), .Z(n58916) );
  NANDN U38281 ( .A(n18955), .B(n58916), .Z(n18956) );
  NAND U38282 ( .A(n18957), .B(n18956), .Z(n18958) );
  AND U38283 ( .A(n58917), .B(n18958), .Z(n18959) );
  ANDN U38284 ( .B(n58919), .A(n18959), .Z(n18960) );
  NAND U38285 ( .A(n23305), .B(n18960), .Z(n18961) );
  NANDN U38286 ( .A(n58920), .B(n18961), .Z(n18962) );
  AND U38287 ( .A(n23303), .B(n18962), .Z(n18963) );
  NANDN U38288 ( .A(x[6301]), .B(y[6301]), .Z(n58921) );
  AND U38289 ( .A(n18963), .B(n58921), .Z(n18965) );
  NANDN U38290 ( .A(y[6302]), .B(x[6302]), .Z(n18964) );
  NANDN U38291 ( .A(y[6303]), .B(x[6303]), .Z(n45925) );
  NAND U38292 ( .A(n18964), .B(n45925), .Z(n58923) );
  OR U38293 ( .A(n18965), .B(n58923), .Z(n18966) );
  AND U38294 ( .A(n45926), .B(n18966), .Z(n18967) );
  NANDN U38295 ( .A(x[6303]), .B(y[6303]), .Z(n58924) );
  AND U38296 ( .A(n18967), .B(n58924), .Z(n18969) );
  NANDN U38297 ( .A(y[6304]), .B(x[6304]), .Z(n18968) );
  NANDN U38298 ( .A(y[6305]), .B(x[6305]), .Z(n23300) );
  AND U38299 ( .A(n18968), .B(n23300), .Z(n58926) );
  NANDN U38300 ( .A(n18969), .B(n58926), .Z(n18970) );
  NAND U38301 ( .A(n18971), .B(n18970), .Z(n18972) );
  AND U38302 ( .A(n58929), .B(n18972), .Z(n18973) );
  ANDN U38303 ( .B(n51106), .A(n18973), .Z(n18974) );
  NAND U38304 ( .A(n45936), .B(n18974), .Z(n18975) );
  NANDN U38305 ( .A(n51104), .B(n18975), .Z(n18976) );
  AND U38306 ( .A(n23299), .B(n18976), .Z(n18977) );
  ANDN U38307 ( .B(y[6309]), .A(x[6309]), .Z(n58930) );
  ANDN U38308 ( .B(n18977), .A(n58930), .Z(n18979) );
  NANDN U38309 ( .A(y[6310]), .B(x[6310]), .Z(n18978) );
  NANDN U38310 ( .A(y[6311]), .B(x[6311]), .Z(n45946) );
  NAND U38311 ( .A(n18978), .B(n45946), .Z(n58932) );
  OR U38312 ( .A(n18979), .B(n58932), .Z(n18980) );
  AND U38313 ( .A(n45947), .B(n18980), .Z(n18981) );
  NANDN U38314 ( .A(n45943), .B(n18981), .Z(n18982) );
  NAND U38315 ( .A(n58935), .B(n18982), .Z(n18983) );
  NANDN U38316 ( .A(n51102), .B(n18983), .Z(n18984) );
  XNOR U38317 ( .A(x[6314]), .B(y[6314]), .Z(n23297) );
  NANDN U38318 ( .A(n18984), .B(n23297), .Z(n18985) );
  AND U38319 ( .A(n58936), .B(n18985), .Z(n18986) );
  ANDN U38320 ( .B(n58938), .A(n18986), .Z(n18987) );
  NAND U38321 ( .A(n45957), .B(n18987), .Z(n18988) );
  NANDN U38322 ( .A(n58939), .B(n18988), .Z(n18989) );
  AND U38323 ( .A(n23295), .B(n18989), .Z(n18990) );
  ANDN U38324 ( .B(y[6317]), .A(x[6317]), .Z(n58940) );
  ANDN U38325 ( .B(n18990), .A(n58940), .Z(n18992) );
  NANDN U38326 ( .A(y[6318]), .B(x[6318]), .Z(n18991) );
  NANDN U38327 ( .A(y[6319]), .B(x[6319]), .Z(n45966) );
  NAND U38328 ( .A(n18991), .B(n45966), .Z(n58943) );
  OR U38329 ( .A(n18992), .B(n58943), .Z(n18993) );
  AND U38330 ( .A(n45967), .B(n18993), .Z(n18994) );
  NANDN U38331 ( .A(x[6319]), .B(y[6319]), .Z(n58944) );
  AND U38332 ( .A(n18994), .B(n58944), .Z(n18996) );
  NANDN U38333 ( .A(y[6320]), .B(x[6320]), .Z(n18995) );
  NANDN U38334 ( .A(y[6321]), .B(x[6321]), .Z(n23292) );
  AND U38335 ( .A(n18995), .B(n23292), .Z(n58946) );
  NANDN U38336 ( .A(n18996), .B(n58946), .Z(n18997) );
  NAND U38337 ( .A(n18998), .B(n18997), .Z(n18999) );
  AND U38338 ( .A(n58947), .B(n18999), .Z(n19000) );
  ANDN U38339 ( .B(n58949), .A(n19000), .Z(n19001) );
  NAND U38340 ( .A(n45977), .B(n19001), .Z(n19002) );
  NANDN U38341 ( .A(n58950), .B(n19002), .Z(n19003) );
  AND U38342 ( .A(n23291), .B(n19003), .Z(n19004) );
  NANDN U38343 ( .A(n58951), .B(n19004), .Z(n19005) );
  NANDN U38344 ( .A(n58953), .B(n19005), .Z(n19006) );
  AND U38345 ( .A(n58954), .B(n19006), .Z(n19007) );
  OR U38346 ( .A(n58955), .B(n19007), .Z(n19008) );
  NAND U38347 ( .A(n58956), .B(n19008), .Z(n19009) );
  NANDN U38348 ( .A(n58958), .B(n19009), .Z(n19010) );
  AND U38349 ( .A(n58959), .B(n19010), .Z(n19011) );
  NANDN U38350 ( .A(y[6332]), .B(x[6332]), .Z(n23279) );
  NANDN U38351 ( .A(y[6333]), .B(x[6333]), .Z(n23278) );
  NAND U38352 ( .A(n23279), .B(n23278), .Z(n58960) );
  OR U38353 ( .A(n19011), .B(n58960), .Z(n19012) );
  AND U38354 ( .A(n58961), .B(n19012), .Z(n19013) );
  OR U38355 ( .A(n58962), .B(n19013), .Z(n19014) );
  NAND U38356 ( .A(n58963), .B(n19014), .Z(n19015) );
  NANDN U38357 ( .A(n58964), .B(n19015), .Z(n19016) );
  AND U38358 ( .A(n58965), .B(n19016), .Z(n19017) );
  NANDN U38359 ( .A(y[6338]), .B(x[6338]), .Z(n23271) );
  NANDN U38360 ( .A(y[6339]), .B(x[6339]), .Z(n23268) );
  NAND U38361 ( .A(n23271), .B(n23268), .Z(n58966) );
  OR U38362 ( .A(n19017), .B(n58966), .Z(n19018) );
  AND U38363 ( .A(n19019), .B(n19018), .Z(n19021) );
  NANDN U38364 ( .A(y[6340]), .B(x[6340]), .Z(n19020) );
  NANDN U38365 ( .A(y[6341]), .B(x[6341]), .Z(n23267) );
  NAND U38366 ( .A(n19020), .B(n23267), .Z(n58967) );
  OR U38367 ( .A(n19021), .B(n58967), .Z(n19022) );
  NAND U38368 ( .A(n58968), .B(n19022), .Z(n19023) );
  NANDN U38369 ( .A(n58969), .B(n19023), .Z(n19024) );
  NANDN U38370 ( .A(x[6343]), .B(y[6343]), .Z(n23264) );
  NANDN U38371 ( .A(x[6344]), .B(y[6344]), .Z(n46027) );
  AND U38372 ( .A(n23264), .B(n46027), .Z(n58970) );
  AND U38373 ( .A(n19024), .B(n58970), .Z(n19025) );
  NANDN U38374 ( .A(y[6344]), .B(x[6344]), .Z(n23262) );
  NANDN U38375 ( .A(y[6345]), .B(x[6345]), .Z(n23261) );
  NAND U38376 ( .A(n23262), .B(n23261), .Z(n51097) );
  OR U38377 ( .A(n19025), .B(n51097), .Z(n19026) );
  NAND U38378 ( .A(n58972), .B(n19026), .Z(n19027) );
  NANDN U38379 ( .A(n58973), .B(n19027), .Z(n19028) );
  AND U38380 ( .A(n46034), .B(n19028), .Z(n19029) );
  NANDN U38381 ( .A(x[6347]), .B(y[6347]), .Z(n58977) );
  NAND U38382 ( .A(n19029), .B(n58977), .Z(n19030) );
  NANDN U38383 ( .A(n58978), .B(n19030), .Z(n19031) );
  AND U38384 ( .A(n23258), .B(n19031), .Z(n19032) );
  ANDN U38385 ( .B(y[6349]), .A(x[6349]), .Z(n58979) );
  ANDN U38386 ( .B(n19032), .A(n58979), .Z(n19033) );
  OR U38387 ( .A(n58981), .B(n19033), .Z(n19034) );
  NAND U38388 ( .A(n19035), .B(n19034), .Z(n19036) );
  AND U38389 ( .A(n58982), .B(n19036), .Z(n19037) );
  NOR U38390 ( .A(n58984), .B(n19037), .Z(n19038) );
  NAND U38391 ( .A(n23256), .B(n19038), .Z(n19039) );
  NANDN U38392 ( .A(n58985), .B(n19039), .Z(n19040) );
  AND U38393 ( .A(n46055), .B(n19040), .Z(n19041) );
  NANDN U38394 ( .A(n46051), .B(n19041), .Z(n19042) );
  NAND U38395 ( .A(n58988), .B(n19042), .Z(n19043) );
  NAND U38396 ( .A(n23254), .B(n19043), .Z(n19044) );
  ANDN U38397 ( .B(y[6357]), .A(x[6357]), .Z(n58989) );
  OR U38398 ( .A(n19044), .B(n58989), .Z(n19045) );
  NAND U38399 ( .A(n58992), .B(n19045), .Z(n19047) );
  XNOR U38400 ( .A(x[6360]), .B(y[6360]), .Z(n46065) );
  NANDN U38401 ( .A(x[6359]), .B(y[6359]), .Z(n51094) );
  NAND U38402 ( .A(n46065), .B(n51094), .Z(n19046) );
  ANDN U38403 ( .B(n19047), .A(n19046), .Z(n19048) );
  OR U38404 ( .A(n58993), .B(n19048), .Z(n19049) );
  NAND U38405 ( .A(n58994), .B(n19049), .Z(n19050) );
  NANDN U38406 ( .A(n58995), .B(n19050), .Z(n19051) );
  AND U38407 ( .A(n23248), .B(n19051), .Z(n19052) );
  NANDN U38408 ( .A(x[6363]), .B(y[6363]), .Z(n58996) );
  AND U38409 ( .A(n19052), .B(n58996), .Z(n19054) );
  NANDN U38410 ( .A(y[6364]), .B(x[6364]), .Z(n19053) );
  NANDN U38411 ( .A(y[6365]), .B(x[6365]), .Z(n23245) );
  NAND U38412 ( .A(n19053), .B(n23245), .Z(n58998) );
  OR U38413 ( .A(n19054), .B(n58998), .Z(n19055) );
  AND U38414 ( .A(n23246), .B(n19055), .Z(n19056) );
  ANDN U38415 ( .B(y[6365]), .A(x[6365]), .Z(n51091) );
  ANDN U38416 ( .B(n19056), .A(n51091), .Z(n19058) );
  ANDN U38417 ( .B(x[6367]), .A(y[6367]), .Z(n46086) );
  NANDN U38418 ( .A(y[6366]), .B(x[6366]), .Z(n19057) );
  NANDN U38419 ( .A(n46086), .B(n19057), .Z(n58999) );
  OR U38420 ( .A(n19058), .B(n58999), .Z(n19059) );
  NAND U38421 ( .A(n59000), .B(n19059), .Z(n19060) );
  AND U38422 ( .A(n59001), .B(n19060), .Z(n19061) );
  NOR U38423 ( .A(n23243), .B(n19061), .Z(n19062) );
  NAND U38424 ( .A(n23242), .B(n19062), .Z(n19063) );
  NANDN U38425 ( .A(n59004), .B(n19063), .Z(n19064) );
  AND U38426 ( .A(n23240), .B(n19064), .Z(n19065) );
  NANDN U38427 ( .A(n46091), .B(n19065), .Z(n19066) );
  NAND U38428 ( .A(n59007), .B(n19066), .Z(n19067) );
  NANDN U38429 ( .A(n51088), .B(n19067), .Z(n19068) );
  NANDN U38430 ( .A(y[6374]), .B(x[6374]), .Z(n23236) );
  NANDN U38431 ( .A(y[6375]), .B(x[6375]), .Z(n23232) );
  AND U38432 ( .A(n23236), .B(n23232), .Z(n51087) );
  AND U38433 ( .A(n19068), .B(n51087), .Z(n19069) );
  NOR U38434 ( .A(n23234), .B(n19069), .Z(n19070) );
  NAND U38435 ( .A(n23233), .B(n19070), .Z(n19071) );
  NANDN U38436 ( .A(n59010), .B(n19071), .Z(n19072) );
  AND U38437 ( .A(n23230), .B(n19072), .Z(n19073) );
  NAND U38438 ( .A(n23231), .B(n19073), .Z(n19074) );
  NANDN U38439 ( .A(n59011), .B(n19074), .Z(n19075) );
  AND U38440 ( .A(n46111), .B(n19075), .Z(n19076) );
  NANDN U38441 ( .A(x[6379]), .B(y[6379]), .Z(n59012) );
  AND U38442 ( .A(n19076), .B(n59012), .Z(n19078) );
  NANDN U38443 ( .A(y[6380]), .B(x[6380]), .Z(n19077) );
  NANDN U38444 ( .A(y[6381]), .B(x[6381]), .Z(n23227) );
  AND U38445 ( .A(n19077), .B(n23227), .Z(n51084) );
  NANDN U38446 ( .A(n19078), .B(n51084), .Z(n19079) );
  NAND U38447 ( .A(n19080), .B(n19079), .Z(n19081) );
  NAND U38448 ( .A(n59018), .B(n19081), .Z(n19082) );
  AND U38449 ( .A(n46121), .B(n19082), .Z(n19083) );
  NAND U38450 ( .A(n59019), .B(n19083), .Z(n19084) );
  NANDN U38451 ( .A(n59021), .B(n19084), .Z(n19085) );
  AND U38452 ( .A(n23226), .B(n19085), .Z(n19086) );
  NANDN U38453 ( .A(n51082), .B(n19086), .Z(n19087) );
  NANDN U38454 ( .A(n59022), .B(n19087), .Z(n19088) );
  AND U38455 ( .A(n46131), .B(n19088), .Z(n19089) );
  NANDN U38456 ( .A(x[6387]), .B(y[6387]), .Z(n59023) );
  AND U38457 ( .A(n19089), .B(n59023), .Z(n19090) );
  OR U38458 ( .A(n59025), .B(n19090), .Z(n19091) );
  NAND U38459 ( .A(n19092), .B(n19091), .Z(n19094) );
  NANDN U38460 ( .A(y[6390]), .B(x[6390]), .Z(n19093) );
  NANDN U38461 ( .A(y[6391]), .B(x[6391]), .Z(n46141) );
  AND U38462 ( .A(n19093), .B(n46141), .Z(n59028) );
  AND U38463 ( .A(n19094), .B(n59028), .Z(n19095) );
  NOR U38464 ( .A(n46138), .B(n19095), .Z(n19096) );
  NAND U38465 ( .A(n46142), .B(n19096), .Z(n19097) );
  NANDN U38466 ( .A(n59033), .B(n19097), .Z(n19098) );
  AND U38467 ( .A(n23222), .B(n19098), .Z(n19099) );
  NANDN U38468 ( .A(n51080), .B(n19099), .Z(n19100) );
  NANDN U38469 ( .A(n59034), .B(n19100), .Z(n19101) );
  AND U38470 ( .A(n46152), .B(n19101), .Z(n19102) );
  NANDN U38471 ( .A(x[6395]), .B(y[6395]), .Z(n51078) );
  AND U38472 ( .A(n19102), .B(n51078), .Z(n19104) );
  NANDN U38473 ( .A(y[6396]), .B(x[6396]), .Z(n19103) );
  NANDN U38474 ( .A(y[6397]), .B(x[6397]), .Z(n23219) );
  NAND U38475 ( .A(n19103), .B(n23219), .Z(n51077) );
  OR U38476 ( .A(n19104), .B(n51077), .Z(n19105) );
  NAND U38477 ( .A(n19106), .B(n19105), .Z(n19108) );
  NANDN U38478 ( .A(y[6398]), .B(x[6398]), .Z(n19107) );
  NANDN U38479 ( .A(y[6399]), .B(x[6399]), .Z(n23217) );
  AND U38480 ( .A(n19107), .B(n23217), .Z(n59037) );
  AND U38481 ( .A(n19108), .B(n59037), .Z(n19109) );
  NOR U38482 ( .A(n46159), .B(n19109), .Z(n19110) );
  NAND U38483 ( .A(n23218), .B(n19110), .Z(n19111) );
  NANDN U38484 ( .A(n59040), .B(n19111), .Z(n19112) );
  AND U38485 ( .A(n23216), .B(n19112), .Z(n19113) );
  NANDN U38486 ( .A(x[6401]), .B(y[6401]), .Z(n51075) );
  NAND U38487 ( .A(n19113), .B(n51075), .Z(n19114) );
  NANDN U38488 ( .A(n59041), .B(n19114), .Z(n19115) );
  AND U38489 ( .A(n46171), .B(n19115), .Z(n19116) );
  NANDN U38490 ( .A(x[6403]), .B(y[6403]), .Z(n59044) );
  AND U38491 ( .A(n19116), .B(n59044), .Z(n19117) );
  OR U38492 ( .A(n59047), .B(n19117), .Z(n19118) );
  NAND U38493 ( .A(n19119), .B(n19118), .Z(n19120) );
  AND U38494 ( .A(n59049), .B(n19120), .Z(n19121) );
  ANDN U38495 ( .B(n59050), .A(n19121), .Z(n19122) );
  NAND U38496 ( .A(n46181), .B(n19122), .Z(n19123) );
  NANDN U38497 ( .A(n59052), .B(n19123), .Z(n19124) );
  AND U38498 ( .A(n23212), .B(n19124), .Z(n19125) );
  NANDN U38499 ( .A(n51072), .B(n19125), .Z(n19126) );
  NANDN U38500 ( .A(n59053), .B(n19126), .Z(n19127) );
  AND U38501 ( .A(n23210), .B(n19127), .Z(n19128) );
  NANDN U38502 ( .A(x[6411]), .B(y[6411]), .Z(n59055) );
  AND U38503 ( .A(n19128), .B(n59055), .Z(n19129) );
  OR U38504 ( .A(n59056), .B(n19129), .Z(n19130) );
  NAND U38505 ( .A(n19131), .B(n19130), .Z(n19133) );
  NANDN U38506 ( .A(y[6414]), .B(x[6414]), .Z(n19132) );
  NANDN U38507 ( .A(y[6415]), .B(x[6415]), .Z(n46199) );
  AND U38508 ( .A(n19132), .B(n46199), .Z(n59060) );
  AND U38509 ( .A(n19133), .B(n59060), .Z(n19134) );
  NOR U38510 ( .A(n46196), .B(n19134), .Z(n19135) );
  NAND U38511 ( .A(n46200), .B(n19135), .Z(n19136) );
  NANDN U38512 ( .A(n59064), .B(n19136), .Z(n19137) );
  AND U38513 ( .A(n23206), .B(n19137), .Z(n19138) );
  NANDN U38514 ( .A(n51070), .B(n19138), .Z(n19139) );
  NANDN U38515 ( .A(n59065), .B(n19139), .Z(n19140) );
  XOR U38516 ( .A(x[6420]), .B(y[6420]), .Z(n46212) );
  ANDN U38517 ( .B(n19140), .A(n46212), .Z(n19141) );
  NANDN U38518 ( .A(x[6419]), .B(y[6419]), .Z(n59066) );
  AND U38519 ( .A(n19141), .B(n59066), .Z(n19143) );
  NANDN U38520 ( .A(y[6420]), .B(x[6420]), .Z(n19142) );
  NANDN U38521 ( .A(y[6421]), .B(x[6421]), .Z(n23202) );
  AND U38522 ( .A(n19142), .B(n23202), .Z(n51069) );
  NANDN U38523 ( .A(n19143), .B(n51069), .Z(n19144) );
  NAND U38524 ( .A(n19145), .B(n19144), .Z(n19146) );
  NAND U38525 ( .A(n59070), .B(n19146), .Z(n19147) );
  AND U38526 ( .A(n23201), .B(n19147), .Z(n19148) );
  NAND U38527 ( .A(n59071), .B(n19148), .Z(n19149) );
  NANDN U38528 ( .A(n59074), .B(n19149), .Z(n19150) );
  AND U38529 ( .A(n23199), .B(n19150), .Z(n19151) );
  NANDN U38530 ( .A(x[6425]), .B(y[6425]), .Z(n51067) );
  NAND U38531 ( .A(n19151), .B(n51067), .Z(n19152) );
  NANDN U38532 ( .A(n59075), .B(n19152), .Z(n19153) );
  AND U38533 ( .A(n23197), .B(n19153), .Z(n19154) );
  NANDN U38534 ( .A(x[6427]), .B(y[6427]), .Z(n59077) );
  AND U38535 ( .A(n19154), .B(n59077), .Z(n19156) );
  NANDN U38536 ( .A(y[6428]), .B(x[6428]), .Z(n19155) );
  NANDN U38537 ( .A(y[6429]), .B(x[6429]), .Z(n23193) );
  NAND U38538 ( .A(n19155), .B(n23193), .Z(n59078) );
  OR U38539 ( .A(n19156), .B(n59078), .Z(n19157) );
  NAND U38540 ( .A(n59079), .B(n19157), .Z(n19159) );
  NANDN U38541 ( .A(y[6430]), .B(x[6430]), .Z(n19158) );
  NANDN U38542 ( .A(y[6431]), .B(x[6431]), .Z(n23191) );
  AND U38543 ( .A(n19158), .B(n23191), .Z(n59080) );
  AND U38544 ( .A(n19159), .B(n59080), .Z(n19161) );
  XNOR U38545 ( .A(x[6432]), .B(y[6432]), .Z(n23192) );
  ANDN U38546 ( .B(y[6431]), .A(x[6431]), .Z(n46233) );
  ANDN U38547 ( .B(n23192), .A(n46233), .Z(n19160) );
  NANDN U38548 ( .A(n19161), .B(n19160), .Z(n19163) );
  NANDN U38549 ( .A(y[6432]), .B(x[6432]), .Z(n19162) );
  NANDN U38550 ( .A(y[6433]), .B(x[6433]), .Z(n23189) );
  AND U38551 ( .A(n19162), .B(n23189), .Z(n59081) );
  AND U38552 ( .A(n19163), .B(n59081), .Z(n19164) );
  NANDN U38553 ( .A(x[6433]), .B(y[6433]), .Z(n23190) );
  NANDN U38554 ( .A(x[6434]), .B(y[6434]), .Z(n23187) );
  NAND U38555 ( .A(n23190), .B(n23187), .Z(n51064) );
  OR U38556 ( .A(n19164), .B(n51064), .Z(n19165) );
  NAND U38557 ( .A(n51063), .B(n19165), .Z(n19166) );
  NANDN U38558 ( .A(n59082), .B(n19166), .Z(n19167) );
  AND U38559 ( .A(n59085), .B(n19167), .Z(n19168) );
  NANDN U38560 ( .A(x[6437]), .B(y[6437]), .Z(n46247) );
  NANDN U38561 ( .A(x[6438]), .B(y[6438]), .Z(n23184) );
  NAND U38562 ( .A(n46247), .B(n23184), .Z(n51062) );
  OR U38563 ( .A(n19168), .B(n51062), .Z(n19169) );
  NAND U38564 ( .A(n59086), .B(n19169), .Z(n19170) );
  NAND U38565 ( .A(n23182), .B(n19170), .Z(n19171) );
  ANDN U38566 ( .B(y[6439]), .A(x[6439]), .Z(n23183) );
  OR U38567 ( .A(n19171), .B(n23183), .Z(n19172) );
  NAND U38568 ( .A(n59089), .B(n19172), .Z(n19174) );
  XNOR U38569 ( .A(x[6442]), .B(y[6442]), .Z(n23180) );
  NANDN U38570 ( .A(x[6441]), .B(y[6441]), .Z(n59090) );
  NAND U38571 ( .A(n23180), .B(n59090), .Z(n19173) );
  ANDN U38572 ( .B(n19174), .A(n19173), .Z(n19175) );
  OR U38573 ( .A(n59092), .B(n19175), .Z(n19176) );
  NAND U38574 ( .A(n59093), .B(n19176), .Z(n19177) );
  NANDN U38575 ( .A(n59094), .B(n19177), .Z(n19178) );
  AND U38576 ( .A(n59095), .B(n19178), .Z(n19179) );
  OR U38577 ( .A(n59096), .B(n19179), .Z(n19180) );
  NAND U38578 ( .A(n19181), .B(n19180), .Z(n19183) );
  NANDN U38579 ( .A(y[6448]), .B(x[6448]), .Z(n19182) );
  NANDN U38580 ( .A(y[6449]), .B(x[6449]), .Z(n23168) );
  AND U38581 ( .A(n19182), .B(n23168), .Z(n59099) );
  AND U38582 ( .A(n19183), .B(n59099), .Z(n19184) );
  NOR U38583 ( .A(n46276), .B(n19184), .Z(n19185) );
  NAND U38584 ( .A(n23169), .B(n19185), .Z(n19186) );
  NANDN U38585 ( .A(n59102), .B(n19186), .Z(n19187) );
  XOR U38586 ( .A(x[6452]), .B(y[6452]), .Z(n46284) );
  ANDN U38587 ( .B(n19187), .A(n46284), .Z(n19188) );
  NANDN U38588 ( .A(x[6451]), .B(y[6451]), .Z(n59103) );
  AND U38589 ( .A(n19188), .B(n59103), .Z(n19189) );
  ANDN U38590 ( .B(n59106), .A(n19189), .Z(n19190) );
  OR U38591 ( .A(n59107), .B(n19190), .Z(n19191) );
  NAND U38592 ( .A(n59108), .B(n19191), .Z(n19192) );
  NANDN U38593 ( .A(n59109), .B(n19192), .Z(n19193) );
  NAND U38594 ( .A(n59110), .B(n19193), .Z(n19194) );
  AND U38595 ( .A(n23160), .B(n19194), .Z(n19195) );
  NAND U38596 ( .A(n59112), .B(n19195), .Z(n19196) );
  NANDN U38597 ( .A(n59113), .B(n19196), .Z(n19197) );
  AND U38598 ( .A(n23158), .B(n19197), .Z(n19198) );
  NANDN U38599 ( .A(x[6459]), .B(y[6459]), .Z(n59114) );
  AND U38600 ( .A(n19198), .B(n59114), .Z(n19200) );
  NANDN U38601 ( .A(y[6460]), .B(x[6460]), .Z(n19199) );
  NANDN U38602 ( .A(y[6461]), .B(x[6461]), .Z(n23155) );
  NAND U38603 ( .A(n19199), .B(n23155), .Z(n59116) );
  OR U38604 ( .A(n19200), .B(n59116), .Z(n19201) );
  AND U38605 ( .A(n23156), .B(n19201), .Z(n19202) );
  NANDN U38606 ( .A(x[6461]), .B(y[6461]), .Z(n59117) );
  AND U38607 ( .A(n19202), .B(n59117), .Z(n19204) );
  NANDN U38608 ( .A(y[6462]), .B(x[6462]), .Z(n19203) );
  NANDN U38609 ( .A(y[6463]), .B(x[6463]), .Z(n23152) );
  AND U38610 ( .A(n19203), .B(n23152), .Z(n59119) );
  NANDN U38611 ( .A(n19204), .B(n59119), .Z(n19205) );
  NAND U38612 ( .A(n19206), .B(n19205), .Z(n19207) );
  AND U38613 ( .A(n59121), .B(n19207), .Z(n19208) );
  ANDN U38614 ( .B(n59123), .A(n19208), .Z(n19209) );
  NAND U38615 ( .A(n23151), .B(n19209), .Z(n19210) );
  NANDN U38616 ( .A(n59124), .B(n19210), .Z(n19211) );
  AND U38617 ( .A(n23149), .B(n19211), .Z(n19212) );
  NANDN U38618 ( .A(x[6467]), .B(y[6467]), .Z(n59125) );
  AND U38619 ( .A(n19212), .B(n59125), .Z(n19214) );
  NANDN U38620 ( .A(y[6468]), .B(x[6468]), .Z(n19213) );
  NANDN U38621 ( .A(y[6469]), .B(x[6469]), .Z(n23146) );
  NAND U38622 ( .A(n19213), .B(n23146), .Z(n59127) );
  OR U38623 ( .A(n19214), .B(n59127), .Z(n19215) );
  AND U38624 ( .A(n23147), .B(n19215), .Z(n19216) );
  NANDN U38625 ( .A(x[6469]), .B(y[6469]), .Z(n59128) );
  AND U38626 ( .A(n19216), .B(n59128), .Z(n19218) );
  NANDN U38627 ( .A(y[6470]), .B(x[6470]), .Z(n19217) );
  ANDN U38628 ( .B(x[6471]), .A(y[6471]), .Z(n46328) );
  ANDN U38629 ( .B(n19217), .A(n46328), .Z(n59130) );
  NANDN U38630 ( .A(n19218), .B(n59130), .Z(n19219) );
  NAND U38631 ( .A(n19220), .B(n19219), .Z(n19221) );
  AND U38632 ( .A(n59131), .B(n19221), .Z(n19222) );
  ANDN U38633 ( .B(n59133), .A(n19222), .Z(n19223) );
  NAND U38634 ( .A(n23145), .B(n19223), .Z(n19224) );
  NANDN U38635 ( .A(n59134), .B(n19224), .Z(n19225) );
  AND U38636 ( .A(n23143), .B(n19225), .Z(n19226) );
  NANDN U38637 ( .A(x[6475]), .B(y[6475]), .Z(n59136) );
  AND U38638 ( .A(n19226), .B(n59136), .Z(n19228) );
  NANDN U38639 ( .A(y[6476]), .B(x[6476]), .Z(n19227) );
  NANDN U38640 ( .A(y[6477]), .B(x[6477]), .Z(n23140) );
  NAND U38641 ( .A(n19227), .B(n23140), .Z(n59139) );
  OR U38642 ( .A(n19228), .B(n59139), .Z(n19229) );
  AND U38643 ( .A(n23141), .B(n19229), .Z(n19230) );
  NANDN U38644 ( .A(x[6477]), .B(y[6477]), .Z(n59142) );
  NAND U38645 ( .A(n19230), .B(n59142), .Z(n19231) );
  AND U38646 ( .A(n59145), .B(n19231), .Z(n19232) );
  OR U38647 ( .A(n19233), .B(n19232), .Z(n19234) );
  NAND U38648 ( .A(n59150), .B(n19234), .Z(n19235) );
  NANDN U38649 ( .A(n19236), .B(n19235), .Z(n19237) );
  NAND U38650 ( .A(n59156), .B(n19237), .Z(n19238) );
  AND U38651 ( .A(n23136), .B(n19238), .Z(n19239) );
  NANDN U38652 ( .A(x[6483]), .B(y[6483]), .Z(n59158) );
  AND U38653 ( .A(n19239), .B(n59158), .Z(n19240) );
  OR U38654 ( .A(n59161), .B(n19240), .Z(n19241) );
  NAND U38655 ( .A(n19242), .B(n19241), .Z(n19243) );
  NANDN U38656 ( .A(n59168), .B(n19243), .Z(n19244) );
  AND U38657 ( .A(n23132), .B(n19244), .Z(n19245) );
  NANDN U38658 ( .A(x[6487]), .B(y[6487]), .Z(n51052) );
  NAND U38659 ( .A(n19245), .B(n51052), .Z(n19246) );
  AND U38660 ( .A(n59172), .B(n19246), .Z(n19248) );
  XNOR U38661 ( .A(x[6490]), .B(y[6490]), .Z(n23130) );
  NANDN U38662 ( .A(x[6489]), .B(y[6489]), .Z(n59175) );
  AND U38663 ( .A(n23130), .B(n59175), .Z(n19247) );
  NANDN U38664 ( .A(n19248), .B(n19247), .Z(n19249) );
  NANDN U38665 ( .A(n59176), .B(n19249), .Z(n19250) );
  AND U38666 ( .A(n23128), .B(n19250), .Z(n19251) );
  NANDN U38667 ( .A(x[6491]), .B(y[6491]), .Z(n59177) );
  NAND U38668 ( .A(n19251), .B(n59177), .Z(n19253) );
  NANDN U38669 ( .A(y[6492]), .B(x[6492]), .Z(n19252) );
  NANDN U38670 ( .A(y[6493]), .B(x[6493]), .Z(n23125) );
  AND U38671 ( .A(n19252), .B(n23125), .Z(n59179) );
  AND U38672 ( .A(n19253), .B(n59179), .Z(n19254) );
  OR U38673 ( .A(n19255), .B(n19254), .Z(n19256) );
  XNOR U38674 ( .A(x[6498]), .B(y[6498]), .Z(n23122) );
  NANDN U38675 ( .A(x[6497]), .B(y[6497]), .Z(n59185) );
  NANDN U38676 ( .A(x[6501]), .B(y[6501]), .Z(n59191) );
  XNOR U38677 ( .A(y[6504]), .B(x[6504]), .Z(n46396) );
  NANDN U38678 ( .A(x[6503]), .B(y[6503]), .Z(n51048) );
  AND U38679 ( .A(n23114), .B(n19257), .Z(n19258) );
  NANDN U38680 ( .A(x[6507]), .B(y[6507]), .Z(n59198) );
  AND U38681 ( .A(n19258), .B(n59198), .Z(n19260) );
  NANDN U38682 ( .A(y[6508]), .B(x[6508]), .Z(n19259) );
  NANDN U38683 ( .A(y[6509]), .B(x[6509]), .Z(n23111) );
  AND U38684 ( .A(n19259), .B(n23111), .Z(n59200) );
  NANDN U38685 ( .A(n19260), .B(n59200), .Z(n19261) );
  NAND U38686 ( .A(n19262), .B(n19261), .Z(n19263) );
  NAND U38687 ( .A(n59203), .B(n19263), .Z(n19264) );
  AND U38688 ( .A(n23110), .B(n19264), .Z(n19265) );
  NANDN U38689 ( .A(x[6511]), .B(y[6511]), .Z(n51046) );
  AND U38690 ( .A(n19265), .B(n51046), .Z(n19267) );
  NANDN U38691 ( .A(y[6512]), .B(x[6512]), .Z(n19266) );
  NANDN U38692 ( .A(y[6513]), .B(x[6513]), .Z(n23107) );
  NAND U38693 ( .A(n19266), .B(n23107), .Z(n59206) );
  OR U38694 ( .A(n19267), .B(n59206), .Z(n19268) );
  AND U38695 ( .A(n19269), .B(n19268), .Z(n19271) );
  NANDN U38696 ( .A(y[6514]), .B(x[6514]), .Z(n19270) );
  NANDN U38697 ( .A(y[6515]), .B(x[6515]), .Z(n23105) );
  AND U38698 ( .A(n19270), .B(n23105), .Z(n51045) );
  NANDN U38699 ( .A(n19271), .B(n51045), .Z(n19272) );
  AND U38700 ( .A(n23106), .B(n19272), .Z(n19273) );
  NANDN U38701 ( .A(x[6515]), .B(y[6515]), .Z(n59210) );
  NAND U38702 ( .A(n19273), .B(n59210), .Z(n19274) );
  NAND U38703 ( .A(n59212), .B(n19274), .Z(n19275) );
  AND U38704 ( .A(n23104), .B(n19275), .Z(n19276) );
  NAND U38705 ( .A(n59213), .B(n19276), .Z(n19277) );
  NANDN U38706 ( .A(n59215), .B(n19277), .Z(n19278) );
  AND U38707 ( .A(n23102), .B(n19278), .Z(n19279) );
  NANDN U38708 ( .A(x[6519]), .B(y[6519]), .Z(n51043) );
  NAND U38709 ( .A(n19279), .B(n51043), .Z(n19280) );
  AND U38710 ( .A(n59216), .B(n19280), .Z(n19282) );
  XNOR U38711 ( .A(x[6522]), .B(y[6522]), .Z(n23100) );
  NANDN U38712 ( .A(x[6521]), .B(y[6521]), .Z(n59218) );
  AND U38713 ( .A(n23100), .B(n59218), .Z(n19281) );
  NANDN U38714 ( .A(n19282), .B(n19281), .Z(n19283) );
  NANDN U38715 ( .A(n59219), .B(n19283), .Z(n19284) );
  AND U38716 ( .A(n23098), .B(n19284), .Z(n19285) );
  NANDN U38717 ( .A(x[6523]), .B(y[6523]), .Z(n59221) );
  NAND U38718 ( .A(n19285), .B(n59221), .Z(n19286) );
  AND U38719 ( .A(n59223), .B(n19286), .Z(n19287) );
  OR U38720 ( .A(n19288), .B(n19287), .Z(n19289) );
  NAND U38721 ( .A(n59226), .B(n19289), .Z(n19290) );
  NANDN U38722 ( .A(n19291), .B(n19290), .Z(n19292) );
  NAND U38723 ( .A(n59227), .B(n19292), .Z(n19293) );
  AND U38724 ( .A(n59228), .B(n19293), .Z(n19294) );
  OR U38725 ( .A(n59229), .B(n19294), .Z(n19295) );
  NAND U38726 ( .A(n59230), .B(n19295), .Z(n19296) );
  NANDN U38727 ( .A(n59231), .B(n19296), .Z(n19297) );
  AND U38728 ( .A(n23086), .B(n19297), .Z(n19298) );
  NANDN U38729 ( .A(x[6533]), .B(y[6533]), .Z(n51039) );
  NAND U38730 ( .A(n19298), .B(n51039), .Z(n19299) );
  AND U38731 ( .A(n59232), .B(n19299), .Z(n19300) );
  OR U38732 ( .A(n19301), .B(n19300), .Z(n19302) );
  NAND U38733 ( .A(n51038), .B(n19302), .Z(n19303) );
  NANDN U38734 ( .A(n19304), .B(n19303), .Z(n19305) );
  NAND U38735 ( .A(n59238), .B(n19305), .Z(n19306) );
  AND U38736 ( .A(n23080), .B(n19306), .Z(n19307) );
  NANDN U38737 ( .A(x[6539]), .B(y[6539]), .Z(n59239) );
  AND U38738 ( .A(n19307), .B(n59239), .Z(n19308) );
  OR U38739 ( .A(n59241), .B(n19308), .Z(n19309) );
  NAND U38740 ( .A(n19310), .B(n19309), .Z(n19311) );
  NANDN U38741 ( .A(n59242), .B(n19311), .Z(n19312) );
  AND U38742 ( .A(n23076), .B(n19312), .Z(n19313) );
  NANDN U38743 ( .A(n59243), .B(n19313), .Z(n19315) );
  NANDN U38744 ( .A(y[6544]), .B(x[6544]), .Z(n19314) );
  NANDN U38745 ( .A(y[6545]), .B(x[6545]), .Z(n23073) );
  AND U38746 ( .A(n19314), .B(n23073), .Z(n51035) );
  AND U38747 ( .A(n19315), .B(n51035), .Z(n19316) );
  OR U38748 ( .A(n19317), .B(n19316), .Z(n19318) );
  NAND U38749 ( .A(n59246), .B(n19318), .Z(n19319) );
  NANDN U38750 ( .A(n59248), .B(n19319), .Z(n19320) );
  NAND U38751 ( .A(n59249), .B(n19320), .Z(n19321) );
  AND U38752 ( .A(n23070), .B(n19321), .Z(n19322) );
  NANDN U38753 ( .A(x[6549]), .B(y[6549]), .Z(n59251) );
  AND U38754 ( .A(n19322), .B(n59251), .Z(n19324) );
  NANDN U38755 ( .A(y[6550]), .B(x[6550]), .Z(n19323) );
  NANDN U38756 ( .A(y[6551]), .B(x[6551]), .Z(n23067) );
  NAND U38757 ( .A(n19323), .B(n23067), .Z(n59252) );
  OR U38758 ( .A(n19324), .B(n59252), .Z(n19325) );
  NAND U38759 ( .A(n19326), .B(n19325), .Z(n19327) );
  NAND U38760 ( .A(n59255), .B(n19327), .Z(n19328) );
  AND U38761 ( .A(n23066), .B(n19328), .Z(n19329) );
  NANDN U38762 ( .A(x[6553]), .B(y[6553]), .Z(n59256) );
  AND U38763 ( .A(n19329), .B(n59256), .Z(n19330) );
  OR U38764 ( .A(n59258), .B(n19330), .Z(n19331) );
  NAND U38765 ( .A(n19332), .B(n19331), .Z(n19333) );
  NANDN U38766 ( .A(n59259), .B(n19333), .Z(n19334) );
  AND U38767 ( .A(n23064), .B(n19334), .Z(n19335) );
  NANDN U38768 ( .A(x[6557]), .B(y[6557]), .Z(n59261) );
  AND U38769 ( .A(n19335), .B(n59261), .Z(n19336) );
  OR U38770 ( .A(n59262), .B(n19336), .Z(n19337) );
  NAND U38771 ( .A(n19338), .B(n19337), .Z(n19339) );
  NANDN U38772 ( .A(n59266), .B(n19339), .Z(n19340) );
  NAND U38773 ( .A(n59267), .B(n19340), .Z(n19341) );
  NAND U38774 ( .A(n59268), .B(n19341), .Z(n19342) );
  NAND U38775 ( .A(n59269), .B(n19342), .Z(n19343) );
  NANDN U38776 ( .A(y[6564]), .B(x[6564]), .Z(n23057) );
  NANDN U38777 ( .A(y[6565]), .B(x[6565]), .Z(n23053) );
  AND U38778 ( .A(n23057), .B(n23053), .Z(n51031) );
  AND U38779 ( .A(n19343), .B(n51031), .Z(n19344) );
  NOR U38780 ( .A(n23055), .B(n19344), .Z(n19345) );
  NAND U38781 ( .A(n23054), .B(n19345), .Z(n19346) );
  NANDN U38782 ( .A(n59272), .B(n19346), .Z(n19347) );
  AND U38783 ( .A(n23051), .B(n19347), .Z(n19348) );
  NANDN U38784 ( .A(n51029), .B(n19348), .Z(n19349) );
  AND U38785 ( .A(n59273), .B(n19349), .Z(n19351) );
  XNOR U38786 ( .A(x[6570]), .B(y[6570]), .Z(n23049) );
  NANDN U38787 ( .A(x[6569]), .B(y[6569]), .Z(n59275) );
  AND U38788 ( .A(n23049), .B(n59275), .Z(n19350) );
  NANDN U38789 ( .A(n19351), .B(n19350), .Z(n19352) );
  NANDN U38790 ( .A(n59276), .B(n19352), .Z(n19353) );
  AND U38791 ( .A(n23047), .B(n19353), .Z(n19354) );
  NANDN U38792 ( .A(x[6571]), .B(y[6571]), .Z(n59277) );
  NAND U38793 ( .A(n19354), .B(n59277), .Z(n19355) );
  NAND U38794 ( .A(n59280), .B(n19355), .Z(n19356) );
  AND U38795 ( .A(n46549), .B(n19356), .Z(n19357) );
  NANDN U38796 ( .A(x[6573]), .B(y[6573]), .Z(n59281) );
  AND U38797 ( .A(n19357), .B(n59281), .Z(n19359) );
  NANDN U38798 ( .A(y[6574]), .B(x[6574]), .Z(n19358) );
  ANDN U38799 ( .B(x[6575]), .A(y[6575]), .Z(n46556) );
  ANDN U38800 ( .B(n19358), .A(n46556), .Z(n59283) );
  NANDN U38801 ( .A(n19359), .B(n59283), .Z(n19360) );
  NAND U38802 ( .A(n19361), .B(n19360), .Z(n19362) );
  NAND U38803 ( .A(n59284), .B(n19362), .Z(n19363) );
  AND U38804 ( .A(n23045), .B(n19363), .Z(n19364) );
  NANDN U38805 ( .A(x[6577]), .B(y[6577]), .Z(n59286) );
  AND U38806 ( .A(n19364), .B(n59286), .Z(n19366) );
  NANDN U38807 ( .A(y[6578]), .B(x[6578]), .Z(n19365) );
  NANDN U38808 ( .A(y[6579]), .B(x[6579]), .Z(n23042) );
  NAND U38809 ( .A(n19365), .B(n23042), .Z(n59287) );
  OR U38810 ( .A(n19366), .B(n59287), .Z(n19367) );
  NAND U38811 ( .A(n19368), .B(n19367), .Z(n19369) );
  NAND U38812 ( .A(n59290), .B(n19369), .Z(n19370) );
  AND U38813 ( .A(n23041), .B(n19370), .Z(n19371) );
  NANDN U38814 ( .A(x[6581]), .B(y[6581]), .Z(n59291) );
  AND U38815 ( .A(n19371), .B(n59291), .Z(n19372) );
  OR U38816 ( .A(n59293), .B(n19372), .Z(n19373) );
  NAND U38817 ( .A(n19374), .B(n19373), .Z(n19375) );
  NANDN U38818 ( .A(n59296), .B(n19375), .Z(n19376) );
  AND U38819 ( .A(n23039), .B(n19376), .Z(n19377) );
  NANDN U38820 ( .A(x[6585]), .B(y[6585]), .Z(n59298) );
  NAND U38821 ( .A(n19377), .B(n59298), .Z(n19379) );
  NANDN U38822 ( .A(y[6586]), .B(x[6586]), .Z(n19378) );
  NANDN U38823 ( .A(y[6587]), .B(x[6587]), .Z(n23036) );
  AND U38824 ( .A(n19378), .B(n23036), .Z(n51024) );
  AND U38825 ( .A(n19379), .B(n51024), .Z(n19381) );
  XNOR U38826 ( .A(x[6588]), .B(y[6588]), .Z(n23037) );
  NANDN U38827 ( .A(x[6587]), .B(y[6587]), .Z(n59299) );
  AND U38828 ( .A(n23037), .B(n59299), .Z(n19380) );
  NANDN U38829 ( .A(n19381), .B(n19380), .Z(n19382) );
  NANDN U38830 ( .A(n59301), .B(n19382), .Z(n19383) );
  AND U38831 ( .A(n23035), .B(n19383), .Z(n19384) );
  NANDN U38832 ( .A(x[6589]), .B(y[6589]), .Z(n59302) );
  NAND U38833 ( .A(n19384), .B(n59302), .Z(n19386) );
  NANDN U38834 ( .A(y[6590]), .B(x[6590]), .Z(n19385) );
  NANDN U38835 ( .A(y[6591]), .B(x[6591]), .Z(n23032) );
  AND U38836 ( .A(n19385), .B(n23032), .Z(n59304) );
  AND U38837 ( .A(n19386), .B(n59304), .Z(n19387) );
  OR U38838 ( .A(n19388), .B(n19387), .Z(n19389) );
  NAND U38839 ( .A(n59305), .B(n19389), .Z(n19390) );
  NANDN U38840 ( .A(n19391), .B(n19390), .Z(n19392) );
  NAND U38841 ( .A(n59309), .B(n19392), .Z(n19393) );
  AND U38842 ( .A(n23029), .B(n19393), .Z(n19394) );
  NANDN U38843 ( .A(x[6595]), .B(y[6595]), .Z(n59310) );
  AND U38844 ( .A(n19394), .B(n59310), .Z(n19395) );
  OR U38845 ( .A(n59312), .B(n19395), .Z(n19396) );
  NAND U38846 ( .A(n19397), .B(n19396), .Z(n19398) );
  NANDN U38847 ( .A(n59315), .B(n19398), .Z(n19399) );
  AND U38848 ( .A(n23025), .B(n19399), .Z(n19400) );
  NANDN U38849 ( .A(x[6599]), .B(y[6599]), .Z(n51020) );
  NAND U38850 ( .A(n19400), .B(n51020), .Z(n19401) );
  AND U38851 ( .A(n59316), .B(n19401), .Z(n19403) );
  XNOR U38852 ( .A(x[6602]), .B(y[6602]), .Z(n23023) );
  NANDN U38853 ( .A(x[6601]), .B(y[6601]), .Z(n59318) );
  AND U38854 ( .A(n23023), .B(n59318), .Z(n19402) );
  NANDN U38855 ( .A(n19403), .B(n19402), .Z(n19404) );
  NANDN U38856 ( .A(n59319), .B(n19404), .Z(n19405) );
  AND U38857 ( .A(n23021), .B(n19405), .Z(n19406) );
  NANDN U38858 ( .A(x[6603]), .B(y[6603]), .Z(n59320) );
  NAND U38859 ( .A(n19406), .B(n59320), .Z(n19407) );
  NAND U38860 ( .A(n59322), .B(n19407), .Z(n19408) );
  AND U38861 ( .A(n23019), .B(n19408), .Z(n19409) );
  NANDN U38862 ( .A(x[6605]), .B(y[6605]), .Z(n59323) );
  AND U38863 ( .A(n19409), .B(n59323), .Z(n19411) );
  NANDN U38864 ( .A(y[6606]), .B(x[6606]), .Z(n19410) );
  ANDN U38865 ( .B(x[6607]), .A(y[6607]), .Z(n46625) );
  ANDN U38866 ( .B(n19410), .A(n46625), .Z(n59325) );
  NANDN U38867 ( .A(n19411), .B(n59325), .Z(n19412) );
  NAND U38868 ( .A(n19413), .B(n19412), .Z(n19414) );
  AND U38869 ( .A(n59329), .B(n19414), .Z(n19415) );
  OR U38870 ( .A(n19416), .B(n19415), .Z(n19417) );
  NAND U38871 ( .A(n59330), .B(n19417), .Z(n19418) );
  NANDN U38872 ( .A(n19419), .B(n19418), .Z(n19420) );
  NAND U38873 ( .A(n59333), .B(n19420), .Z(n19421) );
  AND U38874 ( .A(n23013), .B(n19421), .Z(n19422) );
  NANDN U38875 ( .A(n51016), .B(n19422), .Z(n19424) );
  NANDN U38876 ( .A(y[6614]), .B(x[6614]), .Z(n19423) );
  NANDN U38877 ( .A(y[6615]), .B(x[6615]), .Z(n46643) );
  AND U38878 ( .A(n19423), .B(n46643), .Z(n51015) );
  AND U38879 ( .A(n19424), .B(n51015), .Z(n19426) );
  XNOR U38880 ( .A(x[6616]), .B(y[6616]), .Z(n46644) );
  NANDN U38881 ( .A(x[6615]), .B(y[6615]), .Z(n59334) );
  AND U38882 ( .A(n46644), .B(n59334), .Z(n19425) );
  NANDN U38883 ( .A(n19426), .B(n19425), .Z(n19427) );
  NAND U38884 ( .A(n59336), .B(n19427), .Z(n19428) );
  AND U38885 ( .A(n23011), .B(n19428), .Z(n19429) );
  NANDN U38886 ( .A(n59337), .B(n19429), .Z(n19430) );
  NAND U38887 ( .A(n59340), .B(n19430), .Z(n19431) );
  NAND U38888 ( .A(n23008), .B(n19431), .Z(n19432) );
  ANDN U38889 ( .B(y[6619]), .A(x[6619]), .Z(n23009) );
  OR U38890 ( .A(n19432), .B(n23009), .Z(n19433) );
  NAND U38891 ( .A(n59343), .B(n19433), .Z(n19434) );
  NANDN U38892 ( .A(n51014), .B(n19434), .Z(n19435) );
  NAND U38893 ( .A(n59344), .B(n19435), .Z(n19436) );
  NAND U38894 ( .A(n59345), .B(n19436), .Z(n19437) );
  NANDN U38895 ( .A(y[6624]), .B(x[6624]), .Z(n23000) );
  NANDN U38896 ( .A(y[6625]), .B(x[6625]), .Z(n22996) );
  AND U38897 ( .A(n23000), .B(n22996), .Z(n59346) );
  AND U38898 ( .A(n19437), .B(n59346), .Z(n19438) );
  NOR U38899 ( .A(n22998), .B(n19438), .Z(n19439) );
  NAND U38900 ( .A(n22997), .B(n19439), .Z(n19440) );
  NAND U38901 ( .A(n59349), .B(n19440), .Z(n19441) );
  AND U38902 ( .A(n59350), .B(n19441), .Z(n19442) );
  NANDN U38903 ( .A(y[6628]), .B(x[6628]), .Z(n22994) );
  NANDN U38904 ( .A(y[6629]), .B(x[6629]), .Z(n22991) );
  NAND U38905 ( .A(n22994), .B(n22991), .Z(n59351) );
  OR U38906 ( .A(n19442), .B(n59351), .Z(n19443) );
  AND U38907 ( .A(n22992), .B(n19443), .Z(n19444) );
  NANDN U38908 ( .A(x[6629]), .B(y[6629]), .Z(n51012) );
  AND U38909 ( .A(n19444), .B(n51012), .Z(n19446) );
  NANDN U38910 ( .A(y[6630]), .B(x[6630]), .Z(n19445) );
  NANDN U38911 ( .A(y[6631]), .B(x[6631]), .Z(n22989) );
  AND U38912 ( .A(n19445), .B(n22989), .Z(n59352) );
  NANDN U38913 ( .A(n19446), .B(n59352), .Z(n19447) );
  NAND U38914 ( .A(n59353), .B(n19447), .Z(n19448) );
  NANDN U38915 ( .A(n59355), .B(n19448), .Z(n19449) );
  NAND U38916 ( .A(n59356), .B(n19449), .Z(n19450) );
  NAND U38917 ( .A(n59357), .B(n19450), .Z(n19451) );
  AND U38918 ( .A(n22983), .B(n19451), .Z(n19452) );
  NANDN U38919 ( .A(x[6635]), .B(y[6635]), .Z(n59358) );
  NAND U38920 ( .A(n19452), .B(n59358), .Z(n19453) );
  NAND U38921 ( .A(n59360), .B(n19453), .Z(n19454) );
  AND U38922 ( .A(n22981), .B(n19454), .Z(n19455) );
  NANDN U38923 ( .A(n59361), .B(n19455), .Z(n19456) );
  NAND U38924 ( .A(n59363), .B(n19456), .Z(n19457) );
  AND U38925 ( .A(n46696), .B(n19457), .Z(n19458) );
  NANDN U38926 ( .A(x[6639]), .B(y[6639]), .Z(n51010) );
  AND U38927 ( .A(n19458), .B(n51010), .Z(n19460) );
  NANDN U38928 ( .A(y[6640]), .B(x[6640]), .Z(n19459) );
  NANDN U38929 ( .A(y[6641]), .B(x[6641]), .Z(n22978) );
  AND U38930 ( .A(n19459), .B(n22978), .Z(n59364) );
  NANDN U38931 ( .A(n19460), .B(n59364), .Z(n19461) );
  NAND U38932 ( .A(n19462), .B(n19461), .Z(n19463) );
  NAND U38933 ( .A(n59367), .B(n19463), .Z(n19464) );
  AND U38934 ( .A(n46706), .B(n19464), .Z(n19465) );
  NANDN U38935 ( .A(x[6643]), .B(y[6643]), .Z(n51009) );
  AND U38936 ( .A(n19465), .B(n51009), .Z(n19467) );
  NANDN U38937 ( .A(y[6644]), .B(x[6644]), .Z(n19466) );
  NANDN U38938 ( .A(y[6645]), .B(x[6645]), .Z(n22976) );
  NAND U38939 ( .A(n19466), .B(n22976), .Z(n59369) );
  OR U38940 ( .A(n19467), .B(n59369), .Z(n19468) );
  NAND U38941 ( .A(n19469), .B(n19468), .Z(n19470) );
  NAND U38942 ( .A(n59372), .B(n19470), .Z(n19471) );
  AND U38943 ( .A(n46716), .B(n19471), .Z(n19472) );
  NANDN U38944 ( .A(x[6647]), .B(y[6647]), .Z(n51007) );
  AND U38945 ( .A(n19472), .B(n51007), .Z(n19474) );
  NANDN U38946 ( .A(y[6648]), .B(x[6648]), .Z(n19473) );
  NANDN U38947 ( .A(y[6649]), .B(x[6649]), .Z(n22973) );
  NAND U38948 ( .A(n19473), .B(n22973), .Z(n51005) );
  OR U38949 ( .A(n19474), .B(n51005), .Z(n19475) );
  NAND U38950 ( .A(n59373), .B(n19475), .Z(n19476) );
  NAND U38951 ( .A(n59374), .B(n19476), .Z(n19477) );
  NAND U38952 ( .A(n59375), .B(n19477), .Z(n19478) );
  NAND U38953 ( .A(n59376), .B(n19478), .Z(n19479) );
  AND U38954 ( .A(n59377), .B(n19479), .Z(n19480) );
  OR U38955 ( .A(n59378), .B(n19480), .Z(n19481) );
  NAND U38956 ( .A(n19482), .B(n19481), .Z(n19483) );
  NAND U38957 ( .A(n59381), .B(n19483), .Z(n19484) );
  AND U38958 ( .A(n22963), .B(n19484), .Z(n19485) );
  ANDN U38959 ( .B(y[6657]), .A(x[6657]), .Z(n59382) );
  ANDN U38960 ( .B(n19485), .A(n59382), .Z(n19487) );
  NANDN U38961 ( .A(y[6658]), .B(x[6658]), .Z(n19486) );
  NANDN U38962 ( .A(y[6659]), .B(x[6659]), .Z(n46743) );
  NAND U38963 ( .A(n19486), .B(n46743), .Z(n59384) );
  OR U38964 ( .A(n19487), .B(n59384), .Z(n19488) );
  NAND U38965 ( .A(n19489), .B(n19488), .Z(n19490) );
  NAND U38966 ( .A(n59387), .B(n19490), .Z(n19491) );
  AND U38967 ( .A(n22961), .B(n19491), .Z(n19492) );
  ANDN U38968 ( .B(y[6661]), .A(x[6661]), .Z(n59388) );
  ANDN U38969 ( .B(n19492), .A(n59388), .Z(n19494) );
  NANDN U38970 ( .A(y[6662]), .B(x[6662]), .Z(n19493) );
  NANDN U38971 ( .A(y[6663]), .B(x[6663]), .Z(n46754) );
  AND U38972 ( .A(n19493), .B(n46754), .Z(n59390) );
  NANDN U38973 ( .A(n19494), .B(n59390), .Z(n19495) );
  NAND U38974 ( .A(n19496), .B(n19495), .Z(n19497) );
  NAND U38975 ( .A(n50999), .B(n19497), .Z(n19498) );
  AND U38976 ( .A(n22959), .B(n19498), .Z(n19499) );
  NANDN U38977 ( .A(n59391), .B(n19499), .Z(n19501) );
  NANDN U38978 ( .A(y[6666]), .B(x[6666]), .Z(n19500) );
  NANDN U38979 ( .A(y[6667]), .B(x[6667]), .Z(n46764) );
  AND U38980 ( .A(n19500), .B(n46764), .Z(n59393) );
  AND U38981 ( .A(n19501), .B(n59393), .Z(n19503) );
  XNOR U38982 ( .A(x[6668]), .B(y[6668]), .Z(n46765) );
  NANDN U38983 ( .A(x[6667]), .B(y[6667]), .Z(n50998) );
  AND U38984 ( .A(n46765), .B(n50998), .Z(n19502) );
  NANDN U38985 ( .A(n19503), .B(n19502), .Z(n19504) );
  NANDN U38986 ( .A(n59394), .B(n19504), .Z(n19505) );
  AND U38987 ( .A(n22957), .B(n19505), .Z(n19506) );
  NANDN U38988 ( .A(n50995), .B(n19506), .Z(n19507) );
  NAND U38989 ( .A(n59396), .B(n19507), .Z(n19508) );
  AND U38990 ( .A(n59397), .B(n19508), .Z(n19509) );
  NANDN U38991 ( .A(y[6672]), .B(x[6672]), .Z(n22953) );
  NANDN U38992 ( .A(y[6673]), .B(x[6673]), .Z(n22950) );
  NAND U38993 ( .A(n22953), .B(n22950), .Z(n59398) );
  OR U38994 ( .A(n19509), .B(n59398), .Z(n19510) );
  NAND U38995 ( .A(n59399), .B(n19510), .Z(n19511) );
  NAND U38996 ( .A(n59400), .B(n19511), .Z(n19512) );
  AND U38997 ( .A(n22947), .B(n19512), .Z(n19513) );
  NANDN U38998 ( .A(x[6675]), .B(y[6675]), .Z(n59401) );
  AND U38999 ( .A(n19513), .B(n59401), .Z(n19515) );
  NANDN U39000 ( .A(y[6676]), .B(x[6676]), .Z(n19514) );
  NANDN U39001 ( .A(y[6677]), .B(x[6677]), .Z(n22944) );
  AND U39002 ( .A(n19514), .B(n22944), .Z(n59403) );
  NANDN U39003 ( .A(n19515), .B(n59403), .Z(n19516) );
  NAND U39004 ( .A(n19517), .B(n19516), .Z(n19518) );
  NAND U39005 ( .A(n59406), .B(n19518), .Z(n19519) );
  AND U39006 ( .A(n22943), .B(n19519), .Z(n19520) );
  NANDN U39007 ( .A(x[6679]), .B(y[6679]), .Z(n50993) );
  AND U39008 ( .A(n19520), .B(n50993), .Z(n19522) );
  NANDN U39009 ( .A(y[6680]), .B(x[6680]), .Z(n19521) );
  NANDN U39010 ( .A(y[6681]), .B(x[6681]), .Z(n22940) );
  AND U39011 ( .A(n19521), .B(n22940), .Z(n59407) );
  NANDN U39012 ( .A(n19522), .B(n59407), .Z(n19523) );
  NAND U39013 ( .A(n19524), .B(n19523), .Z(n19525) );
  NANDN U39014 ( .A(n59410), .B(n19525), .Z(n19526) );
  AND U39015 ( .A(n46799), .B(n19526), .Z(n19527) );
  NANDN U39016 ( .A(x[6683]), .B(y[6683]), .Z(n50992) );
  AND U39017 ( .A(n19527), .B(n50992), .Z(n19528) );
  OR U39018 ( .A(n59413), .B(n19528), .Z(n19529) );
  NAND U39019 ( .A(n19530), .B(n19529), .Z(n19531) );
  NANDN U39020 ( .A(n59416), .B(n19531), .Z(n19532) );
  AND U39021 ( .A(n22937), .B(n19532), .Z(n19533) );
  NANDN U39022 ( .A(x[6687]), .B(y[6687]), .Z(n50989) );
  NAND U39023 ( .A(n19533), .B(n50989), .Z(n19534) );
  NAND U39024 ( .A(n59417), .B(n19534), .Z(n19535) );
  AND U39025 ( .A(n22935), .B(n19535), .Z(n19536) );
  NANDN U39026 ( .A(x[6689]), .B(y[6689]), .Z(n50987) );
  AND U39027 ( .A(n19536), .B(n50987), .Z(n19538) );
  NANDN U39028 ( .A(y[6690]), .B(x[6690]), .Z(n19537) );
  NANDN U39029 ( .A(y[6691]), .B(x[6691]), .Z(n46816) );
  AND U39030 ( .A(n19537), .B(n46816), .Z(n59418) );
  NANDN U39031 ( .A(n19538), .B(n59418), .Z(n19539) );
  NAND U39032 ( .A(n19540), .B(n19539), .Z(n19541) );
  NAND U39033 ( .A(n59421), .B(n19541), .Z(n19542) );
  AND U39034 ( .A(n22933), .B(n19542), .Z(n19543) );
  ANDN U39035 ( .B(y[6693]), .A(x[6693]), .Z(n50985) );
  ANDN U39036 ( .B(n19543), .A(n50985), .Z(n19545) );
  NANDN U39037 ( .A(y[6694]), .B(x[6694]), .Z(n19544) );
  NANDN U39038 ( .A(y[6695]), .B(x[6695]), .Z(n46826) );
  AND U39039 ( .A(n19544), .B(n46826), .Z(n59422) );
  NANDN U39040 ( .A(n19545), .B(n59422), .Z(n19546) );
  AND U39041 ( .A(n19547), .B(n19546), .Z(n19549) );
  NANDN U39042 ( .A(y[6696]), .B(x[6696]), .Z(n19548) );
  NANDN U39043 ( .A(y[6697]), .B(x[6697]), .Z(n22930) );
  NAND U39044 ( .A(n19548), .B(n22930), .Z(n59426) );
  OR U39045 ( .A(n19549), .B(n59426), .Z(n19550) );
  NAND U39046 ( .A(n19551), .B(n19550), .Z(n19553) );
  NANDN U39047 ( .A(y[6698]), .B(x[6698]), .Z(n19552) );
  NANDN U39048 ( .A(y[6699]), .B(x[6699]), .Z(n46836) );
  AND U39049 ( .A(n19552), .B(n46836), .Z(n50984) );
  AND U39050 ( .A(n19553), .B(n50984), .Z(n19555) );
  XNOR U39051 ( .A(x[6700]), .B(y[6700]), .Z(n46837) );
  NANDN U39052 ( .A(x[6699]), .B(y[6699]), .Z(n59429) );
  AND U39053 ( .A(n46837), .B(n59429), .Z(n19554) );
  NANDN U39054 ( .A(n19555), .B(n19554), .Z(n19556) );
  NAND U39055 ( .A(n59431), .B(n19556), .Z(n19557) );
  AND U39056 ( .A(n22929), .B(n19557), .Z(n19558) );
  NANDN U39057 ( .A(n59432), .B(n19558), .Z(n19559) );
  NAND U39058 ( .A(n59434), .B(n19559), .Z(n19560) );
  AND U39059 ( .A(n46847), .B(n19560), .Z(n19561) );
  NANDN U39060 ( .A(x[6703]), .B(y[6703]), .Z(n59435) );
  AND U39061 ( .A(n19561), .B(n59435), .Z(n19563) );
  NANDN U39062 ( .A(y[6704]), .B(x[6704]), .Z(n19562) );
  NANDN U39063 ( .A(y[6705]), .B(x[6705]), .Z(n22926) );
  AND U39064 ( .A(n19562), .B(n22926), .Z(n59437) );
  NANDN U39065 ( .A(n19563), .B(n59437), .Z(n19564) );
  NAND U39066 ( .A(n19565), .B(n19564), .Z(n19566) );
  NAND U39067 ( .A(n59440), .B(n19566), .Z(n19567) );
  AND U39068 ( .A(n46857), .B(n19567), .Z(n19568) );
  NANDN U39069 ( .A(x[6707]), .B(y[6707]), .Z(n50982) );
  AND U39070 ( .A(n19568), .B(n50982), .Z(n19570) );
  NANDN U39071 ( .A(y[6708]), .B(x[6708]), .Z(n19569) );
  NANDN U39072 ( .A(y[6709]), .B(x[6709]), .Z(n22924) );
  AND U39073 ( .A(n19569), .B(n22924), .Z(n59442) );
  NANDN U39074 ( .A(n19570), .B(n59442), .Z(n19571) );
  NAND U39075 ( .A(n19572), .B(n19571), .Z(n19573) );
  NAND U39076 ( .A(n59445), .B(n19573), .Z(n19574) );
  AND U39077 ( .A(n46867), .B(n19574), .Z(n19575) );
  NANDN U39078 ( .A(x[6711]), .B(y[6711]), .Z(n50981) );
  AND U39079 ( .A(n19575), .B(n50981), .Z(n19576) );
  OR U39080 ( .A(n59446), .B(n19576), .Z(n19577) );
  NAND U39081 ( .A(n19578), .B(n19577), .Z(n19579) );
  NANDN U39082 ( .A(n59449), .B(n19579), .Z(n19580) );
  AND U39083 ( .A(n22921), .B(n19580), .Z(n19581) );
  NANDN U39084 ( .A(x[6715]), .B(y[6715]), .Z(n50978) );
  NAND U39085 ( .A(n19581), .B(n50978), .Z(n19582) );
  AND U39086 ( .A(n59450), .B(n19582), .Z(n19583) );
  OR U39087 ( .A(n59451), .B(n19583), .Z(n19584) );
  NAND U39088 ( .A(n59453), .B(n19584), .Z(n19585) );
  NANDN U39089 ( .A(n22915), .B(n19585), .Z(n19586) );
  XNOR U39090 ( .A(x[6720]), .B(y[6720]), .Z(n46885) );
  NANDN U39091 ( .A(n19586), .B(n46885), .Z(n19587) );
  NAND U39092 ( .A(n59456), .B(n19587), .Z(n19588) );
  AND U39093 ( .A(n22914), .B(n19588), .Z(n19589) );
  ANDN U39094 ( .B(y[6721]), .A(x[6721]), .Z(n50976) );
  ANDN U39095 ( .B(n19589), .A(n50976), .Z(n19591) );
  NANDN U39096 ( .A(y[6722]), .B(x[6722]), .Z(n19590) );
  NANDN U39097 ( .A(y[6723]), .B(x[6723]), .Z(n22911) );
  NAND U39098 ( .A(n19590), .B(n22911), .Z(n59457) );
  OR U39099 ( .A(n19591), .B(n59457), .Z(n19592) );
  NAND U39100 ( .A(n19593), .B(n19592), .Z(n19594) );
  NAND U39101 ( .A(n59460), .B(n19594), .Z(n19595) );
  AND U39102 ( .A(n22910), .B(n19595), .Z(n19596) );
  NANDN U39103 ( .A(x[6725]), .B(y[6725]), .Z(n59461) );
  AND U39104 ( .A(n19596), .B(n59461), .Z(n19597) );
  OR U39105 ( .A(n59463), .B(n19597), .Z(n19598) );
  NAND U39106 ( .A(n19599), .B(n19598), .Z(n19600) );
  NAND U39107 ( .A(n59466), .B(n19600), .Z(n19601) );
  AND U39108 ( .A(n22908), .B(n19601), .Z(n19602) );
  NANDN U39109 ( .A(n59467), .B(n19602), .Z(n19603) );
  AND U39110 ( .A(n59469), .B(n19603), .Z(n19605) );
  XNOR U39111 ( .A(x[6732]), .B(y[6732]), .Z(n46913) );
  NANDN U39112 ( .A(x[6731]), .B(y[6731]), .Z(n50973) );
  AND U39113 ( .A(n46913), .B(n50973), .Z(n19604) );
  NANDN U39114 ( .A(n19605), .B(n19604), .Z(n19606) );
  NANDN U39115 ( .A(n50972), .B(n19606), .Z(n19607) );
  AND U39116 ( .A(n22906), .B(n19607), .Z(n19608) );
  NANDN U39117 ( .A(n59471), .B(n19608), .Z(n19609) );
  NAND U39118 ( .A(n59473), .B(n19609), .Z(n19610) );
  AND U39119 ( .A(n59474), .B(n19610), .Z(n19611) );
  OR U39120 ( .A(n59475), .B(n19611), .Z(n19612) );
  NAND U39121 ( .A(n19613), .B(n19612), .Z(n19614) );
  NAND U39122 ( .A(n59478), .B(n19614), .Z(n19615) );
  AND U39123 ( .A(n46932), .B(n19615), .Z(n19616) );
  NANDN U39124 ( .A(x[6739]), .B(y[6739]), .Z(n59479) );
  AND U39125 ( .A(n19616), .B(n59479), .Z(n19618) );
  NANDN U39126 ( .A(y[6740]), .B(x[6740]), .Z(n19617) );
  NANDN U39127 ( .A(y[6741]), .B(x[6741]), .Z(n22897) );
  NAND U39128 ( .A(n19617), .B(n22897), .Z(n59481) );
  OR U39129 ( .A(n19618), .B(n59481), .Z(n19619) );
  NAND U39130 ( .A(n19620), .B(n19619), .Z(n19621) );
  NAND U39131 ( .A(n59482), .B(n19621), .Z(n19622) );
  AND U39132 ( .A(n46942), .B(n19622), .Z(n19623) );
  NANDN U39133 ( .A(x[6743]), .B(y[6743]), .Z(n59483) );
  AND U39134 ( .A(n19623), .B(n59483), .Z(n19625) );
  NANDN U39135 ( .A(y[6744]), .B(x[6744]), .Z(n19624) );
  NANDN U39136 ( .A(y[6745]), .B(x[6745]), .Z(n22895) );
  NAND U39137 ( .A(n19624), .B(n22895), .Z(n59486) );
  OR U39138 ( .A(n19625), .B(n59486), .Z(n19626) );
  NAND U39139 ( .A(n19627), .B(n19626), .Z(n19628) );
  NANDN U39140 ( .A(n59489), .B(n19628), .Z(n19629) );
  AND U39141 ( .A(n46952), .B(n19629), .Z(n19630) );
  NANDN U39142 ( .A(x[6747]), .B(y[6747]), .Z(n59490) );
  AND U39143 ( .A(n19630), .B(n59490), .Z(n19632) );
  NANDN U39144 ( .A(y[6748]), .B(x[6748]), .Z(n19631) );
  NANDN U39145 ( .A(y[6749]), .B(x[6749]), .Z(n22893) );
  AND U39146 ( .A(n19631), .B(n22893), .Z(n59492) );
  NANDN U39147 ( .A(n19632), .B(n59492), .Z(n19633) );
  AND U39148 ( .A(n22894), .B(n19633), .Z(n19634) );
  NANDN U39149 ( .A(n59493), .B(n19634), .Z(n19635) );
  NAND U39150 ( .A(n59495), .B(n19635), .Z(n19636) );
  NAND U39151 ( .A(n59496), .B(n19636), .Z(n19637) );
  NAND U39152 ( .A(n59497), .B(n19637), .Z(n19638) );
  AND U39153 ( .A(n22888), .B(n19638), .Z(n19639) );
  NANDN U39154 ( .A(x[6753]), .B(y[6753]), .Z(n59498) );
  AND U39155 ( .A(n19639), .B(n59498), .Z(n19641) );
  NANDN U39156 ( .A(y[6754]), .B(x[6754]), .Z(n19640) );
  NANDN U39157 ( .A(y[6755]), .B(x[6755]), .Z(n46969) );
  AND U39158 ( .A(n19640), .B(n46969), .Z(n59500) );
  NANDN U39159 ( .A(n19641), .B(n59500), .Z(n19642) );
  AND U39160 ( .A(n46970), .B(n19642), .Z(n19643) );
  NAND U39161 ( .A(n50969), .B(n19643), .Z(n19644) );
  NANDN U39162 ( .A(n59503), .B(n19644), .Z(n19645) );
  AND U39163 ( .A(n22886), .B(n19645), .Z(n19646) );
  NANDN U39164 ( .A(n59504), .B(n19646), .Z(n19647) );
  AND U39165 ( .A(n59506), .B(n19647), .Z(n19649) );
  XNOR U39166 ( .A(x[6760]), .B(y[6760]), .Z(n46980) );
  NANDN U39167 ( .A(x[6759]), .B(y[6759]), .Z(n59507) );
  AND U39168 ( .A(n46980), .B(n59507), .Z(n19648) );
  NANDN U39169 ( .A(n19649), .B(n19648), .Z(n19650) );
  NANDN U39170 ( .A(n59508), .B(n19650), .Z(n19651) );
  AND U39171 ( .A(n22884), .B(n19651), .Z(n19652) );
  NANDN U39172 ( .A(n59509), .B(n19652), .Z(n19653) );
  AND U39173 ( .A(n59511), .B(n19653), .Z(n19654) );
  OR U39174 ( .A(n19655), .B(n19654), .Z(n19656) );
  NAND U39175 ( .A(n59514), .B(n19656), .Z(n19657) );
  NANDN U39176 ( .A(n19658), .B(n19657), .Z(n19659) );
  NAND U39177 ( .A(n59516), .B(n19659), .Z(n19660) );
  AND U39178 ( .A(n47000), .B(n19660), .Z(n19661) );
  NANDN U39179 ( .A(x[6767]), .B(y[6767]), .Z(n59517) );
  AND U39180 ( .A(n19661), .B(n59517), .Z(n19662) );
  OR U39181 ( .A(n59519), .B(n19662), .Z(n19663) );
  NAND U39182 ( .A(n19664), .B(n19663), .Z(n19665) );
  NANDN U39183 ( .A(n59520), .B(n19665), .Z(n19666) );
  AND U39184 ( .A(n22877), .B(n19666), .Z(n19667) );
  NANDN U39185 ( .A(x[6771]), .B(y[6771]), .Z(n59521) );
  NAND U39186 ( .A(n19667), .B(n59521), .Z(n19668) );
  AND U39187 ( .A(n59523), .B(n19668), .Z(n19670) );
  XNOR U39188 ( .A(x[6774]), .B(y[6774]), .Z(n22875) );
  NANDN U39189 ( .A(x[6773]), .B(y[6773]), .Z(n59524) );
  AND U39190 ( .A(n22875), .B(n59524), .Z(n19669) );
  NANDN U39191 ( .A(n19670), .B(n19669), .Z(n19671) );
  NANDN U39192 ( .A(n59526), .B(n19671), .Z(n19672) );
  AND U39193 ( .A(n47018), .B(n19672), .Z(n19673) );
  NANDN U39194 ( .A(x[6775]), .B(y[6775]), .Z(n59527) );
  NAND U39195 ( .A(n19673), .B(n59527), .Z(n19674) );
  NAND U39196 ( .A(n59529), .B(n19674), .Z(n19675) );
  AND U39197 ( .A(n22873), .B(n19675), .Z(n19676) );
  ANDN U39198 ( .B(y[6777]), .A(x[6777]), .Z(n59530) );
  ANDN U39199 ( .B(n19676), .A(n59530), .Z(n19678) );
  NANDN U39200 ( .A(y[6778]), .B(x[6778]), .Z(n19677) );
  NANDN U39201 ( .A(y[6779]), .B(x[6779]), .Z(n47027) );
  AND U39202 ( .A(n19677), .B(n47027), .Z(n59532) );
  NANDN U39203 ( .A(n19678), .B(n59532), .Z(n19679) );
  NAND U39204 ( .A(n19680), .B(n19679), .Z(n19681) );
  NAND U39205 ( .A(n59535), .B(n19681), .Z(n19682) );
  AND U39206 ( .A(n22871), .B(n19682), .Z(n19683) );
  ANDN U39207 ( .B(y[6781]), .A(x[6781]), .Z(n59536) );
  ANDN U39208 ( .B(n19683), .A(n59536), .Z(n19685) );
  NANDN U39209 ( .A(y[6782]), .B(x[6782]), .Z(n19684) );
  NANDN U39210 ( .A(y[6783]), .B(x[6783]), .Z(n47037) );
  NAND U39211 ( .A(n19684), .B(n47037), .Z(n59538) );
  OR U39212 ( .A(n19685), .B(n59538), .Z(n19686) );
  NAND U39213 ( .A(n19687), .B(n19686), .Z(n19688) );
  NAND U39214 ( .A(n59539), .B(n19688), .Z(n19689) );
  AND U39215 ( .A(n22869), .B(n19689), .Z(n19690) );
  ANDN U39216 ( .B(y[6785]), .A(x[6785]), .Z(n59540) );
  ANDN U39217 ( .B(n19690), .A(n59540), .Z(n19692) );
  NANDN U39218 ( .A(y[6786]), .B(x[6786]), .Z(n19691) );
  NANDN U39219 ( .A(y[6787]), .B(x[6787]), .Z(n47047) );
  AND U39220 ( .A(n19691), .B(n47047), .Z(n59542) );
  NANDN U39221 ( .A(n19692), .B(n59542), .Z(n19693) );
  NAND U39222 ( .A(n19694), .B(n19693), .Z(n19695) );
  NANDN U39223 ( .A(n59544), .B(n19695), .Z(n19696) );
  AND U39224 ( .A(n22867), .B(n19696), .Z(n19697) );
  NANDN U39225 ( .A(n59545), .B(n19697), .Z(n19698) );
  AND U39226 ( .A(n59547), .B(n19698), .Z(n19700) );
  XNOR U39227 ( .A(x[6792]), .B(y[6792]), .Z(n22865) );
  NANDN U39228 ( .A(x[6791]), .B(y[6791]), .Z(n59548) );
  AND U39229 ( .A(n22865), .B(n59548), .Z(n19699) );
  NANDN U39230 ( .A(n19700), .B(n19699), .Z(n19701) );
  NANDN U39231 ( .A(n59552), .B(n19701), .Z(n19702) );
  AND U39232 ( .A(n22863), .B(n19702), .Z(n19703) );
  NANDN U39233 ( .A(x[6793]), .B(y[6793]), .Z(n50957) );
  NAND U39234 ( .A(n19703), .B(n50957), .Z(n19704) );
  AND U39235 ( .A(n59553), .B(n19704), .Z(n19705) );
  OR U39236 ( .A(n19706), .B(n19705), .Z(n19707) );
  NAND U39237 ( .A(n59556), .B(n19707), .Z(n19708) );
  NANDN U39238 ( .A(n19709), .B(n19708), .Z(n19710) );
  NAND U39239 ( .A(n59557), .B(n19710), .Z(n19711) );
  AND U39240 ( .A(n47076), .B(n19711), .Z(n19712) );
  NANDN U39241 ( .A(x[6799]), .B(y[6799]), .Z(n59558) );
  NAND U39242 ( .A(n19712), .B(n59558), .Z(n19713) );
  AND U39243 ( .A(n59560), .B(n19713), .Z(n19714) );
  NOR U39244 ( .A(n59561), .B(n19714), .Z(n19715) );
  NAND U39245 ( .A(n22859), .B(n19715), .Z(n19716) );
  NANDN U39246 ( .A(n59564), .B(n19716), .Z(n19717) );
  AND U39247 ( .A(n47086), .B(n19717), .Z(n19718) );
  NANDN U39248 ( .A(x[6803]), .B(y[6803]), .Z(n59565) );
  AND U39249 ( .A(n19718), .B(n59565), .Z(n19720) );
  NANDN U39250 ( .A(y[6805]), .B(x[6805]), .Z(n47092) );
  NANDN U39251 ( .A(y[6804]), .B(x[6804]), .Z(n19719) );
  AND U39252 ( .A(n47092), .B(n19719), .Z(n59567) );
  NANDN U39253 ( .A(n19720), .B(n59567), .Z(n19721) );
  AND U39254 ( .A(n59568), .B(n19721), .Z(n19724) );
  NANDN U39255 ( .A(y[6806]), .B(x[6806]), .Z(n19723) );
  NANDN U39256 ( .A(y[6807]), .B(x[6807]), .Z(n19722) );
  AND U39257 ( .A(n19723), .B(n19722), .Z(n59569) );
  NANDN U39258 ( .A(n19724), .B(n59569), .Z(n19725) );
  NAND U39259 ( .A(n59570), .B(n19725), .Z(n19726) );
  NANDN U39260 ( .A(n50953), .B(n19726), .Z(n19727) );
  AND U39261 ( .A(n22855), .B(n19727), .Z(n19728) );
  NANDN U39262 ( .A(n59571), .B(n19728), .Z(n19729) );
  AND U39263 ( .A(n59573), .B(n19729), .Z(n19731) );
  XNOR U39264 ( .A(x[6812]), .B(y[6812]), .Z(n47107) );
  NANDN U39265 ( .A(x[6811]), .B(y[6811]), .Z(n59574) );
  AND U39266 ( .A(n47107), .B(n59574), .Z(n19730) );
  NANDN U39267 ( .A(n19731), .B(n19730), .Z(n19732) );
  NANDN U39268 ( .A(n59576), .B(n19732), .Z(n19733) );
  AND U39269 ( .A(n22853), .B(n19733), .Z(n19734) );
  NANDN U39270 ( .A(n59577), .B(n19734), .Z(n19735) );
  AND U39271 ( .A(n59579), .B(n19735), .Z(n19737) );
  XNOR U39272 ( .A(x[6816]), .B(y[6816]), .Z(n22851) );
  NANDN U39273 ( .A(x[6815]), .B(y[6815]), .Z(n59581) );
  AND U39274 ( .A(n22851), .B(n59581), .Z(n19736) );
  NANDN U39275 ( .A(n19737), .B(n19736), .Z(n19738) );
  NANDN U39276 ( .A(n59583), .B(n19738), .Z(n19739) );
  AND U39277 ( .A(n59584), .B(n19739), .Z(n19740) );
  NAND U39278 ( .A(n22849), .B(n19740), .Z(n19741) );
  NAND U39279 ( .A(n59586), .B(n19741), .Z(n19742) );
  AND U39280 ( .A(n47125), .B(n19742), .Z(n19743) );
  NANDN U39281 ( .A(x[6819]), .B(y[6819]), .Z(n59587) );
  AND U39282 ( .A(n19743), .B(n59587), .Z(n19745) );
  NANDN U39283 ( .A(y[6820]), .B(x[6820]), .Z(n19744) );
  NANDN U39284 ( .A(y[6821]), .B(x[6821]), .Z(n22845) );
  NAND U39285 ( .A(n19744), .B(n22845), .Z(n59589) );
  OR U39286 ( .A(n19745), .B(n59589), .Z(n19746) );
  NAND U39287 ( .A(n19747), .B(n19746), .Z(n19748) );
  NAND U39288 ( .A(n59590), .B(n19748), .Z(n19749) );
  AND U39289 ( .A(n47135), .B(n19749), .Z(n19750) );
  NANDN U39290 ( .A(x[6823]), .B(y[6823]), .Z(n59591) );
  AND U39291 ( .A(n19750), .B(n59591), .Z(n19751) );
  OR U39292 ( .A(n59593), .B(n19751), .Z(n19752) );
  NAND U39293 ( .A(n19753), .B(n19752), .Z(n19754) );
  NANDN U39294 ( .A(n59596), .B(n19754), .Z(n19755) );
  AND U39295 ( .A(n47145), .B(n19755), .Z(n19756) );
  NANDN U39296 ( .A(x[6827]), .B(y[6827]), .Z(n59598) );
  NAND U39297 ( .A(n19756), .B(n59598), .Z(n19757) );
  AND U39298 ( .A(n59600), .B(n19757), .Z(n19759) );
  XNOR U39299 ( .A(x[6830]), .B(y[6830]), .Z(n22842) );
  ANDN U39300 ( .B(y[6829]), .A(x[6829]), .Z(n59601) );
  ANDN U39301 ( .B(n22842), .A(n59601), .Z(n19758) );
  NANDN U39302 ( .A(n19759), .B(n19758), .Z(n19760) );
  NANDN U39303 ( .A(n59603), .B(n19760), .Z(n19761) );
  AND U39304 ( .A(n47156), .B(n19761), .Z(n19762) );
  NANDN U39305 ( .A(n50950), .B(n19762), .Z(n19763) );
  NAND U39306 ( .A(n59604), .B(n19763), .Z(n19764) );
  AND U39307 ( .A(n22840), .B(n19764), .Z(n19765) );
  ANDN U39308 ( .B(y[6833]), .A(x[6833]), .Z(n59605) );
  ANDN U39309 ( .B(n19765), .A(n59605), .Z(n19767) );
  NANDN U39310 ( .A(y[6834]), .B(x[6834]), .Z(n19766) );
  NANDN U39311 ( .A(y[6835]), .B(x[6835]), .Z(n47166) );
  AND U39312 ( .A(n19766), .B(n47166), .Z(n59607) );
  NANDN U39313 ( .A(n19767), .B(n59607), .Z(n19768) );
  NAND U39314 ( .A(n19769), .B(n19768), .Z(n19770) );
  NAND U39315 ( .A(n59608), .B(n19770), .Z(n19771) );
  AND U39316 ( .A(n59609), .B(n19771), .Z(n19773) );
  NANDN U39317 ( .A(y[6838]), .B(x[6838]), .Z(n19772) );
  NANDN U39318 ( .A(y[6839]), .B(x[6839]), .Z(n47177) );
  NAND U39319 ( .A(n19772), .B(n47177), .Z(n59610) );
  OR U39320 ( .A(n19773), .B(n59610), .Z(n19774) );
  NAND U39321 ( .A(n19775), .B(n19774), .Z(n19776) );
  NANDN U39322 ( .A(n50944), .B(n19776), .Z(n19777) );
  AND U39323 ( .A(n22835), .B(n19777), .Z(n19778) );
  NANDN U39324 ( .A(n50943), .B(n19778), .Z(n19779) );
  NAND U39325 ( .A(n59613), .B(n19779), .Z(n19780) );
  AND U39326 ( .A(n22833), .B(n19780), .Z(n19781) );
  NANDN U39327 ( .A(x[6843]), .B(y[6843]), .Z(n59614) );
  NAND U39328 ( .A(n19781), .B(n59614), .Z(n19782) );
  NANDN U39329 ( .A(n59616), .B(n19782), .Z(n19783) );
  AND U39330 ( .A(n22831), .B(n19783), .Z(n19784) );
  NANDN U39331 ( .A(x[6845]), .B(y[6845]), .Z(n50940) );
  NAND U39332 ( .A(n19784), .B(n50940), .Z(n19786) );
  NANDN U39333 ( .A(y[6846]), .B(x[6846]), .Z(n19785) );
  NANDN U39334 ( .A(y[6847]), .B(x[6847]), .Z(n47195) );
  AND U39335 ( .A(n19785), .B(n47195), .Z(n50939) );
  AND U39336 ( .A(n19786), .B(n50939), .Z(n19787) );
  OR U39337 ( .A(n19788), .B(n19787), .Z(n19789) );
  NAND U39338 ( .A(n59619), .B(n19789), .Z(n19790) );
  NANDN U39339 ( .A(n19791), .B(n19790), .Z(n19792) );
  NAND U39340 ( .A(n59622), .B(n19792), .Z(n19793) );
  AND U39341 ( .A(n22827), .B(n19793), .Z(n19794) );
  NANDN U39342 ( .A(x[6851]), .B(y[6851]), .Z(n59623) );
  AND U39343 ( .A(n19794), .B(n59623), .Z(n19796) );
  NANDN U39344 ( .A(y[6852]), .B(x[6852]), .Z(n19795) );
  NANDN U39345 ( .A(y[6853]), .B(x[6853]), .Z(n22824) );
  AND U39346 ( .A(n19795), .B(n22824), .Z(n59626) );
  NANDN U39347 ( .A(n19796), .B(n59626), .Z(n19797) );
  NAND U39348 ( .A(n59627), .B(n19797), .Z(n19798) );
  NANDN U39349 ( .A(n59628), .B(n19798), .Z(n19799) );
  AND U39350 ( .A(n22822), .B(n19799), .Z(n19800) );
  NANDN U39351 ( .A(x[6855]), .B(y[6855]), .Z(n50937) );
  AND U39352 ( .A(n19800), .B(n50937), .Z(n19802) );
  NANDN U39353 ( .A(y[6856]), .B(x[6856]), .Z(n19801) );
  NANDN U39354 ( .A(y[6857]), .B(x[6857]), .Z(n22819) );
  AND U39355 ( .A(n19801), .B(n22819), .Z(n59629) );
  NANDN U39356 ( .A(n19802), .B(n59629), .Z(n19803) );
  AND U39357 ( .A(n59630), .B(n19803), .Z(n19804) );
  NAND U39358 ( .A(n22820), .B(n19804), .Z(n19805) );
  NANDN U39359 ( .A(n59632), .B(n19805), .Z(n19806) );
  NAND U39360 ( .A(n19807), .B(n19806), .Z(n19808) );
  NAND U39361 ( .A(n59633), .B(n19808), .Z(n19809) );
  AND U39362 ( .A(n22818), .B(n19809), .Z(n19810) );
  ANDN U39363 ( .B(y[6861]), .A(x[6861]), .Z(n59634) );
  ANDN U39364 ( .B(n19810), .A(n59634), .Z(n19812) );
  NANDN U39365 ( .A(y[6862]), .B(x[6862]), .Z(n19811) );
  NANDN U39366 ( .A(y[6863]), .B(x[6863]), .Z(n22815) );
  AND U39367 ( .A(n19811), .B(n22815), .Z(n59636) );
  NANDN U39368 ( .A(n19812), .B(n59636), .Z(n19813) );
  NAND U39369 ( .A(n19814), .B(n19813), .Z(n19815) );
  NANDN U39370 ( .A(n59639), .B(n19815), .Z(n19816) );
  AND U39371 ( .A(n22814), .B(n19816), .Z(n19817) );
  NANDN U39372 ( .A(x[6865]), .B(y[6865]), .Z(n59641) );
  NAND U39373 ( .A(n19817), .B(n59641), .Z(n19818) );
  AND U39374 ( .A(n59643), .B(n19818), .Z(n19820) );
  XNOR U39375 ( .A(x[6868]), .B(y[6868]), .Z(n47241) );
  NANDN U39376 ( .A(x[6867]), .B(y[6867]), .Z(n59644) );
  AND U39377 ( .A(n47241), .B(n59644), .Z(n19819) );
  NANDN U39378 ( .A(n19820), .B(n19819), .Z(n19821) );
  NANDN U39379 ( .A(n59646), .B(n19821), .Z(n19822) );
  AND U39380 ( .A(n22812), .B(n19822), .Z(n19823) );
  NANDN U39381 ( .A(x[6869]), .B(y[6869]), .Z(n50934) );
  NAND U39382 ( .A(n19823), .B(n50934), .Z(n19824) );
  AND U39383 ( .A(n59647), .B(n19824), .Z(n19825) );
  OR U39384 ( .A(n19826), .B(n19825), .Z(n19827) );
  NAND U39385 ( .A(n59650), .B(n19827), .Z(n19828) );
  NANDN U39386 ( .A(n19829), .B(n19828), .Z(n19830) );
  NAND U39387 ( .A(n59651), .B(n19830), .Z(n19831) );
  AND U39388 ( .A(n22808), .B(n19831), .Z(n19832) );
  NANDN U39389 ( .A(x[6875]), .B(y[6875]), .Z(n59652) );
  AND U39390 ( .A(n19832), .B(n59652), .Z(n19834) );
  NANDN U39391 ( .A(y[6876]), .B(x[6876]), .Z(n19833) );
  NANDN U39392 ( .A(y[6877]), .B(x[6877]), .Z(n22805) );
  AND U39393 ( .A(n19833), .B(n22805), .Z(n59655) );
  NANDN U39394 ( .A(n19834), .B(n59655), .Z(n19835) );
  NAND U39395 ( .A(n19836), .B(n19835), .Z(n19837) );
  NANDN U39396 ( .A(n59658), .B(n19837), .Z(n19838) );
  AND U39397 ( .A(n47269), .B(n19838), .Z(n19839) );
  NANDN U39398 ( .A(x[6879]), .B(y[6879]), .Z(n59659) );
  NAND U39399 ( .A(n19839), .B(n59659), .Z(n19840) );
  AND U39400 ( .A(n59661), .B(n19840), .Z(n19842) );
  XNOR U39401 ( .A(x[6882]), .B(y[6882]), .Z(n22804) );
  ANDN U39402 ( .B(y[6881]), .A(x[6881]), .Z(n59662) );
  ANDN U39403 ( .B(n22804), .A(n59662), .Z(n19841) );
  NANDN U39404 ( .A(n19842), .B(n19841), .Z(n19843) );
  NANDN U39405 ( .A(n59664), .B(n19843), .Z(n19844) );
  AND U39406 ( .A(n47280), .B(n19844), .Z(n19845) );
  NANDN U39407 ( .A(n50930), .B(n19845), .Z(n19846) );
  NAND U39408 ( .A(n59665), .B(n19846), .Z(n19847) );
  AND U39409 ( .A(n22802), .B(n19847), .Z(n19848) );
  ANDN U39410 ( .B(y[6885]), .A(x[6885]), .Z(n59666) );
  ANDN U39411 ( .B(n19848), .A(n59666), .Z(n19850) );
  NANDN U39412 ( .A(y[6886]), .B(x[6886]), .Z(n19849) );
  NANDN U39413 ( .A(y[6887]), .B(x[6887]), .Z(n47290) );
  AND U39414 ( .A(n19849), .B(n47290), .Z(n59668) );
  NANDN U39415 ( .A(n19850), .B(n59668), .Z(n19851) );
  NAND U39416 ( .A(n19852), .B(n19851), .Z(n19854) );
  NANDN U39417 ( .A(y[6888]), .B(x[6888]), .Z(n19853) );
  NANDN U39418 ( .A(y[6889]), .B(x[6889]), .Z(n22799) );
  AND U39419 ( .A(n19853), .B(n22799), .Z(n50926) );
  AND U39420 ( .A(n19854), .B(n50926), .Z(n19856) );
  XNOR U39421 ( .A(x[6890]), .B(y[6890]), .Z(n22800) );
  ANDN U39422 ( .B(y[6889]), .A(x[6889]), .Z(n59671) );
  ANDN U39423 ( .B(n22800), .A(n59671), .Z(n19855) );
  NANDN U39424 ( .A(n19856), .B(n19855), .Z(n19857) );
  NAND U39425 ( .A(n59673), .B(n19857), .Z(n19858) );
  AND U39426 ( .A(n47301), .B(n19858), .Z(n19859) );
  NANDN U39427 ( .A(x[6891]), .B(y[6891]), .Z(n59674) );
  NAND U39428 ( .A(n19859), .B(n59674), .Z(n19860) );
  NANDN U39429 ( .A(n59675), .B(n19860), .Z(n19861) );
  AND U39430 ( .A(n22798), .B(n19861), .Z(n19862) );
  NANDN U39431 ( .A(n59676), .B(n19862), .Z(n19863) );
  AND U39432 ( .A(n59678), .B(n19863), .Z(n19864) );
  OR U39433 ( .A(n19865), .B(n19864), .Z(n19866) );
  NAND U39434 ( .A(n59681), .B(n19866), .Z(n19867) );
  NANDN U39435 ( .A(n19868), .B(n19867), .Z(n19869) );
  NAND U39436 ( .A(n59682), .B(n19869), .Z(n19870) );
  AND U39437 ( .A(n47321), .B(n19870), .Z(n19871) );
  NANDN U39438 ( .A(x[6899]), .B(y[6899]), .Z(n59683) );
  AND U39439 ( .A(n19871), .B(n59683), .Z(n19872) );
  OR U39440 ( .A(n59687), .B(n19872), .Z(n19873) );
  NAND U39441 ( .A(n59688), .B(n19873), .Z(n19874) );
  NANDN U39442 ( .A(n59689), .B(n19874), .Z(n19875) );
  AND U39443 ( .A(n47331), .B(n19875), .Z(n19876) );
  NANDN U39444 ( .A(x[6903]), .B(y[6903]), .Z(n59690) );
  NAND U39445 ( .A(n19876), .B(n59690), .Z(n19877) );
  NAND U39446 ( .A(n59692), .B(n19877), .Z(n19878) );
  AND U39447 ( .A(n22789), .B(n19878), .Z(n19879) );
  NANDN U39448 ( .A(x[6905]), .B(y[6905]), .Z(n22790) );
  AND U39449 ( .A(n19879), .B(n22790), .Z(n19881) );
  NANDN U39450 ( .A(y[6906]), .B(x[6906]), .Z(n19880) );
  NANDN U39451 ( .A(y[6907]), .B(x[6907]), .Z(n47341) );
  NAND U39452 ( .A(n19880), .B(n47341), .Z(n59693) );
  OR U39453 ( .A(n19881), .B(n59693), .Z(n19882) );
  AND U39454 ( .A(n47342), .B(n19882), .Z(n19883) );
  NANDN U39455 ( .A(n59695), .B(n19883), .Z(n19885) );
  NANDN U39456 ( .A(y[6908]), .B(x[6908]), .Z(n19884) );
  NANDN U39457 ( .A(y[6909]), .B(x[6909]), .Z(n22786) );
  AND U39458 ( .A(n19884), .B(n22786), .Z(n50920) );
  AND U39459 ( .A(n19885), .B(n50920), .Z(n19886) );
  OR U39460 ( .A(n19887), .B(n19886), .Z(n19888) );
  NAND U39461 ( .A(n59698), .B(n19888), .Z(n19889) );
  NANDN U39462 ( .A(n19890), .B(n19889), .Z(n19891) );
  NAND U39463 ( .A(n59703), .B(n19891), .Z(n19892) );
  AND U39464 ( .A(n22785), .B(n19892), .Z(n19893) );
  ANDN U39465 ( .B(y[6913]), .A(x[6913]), .Z(n50918) );
  ANDN U39466 ( .B(n19893), .A(n50918), .Z(n19895) );
  NANDN U39467 ( .A(y[6914]), .B(x[6914]), .Z(n19894) );
  NANDN U39468 ( .A(y[6915]), .B(x[6915]), .Z(n47361) );
  NAND U39469 ( .A(n19894), .B(n47361), .Z(n59704) );
  OR U39470 ( .A(n19895), .B(n59704), .Z(n19896) );
  NAND U39471 ( .A(n19897), .B(n19896), .Z(n19898) );
  NANDN U39472 ( .A(n59707), .B(n19898), .Z(n19899) );
  AND U39473 ( .A(n22783), .B(n19899), .Z(n19900) );
  NANDN U39474 ( .A(n59708), .B(n19900), .Z(n19902) );
  NANDN U39475 ( .A(y[6918]), .B(x[6918]), .Z(n19901) );
  NANDN U39476 ( .A(y[6919]), .B(x[6919]), .Z(n47371) );
  AND U39477 ( .A(n19901), .B(n47371), .Z(n59710) );
  AND U39478 ( .A(n19902), .B(n59710), .Z(n19904) );
  XNOR U39479 ( .A(x[6920]), .B(y[6920]), .Z(n47372) );
  NANDN U39480 ( .A(x[6919]), .B(y[6919]), .Z(n59711) );
  AND U39481 ( .A(n47372), .B(n59711), .Z(n19903) );
  NANDN U39482 ( .A(n19904), .B(n19903), .Z(n19905) );
  NAND U39483 ( .A(n59713), .B(n19905), .Z(n19906) );
  AND U39484 ( .A(n22781), .B(n19906), .Z(n19907) );
  NANDN U39485 ( .A(n59714), .B(n19907), .Z(n19908) );
  AND U39486 ( .A(n59716), .B(n19908), .Z(n19910) );
  XNOR U39487 ( .A(x[6924]), .B(y[6924]), .Z(n47382) );
  NANDN U39488 ( .A(x[6923]), .B(y[6923]), .Z(n50915) );
  AND U39489 ( .A(n47382), .B(n50915), .Z(n19909) );
  NANDN U39490 ( .A(n19910), .B(n19909), .Z(n19911) );
  NAND U39491 ( .A(n59718), .B(n19911), .Z(n19912) );
  ANDN U39492 ( .B(y[6925]), .A(x[6925]), .Z(n59719) );
  ANDN U39493 ( .B(n19912), .A(n59719), .Z(n19913) );
  NAND U39494 ( .A(n22779), .B(n19913), .Z(n19914) );
  NAND U39495 ( .A(n59721), .B(n19914), .Z(n19915) );
  AND U39496 ( .A(n22777), .B(n19915), .Z(n19916) );
  NANDN U39497 ( .A(x[6927]), .B(y[6927]), .Z(n50913) );
  AND U39498 ( .A(n19916), .B(n50913), .Z(n19917) );
  OR U39499 ( .A(n59722), .B(n19917), .Z(n19918) );
  NAND U39500 ( .A(n19919), .B(n19918), .Z(n19920) );
  NAND U39501 ( .A(n59725), .B(n19920), .Z(n19921) );
  AND U39502 ( .A(n47400), .B(n19921), .Z(n19922) );
  NANDN U39503 ( .A(x[6931]), .B(y[6931]), .Z(n59726) );
  NAND U39504 ( .A(n19922), .B(n59726), .Z(n19924) );
  NANDN U39505 ( .A(y[6932]), .B(x[6932]), .Z(n19923) );
  NANDN U39506 ( .A(y[6933]), .B(x[6933]), .Z(n22772) );
  AND U39507 ( .A(n19923), .B(n22772), .Z(n50911) );
  AND U39508 ( .A(n19924), .B(n50911), .Z(n19926) );
  XNOR U39509 ( .A(x[6934]), .B(y[6934]), .Z(n22773) );
  ANDN U39510 ( .B(y[6933]), .A(x[6933]), .Z(n59727) );
  ANDN U39511 ( .B(n22773), .A(n59727), .Z(n19925) );
  NANDN U39512 ( .A(n19926), .B(n19925), .Z(n19927) );
  NAND U39513 ( .A(n59729), .B(n19927), .Z(n19928) );
  AND U39514 ( .A(n47410), .B(n19928), .Z(n19929) );
  NANDN U39515 ( .A(x[6935]), .B(y[6935]), .Z(n59731) );
  NAND U39516 ( .A(n19929), .B(n59731), .Z(n19930) );
  NAND U39517 ( .A(n59734), .B(n19930), .Z(n19931) );
  NAND U39518 ( .A(n22771), .B(n19931), .Z(n19932) );
  ANDN U39519 ( .B(y[6937]), .A(x[6937]), .Z(n50910) );
  OR U39520 ( .A(n19932), .B(n50910), .Z(n19933) );
  NAND U39521 ( .A(n59735), .B(n19933), .Z(n19934) );
  NAND U39522 ( .A(n59736), .B(n19934), .Z(n19935) );
  NAND U39523 ( .A(n59737), .B(n19935), .Z(n19936) );
  AND U39524 ( .A(n22768), .B(n19936), .Z(n19937) );
  NANDN U39525 ( .A(x[6941]), .B(y[6941]), .Z(n59739) );
  AND U39526 ( .A(n19937), .B(n59739), .Z(n19939) );
  NANDN U39527 ( .A(y[6942]), .B(x[6942]), .Z(n19938) );
  NANDN U39528 ( .A(y[6943]), .B(x[6943]), .Z(n47430) );
  NAND U39529 ( .A(n19938), .B(n47430), .Z(n59740) );
  OR U39530 ( .A(n19939), .B(n59740), .Z(n19940) );
  NAND U39531 ( .A(n19941), .B(n19940), .Z(n19942) );
  NAND U39532 ( .A(n59743), .B(n19942), .Z(n19943) );
  AND U39533 ( .A(n22766), .B(n19943), .Z(n19944) );
  ANDN U39534 ( .B(y[6945]), .A(x[6945]), .Z(n59744) );
  ANDN U39535 ( .B(n19944), .A(n59744), .Z(n19945) );
  OR U39536 ( .A(n59746), .B(n19945), .Z(n19946) );
  NAND U39537 ( .A(n19947), .B(n19946), .Z(n19948) );
  NAND U39538 ( .A(n59750), .B(n19948), .Z(n19949) );
  AND U39539 ( .A(n22764), .B(n19949), .Z(n19950) );
  NANDN U39540 ( .A(n59751), .B(n19950), .Z(n19951) );
  AND U39541 ( .A(n59753), .B(n19951), .Z(n19953) );
  XNOR U39542 ( .A(x[6952]), .B(y[6952]), .Z(n47451) );
  NANDN U39543 ( .A(x[6951]), .B(y[6951]), .Z(n50907) );
  AND U39544 ( .A(n47451), .B(n50907), .Z(n19952) );
  NANDN U39545 ( .A(n19953), .B(n19952), .Z(n19954) );
  NAND U39546 ( .A(n59754), .B(n19954), .Z(n19955) );
  AND U39547 ( .A(n22762), .B(n19955), .Z(n19956) );
  NANDN U39548 ( .A(n59755), .B(n19956), .Z(n19957) );
  NAND U39549 ( .A(n59757), .B(n19957), .Z(n19958) );
  AND U39550 ( .A(n59758), .B(n19958), .Z(n19959) );
  OR U39551 ( .A(n59759), .B(n19959), .Z(n19960) );
  NAND U39552 ( .A(n19961), .B(n19960), .Z(n19962) );
  NAND U39553 ( .A(n59762), .B(n19962), .Z(n19963) );
  AND U39554 ( .A(n47472), .B(n19963), .Z(n19964) );
  NANDN U39555 ( .A(x[6959]), .B(y[6959]), .Z(n50906) );
  AND U39556 ( .A(n19964), .B(n50906), .Z(n19966) );
  NANDN U39557 ( .A(y[6960]), .B(x[6960]), .Z(n19965) );
  NANDN U39558 ( .A(y[6961]), .B(x[6961]), .Z(n22756) );
  NAND U39559 ( .A(n19965), .B(n22756), .Z(n50904) );
  OR U39560 ( .A(n19966), .B(n50904), .Z(n19967) );
  NAND U39561 ( .A(n19968), .B(n19967), .Z(n19969) );
  NAND U39562 ( .A(n59764), .B(n19969), .Z(n19970) );
  AND U39563 ( .A(n47482), .B(n19970), .Z(n19971) );
  NANDN U39564 ( .A(x[6963]), .B(y[6963]), .Z(n59765) );
  AND U39565 ( .A(n19971), .B(n59765), .Z(n19972) );
  OR U39566 ( .A(n59767), .B(n19972), .Z(n19973) );
  NAND U39567 ( .A(n19974), .B(n19973), .Z(n19975) );
  NANDN U39568 ( .A(n59768), .B(n19975), .Z(n19976) );
  AND U39569 ( .A(n47492), .B(n19976), .Z(n19977) );
  NANDN U39570 ( .A(x[6967]), .B(y[6967]), .Z(n59769) );
  AND U39571 ( .A(n19977), .B(n59769), .Z(n19979) );
  NANDN U39572 ( .A(y[6968]), .B(x[6968]), .Z(n19978) );
  NANDN U39573 ( .A(y[6969]), .B(x[6969]), .Z(n22752) );
  AND U39574 ( .A(n19978), .B(n22752), .Z(n59771) );
  NANDN U39575 ( .A(n19979), .B(n59771), .Z(n19980) );
  NAND U39576 ( .A(n19981), .B(n19980), .Z(n19982) );
  NANDN U39577 ( .A(n59774), .B(n19982), .Z(n19983) );
  AND U39578 ( .A(n47502), .B(n19983), .Z(n19984) );
  NANDN U39579 ( .A(x[6971]), .B(y[6971]), .Z(n59775) );
  NAND U39580 ( .A(n19984), .B(n59775), .Z(n19985) );
  NAND U39581 ( .A(n59778), .B(n19985), .Z(n19986) );
  AND U39582 ( .A(n22751), .B(n19986), .Z(n19987) );
  ANDN U39583 ( .B(y[6973]), .A(x[6973]), .Z(n59779) );
  ANDN U39584 ( .B(n19987), .A(n59779), .Z(n19989) );
  NANDN U39585 ( .A(y[6974]), .B(x[6974]), .Z(n19988) );
  NANDN U39586 ( .A(y[6975]), .B(x[6975]), .Z(n22748) );
  NAND U39587 ( .A(n19988), .B(n22748), .Z(n59781) );
  OR U39588 ( .A(n19989), .B(n59781), .Z(n19990) );
  NAND U39589 ( .A(n19991), .B(n19990), .Z(n19992) );
  NAND U39590 ( .A(n59782), .B(n19992), .Z(n19993) );
  AND U39591 ( .A(n22747), .B(n19993), .Z(n19994) );
  NANDN U39592 ( .A(x[6977]), .B(y[6977]), .Z(n59783) );
  AND U39593 ( .A(n19994), .B(n59783), .Z(n19996) );
  NANDN U39594 ( .A(y[6978]), .B(x[6978]), .Z(n19995) );
  NANDN U39595 ( .A(y[6979]), .B(x[6979]), .Z(n47519) );
  NAND U39596 ( .A(n19995), .B(n47519), .Z(n59785) );
  OR U39597 ( .A(n19996), .B(n59785), .Z(n19997) );
  AND U39598 ( .A(n19998), .B(n19997), .Z(n19999) );
  OR U39599 ( .A(n59786), .B(n19999), .Z(n20000) );
  NAND U39600 ( .A(n20001), .B(n20000), .Z(n20002) );
  AND U39601 ( .A(n59789), .B(n20002), .Z(n20004) );
  XNOR U39602 ( .A(x[6984]), .B(y[6984]), .Z(n47530) );
  NANDN U39603 ( .A(x[6983]), .B(y[6983]), .Z(n59790) );
  AND U39604 ( .A(n47530), .B(n59790), .Z(n20003) );
  NANDN U39605 ( .A(n20004), .B(n20003), .Z(n20005) );
  NANDN U39606 ( .A(n59793), .B(n20005), .Z(n20006) );
  AND U39607 ( .A(n22743), .B(n20006), .Z(n20007) );
  NANDN U39608 ( .A(n59794), .B(n20007), .Z(n20008) );
  NAND U39609 ( .A(n59796), .B(n20008), .Z(n20009) );
  AND U39610 ( .A(n47540), .B(n20009), .Z(n20010) );
  NANDN U39611 ( .A(x[6987]), .B(y[6987]), .Z(n59797) );
  AND U39612 ( .A(n20010), .B(n59797), .Z(n20012) );
  NANDN U39613 ( .A(y[6988]), .B(x[6988]), .Z(n20011) );
  NANDN U39614 ( .A(y[6989]), .B(x[6989]), .Z(n22740) );
  AND U39615 ( .A(n20011), .B(n22740), .Z(n59799) );
  NANDN U39616 ( .A(n20012), .B(n59799), .Z(n20013) );
  NAND U39617 ( .A(n20014), .B(n20013), .Z(n20015) );
  AND U39618 ( .A(n59800), .B(n20015), .Z(n20017) );
  XNOR U39619 ( .A(x[6992]), .B(y[6992]), .Z(n47550) );
  NANDN U39620 ( .A(x[6991]), .B(y[6991]), .Z(n59801) );
  AND U39621 ( .A(n47550), .B(n59801), .Z(n20016) );
  NANDN U39622 ( .A(n20017), .B(n20016), .Z(n20018) );
  NANDN U39623 ( .A(n59803), .B(n20018), .Z(n20019) );
  AND U39624 ( .A(n22739), .B(n20019), .Z(n20020) );
  NANDN U39625 ( .A(x[6995]), .B(y[6995]), .Z(n59806) );
  NANDN U39626 ( .A(x[6997]), .B(y[6997]), .Z(n22735) );
  NANDN U39627 ( .A(x[6998]), .B(y[6998]), .Z(n22732) );
  AND U39628 ( .A(n22735), .B(n22732), .Z(n50889) );
  ANDN U39629 ( .B(x[6999]), .A(y[6999]), .Z(n47568) );
  NANDN U39630 ( .A(y[6998]), .B(x[6998]), .Z(n22733) );
  NANDN U39631 ( .A(n47568), .B(n22733), .Z(n59808) );
  NANDN U39632 ( .A(x[7001]), .B(y[7001]), .Z(n59812) );
  NANDN U39633 ( .A(y[7002]), .B(x[7002]), .Z(n20021) );
  NANDN U39634 ( .A(y[7003]), .B(x[7003]), .Z(n22728) );
  NAND U39635 ( .A(n20021), .B(n22728), .Z(n59814) );
  NANDN U39636 ( .A(x[7005]), .B(y[7005]), .Z(n50887) );
  NANDN U39637 ( .A(y[7006]), .B(x[7006]), .Z(n20022) );
  NANDN U39638 ( .A(y[7007]), .B(x[7007]), .Z(n47585) );
  NAND U39639 ( .A(n20022), .B(n47585), .Z(n59818) );
  NAND U39640 ( .A(n20024), .B(n20023), .Z(n20025) );
  NANDN U39641 ( .A(n59824), .B(n20025), .Z(n20026) );
  AND U39642 ( .A(n22725), .B(n20026), .Z(n20027) );
  NANDN U39643 ( .A(n59825), .B(n20027), .Z(n20029) );
  NANDN U39644 ( .A(y[7010]), .B(x[7010]), .Z(n20028) );
  NANDN U39645 ( .A(y[7011]), .B(x[7011]), .Z(n47595) );
  AND U39646 ( .A(n20028), .B(n47595), .Z(n59827) );
  AND U39647 ( .A(n20029), .B(n59827), .Z(n20031) );
  XNOR U39648 ( .A(x[7012]), .B(y[7012]), .Z(n47596) );
  NANDN U39649 ( .A(x[7011]), .B(y[7011]), .Z(n59828) );
  AND U39650 ( .A(n47596), .B(n59828), .Z(n20030) );
  NANDN U39651 ( .A(n20031), .B(n20030), .Z(n20032) );
  NAND U39652 ( .A(n59830), .B(n20032), .Z(n20033) );
  AND U39653 ( .A(n22723), .B(n20033), .Z(n20034) );
  ANDN U39654 ( .B(y[7013]), .A(x[7013]), .Z(n59831) );
  ANDN U39655 ( .B(n20034), .A(n59831), .Z(n20036) );
  NANDN U39656 ( .A(y[7014]), .B(x[7014]), .Z(n20035) );
  NANDN U39657 ( .A(y[7015]), .B(x[7015]), .Z(n47605) );
  AND U39658 ( .A(n20035), .B(n47605), .Z(n59833) );
  NANDN U39659 ( .A(n20036), .B(n59833), .Z(n20037) );
  NAND U39660 ( .A(n20038), .B(n20037), .Z(n20039) );
  NAND U39661 ( .A(n59834), .B(n20039), .Z(n20040) );
  AND U39662 ( .A(n22721), .B(n20040), .Z(n20041) );
  NANDN U39663 ( .A(n59835), .B(n20041), .Z(n20042) );
  NANDN U39664 ( .A(n59837), .B(n20042), .Z(n20043) );
  AND U39665 ( .A(n47616), .B(n20043), .Z(n20044) );
  NANDN U39666 ( .A(x[7019]), .B(y[7019]), .Z(n50884) );
  NAND U39667 ( .A(n20044), .B(n50884), .Z(n20046) );
  NANDN U39668 ( .A(y[7020]), .B(x[7020]), .Z(n20045) );
  NANDN U39669 ( .A(y[7021]), .B(x[7021]), .Z(n22718) );
  AND U39670 ( .A(n20045), .B(n22718), .Z(n50881) );
  AND U39671 ( .A(n20046), .B(n50881), .Z(n20048) );
  XNOR U39672 ( .A(x[7022]), .B(y[7022]), .Z(n22719) );
  ANDN U39673 ( .B(y[7021]), .A(x[7021]), .Z(n59839) );
  ANDN U39674 ( .B(n22719), .A(n59839), .Z(n20047) );
  NANDN U39675 ( .A(n20048), .B(n20047), .Z(n20049) );
  NAND U39676 ( .A(n59841), .B(n20049), .Z(n20050) );
  AND U39677 ( .A(n47626), .B(n20050), .Z(n20051) );
  NANDN U39678 ( .A(x[7023]), .B(y[7023]), .Z(n59842) );
  NAND U39679 ( .A(n20051), .B(n59842), .Z(n20053) );
  NANDN U39680 ( .A(y[7024]), .B(x[7024]), .Z(n20052) );
  NANDN U39681 ( .A(y[7025]), .B(x[7025]), .Z(n22716) );
  AND U39682 ( .A(n20052), .B(n22716), .Z(n50879) );
  AND U39683 ( .A(n20053), .B(n50879), .Z(n20054) );
  OR U39684 ( .A(n20055), .B(n20054), .Z(n20056) );
  NAND U39685 ( .A(n59845), .B(n20056), .Z(n20057) );
  NANDN U39686 ( .A(n20058), .B(n20057), .Z(n20059) );
  NAND U39687 ( .A(n59848), .B(n20059), .Z(n20060) );
  AND U39688 ( .A(n22714), .B(n20060), .Z(n20061) );
  NANDN U39689 ( .A(x[7029]), .B(y[7029]), .Z(n22715) );
  AND U39690 ( .A(n20061), .B(n22715), .Z(n20063) );
  NANDN U39691 ( .A(y[7030]), .B(x[7030]), .Z(n20062) );
  NANDN U39692 ( .A(y[7031]), .B(x[7031]), .Z(n47645) );
  AND U39693 ( .A(n20062), .B(n47645), .Z(n59850) );
  NANDN U39694 ( .A(n20063), .B(n59850), .Z(n20064) );
  NAND U39695 ( .A(n20065), .B(n20064), .Z(n20066) );
  NANDN U39696 ( .A(n59853), .B(n20066), .Z(n20067) );
  AND U39697 ( .A(n22712), .B(n20067), .Z(n20068) );
  NANDN U39698 ( .A(n50875), .B(n20068), .Z(n20070) );
  NANDN U39699 ( .A(y[7034]), .B(x[7034]), .Z(n20069) );
  NANDN U39700 ( .A(y[7035]), .B(x[7035]), .Z(n47655) );
  AND U39701 ( .A(n20069), .B(n47655), .Z(n50874) );
  AND U39702 ( .A(n20070), .B(n50874), .Z(n20072) );
  XNOR U39703 ( .A(x[7036]), .B(y[7036]), .Z(n47656) );
  NANDN U39704 ( .A(x[7035]), .B(y[7035]), .Z(n59854) );
  AND U39705 ( .A(n47656), .B(n59854), .Z(n20071) );
  NANDN U39706 ( .A(n20072), .B(n20071), .Z(n20073) );
  NAND U39707 ( .A(n59856), .B(n20073), .Z(n20074) );
  AND U39708 ( .A(n22710), .B(n20074), .Z(n20075) );
  NANDN U39709 ( .A(n59857), .B(n20075), .Z(n20076) );
  NAND U39710 ( .A(n59859), .B(n20076), .Z(n20077) );
  NAND U39711 ( .A(n47667), .B(n20077), .Z(n20078) );
  ANDN U39712 ( .B(y[7039]), .A(x[7039]), .Z(n47663) );
  OR U39713 ( .A(n20078), .B(n47663), .Z(n20079) );
  NAND U39714 ( .A(n59862), .B(n20079), .Z(n20080) );
  NANDN U39715 ( .A(n59863), .B(n20080), .Z(n20081) );
  NAND U39716 ( .A(n59864), .B(n20081), .Z(n20082) );
  AND U39717 ( .A(n47678), .B(n20082), .Z(n20083) );
  NANDN U39718 ( .A(x[7043]), .B(y[7043]), .Z(n50873) );
  AND U39719 ( .A(n20083), .B(n50873), .Z(n20085) );
  NANDN U39720 ( .A(y[7044]), .B(x[7044]), .Z(n20084) );
  NANDN U39721 ( .A(y[7045]), .B(x[7045]), .Z(n22704) );
  AND U39722 ( .A(n20084), .B(n22704), .Z(n59866) );
  NANDN U39723 ( .A(n20085), .B(n59866), .Z(n20086) );
  NAND U39724 ( .A(n20087), .B(n20086), .Z(n20088) );
  NAND U39725 ( .A(n59869), .B(n20088), .Z(n20089) );
  AND U39726 ( .A(n22703), .B(n20089), .Z(n20090) );
  NANDN U39727 ( .A(x[7047]), .B(y[7047]), .Z(n59870) );
  AND U39728 ( .A(n20090), .B(n59870), .Z(n20092) );
  NANDN U39729 ( .A(y[7048]), .B(x[7048]), .Z(n20091) );
  NANDN U39730 ( .A(y[7049]), .B(x[7049]), .Z(n22700) );
  AND U39731 ( .A(n20091), .B(n22700), .Z(n50871) );
  NANDN U39732 ( .A(n20092), .B(n50871), .Z(n20093) );
  NAND U39733 ( .A(n20094), .B(n20093), .Z(n20095) );
  NAND U39734 ( .A(n59874), .B(n20095), .Z(n20096) );
  AND U39735 ( .A(n47696), .B(n20096), .Z(n20097) );
  NANDN U39736 ( .A(x[7051]), .B(y[7051]), .Z(n59875) );
  NAND U39737 ( .A(n20097), .B(n59875), .Z(n20099) );
  NANDN U39738 ( .A(y[7052]), .B(x[7052]), .Z(n20098) );
  NANDN U39739 ( .A(y[7053]), .B(x[7053]), .Z(n22698) );
  AND U39740 ( .A(n20098), .B(n22698), .Z(n50869) );
  AND U39741 ( .A(n20099), .B(n50869), .Z(n20101) );
  XNOR U39742 ( .A(x[7054]), .B(y[7054]), .Z(n22699) );
  ANDN U39743 ( .B(y[7053]), .A(x[7053]), .Z(n59877) );
  ANDN U39744 ( .B(n22699), .A(n59877), .Z(n20100) );
  NANDN U39745 ( .A(n20101), .B(n20100), .Z(n20102) );
  NAND U39746 ( .A(n59879), .B(n20102), .Z(n20103) );
  AND U39747 ( .A(n22697), .B(n20103), .Z(n20104) );
  NANDN U39748 ( .A(x[7055]), .B(y[7055]), .Z(n59880) );
  NAND U39749 ( .A(n20104), .B(n59880), .Z(n20105) );
  NAND U39750 ( .A(n59882), .B(n20105), .Z(n20106) );
  AND U39751 ( .A(n59883), .B(n20106), .Z(n20108) );
  NANDN U39752 ( .A(y[7058]), .B(x[7058]), .Z(n20107) );
  NANDN U39753 ( .A(y[7059]), .B(x[7059]), .Z(n22691) );
  AND U39754 ( .A(n20107), .B(n22691), .Z(n59884) );
  NANDN U39755 ( .A(n20108), .B(n59884), .Z(n20109) );
  NAND U39756 ( .A(n20110), .B(n20109), .Z(n20112) );
  NANDN U39757 ( .A(y[7060]), .B(x[7060]), .Z(n20111) );
  NANDN U39758 ( .A(y[7061]), .B(x[7061]), .Z(n22689) );
  AND U39759 ( .A(n20111), .B(n22689), .Z(n59887) );
  AND U39760 ( .A(n20112), .B(n59887), .Z(n20113) );
  ANDN U39761 ( .B(n22690), .A(n20113), .Z(n20114) );
  NANDN U39762 ( .A(x[7061]), .B(y[7061]), .Z(n50867) );
  AND U39763 ( .A(n20114), .B(n50867), .Z(n20115) );
  OR U39764 ( .A(n59888), .B(n20115), .Z(n20116) );
  NAND U39765 ( .A(n20117), .B(n20116), .Z(n20118) );
  NAND U39766 ( .A(n59892), .B(n20118), .Z(n20119) );
  AND U39767 ( .A(n22688), .B(n20119), .Z(n20120) );
  NANDN U39768 ( .A(n59893), .B(n20120), .Z(n20121) );
  NAND U39769 ( .A(n59895), .B(n20121), .Z(n20122) );
  AND U39770 ( .A(n47733), .B(n20122), .Z(n20123) );
  NANDN U39771 ( .A(x[7067]), .B(y[7067]), .Z(n59896) );
  NAND U39772 ( .A(n20123), .B(n59896), .Z(n20124) );
  NAND U39773 ( .A(n59898), .B(n20124), .Z(n20125) );
  AND U39774 ( .A(n22686), .B(n20125), .Z(n20126) );
  NANDN U39775 ( .A(n59899), .B(n20126), .Z(n20127) );
  AND U39776 ( .A(n59901), .B(n20127), .Z(n20128) );
  OR U39777 ( .A(n20129), .B(n20128), .Z(n20130) );
  NAND U39778 ( .A(n59902), .B(n20130), .Z(n20131) );
  NANDN U39779 ( .A(n20132), .B(n20131), .Z(n20133) );
  NAND U39780 ( .A(n59905), .B(n20133), .Z(n20134) );
  AND U39781 ( .A(n47753), .B(n20134), .Z(n20135) );
  NANDN U39782 ( .A(x[7075]), .B(y[7075]), .Z(n50864) );
  AND U39783 ( .A(n20135), .B(n50864), .Z(n20136) );
  OR U39784 ( .A(n59907), .B(n20136), .Z(n20137) );
  NAND U39785 ( .A(n20138), .B(n20137), .Z(n20139) );
  NAND U39786 ( .A(n59910), .B(n20139), .Z(n20140) );
  AND U39787 ( .A(n22680), .B(n20140), .Z(n20141) );
  NANDN U39788 ( .A(x[7079]), .B(y[7079]), .Z(n59911) );
  NAND U39789 ( .A(n20141), .B(n59911), .Z(n20143) );
  NANDN U39790 ( .A(y[7080]), .B(x[7080]), .Z(n20142) );
  NANDN U39791 ( .A(y[7081]), .B(x[7081]), .Z(n22677) );
  AND U39792 ( .A(n20142), .B(n22677), .Z(n50862) );
  AND U39793 ( .A(n20143), .B(n50862), .Z(n20145) );
  XNOR U39794 ( .A(x[7082]), .B(y[7082]), .Z(n22678) );
  NANDN U39795 ( .A(x[7081]), .B(y[7081]), .Z(n59913) );
  AND U39796 ( .A(n22678), .B(n59913), .Z(n20144) );
  NANDN U39797 ( .A(n20145), .B(n20144), .Z(n20146) );
  NANDN U39798 ( .A(n59915), .B(n20146), .Z(n20147) );
  AND U39799 ( .A(n47771), .B(n20147), .Z(n20148) );
  NANDN U39800 ( .A(x[7083]), .B(y[7083]), .Z(n50861) );
  NAND U39801 ( .A(n20148), .B(n50861), .Z(n20149) );
  AND U39802 ( .A(n59916), .B(n20149), .Z(n20150) );
  OR U39803 ( .A(n20151), .B(n20150), .Z(n20152) );
  NAND U39804 ( .A(n50859), .B(n20152), .Z(n20153) );
  NANDN U39805 ( .A(n20154), .B(n20153), .Z(n20155) );
  NAND U39806 ( .A(n59922), .B(n20155), .Z(n20156) );
  AND U39807 ( .A(n22674), .B(n20156), .Z(n20157) );
  ANDN U39808 ( .B(y[7089]), .A(x[7089]), .Z(n59923) );
  ANDN U39809 ( .B(n20157), .A(n59923), .Z(n20159) );
  NANDN U39810 ( .A(y[7090]), .B(x[7090]), .Z(n20158) );
  NANDN U39811 ( .A(y[7091]), .B(x[7091]), .Z(n22671) );
  NAND U39812 ( .A(n20158), .B(n22671), .Z(n50858) );
  OR U39813 ( .A(n20159), .B(n50858), .Z(n20160) );
  NAND U39814 ( .A(n20161), .B(n20160), .Z(n20162) );
  NAND U39815 ( .A(n59927), .B(n20162), .Z(n20163) );
  NAND U39816 ( .A(n59928), .B(n20163), .Z(n20164) );
  NAND U39817 ( .A(n59929), .B(n20164), .Z(n20165) );
  AND U39818 ( .A(n47799), .B(n20165), .Z(n20166) );
  NANDN U39819 ( .A(x[7095]), .B(y[7095]), .Z(n50857) );
  AND U39820 ( .A(n20166), .B(n50857), .Z(n20168) );
  NANDN U39821 ( .A(y[7096]), .B(x[7096]), .Z(n20167) );
  NANDN U39822 ( .A(y[7097]), .B(x[7097]), .Z(n22665) );
  AND U39823 ( .A(n20167), .B(n22665), .Z(n59930) );
  NANDN U39824 ( .A(n20168), .B(n59930), .Z(n20169) );
  AND U39825 ( .A(n22666), .B(n20169), .Z(n20170) );
  NANDN U39826 ( .A(n59931), .B(n20170), .Z(n20172) );
  NANDN U39827 ( .A(y[7098]), .B(x[7098]), .Z(n20171) );
  NANDN U39828 ( .A(y[7099]), .B(x[7099]), .Z(n47808) );
  AND U39829 ( .A(n20171), .B(n47808), .Z(n59933) );
  AND U39830 ( .A(n20172), .B(n59933), .Z(n20173) );
  OR U39831 ( .A(n20174), .B(n20173), .Z(n20175) );
  NAND U39832 ( .A(n50852), .B(n20175), .Z(n20176) );
  NANDN U39833 ( .A(n20177), .B(n20176), .Z(n20178) );
  NAND U39834 ( .A(n59938), .B(n20178), .Z(n20179) );
  AND U39835 ( .A(n47819), .B(n20179), .Z(n20180) );
  NANDN U39836 ( .A(x[7103]), .B(y[7103]), .Z(n59939) );
  AND U39837 ( .A(n20180), .B(n59939), .Z(n20181) );
  OR U39838 ( .A(n59940), .B(n20181), .Z(n20182) );
  NAND U39839 ( .A(n20183), .B(n20182), .Z(n20184) );
  NAND U39840 ( .A(n59943), .B(n20184), .Z(n20185) );
  AND U39841 ( .A(n47829), .B(n20185), .Z(n20186) );
  NANDN U39842 ( .A(x[7107]), .B(y[7107]), .Z(n59944) );
  NAND U39843 ( .A(n20186), .B(n59944), .Z(n20187) );
  AND U39844 ( .A(n59946), .B(n20187), .Z(n20189) );
  XNOR U39845 ( .A(x[7110]), .B(y[7110]), .Z(n22659) );
  NANDN U39846 ( .A(x[7109]), .B(y[7109]), .Z(n22660) );
  AND U39847 ( .A(n22659), .B(n22660), .Z(n20188) );
  NANDN U39848 ( .A(n20189), .B(n20188), .Z(n20190) );
  NANDN U39849 ( .A(n50848), .B(n20190), .Z(n20191) );
  AND U39850 ( .A(n47839), .B(n20191), .Z(n20192) );
  NANDN U39851 ( .A(x[7111]), .B(y[7111]), .Z(n59949) );
  NAND U39852 ( .A(n20192), .B(n59949), .Z(n20193) );
  AND U39853 ( .A(n59951), .B(n20193), .Z(n20194) );
  OR U39854 ( .A(n20195), .B(n20194), .Z(n20196) );
  NAND U39855 ( .A(n50847), .B(n20196), .Z(n20197) );
  NANDN U39856 ( .A(n20198), .B(n20197), .Z(n20199) );
  NAND U39857 ( .A(n59956), .B(n20199), .Z(n20200) );
  AND U39858 ( .A(n22655), .B(n20200), .Z(n20201) );
  ANDN U39859 ( .B(y[7117]), .A(x[7117]), .Z(n59957) );
  ANDN U39860 ( .B(n20201), .A(n59957), .Z(n20202) );
  OR U39861 ( .A(n59959), .B(n20202), .Z(n20203) );
  NAND U39862 ( .A(n20204), .B(n20203), .Z(n20205) );
  NAND U39863 ( .A(n59962), .B(n20205), .Z(n20206) );
  AND U39864 ( .A(n22653), .B(n20206), .Z(n20207) );
  NANDN U39865 ( .A(n59963), .B(n20207), .Z(n20208) );
  AND U39866 ( .A(n59965), .B(n20208), .Z(n20210) );
  XNOR U39867 ( .A(x[7124]), .B(y[7124]), .Z(n22651) );
  NANDN U39868 ( .A(x[7123]), .B(y[7123]), .Z(n50844) );
  AND U39869 ( .A(n22651), .B(n50844), .Z(n20209) );
  NANDN U39870 ( .A(n20210), .B(n20209), .Z(n20211) );
  NAND U39871 ( .A(n59967), .B(n20211), .Z(n20212) );
  AND U39872 ( .A(n22649), .B(n20212), .Z(n20213) );
  NANDN U39873 ( .A(n59968), .B(n20213), .Z(n20214) );
  NAND U39874 ( .A(n59970), .B(n20214), .Z(n20215) );
  AND U39875 ( .A(n47878), .B(n20215), .Z(n20216) );
  NANDN U39876 ( .A(n47874), .B(n20216), .Z(n20217) );
  NAND U39877 ( .A(n50843), .B(n20217), .Z(n20218) );
  NAND U39878 ( .A(n22647), .B(n20218), .Z(n20219) );
  ANDN U39879 ( .B(y[7129]), .A(x[7129]), .Z(n59973) );
  OR U39880 ( .A(n20219), .B(n59973), .Z(n20220) );
  NAND U39881 ( .A(n59975), .B(n20220), .Z(n20221) );
  AND U39882 ( .A(n47888), .B(n20221), .Z(n20222) );
  NANDN U39883 ( .A(x[7131]), .B(y[7131]), .Z(n59976) );
  AND U39884 ( .A(n20222), .B(n59976), .Z(n20224) );
  NANDN U39885 ( .A(y[7132]), .B(x[7132]), .Z(n20223) );
  NANDN U39886 ( .A(y[7133]), .B(x[7133]), .Z(n22644) );
  NAND U39887 ( .A(n20223), .B(n22644), .Z(n59977) );
  OR U39888 ( .A(n20224), .B(n59977), .Z(n20225) );
  NANDN U39889 ( .A(x[7135]), .B(y[7135]), .Z(n59982) );
  NANDN U39890 ( .A(y[7136]), .B(x[7136]), .Z(n20227) );
  NANDN U39891 ( .A(y[7137]), .B(x[7137]), .Z(n22641) );
  NAND U39892 ( .A(n20227), .B(n22641), .Z(n50841) );
  NANDN U39893 ( .A(x[7139]), .B(y[7139]), .Z(n59987) );
  ANDN U39894 ( .B(y[7141]), .A(x[7141]), .Z(n50839) );
  NANDN U39895 ( .A(x[7145]), .B(y[7145]), .Z(n50837) );
  NANDN U39896 ( .A(y[7146]), .B(x[7146]), .Z(n20228) );
  NANDN U39897 ( .A(y[7147]), .B(x[7147]), .Z(n47925) );
  NAND U39898 ( .A(n20228), .B(n47925), .Z(n50836) );
  OR U39899 ( .A(n20229), .B(n50836), .Z(n20230) );
  AND U39900 ( .A(n47926), .B(n20230), .Z(n20231) );
  NANDN U39901 ( .A(x[7147]), .B(y[7147]), .Z(n50835) );
  NAND U39902 ( .A(n20231), .B(n50835), .Z(n20232) );
  AND U39903 ( .A(n59994), .B(n20232), .Z(n20233) );
  OR U39904 ( .A(n20234), .B(n20233), .Z(n20235) );
  NAND U39905 ( .A(n59997), .B(n20235), .Z(n20236) );
  NANDN U39906 ( .A(n20237), .B(n20236), .Z(n20238) );
  NAND U39907 ( .A(n59998), .B(n20238), .Z(n20239) );
  AND U39908 ( .A(n22630), .B(n20239), .Z(n20240) );
  ANDN U39909 ( .B(y[7153]), .A(x[7153]), .Z(n59999) );
  ANDN U39910 ( .B(n20240), .A(n59999), .Z(n20242) );
  NANDN U39911 ( .A(y[7154]), .B(x[7154]), .Z(n20241) );
  NANDN U39912 ( .A(y[7155]), .B(x[7155]), .Z(n22627) );
  NAND U39913 ( .A(n20241), .B(n22627), .Z(n60001) );
  OR U39914 ( .A(n20242), .B(n60001), .Z(n20243) );
  NAND U39915 ( .A(n20244), .B(n20243), .Z(n20245) );
  NANDN U39916 ( .A(n50829), .B(n20245), .Z(n20246) );
  AND U39917 ( .A(n22626), .B(n20246), .Z(n20247) );
  NANDN U39918 ( .A(x[7157]), .B(y[7157]), .Z(n50827) );
  NAND U39919 ( .A(n20247), .B(n50827), .Z(n20248) );
  AND U39920 ( .A(n60003), .B(n20248), .Z(n20249) );
  XNOR U39921 ( .A(y[7160]), .B(x[7160]), .Z(n47955) );
  NANDN U39922 ( .A(x[7159]), .B(y[7159]), .Z(n47951) );
  AND U39923 ( .A(n47955), .B(n47951), .Z(n60004) );
  NANDN U39924 ( .A(n20249), .B(n60004), .Z(n20250) );
  NAND U39925 ( .A(n60005), .B(n20250), .Z(n20251) );
  AND U39926 ( .A(n22623), .B(n20251), .Z(n20252) );
  NANDN U39927 ( .A(x[7161]), .B(y[7161]), .Z(n60007) );
  NAND U39928 ( .A(n20252), .B(n60007), .Z(n20254) );
  NANDN U39929 ( .A(y[7162]), .B(x[7162]), .Z(n20253) );
  NANDN U39930 ( .A(y[7163]), .B(x[7163]), .Z(n47964) );
  AND U39931 ( .A(n20253), .B(n47964), .Z(n50826) );
  AND U39932 ( .A(n20254), .B(n50826), .Z(n20255) );
  ANDN U39933 ( .B(n47965), .A(n20255), .Z(n20256) );
  NANDN U39934 ( .A(x[7163]), .B(y[7163]), .Z(n60008) );
  AND U39935 ( .A(n20256), .B(n60008), .Z(n20258) );
  NANDN U39936 ( .A(y[7164]), .B(x[7164]), .Z(n20257) );
  NANDN U39937 ( .A(y[7165]), .B(x[7165]), .Z(n22620) );
  AND U39938 ( .A(n20257), .B(n22620), .Z(n60010) );
  NANDN U39939 ( .A(n20258), .B(n60010), .Z(n20259) );
  NAND U39940 ( .A(n20260), .B(n20259), .Z(n20261) );
  NAND U39941 ( .A(n60013), .B(n20261), .Z(n20262) );
  AND U39942 ( .A(n47975), .B(n20262), .Z(n20263) );
  NANDN U39943 ( .A(x[7167]), .B(y[7167]), .Z(n60014) );
  AND U39944 ( .A(n20263), .B(n60014), .Z(n20265) );
  NANDN U39945 ( .A(y[7168]), .B(x[7168]), .Z(n20264) );
  NANDN U39946 ( .A(y[7169]), .B(x[7169]), .Z(n22618) );
  AND U39947 ( .A(n20264), .B(n22618), .Z(n60017) );
  NANDN U39948 ( .A(n20265), .B(n60017), .Z(n20266) );
  NAND U39949 ( .A(n20267), .B(n20266), .Z(n20268) );
  NAND U39950 ( .A(n60020), .B(n20268), .Z(n20269) );
  AND U39951 ( .A(n47986), .B(n20269), .Z(n20270) );
  NANDN U39952 ( .A(n50825), .B(n20270), .Z(n20271) );
  AND U39953 ( .A(n60021), .B(n20271), .Z(n20272) );
  NOR U39954 ( .A(n60022), .B(n20272), .Z(n20273) );
  NAND U39955 ( .A(n22617), .B(n20273), .Z(n20274) );
  NANDN U39956 ( .A(n60024), .B(n20274), .Z(n20275) );
  XOR U39957 ( .A(x[7176]), .B(y[7176]), .Z(n47996) );
  ANDN U39958 ( .B(n20275), .A(n47996), .Z(n20276) );
  NANDN U39959 ( .A(x[7175]), .B(y[7175]), .Z(n50822) );
  NAND U39960 ( .A(n20276), .B(n50822), .Z(n20278) );
  NANDN U39961 ( .A(y[7176]), .B(x[7176]), .Z(n20277) );
  NANDN U39962 ( .A(y[7177]), .B(x[7177]), .Z(n22614) );
  AND U39963 ( .A(n20277), .B(n22614), .Z(n50821) );
  AND U39964 ( .A(n20278), .B(n50821), .Z(n20280) );
  XNOR U39965 ( .A(x[7178]), .B(y[7178]), .Z(n22615) );
  NANDN U39966 ( .A(x[7177]), .B(y[7177]), .Z(n60025) );
  AND U39967 ( .A(n22615), .B(n60025), .Z(n20279) );
  NANDN U39968 ( .A(n20280), .B(n20279), .Z(n20281) );
  NAND U39969 ( .A(n60027), .B(n20281), .Z(n20282) );
  AND U39970 ( .A(n22613), .B(n20282), .Z(n20283) );
  NANDN U39971 ( .A(x[7179]), .B(y[7179]), .Z(n60028) );
  NAND U39972 ( .A(n20283), .B(n60028), .Z(n20285) );
  NANDN U39973 ( .A(y[7180]), .B(x[7180]), .Z(n20284) );
  NANDN U39974 ( .A(y[7181]), .B(x[7181]), .Z(n22610) );
  AND U39975 ( .A(n20284), .B(n22610), .Z(n50820) );
  AND U39976 ( .A(n20285), .B(n50820), .Z(n20286) );
  OR U39977 ( .A(n20287), .B(n20286), .Z(n20288) );
  NAND U39978 ( .A(n60034), .B(n20288), .Z(n20289) );
  NANDN U39979 ( .A(n20290), .B(n20289), .Z(n20291) );
  NAND U39980 ( .A(n60037), .B(n20291), .Z(n20292) );
  AND U39981 ( .A(n22608), .B(n20292), .Z(n20293) );
  NANDN U39982 ( .A(x[7185]), .B(y[7185]), .Z(n22609) );
  AND U39983 ( .A(n20293), .B(n22609), .Z(n20295) );
  NANDN U39984 ( .A(y[7186]), .B(x[7186]), .Z(n20294) );
  NANDN U39985 ( .A(y[7187]), .B(x[7187]), .Z(n48023) );
  AND U39986 ( .A(n20294), .B(n48023), .Z(n60038) );
  NANDN U39987 ( .A(n20295), .B(n60038), .Z(n20296) );
  NAND U39988 ( .A(n20297), .B(n20296), .Z(n20298) );
  NANDN U39989 ( .A(n60041), .B(n20298), .Z(n20299) );
  NAND U39990 ( .A(n60042), .B(n20299), .Z(n20300) );
  NAND U39991 ( .A(n60043), .B(n20300), .Z(n20301) );
  AND U39992 ( .A(n60044), .B(n20301), .Z(n20302) );
  NANDN U39993 ( .A(y[7192]), .B(x[7192]), .Z(n22600) );
  NANDN U39994 ( .A(y[7193]), .B(x[7193]), .Z(n22598) );
  AND U39995 ( .A(n22600), .B(n22598), .Z(n60045) );
  NANDN U39996 ( .A(n20302), .B(n60045), .Z(n20303) );
  NAND U39997 ( .A(n20304), .B(n20303), .Z(n20305) );
  AND U39998 ( .A(n60049), .B(n20305), .Z(n20307) );
  XNOR U39999 ( .A(x[7196]), .B(y[7196]), .Z(n48043) );
  NANDN U40000 ( .A(x[7195]), .B(y[7195]), .Z(n50816) );
  AND U40001 ( .A(n48043), .B(n50816), .Z(n20306) );
  NANDN U40002 ( .A(n20307), .B(n20306), .Z(n20308) );
  NAND U40003 ( .A(n60050), .B(n20308), .Z(n20309) );
  ANDN U40004 ( .B(y[7197]), .A(x[7197]), .Z(n60051) );
  ANDN U40005 ( .B(n20309), .A(n60051), .Z(n20310) );
  NAND U40006 ( .A(n22597), .B(n20310), .Z(n20311) );
  NANDN U40007 ( .A(n60053), .B(n20311), .Z(n20312) );
  AND U40008 ( .A(n48053), .B(n20312), .Z(n20313) );
  NANDN U40009 ( .A(x[7199]), .B(y[7199]), .Z(n50815) );
  NAND U40010 ( .A(n20313), .B(n50815), .Z(n20315) );
  NANDN U40011 ( .A(y[7200]), .B(x[7200]), .Z(n20314) );
  NANDN U40012 ( .A(y[7201]), .B(x[7201]), .Z(n22594) );
  AND U40013 ( .A(n20314), .B(n22594), .Z(n50813) );
  AND U40014 ( .A(n20315), .B(n50813), .Z(n20316) );
  NANDN U40015 ( .A(x[7202]), .B(y[7202]), .Z(n22592) );
  ANDN U40016 ( .B(y[7201]), .A(x[7201]), .Z(n22595) );
  ANDN U40017 ( .B(n22592), .A(n22595), .Z(n60054) );
  NANDN U40018 ( .A(n20316), .B(n60054), .Z(n20317) );
  NAND U40019 ( .A(n60055), .B(n20317), .Z(n20318) );
  NAND U40020 ( .A(n22590), .B(n20318), .Z(n20319) );
  ANDN U40021 ( .B(y[7203]), .A(x[7203]), .Z(n22591) );
  OR U40022 ( .A(n20319), .B(n22591), .Z(n20320) );
  NAND U40023 ( .A(n60057), .B(n20320), .Z(n20321) );
  NAND U40024 ( .A(n60059), .B(n20321), .Z(n20322) );
  AND U40025 ( .A(n60060), .B(n20322), .Z(n20323) );
  NANDN U40026 ( .A(x[7207]), .B(y[7207]), .Z(n22585) );
  ANDN U40027 ( .B(y[7208]), .A(x[7208]), .Z(n48074) );
  ANDN U40028 ( .B(n22585), .A(n48074), .Z(n60061) );
  NANDN U40029 ( .A(n20323), .B(n60061), .Z(n20324) );
  NAND U40030 ( .A(n60062), .B(n20324), .Z(n20325) );
  NAND U40031 ( .A(n60064), .B(n20325), .Z(n20326) );
  XNOR U40032 ( .A(x[7210]), .B(y[7210]), .Z(n22582) );
  NANDN U40033 ( .A(n20326), .B(n22582), .Z(n20327) );
  NAND U40034 ( .A(n60065), .B(n20327), .Z(n20328) );
  AND U40035 ( .A(n48081), .B(n20328), .Z(n20329) );
  NANDN U40036 ( .A(x[7211]), .B(y[7211]), .Z(n60066) );
  AND U40037 ( .A(n20329), .B(n60066), .Z(n20331) );
  NANDN U40038 ( .A(y[7212]), .B(x[7212]), .Z(n20330) );
  NANDN U40039 ( .A(y[7213]), .B(x[7213]), .Z(n22579) );
  AND U40040 ( .A(n20330), .B(n22579), .Z(n60068) );
  NANDN U40041 ( .A(n20331), .B(n60068), .Z(n20332) );
  NAND U40042 ( .A(n20333), .B(n20332), .Z(n20334) );
  NAND U40043 ( .A(n50811), .B(n20334), .Z(n20335) );
  AND U40044 ( .A(n48091), .B(n20335), .Z(n20336) );
  NANDN U40045 ( .A(x[7215]), .B(y[7215]), .Z(n60071) );
  NAND U40046 ( .A(n20336), .B(n60071), .Z(n20337) );
  AND U40047 ( .A(n60073), .B(n20337), .Z(n20338) );
  NOR U40048 ( .A(n60074), .B(n20338), .Z(n20339) );
  NAND U40049 ( .A(n22578), .B(n20339), .Z(n20340) );
  NANDN U40050 ( .A(n60077), .B(n20340), .Z(n20341) );
  AND U40051 ( .A(n48102), .B(n20341), .Z(n20342) );
  NANDN U40052 ( .A(n50810), .B(n20342), .Z(n20343) );
  AND U40053 ( .A(n60078), .B(n20343), .Z(n20345) );
  XNOR U40054 ( .A(x[7222]), .B(y[7222]), .Z(n22576) );
  ANDN U40055 ( .B(y[7221]), .A(x[7221]), .Z(n60079) );
  ANDN U40056 ( .B(n22576), .A(n60079), .Z(n20344) );
  NANDN U40057 ( .A(n20345), .B(n20344), .Z(n20346) );
  NANDN U40058 ( .A(n60081), .B(n20346), .Z(n20347) );
  AND U40059 ( .A(n48112), .B(n20347), .Z(n20348) );
  NANDN U40060 ( .A(x[7223]), .B(y[7223]), .Z(n50808) );
  NAND U40061 ( .A(n20348), .B(n50808), .Z(n20350) );
  NANDN U40062 ( .A(y[7224]), .B(x[7224]), .Z(n20349) );
  NANDN U40063 ( .A(y[7225]), .B(x[7225]), .Z(n22573) );
  AND U40064 ( .A(n20349), .B(n22573), .Z(n50806) );
  AND U40065 ( .A(n20350), .B(n50806), .Z(n20351) );
  OR U40066 ( .A(n20352), .B(n20351), .Z(n20353) );
  NAND U40067 ( .A(n60084), .B(n20353), .Z(n20354) );
  NANDN U40068 ( .A(n20355), .B(n20354), .Z(n20357) );
  NANDN U40069 ( .A(y[7228]), .B(x[7228]), .Z(n20356) );
  NANDN U40070 ( .A(y[7229]), .B(x[7229]), .Z(n22571) );
  AND U40071 ( .A(n20356), .B(n22571), .Z(n50804) );
  AND U40072 ( .A(n20357), .B(n50804), .Z(n20359) );
  XNOR U40073 ( .A(x[7230]), .B(y[7230]), .Z(n22572) );
  ANDN U40074 ( .B(y[7229]), .A(x[7229]), .Z(n60087) );
  ANDN U40075 ( .B(n22572), .A(n60087), .Z(n20358) );
  NANDN U40076 ( .A(n20359), .B(n20358), .Z(n20360) );
  NAND U40077 ( .A(n60089), .B(n20360), .Z(n20361) );
  AND U40078 ( .A(n20362), .B(n20361), .Z(n20364) );
  NANDN U40079 ( .A(y[7232]), .B(x[7232]), .Z(n20363) );
  NANDN U40080 ( .A(y[7233]), .B(x[7233]), .Z(n22568) );
  NAND U40081 ( .A(n20363), .B(n22568), .Z(n60092) );
  OR U40082 ( .A(n20364), .B(n60092), .Z(n20365) );
  AND U40083 ( .A(n22569), .B(n20365), .Z(n20366) );
  NANDN U40084 ( .A(n50802), .B(n20366), .Z(n20367) );
  AND U40085 ( .A(n60093), .B(n20367), .Z(n20368) );
  OR U40086 ( .A(n20369), .B(n20368), .Z(n20370) );
  NAND U40087 ( .A(n60096), .B(n20370), .Z(n20371) );
  NANDN U40088 ( .A(n20372), .B(n20371), .Z(n20373) );
  NAND U40089 ( .A(n60097), .B(n20373), .Z(n20374) );
  AND U40090 ( .A(n48150), .B(n20374), .Z(n20375) );
  NANDN U40091 ( .A(x[7239]), .B(y[7239]), .Z(n60098) );
  AND U40092 ( .A(n20375), .B(n60098), .Z(n20377) );
  NANDN U40093 ( .A(y[7240]), .B(x[7240]), .Z(n20376) );
  NANDN U40094 ( .A(y[7241]), .B(x[7241]), .Z(n22562) );
  AND U40095 ( .A(n20376), .B(n22562), .Z(n60101) );
  NANDN U40096 ( .A(n20377), .B(n60101), .Z(n20378) );
  NAND U40097 ( .A(n20379), .B(n20378), .Z(n20380) );
  NANDN U40098 ( .A(n60104), .B(n20380), .Z(n20381) );
  AND U40099 ( .A(n22561), .B(n20381), .Z(n20382) );
  NANDN U40100 ( .A(x[7243]), .B(y[7243]), .Z(n60105) );
  NAND U40101 ( .A(n20382), .B(n60105), .Z(n20383) );
  AND U40102 ( .A(n60107), .B(n20383), .Z(n20384) );
  XNOR U40103 ( .A(y[7246]), .B(x[7246]), .Z(n22558) );
  NANDN U40104 ( .A(x[7245]), .B(y[7245]), .Z(n22559) );
  NAND U40105 ( .A(n22558), .B(n22559), .Z(n60108) );
  OR U40106 ( .A(n20384), .B(n60108), .Z(n20385) );
  NAND U40107 ( .A(n60109), .B(n20385), .Z(n20386) );
  AND U40108 ( .A(n48169), .B(n20386), .Z(n20387) );
  NANDN U40109 ( .A(x[7247]), .B(y[7247]), .Z(n50799) );
  NAND U40110 ( .A(n20387), .B(n50799), .Z(n20388) );
  NAND U40111 ( .A(n60110), .B(n20388), .Z(n20389) );
  AND U40112 ( .A(n22556), .B(n20389), .Z(n20390) );
  ANDN U40113 ( .B(y[7249]), .A(x[7249]), .Z(n60111) );
  ANDN U40114 ( .B(n20390), .A(n60111), .Z(n20392) );
  NANDN U40115 ( .A(y[7250]), .B(x[7250]), .Z(n20391) );
  NANDN U40116 ( .A(y[7251]), .B(x[7251]), .Z(n48179) );
  AND U40117 ( .A(n20391), .B(n48179), .Z(n50797) );
  NANDN U40118 ( .A(n20392), .B(n50797), .Z(n20393) );
  NAND U40119 ( .A(n20394), .B(n20393), .Z(n20395) );
  NAND U40120 ( .A(n60115), .B(n20395), .Z(n20396) );
  AND U40121 ( .A(n22554), .B(n20396), .Z(n20397) );
  ANDN U40122 ( .B(y[7253]), .A(x[7253]), .Z(n60116) );
  ANDN U40123 ( .B(n20397), .A(n60116), .Z(n20399) );
  NANDN U40124 ( .A(y[7254]), .B(x[7254]), .Z(n20398) );
  NANDN U40125 ( .A(y[7255]), .B(x[7255]), .Z(n48189) );
  NAND U40126 ( .A(n20398), .B(n48189), .Z(n60118) );
  OR U40127 ( .A(n20399), .B(n60118), .Z(n20400) );
  NAND U40128 ( .A(n20401), .B(n20400), .Z(n20402) );
  NAND U40129 ( .A(n60121), .B(n20402), .Z(n20403) );
  AND U40130 ( .A(n22552), .B(n20403), .Z(n20404) );
  ANDN U40131 ( .B(y[7257]), .A(x[7257]), .Z(n60122) );
  ANDN U40132 ( .B(n20404), .A(n60122), .Z(n20406) );
  NANDN U40133 ( .A(y[7258]), .B(x[7258]), .Z(n20405) );
  NANDN U40134 ( .A(y[7259]), .B(x[7259]), .Z(n48199) );
  AND U40135 ( .A(n20405), .B(n48199), .Z(n60124) );
  NANDN U40136 ( .A(n20406), .B(n60124), .Z(n20407) );
  NAND U40137 ( .A(n20408), .B(n20407), .Z(n20409) );
  NANDN U40138 ( .A(n60127), .B(n20409), .Z(n20410) );
  NAND U40139 ( .A(n60128), .B(n20410), .Z(n20411) );
  NAND U40140 ( .A(n60129), .B(n20411), .Z(n20412) );
  AND U40141 ( .A(n22547), .B(n20412), .Z(n20413) );
  NANDN U40142 ( .A(x[7263]), .B(y[7263]), .Z(n60130) );
  NAND U40143 ( .A(n20413), .B(n60130), .Z(n20414) );
  NANDN U40144 ( .A(n60133), .B(n20414), .Z(n20415) );
  AND U40145 ( .A(n22545), .B(n20415), .Z(n20416) );
  NANDN U40146 ( .A(n50794), .B(n20416), .Z(n20417) );
  NAND U40147 ( .A(n60135), .B(n20417), .Z(n20418) );
  AND U40148 ( .A(n48219), .B(n20418), .Z(n20419) );
  NANDN U40149 ( .A(x[7267]), .B(y[7267]), .Z(n50791) );
  AND U40150 ( .A(n20419), .B(n50791), .Z(n20421) );
  NANDN U40151 ( .A(y[7268]), .B(x[7268]), .Z(n20420) );
  NANDN U40152 ( .A(y[7269]), .B(x[7269]), .Z(n22542) );
  AND U40153 ( .A(n20420), .B(n22542), .Z(n60136) );
  NANDN U40154 ( .A(n20421), .B(n60136), .Z(n20422) );
  NAND U40155 ( .A(n20423), .B(n20422), .Z(n20424) );
  NAND U40156 ( .A(n60139), .B(n20424), .Z(n20425) );
  AND U40157 ( .A(n48229), .B(n20425), .Z(n20426) );
  NANDN U40158 ( .A(x[7271]), .B(y[7271]), .Z(n50790) );
  AND U40159 ( .A(n20426), .B(n50790), .Z(n20428) );
  NANDN U40160 ( .A(y[7272]), .B(x[7272]), .Z(n20427) );
  NANDN U40161 ( .A(y[7273]), .B(x[7273]), .Z(n22540) );
  NAND U40162 ( .A(n20427), .B(n22540), .Z(n60140) );
  OR U40163 ( .A(n20428), .B(n60140), .Z(n20429) );
  NAND U40164 ( .A(n20430), .B(n20429), .Z(n20431) );
  AND U40165 ( .A(n60143), .B(n20431), .Z(n20433) );
  XNOR U40166 ( .A(x[7276]), .B(y[7276]), .Z(n48239) );
  NANDN U40167 ( .A(x[7275]), .B(y[7275]), .Z(n60144) );
  AND U40168 ( .A(n48239), .B(n60144), .Z(n20432) );
  NANDN U40169 ( .A(n20433), .B(n20432), .Z(n20434) );
  NANDN U40170 ( .A(n60146), .B(n20434), .Z(n20435) );
  AND U40171 ( .A(n22539), .B(n20435), .Z(n20436) );
  NANDN U40172 ( .A(n60147), .B(n20436), .Z(n20437) );
  NAND U40173 ( .A(n60149), .B(n20437), .Z(n20438) );
  AND U40174 ( .A(n48249), .B(n20438), .Z(n20439) );
  NANDN U40175 ( .A(x[7279]), .B(y[7279]), .Z(n60150) );
  NAND U40176 ( .A(n20439), .B(n60150), .Z(n20440) );
  NAND U40177 ( .A(n60152), .B(n20440), .Z(n20441) );
  AND U40178 ( .A(n22536), .B(n20441), .Z(n20442) );
  NANDN U40179 ( .A(x[7281]), .B(y[7281]), .Z(n22537) );
  AND U40180 ( .A(n20442), .B(n22537), .Z(n20444) );
  NANDN U40181 ( .A(y[7282]), .B(x[7282]), .Z(n20443) );
  NANDN U40182 ( .A(y[7283]), .B(x[7283]), .Z(n22533) );
  AND U40183 ( .A(n20443), .B(n22533), .Z(n60153) );
  NANDN U40184 ( .A(n20444), .B(n60153), .Z(n20445) );
  NAND U40185 ( .A(n20446), .B(n20445), .Z(n20447) );
  NAND U40186 ( .A(n60156), .B(n20447), .Z(n20448) );
  AND U40187 ( .A(n60157), .B(n20448), .Z(n20449) );
  OR U40188 ( .A(n60158), .B(n20449), .Z(n20450) );
  NAND U40189 ( .A(n60159), .B(n20450), .Z(n20451) );
  NAND U40190 ( .A(n60160), .B(n20451), .Z(n20452) );
  AND U40191 ( .A(n22524), .B(n20452), .Z(n20453) );
  NANDN U40192 ( .A(x[7289]), .B(y[7289]), .Z(n60161) );
  NAND U40193 ( .A(n20453), .B(n60161), .Z(n20454) );
  AND U40194 ( .A(n60164), .B(n20454), .Z(n20455) );
  OR U40195 ( .A(n20456), .B(n20455), .Z(n20457) );
  NAND U40196 ( .A(n60165), .B(n20457), .Z(n20458) );
  NANDN U40197 ( .A(n20459), .B(n20458), .Z(n20460) );
  NAND U40198 ( .A(n60167), .B(n20460), .Z(n20461) );
  NANDN U40199 ( .A(x[7295]), .B(y[7295]), .Z(n22520) );
  NANDN U40200 ( .A(x[7296]), .B(y[7296]), .Z(n22517) );
  AND U40201 ( .A(n22520), .B(n22517), .Z(n50782) );
  AND U40202 ( .A(n20461), .B(n50782), .Z(n20462) );
  NANDN U40203 ( .A(y[7296]), .B(x[7296]), .Z(n22518) );
  NANDN U40204 ( .A(y[7297]), .B(x[7297]), .Z(n22515) );
  AND U40205 ( .A(n22518), .B(n22515), .Z(n60168) );
  NANDN U40206 ( .A(n20462), .B(n60168), .Z(n20463) );
  NAND U40207 ( .A(n60169), .B(n20463), .Z(n20464) );
  NANDN U40208 ( .A(n60170), .B(n20464), .Z(n20465) );
  AND U40209 ( .A(n48294), .B(n20465), .Z(n20466) );
  NANDN U40210 ( .A(x[7299]), .B(y[7299]), .Z(n50781) );
  NAND U40211 ( .A(n20466), .B(n50781), .Z(n20467) );
  AND U40212 ( .A(n60171), .B(n20467), .Z(n20468) );
  OR U40213 ( .A(n20469), .B(n20468), .Z(n20470) );
  NAND U40214 ( .A(n60173), .B(n20470), .Z(n20471) );
  NANDN U40215 ( .A(n20472), .B(n20471), .Z(n20473) );
  NAND U40216 ( .A(n60176), .B(n20473), .Z(n20474) );
  AND U40217 ( .A(n22510), .B(n20474), .Z(n20475) );
  ANDN U40218 ( .B(y[7305]), .A(x[7305]), .Z(n50776) );
  ANDN U40219 ( .B(n20475), .A(n50776), .Z(n20476) );
  OR U40220 ( .A(n60177), .B(n20476), .Z(n20477) );
  NAND U40221 ( .A(n20478), .B(n20477), .Z(n20479) );
  NAND U40222 ( .A(n60180), .B(n20479), .Z(n20480) );
  AND U40223 ( .A(n22508), .B(n20480), .Z(n20481) );
  NANDN U40224 ( .A(x[7309]), .B(y[7309]), .Z(n60181) );
  NAND U40225 ( .A(n20481), .B(n60181), .Z(n20482) );
  AND U40226 ( .A(n60183), .B(n20482), .Z(n20484) );
  NANDN U40227 ( .A(x[7311]), .B(y[7311]), .Z(n60184) );
  XOR U40228 ( .A(x[7312]), .B(y[7312]), .Z(n48324) );
  ANDN U40229 ( .B(n60184), .A(n48324), .Z(n20483) );
  NANDN U40230 ( .A(n20484), .B(n20483), .Z(n20485) );
  NAND U40231 ( .A(n60186), .B(n20485), .Z(n20486) );
  AND U40232 ( .A(n22506), .B(n20486), .Z(n20487) );
  NANDN U40233 ( .A(x[7313]), .B(y[7313]), .Z(n60187) );
  NAND U40234 ( .A(n20487), .B(n60187), .Z(n20488) );
  NAND U40235 ( .A(n60190), .B(n20488), .Z(n20489) );
  AND U40236 ( .A(n22504), .B(n20489), .Z(n20490) );
  NANDN U40237 ( .A(x[7315]), .B(y[7315]), .Z(n50774) );
  AND U40238 ( .A(n20490), .B(n50774), .Z(n20492) );
  NANDN U40239 ( .A(y[7316]), .B(x[7316]), .Z(n20491) );
  NANDN U40240 ( .A(y[7317]), .B(x[7317]), .Z(n22500) );
  AND U40241 ( .A(n20491), .B(n22500), .Z(n60191) );
  NANDN U40242 ( .A(n20492), .B(n60191), .Z(n20493) );
  NAND U40243 ( .A(n20494), .B(n20493), .Z(n20495) );
  NAND U40244 ( .A(n60194), .B(n20495), .Z(n20496) );
  AND U40245 ( .A(n48342), .B(n20496), .Z(n20497) );
  NANDN U40246 ( .A(x[7319]), .B(y[7319]), .Z(n50773) );
  AND U40247 ( .A(n20497), .B(n50773), .Z(n20499) );
  NANDN U40248 ( .A(y[7320]), .B(x[7320]), .Z(n20498) );
  NANDN U40249 ( .A(y[7321]), .B(x[7321]), .Z(n22498) );
  NAND U40250 ( .A(n20498), .B(n22498), .Z(n60195) );
  OR U40251 ( .A(n20499), .B(n60195), .Z(n20500) );
  AND U40252 ( .A(n20501), .B(n20500), .Z(n20503) );
  NANDN U40253 ( .A(y[7322]), .B(x[7322]), .Z(n20502) );
  NANDN U40254 ( .A(y[7323]), .B(x[7323]), .Z(n48351) );
  AND U40255 ( .A(n20502), .B(n48351), .Z(n60198) );
  NANDN U40256 ( .A(n20503), .B(n60198), .Z(n20504) );
  AND U40257 ( .A(n48352), .B(n20504), .Z(n20505) );
  NANDN U40258 ( .A(x[7323]), .B(y[7323]), .Z(n60199) );
  NAND U40259 ( .A(n20505), .B(n60199), .Z(n20506) );
  NAND U40260 ( .A(n60200), .B(n20506), .Z(n20507) );
  ANDN U40261 ( .B(y[7325]), .A(x[7325]), .Z(n60201) );
  ANDN U40262 ( .B(n20507), .A(n60201), .Z(n20508) );
  XNOR U40263 ( .A(x[7326]), .B(y[7326]), .Z(n22497) );
  NAND U40264 ( .A(n20508), .B(n22497), .Z(n20509) );
  NAND U40265 ( .A(n60204), .B(n20509), .Z(n20510) );
  AND U40266 ( .A(n48362), .B(n20510), .Z(n20511) );
  NANDN U40267 ( .A(x[7327]), .B(y[7327]), .Z(n60205) );
  AND U40268 ( .A(n20511), .B(n60205), .Z(n20513) );
  NANDN U40269 ( .A(y[7328]), .B(x[7328]), .Z(n20512) );
  NANDN U40270 ( .A(y[7329]), .B(x[7329]), .Z(n22493) );
  AND U40271 ( .A(n20512), .B(n22493), .Z(n60207) );
  NANDN U40272 ( .A(n20513), .B(n60207), .Z(n20514) );
  AND U40273 ( .A(n22494), .B(n20514), .Z(n20515) );
  NANDN U40274 ( .A(x[7329]), .B(y[7329]), .Z(n22495) );
  AND U40275 ( .A(n20515), .B(n22495), .Z(n20517) );
  NANDN U40276 ( .A(y[7330]), .B(x[7330]), .Z(n20516) );
  NANDN U40277 ( .A(y[7331]), .B(x[7331]), .Z(n48371) );
  AND U40278 ( .A(n20516), .B(n48371), .Z(n60208) );
  NANDN U40279 ( .A(n20517), .B(n60208), .Z(n20518) );
  AND U40280 ( .A(n48372), .B(n20518), .Z(n20519) );
  NANDN U40281 ( .A(x[7331]), .B(y[7331]), .Z(n60209) );
  NAND U40282 ( .A(n20519), .B(n60209), .Z(n20520) );
  NAND U40283 ( .A(n60211), .B(n20520), .Z(n20521) );
  AND U40284 ( .A(n22492), .B(n20521), .Z(n20522) );
  ANDN U40285 ( .B(y[7333]), .A(x[7333]), .Z(n50767) );
  ANDN U40286 ( .B(n20522), .A(n50767), .Z(n20524) );
  NANDN U40287 ( .A(y[7334]), .B(x[7334]), .Z(n20523) );
  NANDN U40288 ( .A(y[7335]), .B(x[7335]), .Z(n48382) );
  AND U40289 ( .A(n20523), .B(n48382), .Z(n50766) );
  NANDN U40290 ( .A(n20524), .B(n50766), .Z(n20525) );
  NAND U40291 ( .A(n20526), .B(n20525), .Z(n20527) );
  NAND U40292 ( .A(n60214), .B(n20527), .Z(n20528) );
  AND U40293 ( .A(n22490), .B(n20528), .Z(n20529) );
  ANDN U40294 ( .B(y[7337]), .A(x[7337]), .Z(n60215) );
  ANDN U40295 ( .B(n20529), .A(n60215), .Z(n20531) );
  NANDN U40296 ( .A(y[7338]), .B(x[7338]), .Z(n20530) );
  NANDN U40297 ( .A(y[7339]), .B(x[7339]), .Z(n22487) );
  NAND U40298 ( .A(n20530), .B(n22487), .Z(n60218) );
  OR U40299 ( .A(n20531), .B(n60218), .Z(n20532) );
  NAND U40300 ( .A(n20533), .B(n20532), .Z(n20534) );
  NAND U40301 ( .A(n60221), .B(n20534), .Z(n20535) );
  AND U40302 ( .A(n22486), .B(n20535), .Z(n20536) );
  NANDN U40303 ( .A(x[7341]), .B(y[7341]), .Z(n60222) );
  AND U40304 ( .A(n20536), .B(n60222), .Z(n20538) );
  NANDN U40305 ( .A(y[7342]), .B(x[7342]), .Z(n20537) );
  NANDN U40306 ( .A(y[7343]), .B(x[7343]), .Z(n48400) );
  NAND U40307 ( .A(n20537), .B(n48400), .Z(n60224) );
  OR U40308 ( .A(n20538), .B(n60224), .Z(n20539) );
  NAND U40309 ( .A(n20540), .B(n20539), .Z(n20541) );
  NAND U40310 ( .A(n60225), .B(n20541), .Z(n20542) );
  AND U40311 ( .A(n22484), .B(n20542), .Z(n20543) );
  NANDN U40312 ( .A(n60226), .B(n20543), .Z(n20545) );
  NANDN U40313 ( .A(y[7346]), .B(x[7346]), .Z(n20544) );
  NANDN U40314 ( .A(y[7347]), .B(x[7347]), .Z(n22480) );
  AND U40315 ( .A(n20544), .B(n22480), .Z(n60228) );
  AND U40316 ( .A(n20545), .B(n60228), .Z(n20546) );
  XNOR U40317 ( .A(y[7348]), .B(x[7348]), .Z(n22481) );
  NANDN U40318 ( .A(x[7347]), .B(y[7347]), .Z(n22482) );
  NAND U40319 ( .A(n22481), .B(n22482), .Z(n50763) );
  OR U40320 ( .A(n20546), .B(n50763), .Z(n20547) );
  NAND U40321 ( .A(n50762), .B(n20547), .Z(n20548) );
  AND U40322 ( .A(n22478), .B(n20548), .Z(n20549) );
  NANDN U40323 ( .A(x[7349]), .B(y[7349]), .Z(n60230) );
  NAND U40324 ( .A(n20549), .B(n60230), .Z(n20550) );
  NAND U40325 ( .A(n60232), .B(n20550), .Z(n20551) );
  AND U40326 ( .A(n48419), .B(n20551), .Z(n20552) );
  NANDN U40327 ( .A(x[7351]), .B(y[7351]), .Z(n60233) );
  AND U40328 ( .A(n20552), .B(n60233), .Z(n20554) );
  NANDN U40329 ( .A(y[7352]), .B(x[7352]), .Z(n20553) );
  NANDN U40330 ( .A(y[7353]), .B(x[7353]), .Z(n22475) );
  AND U40331 ( .A(n20553), .B(n22475), .Z(n60235) );
  NANDN U40332 ( .A(n20554), .B(n60235), .Z(n20555) );
  NAND U40333 ( .A(n20556), .B(n20555), .Z(n20557) );
  NAND U40334 ( .A(n60236), .B(n20557), .Z(n20558) );
  AND U40335 ( .A(n48429), .B(n20558), .Z(n20559) );
  NANDN U40336 ( .A(x[7355]), .B(y[7355]), .Z(n60237) );
  AND U40337 ( .A(n20559), .B(n60237), .Z(n20561) );
  NANDN U40338 ( .A(y[7356]), .B(x[7356]), .Z(n20560) );
  NANDN U40339 ( .A(y[7357]), .B(x[7357]), .Z(n22473) );
  NAND U40340 ( .A(n20560), .B(n22473), .Z(n60239) );
  OR U40341 ( .A(n20561), .B(n60239), .Z(n20562) );
  NAND U40342 ( .A(n20563), .B(n20562), .Z(n20564) );
  NAND U40343 ( .A(n60243), .B(n20564), .Z(n20565) );
  AND U40344 ( .A(n22472), .B(n20565), .Z(n20566) );
  NANDN U40345 ( .A(x[7359]), .B(y[7359]), .Z(n60244) );
  AND U40346 ( .A(n20566), .B(n60244), .Z(n20568) );
  NANDN U40347 ( .A(y[7360]), .B(x[7360]), .Z(n20567) );
  NANDN U40348 ( .A(y[7361]), .B(x[7361]), .Z(n22469) );
  NAND U40349 ( .A(n20567), .B(n22469), .Z(n60246) );
  OR U40350 ( .A(n20568), .B(n60246), .Z(n20569) );
  NAND U40351 ( .A(n20570), .B(n20569), .Z(n20571) );
  NANDN U40352 ( .A(n50759), .B(n20571), .Z(n20572) );
  NAND U40353 ( .A(n60249), .B(n20572), .Z(n20573) );
  NAND U40354 ( .A(n60250), .B(n20573), .Z(n20574) );
  AND U40355 ( .A(n22467), .B(n20574), .Z(n20575) );
  NANDN U40356 ( .A(n60251), .B(n20575), .Z(n20576) );
  NANDN U40357 ( .A(n60253), .B(n20576), .Z(n20577) );
  AND U40358 ( .A(n48458), .B(n20577), .Z(n20578) );
  NANDN U40359 ( .A(x[7367]), .B(y[7367]), .Z(n50758) );
  NAND U40360 ( .A(n20578), .B(n50758), .Z(n20579) );
  NAND U40361 ( .A(n60254), .B(n20579), .Z(n20580) );
  AND U40362 ( .A(n22465), .B(n20580), .Z(n20581) );
  ANDN U40363 ( .B(y[7369]), .A(x[7369]), .Z(n60255) );
  ANDN U40364 ( .B(n20581), .A(n60255), .Z(n20583) );
  NANDN U40365 ( .A(y[7370]), .B(x[7370]), .Z(n20582) );
  NANDN U40366 ( .A(y[7371]), .B(x[7371]), .Z(n48468) );
  AND U40367 ( .A(n20582), .B(n48468), .Z(n60258) );
  NANDN U40368 ( .A(n20583), .B(n60258), .Z(n20584) );
  NAND U40369 ( .A(n20585), .B(n20584), .Z(n20586) );
  NAND U40370 ( .A(n60260), .B(n20586), .Z(n20587) );
  AND U40371 ( .A(n22463), .B(n20587), .Z(n20588) );
  ANDN U40372 ( .B(y[7373]), .A(x[7373]), .Z(n50753) );
  ANDN U40373 ( .B(n20588), .A(n50753), .Z(n20590) );
  NANDN U40374 ( .A(y[7374]), .B(x[7374]), .Z(n20589) );
  NANDN U40375 ( .A(y[7375]), .B(x[7375]), .Z(n48478) );
  NAND U40376 ( .A(n20589), .B(n48478), .Z(n60261) );
  OR U40377 ( .A(n20590), .B(n60261), .Z(n20591) );
  NAND U40378 ( .A(n20592), .B(n20591), .Z(n20593) );
  NAND U40379 ( .A(n60262), .B(n20593), .Z(n20594) );
  AND U40380 ( .A(n22460), .B(n20594), .Z(n20595) );
  NANDN U40381 ( .A(x[7377]), .B(y[7377]), .Z(n22461) );
  AND U40382 ( .A(n20595), .B(n22461), .Z(n20597) );
  NANDN U40383 ( .A(y[7378]), .B(x[7378]), .Z(n20596) );
  NANDN U40384 ( .A(y[7379]), .B(x[7379]), .Z(n22457) );
  NAND U40385 ( .A(n20596), .B(n22457), .Z(n50750) );
  OR U40386 ( .A(n20597), .B(n50750), .Z(n20598) );
  NAND U40387 ( .A(n20599), .B(n20598), .Z(n20600) );
  NAND U40388 ( .A(n60268), .B(n20600), .Z(n20601) );
  NAND U40389 ( .A(n60269), .B(n20601), .Z(n20602) );
  NAND U40390 ( .A(n60270), .B(n20602), .Z(n20603) );
  AND U40391 ( .A(n48497), .B(n20603), .Z(n20604) );
  NANDN U40392 ( .A(x[7383]), .B(y[7383]), .Z(n50749) );
  NAND U40393 ( .A(n20604), .B(n50749), .Z(n20605) );
  NAND U40394 ( .A(n60271), .B(n20605), .Z(n20606) );
  AND U40395 ( .A(n22452), .B(n20606), .Z(n20607) );
  NANDN U40396 ( .A(n60272), .B(n20607), .Z(n20608) );
  NAND U40397 ( .A(n60274), .B(n20608), .Z(n20609) );
  AND U40398 ( .A(n48507), .B(n20609), .Z(n20610) );
  NANDN U40399 ( .A(x[7387]), .B(y[7387]), .Z(n50747) );
  AND U40400 ( .A(n20610), .B(n50747), .Z(n20612) );
  NANDN U40401 ( .A(y[7388]), .B(x[7388]), .Z(n20611) );
  NANDN U40402 ( .A(y[7389]), .B(x[7389]), .Z(n22449) );
  AND U40403 ( .A(n20611), .B(n22449), .Z(n50745) );
  NANDN U40404 ( .A(n20612), .B(n50745), .Z(n20613) );
  NAND U40405 ( .A(n20614), .B(n20613), .Z(n20615) );
  NAND U40406 ( .A(n60277), .B(n20615), .Z(n20616) );
  NANDN U40407 ( .A(x[7391]), .B(y[7391]), .Z(n48514) );
  NANDN U40408 ( .A(x[7392]), .B(y[7392]), .Z(n22446) );
  AND U40409 ( .A(n48514), .B(n22446), .Z(n60278) );
  AND U40410 ( .A(n20616), .B(n60278), .Z(n20617) );
  NANDN U40411 ( .A(y[7392]), .B(x[7392]), .Z(n22447) );
  NANDN U40412 ( .A(y[7393]), .B(x[7393]), .Z(n22444) );
  NAND U40413 ( .A(n22447), .B(n22444), .Z(n50744) );
  OR U40414 ( .A(n20617), .B(n50744), .Z(n20618) );
  NAND U40415 ( .A(n20619), .B(n20618), .Z(n20620) );
  NAND U40416 ( .A(n60281), .B(n20620), .Z(n20621) );
  NAND U40417 ( .A(n60282), .B(n20621), .Z(n20622) );
  AND U40418 ( .A(n60283), .B(n20622), .Z(n20623) );
  OR U40419 ( .A(n20624), .B(n20623), .Z(n20625) );
  NAND U40420 ( .A(n50742), .B(n20625), .Z(n20626) );
  NANDN U40421 ( .A(n20627), .B(n20626), .Z(n20628) );
  AND U40422 ( .A(n60288), .B(n20628), .Z(n20629) );
  NOR U40423 ( .A(n60289), .B(n20629), .Z(n20630) );
  NAND U40424 ( .A(n22437), .B(n20630), .Z(n20631) );
  NANDN U40425 ( .A(n60291), .B(n20631), .Z(n20632) );
  AND U40426 ( .A(n48544), .B(n20632), .Z(n20633) );
  NANDN U40427 ( .A(x[7403]), .B(y[7403]), .Z(n60293) );
  NAND U40428 ( .A(n20633), .B(n60293), .Z(n20634) );
  NANDN U40429 ( .A(n60296), .B(n20634), .Z(n20635) );
  AND U40430 ( .A(n22435), .B(n20635), .Z(n20636) );
  NANDN U40431 ( .A(n60297), .B(n20636), .Z(n20637) );
  NAND U40432 ( .A(n60299), .B(n20637), .Z(n20638) );
  AND U40433 ( .A(n48554), .B(n20638), .Z(n20639) );
  NANDN U40434 ( .A(x[7407]), .B(y[7407]), .Z(n50741) );
  AND U40435 ( .A(n20639), .B(n50741), .Z(n20641) );
  NANDN U40436 ( .A(y[7408]), .B(x[7408]), .Z(n20640) );
  NANDN U40437 ( .A(y[7409]), .B(x[7409]), .Z(n22432) );
  AND U40438 ( .A(n20640), .B(n22432), .Z(n60300) );
  NANDN U40439 ( .A(n20641), .B(n60300), .Z(n20642) );
  NAND U40440 ( .A(n20643), .B(n20642), .Z(n20644) );
  NAND U40441 ( .A(n60303), .B(n20644), .Z(n20645) );
  AND U40442 ( .A(n48564), .B(n20645), .Z(n20646) );
  NANDN U40443 ( .A(x[7411]), .B(y[7411]), .Z(n60304) );
  AND U40444 ( .A(n20646), .B(n60304), .Z(n20648) );
  NANDN U40445 ( .A(y[7412]), .B(x[7412]), .Z(n20647) );
  NANDN U40446 ( .A(y[7413]), .B(x[7413]), .Z(n22430) );
  NAND U40447 ( .A(n20647), .B(n22430), .Z(n60306) );
  OR U40448 ( .A(n20648), .B(n60306), .Z(n20649) );
  NAND U40449 ( .A(n20650), .B(n20649), .Z(n20651) );
  NAND U40450 ( .A(n60310), .B(n20651), .Z(n20652) );
  AND U40451 ( .A(n48574), .B(n20652), .Z(n20653) );
  NANDN U40452 ( .A(x[7415]), .B(y[7415]), .Z(n60311) );
  AND U40453 ( .A(n20653), .B(n60311), .Z(n20655) );
  NANDN U40454 ( .A(y[7416]), .B(x[7416]), .Z(n20654) );
  NANDN U40455 ( .A(y[7417]), .B(x[7417]), .Z(n22428) );
  NAND U40456 ( .A(n20654), .B(n22428), .Z(n50739) );
  OR U40457 ( .A(n20655), .B(n50739), .Z(n20656) );
  NAND U40458 ( .A(n20657), .B(n20656), .Z(n20658) );
  NANDN U40459 ( .A(n60315), .B(n20658), .Z(n20659) );
  AND U40460 ( .A(n48584), .B(n20659), .Z(n20660) );
  NANDN U40461 ( .A(x[7419]), .B(y[7419]), .Z(n50738) );
  NAND U40462 ( .A(n20660), .B(n50738), .Z(n20662) );
  NANDN U40463 ( .A(y[7420]), .B(x[7420]), .Z(n20661) );
  NANDN U40464 ( .A(y[7421]), .B(x[7421]), .Z(n22426) );
  AND U40465 ( .A(n20661), .B(n22426), .Z(n50736) );
  AND U40466 ( .A(n20662), .B(n50736), .Z(n20664) );
  XNOR U40467 ( .A(x[7422]), .B(y[7422]), .Z(n22427) );
  ANDN U40468 ( .B(y[7421]), .A(x[7421]), .Z(n60317) );
  ANDN U40469 ( .B(n22427), .A(n60317), .Z(n20663) );
  NANDN U40470 ( .A(n20664), .B(n20663), .Z(n20665) );
  NANDN U40471 ( .A(n60318), .B(n20665), .Z(n20666) );
  AND U40472 ( .A(n22425), .B(n20666), .Z(n20667) );
  NANDN U40473 ( .A(x[7423]), .B(y[7423]), .Z(n60319) );
  NAND U40474 ( .A(n20667), .B(n60319), .Z(n20668) );
  AND U40475 ( .A(n60321), .B(n20668), .Z(n20669) );
  ANDN U40476 ( .B(n22423), .A(n20669), .Z(n20670) );
  NANDN U40477 ( .A(x[7425]), .B(y[7425]), .Z(n50734) );
  AND U40478 ( .A(n20670), .B(n50734), .Z(n20672) );
  NANDN U40479 ( .A(y[7426]), .B(x[7426]), .Z(n20671) );
  NANDN U40480 ( .A(y[7427]), .B(x[7427]), .Z(n22420) );
  AND U40481 ( .A(n20671), .B(n22420), .Z(n60324) );
  NANDN U40482 ( .A(n20672), .B(n60324), .Z(n20673) );
  NAND U40483 ( .A(n20674), .B(n20673), .Z(n20675) );
  NAND U40484 ( .A(n60325), .B(n20675), .Z(n20676) );
  AND U40485 ( .A(n22419), .B(n20676), .Z(n20677) );
  NANDN U40486 ( .A(x[7429]), .B(y[7429]), .Z(n60326) );
  AND U40487 ( .A(n20677), .B(n60326), .Z(n20678) );
  OR U40488 ( .A(n60328), .B(n20678), .Z(n20679) );
  NAND U40489 ( .A(n20680), .B(n20679), .Z(n20681) );
  NANDN U40490 ( .A(n60329), .B(n20681), .Z(n20682) );
  AND U40491 ( .A(n22417), .B(n20682), .Z(n20683) );
  NANDN U40492 ( .A(n60330), .B(n20683), .Z(n20684) );
  AND U40493 ( .A(n60332), .B(n20684), .Z(n20686) );
  XNOR U40494 ( .A(x[7436]), .B(y[7436]), .Z(n22415) );
  NANDN U40495 ( .A(x[7435]), .B(y[7435]), .Z(n60333) );
  AND U40496 ( .A(n22415), .B(n60333), .Z(n20685) );
  NANDN U40497 ( .A(n20686), .B(n20685), .Z(n20687) );
  NANDN U40498 ( .A(n60335), .B(n20687), .Z(n20688) );
  AND U40499 ( .A(n22413), .B(n20688), .Z(n20689) );
  NANDN U40500 ( .A(x[7437]), .B(y[7437]), .Z(n60336) );
  NAND U40501 ( .A(n20689), .B(n60336), .Z(n20690) );
  NAND U40502 ( .A(n60339), .B(n20690), .Z(n20691) );
  AND U40503 ( .A(n48629), .B(n20691), .Z(n20692) );
  NANDN U40504 ( .A(x[7439]), .B(y[7439]), .Z(n60340) );
  AND U40505 ( .A(n20692), .B(n60340), .Z(n20694) );
  NANDN U40506 ( .A(y[7440]), .B(x[7440]), .Z(n20693) );
  NANDN U40507 ( .A(y[7441]), .B(x[7441]), .Z(n22410) );
  AND U40508 ( .A(n20693), .B(n22410), .Z(n60342) );
  NANDN U40509 ( .A(n20694), .B(n60342), .Z(n20695) );
  NAND U40510 ( .A(n20696), .B(n20695), .Z(n20697) );
  NAND U40511 ( .A(n60343), .B(n20697), .Z(n20698) );
  AND U40512 ( .A(n48639), .B(n20698), .Z(n20699) );
  NANDN U40513 ( .A(x[7443]), .B(y[7443]), .Z(n60344) );
  AND U40514 ( .A(n20699), .B(n60344), .Z(n20701) );
  NANDN U40515 ( .A(y[7444]), .B(x[7444]), .Z(n20700) );
  NANDN U40516 ( .A(y[7445]), .B(x[7445]), .Z(n22408) );
  NAND U40517 ( .A(n20700), .B(n22408), .Z(n60346) );
  OR U40518 ( .A(n20701), .B(n60346), .Z(n20702) );
  AND U40519 ( .A(n20703), .B(n20702), .Z(n20705) );
  NANDN U40520 ( .A(y[7446]), .B(x[7446]), .Z(n20704) );
  NANDN U40521 ( .A(y[7447]), .B(x[7447]), .Z(n48649) );
  AND U40522 ( .A(n20704), .B(n48649), .Z(n50725) );
  NANDN U40523 ( .A(n20705), .B(n50725), .Z(n20706) );
  NAND U40524 ( .A(n20707), .B(n20706), .Z(n20708) );
  NAND U40525 ( .A(n60349), .B(n20708), .Z(n20709) );
  AND U40526 ( .A(n60350), .B(n20709), .Z(n20711) );
  NANDN U40527 ( .A(y[7450]), .B(x[7450]), .Z(n20710) );
  NANDN U40528 ( .A(y[7451]), .B(x[7451]), .Z(n48660) );
  AND U40529 ( .A(n20710), .B(n48660), .Z(n60352) );
  NANDN U40530 ( .A(n20711), .B(n60352), .Z(n20712) );
  NAND U40531 ( .A(n20713), .B(n20712), .Z(n20714) );
  AND U40532 ( .A(n60355), .B(n20714), .Z(n20716) );
  XNOR U40533 ( .A(x[7454]), .B(y[7454]), .Z(n22404) );
  ANDN U40534 ( .B(y[7453]), .A(x[7453]), .Z(n60356) );
  ANDN U40535 ( .B(n22404), .A(n60356), .Z(n20715) );
  NANDN U40536 ( .A(n20716), .B(n20715), .Z(n20717) );
  AND U40537 ( .A(n60358), .B(n20717), .Z(n20718) );
  ANDN U40538 ( .B(n60360), .A(n20718), .Z(n20719) );
  NAND U40539 ( .A(n48671), .B(n20719), .Z(n20720) );
  NANDN U40540 ( .A(n60361), .B(n20720), .Z(n20721) );
  AND U40541 ( .A(n22402), .B(n20721), .Z(n20722) );
  NANDN U40542 ( .A(n60362), .B(n20722), .Z(n20723) );
  AND U40543 ( .A(n60364), .B(n20723), .Z(n20725) );
  XNOR U40544 ( .A(x[7460]), .B(y[7460]), .Z(n48681) );
  NANDN U40545 ( .A(x[7459]), .B(y[7459]), .Z(n60365) );
  AND U40546 ( .A(n48681), .B(n60365), .Z(n20724) );
  NANDN U40547 ( .A(n20725), .B(n20724), .Z(n20726) );
  NANDN U40548 ( .A(n60367), .B(n20726), .Z(n20727) );
  AND U40549 ( .A(n22400), .B(n20727), .Z(n20728) );
  NANDN U40550 ( .A(x[7461]), .B(y[7461]), .Z(n50723) );
  NAND U40551 ( .A(n20728), .B(n50723), .Z(n20729) );
  NAND U40552 ( .A(n60370), .B(n20729), .Z(n20730) );
  NAND U40553 ( .A(n22397), .B(n20730), .Z(n20731) );
  ANDN U40554 ( .B(y[7463]), .A(x[7463]), .Z(n22398) );
  OR U40555 ( .A(n20731), .B(n22398), .Z(n20732) );
  NAND U40556 ( .A(n60373), .B(n20732), .Z(n20733) );
  NANDN U40557 ( .A(n50722), .B(n20733), .Z(n20734) );
  NAND U40558 ( .A(n60374), .B(n20734), .Z(n20735) );
  NAND U40559 ( .A(n60375), .B(n20735), .Z(n20736) );
  AND U40560 ( .A(n60376), .B(n20736), .Z(n20737) );
  NOR U40561 ( .A(n22391), .B(n20737), .Z(n20738) );
  NAND U40562 ( .A(n22390), .B(n20738), .Z(n20739) );
  NANDN U40563 ( .A(n60379), .B(n20739), .Z(n20740) );
  AND U40564 ( .A(n48712), .B(n20740), .Z(n20741) );
  NANDN U40565 ( .A(n50721), .B(n20741), .Z(n20742) );
  AND U40566 ( .A(n60380), .B(n20742), .Z(n20744) );
  XNOR U40567 ( .A(x[7474]), .B(y[7474]), .Z(n22388) );
  ANDN U40568 ( .B(y[7473]), .A(x[7473]), .Z(n60381) );
  ANDN U40569 ( .B(n22388), .A(n60381), .Z(n20743) );
  NANDN U40570 ( .A(n20744), .B(n20743), .Z(n20745) );
  NANDN U40571 ( .A(n60384), .B(n20745), .Z(n20746) );
  AND U40572 ( .A(n48722), .B(n20746), .Z(n20747) );
  NANDN U40573 ( .A(x[7475]), .B(y[7475]), .Z(n50719) );
  AND U40574 ( .A(n20747), .B(n50719), .Z(n20749) );
  NANDN U40575 ( .A(y[7476]), .B(x[7476]), .Z(n20748) );
  NANDN U40576 ( .A(y[7477]), .B(x[7477]), .Z(n22385) );
  AND U40577 ( .A(n20748), .B(n22385), .Z(n50717) );
  NANDN U40578 ( .A(n20749), .B(n50717), .Z(n20750) );
  AND U40579 ( .A(n60385), .B(n20750), .Z(n20751) );
  NANDN U40580 ( .A(y[7478]), .B(x[7478]), .Z(n22384) );
  NANDN U40581 ( .A(y[7479]), .B(x[7479]), .Z(n22381) );
  NAND U40582 ( .A(n22384), .B(n22381), .Z(n60386) );
  OR U40583 ( .A(n20751), .B(n60386), .Z(n20752) );
  NAND U40584 ( .A(n20753), .B(n20752), .Z(n20754) );
  NANDN U40585 ( .A(n50714), .B(n20754), .Z(n20755) );
  AND U40586 ( .A(n22380), .B(n20755), .Z(n20756) );
  NANDN U40587 ( .A(x[7481]), .B(y[7481]), .Z(n50713) );
  AND U40588 ( .A(n20756), .B(n50713), .Z(n20758) );
  NANDN U40589 ( .A(y[7482]), .B(x[7482]), .Z(n20757) );
  NANDN U40590 ( .A(y[7483]), .B(x[7483]), .Z(n22378) );
  AND U40591 ( .A(n20757), .B(n22378), .Z(n60387) );
  NANDN U40592 ( .A(n20758), .B(n60387), .Z(n20759) );
  AND U40593 ( .A(n60388), .B(n20759), .Z(n20760) );
  NANDN U40594 ( .A(y[7484]), .B(x[7484]), .Z(n22377) );
  NANDN U40595 ( .A(y[7485]), .B(x[7485]), .Z(n22374) );
  NAND U40596 ( .A(n22377), .B(n22374), .Z(n60389) );
  OR U40597 ( .A(n20760), .B(n60389), .Z(n20761) );
  NAND U40598 ( .A(n60390), .B(n20761), .Z(n20762) );
  NAND U40599 ( .A(n60392), .B(n20762), .Z(n20763) );
  AND U40600 ( .A(n60393), .B(n20763), .Z(n20764) );
  NANDN U40601 ( .A(y[7488]), .B(x[7488]), .Z(n22369) );
  NANDN U40602 ( .A(y[7489]), .B(x[7489]), .Z(n22368) );
  AND U40603 ( .A(n22369), .B(n22368), .Z(n60394) );
  NANDN U40604 ( .A(n20764), .B(n60394), .Z(n20765) );
  NAND U40605 ( .A(n60395), .B(n20765), .Z(n20766) );
  NANDN U40606 ( .A(n60396), .B(n20766), .Z(n20767) );
  NAND U40607 ( .A(n60397), .B(n20767), .Z(n20768) );
  NAND U40608 ( .A(n60398), .B(n20768), .Z(n20769) );
  AND U40609 ( .A(n60399), .B(n20769), .Z(n20770) );
  NANDN U40610 ( .A(y[7494]), .B(x[7494]), .Z(n22359) );
  NANDN U40611 ( .A(y[7495]), .B(x[7495]), .Z(n22356) );
  AND U40612 ( .A(n22359), .B(n22356), .Z(n60400) );
  NANDN U40613 ( .A(n20770), .B(n60400), .Z(n20771) );
  NAND U40614 ( .A(n60401), .B(n20771), .Z(n20772) );
  NANDN U40615 ( .A(n60402), .B(n20772), .Z(n20773) );
  AND U40616 ( .A(n22354), .B(n20773), .Z(n20774) );
  NANDN U40617 ( .A(x[7497]), .B(y[7497]), .Z(n50711) );
  NAND U40618 ( .A(n20774), .B(n50711), .Z(n20775) );
  AND U40619 ( .A(n60403), .B(n20775), .Z(n20777) );
  XNOR U40620 ( .A(x[7500]), .B(y[7500]), .Z(n48776) );
  NANDN U40621 ( .A(x[7499]), .B(y[7499]), .Z(n60404) );
  AND U40622 ( .A(n48776), .B(n60404), .Z(n20776) );
  NANDN U40623 ( .A(n20777), .B(n20776), .Z(n20778) );
  NANDN U40624 ( .A(n60406), .B(n20778), .Z(n20779) );
  AND U40625 ( .A(n22352), .B(n20779), .Z(n20780) );
  NANDN U40626 ( .A(n50708), .B(n20780), .Z(n20782) );
  NANDN U40627 ( .A(y[7502]), .B(x[7502]), .Z(n20781) );
  NANDN U40628 ( .A(y[7503]), .B(x[7503]), .Z(n48785) );
  AND U40629 ( .A(n20781), .B(n48785), .Z(n50707) );
  AND U40630 ( .A(n20782), .B(n50707), .Z(n20783) );
  OR U40631 ( .A(n20784), .B(n20783), .Z(n20785) );
  NAND U40632 ( .A(n60410), .B(n20785), .Z(n20786) );
  NANDN U40633 ( .A(n20787), .B(n20786), .Z(n20788) );
  NAND U40634 ( .A(n60413), .B(n20788), .Z(n20789) );
  AND U40635 ( .A(n48796), .B(n20789), .Z(n20790) );
  NANDN U40636 ( .A(x[7507]), .B(y[7507]), .Z(n60414) );
  AND U40637 ( .A(n20790), .B(n60414), .Z(n20791) );
  OR U40638 ( .A(n60416), .B(n20791), .Z(n20792) );
  NAND U40639 ( .A(n20793), .B(n20792), .Z(n20794) );
  NANDN U40640 ( .A(n60417), .B(n20794), .Z(n20795) );
  AND U40641 ( .A(n48807), .B(n20795), .Z(n20796) );
  NANDN U40642 ( .A(n60419), .B(n20796), .Z(n20798) );
  NANDN U40643 ( .A(y[7512]), .B(x[7512]), .Z(n20797) );
  NANDN U40644 ( .A(y[7513]), .B(x[7513]), .Z(n22345) );
  AND U40645 ( .A(n20797), .B(n22345), .Z(n50704) );
  AND U40646 ( .A(n20798), .B(n50704), .Z(n20800) );
  XNOR U40647 ( .A(x[7514]), .B(y[7514]), .Z(n22346) );
  ANDN U40648 ( .B(y[7513]), .A(x[7513]), .Z(n60421) );
  ANDN U40649 ( .B(n22346), .A(n60421), .Z(n20799) );
  NANDN U40650 ( .A(n20800), .B(n20799), .Z(n20801) );
  NANDN U40651 ( .A(n60423), .B(n20801), .Z(n20802) );
  AND U40652 ( .A(n48817), .B(n20802), .Z(n20803) );
  NANDN U40653 ( .A(x[7515]), .B(y[7515]), .Z(n60424) );
  NAND U40654 ( .A(n20803), .B(n60424), .Z(n20804) );
  NAND U40655 ( .A(n60426), .B(n20804), .Z(n20805) );
  AND U40656 ( .A(n22344), .B(n20805), .Z(n20806) );
  NANDN U40657 ( .A(n50702), .B(n20806), .Z(n20807) );
  NAND U40658 ( .A(n60427), .B(n20807), .Z(n20808) );
  NANDN U40659 ( .A(x[7519]), .B(y[7519]), .Z(n60429) );
  AND U40660 ( .A(n20808), .B(n60429), .Z(n20809) );
  NAND U40661 ( .A(n48827), .B(n20809), .Z(n20810) );
  NAND U40662 ( .A(n60430), .B(n20810), .Z(n20811) );
  AND U40663 ( .A(n22342), .B(n20811), .Z(n20812) );
  ANDN U40664 ( .B(y[7521]), .A(x[7521]), .Z(n60431) );
  ANDN U40665 ( .B(n20812), .A(n60431), .Z(n20814) );
  NANDN U40666 ( .A(y[7522]), .B(x[7522]), .Z(n20813) );
  NANDN U40667 ( .A(y[7523]), .B(x[7523]), .Z(n48836) );
  NAND U40668 ( .A(n20813), .B(n48836), .Z(n60433) );
  OR U40669 ( .A(n20814), .B(n60433), .Z(n20815) );
  NAND U40670 ( .A(n20816), .B(n20815), .Z(n20817) );
  NAND U40671 ( .A(n60437), .B(n20817), .Z(n20818) );
  AND U40672 ( .A(n22340), .B(n20818), .Z(n20819) );
  ANDN U40673 ( .B(y[7525]), .A(x[7525]), .Z(n60438) );
  ANDN U40674 ( .B(n20819), .A(n60438), .Z(n20821) );
  NANDN U40675 ( .A(y[7526]), .B(x[7526]), .Z(n20820) );
  NANDN U40676 ( .A(y[7527]), .B(x[7527]), .Z(n48846) );
  NAND U40677 ( .A(n20820), .B(n48846), .Z(n60440) );
  OR U40678 ( .A(n20821), .B(n60440), .Z(n20822) );
  NAND U40679 ( .A(n20823), .B(n20822), .Z(n20824) );
  NAND U40680 ( .A(n60441), .B(n20824), .Z(n20825) );
  AND U40681 ( .A(n22338), .B(n20825), .Z(n20826) );
  NANDN U40682 ( .A(n60442), .B(n20826), .Z(n20828) );
  NANDN U40683 ( .A(y[7530]), .B(x[7530]), .Z(n20827) );
  NANDN U40684 ( .A(y[7531]), .B(x[7531]), .Z(n48856) );
  AND U40685 ( .A(n20827), .B(n48856), .Z(n60444) );
  AND U40686 ( .A(n20828), .B(n60444), .Z(n20830) );
  XNOR U40687 ( .A(x[7532]), .B(y[7532]), .Z(n48857) );
  NANDN U40688 ( .A(x[7531]), .B(y[7531]), .Z(n50699) );
  AND U40689 ( .A(n48857), .B(n50699), .Z(n20829) );
  NANDN U40690 ( .A(n20830), .B(n20829), .Z(n20831) );
  NANDN U40691 ( .A(n60445), .B(n20831), .Z(n20832) );
  AND U40692 ( .A(n22336), .B(n20832), .Z(n20833) );
  NANDN U40693 ( .A(n60446), .B(n20833), .Z(n20834) );
  NAND U40694 ( .A(n60448), .B(n20834), .Z(n20835) );
  AND U40695 ( .A(n48867), .B(n20835), .Z(n20836) );
  NANDN U40696 ( .A(x[7535]), .B(y[7535]), .Z(n60450) );
  AND U40697 ( .A(n20836), .B(n60450), .Z(n20838) );
  NANDN U40698 ( .A(y[7536]), .B(x[7536]), .Z(n20837) );
  NANDN U40699 ( .A(y[7537]), .B(x[7537]), .Z(n22333) );
  AND U40700 ( .A(n20837), .B(n22333), .Z(n50697) );
  NANDN U40701 ( .A(n20838), .B(n50697), .Z(n20839) );
  NAND U40702 ( .A(n20840), .B(n20839), .Z(n20841) );
  NAND U40703 ( .A(n60454), .B(n20841), .Z(n20842) );
  AND U40704 ( .A(n48877), .B(n20842), .Z(n20843) );
  NANDN U40705 ( .A(x[7539]), .B(y[7539]), .Z(n60455) );
  AND U40706 ( .A(n20843), .B(n60455), .Z(n20845) );
  NANDN U40707 ( .A(y[7540]), .B(x[7540]), .Z(n20844) );
  NANDN U40708 ( .A(y[7541]), .B(x[7541]), .Z(n22330) );
  NAND U40709 ( .A(n20844), .B(n22330), .Z(n60457) );
  OR U40710 ( .A(n20845), .B(n60457), .Z(n20846) );
  NAND U40711 ( .A(n20847), .B(n20846), .Z(n20848) );
  NAND U40712 ( .A(n60458), .B(n20848), .Z(n20849) );
  AND U40713 ( .A(n48887), .B(n20849), .Z(n20850) );
  NANDN U40714 ( .A(x[7543]), .B(y[7543]), .Z(n60459) );
  NAND U40715 ( .A(n20850), .B(n60459), .Z(n20852) );
  NANDN U40716 ( .A(y[7544]), .B(x[7544]), .Z(n20851) );
  NANDN U40717 ( .A(y[7545]), .B(x[7545]), .Z(n22328) );
  AND U40718 ( .A(n20851), .B(n22328), .Z(n60461) );
  AND U40719 ( .A(n20852), .B(n60461), .Z(n20854) );
  XNOR U40720 ( .A(x[7546]), .B(y[7546]), .Z(n22329) );
  ANDN U40721 ( .B(y[7545]), .A(x[7545]), .Z(n50693) );
  ANDN U40722 ( .B(n22329), .A(n50693), .Z(n20853) );
  NANDN U40723 ( .A(n20854), .B(n20853), .Z(n20855) );
  NANDN U40724 ( .A(n60464), .B(n20855), .Z(n20856) );
  AND U40725 ( .A(n48897), .B(n20856), .Z(n20857) );
  NANDN U40726 ( .A(x[7547]), .B(y[7547]), .Z(n60465) );
  NAND U40727 ( .A(n20857), .B(n60465), .Z(n20858) );
  AND U40728 ( .A(n60467), .B(n20858), .Z(n20859) );
  OR U40729 ( .A(n20860), .B(n20859), .Z(n20861) );
  NAND U40730 ( .A(n50692), .B(n20861), .Z(n20862) );
  NANDN U40731 ( .A(n20863), .B(n20862), .Z(n20864) );
  NAND U40732 ( .A(n60472), .B(n20864), .Z(n20865) );
  AND U40733 ( .A(n22325), .B(n20865), .Z(n20866) );
  ANDN U40734 ( .B(y[7553]), .A(x[7553]), .Z(n60473) );
  ANDN U40735 ( .B(n20866), .A(n60473), .Z(n20867) );
  OR U40736 ( .A(n60475), .B(n20867), .Z(n20868) );
  NAND U40737 ( .A(n20869), .B(n20868), .Z(n20870) );
  NAND U40738 ( .A(n60476), .B(n20870), .Z(n20871) );
  AND U40739 ( .A(n22323), .B(n20871), .Z(n20872) );
  NANDN U40740 ( .A(n60477), .B(n20872), .Z(n20874) );
  NANDN U40741 ( .A(y[7558]), .B(x[7558]), .Z(n20873) );
  NANDN U40742 ( .A(y[7559]), .B(x[7559]), .Z(n48926) );
  AND U40743 ( .A(n20873), .B(n48926), .Z(n60480) );
  AND U40744 ( .A(n20874), .B(n60480), .Z(n20876) );
  XNOR U40745 ( .A(x[7560]), .B(y[7560]), .Z(n48927) );
  NANDN U40746 ( .A(x[7559]), .B(y[7559]), .Z(n50689) );
  AND U40747 ( .A(n48927), .B(n50689), .Z(n20875) );
  NANDN U40748 ( .A(n20876), .B(n20875), .Z(n20877) );
  NANDN U40749 ( .A(n60482), .B(n20877), .Z(n20878) );
  AND U40750 ( .A(n22321), .B(n20878), .Z(n20879) );
  NANDN U40751 ( .A(n60483), .B(n20879), .Z(n20880) );
  NAND U40752 ( .A(n60485), .B(n20880), .Z(n20881) );
  AND U40753 ( .A(n48937), .B(n20881), .Z(n20882) );
  NANDN U40754 ( .A(x[7563]), .B(y[7563]), .Z(n60486) );
  AND U40755 ( .A(n20882), .B(n60486), .Z(n20884) );
  NANDN U40756 ( .A(y[7564]), .B(x[7564]), .Z(n20883) );
  NANDN U40757 ( .A(y[7565]), .B(x[7565]), .Z(n22318) );
  AND U40758 ( .A(n20883), .B(n22318), .Z(n50687) );
  NANDN U40759 ( .A(n20884), .B(n50687), .Z(n20885) );
  NAND U40760 ( .A(n20886), .B(n20885), .Z(n20887) );
  AND U40761 ( .A(n60490), .B(n20887), .Z(n20888) );
  ANDN U40762 ( .B(n60492), .A(n20888), .Z(n20889) );
  NAND U40763 ( .A(n48947), .B(n20889), .Z(n20890) );
  NANDN U40764 ( .A(n60493), .B(n20890), .Z(n20891) );
  AND U40765 ( .A(n22317), .B(n20891), .Z(n20892) );
  NANDN U40766 ( .A(n60496), .B(n20892), .Z(n20893) );
  NANDN U40767 ( .A(n60497), .B(n20893), .Z(n20894) );
  AND U40768 ( .A(n48957), .B(n20894), .Z(n20895) );
  NANDN U40769 ( .A(x[7571]), .B(y[7571]), .Z(n60498) );
  AND U40770 ( .A(n20895), .B(n60498), .Z(n20897) );
  NANDN U40771 ( .A(y[7572]), .B(x[7572]), .Z(n20896) );
  NANDN U40772 ( .A(y[7573]), .B(x[7573]), .Z(n22314) );
  NAND U40773 ( .A(n20896), .B(n22314), .Z(n60500) );
  OR U40774 ( .A(n20897), .B(n60500), .Z(n20898) );
  NAND U40775 ( .A(n60501), .B(n20898), .Z(n20899) );
  NANDN U40776 ( .A(n50686), .B(n20899), .Z(n20900) );
  AND U40777 ( .A(n22311), .B(n20900), .Z(n20901) );
  NAND U40778 ( .A(n50685), .B(n20901), .Z(n20902) );
  NAND U40779 ( .A(n60503), .B(n20902), .Z(n20903) );
  AND U40780 ( .A(n22309), .B(n20903), .Z(n20904) );
  ANDN U40781 ( .B(y[7577]), .A(x[7577]), .Z(n60504) );
  ANDN U40782 ( .B(n20904), .A(n60504), .Z(n20905) );
  OR U40783 ( .A(n60506), .B(n20905), .Z(n20906) );
  NAND U40784 ( .A(n60507), .B(n20906), .Z(n20907) );
  NANDN U40785 ( .A(n60508), .B(n20907), .Z(n20908) );
  AND U40786 ( .A(n60510), .B(n20908), .Z(n20910) );
  NAND U40787 ( .A(n20910), .B(n20909), .Z(n20911) );
  NANDN U40788 ( .A(n60512), .B(n20911), .Z(n20912) );
  AND U40789 ( .A(n48984), .B(n20912), .Z(n20913) );
  NANDN U40790 ( .A(x[7583]), .B(y[7583]), .Z(n50684) );
  NAND U40791 ( .A(n20913), .B(n50684), .Z(n20914) );
  AND U40792 ( .A(n60513), .B(n20914), .Z(n20916) );
  XNOR U40793 ( .A(x[7586]), .B(y[7586]), .Z(n22302) );
  ANDN U40794 ( .B(y[7585]), .A(x[7585]), .Z(n50682) );
  ANDN U40795 ( .B(n22302), .A(n50682), .Z(n20915) );
  NANDN U40796 ( .A(n20916), .B(n20915), .Z(n20917) );
  NAND U40797 ( .A(n60514), .B(n20917), .Z(n20918) );
  AND U40798 ( .A(n48994), .B(n20918), .Z(n20919) );
  NANDN U40799 ( .A(x[7587]), .B(y[7587]), .Z(n60515) );
  NAND U40800 ( .A(n20919), .B(n60515), .Z(n20920) );
  NAND U40801 ( .A(n60517), .B(n20920), .Z(n20921) );
  AND U40802 ( .A(n22300), .B(n20921), .Z(n20922) );
  ANDN U40803 ( .B(y[7589]), .A(x[7589]), .Z(n50679) );
  ANDN U40804 ( .B(n20922), .A(n50679), .Z(n20924) );
  NANDN U40805 ( .A(y[7590]), .B(x[7590]), .Z(n20923) );
  NANDN U40806 ( .A(y[7591]), .B(x[7591]), .Z(n49004) );
  AND U40807 ( .A(n20923), .B(n49004), .Z(n50678) );
  NANDN U40808 ( .A(n20924), .B(n50678), .Z(n20925) );
  NAND U40809 ( .A(n20926), .B(n20925), .Z(n20927) );
  NAND U40810 ( .A(n60521), .B(n20927), .Z(n20928) );
  AND U40811 ( .A(n22298), .B(n20928), .Z(n20929) );
  ANDN U40812 ( .B(y[7593]), .A(x[7593]), .Z(n60522) );
  ANDN U40813 ( .B(n20929), .A(n60522), .Z(n20931) );
  NANDN U40814 ( .A(y[7594]), .B(x[7594]), .Z(n20930) );
  NANDN U40815 ( .A(y[7595]), .B(x[7595]), .Z(n49014) );
  NAND U40816 ( .A(n20930), .B(n49014), .Z(n60524) );
  OR U40817 ( .A(n20931), .B(n60524), .Z(n20932) );
  NAND U40818 ( .A(n20933), .B(n20932), .Z(n20934) );
  NAND U40819 ( .A(n60527), .B(n20934), .Z(n20935) );
  AND U40820 ( .A(n22296), .B(n20935), .Z(n20936) );
  ANDN U40821 ( .B(y[7597]), .A(x[7597]), .Z(n60528) );
  ANDN U40822 ( .B(n20936), .A(n60528), .Z(n20938) );
  NANDN U40823 ( .A(y[7598]), .B(x[7598]), .Z(n20937) );
  NANDN U40824 ( .A(y[7599]), .B(x[7599]), .Z(n49024) );
  NAND U40825 ( .A(n20937), .B(n49024), .Z(n60530) );
  OR U40826 ( .A(n20938), .B(n60530), .Z(n20939) );
  NAND U40827 ( .A(n20940), .B(n20939), .Z(n20941) );
  NAND U40828 ( .A(n60531), .B(n20941), .Z(n20942) );
  AND U40829 ( .A(n22294), .B(n20942), .Z(n20943) );
  NANDN U40830 ( .A(n60532), .B(n20943), .Z(n20945) );
  NANDN U40831 ( .A(y[7602]), .B(x[7602]), .Z(n20944) );
  NANDN U40832 ( .A(y[7603]), .B(x[7603]), .Z(n49034) );
  AND U40833 ( .A(n20944), .B(n49034), .Z(n60534) );
  AND U40834 ( .A(n20945), .B(n60534), .Z(n20947) );
  XNOR U40835 ( .A(x[7604]), .B(y[7604]), .Z(n49035) );
  NANDN U40836 ( .A(x[7603]), .B(y[7603]), .Z(n50675) );
  AND U40837 ( .A(n49035), .B(n50675), .Z(n20946) );
  NANDN U40838 ( .A(n20947), .B(n20946), .Z(n20948) );
  NANDN U40839 ( .A(n60537), .B(n20948), .Z(n20949) );
  AND U40840 ( .A(n22292), .B(n20949), .Z(n20950) );
  NANDN U40841 ( .A(n60538), .B(n20950), .Z(n20951) );
  AND U40842 ( .A(n60540), .B(n20951), .Z(n20952) );
  NOR U40843 ( .A(n49042), .B(n20952), .Z(n20953) );
  NAND U40844 ( .A(n49046), .B(n20953), .Z(n20954) );
  NANDN U40845 ( .A(n60542), .B(n20954), .Z(n20955) );
  AND U40846 ( .A(n22290), .B(n20955), .Z(n20956) );
  NANDN U40847 ( .A(n60543), .B(n20956), .Z(n20957) );
  NAND U40848 ( .A(n60545), .B(n20957), .Z(n20958) );
  AND U40849 ( .A(n49056), .B(n20958), .Z(n20959) );
  NANDN U40850 ( .A(x[7611]), .B(y[7611]), .Z(n60546) );
  NAND U40851 ( .A(n20959), .B(n60546), .Z(n20960) );
  AND U40852 ( .A(n60548), .B(n20960), .Z(n20962) );
  XNOR U40853 ( .A(x[7614]), .B(y[7614]), .Z(n22287) );
  NANDN U40854 ( .A(x[7613]), .B(y[7613]), .Z(n22288) );
  AND U40855 ( .A(n22287), .B(n22288), .Z(n20961) );
  NANDN U40856 ( .A(n20962), .B(n20961), .Z(n20963) );
  NAND U40857 ( .A(n60549), .B(n20963), .Z(n20964) );
  AND U40858 ( .A(n49066), .B(n20964), .Z(n20965) );
  NANDN U40859 ( .A(x[7615]), .B(y[7615]), .Z(n60550) );
  NAND U40860 ( .A(n20965), .B(n60550), .Z(n20966) );
  NAND U40861 ( .A(n60552), .B(n20966), .Z(n20967) );
  NAND U40862 ( .A(n22285), .B(n20967), .Z(n20968) );
  ANDN U40863 ( .B(y[7617]), .A(x[7617]), .Z(n50668) );
  OR U40864 ( .A(n20968), .B(n50668), .Z(n20969) );
  NAND U40865 ( .A(n50667), .B(n20969), .Z(n20970) );
  NAND U40866 ( .A(n60554), .B(n20970), .Z(n20971) );
  NAND U40867 ( .A(n60555), .B(n20971), .Z(n20972) );
  AND U40868 ( .A(n22279), .B(n20972), .Z(n20973) );
  NANDN U40869 ( .A(x[7621]), .B(y[7621]), .Z(n50665) );
  AND U40870 ( .A(n20973), .B(n50665), .Z(n20975) );
  NANDN U40871 ( .A(y[7622]), .B(x[7622]), .Z(n20974) );
  NANDN U40872 ( .A(y[7623]), .B(x[7623]), .Z(n49083) );
  NAND U40873 ( .A(n20974), .B(n49083), .Z(n50664) );
  OR U40874 ( .A(n20975), .B(n50664), .Z(n20976) );
  AND U40875 ( .A(n20977), .B(n20976), .Z(n20979) );
  NANDN U40876 ( .A(y[7624]), .B(x[7624]), .Z(n20978) );
  NANDN U40877 ( .A(y[7625]), .B(x[7625]), .Z(n22276) );
  AND U40878 ( .A(n20978), .B(n22276), .Z(n60556) );
  NANDN U40879 ( .A(n20979), .B(n60556), .Z(n20980) );
  NAND U40880 ( .A(n20981), .B(n20980), .Z(n20982) );
  NAND U40881 ( .A(n60559), .B(n20982), .Z(n20983) );
  AND U40882 ( .A(n22275), .B(n20983), .Z(n20984) );
  NANDN U40883 ( .A(x[7627]), .B(y[7627]), .Z(n50660) );
  AND U40884 ( .A(n20984), .B(n50660), .Z(n20985) );
  OR U40885 ( .A(n60561), .B(n20985), .Z(n20986) );
  AND U40886 ( .A(n22273), .B(n20986), .Z(n20987) );
  NANDN U40887 ( .A(x[7629]), .B(y[7629]), .Z(n60562) );
  NAND U40888 ( .A(n20987), .B(n60562), .Z(n20988) );
  AND U40889 ( .A(n60564), .B(n20988), .Z(n20989) );
  NANDN U40890 ( .A(x[7631]), .B(y[7631]), .Z(n60565) );
  NANDN U40891 ( .A(n20989), .B(n60565), .Z(n20990) );
  XNOR U40892 ( .A(x[7632]), .B(y[7632]), .Z(n49102) );
  NANDN U40893 ( .A(n20990), .B(n49102), .Z(n20991) );
  NAND U40894 ( .A(n50658), .B(n20991), .Z(n20992) );
  NANDN U40895 ( .A(n20993), .B(n20992), .Z(n20994) );
  NAND U40896 ( .A(n60567), .B(n20994), .Z(n20995) );
  AND U40897 ( .A(n22269), .B(n20995), .Z(n20996) );
  NANDN U40898 ( .A(x[7635]), .B(y[7635]), .Z(n60568) );
  AND U40899 ( .A(n20996), .B(n60568), .Z(n20997) );
  OR U40900 ( .A(n60570), .B(n20997), .Z(n20998) );
  NAND U40901 ( .A(n20999), .B(n20998), .Z(n21000) );
  NANDN U40902 ( .A(n60571), .B(n21000), .Z(n21001) );
  AND U40903 ( .A(n49120), .B(n21001), .Z(n21002) );
  NANDN U40904 ( .A(x[7639]), .B(y[7639]), .Z(n60572) );
  NAND U40905 ( .A(n21002), .B(n60572), .Z(n21003) );
  AND U40906 ( .A(n60575), .B(n21003), .Z(n21004) );
  NOR U40907 ( .A(n60576), .B(n21004), .Z(n21005) );
  NAND U40908 ( .A(n22265), .B(n21005), .Z(n21006) );
  NANDN U40909 ( .A(n60578), .B(n21006), .Z(n21007) );
  AND U40910 ( .A(n49131), .B(n21007), .Z(n21008) );
  NANDN U40911 ( .A(n60580), .B(n21008), .Z(n21010) );
  NANDN U40912 ( .A(y[7644]), .B(x[7644]), .Z(n21009) );
  NANDN U40913 ( .A(y[7645]), .B(x[7645]), .Z(n22262) );
  AND U40914 ( .A(n21009), .B(n22262), .Z(n50654) );
  AND U40915 ( .A(n21010), .B(n50654), .Z(n21011) );
  OR U40916 ( .A(n21012), .B(n21011), .Z(n21013) );
  NAND U40917 ( .A(n60583), .B(n21013), .Z(n21014) );
  NANDN U40918 ( .A(n21015), .B(n21014), .Z(n21016) );
  NAND U40919 ( .A(n60584), .B(n21016), .Z(n21017) );
  AND U40920 ( .A(n22261), .B(n21017), .Z(n21018) );
  ANDN U40921 ( .B(y[7649]), .A(x[7649]), .Z(n60585) );
  ANDN U40922 ( .B(n21018), .A(n60585), .Z(n21020) );
  NANDN U40923 ( .A(y[7650]), .B(x[7650]), .Z(n21019) );
  NANDN U40924 ( .A(y[7651]), .B(x[7651]), .Z(n49150) );
  NAND U40925 ( .A(n21019), .B(n49150), .Z(n60588) );
  OR U40926 ( .A(n21020), .B(n60588), .Z(n21021) );
  NAND U40927 ( .A(n21022), .B(n21021), .Z(n21023) );
  NANDN U40928 ( .A(n60593), .B(n21023), .Z(n21024) );
  AND U40929 ( .A(n22259), .B(n21024), .Z(n21025) );
  NANDN U40930 ( .A(n60594), .B(n21025), .Z(n21026) );
  AND U40931 ( .A(n60596), .B(n21026), .Z(n21028) );
  XNOR U40932 ( .A(x[7656]), .B(y[7656]), .Z(n49161) );
  NANDN U40933 ( .A(x[7655]), .B(y[7655]), .Z(n60597) );
  AND U40934 ( .A(n49161), .B(n60597), .Z(n21027) );
  NANDN U40935 ( .A(n21028), .B(n21027), .Z(n21029) );
  NANDN U40936 ( .A(n50651), .B(n21029), .Z(n21030) );
  AND U40937 ( .A(n22256), .B(n21030), .Z(n21031) );
  NANDN U40938 ( .A(x[7657]), .B(y[7657]), .Z(n22257) );
  AND U40939 ( .A(n21031), .B(n22257), .Z(n21033) );
  NANDN U40940 ( .A(y[7658]), .B(x[7658]), .Z(n21032) );
  NANDN U40941 ( .A(y[7659]), .B(x[7659]), .Z(n49171) );
  AND U40942 ( .A(n21032), .B(n49171), .Z(n60601) );
  NANDN U40943 ( .A(n21033), .B(n60601), .Z(n21034) );
  NAND U40944 ( .A(n21035), .B(n21034), .Z(n21036) );
  NAND U40945 ( .A(n60602), .B(n21036), .Z(n21037) );
  AND U40946 ( .A(n22254), .B(n21037), .Z(n21038) );
  NANDN U40947 ( .A(n60605), .B(n21038), .Z(n21039) );
  NANDN U40948 ( .A(n60606), .B(n21039), .Z(n21040) );
  AND U40949 ( .A(n49182), .B(n21040), .Z(n21041) );
  NANDN U40950 ( .A(x[7663]), .B(y[7663]), .Z(n60607) );
  NAND U40951 ( .A(n21041), .B(n60607), .Z(n21042) );
  AND U40952 ( .A(n60609), .B(n21042), .Z(n21044) );
  XNOR U40953 ( .A(x[7666]), .B(y[7666]), .Z(n22252) );
  ANDN U40954 ( .B(y[7665]), .A(x[7665]), .Z(n50648) );
  ANDN U40955 ( .B(n22252), .A(n50648), .Z(n21043) );
  NANDN U40956 ( .A(n21044), .B(n21043), .Z(n21045) );
  NANDN U40957 ( .A(n50646), .B(n21045), .Z(n21046) );
  AND U40958 ( .A(n49192), .B(n21046), .Z(n21047) );
  NANDN U40959 ( .A(x[7667]), .B(y[7667]), .Z(n50645) );
  NAND U40960 ( .A(n21047), .B(n50645), .Z(n21048) );
  NAND U40961 ( .A(n60610), .B(n21048), .Z(n21049) );
  AND U40962 ( .A(n60611), .B(n21049), .Z(n21050) );
  NANDN U40963 ( .A(y[7670]), .B(x[7670]), .Z(n22248) );
  NANDN U40964 ( .A(y[7671]), .B(x[7671]), .Z(n22245) );
  NAND U40965 ( .A(n22248), .B(n22245), .Z(n60612) );
  OR U40966 ( .A(n21050), .B(n60612), .Z(n21051) );
  NAND U40967 ( .A(n60613), .B(n21051), .Z(n21052) );
  NAND U40968 ( .A(n60614), .B(n21052), .Z(n21053) );
  NAND U40969 ( .A(n60615), .B(n21053), .Z(n21054) );
  AND U40970 ( .A(n60616), .B(n21054), .Z(n21055) );
  NOR U40971 ( .A(n22240), .B(n21055), .Z(n21056) );
  NAND U40972 ( .A(n22239), .B(n21056), .Z(n21057) );
  NANDN U40973 ( .A(n60620), .B(n21057), .Z(n21058) );
  AND U40974 ( .A(n22237), .B(n21058), .Z(n21059) );
  NANDN U40975 ( .A(x[7677]), .B(y[7677]), .Z(n50642) );
  NAND U40976 ( .A(n21059), .B(n50642), .Z(n21060) );
  AND U40977 ( .A(n60621), .B(n21060), .Z(n21062) );
  XNOR U40978 ( .A(x[7680]), .B(y[7680]), .Z(n49220) );
  NANDN U40979 ( .A(x[7679]), .B(y[7679]), .Z(n60622) );
  AND U40980 ( .A(n49220), .B(n60622), .Z(n21061) );
  NANDN U40981 ( .A(n21062), .B(n21061), .Z(n21063) );
  NANDN U40982 ( .A(n60624), .B(n21063), .Z(n21064) );
  AND U40983 ( .A(n22235), .B(n21064), .Z(n21065) );
  ANDN U40984 ( .B(y[7681]), .A(x[7681]), .Z(n50640) );
  ANDN U40985 ( .B(n21065), .A(n50640), .Z(n21067) );
  NANDN U40986 ( .A(y[7682]), .B(x[7682]), .Z(n21066) );
  NANDN U40987 ( .A(y[7683]), .B(x[7683]), .Z(n22232) );
  AND U40988 ( .A(n21066), .B(n22232), .Z(n50639) );
  NANDN U40989 ( .A(n21067), .B(n50639), .Z(n21068) );
  AND U40990 ( .A(n60625), .B(n21068), .Z(n21069) );
  NANDN U40991 ( .A(y[7684]), .B(x[7684]), .Z(n22231) );
  NANDN U40992 ( .A(y[7685]), .B(x[7685]), .Z(n22228) );
  NAND U40993 ( .A(n22231), .B(n22228), .Z(n60626) );
  OR U40994 ( .A(n21069), .B(n60626), .Z(n21070) );
  NAND U40995 ( .A(n21071), .B(n21070), .Z(n21072) );
  NANDN U40996 ( .A(n50636), .B(n21072), .Z(n21073) );
  AND U40997 ( .A(n49238), .B(n21073), .Z(n21074) );
  NANDN U40998 ( .A(x[7687]), .B(y[7687]), .Z(n50634) );
  AND U40999 ( .A(n21074), .B(n50634), .Z(n21076) );
  NANDN U41000 ( .A(y[7688]), .B(x[7688]), .Z(n21075) );
  NANDN U41001 ( .A(y[7689]), .B(x[7689]), .Z(n22226) );
  AND U41002 ( .A(n21075), .B(n22226), .Z(n60628) );
  NANDN U41003 ( .A(n21076), .B(n60628), .Z(n21077) );
  AND U41004 ( .A(n22227), .B(n21077), .Z(n21078) );
  ANDN U41005 ( .B(y[7689]), .A(x[7689]), .Z(n60629) );
  ANDN U41006 ( .B(n21078), .A(n60629), .Z(n21080) );
  NANDN U41007 ( .A(y[7690]), .B(x[7690]), .Z(n21079) );
  NANDN U41008 ( .A(y[7691]), .B(x[7691]), .Z(n49248) );
  NAND U41009 ( .A(n21079), .B(n49248), .Z(n60631) );
  OR U41010 ( .A(n21080), .B(n60631), .Z(n21081) );
  AND U41011 ( .A(n49249), .B(n21081), .Z(n21082) );
  NANDN U41012 ( .A(n60633), .B(n21082), .Z(n21084) );
  NANDN U41013 ( .A(y[7692]), .B(x[7692]), .Z(n21083) );
  NANDN U41014 ( .A(y[7693]), .B(x[7693]), .Z(n22224) );
  AND U41015 ( .A(n21083), .B(n22224), .Z(n50632) );
  AND U41016 ( .A(n21084), .B(n50632), .Z(n21085) );
  OR U41017 ( .A(n21086), .B(n21085), .Z(n21087) );
  NAND U41018 ( .A(n60636), .B(n21087), .Z(n21088) );
  NANDN U41019 ( .A(n21089), .B(n21088), .Z(n21090) );
  NAND U41020 ( .A(n60637), .B(n21090), .Z(n21091) );
  NAND U41021 ( .A(n60638), .B(n21091), .Z(n21092) );
  AND U41022 ( .A(n60639), .B(n21092), .Z(n21093) );
  NOR U41023 ( .A(n22219), .B(n21093), .Z(n21094) );
  NAND U41024 ( .A(n49269), .B(n21094), .Z(n21095) );
  NANDN U41025 ( .A(n60644), .B(n21095), .Z(n21096) );
  AND U41026 ( .A(n22218), .B(n21096), .Z(n21097) );
  NANDN U41027 ( .A(n50628), .B(n21097), .Z(n21099) );
  NANDN U41028 ( .A(y[7702]), .B(x[7702]), .Z(n21098) );
  NANDN U41029 ( .A(y[7703]), .B(x[7703]), .Z(n49278) );
  AND U41030 ( .A(n21098), .B(n49278), .Z(n50627) );
  AND U41031 ( .A(n21099), .B(n50627), .Z(n21101) );
  XNOR U41032 ( .A(x[7704]), .B(y[7704]), .Z(n49279) );
  NANDN U41033 ( .A(x[7703]), .B(y[7703]), .Z(n60645) );
  AND U41034 ( .A(n49279), .B(n60645), .Z(n21100) );
  NANDN U41035 ( .A(n21101), .B(n21100), .Z(n21102) );
  NAND U41036 ( .A(n60647), .B(n21102), .Z(n21103) );
  AND U41037 ( .A(n22216), .B(n21103), .Z(n21104) );
  NANDN U41038 ( .A(n60648), .B(n21104), .Z(n21105) );
  NAND U41039 ( .A(n60650), .B(n21105), .Z(n21106) );
  AND U41040 ( .A(n49289), .B(n21106), .Z(n21107) );
  NANDN U41041 ( .A(x[7707]), .B(y[7707]), .Z(n60651) );
  AND U41042 ( .A(n21107), .B(n60651), .Z(n21109) );
  NANDN U41043 ( .A(y[7708]), .B(x[7708]), .Z(n21108) );
  NANDN U41044 ( .A(y[7709]), .B(x[7709]), .Z(n22213) );
  AND U41045 ( .A(n21108), .B(n22213), .Z(n60653) );
  NANDN U41046 ( .A(n21109), .B(n60653), .Z(n21110) );
  NAND U41047 ( .A(n21111), .B(n21110), .Z(n21112) );
  NAND U41048 ( .A(n60656), .B(n21112), .Z(n21113) );
  AND U41049 ( .A(n49299), .B(n21113), .Z(n21114) );
  NANDN U41050 ( .A(x[7711]), .B(y[7711]), .Z(n50624) );
  AND U41051 ( .A(n21114), .B(n50624), .Z(n21116) );
  NANDN U41052 ( .A(y[7712]), .B(x[7712]), .Z(n21115) );
  NANDN U41053 ( .A(y[7713]), .B(x[7713]), .Z(n22211) );
  AND U41054 ( .A(n21115), .B(n22211), .Z(n60658) );
  NANDN U41055 ( .A(n21116), .B(n60658), .Z(n21117) );
  NAND U41056 ( .A(n21118), .B(n21117), .Z(n21119) );
  NAND U41057 ( .A(n60661), .B(n21119), .Z(n21120) );
  AND U41058 ( .A(n22210), .B(n21120), .Z(n21121) );
  NANDN U41059 ( .A(x[7715]), .B(y[7715]), .Z(n50622) );
  AND U41060 ( .A(n21121), .B(n50622), .Z(n21122) );
  OR U41061 ( .A(n60662), .B(n21122), .Z(n21123) );
  NAND U41062 ( .A(n21124), .B(n21123), .Z(n21125) );
  NAND U41063 ( .A(n60665), .B(n21125), .Z(n21126) );
  AND U41064 ( .A(n49317), .B(n21126), .Z(n21127) );
  NANDN U41065 ( .A(x[7719]), .B(y[7719]), .Z(n60666) );
  AND U41066 ( .A(n21127), .B(n60666), .Z(n21128) );
  OR U41067 ( .A(n60667), .B(n21128), .Z(n21129) );
  NAND U41068 ( .A(n21130), .B(n21129), .Z(n21131) );
  NAND U41069 ( .A(n60670), .B(n21131), .Z(n21132) );
  AND U41070 ( .A(n49327), .B(n21132), .Z(n21133) );
  NANDN U41071 ( .A(x[7723]), .B(y[7723]), .Z(n60671) );
  NAND U41072 ( .A(n21133), .B(n60671), .Z(n21134) );
  NAND U41073 ( .A(n60674), .B(n21134), .Z(n21135) );
  AND U41074 ( .A(n22203), .B(n21135), .Z(n21136) );
  NANDN U41075 ( .A(x[7725]), .B(y[7725]), .Z(n22204) );
  AND U41076 ( .A(n21136), .B(n22204), .Z(n21138) );
  NANDN U41077 ( .A(y[7726]), .B(x[7726]), .Z(n21137) );
  NANDN U41078 ( .A(y[7727]), .B(x[7727]), .Z(n22200) );
  AND U41079 ( .A(n21137), .B(n22200), .Z(n60679) );
  NANDN U41080 ( .A(n21138), .B(n60679), .Z(n21139) );
  NAND U41081 ( .A(n21140), .B(n21139), .Z(n21141) );
  NAND U41082 ( .A(n60684), .B(n21141), .Z(n21142) );
  AND U41083 ( .A(n22199), .B(n21142), .Z(n21143) );
  NANDN U41084 ( .A(x[7729]), .B(y[7729]), .Z(n50617) );
  AND U41085 ( .A(n21143), .B(n50617), .Z(n21145) );
  NANDN U41086 ( .A(y[7730]), .B(x[7730]), .Z(n21144) );
  NANDN U41087 ( .A(y[7731]), .B(x[7731]), .Z(n49344) );
  NAND U41088 ( .A(n21144), .B(n49344), .Z(n60689) );
  OR U41089 ( .A(n21145), .B(n60689), .Z(n21146) );
  NAND U41090 ( .A(n21147), .B(n21146), .Z(n21148) );
  AND U41091 ( .A(n60695), .B(n21148), .Z(n21150) );
  XNOR U41092 ( .A(x[7734]), .B(y[7734]), .Z(n22197) );
  ANDN U41093 ( .B(y[7733]), .A(x[7733]), .Z(n60696) );
  ANDN U41094 ( .B(n22197), .A(n60696), .Z(n21149) );
  NANDN U41095 ( .A(n21150), .B(n21149), .Z(n21151) );
  NAND U41096 ( .A(n60701), .B(n21151), .Z(n21152) );
  AND U41097 ( .A(n49355), .B(n21152), .Z(n21153) );
  NAND U41098 ( .A(n60703), .B(n21153), .Z(n21154) );
  NAND U41099 ( .A(n60707), .B(n21154), .Z(n21155) );
  AND U41100 ( .A(n22195), .B(n21155), .Z(n21156) );
  NANDN U41101 ( .A(n60708), .B(n21156), .Z(n21157) );
  AND U41102 ( .A(n60711), .B(n21157), .Z(n21159) );
  XNOR U41103 ( .A(x[7740]), .B(y[7740]), .Z(n49365) );
  NANDN U41104 ( .A(x[7739]), .B(y[7739]), .Z(n50615) );
  AND U41105 ( .A(n49365), .B(n50615), .Z(n21158) );
  NANDN U41106 ( .A(n21159), .B(n21158), .Z(n21160) );
  NAND U41107 ( .A(n60712), .B(n21160), .Z(n21161) );
  AND U41108 ( .A(n22193), .B(n21161), .Z(n21162) );
  NANDN U41109 ( .A(n60713), .B(n21162), .Z(n21164) );
  NANDN U41110 ( .A(y[7742]), .B(x[7742]), .Z(n21163) );
  NANDN U41111 ( .A(y[7743]), .B(x[7743]), .Z(n49374) );
  AND U41112 ( .A(n21163), .B(n49374), .Z(n60715) );
  AND U41113 ( .A(n21164), .B(n60715), .Z(n21165) );
  OR U41114 ( .A(n21166), .B(n21165), .Z(n21167) );
  NAND U41115 ( .A(n50612), .B(n21167), .Z(n21168) );
  NANDN U41116 ( .A(n21169), .B(n21168), .Z(n21170) );
  NAND U41117 ( .A(n60718), .B(n21170), .Z(n21171) );
  AND U41118 ( .A(n49385), .B(n21171), .Z(n21172) );
  NANDN U41119 ( .A(x[7747]), .B(y[7747]), .Z(n60719) );
  AND U41120 ( .A(n21172), .B(n60719), .Z(n21173) );
  OR U41121 ( .A(n60721), .B(n21173), .Z(n21174) );
  NAND U41122 ( .A(n21175), .B(n21174), .Z(n21176) );
  NAND U41123 ( .A(n60724), .B(n21176), .Z(n21177) );
  AND U41124 ( .A(n49395), .B(n21177), .Z(n21178) );
  NANDN U41125 ( .A(x[7751]), .B(y[7751]), .Z(n60725) );
  NAND U41126 ( .A(n21178), .B(n60725), .Z(n21179) );
  AND U41127 ( .A(n60727), .B(n21179), .Z(n21181) );
  XNOR U41128 ( .A(x[7754]), .B(y[7754]), .Z(n22186) );
  NANDN U41129 ( .A(x[7753]), .B(y[7753]), .Z(n22187) );
  AND U41130 ( .A(n22186), .B(n22187), .Z(n21180) );
  NANDN U41131 ( .A(n21181), .B(n21180), .Z(n21182) );
  NAND U41132 ( .A(n60728), .B(n21182), .Z(n21183) );
  AND U41133 ( .A(n49405), .B(n21183), .Z(n21184) );
  NANDN U41134 ( .A(x[7755]), .B(y[7755]), .Z(n60729) );
  NAND U41135 ( .A(n21184), .B(n60729), .Z(n21185) );
  NAND U41136 ( .A(n60731), .B(n21185), .Z(n21186) );
  AND U41137 ( .A(n22184), .B(n21186), .Z(n21187) );
  ANDN U41138 ( .B(y[7757]), .A(x[7757]), .Z(n50607) );
  ANDN U41139 ( .B(n21187), .A(n50607), .Z(n21189) );
  NANDN U41140 ( .A(y[7758]), .B(x[7758]), .Z(n21188) );
  NANDN U41141 ( .A(y[7759]), .B(x[7759]), .Z(n49415) );
  AND U41142 ( .A(n21188), .B(n49415), .Z(n50606) );
  NANDN U41143 ( .A(n21189), .B(n50606), .Z(n21190) );
  NAND U41144 ( .A(n21191), .B(n21190), .Z(n21192) );
  NAND U41145 ( .A(n60735), .B(n21192), .Z(n21193) );
  AND U41146 ( .A(n22182), .B(n21193), .Z(n21194) );
  ANDN U41147 ( .B(y[7761]), .A(x[7761]), .Z(n60736) );
  ANDN U41148 ( .B(n21194), .A(n60736), .Z(n21196) );
  NANDN U41149 ( .A(y[7762]), .B(x[7762]), .Z(n21195) );
  NANDN U41150 ( .A(y[7763]), .B(x[7763]), .Z(n49425) );
  NAND U41151 ( .A(n21195), .B(n49425), .Z(n60738) );
  OR U41152 ( .A(n21196), .B(n60738), .Z(n21197) );
  NAND U41153 ( .A(n21198), .B(n21197), .Z(n21199) );
  NAND U41154 ( .A(n60741), .B(n21199), .Z(n21200) );
  AND U41155 ( .A(n60742), .B(n21200), .Z(n21201) );
  NANDN U41156 ( .A(y[7766]), .B(x[7766]), .Z(n22178) );
  NANDN U41157 ( .A(y[7767]), .B(x[7767]), .Z(n22174) );
  AND U41158 ( .A(n22178), .B(n22174), .Z(n60743) );
  NANDN U41159 ( .A(n21201), .B(n60743), .Z(n21202) );
  NAND U41160 ( .A(n21203), .B(n21202), .Z(n21204) );
  NAND U41161 ( .A(n60744), .B(n21204), .Z(n21205) );
  NAND U41162 ( .A(n60745), .B(n21205), .Z(n21206) );
  NANDN U41163 ( .A(y[7770]), .B(x[7770]), .Z(n22172) );
  NANDN U41164 ( .A(y[7771]), .B(x[7771]), .Z(n22169) );
  AND U41165 ( .A(n22172), .B(n22169), .Z(n60746) );
  AND U41166 ( .A(n21206), .B(n60746), .Z(n21207) );
  ANDN U41167 ( .B(y[7772]), .A(x[7772]), .Z(n49447) );
  NANDN U41168 ( .A(x[7771]), .B(y[7771]), .Z(n22170) );
  NANDN U41169 ( .A(n49447), .B(n22170), .Z(n50603) );
  OR U41170 ( .A(n21207), .B(n50603), .Z(n21208) );
  NAND U41171 ( .A(n50602), .B(n21208), .Z(n21209) );
  NANDN U41172 ( .A(n21210), .B(n21209), .Z(n21211) );
  NAND U41173 ( .A(n60750), .B(n21211), .Z(n21212) );
  AND U41174 ( .A(n49454), .B(n21212), .Z(n21213) );
  NANDN U41175 ( .A(x[7775]), .B(y[7775]), .Z(n60751) );
  AND U41176 ( .A(n21213), .B(n60751), .Z(n21215) );
  NANDN U41177 ( .A(y[7776]), .B(x[7776]), .Z(n21214) );
  NANDN U41178 ( .A(y[7777]), .B(x[7777]), .Z(n22163) );
  NAND U41179 ( .A(n21214), .B(n22163), .Z(n60753) );
  OR U41180 ( .A(n21215), .B(n60753), .Z(n21216) );
  NAND U41181 ( .A(n21217), .B(n21216), .Z(n21218) );
  NAND U41182 ( .A(n60754), .B(n21218), .Z(n21219) );
  AND U41183 ( .A(n49464), .B(n21219), .Z(n21220) );
  NANDN U41184 ( .A(x[7779]), .B(y[7779]), .Z(n60755) );
  NAND U41185 ( .A(n21220), .B(n60755), .Z(n21222) );
  NANDN U41186 ( .A(y[7780]), .B(x[7780]), .Z(n21221) );
  NANDN U41187 ( .A(y[7781]), .B(x[7781]), .Z(n22161) );
  AND U41188 ( .A(n21221), .B(n22161), .Z(n60757) );
  AND U41189 ( .A(n21222), .B(n60757), .Z(n21224) );
  XNOR U41190 ( .A(x[7782]), .B(y[7782]), .Z(n22162) );
  ANDN U41191 ( .B(y[7781]), .A(x[7781]), .Z(n50598) );
  ANDN U41192 ( .B(n22162), .A(n50598), .Z(n21223) );
  NANDN U41193 ( .A(n21224), .B(n21223), .Z(n21225) );
  NANDN U41194 ( .A(n60758), .B(n21225), .Z(n21226) );
  AND U41195 ( .A(n49474), .B(n21226), .Z(n21227) );
  NANDN U41196 ( .A(x[7783]), .B(y[7783]), .Z(n60760) );
  NAND U41197 ( .A(n21227), .B(n60760), .Z(n21228) );
  NAND U41198 ( .A(n60762), .B(n21228), .Z(n21229) );
  AND U41199 ( .A(n22160), .B(n21229), .Z(n21230) );
  ANDN U41200 ( .B(y[7785]), .A(x[7785]), .Z(n50596) );
  ANDN U41201 ( .B(n21230), .A(n50596), .Z(n21232) );
  NANDN U41202 ( .A(y[7786]), .B(x[7786]), .Z(n21231) );
  NANDN U41203 ( .A(y[7787]), .B(x[7787]), .Z(n49484) );
  AND U41204 ( .A(n21231), .B(n49484), .Z(n60763) );
  NANDN U41205 ( .A(n21232), .B(n60763), .Z(n21233) );
  NAND U41206 ( .A(n21234), .B(n21233), .Z(n21235) );
  AND U41207 ( .A(n60764), .B(n21235), .Z(n21236) );
  NOR U41208 ( .A(n60765), .B(n21236), .Z(n21237) );
  NAND U41209 ( .A(n22158), .B(n21237), .Z(n21238) );
  NANDN U41210 ( .A(n60767), .B(n21238), .Z(n21239) );
  AND U41211 ( .A(n49495), .B(n21239), .Z(n21240) );
  NANDN U41212 ( .A(x[7791]), .B(y[7791]), .Z(n50593) );
  NAND U41213 ( .A(n21240), .B(n50593), .Z(n21241) );
  NANDN U41214 ( .A(n60768), .B(n21241), .Z(n21242) );
  AND U41215 ( .A(n22156), .B(n21242), .Z(n21243) );
  NANDN U41216 ( .A(n60769), .B(n21243), .Z(n21244) );
  NAND U41217 ( .A(n60772), .B(n21244), .Z(n21245) );
  AND U41218 ( .A(n49505), .B(n21245), .Z(n21246) );
  NANDN U41219 ( .A(x[7795]), .B(y[7795]), .Z(n60773) );
  AND U41220 ( .A(n21246), .B(n60773), .Z(n21248) );
  NANDN U41221 ( .A(y[7796]), .B(x[7796]), .Z(n21247) );
  NANDN U41222 ( .A(y[7797]), .B(x[7797]), .Z(n22153) );
  AND U41223 ( .A(n21247), .B(n22153), .Z(n50591) );
  NANDN U41224 ( .A(n21248), .B(n50591), .Z(n21249) );
  NAND U41225 ( .A(n21250), .B(n21249), .Z(n21251) );
  NAND U41226 ( .A(n60777), .B(n21251), .Z(n21252) );
  AND U41227 ( .A(n49515), .B(n21252), .Z(n21253) );
  NANDN U41228 ( .A(x[7799]), .B(y[7799]), .Z(n50590) );
  AND U41229 ( .A(n21253), .B(n50590), .Z(n21255) );
  NANDN U41230 ( .A(y[7800]), .B(x[7800]), .Z(n21254) );
  NANDN U41231 ( .A(y[7801]), .B(x[7801]), .Z(n22151) );
  NAND U41232 ( .A(n21254), .B(n22151), .Z(n50588) );
  OR U41233 ( .A(n21255), .B(n50588), .Z(n21256) );
  NAND U41234 ( .A(n21257), .B(n21256), .Z(n21258) );
  NAND U41235 ( .A(n60778), .B(n21258), .Z(n21259) );
  AND U41236 ( .A(n49525), .B(n21259), .Z(n21260) );
  NANDN U41237 ( .A(x[7803]), .B(y[7803]), .Z(n60779) );
  AND U41238 ( .A(n21260), .B(n60779), .Z(n21262) );
  NANDN U41239 ( .A(y[7804]), .B(x[7804]), .Z(n21261) );
  NANDN U41240 ( .A(y[7805]), .B(x[7805]), .Z(n22149) );
  NAND U41241 ( .A(n21261), .B(n22149), .Z(n60781) );
  OR U41242 ( .A(n21262), .B(n60781), .Z(n21263) );
  NAND U41243 ( .A(n21264), .B(n21263), .Z(n21265) );
  NANDN U41244 ( .A(n60789), .B(n21265), .Z(n21266) );
  AND U41245 ( .A(n49535), .B(n21266), .Z(n21267) );
  NANDN U41246 ( .A(x[7807]), .B(y[7807]), .Z(n60791) );
  NAND U41247 ( .A(n21267), .B(n60791), .Z(n21268) );
  AND U41248 ( .A(n60795), .B(n21268), .Z(n21270) );
  XNOR U41249 ( .A(x[7810]), .B(y[7810]), .Z(n22148) );
  ANDN U41250 ( .B(y[7809]), .A(x[7809]), .Z(n60796) );
  ANDN U41251 ( .B(n22148), .A(n60796), .Z(n21269) );
  NANDN U41252 ( .A(n21270), .B(n21269), .Z(n21271) );
  NANDN U41253 ( .A(n60801), .B(n21271), .Z(n21272) );
  AND U41254 ( .A(n49545), .B(n21272), .Z(n21273) );
  NANDN U41255 ( .A(x[7811]), .B(y[7811]), .Z(n60803) );
  NAND U41256 ( .A(n21273), .B(n60803), .Z(n21274) );
  AND U41257 ( .A(n60807), .B(n21274), .Z(n21275) );
  ANDN U41258 ( .B(n22146), .A(n21275), .Z(n21276) );
  ANDN U41259 ( .B(y[7813]), .A(x[7813]), .Z(n60808) );
  ANDN U41260 ( .B(n21276), .A(n60808), .Z(n21278) );
  NANDN U41261 ( .A(y[7814]), .B(x[7814]), .Z(n21277) );
  NANDN U41262 ( .A(y[7815]), .B(x[7815]), .Z(n22143) );
  AND U41263 ( .A(n21277), .B(n22143), .Z(n60812) );
  NANDN U41264 ( .A(n21278), .B(n60812), .Z(n21279) );
  NAND U41265 ( .A(n21280), .B(n21279), .Z(n21281) );
  NAND U41266 ( .A(n60817), .B(n21281), .Z(n21282) );
  AND U41267 ( .A(n22142), .B(n21282), .Z(n21283) );
  NANDN U41268 ( .A(x[7817]), .B(y[7817]), .Z(n60819) );
  AND U41269 ( .A(n21283), .B(n60819), .Z(n21284) );
  OR U41270 ( .A(n60823), .B(n21284), .Z(n21285) );
  NAND U41271 ( .A(n21286), .B(n21285), .Z(n21287) );
  NANDN U41272 ( .A(n60824), .B(n21287), .Z(n21288) );
  AND U41273 ( .A(n22140), .B(n21288), .Z(n21289) );
  ANDN U41274 ( .B(y[7821]), .A(x[7821]), .Z(n60825) );
  ANDN U41275 ( .B(n21289), .A(n60825), .Z(n21291) );
  NANDN U41276 ( .A(y[7822]), .B(x[7822]), .Z(n21290) );
  NANDN U41277 ( .A(y[7823]), .B(x[7823]), .Z(n49572) );
  AND U41278 ( .A(n21290), .B(n49572), .Z(n60827) );
  NANDN U41279 ( .A(n21291), .B(n60827), .Z(n21292) );
  NAND U41280 ( .A(n21293), .B(n21292), .Z(n21294) );
  NANDN U41281 ( .A(n60829), .B(n21294), .Z(n21295) );
  AND U41282 ( .A(n22138), .B(n21295), .Z(n21296) );
  NANDN U41283 ( .A(n60830), .B(n21296), .Z(n21297) );
  NAND U41284 ( .A(n60832), .B(n21297), .Z(n21298) );
  AND U41285 ( .A(n49583), .B(n21298), .Z(n21299) );
  NANDN U41286 ( .A(x[7827]), .B(y[7827]), .Z(n60833) );
  AND U41287 ( .A(n21299), .B(n60833), .Z(n21301) );
  NANDN U41288 ( .A(y[7828]), .B(x[7828]), .Z(n21300) );
  NANDN U41289 ( .A(y[7829]), .B(x[7829]), .Z(n22134) );
  NAND U41290 ( .A(n21300), .B(n22134), .Z(n60835) );
  OR U41291 ( .A(n21301), .B(n60835), .Z(n21302) );
  NAND U41292 ( .A(n21303), .B(n21302), .Z(n21304) );
  NAND U41293 ( .A(n60837), .B(n21304), .Z(n21305) );
  AND U41294 ( .A(n49593), .B(n21305), .Z(n21306) );
  NANDN U41295 ( .A(x[7831]), .B(y[7831]), .Z(n60840) );
  AND U41296 ( .A(n21306), .B(n60840), .Z(n21308) );
  NANDN U41297 ( .A(y[7832]), .B(x[7832]), .Z(n21307) );
  NANDN U41298 ( .A(y[7833]), .B(x[7833]), .Z(n22132) );
  NAND U41299 ( .A(n21307), .B(n22132), .Z(n60841) );
  OR U41300 ( .A(n21308), .B(n60841), .Z(n21309) );
  AND U41301 ( .A(n21310), .B(n21309), .Z(n21311) );
  OR U41302 ( .A(n60842), .B(n21311), .Z(n21312) );
  NAND U41303 ( .A(n21313), .B(n21312), .Z(n21314) );
  AND U41304 ( .A(n60845), .B(n21314), .Z(n21316) );
  XNOR U41305 ( .A(x[7838]), .B(y[7838]), .Z(n22129) );
  NANDN U41306 ( .A(x[7837]), .B(y[7837]), .Z(n60846) );
  AND U41307 ( .A(n22129), .B(n60846), .Z(n21315) );
  NANDN U41308 ( .A(n21316), .B(n21315), .Z(n21317) );
  NANDN U41309 ( .A(n60848), .B(n21317), .Z(n21318) );
  AND U41310 ( .A(n49612), .B(n21318), .Z(n21319) );
  NANDN U41311 ( .A(n50575), .B(n21319), .Z(n21320) );
  NAND U41312 ( .A(n60849), .B(n21320), .Z(n21321) );
  AND U41313 ( .A(n22127), .B(n21321), .Z(n21322) );
  ANDN U41314 ( .B(y[7841]), .A(x[7841]), .Z(n60850) );
  ANDN U41315 ( .B(n21322), .A(n60850), .Z(n21324) );
  NANDN U41316 ( .A(y[7842]), .B(x[7842]), .Z(n21323) );
  NANDN U41317 ( .A(y[7843]), .B(x[7843]), .Z(n22124) );
  AND U41318 ( .A(n21323), .B(n22124), .Z(n60852) );
  NANDN U41319 ( .A(n21324), .B(n60852), .Z(n21325) );
  NAND U41320 ( .A(n21326), .B(n21325), .Z(n21327) );
  NAND U41321 ( .A(n60855), .B(n21327), .Z(n21328) );
  AND U41322 ( .A(n22123), .B(n21328), .Z(n21329) );
  ANDN U41323 ( .B(y[7845]), .A(x[7845]), .Z(n60856) );
  ANDN U41324 ( .B(n21329), .A(n60856), .Z(n21331) );
  NANDN U41325 ( .A(y[7846]), .B(x[7846]), .Z(n21330) );
  NANDN U41326 ( .A(y[7847]), .B(x[7847]), .Z(n49630) );
  AND U41327 ( .A(n21330), .B(n49630), .Z(n60858) );
  NANDN U41328 ( .A(n21331), .B(n60858), .Z(n21332) );
  NAND U41329 ( .A(n21333), .B(n21332), .Z(n21334) );
  NAND U41330 ( .A(n60860), .B(n21334), .Z(n21335) );
  AND U41331 ( .A(n22121), .B(n21335), .Z(n21336) );
  ANDN U41332 ( .B(y[7849]), .A(x[7849]), .Z(n60861) );
  ANDN U41333 ( .B(n21336), .A(n60861), .Z(n21338) );
  NANDN U41334 ( .A(y[7850]), .B(x[7850]), .Z(n21337) );
  NANDN U41335 ( .A(y[7851]), .B(x[7851]), .Z(n49640) );
  AND U41336 ( .A(n21337), .B(n49640), .Z(n60863) );
  NANDN U41337 ( .A(n21338), .B(n60863), .Z(n21339) );
  NAND U41338 ( .A(n21340), .B(n21339), .Z(n21341) );
  NANDN U41339 ( .A(n60866), .B(n21341), .Z(n21342) );
  AND U41340 ( .A(n22119), .B(n21342), .Z(n21343) );
  NANDN U41341 ( .A(n50569), .B(n21343), .Z(n21345) );
  NANDN U41342 ( .A(y[7854]), .B(x[7854]), .Z(n21344) );
  NANDN U41343 ( .A(y[7855]), .B(x[7855]), .Z(n49650) );
  AND U41344 ( .A(n21344), .B(n49650), .Z(n60867) );
  AND U41345 ( .A(n21345), .B(n60867), .Z(n21347) );
  XNOR U41346 ( .A(x[7856]), .B(y[7856]), .Z(n49651) );
  NANDN U41347 ( .A(x[7855]), .B(y[7855]), .Z(n60870) );
  AND U41348 ( .A(n49651), .B(n60870), .Z(n21346) );
  NANDN U41349 ( .A(n21347), .B(n21346), .Z(n21348) );
  NANDN U41350 ( .A(n60872), .B(n21348), .Z(n21349) );
  AND U41351 ( .A(n22117), .B(n21349), .Z(n21350) );
  NANDN U41352 ( .A(n60874), .B(n21350), .Z(n21351) );
  NAND U41353 ( .A(n60875), .B(n21351), .Z(n21352) );
  NAND U41354 ( .A(n22115), .B(n21352), .Z(n21353) );
  NANDN U41355 ( .A(x[7859]), .B(y[7859]), .Z(n60877) );
  NANDN U41356 ( .A(n21353), .B(n60877), .Z(n21354) );
  NAND U41357 ( .A(n50568), .B(n21354), .Z(n21355) );
  NANDN U41358 ( .A(n60878), .B(n21355), .Z(n21356) );
  NAND U41359 ( .A(n60879), .B(n21356), .Z(n21357) );
  XOR U41360 ( .A(x[7864]), .B(y[7864]), .Z(n49669) );
  ANDN U41361 ( .B(n21357), .A(n49669), .Z(n21358) );
  NANDN U41362 ( .A(x[7863]), .B(y[7863]), .Z(n50566) );
  AND U41363 ( .A(n21358), .B(n50566), .Z(n21359) );
  OR U41364 ( .A(n60880), .B(n21359), .Z(n21360) );
  NAND U41365 ( .A(n60881), .B(n21360), .Z(n21361) );
  NANDN U41366 ( .A(n60882), .B(n21361), .Z(n21362) );
  NAND U41367 ( .A(n60885), .B(n21362), .Z(n21363) );
  NAND U41368 ( .A(n60886), .B(n21363), .Z(n21364) );
  AND U41369 ( .A(n22100), .B(n21364), .Z(n21365) );
  NANDN U41370 ( .A(n22101), .B(n21365), .Z(n21366) );
  NAND U41371 ( .A(n60887), .B(n21366), .Z(n21367) );
  NANDN U41372 ( .A(n50563), .B(n21367), .Z(n21368) );
  NAND U41373 ( .A(n60888), .B(n21368), .Z(n21369) );
  AND U41374 ( .A(n22095), .B(n21369), .Z(n21370) );
  NANDN U41375 ( .A(x[7873]), .B(y[7873]), .Z(n60889) );
  AND U41376 ( .A(n21370), .B(n60889), .Z(n21371) );
  OR U41377 ( .A(n60891), .B(n21371), .Z(n21372) );
  NAND U41378 ( .A(n60892), .B(n21372), .Z(n21373) );
  NAND U41379 ( .A(n60893), .B(n21373), .Z(n21374) );
  AND U41380 ( .A(n22090), .B(n21374), .Z(n21375) );
  NANDN U41381 ( .A(x[7877]), .B(y[7877]), .Z(n60894) );
  NAND U41382 ( .A(n21375), .B(n60894), .Z(n21377) );
  NANDN U41383 ( .A(y[7878]), .B(x[7878]), .Z(n21376) );
  NANDN U41384 ( .A(y[7879]), .B(x[7879]), .Z(n22087) );
  AND U41385 ( .A(n21376), .B(n22087), .Z(n60896) );
  AND U41386 ( .A(n21377), .B(n60896), .Z(n21378) );
  NANDN U41387 ( .A(x[7879]), .B(y[7879]), .Z(n22088) );
  NANDN U41388 ( .A(x[7880]), .B(y[7880]), .Z(n22085) );
  NAND U41389 ( .A(n22088), .B(n22085), .Z(n50562) );
  OR U41390 ( .A(n21378), .B(n50562), .Z(n21379) );
  NAND U41391 ( .A(n50561), .B(n21379), .Z(n21380) );
  NAND U41392 ( .A(n60899), .B(n21380), .Z(n21381) );
  NAND U41393 ( .A(n60900), .B(n21381), .Z(n21382) );
  AND U41394 ( .A(n49713), .B(n21382), .Z(n21383) );
  NANDN U41395 ( .A(x[7883]), .B(y[7883]), .Z(n60901) );
  NAND U41396 ( .A(n21383), .B(n60901), .Z(n21384) );
  AND U41397 ( .A(n60903), .B(n21384), .Z(n21385) );
  NOR U41398 ( .A(n50560), .B(n21385), .Z(n21386) );
  NAND U41399 ( .A(n22080), .B(n21386), .Z(n21387) );
  NAND U41400 ( .A(n60904), .B(n21387), .Z(n21388) );
  AND U41401 ( .A(n49723), .B(n21388), .Z(n21389) );
  NANDN U41402 ( .A(x[7887]), .B(y[7887]), .Z(n60905) );
  NAND U41403 ( .A(n21389), .B(n60905), .Z(n21390) );
  NAND U41404 ( .A(n60907), .B(n21390), .Z(n21391) );
  AND U41405 ( .A(n22078), .B(n21391), .Z(n21392) );
  NANDN U41406 ( .A(n50557), .B(n21392), .Z(n21393) );
  NANDN U41407 ( .A(n60908), .B(n21393), .Z(n21394) );
  AND U41408 ( .A(n22076), .B(n21394), .Z(n21395) );
  NANDN U41409 ( .A(x[7891]), .B(y[7891]), .Z(n60910) );
  NAND U41410 ( .A(n21395), .B(n60910), .Z(n21396) );
  AND U41411 ( .A(n60912), .B(n21396), .Z(n21397) );
  ANDN U41412 ( .B(n22074), .A(n21397), .Z(n21398) );
  NANDN U41413 ( .A(x[7893]), .B(y[7893]), .Z(n60913) );
  AND U41414 ( .A(n21398), .B(n60913), .Z(n21400) );
  NANDN U41415 ( .A(y[7894]), .B(x[7894]), .Z(n21399) );
  NANDN U41416 ( .A(y[7895]), .B(x[7895]), .Z(n49741) );
  AND U41417 ( .A(n21399), .B(n49741), .Z(n50556) );
  NANDN U41418 ( .A(n21400), .B(n50556), .Z(n21401) );
  NAND U41419 ( .A(n21402), .B(n21401), .Z(n21403) );
  NAND U41420 ( .A(n60917), .B(n21403), .Z(n21404) );
  AND U41421 ( .A(n22072), .B(n21404), .Z(n21405) );
  ANDN U41422 ( .B(y[7897]), .A(x[7897]), .Z(n60918) );
  ANDN U41423 ( .B(n21405), .A(n60918), .Z(n21407) );
  NANDN U41424 ( .A(y[7898]), .B(x[7898]), .Z(n21406) );
  NANDN U41425 ( .A(y[7899]), .B(x[7899]), .Z(n49751) );
  NAND U41426 ( .A(n21406), .B(n49751), .Z(n60920) );
  OR U41427 ( .A(n21407), .B(n60920), .Z(n21408) );
  NAND U41428 ( .A(n21409), .B(n21408), .Z(n21410) );
  NAND U41429 ( .A(n60921), .B(n21410), .Z(n21411) );
  AND U41430 ( .A(n22070), .B(n21411), .Z(n21412) );
  NANDN U41431 ( .A(n60922), .B(n21412), .Z(n21414) );
  NANDN U41432 ( .A(y[7902]), .B(x[7902]), .Z(n21413) );
  NANDN U41433 ( .A(y[7903]), .B(x[7903]), .Z(n49761) );
  AND U41434 ( .A(n21413), .B(n49761), .Z(n60924) );
  AND U41435 ( .A(n21414), .B(n60924), .Z(n21416) );
  XNOR U41436 ( .A(x[7904]), .B(y[7904]), .Z(n49762) );
  NANDN U41437 ( .A(x[7903]), .B(y[7903]), .Z(n50553) );
  AND U41438 ( .A(n49762), .B(n50553), .Z(n21415) );
  NANDN U41439 ( .A(n21416), .B(n21415), .Z(n21417) );
  NANDN U41440 ( .A(n60927), .B(n21417), .Z(n21418) );
  AND U41441 ( .A(n22068), .B(n21418), .Z(n21419) );
  NANDN U41442 ( .A(n60928), .B(n21419), .Z(n21420) );
  AND U41443 ( .A(n60930), .B(n21420), .Z(n21421) );
  OR U41444 ( .A(n21422), .B(n21421), .Z(n21423) );
  NAND U41445 ( .A(n50550), .B(n21423), .Z(n21424) );
  NANDN U41446 ( .A(n21425), .B(n21424), .Z(n21426) );
  NAND U41447 ( .A(n60934), .B(n21426), .Z(n21427) );
  AND U41448 ( .A(n49782), .B(n21427), .Z(n21428) );
  NANDN U41449 ( .A(x[7911]), .B(y[7911]), .Z(n60935) );
  AND U41450 ( .A(n21428), .B(n60935), .Z(n21430) );
  NANDN U41451 ( .A(y[7912]), .B(x[7912]), .Z(n21429) );
  NANDN U41452 ( .A(y[7913]), .B(x[7913]), .Z(n22062) );
  NAND U41453 ( .A(n21429), .B(n22062), .Z(n60937) );
  OR U41454 ( .A(n21430), .B(n60937), .Z(n21431) );
  NAND U41455 ( .A(n21432), .B(n21431), .Z(n21433) );
  NAND U41456 ( .A(n60940), .B(n21433), .Z(n21434) );
  AND U41457 ( .A(n49792), .B(n21434), .Z(n21435) );
  NANDN U41458 ( .A(x[7915]), .B(y[7915]), .Z(n60941) );
  NAND U41459 ( .A(n21435), .B(n60941), .Z(n21437) );
  NANDN U41460 ( .A(y[7916]), .B(x[7916]), .Z(n21436) );
  NANDN U41461 ( .A(y[7917]), .B(x[7917]), .Z(n22060) );
  AND U41462 ( .A(n21436), .B(n22060), .Z(n60943) );
  AND U41463 ( .A(n21437), .B(n60943), .Z(n21439) );
  XNOR U41464 ( .A(x[7918]), .B(y[7918]), .Z(n22061) );
  ANDN U41465 ( .B(y[7917]), .A(x[7917]), .Z(n50546) );
  ANDN U41466 ( .B(n22061), .A(n50546), .Z(n21438) );
  NANDN U41467 ( .A(n21439), .B(n21438), .Z(n21440) );
  NANDN U41468 ( .A(n60944), .B(n21440), .Z(n21441) );
  AND U41469 ( .A(n49802), .B(n21441), .Z(n21442) );
  NANDN U41470 ( .A(x[7919]), .B(y[7919]), .Z(n60945) );
  NAND U41471 ( .A(n21442), .B(n60945), .Z(n21443) );
  NAND U41472 ( .A(n60947), .B(n21443), .Z(n21444) );
  AND U41473 ( .A(n22059), .B(n21444), .Z(n21445) );
  ANDN U41474 ( .B(y[7921]), .A(x[7921]), .Z(n60948) );
  ANDN U41475 ( .B(n21445), .A(n60948), .Z(n21447) );
  NANDN U41476 ( .A(y[7922]), .B(x[7922]), .Z(n21446) );
  NANDN U41477 ( .A(y[7923]), .B(x[7923]), .Z(n49812) );
  AND U41478 ( .A(n21446), .B(n49812), .Z(n50545) );
  NANDN U41479 ( .A(n21447), .B(n50545), .Z(n21448) );
  NAND U41480 ( .A(n21449), .B(n21448), .Z(n21450) );
  AND U41481 ( .A(n60952), .B(n21450), .Z(n21452) );
  XNOR U41482 ( .A(x[7926]), .B(y[7926]), .Z(n22057) );
  ANDN U41483 ( .B(y[7925]), .A(x[7925]), .Z(n60953) );
  ANDN U41484 ( .B(n22057), .A(n60953), .Z(n21451) );
  NANDN U41485 ( .A(n21452), .B(n21451), .Z(n21453) );
  NANDN U41486 ( .A(n60956), .B(n21453), .Z(n21454) );
  AND U41487 ( .A(n49823), .B(n21454), .Z(n21455) );
  NAND U41488 ( .A(n50543), .B(n21455), .Z(n21456) );
  NAND U41489 ( .A(n60957), .B(n21456), .Z(n21457) );
  AND U41490 ( .A(n22055), .B(n21457), .Z(n21458) );
  NANDN U41491 ( .A(n60958), .B(n21458), .Z(n21460) );
  NANDN U41492 ( .A(y[7930]), .B(x[7930]), .Z(n21459) );
  NANDN U41493 ( .A(y[7931]), .B(x[7931]), .Z(n49832) );
  AND U41494 ( .A(n21459), .B(n49832), .Z(n60960) );
  AND U41495 ( .A(n21460), .B(n60960), .Z(n21461) );
  OR U41496 ( .A(n21462), .B(n21461), .Z(n21463) );
  NAND U41497 ( .A(n50540), .B(n21463), .Z(n21464) );
  NANDN U41498 ( .A(n21465), .B(n21464), .Z(n21466) );
  NAND U41499 ( .A(n60963), .B(n21466), .Z(n21467) );
  AND U41500 ( .A(n49843), .B(n21467), .Z(n21468) );
  NANDN U41501 ( .A(x[7935]), .B(y[7935]), .Z(n60965) );
  AND U41502 ( .A(n21468), .B(n60965), .Z(n21469) );
  OR U41503 ( .A(n60966), .B(n21469), .Z(n21470) );
  NAND U41504 ( .A(n21471), .B(n21470), .Z(n21472) );
  NAND U41505 ( .A(n60969), .B(n21472), .Z(n21473) );
  AND U41506 ( .A(n49853), .B(n21473), .Z(n21474) );
  NANDN U41507 ( .A(x[7939]), .B(y[7939]), .Z(n60970) );
  NAND U41508 ( .A(n21474), .B(n60970), .Z(n21475) );
  AND U41509 ( .A(n60972), .B(n21475), .Z(n21477) );
  XNOR U41510 ( .A(x[7942]), .B(y[7942]), .Z(n22048) );
  NANDN U41511 ( .A(x[7941]), .B(y[7941]), .Z(n22049) );
  AND U41512 ( .A(n22048), .B(n22049), .Z(n21476) );
  NANDN U41513 ( .A(n21477), .B(n21476), .Z(n21478) );
  NAND U41514 ( .A(n60973), .B(n21478), .Z(n21479) );
  AND U41515 ( .A(n22046), .B(n21479), .Z(n21480) );
  NANDN U41516 ( .A(x[7943]), .B(y[7943]), .Z(n60974) );
  NAND U41517 ( .A(n21480), .B(n60974), .Z(n21481) );
  NAND U41518 ( .A(n60976), .B(n21481), .Z(n21482) );
  AND U41519 ( .A(n22044), .B(n21482), .Z(n21483) );
  NANDN U41520 ( .A(x[7945]), .B(y[7945]), .Z(n50535) );
  AND U41521 ( .A(n21483), .B(n50535), .Z(n21485) );
  NANDN U41522 ( .A(y[7946]), .B(x[7946]), .Z(n21484) );
  NANDN U41523 ( .A(y[7947]), .B(x[7947]), .Z(n49871) );
  AND U41524 ( .A(n21484), .B(n49871), .Z(n50534) );
  NANDN U41525 ( .A(n21485), .B(n50534), .Z(n21486) );
  NAND U41526 ( .A(n21487), .B(n21486), .Z(n21488) );
  AND U41527 ( .A(n60980), .B(n21488), .Z(n21490) );
  XNOR U41528 ( .A(x[7950]), .B(y[7950]), .Z(n22042) );
  ANDN U41529 ( .B(y[7949]), .A(x[7949]), .Z(n60981) );
  ANDN U41530 ( .B(n22042), .A(n60981), .Z(n21489) );
  NANDN U41531 ( .A(n21490), .B(n21489), .Z(n21492) );
  NANDN U41532 ( .A(y[7950]), .B(x[7950]), .Z(n21491) );
  NANDN U41533 ( .A(y[7951]), .B(x[7951]), .Z(n22039) );
  AND U41534 ( .A(n21491), .B(n22039), .Z(n50532) );
  AND U41535 ( .A(n21492), .B(n50532), .Z(n21493) );
  NOR U41536 ( .A(n49879), .B(n21493), .Z(n21494) );
  NAND U41537 ( .A(n22040), .B(n21494), .Z(n21495) );
  NAND U41538 ( .A(n60984), .B(n21495), .Z(n21496) );
  AND U41539 ( .A(n22038), .B(n21496), .Z(n21497) );
  NANDN U41540 ( .A(n60985), .B(n21497), .Z(n21498) );
  AND U41541 ( .A(n60987), .B(n21498), .Z(n21499) );
  OR U41542 ( .A(n21500), .B(n21499), .Z(n21501) );
  NAND U41543 ( .A(n60988), .B(n21501), .Z(n21502) );
  NAND U41544 ( .A(n60989), .B(n21502), .Z(n21503) );
  NAND U41545 ( .A(n60990), .B(n21503), .Z(n21504) );
  AND U41546 ( .A(n22032), .B(n21504), .Z(n21505) );
  NANDN U41547 ( .A(x[7959]), .B(y[7959]), .Z(n60992) );
  AND U41548 ( .A(n21505), .B(n60992), .Z(n21506) );
  OR U41549 ( .A(n60995), .B(n21506), .Z(n21507) );
  NAND U41550 ( .A(n21508), .B(n21507), .Z(n21509) );
  NAND U41551 ( .A(n60998), .B(n21509), .Z(n21510) );
  AND U41552 ( .A(n49909), .B(n21510), .Z(n21511) );
  NANDN U41553 ( .A(x[7963]), .B(y[7963]), .Z(n50529) );
  AND U41554 ( .A(n21511), .B(n50529), .Z(n21513) );
  NANDN U41555 ( .A(y[7964]), .B(x[7964]), .Z(n21512) );
  NANDN U41556 ( .A(y[7965]), .B(x[7965]), .Z(n22027) );
  NAND U41557 ( .A(n21512), .B(n22027), .Z(n50527) );
  OR U41558 ( .A(n21513), .B(n50527), .Z(n21514) );
  NAND U41559 ( .A(n60999), .B(n21514), .Z(n21515) );
  NAND U41560 ( .A(n61000), .B(n21515), .Z(n21516) );
  NAND U41561 ( .A(n61001), .B(n21516), .Z(n21517) );
  NAND U41562 ( .A(n61002), .B(n21517), .Z(n21518) );
  AND U41563 ( .A(n22021), .B(n21518), .Z(n21519) );
  NANDN U41564 ( .A(x[7969]), .B(y[7969]), .Z(n61004) );
  AND U41565 ( .A(n21519), .B(n61004), .Z(n21521) );
  NANDN U41566 ( .A(y[7970]), .B(x[7970]), .Z(n21520) );
  NANDN U41567 ( .A(y[7971]), .B(x[7971]), .Z(n49928) );
  AND U41568 ( .A(n21520), .B(n49928), .Z(n50526) );
  NANDN U41569 ( .A(n21521), .B(n50526), .Z(n21522) );
  NAND U41570 ( .A(n21523), .B(n21522), .Z(n21524) );
  NAND U41571 ( .A(n61008), .B(n21524), .Z(n21525) );
  AND U41572 ( .A(n22019), .B(n21525), .Z(n21526) );
  ANDN U41573 ( .B(y[7973]), .A(x[7973]), .Z(n61009) );
  ANDN U41574 ( .B(n21526), .A(n61009), .Z(n21527) );
  OR U41575 ( .A(n61011), .B(n21527), .Z(n21528) );
  NAND U41576 ( .A(n21529), .B(n21528), .Z(n21530) );
  NAND U41577 ( .A(n61014), .B(n21530), .Z(n21531) );
  AND U41578 ( .A(n22017), .B(n21531), .Z(n21532) );
  ANDN U41579 ( .B(y[7977]), .A(x[7977]), .Z(n61015) );
  ANDN U41580 ( .B(n21532), .A(n61015), .Z(n21534) );
  NANDN U41581 ( .A(y[7978]), .B(x[7978]), .Z(n21533) );
  NANDN U41582 ( .A(y[7979]), .B(x[7979]), .Z(n22014) );
  AND U41583 ( .A(n21533), .B(n22014), .Z(n61017) );
  NANDN U41584 ( .A(n21534), .B(n61017), .Z(n21535) );
  AND U41585 ( .A(n22015), .B(n21535), .Z(n21536) );
  NANDN U41586 ( .A(x[7979]), .B(y[7979]), .Z(n50524) );
  AND U41587 ( .A(n21536), .B(n50524), .Z(n21538) );
  NANDN U41588 ( .A(y[7980]), .B(x[7980]), .Z(n21537) );
  NANDN U41589 ( .A(y[7981]), .B(x[7981]), .Z(n22012) );
  AND U41590 ( .A(n21537), .B(n22012), .Z(n61018) );
  NANDN U41591 ( .A(n21538), .B(n61018), .Z(n21539) );
  AND U41592 ( .A(n22013), .B(n21539), .Z(n21540) );
  NANDN U41593 ( .A(x[7981]), .B(y[7981]), .Z(n61019) );
  NAND U41594 ( .A(n21540), .B(n61019), .Z(n21541) );
  NAND U41595 ( .A(n61021), .B(n21541), .Z(n21542) );
  AND U41596 ( .A(n49957), .B(n21542), .Z(n21543) );
  NANDN U41597 ( .A(x[7983]), .B(y[7983]), .Z(n50523) );
  AND U41598 ( .A(n21543), .B(n50523), .Z(n21545) );
  NANDN U41599 ( .A(y[7984]), .B(x[7984]), .Z(n21544) );
  NANDN U41600 ( .A(y[7985]), .B(x[7985]), .Z(n22010) );
  AND U41601 ( .A(n21544), .B(n22010), .Z(n50521) );
  NANDN U41602 ( .A(n21545), .B(n50521), .Z(n21546) );
  NAND U41603 ( .A(n21547), .B(n21546), .Z(n21548) );
  NAND U41604 ( .A(n61026), .B(n21548), .Z(n21549) );
  AND U41605 ( .A(n49967), .B(n21549), .Z(n21550) );
  NANDN U41606 ( .A(x[7987]), .B(y[7987]), .Z(n61027) );
  AND U41607 ( .A(n21550), .B(n61027), .Z(n21552) );
  NANDN U41608 ( .A(y[7988]), .B(x[7988]), .Z(n21551) );
  NANDN U41609 ( .A(y[7989]), .B(x[7989]), .Z(n22008) );
  NAND U41610 ( .A(n21551), .B(n22008), .Z(n61028) );
  OR U41611 ( .A(n21552), .B(n61028), .Z(n21553) );
  NAND U41612 ( .A(n21554), .B(n21553), .Z(n21555) );
  NAND U41613 ( .A(n61031), .B(n21555), .Z(n21556) );
  AND U41614 ( .A(n22007), .B(n21556), .Z(n21557) );
  NANDN U41615 ( .A(x[7991]), .B(y[7991]), .Z(n61032) );
  AND U41616 ( .A(n21557), .B(n61032), .Z(n21559) );
  NANDN U41617 ( .A(y[7992]), .B(x[7992]), .Z(n21558) );
  NANDN U41618 ( .A(y[7993]), .B(x[7993]), .Z(n22004) );
  NAND U41619 ( .A(n21558), .B(n22004), .Z(n61034) );
  OR U41620 ( .A(n21559), .B(n61034), .Z(n21560) );
  NAND U41621 ( .A(n21561), .B(n21560), .Z(n21562) );
  NAND U41622 ( .A(n61035), .B(n21562), .Z(n21563) );
  AND U41623 ( .A(n49985), .B(n21563), .Z(n21564) );
  NANDN U41624 ( .A(x[7995]), .B(y[7995]), .Z(n61037) );
  NAND U41625 ( .A(n21564), .B(n61037), .Z(n21566) );
  NANDN U41626 ( .A(y[7996]), .B(x[7996]), .Z(n21565) );
  NANDN U41627 ( .A(y[7997]), .B(x[7997]), .Z(n22002) );
  AND U41628 ( .A(n21565), .B(n22002), .Z(n61040) );
  AND U41629 ( .A(n21566), .B(n61040), .Z(n21568) );
  XNOR U41630 ( .A(x[7998]), .B(y[7998]), .Z(n22003) );
  ANDN U41631 ( .B(y[7997]), .A(x[7997]), .Z(n50516) );
  ANDN U41632 ( .B(n22003), .A(n50516), .Z(n21567) );
  NANDN U41633 ( .A(n21568), .B(n21567), .Z(n21569) );
  NANDN U41634 ( .A(n61041), .B(n21569), .Z(n21570) );
  XOR U41635 ( .A(x[8000]), .B(y[8000]), .Z(n49997) );
  ANDN U41636 ( .B(n21570), .A(n49997), .Z(n21571) );
  NANDN U41637 ( .A(x[7999]), .B(y[7999]), .Z(n61042) );
  AND U41638 ( .A(n21571), .B(n61042), .Z(n21573) );
  NANDN U41639 ( .A(y[8000]), .B(x[8000]), .Z(n21572) );
  NANDN U41640 ( .A(y[8001]), .B(x[8001]), .Z(n22000) );
  AND U41641 ( .A(n21572), .B(n22000), .Z(n61044) );
  NANDN U41642 ( .A(n21573), .B(n61044), .Z(n21574) );
  AND U41643 ( .A(n22001), .B(n21574), .Z(n21575) );
  NANDN U41644 ( .A(x[8001]), .B(y[8001]), .Z(n61045) );
  AND U41645 ( .A(n21575), .B(n61045), .Z(n21577) );
  NANDN U41646 ( .A(y[8002]), .B(x[8002]), .Z(n21576) );
  NANDN U41647 ( .A(y[8003]), .B(x[8003]), .Z(n21998) );
  NAND U41648 ( .A(n21576), .B(n21998), .Z(n61047) );
  OR U41649 ( .A(n21577), .B(n61047), .Z(n21578) );
  NAND U41650 ( .A(n21579), .B(n21578), .Z(n21580) );
  NAND U41651 ( .A(n61050), .B(n21580), .Z(n21581) );
  AND U41652 ( .A(n21997), .B(n21581), .Z(n21582) );
  NANDN U41653 ( .A(x[8005]), .B(y[8005]), .Z(n61051) );
  AND U41654 ( .A(n21582), .B(n61051), .Z(n21584) );
  NANDN U41655 ( .A(y[8006]), .B(x[8006]), .Z(n21583) );
  NANDN U41656 ( .A(y[8007]), .B(x[8007]), .Z(n50012) );
  NAND U41657 ( .A(n21583), .B(n50012), .Z(n61053) );
  OR U41658 ( .A(n21584), .B(n61053), .Z(n21585) );
  NAND U41659 ( .A(n21586), .B(n21585), .Z(n21587) );
  NAND U41660 ( .A(n61056), .B(n21587), .Z(n21588) );
  AND U41661 ( .A(n21995), .B(n21588), .Z(n21589) );
  NANDN U41662 ( .A(n61057), .B(n21589), .Z(n21591) );
  NANDN U41663 ( .A(y[8010]), .B(x[8010]), .Z(n21590) );
  NANDN U41664 ( .A(y[8011]), .B(x[8011]), .Z(n50022) );
  AND U41665 ( .A(n21590), .B(n50022), .Z(n61059) );
  AND U41666 ( .A(n21591), .B(n61059), .Z(n21593) );
  XNOR U41667 ( .A(x[8012]), .B(y[8012]), .Z(n50023) );
  NANDN U41668 ( .A(x[8011]), .B(y[8011]), .Z(n50513) );
  AND U41669 ( .A(n50023), .B(n50513), .Z(n21592) );
  NANDN U41670 ( .A(n21593), .B(n21592), .Z(n21594) );
  NANDN U41671 ( .A(n61060), .B(n21594), .Z(n21595) );
  AND U41672 ( .A(n21993), .B(n21595), .Z(n21596) );
  NANDN U41673 ( .A(n61061), .B(n21596), .Z(n21597) );
  NAND U41674 ( .A(n61063), .B(n21597), .Z(n21598) );
  AND U41675 ( .A(n50033), .B(n21598), .Z(n21599) );
  NANDN U41676 ( .A(x[8015]), .B(y[8015]), .Z(n61064) );
  AND U41677 ( .A(n21599), .B(n61064), .Z(n21601) );
  NANDN U41678 ( .A(y[8016]), .B(x[8016]), .Z(n21600) );
  NANDN U41679 ( .A(y[8017]), .B(x[8017]), .Z(n21990) );
  AND U41680 ( .A(n21600), .B(n21990), .Z(n50511) );
  NANDN U41681 ( .A(n21601), .B(n50511), .Z(n21602) );
  NAND U41682 ( .A(n21603), .B(n21602), .Z(n21604) );
  NAND U41683 ( .A(n61069), .B(n21604), .Z(n21605) );
  AND U41684 ( .A(n50043), .B(n21605), .Z(n21606) );
  NANDN U41685 ( .A(x[8019]), .B(y[8019]), .Z(n61070) );
  AND U41686 ( .A(n21606), .B(n61070), .Z(n21608) );
  NANDN U41687 ( .A(y[8020]), .B(x[8020]), .Z(n21607) );
  NANDN U41688 ( .A(y[8021]), .B(x[8021]), .Z(n21987) );
  NAND U41689 ( .A(n21607), .B(n21987), .Z(n61072) );
  OR U41690 ( .A(n21608), .B(n61072), .Z(n21609) );
  AND U41691 ( .A(n21610), .B(n21609), .Z(n21612) );
  NANDN U41692 ( .A(y[8022]), .B(x[8022]), .Z(n21611) );
  NANDN U41693 ( .A(y[8023]), .B(x[8023]), .Z(n50053) );
  AND U41694 ( .A(n21611), .B(n50053), .Z(n61073) );
  NANDN U41695 ( .A(n21612), .B(n61073), .Z(n21613) );
  NAND U41696 ( .A(n21614), .B(n21613), .Z(n21615) );
  NAND U41697 ( .A(n61076), .B(n21615), .Z(n21616) );
  AND U41698 ( .A(n21986), .B(n21616), .Z(n21617) );
  ANDN U41699 ( .B(y[8025]), .A(x[8025]), .Z(n50507) );
  ANDN U41700 ( .B(n21617), .A(n50507), .Z(n21618) );
  OR U41701 ( .A(n61077), .B(n21618), .Z(n21619) );
  AND U41702 ( .A(n50064), .B(n21619), .Z(n21620) );
  NANDN U41703 ( .A(x[8027]), .B(y[8027]), .Z(n61078) );
  NAND U41704 ( .A(n21620), .B(n61078), .Z(n21621) );
  AND U41705 ( .A(n61080), .B(n21621), .Z(n21622) );
  ANDN U41706 ( .B(y[8029]), .A(x[8029]), .Z(n61081) );
  OR U41707 ( .A(n21622), .B(n61081), .Z(n21623) );
  XNOR U41708 ( .A(x[8030]), .B(y[8030]), .Z(n21984) );
  NANDN U41709 ( .A(n21623), .B(n21984), .Z(n21624) );
  NAND U41710 ( .A(n50506), .B(n21624), .Z(n21625) );
  NANDN U41711 ( .A(n21626), .B(n21625), .Z(n21627) );
  NAND U41712 ( .A(n61086), .B(n21627), .Z(n21628) );
  AND U41713 ( .A(n21982), .B(n21628), .Z(n21629) );
  ANDN U41714 ( .B(y[8033]), .A(x[8033]), .Z(n61087) );
  ANDN U41715 ( .B(n21629), .A(n61087), .Z(n21631) );
  NANDN U41716 ( .A(y[8034]), .B(x[8034]), .Z(n21630) );
  NANDN U41717 ( .A(y[8035]), .B(x[8035]), .Z(n50083) );
  NAND U41718 ( .A(n21630), .B(n50083), .Z(n61089) );
  OR U41719 ( .A(n21631), .B(n61089), .Z(n21632) );
  NAND U41720 ( .A(n21633), .B(n21632), .Z(n21634) );
  NAND U41721 ( .A(n61090), .B(n21634), .Z(n21635) );
  AND U41722 ( .A(n21980), .B(n21635), .Z(n21636) );
  NANDN U41723 ( .A(n61091), .B(n21636), .Z(n21638) );
  NANDN U41724 ( .A(y[8038]), .B(x[8038]), .Z(n21637) );
  NANDN U41725 ( .A(y[8039]), .B(x[8039]), .Z(n50094) );
  AND U41726 ( .A(n21637), .B(n50094), .Z(n61093) );
  AND U41727 ( .A(n21638), .B(n61093), .Z(n21639) );
  NOR U41728 ( .A(n50091), .B(n21639), .Z(n21640) );
  NAND U41729 ( .A(n50095), .B(n21640), .Z(n21641) );
  NANDN U41730 ( .A(n61094), .B(n21641), .Z(n21642) );
  AND U41731 ( .A(n21978), .B(n21642), .Z(n21643) );
  NANDN U41732 ( .A(n61095), .B(n21643), .Z(n21644) );
  AND U41733 ( .A(n61098), .B(n21644), .Z(n21645) );
  OR U41734 ( .A(n21646), .B(n21645), .Z(n21647) );
  NAND U41735 ( .A(n50500), .B(n21647), .Z(n21648) );
  NANDN U41736 ( .A(n21649), .B(n21648), .Z(n21650) );
  NAND U41737 ( .A(n61102), .B(n21650), .Z(n21651) );
  AND U41738 ( .A(n50115), .B(n21651), .Z(n21652) );
  NANDN U41739 ( .A(x[8047]), .B(y[8047]), .Z(n61103) );
  AND U41740 ( .A(n21652), .B(n61103), .Z(n21654) );
  NANDN U41741 ( .A(y[8048]), .B(x[8048]), .Z(n21653) );
  NANDN U41742 ( .A(y[8049]), .B(x[8049]), .Z(n21972) );
  NAND U41743 ( .A(n21653), .B(n21972), .Z(n61105) );
  OR U41744 ( .A(n21654), .B(n61105), .Z(n21655) );
  NAND U41745 ( .A(n21656), .B(n21655), .Z(n21657) );
  NAND U41746 ( .A(n61106), .B(n21657), .Z(n21658) );
  AND U41747 ( .A(n21971), .B(n21658), .Z(n21659) );
  NANDN U41748 ( .A(x[8051]), .B(y[8051]), .Z(n61107) );
  NAND U41749 ( .A(n21659), .B(n61107), .Z(n21661) );
  NANDN U41750 ( .A(y[8052]), .B(x[8052]), .Z(n21660) );
  NANDN U41751 ( .A(y[8053]), .B(x[8053]), .Z(n21969) );
  AND U41752 ( .A(n21660), .B(n21969), .Z(n61109) );
  AND U41753 ( .A(n21661), .B(n61109), .Z(n21662) );
  NANDN U41754 ( .A(x[8053]), .B(y[8053]), .Z(n50126) );
  NANDN U41755 ( .A(x[8054]), .B(y[8054]), .Z(n50132) );
  NAND U41756 ( .A(n50126), .B(n50132), .Z(n50497) );
  OR U41757 ( .A(n21662), .B(n50497), .Z(n21663) );
  NAND U41758 ( .A(n50496), .B(n21663), .Z(n21664) );
  NANDN U41759 ( .A(n50131), .B(n21664), .Z(n21665) );
  XNOR U41760 ( .A(x[8056]), .B(y[8056]), .Z(n21967) );
  NANDN U41761 ( .A(n21665), .B(n21967), .Z(n21666) );
  NAND U41762 ( .A(n61114), .B(n21666), .Z(n21667) );
  AND U41763 ( .A(n21965), .B(n21667), .Z(n21668) );
  NANDN U41764 ( .A(x[8057]), .B(y[8057]), .Z(n61115) );
  AND U41765 ( .A(n21668), .B(n61115), .Z(n21670) );
  NANDN U41766 ( .A(y[8058]), .B(x[8058]), .Z(n21669) );
  NANDN U41767 ( .A(y[8059]), .B(x[8059]), .Z(n21962) );
  NAND U41768 ( .A(n21669), .B(n21962), .Z(n50495) );
  OR U41769 ( .A(n21670), .B(n50495), .Z(n21671) );
  NAND U41770 ( .A(n50494), .B(n21671), .Z(n21672) );
  NAND U41771 ( .A(n61117), .B(n21672), .Z(n21673) );
  AND U41772 ( .A(n21959), .B(n21673), .Z(n21674) );
  NANDN U41773 ( .A(x[8061]), .B(y[8061]), .Z(n61118) );
  AND U41774 ( .A(n21674), .B(n61118), .Z(n21676) );
  NANDN U41775 ( .A(y[8062]), .B(x[8062]), .Z(n21675) );
  NANDN U41776 ( .A(y[8063]), .B(x[8063]), .Z(n50152) );
  AND U41777 ( .A(n21675), .B(n50152), .Z(n61120) );
  NANDN U41778 ( .A(n21676), .B(n61120), .Z(n21677) );
  NAND U41779 ( .A(n21678), .B(n21677), .Z(n21679) );
  NAND U41780 ( .A(n50491), .B(n21679), .Z(n21680) );
  NAND U41781 ( .A(n61123), .B(n21680), .Z(n21681) );
  NANDN U41782 ( .A(n61124), .B(n21681), .Z(n21682) );
  AND U41783 ( .A(n50163), .B(n21682), .Z(n21683) );
  NANDN U41784 ( .A(x[8067]), .B(y[8067]), .Z(n50490) );
  NAND U41785 ( .A(n21683), .B(n50490), .Z(n21684) );
  AND U41786 ( .A(n61125), .B(n21684), .Z(n21686) );
  XNOR U41787 ( .A(x[8070]), .B(y[8070]), .Z(n21953) );
  ANDN U41788 ( .B(y[8069]), .A(x[8069]), .Z(n50488) );
  ANDN U41789 ( .B(n21953), .A(n50488), .Z(n21685) );
  NANDN U41790 ( .A(n21686), .B(n21685), .Z(n21687) );
  NAND U41791 ( .A(n61126), .B(n21687), .Z(n21688) );
  AND U41792 ( .A(n50173), .B(n21688), .Z(n21689) );
  NANDN U41793 ( .A(x[8071]), .B(y[8071]), .Z(n61127) );
  NAND U41794 ( .A(n21689), .B(n61127), .Z(n21691) );
  NANDN U41795 ( .A(y[8072]), .B(x[8072]), .Z(n21690) );
  NANDN U41796 ( .A(y[8073]), .B(x[8073]), .Z(n21950) );
  AND U41797 ( .A(n21690), .B(n21950), .Z(n61129) );
  AND U41798 ( .A(n21691), .B(n61129), .Z(n21693) );
  XNOR U41799 ( .A(x[8074]), .B(y[8074]), .Z(n21951) );
  ANDN U41800 ( .B(y[8073]), .A(x[8073]), .Z(n50485) );
  ANDN U41801 ( .B(n21951), .A(n50485), .Z(n21692) );
  NANDN U41802 ( .A(n21693), .B(n21692), .Z(n21694) );
  NANDN U41803 ( .A(n61131), .B(n21694), .Z(n21695) );
  AND U41804 ( .A(n61132), .B(n21695), .Z(n21696) );
  NAND U41805 ( .A(n21949), .B(n21696), .Z(n21697) );
  NAND U41806 ( .A(n61134), .B(n21697), .Z(n21698) );
  NANDN U41807 ( .A(x[8077]), .B(y[8077]), .Z(n21947) );
  NANDN U41808 ( .A(x[8078]), .B(y[8078]), .Z(n21944) );
  AND U41809 ( .A(n21947), .B(n21944), .Z(n61135) );
  AND U41810 ( .A(n21698), .B(n61135), .Z(n21699) );
  ANDN U41811 ( .B(x[8079]), .A(y[8079]), .Z(n50193) );
  NANDN U41812 ( .A(y[8078]), .B(x[8078]), .Z(n21945) );
  NANDN U41813 ( .A(n50193), .B(n21945), .Z(n50484) );
  OR U41814 ( .A(n21699), .B(n50484), .Z(n21700) );
  NAND U41815 ( .A(n50483), .B(n21700), .Z(n21701) );
  NAND U41816 ( .A(n61136), .B(n21701), .Z(n21702) );
  AND U41817 ( .A(n21941), .B(n21702), .Z(n21703) );
  NANDN U41818 ( .A(x[8081]), .B(y[8081]), .Z(n61137) );
  NAND U41819 ( .A(n21703), .B(n61137), .Z(n21704) );
  AND U41820 ( .A(n61139), .B(n21704), .Z(n21705) );
  OR U41821 ( .A(n21706), .B(n21705), .Z(n21707) );
  NAND U41822 ( .A(n50480), .B(n21707), .Z(n21708) );
  NANDN U41823 ( .A(n21709), .B(n21708), .Z(n21710) );
  NAND U41824 ( .A(n61143), .B(n21710), .Z(n21711) );
  AND U41825 ( .A(n50211), .B(n21711), .Z(n21712) );
  NANDN U41826 ( .A(x[8087]), .B(y[8087]), .Z(n61144) );
  AND U41827 ( .A(n21712), .B(n61144), .Z(n21714) );
  NANDN U41828 ( .A(y[8088]), .B(x[8088]), .Z(n21713) );
  NANDN U41829 ( .A(y[8089]), .B(x[8089]), .Z(n21935) );
  NAND U41830 ( .A(n21713), .B(n21935), .Z(n61146) );
  OR U41831 ( .A(n21714), .B(n61146), .Z(n21715) );
  NAND U41832 ( .A(n21716), .B(n21715), .Z(n21717) );
  NAND U41833 ( .A(n61147), .B(n21717), .Z(n21718) );
  AND U41834 ( .A(n50221), .B(n21718), .Z(n21719) );
  NANDN U41835 ( .A(x[8091]), .B(y[8091]), .Z(n61148) );
  AND U41836 ( .A(n21719), .B(n61148), .Z(n21720) );
  OR U41837 ( .A(n61150), .B(n21720), .Z(n21721) );
  NAND U41838 ( .A(n21722), .B(n21721), .Z(n21723) );
  NANDN U41839 ( .A(n61151), .B(n21723), .Z(n21724) );
  AND U41840 ( .A(n50231), .B(n21724), .Z(n21725) );
  NANDN U41841 ( .A(x[8095]), .B(y[8095]), .Z(n61152) );
  NAND U41842 ( .A(n21725), .B(n61152), .Z(n21726) );
  AND U41843 ( .A(n61154), .B(n21726), .Z(n21728) );
  XNOR U41844 ( .A(x[8098]), .B(y[8098]), .Z(n21932) );
  ANDN U41845 ( .B(y[8097]), .A(x[8097]), .Z(n61155) );
  ANDN U41846 ( .B(n21932), .A(n61155), .Z(n21727) );
  NANDN U41847 ( .A(n21728), .B(n21727), .Z(n21729) );
  NANDN U41848 ( .A(n61158), .B(n21729), .Z(n21730) );
  AND U41849 ( .A(n50241), .B(n21730), .Z(n21731) );
  NANDN U41850 ( .A(x[8099]), .B(y[8099]), .Z(n61159) );
  NAND U41851 ( .A(n21731), .B(n61159), .Z(n21732) );
  NAND U41852 ( .A(n61160), .B(n21732), .Z(n21733) );
  AND U41853 ( .A(n21930), .B(n21733), .Z(n21734) );
  ANDN U41854 ( .B(y[8101]), .A(x[8101]), .Z(n61161) );
  ANDN U41855 ( .B(n21734), .A(n61161), .Z(n21736) );
  NANDN U41856 ( .A(y[8102]), .B(x[8102]), .Z(n21735) );
  NANDN U41857 ( .A(y[8103]), .B(x[8103]), .Z(n50251) );
  AND U41858 ( .A(n21735), .B(n50251), .Z(n61163) );
  NANDN U41859 ( .A(n21736), .B(n61163), .Z(n21737) );
  NAND U41860 ( .A(n21738), .B(n21737), .Z(n21739) );
  NAND U41861 ( .A(n61164), .B(n21739), .Z(n21740) );
  AND U41862 ( .A(n21928), .B(n21740), .Z(n21741) );
  ANDN U41863 ( .B(y[8105]), .A(x[8105]), .Z(n61165) );
  ANDN U41864 ( .B(n21741), .A(n61165), .Z(n21743) );
  NANDN U41865 ( .A(y[8106]), .B(x[8106]), .Z(n21742) );
  NANDN U41866 ( .A(y[8107]), .B(x[8107]), .Z(n21925) );
  AND U41867 ( .A(n21742), .B(n21925), .Z(n61167) );
  NANDN U41868 ( .A(n21743), .B(n61167), .Z(n21744) );
  NAND U41869 ( .A(n21745), .B(n21744), .Z(n21746) );
  NAND U41870 ( .A(n61170), .B(n21746), .Z(n21747) );
  AND U41871 ( .A(n21924), .B(n21747), .Z(n21748) );
  NANDN U41872 ( .A(x[8109]), .B(y[8109]), .Z(n61171) );
  AND U41873 ( .A(n21748), .B(n61171), .Z(n21750) );
  NANDN U41874 ( .A(y[8110]), .B(x[8110]), .Z(n21749) );
  NANDN U41875 ( .A(y[8111]), .B(x[8111]), .Z(n50269) );
  AND U41876 ( .A(n21749), .B(n50269), .Z(n61174) );
  NANDN U41877 ( .A(n21750), .B(n61174), .Z(n21751) );
  NAND U41878 ( .A(n21752), .B(n21751), .Z(n21753) );
  NANDN U41879 ( .A(n61176), .B(n21753), .Z(n21754) );
  AND U41880 ( .A(n21922), .B(n21754), .Z(n21755) );
  NANDN U41881 ( .A(n61177), .B(n21755), .Z(n21756) );
  AND U41882 ( .A(n61179), .B(n21756), .Z(n21758) );
  XNOR U41883 ( .A(x[8116]), .B(y[8116]), .Z(n50280) );
  NANDN U41884 ( .A(x[8115]), .B(y[8115]), .Z(n50470) );
  AND U41885 ( .A(n50280), .B(n50470), .Z(n21757) );
  NANDN U41886 ( .A(n21758), .B(n21757), .Z(n21759) );
  NAND U41887 ( .A(n61180), .B(n21759), .Z(n21760) );
  AND U41888 ( .A(n21920), .B(n21760), .Z(n21761) );
  NANDN U41889 ( .A(n61182), .B(n21761), .Z(n21763) );
  NANDN U41890 ( .A(y[8118]), .B(x[8118]), .Z(n21762) );
  NANDN U41891 ( .A(y[8119]), .B(x[8119]), .Z(n50290) );
  AND U41892 ( .A(n21762), .B(n50290), .Z(n50469) );
  AND U41893 ( .A(n21763), .B(n50469), .Z(n21764) );
  NOR U41894 ( .A(n50287), .B(n21764), .Z(n21765) );
  NAND U41895 ( .A(n50291), .B(n21765), .Z(n21766) );
  NANDN U41896 ( .A(n61185), .B(n21766), .Z(n21767) );
  AND U41897 ( .A(n21918), .B(n21767), .Z(n21768) );
  NANDN U41898 ( .A(n61187), .B(n21768), .Z(n21769) );
  NAND U41899 ( .A(n61189), .B(n21769), .Z(n21770) );
  AND U41900 ( .A(n50301), .B(n21770), .Z(n21771) );
  NANDN U41901 ( .A(x[8123]), .B(y[8123]), .Z(n50468) );
  AND U41902 ( .A(n21771), .B(n50468), .Z(n21773) );
  NANDN U41903 ( .A(y[8124]), .B(x[8124]), .Z(n21772) );
  NANDN U41904 ( .A(y[8125]), .B(x[8125]), .Z(n21915) );
  NAND U41905 ( .A(n21772), .B(n21915), .Z(n61190) );
  OR U41906 ( .A(n21773), .B(n61190), .Z(n21774) );
  NAND U41907 ( .A(n21775), .B(n21774), .Z(n21776) );
  NANDN U41908 ( .A(n61193), .B(n21776), .Z(n21777) );
  AND U41909 ( .A(n21914), .B(n21777), .Z(n21778) );
  NANDN U41910 ( .A(x[8127]), .B(y[8127]), .Z(n61194) );
  NAND U41911 ( .A(n21778), .B(n61194), .Z(n21780) );
  NANDN U41912 ( .A(y[8128]), .B(x[8128]), .Z(n21779) );
  NANDN U41913 ( .A(y[8129]), .B(x[8129]), .Z(n21911) );
  AND U41914 ( .A(n21779), .B(n21911), .Z(n61196) );
  AND U41915 ( .A(n21780), .B(n61196), .Z(n21782) );
  XNOR U41916 ( .A(x[8130]), .B(y[8130]), .Z(n21912) );
  NANDN U41917 ( .A(x[8129]), .B(y[8129]), .Z(n61197) );
  AND U41918 ( .A(n21912), .B(n61197), .Z(n21781) );
  NANDN U41919 ( .A(n21782), .B(n21781), .Z(n21783) );
  NAND U41920 ( .A(n61199), .B(n21783), .Z(n21784) );
  AND U41921 ( .A(n50319), .B(n21784), .Z(n21785) );
  NANDN U41922 ( .A(x[8131]), .B(y[8131]), .Z(n61201) );
  NAND U41923 ( .A(n21785), .B(n61201), .Z(n21786) );
  NAND U41924 ( .A(n61204), .B(n21786), .Z(n21787) );
  AND U41925 ( .A(n21909), .B(n21787), .Z(n21788) );
  NANDN U41926 ( .A(x[8133]), .B(y[8133]), .Z(n21910) );
  AND U41927 ( .A(n21788), .B(n21910), .Z(n21790) );
  NANDN U41928 ( .A(y[8134]), .B(x[8134]), .Z(n21789) );
  NANDN U41929 ( .A(y[8135]), .B(x[8135]), .Z(n21906) );
  AND U41930 ( .A(n21789), .B(n21906), .Z(n61209) );
  NANDN U41931 ( .A(n21790), .B(n61209), .Z(n21791) );
  NAND U41932 ( .A(n21792), .B(n21791), .Z(n21793) );
  NAND U41933 ( .A(n61214), .B(n21793), .Z(n21794) );
  AND U41934 ( .A(n21905), .B(n21794), .Z(n21795) );
  ANDN U41935 ( .B(y[8137]), .A(x[8137]), .Z(n50463) );
  ANDN U41936 ( .B(n21795), .A(n50463), .Z(n21797) );
  NANDN U41937 ( .A(y[8138]), .B(x[8138]), .Z(n21796) );
  NANDN U41938 ( .A(y[8139]), .B(x[8139]), .Z(n50337) );
  NAND U41939 ( .A(n21796), .B(n50337), .Z(n61219) );
  OR U41940 ( .A(n21797), .B(n61219), .Z(n21798) );
  NAND U41941 ( .A(n21799), .B(n21798), .Z(n21800) );
  AND U41942 ( .A(n61225), .B(n21800), .Z(n21802) );
  XNOR U41943 ( .A(x[8142]), .B(y[8142]), .Z(n21903) );
  ANDN U41944 ( .B(y[8141]), .A(x[8141]), .Z(n61226) );
  ANDN U41945 ( .B(n21903), .A(n61226), .Z(n21801) );
  NANDN U41946 ( .A(n21802), .B(n21801), .Z(n21803) );
  NANDN U41947 ( .A(n61231), .B(n21803), .Z(n21804) );
  AND U41948 ( .A(n50348), .B(n21804), .Z(n21805) );
  NANDN U41949 ( .A(x[8143]), .B(y[8143]), .Z(n61233) );
  NAND U41950 ( .A(n21805), .B(n61233), .Z(n21806) );
  NAND U41951 ( .A(n61237), .B(n21806), .Z(n21807) );
  NANDN U41952 ( .A(n61238), .B(n21807), .Z(n21808) );
  NAND U41953 ( .A(n61240), .B(n21808), .Z(n21809) );
  AND U41954 ( .A(n50358), .B(n21809), .Z(n21810) );
  NANDN U41955 ( .A(x[8147]), .B(y[8147]), .Z(n50461) );
  AND U41956 ( .A(n21810), .B(n50461), .Z(n21812) );
  NANDN U41957 ( .A(y[8148]), .B(x[8148]), .Z(n21811) );
  NANDN U41958 ( .A(y[8149]), .B(x[8149]), .Z(n21898) );
  AND U41959 ( .A(n21811), .B(n21898), .Z(n61241) );
  NANDN U41960 ( .A(n21812), .B(n61241), .Z(n21813) );
  NAND U41961 ( .A(n61242), .B(n21813), .Z(n21814) );
  NANDN U41962 ( .A(n61243), .B(n21814), .Z(n21815) );
  NAND U41963 ( .A(n61244), .B(n21815), .Z(n21816) );
  NANDN U41964 ( .A(y[8152]), .B(x[8152]), .Z(n21893) );
  NANDN U41965 ( .A(y[8153]), .B(x[8153]), .Z(n21892) );
  AND U41966 ( .A(n21893), .B(n21892), .Z(n50460) );
  AND U41967 ( .A(n21816), .B(n50460), .Z(n21817) );
  NANDN U41968 ( .A(x[8154]), .B(y[8154]), .Z(n21890) );
  ANDN U41969 ( .B(y[8153]), .A(x[8153]), .Z(n50370) );
  ANDN U41970 ( .B(n21890), .A(n50370), .Z(n61245) );
  NANDN U41971 ( .A(n21817), .B(n61245), .Z(n21818) );
  NAND U41972 ( .A(n61246), .B(n21818), .Z(n21819) );
  NANDN U41973 ( .A(n61247), .B(n21819), .Z(n21820) );
  NAND U41974 ( .A(n61248), .B(n21820), .Z(n21821) );
  AND U41975 ( .A(n21886), .B(n21821), .Z(n21822) );
  NANDN U41976 ( .A(n50458), .B(n21822), .Z(n21823) );
  NAND U41977 ( .A(n61249), .B(n21823), .Z(n21824) );
  AND U41978 ( .A(n50387), .B(n21824), .Z(n21825) );
  NAND U41979 ( .A(n50455), .B(n21825), .Z(n21826) );
  NANDN U41980 ( .A(n61251), .B(n21826), .Z(n21827) );
  AND U41981 ( .A(n21884), .B(n21827), .Z(n21828) );
  NANDN U41982 ( .A(n50454), .B(n21828), .Z(n21829) );
  AND U41983 ( .A(n61252), .B(n21829), .Z(n21830) );
  NANDN U41984 ( .A(x[8163]), .B(y[8163]), .Z(n50452) );
  NANDN U41985 ( .A(n21830), .B(n50452), .Z(n21831) );
  NAND U41986 ( .A(n61253), .B(n21831), .Z(n21832) );
  NANDN U41987 ( .A(n21833), .B(n21832), .Z(n21834) );
  NAND U41988 ( .A(n61256), .B(n21834), .Z(n21835) );
  AND U41989 ( .A(n21880), .B(n21835), .Z(n21836) );
  NANDN U41990 ( .A(x[8167]), .B(y[8167]), .Z(n50449) );
  AND U41991 ( .A(n21836), .B(n50449), .Z(n21837) );
  OR U41992 ( .A(n61257), .B(n21837), .Z(n21838) );
  NAND U41993 ( .A(n21839), .B(n21838), .Z(n21840) );
  NANDN U41994 ( .A(n50448), .B(n21840), .Z(n21841) );
  AND U41995 ( .A(n21876), .B(n21841), .Z(n21842) );
  NANDN U41996 ( .A(x[8171]), .B(y[8171]), .Z(n61261) );
  AND U41997 ( .A(n21842), .B(n61261), .Z(n21844) );
  NANDN U41998 ( .A(y[8172]), .B(x[8172]), .Z(n21843) );
  NANDN U41999 ( .A(y[8173]), .B(x[8173]), .Z(n21873) );
  NAND U42000 ( .A(n21843), .B(n21873), .Z(n61263) );
  OR U42001 ( .A(n21844), .B(n61263), .Z(n21845) );
  AND U42002 ( .A(n21874), .B(n21845), .Z(n21846) );
  NANDN U42003 ( .A(x[8173]), .B(y[8173]), .Z(n61264) );
  AND U42004 ( .A(n21846), .B(n61264), .Z(n21848) );
  NANDN U42005 ( .A(y[8174]), .B(x[8174]), .Z(n21847) );
  NANDN U42006 ( .A(y[8175]), .B(x[8175]), .Z(n50423) );
  AND U42007 ( .A(n21847), .B(n50423), .Z(n61266) );
  NANDN U42008 ( .A(n21848), .B(n61266), .Z(n21849) );
  NAND U42009 ( .A(n21850), .B(n21849), .Z(n21851) );
  NAND U42010 ( .A(n61269), .B(n21851), .Z(n21852) );
  AND U42011 ( .A(n21872), .B(n21852), .Z(n21853) );
  NANDN U42012 ( .A(x[8177]), .B(y[8177]), .Z(n50447) );
  NAND U42013 ( .A(n21853), .B(n50447), .Z(n21854) );
  AND U42014 ( .A(n61270), .B(n21854), .Z(n21855) );
  XNOR U42015 ( .A(x[8180]), .B(y[8180]), .Z(n50434) );
  NANDN U42016 ( .A(n21855), .B(n50434), .Z(n21856) );
  NANDN U42017 ( .A(n61273), .B(n21856), .Z(n21857) );
  AND U42018 ( .A(n21870), .B(n21857), .Z(n21858) );
  NANDN U42019 ( .A(n50444), .B(n21858), .Z(n21859) );
  NAND U42020 ( .A(n61275), .B(n21859), .Z(n21860) );
  AND U42021 ( .A(n21861), .B(n21860), .Z(n21864) );
  NANDN U42022 ( .A(y[8184]), .B(x[8184]), .Z(n21863) );
  NANDN U42023 ( .A(y[8185]), .B(x[8185]), .Z(n21862) );
  AND U42024 ( .A(n21863), .B(n21862), .Z(n61277) );
  NANDN U42025 ( .A(n21864), .B(n61277), .Z(n21865) );
  NAND U42026 ( .A(n21866), .B(n21865), .Z(n21867) );
  AND U42027 ( .A(n21868), .B(n21867), .Z(n50442) );
  AND U42028 ( .A(n21870), .B(n21869), .Z(n50440) );
  ANDN U42029 ( .B(y[8180]), .A(x[8180]), .Z(n61272) );
  NOR U42030 ( .A(n61272), .B(n50444), .Z(n50438) );
  AND U42031 ( .A(n21872), .B(n21871), .Z(n50430) );
  ANDN U42032 ( .B(y[8176]), .A(x[8176]), .Z(n61268) );
  ANDN U42033 ( .B(n50447), .A(n61268), .Z(n50428) );
  AND U42034 ( .A(n21874), .B(n21873), .Z(n50419) );
  NANDN U42035 ( .A(x[8172]), .B(y[8172]), .Z(n61262) );
  AND U42036 ( .A(n61262), .B(n61264), .Z(n50417) );
  NAND U42037 ( .A(n21876), .B(n21875), .Z(n50415) );
  AND U42038 ( .A(n21878), .B(n21877), .Z(n50411) );
  NANDN U42039 ( .A(x[8168]), .B(y[8168]), .Z(n50450) );
  NAND U42040 ( .A(n50450), .B(n61258), .Z(n50409) );
  AND U42041 ( .A(n21880), .B(n21879), .Z(n50407) );
  NANDN U42042 ( .A(x[8166]), .B(y[8166]), .Z(n61255) );
  NAND U42043 ( .A(n61255), .B(n50449), .Z(n50405) );
  AND U42044 ( .A(n21882), .B(n21881), .Z(n50403) );
  ANDN U42045 ( .B(y[8164]), .A(x[8164]), .Z(n50451) );
  NOR U42046 ( .A(n50451), .B(n61254), .Z(n50401) );
  AND U42047 ( .A(n21884), .B(n21883), .Z(n50393) );
  ANDN U42048 ( .B(y[8160]), .A(x[8160]), .Z(n50456) );
  NOR U42049 ( .A(n50456), .B(n50454), .Z(n50391) );
  AND U42050 ( .A(n21886), .B(n21885), .Z(n50383) );
  AND U42051 ( .A(n21888), .B(n21887), .Z(n50378) );
  NAND U42052 ( .A(n21890), .B(n21889), .Z(n50376) );
  AND U42053 ( .A(n21892), .B(n21891), .Z(n50374) );
  AND U42054 ( .A(n21894), .B(n21893), .Z(n50368) );
  NAND U42055 ( .A(n21896), .B(n21895), .Z(n50366) );
  AND U42056 ( .A(n21898), .B(n21897), .Z(n50364) );
  ANDN U42057 ( .B(y[8148]), .A(x[8148]), .Z(n50462) );
  NOR U42058 ( .A(n50462), .B(n21899), .Z(n50362) );
  XNOR U42059 ( .A(y[8146]), .B(x[8146]), .Z(n21900) );
  AND U42060 ( .A(n21901), .B(n21900), .Z(n50354) );
  NANDN U42061 ( .A(x[8144]), .B(y[8144]), .Z(n61234) );
  ANDN U42062 ( .B(n61234), .A(n61238), .Z(n50352) );
  AND U42063 ( .A(n21903), .B(n21902), .Z(n50344) );
  NANDN U42064 ( .A(x[8140]), .B(y[8140]), .Z(n61222) );
  ANDN U42065 ( .B(n61222), .A(n61226), .Z(n50342) );
  AND U42066 ( .A(n21905), .B(n21904), .Z(n50334) );
  AND U42067 ( .A(n21907), .B(n21906), .Z(n50330) );
  ANDN U42068 ( .B(y[8134]), .A(x[8134]), .Z(n50465) );
  AND U42069 ( .A(n21909), .B(n21908), .Z(n50325) );
  NANDN U42070 ( .A(x[8132]), .B(y[8132]), .Z(n61202) );
  IV U42071 ( .A(n21910), .Z(n50466) );
  ANDN U42072 ( .B(n61202), .A(n50466), .Z(n50323) );
  AND U42073 ( .A(n21912), .B(n21911), .Z(n50315) );
  NANDN U42074 ( .A(x[8128]), .B(y[8128]), .Z(n61195) );
  AND U42075 ( .A(n61195), .B(n61197), .Z(n50313) );
  NAND U42076 ( .A(n21914), .B(n21913), .Z(n50311) );
  NANDN U42077 ( .A(x[8126]), .B(y[8126]), .Z(n61191) );
  AND U42078 ( .A(n61194), .B(n61191), .Z(n50309) );
  AND U42079 ( .A(n21916), .B(n21915), .Z(n50307) );
  ANDN U42080 ( .B(y[8124]), .A(x[8124]), .Z(n50467) );
  ANDN U42081 ( .B(n61192), .A(n50467), .Z(n50305) );
  AND U42082 ( .A(n21918), .B(n21917), .Z(n50297) );
  ANDN U42083 ( .B(y[8120]), .A(x[8120]), .Z(n61184) );
  NOR U42084 ( .A(n61184), .B(n61187), .Z(n50295) );
  AND U42085 ( .A(n21920), .B(n21919), .Z(n50286) );
  ANDN U42086 ( .B(y[8116]), .A(x[8116]), .Z(n50471) );
  NOR U42087 ( .A(n50471), .B(n61182), .Z(n50284) );
  AND U42088 ( .A(n21922), .B(n21921), .Z(n50276) );
  ANDN U42089 ( .B(y[8112]), .A(x[8112]), .Z(n50472) );
  NOR U42090 ( .A(n50472), .B(n61177), .Z(n50274) );
  AND U42091 ( .A(n21924), .B(n21923), .Z(n50266) );
  NAND U42092 ( .A(n21926), .B(n21925), .Z(n50262) );
  NANDN U42093 ( .A(x[8106]), .B(y[8106]), .Z(n61166) );
  AND U42094 ( .A(n21928), .B(n21927), .Z(n50258) );
  NANDN U42095 ( .A(x[8104]), .B(y[8104]), .Z(n50474) );
  ANDN U42096 ( .B(n50474), .A(n61165), .Z(n50256) );
  AND U42097 ( .A(n21930), .B(n21929), .Z(n50247) );
  ANDN U42098 ( .B(y[8100]), .A(x[8100]), .Z(n50475) );
  NOR U42099 ( .A(n50475), .B(n61161), .Z(n50245) );
  AND U42100 ( .A(n21932), .B(n21931), .Z(n50237) );
  NANDN U42101 ( .A(x[8096]), .B(y[8096]), .Z(n61153) );
  ANDN U42102 ( .B(n61153), .A(n61155), .Z(n50235) );
  AND U42103 ( .A(n21934), .B(n21933), .Z(n50227) );
  ANDN U42104 ( .B(y[8092]), .A(x[8092]), .Z(n61149) );
  NOR U42105 ( .A(n61149), .B(n50476), .Z(n50225) );
  AND U42106 ( .A(n21936), .B(n21935), .Z(n50217) );
  NANDN U42107 ( .A(x[8088]), .B(y[8088]), .Z(n61145) );
  IV U42108 ( .A(n21937), .Z(n50478) );
  ANDN U42109 ( .B(n61145), .A(n50478), .Z(n50215) );
  AND U42110 ( .A(n21939), .B(n21938), .Z(n50207) );
  ANDN U42111 ( .B(y[8084]), .A(x[8084]), .Z(n50482) );
  NOR U42112 ( .A(n50482), .B(n61140), .Z(n50205) );
  AND U42113 ( .A(n21941), .B(n21940), .Z(n50197) );
  AND U42114 ( .A(n21942), .B(n61137), .Z(n50195) );
  AND U42115 ( .A(n21944), .B(n21943), .Z(n50189) );
  NAND U42116 ( .A(n21946), .B(n21945), .Z(n50187) );
  NANDN U42117 ( .A(x[8076]), .B(y[8076]), .Z(n61133) );
  AND U42118 ( .A(n61133), .B(n21947), .Z(n50185) );
  NAND U42119 ( .A(n21949), .B(n21948), .Z(n50183) );
  AND U42120 ( .A(n21951), .B(n21950), .Z(n50179) );
  ANDN U42121 ( .B(y[8072]), .A(x[8072]), .Z(n61128) );
  NOR U42122 ( .A(n61128), .B(n50485), .Z(n50177) );
  AND U42123 ( .A(n21953), .B(n21952), .Z(n50169) );
  ANDN U42124 ( .B(y[8068]), .A(x[8068]), .Z(n50489) );
  NOR U42125 ( .A(n50489), .B(n50488), .Z(n50167) );
  AND U42126 ( .A(n21954), .B(n50490), .Z(n50161) );
  AND U42127 ( .A(n21956), .B(n21955), .Z(n50159) );
  NANDN U42128 ( .A(x[8064]), .B(y[8064]), .Z(n50493) );
  ANDN U42129 ( .B(n50493), .A(n21957), .Z(n50157) );
  AND U42130 ( .A(n21959), .B(n21958), .Z(n50148) );
  NAND U42131 ( .A(n21960), .B(n61118), .Z(n50146) );
  AND U42132 ( .A(n21962), .B(n21961), .Z(n50144) );
  NANDN U42133 ( .A(x[8058]), .B(y[8058]), .Z(n61116) );
  NAND U42134 ( .A(n61116), .B(n21963), .Z(n50142) );
  AND U42135 ( .A(n21965), .B(n21964), .Z(n50140) );
  NAND U42136 ( .A(n21967), .B(n21966), .Z(n50136) );
  AND U42137 ( .A(n21969), .B(n21968), .Z(n50130) );
  NAND U42138 ( .A(n21971), .B(n21970), .Z(n50125) );
  NANDN U42139 ( .A(x[8050]), .B(y[8050]), .Z(n50499) );
  AND U42140 ( .A(n21973), .B(n21972), .Z(n50121) );
  NANDN U42141 ( .A(x[8048]), .B(y[8048]), .Z(n61104) );
  IV U42142 ( .A(n21974), .Z(n50498) );
  ANDN U42143 ( .B(n61104), .A(n50498), .Z(n50119) );
  AND U42144 ( .A(n21976), .B(n21975), .Z(n50111) );
  ANDN U42145 ( .B(y[8044]), .A(x[8044]), .Z(n50501) );
  NOR U42146 ( .A(n50501), .B(n61100), .Z(n50109) );
  AND U42147 ( .A(n21978), .B(n21977), .Z(n50101) );
  NANDN U42148 ( .A(x[8040]), .B(y[8040]), .Z(n50503) );
  ANDN U42149 ( .B(n50503), .A(n61095), .Z(n50099) );
  AND U42150 ( .A(n21980), .B(n21979), .Z(n50090) );
  ANDN U42151 ( .B(y[8036]), .A(x[8036]), .Z(n50505) );
  NOR U42152 ( .A(n50505), .B(n61091), .Z(n50088) );
  AND U42153 ( .A(n21982), .B(n21981), .Z(n50080) );
  NANDN U42154 ( .A(x[8032]), .B(y[8032]), .Z(n61085) );
  ANDN U42155 ( .B(n61085), .A(n61087), .Z(n50078) );
  AND U42156 ( .A(n21984), .B(n21983), .Z(n50070) );
  NANDN U42157 ( .A(x[8028]), .B(y[8028]), .Z(n61079) );
  ANDN U42158 ( .B(n61079), .A(n61081), .Z(n50068) );
  AND U42159 ( .A(n21986), .B(n21985), .Z(n50060) );
  ANDN U42160 ( .B(y[8024]), .A(x[8024]), .Z(n61075) );
  NOR U42161 ( .A(n61075), .B(n50507), .Z(n50058) );
  AND U42162 ( .A(n21988), .B(n21987), .Z(n50049) );
  NANDN U42163 ( .A(x[8020]), .B(y[8020]), .Z(n61071) );
  IV U42164 ( .A(n21989), .Z(n50509) );
  ANDN U42165 ( .B(n61071), .A(n50509), .Z(n50047) );
  AND U42166 ( .A(n21991), .B(n21990), .Z(n50039) );
  NANDN U42167 ( .A(x[8016]), .B(y[8016]), .Z(n61065) );
  ANDN U42168 ( .B(n61065), .A(n61066), .Z(n50037) );
  AND U42169 ( .A(n21993), .B(n21992), .Z(n50029) );
  ANDN U42170 ( .B(y[8012]), .A(x[8012]), .Z(n50512) );
  NOR U42171 ( .A(n50512), .B(n61061), .Z(n50027) );
  AND U42172 ( .A(n21995), .B(n21994), .Z(n50019) );
  ANDN U42173 ( .B(y[8008]), .A(x[8008]), .Z(n50515) );
  NOR U42174 ( .A(n50515), .B(n61057), .Z(n50017) );
  AND U42175 ( .A(n21997), .B(n21996), .Z(n50009) );
  NANDN U42176 ( .A(x[8004]), .B(y[8004]), .Z(n61049) );
  AND U42177 ( .A(n61049), .B(n61051), .Z(n50007) );
  NAND U42178 ( .A(n21999), .B(n21998), .Z(n50005) );
  AND U42179 ( .A(n22001), .B(n22000), .Z(n50001) );
  NANDN U42180 ( .A(x[8000]), .B(y[8000]), .Z(n61043) );
  AND U42181 ( .A(n61043), .B(n61045), .Z(n49999) );
  NANDN U42182 ( .A(x[7998]), .B(y[7998]), .Z(n50517) );
  AND U42183 ( .A(n22003), .B(n22002), .Z(n49991) );
  ANDN U42184 ( .B(y[7996]), .A(x[7996]), .Z(n61038) );
  NOR U42185 ( .A(n61038), .B(n50516), .Z(n49989) );
  AND U42186 ( .A(n22005), .B(n22004), .Z(n49981) );
  NANDN U42187 ( .A(x[7992]), .B(y[7992]), .Z(n61033) );
  AND U42188 ( .A(n61033), .B(n50518), .Z(n49979) );
  NAND U42189 ( .A(n22007), .B(n22006), .Z(n49977) );
  AND U42190 ( .A(n22009), .B(n22008), .Z(n49973) );
  ANDN U42191 ( .B(y[7988]), .A(x[7988]), .Z(n50520) );
  NOR U42192 ( .A(n50520), .B(n61029), .Z(n49971) );
  AND U42193 ( .A(n22011), .B(n22010), .Z(n49963) );
  NANDN U42194 ( .A(x[7984]), .B(y[7984]), .Z(n50522) );
  ANDN U42195 ( .B(n50522), .A(n61024), .Z(n49961) );
  AND U42196 ( .A(n22013), .B(n22012), .Z(n49953) );
  NAND U42197 ( .A(n22015), .B(n22014), .Z(n49949) );
  AND U42198 ( .A(n22017), .B(n22016), .Z(n49945) );
  NANDN U42199 ( .A(x[7976]), .B(y[7976]), .Z(n61013) );
  ANDN U42200 ( .B(n61013), .A(n61015), .Z(n49943) );
  AND U42201 ( .A(n22019), .B(n22018), .Z(n49935) );
  NANDN U42202 ( .A(x[7972]), .B(y[7972]), .Z(n61006) );
  ANDN U42203 ( .B(n61006), .A(n61009), .Z(n49933) );
  AND U42204 ( .A(n22021), .B(n22020), .Z(n49924) );
  AND U42205 ( .A(n22023), .B(n22022), .Z(n49919) );
  NAND U42206 ( .A(n22025), .B(n22024), .Z(n49917) );
  AND U42207 ( .A(n22027), .B(n22026), .Z(n49915) );
  ANDN U42208 ( .B(y[7964]), .A(x[7964]), .Z(n50528) );
  NOR U42209 ( .A(n50528), .B(n22028), .Z(n49913) );
  AND U42210 ( .A(n22030), .B(n22029), .Z(n49905) );
  AND U42211 ( .A(n22032), .B(n22031), .Z(n49901) );
  NAND U42212 ( .A(n60992), .B(n22033), .Z(n49899) );
  AND U42213 ( .A(n22035), .B(n22034), .Z(n49897) );
  ANDN U42214 ( .B(y[7956]), .A(x[7956]), .Z(n50531) );
  NOR U42215 ( .A(n50531), .B(n22036), .Z(n49895) );
  AND U42216 ( .A(n22038), .B(n22037), .Z(n49887) );
  AND U42217 ( .A(n22040), .B(n22039), .Z(n49883) );
  ANDN U42218 ( .B(y[7950]), .A(x[7950]), .Z(n50533) );
  AND U42219 ( .A(n22042), .B(n22041), .Z(n49878) );
  NANDN U42220 ( .A(x[7948]), .B(y[7948]), .Z(n60979) );
  ANDN U42221 ( .B(n60979), .A(n60981), .Z(n49876) );
  AND U42222 ( .A(n22044), .B(n22043), .Z(n49867) );
  NANDN U42223 ( .A(x[7944]), .B(y[7944]), .Z(n60975) );
  AND U42224 ( .A(n60975), .B(n50535), .Z(n49865) );
  NAND U42225 ( .A(n22046), .B(n22045), .Z(n49863) );
  NANDN U42226 ( .A(x[7942]), .B(y[7942]), .Z(n50538) );
  AND U42227 ( .A(n60974), .B(n50538), .Z(n49861) );
  AND U42228 ( .A(n22048), .B(n22047), .Z(n49859) );
  NANDN U42229 ( .A(x[7940]), .B(y[7940]), .Z(n60971) );
  IV U42230 ( .A(n22049), .Z(n50537) );
  ANDN U42231 ( .B(n60971), .A(n50537), .Z(n49857) );
  AND U42232 ( .A(n22051), .B(n22050), .Z(n49849) );
  ANDN U42233 ( .B(y[7936]), .A(x[7936]), .Z(n50539) );
  NOR U42234 ( .A(n50539), .B(n60967), .Z(n49847) );
  AND U42235 ( .A(n22053), .B(n22052), .Z(n49839) );
  ANDN U42236 ( .B(y[7932]), .A(x[7932]), .Z(n50541) );
  NOR U42237 ( .A(n50541), .B(n60961), .Z(n49837) );
  AND U42238 ( .A(n22055), .B(n22054), .Z(n49829) );
  ANDN U42239 ( .B(y[7928]), .A(x[7928]), .Z(n50544) );
  NOR U42240 ( .A(n50544), .B(n60958), .Z(n49827) );
  AND U42241 ( .A(n22057), .B(n22056), .Z(n49819) );
  NANDN U42242 ( .A(x[7924]), .B(y[7924]), .Z(n60951) );
  ANDN U42243 ( .B(n60951), .A(n60953), .Z(n49817) );
  AND U42244 ( .A(n22059), .B(n22058), .Z(n49808) );
  NANDN U42245 ( .A(x[7920]), .B(y[7920]), .Z(n60946) );
  ANDN U42246 ( .B(n60946), .A(n60948), .Z(n49806) );
  AND U42247 ( .A(n22061), .B(n22060), .Z(n49798) );
  ANDN U42248 ( .B(y[7916]), .A(x[7916]), .Z(n60942) );
  NOR U42249 ( .A(n60942), .B(n50546), .Z(n49796) );
  AND U42250 ( .A(n22063), .B(n22062), .Z(n49788) );
  NANDN U42251 ( .A(x[7912]), .B(y[7912]), .Z(n60936) );
  IV U42252 ( .A(n22064), .Z(n50548) );
  ANDN U42253 ( .B(n60936), .A(n50548), .Z(n49786) );
  AND U42254 ( .A(n22066), .B(n22065), .Z(n49778) );
  ANDN U42255 ( .B(y[7908]), .A(x[7908]), .Z(n50551) );
  NOR U42256 ( .A(n50551), .B(n60932), .Z(n49776) );
  AND U42257 ( .A(n22068), .B(n22067), .Z(n49768) );
  ANDN U42258 ( .B(y[7904]), .A(x[7904]), .Z(n50552) );
  NOR U42259 ( .A(n50552), .B(n60928), .Z(n49766) );
  AND U42260 ( .A(n22070), .B(n22069), .Z(n49758) );
  ANDN U42261 ( .B(y[7900]), .A(x[7900]), .Z(n50555) );
  NOR U42262 ( .A(n50555), .B(n60922), .Z(n49756) );
  AND U42263 ( .A(n22072), .B(n22071), .Z(n49748) );
  NANDN U42264 ( .A(x[7896]), .B(y[7896]), .Z(n60916) );
  ANDN U42265 ( .B(n60916), .A(n60918), .Z(n49746) );
  AND U42266 ( .A(n22074), .B(n22073), .Z(n49737) );
  NANDN U42267 ( .A(x[7892]), .B(y[7892]), .Z(n60911) );
  AND U42268 ( .A(n60911), .B(n60913), .Z(n49735) );
  NAND U42269 ( .A(n22076), .B(n22075), .Z(n49733) );
  AND U42270 ( .A(n22078), .B(n22077), .Z(n49729) );
  ANDN U42271 ( .B(y[7888]), .A(x[7888]), .Z(n60906) );
  NOR U42272 ( .A(n60906), .B(n50557), .Z(n49727) );
  AND U42273 ( .A(n22080), .B(n22079), .Z(n49719) );
  ANDN U42274 ( .B(y[7884]), .A(x[7884]), .Z(n60902) );
  NOR U42275 ( .A(n60902), .B(n50560), .Z(n49717) );
  AND U42276 ( .A(n22081), .B(n60901), .Z(n49711) );
  AND U42277 ( .A(n22083), .B(n22082), .Z(n49709) );
  NAND U42278 ( .A(n22085), .B(n22084), .Z(n49707) );
  AND U42279 ( .A(n22087), .B(n22086), .Z(n49705) );
  NANDN U42280 ( .A(x[7878]), .B(y[7878]), .Z(n60895) );
  NAND U42281 ( .A(n60895), .B(n22088), .Z(n49703) );
  AND U42282 ( .A(n22090), .B(n22089), .Z(n49701) );
  NAND U42283 ( .A(n22091), .B(n60894), .Z(n49699) );
  AND U42284 ( .A(n22093), .B(n22092), .Z(n49697) );
  ANDN U42285 ( .B(y[7874]), .A(x[7874]), .Z(n60890) );
  AND U42286 ( .A(n22095), .B(n22094), .Z(n49692) );
  NAND U42287 ( .A(n22096), .B(n60889), .Z(n49690) );
  AND U42288 ( .A(n22098), .B(n22097), .Z(n49688) );
  NANDN U42289 ( .A(x[7870]), .B(y[7870]), .Z(n50565) );
  AND U42290 ( .A(n22100), .B(n22099), .Z(n49683) );
  IV U42291 ( .A(n22101), .Z(n50564) );
  NAND U42292 ( .A(n50564), .B(n22102), .Z(n49681) );
  AND U42293 ( .A(n22104), .B(n22103), .Z(n49679) );
  NAND U42294 ( .A(n22106), .B(n22105), .Z(n49677) );
  AND U42295 ( .A(n22108), .B(n22107), .Z(n49675) );
  NANDN U42296 ( .A(x[7864]), .B(y[7864]), .Z(n50567) );
  AND U42297 ( .A(n50567), .B(n22109), .Z(n49673) );
  AND U42298 ( .A(n22110), .B(n50566), .Z(n49667) );
  NAND U42299 ( .A(n22112), .B(n22111), .Z(n49665) );
  NANDN U42300 ( .A(x[7860]), .B(y[7860]), .Z(n60876) );
  AND U42301 ( .A(n22113), .B(n60876), .Z(n49663) );
  NAND U42302 ( .A(n22115), .B(n22114), .Z(n49661) );
  AND U42303 ( .A(n22117), .B(n22116), .Z(n49657) );
  NANDN U42304 ( .A(x[7856]), .B(y[7856]), .Z(n60871) );
  ANDN U42305 ( .B(n60871), .A(n60874), .Z(n49655) );
  AND U42306 ( .A(n22119), .B(n22118), .Z(n49647) );
  ANDN U42307 ( .B(y[7852]), .A(x[7852]), .Z(n60865) );
  NOR U42308 ( .A(n60865), .B(n50569), .Z(n49645) );
  AND U42309 ( .A(n22121), .B(n22120), .Z(n49637) );
  ANDN U42310 ( .B(y[7848]), .A(x[7848]), .Z(n50571) );
  NOR U42311 ( .A(n50571), .B(n60861), .Z(n49635) );
  AND U42312 ( .A(n22123), .B(n22122), .Z(n49627) );
  AND U42313 ( .A(n22125), .B(n22124), .Z(n49623) );
  ANDN U42314 ( .B(y[7842]), .A(x[7842]), .Z(n60851) );
  AND U42315 ( .A(n22127), .B(n22126), .Z(n49618) );
  ANDN U42316 ( .B(y[7840]), .A(x[7840]), .Z(n50574) );
  NOR U42317 ( .A(n50574), .B(n60850), .Z(n49616) );
  AND U42318 ( .A(n22129), .B(n22128), .Z(n49607) );
  NANDN U42319 ( .A(x[7836]), .B(y[7836]), .Z(n60844) );
  AND U42320 ( .A(n60844), .B(n60846), .Z(n49605) );
  NAND U42321 ( .A(n22131), .B(n22130), .Z(n49603) );
  NANDN U42322 ( .A(x[7834]), .B(y[7834]), .Z(n50577) );
  AND U42323 ( .A(n50577), .B(n60843), .Z(n49601) );
  AND U42324 ( .A(n22133), .B(n22132), .Z(n49599) );
  ANDN U42325 ( .B(y[7832]), .A(x[7832]), .Z(n60838) );
  NOR U42326 ( .A(n60838), .B(n50576), .Z(n49597) );
  AND U42327 ( .A(n22135), .B(n22134), .Z(n49589) );
  NANDN U42328 ( .A(x[7828]), .B(y[7828]), .Z(n60834) );
  IV U42329 ( .A(n22136), .Z(n50578) );
  ANDN U42330 ( .B(n60834), .A(n50578), .Z(n49587) );
  AND U42331 ( .A(n22138), .B(n22137), .Z(n49579) );
  ANDN U42332 ( .B(y[7824]), .A(x[7824]), .Z(n50580) );
  NOR U42333 ( .A(n50580), .B(n60830), .Z(n49577) );
  AND U42334 ( .A(n22140), .B(n22139), .Z(n49569) );
  ANDN U42335 ( .B(y[7820]), .A(x[7820]), .Z(n50581) );
  NOR U42336 ( .A(n50581), .B(n60825), .Z(n49567) );
  AND U42337 ( .A(n22142), .B(n22141), .Z(n49559) );
  NAND U42338 ( .A(n22144), .B(n22143), .Z(n49555) );
  NANDN U42339 ( .A(x[7814]), .B(y[7814]), .Z(n60810) );
  AND U42340 ( .A(n22146), .B(n22145), .Z(n49551) );
  NANDN U42341 ( .A(x[7812]), .B(y[7812]), .Z(n60804) );
  ANDN U42342 ( .B(n60804), .A(n60808), .Z(n49549) );
  AND U42343 ( .A(n22148), .B(n22147), .Z(n49541) );
  NANDN U42344 ( .A(x[7808]), .B(y[7808]), .Z(n60792) );
  ANDN U42345 ( .B(n60792), .A(n60796), .Z(n49539) );
  AND U42346 ( .A(n22150), .B(n22149), .Z(n49531) );
  NANDN U42347 ( .A(x[7804]), .B(y[7804]), .Z(n60780) );
  AND U42348 ( .A(n60780), .B(n60785), .Z(n49529) );
  AND U42349 ( .A(n22152), .B(n22151), .Z(n49521) );
  ANDN U42350 ( .B(y[7800]), .A(x[7800]), .Z(n50589) );
  NOR U42351 ( .A(n50589), .B(n50587), .Z(n49519) );
  AND U42352 ( .A(n22154), .B(n22153), .Z(n49511) );
  NANDN U42353 ( .A(x[7796]), .B(y[7796]), .Z(n60774) );
  ANDN U42354 ( .B(n60774), .A(n60775), .Z(n49509) );
  AND U42355 ( .A(n22156), .B(n22155), .Z(n49501) );
  ANDN U42356 ( .B(y[7792]), .A(x[7792]), .Z(n50592) );
  NOR U42357 ( .A(n50592), .B(n60769), .Z(n49499) );
  AND U42358 ( .A(n22158), .B(n22157), .Z(n49491) );
  NANDN U42359 ( .A(x[7788]), .B(y[7788]), .Z(n50595) );
  ANDN U42360 ( .B(n50595), .A(n60765), .Z(n49489) );
  AND U42361 ( .A(n22160), .B(n22159), .Z(n49480) );
  ANDN U42362 ( .B(y[7784]), .A(x[7784]), .Z(n60761) );
  NOR U42363 ( .A(n60761), .B(n50596), .Z(n49478) );
  AND U42364 ( .A(n22162), .B(n22161), .Z(n49470) );
  ANDN U42365 ( .B(y[7780]), .A(x[7780]), .Z(n60756) );
  NOR U42366 ( .A(n60756), .B(n50598), .Z(n49468) );
  AND U42367 ( .A(n22164), .B(n22163), .Z(n49460) );
  NANDN U42368 ( .A(x[7776]), .B(y[7776]), .Z(n60752) );
  IV U42369 ( .A(n22165), .Z(n50600) );
  ANDN U42370 ( .B(n60752), .A(n50600), .Z(n49458) );
  AND U42371 ( .A(n22167), .B(n22166), .Z(n49450) );
  AND U42372 ( .A(n22169), .B(n22168), .Z(n49445) );
  NAND U42373 ( .A(n22171), .B(n22170), .Z(n49443) );
  AND U42374 ( .A(n22173), .B(n22172), .Z(n49441) );
  AND U42375 ( .A(n22175), .B(n22174), .Z(n49436) );
  IV U42376 ( .A(n22176), .Z(n50604) );
  NAND U42377 ( .A(n50604), .B(n22177), .Z(n49434) );
  AND U42378 ( .A(n22179), .B(n22178), .Z(n49432) );
  NANDN U42379 ( .A(x[7764]), .B(y[7764]), .Z(n60740) );
  ANDN U42380 ( .B(n60740), .A(n22180), .Z(n49430) );
  AND U42381 ( .A(n22182), .B(n22181), .Z(n49422) );
  NANDN U42382 ( .A(x[7760]), .B(y[7760]), .Z(n60734) );
  ANDN U42383 ( .B(n60734), .A(n60736), .Z(n49420) );
  AND U42384 ( .A(n22184), .B(n22183), .Z(n49411) );
  ANDN U42385 ( .B(y[7756]), .A(x[7756]), .Z(n60730) );
  NOR U42386 ( .A(n60730), .B(n50607), .Z(n49409) );
  AND U42387 ( .A(n22186), .B(n22185), .Z(n49401) );
  NANDN U42388 ( .A(x[7752]), .B(y[7752]), .Z(n60726) );
  IV U42389 ( .A(n22187), .Z(n50609) );
  ANDN U42390 ( .B(n60726), .A(n50609), .Z(n49399) );
  AND U42391 ( .A(n22189), .B(n22188), .Z(n49391) );
  ANDN U42392 ( .B(y[7748]), .A(x[7748]), .Z(n50611) );
  NOR U42393 ( .A(n50611), .B(n60722), .Z(n49389) );
  AND U42394 ( .A(n22191), .B(n22190), .Z(n49381) );
  ANDN U42395 ( .B(y[7744]), .A(x[7744]), .Z(n50613) );
  NOR U42396 ( .A(n50613), .B(n60716), .Z(n49379) );
  AND U42397 ( .A(n22193), .B(n22192), .Z(n49371) );
  ANDN U42398 ( .B(y[7740]), .A(x[7740]), .Z(n50616) );
  NOR U42399 ( .A(n50616), .B(n60713), .Z(n49369) );
  AND U42400 ( .A(n22195), .B(n22194), .Z(n49361) );
  NANDN U42401 ( .A(x[7736]), .B(y[7736]), .Z(n60704) );
  ANDN U42402 ( .B(n60704), .A(n60708), .Z(n49359) );
  AND U42403 ( .A(n22197), .B(n22196), .Z(n49351) );
  NANDN U42404 ( .A(x[7732]), .B(y[7732]), .Z(n60692) );
  ANDN U42405 ( .B(n60692), .A(n60696), .Z(n49349) );
  AND U42406 ( .A(n22199), .B(n22198), .Z(n49341) );
  NANDN U42407 ( .A(x[7728]), .B(y[7728]), .Z(n60682) );
  AND U42408 ( .A(n60682), .B(n50617), .Z(n49339) );
  NAND U42409 ( .A(n22201), .B(n22200), .Z(n49337) );
  AND U42410 ( .A(n22203), .B(n22202), .Z(n49333) );
  NANDN U42411 ( .A(x[7724]), .B(y[7724]), .Z(n60672) );
  IV U42412 ( .A(n22204), .Z(n50619) );
  ANDN U42413 ( .B(n60672), .A(n50619), .Z(n49331) );
  AND U42414 ( .A(n22206), .B(n22205), .Z(n49323) );
  ANDN U42415 ( .B(y[7720]), .A(x[7720]), .Z(n50621) );
  NOR U42416 ( .A(n50621), .B(n60668), .Z(n49321) );
  AND U42417 ( .A(n22208), .B(n22207), .Z(n49313) );
  NAND U42418 ( .A(n22210), .B(n22209), .Z(n49309) );
  AND U42419 ( .A(n22212), .B(n22211), .Z(n49305) );
  ANDN U42420 ( .B(y[7712]), .A(x[7712]), .Z(n50625) );
  NOR U42421 ( .A(n50625), .B(n60659), .Z(n49303) );
  AND U42422 ( .A(n22214), .B(n22213), .Z(n49295) );
  NANDN U42423 ( .A(x[7708]), .B(y[7708]), .Z(n60652) );
  ANDN U42424 ( .B(n60652), .A(n60654), .Z(n49293) );
  AND U42425 ( .A(n22216), .B(n22215), .Z(n49285) );
  NANDN U42426 ( .A(x[7704]), .B(y[7704]), .Z(n60646) );
  ANDN U42427 ( .B(n60646), .A(n60648), .Z(n49283) );
  AND U42428 ( .A(n22218), .B(n22217), .Z(n49275) );
  ANDN U42429 ( .B(y[7700]), .A(x[7700]), .Z(n60642) );
  NOR U42430 ( .A(n60642), .B(n50628), .Z(n49273) );
  IV U42431 ( .A(n22219), .Z(n60640) );
  AND U42432 ( .A(n22220), .B(n60640), .Z(n49267) );
  AND U42433 ( .A(n22222), .B(n22221), .Z(n49265) );
  ANDN U42434 ( .B(y[7696]), .A(x[7696]), .Z(n50630) );
  NOR U42435 ( .A(n50630), .B(n22223), .Z(n49263) );
  AND U42436 ( .A(n22225), .B(n22224), .Z(n49255) );
  ANDN U42437 ( .B(y[7692]), .A(x[7692]), .Z(n60632) );
  NOR U42438 ( .A(n60632), .B(n60634), .Z(n49253) );
  AND U42439 ( .A(n22227), .B(n22226), .Z(n49244) );
  ANDN U42440 ( .B(y[7688]), .A(x[7688]), .Z(n50633) );
  NOR U42441 ( .A(n50633), .B(n60629), .Z(n49242) );
  AND U42442 ( .A(n22229), .B(n22228), .Z(n49234) );
  NAND U42443 ( .A(n22230), .B(n50637), .Z(n49232) );
  AND U42444 ( .A(n22232), .B(n22231), .Z(n49230) );
  NANDN U42445 ( .A(x[7682]), .B(y[7682]), .Z(n50641) );
  NAND U42446 ( .A(n50641), .B(n22233), .Z(n49228) );
  AND U42447 ( .A(n22235), .B(n22234), .Z(n49226) );
  ANDN U42448 ( .B(y[7680]), .A(x[7680]), .Z(n60623) );
  NOR U42449 ( .A(n60623), .B(n50640), .Z(n49224) );
  AND U42450 ( .A(n22237), .B(n22236), .Z(n49216) );
  NANDN U42451 ( .A(x[7676]), .B(y[7676]), .Z(n60618) );
  AND U42452 ( .A(n60618), .B(n50642), .Z(n49214) );
  NAND U42453 ( .A(n22239), .B(n22238), .Z(n49212) );
  IV U42454 ( .A(n22240), .Z(n60617) );
  AND U42455 ( .A(n22241), .B(n60617), .Z(n49210) );
  AND U42456 ( .A(n22243), .B(n22242), .Z(n49208) );
  AND U42457 ( .A(n22245), .B(n22244), .Z(n49202) );
  NAND U42458 ( .A(n22247), .B(n22246), .Z(n49200) );
  AND U42459 ( .A(n22249), .B(n22248), .Z(n49198) );
  ANDN U42460 ( .B(y[7668]), .A(x[7668]), .Z(n50644) );
  NOR U42461 ( .A(n50644), .B(n22250), .Z(n49196) );
  AND U42462 ( .A(n22252), .B(n22251), .Z(n49188) );
  NANDN U42463 ( .A(x[7664]), .B(y[7664]), .Z(n60608) );
  ANDN U42464 ( .B(n60608), .A(n50648), .Z(n49186) );
  AND U42465 ( .A(n22254), .B(n22253), .Z(n49178) );
  NANDN U42466 ( .A(x[7660]), .B(y[7660]), .Z(n50650) );
  ANDN U42467 ( .B(n50650), .A(n60605), .Z(n49176) );
  AND U42468 ( .A(n22256), .B(n22255), .Z(n49167) );
  IV U42469 ( .A(n22257), .Z(n60599) );
  ANDN U42470 ( .B(y[7656]), .A(x[7656]), .Z(n60598) );
  NOR U42471 ( .A(n60599), .B(n60598), .Z(n49165) );
  AND U42472 ( .A(n22259), .B(n22258), .Z(n49157) );
  ANDN U42473 ( .B(y[7652]), .A(x[7652]), .Z(n60591) );
  NOR U42474 ( .A(n60591), .B(n60594), .Z(n49155) );
  AND U42475 ( .A(n22261), .B(n22260), .Z(n49147) );
  ANDN U42476 ( .B(y[7648]), .A(x[7648]), .Z(n50652) );
  NOR U42477 ( .A(n50652), .B(n60585), .Z(n49145) );
  AND U42478 ( .A(n22263), .B(n22262), .Z(n49137) );
  ANDN U42479 ( .B(y[7644]), .A(x[7644]), .Z(n60579) );
  NOR U42480 ( .A(n60579), .B(n60581), .Z(n49135) );
  AND U42481 ( .A(n22265), .B(n22264), .Z(n49126) );
  NANDN U42482 ( .A(x[7640]), .B(y[7640]), .Z(n60573) );
  ANDN U42483 ( .B(n60573), .A(n60576), .Z(n49124) );
  AND U42484 ( .A(n22267), .B(n22266), .Z(n49116) );
  AND U42485 ( .A(n22269), .B(n22268), .Z(n49112) );
  ANDN U42486 ( .B(y[7634]), .A(x[7634]), .Z(n50657) );
  AND U42487 ( .A(n22271), .B(n22270), .Z(n49108) );
  ANDN U42488 ( .B(y[7632]), .A(x[7632]), .Z(n50659) );
  NOR U42489 ( .A(n50659), .B(n60566), .Z(n49106) );
  AND U42490 ( .A(n22273), .B(n22272), .Z(n49098) );
  NANDN U42491 ( .A(x[7628]), .B(y[7628]), .Z(n50661) );
  AND U42492 ( .A(n50661), .B(n60562), .Z(n49096) );
  NAND U42493 ( .A(n22275), .B(n22274), .Z(n49094) );
  NANDN U42494 ( .A(x[7626]), .B(y[7626]), .Z(n60558) );
  AND U42495 ( .A(n60558), .B(n50660), .Z(n49092) );
  AND U42496 ( .A(n22277), .B(n22276), .Z(n49090) );
  NANDN U42497 ( .A(x[7624]), .B(y[7624]), .Z(n50663) );
  ANDN U42498 ( .B(n50663), .A(n60557), .Z(n49088) );
  AND U42499 ( .A(n22279), .B(n22278), .Z(n49080) );
  NAND U42500 ( .A(n22280), .B(n50665), .Z(n49078) );
  AND U42501 ( .A(n22282), .B(n22281), .Z(n49076) );
  NANDN U42502 ( .A(x[7618]), .B(y[7618]), .Z(n50670) );
  NAND U42503 ( .A(n50670), .B(n22283), .Z(n49074) );
  AND U42504 ( .A(n22285), .B(n22284), .Z(n49072) );
  NANDN U42505 ( .A(x[7616]), .B(y[7616]), .Z(n60551) );
  ANDN U42506 ( .B(n60551), .A(n50668), .Z(n49070) );
  AND U42507 ( .A(n22287), .B(n22286), .Z(n49062) );
  NANDN U42508 ( .A(x[7612]), .B(y[7612]), .Z(n60547) );
  IV U42509 ( .A(n22288), .Z(n50671) );
  ANDN U42510 ( .B(n60547), .A(n50671), .Z(n49060) );
  AND U42511 ( .A(n22290), .B(n22289), .Z(n49052) );
  ANDN U42512 ( .B(y[7608]), .A(x[7608]), .Z(n50673) );
  NOR U42513 ( .A(n50673), .B(n60543), .Z(n49050) );
  AND U42514 ( .A(n22292), .B(n22291), .Z(n49041) );
  ANDN U42515 ( .B(y[7604]), .A(x[7604]), .Z(n50674) );
  NOR U42516 ( .A(n50674), .B(n60538), .Z(n49039) );
  AND U42517 ( .A(n22294), .B(n22293), .Z(n49031) );
  ANDN U42518 ( .B(y[7600]), .A(x[7600]), .Z(n50677) );
  NOR U42519 ( .A(n50677), .B(n60532), .Z(n49029) );
  AND U42520 ( .A(n22296), .B(n22295), .Z(n49021) );
  NANDN U42521 ( .A(x[7596]), .B(y[7596]), .Z(n60526) );
  ANDN U42522 ( .B(n60526), .A(n60528), .Z(n49019) );
  AND U42523 ( .A(n22298), .B(n22297), .Z(n49011) );
  NANDN U42524 ( .A(x[7592]), .B(y[7592]), .Z(n60519) );
  ANDN U42525 ( .B(n60519), .A(n60522), .Z(n49009) );
  AND U42526 ( .A(n22300), .B(n22299), .Z(n49000) );
  ANDN U42527 ( .B(y[7588]), .A(x[7588]), .Z(n60516) );
  NOR U42528 ( .A(n60516), .B(n50679), .Z(n48998) );
  AND U42529 ( .A(n22302), .B(n22301), .Z(n48990) );
  ANDN U42530 ( .B(y[7584]), .A(x[7584]), .Z(n50683) );
  NOR U42531 ( .A(n50683), .B(n50682), .Z(n48988) );
  XNOR U42532 ( .A(x[7582]), .B(y[7582]), .Z(n22304) );
  AND U42533 ( .A(n22304), .B(n22303), .Z(n48980) );
  NAND U42534 ( .A(n22305), .B(n60510), .Z(n48978) );
  AND U42535 ( .A(n22307), .B(n22306), .Z(n48976) );
  ANDN U42536 ( .B(y[7578]), .A(x[7578]), .Z(n60505) );
  AND U42537 ( .A(n22309), .B(n22308), .Z(n48971) );
  AND U42538 ( .A(n22311), .B(n22310), .Z(n48967) );
  NAND U42539 ( .A(n50685), .B(n22312), .Z(n48965) );
  AND U42540 ( .A(n22314), .B(n22313), .Z(n48963) );
  NANDN U42541 ( .A(x[7572]), .B(y[7572]), .Z(n60499) );
  ANDN U42542 ( .B(n60499), .A(n22315), .Z(n48961) );
  AND U42543 ( .A(n22317), .B(n22316), .Z(n48953) );
  ANDN U42544 ( .B(y[7568]), .A(x[7568]), .Z(n60491) );
  NOR U42545 ( .A(n60491), .B(n60496), .Z(n48951) );
  AND U42546 ( .A(n22319), .B(n22318), .Z(n48943) );
  NANDN U42547 ( .A(x[7564]), .B(y[7564]), .Z(n60487) );
  ANDN U42548 ( .B(n60487), .A(n60488), .Z(n48941) );
  AND U42549 ( .A(n22321), .B(n22320), .Z(n48933) );
  ANDN U42550 ( .B(y[7560]), .A(x[7560]), .Z(n50688) );
  NOR U42551 ( .A(n50688), .B(n60483), .Z(n48931) );
  AND U42552 ( .A(n22323), .B(n22322), .Z(n48923) );
  ANDN U42553 ( .B(y[7556]), .A(x[7556]), .Z(n50690) );
  NOR U42554 ( .A(n50690), .B(n60477), .Z(n48921) );
  AND U42555 ( .A(n22325), .B(n22324), .Z(n48913) );
  NANDN U42556 ( .A(x[7552]), .B(y[7552]), .Z(n60471) );
  ANDN U42557 ( .B(n60471), .A(n60473), .Z(n48911) );
  AND U42558 ( .A(n22327), .B(n22326), .Z(n48903) );
  NANDN U42559 ( .A(x[7548]), .B(y[7548]), .Z(n60466) );
  ANDN U42560 ( .B(n60466), .A(n60468), .Z(n48901) );
  AND U42561 ( .A(n22329), .B(n22328), .Z(n48893) );
  ANDN U42562 ( .B(y[7544]), .A(x[7544]), .Z(n60460) );
  NOR U42563 ( .A(n60460), .B(n50693), .Z(n48891) );
  AND U42564 ( .A(n22331), .B(n22330), .Z(n48883) );
  NANDN U42565 ( .A(x[7540]), .B(y[7540]), .Z(n60456) );
  IV U42566 ( .A(n22332), .Z(n50695) );
  ANDN U42567 ( .B(n60456), .A(n50695), .Z(n48881) );
  AND U42568 ( .A(n22334), .B(n22333), .Z(n48873) );
  NANDN U42569 ( .A(x[7536]), .B(y[7536]), .Z(n60451) );
  ANDN U42570 ( .B(n60451), .A(n60452), .Z(n48871) );
  AND U42571 ( .A(n22336), .B(n22335), .Z(n48863) );
  ANDN U42572 ( .B(y[7532]), .A(x[7532]), .Z(n50698) );
  NOR U42573 ( .A(n50698), .B(n60446), .Z(n48861) );
  AND U42574 ( .A(n22338), .B(n22337), .Z(n48853) );
  ANDN U42575 ( .B(y[7528]), .A(x[7528]), .Z(n50701) );
  NOR U42576 ( .A(n50701), .B(n60442), .Z(n48851) );
  AND U42577 ( .A(n22340), .B(n22339), .Z(n48843) );
  NANDN U42578 ( .A(x[7524]), .B(y[7524]), .Z(n60435) );
  ANDN U42579 ( .B(n60435), .A(n60438), .Z(n48841) );
  AND U42580 ( .A(n22342), .B(n22341), .Z(n48833) );
  ANDN U42581 ( .B(y[7520]), .A(x[7520]), .Z(n60428) );
  NOR U42582 ( .A(n60428), .B(n60431), .Z(n48831) );
  AND U42583 ( .A(n22344), .B(n22343), .Z(n48823) );
  ANDN U42584 ( .B(y[7516]), .A(x[7516]), .Z(n60425) );
  NOR U42585 ( .A(n60425), .B(n50702), .Z(n48821) );
  AND U42586 ( .A(n22346), .B(n22345), .Z(n48813) );
  ANDN U42587 ( .B(y[7512]), .A(x[7512]), .Z(n60418) );
  NOR U42588 ( .A(n60418), .B(n60421), .Z(n48811) );
  AND U42589 ( .A(n22348), .B(n22347), .Z(n48802) );
  ANDN U42590 ( .B(y[7508]), .A(x[7508]), .Z(n60415) );
  NOR U42591 ( .A(n60415), .B(n50705), .Z(n48800) );
  AND U42592 ( .A(n22350), .B(n22349), .Z(n48792) );
  NANDN U42593 ( .A(x[7504]), .B(y[7504]), .Z(n60409) );
  ANDN U42594 ( .B(n60409), .A(n60411), .Z(n48790) );
  AND U42595 ( .A(n22352), .B(n22351), .Z(n48782) );
  ANDN U42596 ( .B(y[7500]), .A(x[7500]), .Z(n60405) );
  NOR U42597 ( .A(n60405), .B(n50708), .Z(n48780) );
  AND U42598 ( .A(n22354), .B(n22353), .Z(n48772) );
  AND U42599 ( .A(n22356), .B(n22355), .Z(n48767) );
  NAND U42600 ( .A(n22358), .B(n22357), .Z(n48765) );
  AND U42601 ( .A(n22360), .B(n22359), .Z(n48763) );
  NAND U42602 ( .A(n22362), .B(n22361), .Z(n48761) );
  AND U42603 ( .A(n22364), .B(n22363), .Z(n48759) );
  NAND U42604 ( .A(n22366), .B(n22365), .Z(n48757) );
  AND U42605 ( .A(n22368), .B(n22367), .Z(n48755) );
  AND U42606 ( .A(n22370), .B(n22369), .Z(n48749) );
  NAND U42607 ( .A(n22372), .B(n22371), .Z(n48747) );
  AND U42608 ( .A(n22374), .B(n22373), .Z(n48745) );
  NAND U42609 ( .A(n22376), .B(n22375), .Z(n48743) );
  AND U42610 ( .A(n22378), .B(n22377), .Z(n48741) );
  ANDN U42611 ( .B(y[7482]), .A(x[7482]), .Z(n50712) );
  AND U42612 ( .A(n22380), .B(n22379), .Z(n48736) );
  AND U42613 ( .A(n22382), .B(n22381), .Z(n48732) );
  NAND U42614 ( .A(n22383), .B(n50715), .Z(n48730) );
  AND U42615 ( .A(n22385), .B(n22384), .Z(n48728) );
  ANDN U42616 ( .B(y[7476]), .A(x[7476]), .Z(n50718) );
  NOR U42617 ( .A(n50718), .B(n22386), .Z(n48726) );
  AND U42618 ( .A(n22388), .B(n22387), .Z(n48718) );
  ANDN U42619 ( .B(y[7472]), .A(x[7472]), .Z(n50720) );
  NOR U42620 ( .A(n50720), .B(n60381), .Z(n48716) );
  AND U42621 ( .A(n22390), .B(n22389), .Z(n48707) );
  IV U42622 ( .A(n22391), .Z(n60377) );
  AND U42623 ( .A(n22392), .B(n60377), .Z(n48705) );
  ANDN U42624 ( .B(y[7466]), .A(x[7466]), .Z(n48697) );
  AND U42625 ( .A(n22394), .B(n22393), .Z(n48695) );
  NANDN U42626 ( .A(x[7464]), .B(y[7464]), .Z(n60372) );
  AND U42627 ( .A(n60372), .B(n22395), .Z(n48693) );
  NAND U42628 ( .A(n22397), .B(n22396), .Z(n48691) );
  NANDN U42629 ( .A(x[7462]), .B(y[7462]), .Z(n50724) );
  IV U42630 ( .A(n22398), .Z(n60371) );
  AND U42631 ( .A(n50724), .B(n60371), .Z(n48689) );
  AND U42632 ( .A(n22400), .B(n22399), .Z(n48687) );
  ANDN U42633 ( .B(y[7460]), .A(x[7460]), .Z(n60366) );
  ANDN U42634 ( .B(n50723), .A(n60366), .Z(n48685) );
  AND U42635 ( .A(n22402), .B(n22401), .Z(n48677) );
  ANDN U42636 ( .B(y[7456]), .A(x[7456]), .Z(n60359) );
  NOR U42637 ( .A(n60359), .B(n60362), .Z(n48675) );
  AND U42638 ( .A(n22404), .B(n22403), .Z(n48667) );
  ANDN U42639 ( .B(y[7452]), .A(x[7452]), .Z(n60354) );
  NOR U42640 ( .A(n60354), .B(n60356), .Z(n48665) );
  AND U42641 ( .A(n22406), .B(n22405), .Z(n48656) );
  NANDN U42642 ( .A(x[7448]), .B(y[7448]), .Z(n60348) );
  ANDN U42643 ( .B(n60348), .A(n22407), .Z(n48654) );
  AND U42644 ( .A(n22409), .B(n22408), .Z(n48645) );
  ANDN U42645 ( .B(y[7444]), .A(x[7444]), .Z(n60345) );
  NOR U42646 ( .A(n60345), .B(n50726), .Z(n48643) );
  AND U42647 ( .A(n22411), .B(n22410), .Z(n48635) );
  ANDN U42648 ( .B(y[7440]), .A(x[7440]), .Z(n60341) );
  NOR U42649 ( .A(n60341), .B(n50729), .Z(n48633) );
  AND U42650 ( .A(n22413), .B(n22412), .Z(n48625) );
  NANDN U42651 ( .A(x[7436]), .B(y[7436]), .Z(n60334) );
  AND U42652 ( .A(n60334), .B(n60336), .Z(n48623) );
  NAND U42653 ( .A(n22415), .B(n22414), .Z(n48621) );
  AND U42654 ( .A(n22417), .B(n22416), .Z(n48617) );
  ANDN U42655 ( .B(y[7432]), .A(x[7432]), .Z(n50730) );
  NOR U42656 ( .A(n50730), .B(n60330), .Z(n48615) );
  AND U42657 ( .A(n22419), .B(n22418), .Z(n48607) );
  NANDN U42658 ( .A(x[7428]), .B(y[7428]), .Z(n50732) );
  AND U42659 ( .A(n50732), .B(n60326), .Z(n48605) );
  NAND U42660 ( .A(n22421), .B(n22420), .Z(n48603) );
  AND U42661 ( .A(n22423), .B(n22422), .Z(n48598) );
  NANDN U42662 ( .A(x[7424]), .B(y[7424]), .Z(n60320) );
  NAND U42663 ( .A(n60320), .B(n50734), .Z(n48596) );
  AND U42664 ( .A(n22425), .B(n22424), .Z(n48594) );
  NANDN U42665 ( .A(x[7422]), .B(y[7422]), .Z(n60316) );
  NAND U42666 ( .A(n60316), .B(n60319), .Z(n48592) );
  AND U42667 ( .A(n22427), .B(n22426), .Z(n48590) );
  ANDN U42668 ( .B(y[7420]), .A(x[7420]), .Z(n50737) );
  NOR U42669 ( .A(n50737), .B(n60317), .Z(n48588) );
  AND U42670 ( .A(n22429), .B(n22428), .Z(n48580) );
  NANDN U42671 ( .A(x[7416]), .B(y[7416]), .Z(n60312) );
  AND U42672 ( .A(n60312), .B(n60313), .Z(n48578) );
  AND U42673 ( .A(n22431), .B(n22430), .Z(n48570) );
  ANDN U42674 ( .B(y[7412]), .A(x[7412]), .Z(n60305) );
  NOR U42675 ( .A(n60305), .B(n60307), .Z(n48568) );
  AND U42676 ( .A(n22433), .B(n22432), .Z(n48560) );
  NANDN U42677 ( .A(x[7408]), .B(y[7408]), .Z(n50740) );
  ANDN U42678 ( .B(n50740), .A(n60301), .Z(n48558) );
  AND U42679 ( .A(n22435), .B(n22434), .Z(n48550) );
  ANDN U42680 ( .B(y[7404]), .A(x[7404]), .Z(n60294) );
  NOR U42681 ( .A(n60294), .B(n60297), .Z(n48548) );
  AND U42682 ( .A(n22437), .B(n22436), .Z(n48540) );
  NANDN U42683 ( .A(x[7400]), .B(y[7400]), .Z(n60287) );
  ANDN U42684 ( .B(n60287), .A(n60289), .Z(n48538) );
  AND U42685 ( .A(n22439), .B(n22438), .Z(n48530) );
  NAND U42686 ( .A(n60285), .B(n22440), .Z(n48528) );
  AND U42687 ( .A(n22442), .B(n22441), .Z(n48526) );
  NANDN U42688 ( .A(x[7394]), .B(y[7394]), .Z(n60280) );
  NAND U42689 ( .A(n60280), .B(n22443), .Z(n48524) );
  AND U42690 ( .A(n22445), .B(n22444), .Z(n48522) );
  NAND U42691 ( .A(n50743), .B(n22446), .Z(n48520) );
  AND U42692 ( .A(n22448), .B(n22447), .Z(n48518) );
  NANDN U42693 ( .A(x[7390]), .B(y[7390]), .Z(n60276) );
  AND U42694 ( .A(n22450), .B(n22449), .Z(n48513) );
  NANDN U42695 ( .A(x[7388]), .B(y[7388]), .Z(n50746) );
  ANDN U42696 ( .B(n50746), .A(n60275), .Z(n48511) );
  AND U42697 ( .A(n22452), .B(n22451), .Z(n48503) );
  ANDN U42698 ( .B(y[7384]), .A(x[7384]), .Z(n50748) );
  NOR U42699 ( .A(n50748), .B(n60272), .Z(n48501) );
  AND U42700 ( .A(n22453), .B(n50749), .Z(n48495) );
  AND U42701 ( .A(n22455), .B(n22454), .Z(n48493) );
  NANDN U42702 ( .A(x[7380]), .B(y[7380]), .Z(n60266) );
  NAND U42703 ( .A(n60266), .B(n22456), .Z(n48491) );
  AND U42704 ( .A(n22458), .B(n22457), .Z(n48489) );
  NANDN U42705 ( .A(x[7378]), .B(y[7378]), .Z(n60264) );
  NAND U42706 ( .A(n60264), .B(n60265), .Z(n48487) );
  AND U42707 ( .A(n22460), .B(n22459), .Z(n48485) );
  NANDN U42708 ( .A(x[7376]), .B(y[7376]), .Z(n50752) );
  IV U42709 ( .A(n22461), .Z(n60263) );
  ANDN U42710 ( .B(n50752), .A(n60263), .Z(n48483) );
  AND U42711 ( .A(n22463), .B(n22462), .Z(n48475) );
  NANDN U42712 ( .A(x[7372]), .B(y[7372]), .Z(n50756) );
  ANDN U42713 ( .B(n50756), .A(n50753), .Z(n48473) );
  AND U42714 ( .A(n22465), .B(n22464), .Z(n48464) );
  ANDN U42715 ( .B(y[7368]), .A(x[7368]), .Z(n50757) );
  NOR U42716 ( .A(n50757), .B(n60255), .Z(n48462) );
  AND U42717 ( .A(n22467), .B(n22466), .Z(n48454) );
  ANDN U42718 ( .B(y[7364]), .A(x[7364]), .Z(n22468) );
  NOR U42719 ( .A(n22468), .B(n60251), .Z(n48452) );
  AND U42720 ( .A(n22470), .B(n22469), .Z(n48443) );
  NANDN U42721 ( .A(x[7360]), .B(y[7360]), .Z(n60245) );
  AND U42722 ( .A(n60245), .B(n60247), .Z(n48441) );
  NAND U42723 ( .A(n22472), .B(n22471), .Z(n48439) );
  NANDN U42724 ( .A(x[7358]), .B(y[7358]), .Z(n60240) );
  AND U42725 ( .A(n60244), .B(n60240), .Z(n48437) );
  AND U42726 ( .A(n22474), .B(n22473), .Z(n48435) );
  NANDN U42727 ( .A(x[7356]), .B(y[7356]), .Z(n60238) );
  AND U42728 ( .A(n60238), .B(n60241), .Z(n48433) );
  AND U42729 ( .A(n22476), .B(n22475), .Z(n48425) );
  ANDN U42730 ( .B(y[7352]), .A(x[7352]), .Z(n60234) );
  NOR U42731 ( .A(n60234), .B(n50761), .Z(n48423) );
  AND U42732 ( .A(n22478), .B(n22477), .Z(n48415) );
  NANDN U42733 ( .A(x[7348]), .B(y[7348]), .Z(n22479) );
  NAND U42734 ( .A(n22479), .B(n60230), .Z(n48413) );
  AND U42735 ( .A(n22481), .B(n22480), .Z(n48411) );
  NANDN U42736 ( .A(x[7346]), .B(y[7346]), .Z(n60227) );
  NAND U42737 ( .A(n60227), .B(n22482), .Z(n48409) );
  AND U42738 ( .A(n22484), .B(n22483), .Z(n48407) );
  ANDN U42739 ( .B(y[7344]), .A(x[7344]), .Z(n50765) );
  NOR U42740 ( .A(n50765), .B(n60226), .Z(n48405) );
  AND U42741 ( .A(n22486), .B(n22485), .Z(n48397) );
  NAND U42742 ( .A(n22488), .B(n22487), .Z(n48393) );
  NANDN U42743 ( .A(x[7338]), .B(y[7338]), .Z(n60217) );
  AND U42744 ( .A(n22490), .B(n22489), .Z(n48389) );
  NANDN U42745 ( .A(x[7336]), .B(y[7336]), .Z(n60213) );
  ANDN U42746 ( .B(n60213), .A(n60215), .Z(n48387) );
  AND U42747 ( .A(n22492), .B(n22491), .Z(n48378) );
  ANDN U42748 ( .B(y[7332]), .A(x[7332]), .Z(n60210) );
  NOR U42749 ( .A(n60210), .B(n50767), .Z(n48376) );
  AND U42750 ( .A(n22494), .B(n22493), .Z(n48368) );
  NANDN U42751 ( .A(x[7328]), .B(y[7328]), .Z(n60206) );
  IV U42752 ( .A(n22495), .Z(n50769) );
  ANDN U42753 ( .B(n60206), .A(n50769), .Z(n48366) );
  AND U42754 ( .A(n22497), .B(n22496), .Z(n48358) );
  ANDN U42755 ( .B(y[7324]), .A(x[7324]), .Z(n50771) );
  NOR U42756 ( .A(n50771), .B(n60201), .Z(n48356) );
  AND U42757 ( .A(n22499), .B(n22498), .Z(n48348) );
  ANDN U42758 ( .B(y[7320]), .A(x[7320]), .Z(n50772) );
  NOR U42759 ( .A(n50772), .B(n60196), .Z(n48346) );
  AND U42760 ( .A(n22501), .B(n22500), .Z(n48338) );
  NANDN U42761 ( .A(x[7316]), .B(y[7316]), .Z(n50775) );
  IV U42762 ( .A(n22502), .Z(n60192) );
  AND U42763 ( .A(n50775), .B(n60192), .Z(n48336) );
  NAND U42764 ( .A(n22504), .B(n22503), .Z(n48334) );
  AND U42765 ( .A(n22506), .B(n22505), .Z(n48330) );
  NANDN U42766 ( .A(x[7312]), .B(y[7312]), .Z(n60185) );
  AND U42767 ( .A(n60185), .B(n60187), .Z(n48328) );
  NANDN U42768 ( .A(x[7310]), .B(y[7310]), .Z(n60182) );
  AND U42769 ( .A(n60182), .B(n60184), .Z(n48322) );
  NAND U42770 ( .A(n22508), .B(n22507), .Z(n48320) );
  NANDN U42771 ( .A(x[7308]), .B(y[7308]), .Z(n60179) );
  AND U42772 ( .A(n60179), .B(n60181), .Z(n48318) );
  AND U42773 ( .A(n22510), .B(n22509), .Z(n48310) );
  ANDN U42774 ( .B(y[7304]), .A(x[7304]), .Z(n60175) );
  NOR U42775 ( .A(n60175), .B(n50776), .Z(n48308) );
  AND U42776 ( .A(n22512), .B(n22511), .Z(n48300) );
  ANDN U42777 ( .B(y[7300]), .A(x[7300]), .Z(n50780) );
  NOR U42778 ( .A(n50780), .B(n50779), .Z(n48298) );
  AND U42779 ( .A(n22513), .B(n50781), .Z(n48292) );
  AND U42780 ( .A(n22515), .B(n22514), .Z(n48290) );
  NAND U42781 ( .A(n22517), .B(n22516), .Z(n48288) );
  AND U42782 ( .A(n22519), .B(n22518), .Z(n48286) );
  NANDN U42783 ( .A(x[7294]), .B(y[7294]), .Z(n50783) );
  NAND U42784 ( .A(n50783), .B(n22520), .Z(n48284) );
  AND U42785 ( .A(n22522), .B(n22521), .Z(n48282) );
  ANDN U42786 ( .B(y[7292]), .A(x[7292]), .Z(n50785) );
  NOR U42787 ( .A(n50785), .B(n60166), .Z(n48280) );
  AND U42788 ( .A(n22524), .B(n22523), .Z(n48272) );
  AND U42789 ( .A(n22525), .B(n60161), .Z(n48270) );
  NAND U42790 ( .A(n22527), .B(n22526), .Z(n48268) );
  AND U42791 ( .A(n22529), .B(n22528), .Z(n48266) );
  NAND U42792 ( .A(n22531), .B(n22530), .Z(n48264) );
  NANDN U42793 ( .A(x[7284]), .B(y[7284]), .Z(n60155) );
  AND U42794 ( .A(n60155), .B(n22532), .Z(n48262) );
  NAND U42795 ( .A(n22534), .B(n22533), .Z(n48260) );
  AND U42796 ( .A(n22536), .B(n22535), .Z(n48255) );
  NANDN U42797 ( .A(x[7280]), .B(y[7280]), .Z(n60151) );
  IV U42798 ( .A(n22537), .Z(n50786) );
  ANDN U42799 ( .B(n60151), .A(n50786), .Z(n48253) );
  AND U42800 ( .A(n22539), .B(n22538), .Z(n48245) );
  ANDN U42801 ( .B(y[7276]), .A(x[7276]), .Z(n50788) );
  NOR U42802 ( .A(n50788), .B(n60147), .Z(n48243) );
  AND U42803 ( .A(n22541), .B(n22540), .Z(n48235) );
  ANDN U42804 ( .B(y[7272]), .A(x[7272]), .Z(n50789) );
  NOR U42805 ( .A(n50789), .B(n60141), .Z(n48233) );
  AND U42806 ( .A(n22543), .B(n22542), .Z(n48225) );
  NANDN U42807 ( .A(x[7268]), .B(y[7268]), .Z(n50792) );
  ANDN U42808 ( .B(n50792), .A(n60137), .Z(n48223) );
  AND U42809 ( .A(n22545), .B(n22544), .Z(n48215) );
  AND U42810 ( .A(n22547), .B(n22546), .Z(n48211) );
  ANDN U42811 ( .B(y[7262]), .A(x[7262]), .Z(n48209) );
  AND U42812 ( .A(n22549), .B(n22548), .Z(n48206) );
  ANDN U42813 ( .B(y[7260]), .A(x[7260]), .Z(n60126) );
  NOR U42814 ( .A(n60126), .B(n22550), .Z(n48204) );
  AND U42815 ( .A(n22552), .B(n22551), .Z(n48196) );
  ANDN U42816 ( .B(y[7256]), .A(x[7256]), .Z(n60119) );
  NOR U42817 ( .A(n60119), .B(n60122), .Z(n48194) );
  AND U42818 ( .A(n22554), .B(n22553), .Z(n48186) );
  NANDN U42819 ( .A(x[7252]), .B(y[7252]), .Z(n50796) );
  ANDN U42820 ( .B(n50796), .A(n60116), .Z(n48184) );
  AND U42821 ( .A(n22556), .B(n22555), .Z(n48175) );
  ANDN U42822 ( .B(y[7248]), .A(x[7248]), .Z(n50798) );
  NOR U42823 ( .A(n50798), .B(n60111), .Z(n48173) );
  AND U42824 ( .A(n22558), .B(n22557), .Z(n48164) );
  NANDN U42825 ( .A(x[7244]), .B(y[7244]), .Z(n60106) );
  NAND U42826 ( .A(n60106), .B(n22559), .Z(n48162) );
  AND U42827 ( .A(n22561), .B(n22560), .Z(n48160) );
  NANDN U42828 ( .A(x[7242]), .B(y[7242]), .Z(n60103) );
  NAND U42829 ( .A(n60103), .B(n60105), .Z(n48158) );
  AND U42830 ( .A(n22563), .B(n22562), .Z(n48156) );
  NANDN U42831 ( .A(x[7240]), .B(y[7240]), .Z(n60099) );
  ANDN U42832 ( .B(n60099), .A(n60102), .Z(n48154) );
  AND U42833 ( .A(n22565), .B(n22564), .Z(n48146) );
  NANDN U42834 ( .A(x[7236]), .B(y[7236]), .Z(n60095) );
  AND U42835 ( .A(n60095), .B(n50800), .Z(n48144) );
  NAND U42836 ( .A(n22567), .B(n22566), .Z(n48142) );
  AND U42837 ( .A(n22569), .B(n22568), .Z(n48138) );
  NANDN U42838 ( .A(x[7232]), .B(y[7232]), .Z(n60091) );
  AND U42839 ( .A(n60091), .B(n22570), .Z(n48136) );
  AND U42840 ( .A(n22572), .B(n22571), .Z(n48128) );
  ANDN U42841 ( .B(y[7228]), .A(x[7228]), .Z(n50805) );
  NOR U42842 ( .A(n50805), .B(n60087), .Z(n48126) );
  AND U42843 ( .A(n22574), .B(n22573), .Z(n48118) );
  ANDN U42844 ( .B(y[7224]), .A(x[7224]), .Z(n50807) );
  NOR U42845 ( .A(n50807), .B(n60082), .Z(n48116) );
  AND U42846 ( .A(n22576), .B(n22575), .Z(n48108) );
  ANDN U42847 ( .B(y[7220]), .A(x[7220]), .Z(n50809) );
  NOR U42848 ( .A(n50809), .B(n60079), .Z(n48106) );
  AND U42849 ( .A(n22578), .B(n22577), .Z(n48097) );
  NANDN U42850 ( .A(x[7216]), .B(y[7216]), .Z(n60072) );
  ANDN U42851 ( .B(n60072), .A(n60074), .Z(n48095) );
  AND U42852 ( .A(n22580), .B(n22579), .Z(n48087) );
  NANDN U42853 ( .A(x[7212]), .B(y[7212]), .Z(n60067) );
  ANDN U42854 ( .B(n60067), .A(n60069), .Z(n48085) );
  AND U42855 ( .A(n22582), .B(n22581), .Z(n48077) );
  AND U42856 ( .A(n22584), .B(n22583), .Z(n48072) );
  NAND U42857 ( .A(n22586), .B(n22585), .Z(n48070) );
  AND U42858 ( .A(n22588), .B(n22587), .Z(n48068) );
  AND U42859 ( .A(n22590), .B(n22589), .Z(n48063) );
  IV U42860 ( .A(n22591), .Z(n60056) );
  NAND U42861 ( .A(n60056), .B(n22592), .Z(n48061) );
  AND U42862 ( .A(n22594), .B(n22593), .Z(n48059) );
  ANDN U42863 ( .B(y[7200]), .A(x[7200]), .Z(n50814) );
  NOR U42864 ( .A(n50814), .B(n22595), .Z(n48057) );
  AND U42865 ( .A(n22597), .B(n22596), .Z(n48049) );
  ANDN U42866 ( .B(y[7196]), .A(x[7196]), .Z(n50817) );
  NOR U42867 ( .A(n50817), .B(n60051), .Z(n48047) );
  AND U42868 ( .A(n22599), .B(n22598), .Z(n48039) );
  AND U42869 ( .A(n22601), .B(n22600), .Z(n48034) );
  NAND U42870 ( .A(n22603), .B(n22602), .Z(n48032) );
  AND U42871 ( .A(n22605), .B(n22604), .Z(n48030) );
  ANDN U42872 ( .B(y[7188]), .A(x[7188]), .Z(n60040) );
  NOR U42873 ( .A(n60040), .B(n22606), .Z(n48028) );
  AND U42874 ( .A(n22608), .B(n22607), .Z(n48020) );
  NANDN U42875 ( .A(x[7184]), .B(y[7184]), .Z(n60036) );
  IV U42876 ( .A(n22609), .Z(n50818) );
  ANDN U42877 ( .B(n60036), .A(n50818), .Z(n48018) );
  AND U42878 ( .A(n22611), .B(n22610), .Z(n48010) );
  NANDN U42879 ( .A(x[7180]), .B(y[7180]), .Z(n60029) );
  AND U42880 ( .A(n60029), .B(n60032), .Z(n48008) );
  NAND U42881 ( .A(n22613), .B(n22612), .Z(n48006) );
  AND U42882 ( .A(n22615), .B(n22614), .Z(n48002) );
  NANDN U42883 ( .A(x[7176]), .B(y[7176]), .Z(n50823) );
  AND U42884 ( .A(n50823), .B(n60025), .Z(n48000) );
  NANDN U42885 ( .A(x[7174]), .B(y[7174]), .Z(n60023) );
  AND U42886 ( .A(n22617), .B(n22616), .Z(n47992) );
  ANDN U42887 ( .B(y[7172]), .A(x[7172]), .Z(n50824) );
  NOR U42888 ( .A(n60022), .B(n50824), .Z(n47990) );
  AND U42889 ( .A(n22619), .B(n22618), .Z(n47981) );
  NANDN U42890 ( .A(x[7168]), .B(y[7168]), .Z(n60015) );
  ANDN U42891 ( .B(n60015), .A(n60018), .Z(n47979) );
  AND U42892 ( .A(n22621), .B(n22620), .Z(n47971) );
  NANDN U42893 ( .A(x[7164]), .B(y[7164]), .Z(n60009) );
  ANDN U42894 ( .B(n60009), .A(n60011), .Z(n47969) );
  AND U42895 ( .A(n22623), .B(n22622), .Z(n47961) );
  ANDN U42896 ( .B(y[7160]), .A(x[7160]), .Z(n22624) );
  ANDN U42897 ( .B(n60007), .A(n22624), .Z(n47959) );
  AND U42898 ( .A(n22626), .B(n22625), .Z(n47950) );
  NAND U42899 ( .A(n22628), .B(n22627), .Z(n47946) );
  AND U42900 ( .A(n22630), .B(n22629), .Z(n47942) );
  ANDN U42901 ( .B(y[7152]), .A(x[7152]), .Z(n50832) );
  NOR U42902 ( .A(n50832), .B(n59999), .Z(n47940) );
  AND U42903 ( .A(n22632), .B(n22631), .Z(n47932) );
  ANDN U42904 ( .B(y[7148]), .A(x[7148]), .Z(n50834) );
  NOR U42905 ( .A(n50834), .B(n59995), .Z(n47930) );
  AND U42906 ( .A(n22634), .B(n22633), .Z(n47922) );
  NANDN U42907 ( .A(x[7144]), .B(y[7144]), .Z(n22635) );
  NAND U42908 ( .A(n22635), .B(n50837), .Z(n47920) );
  AND U42909 ( .A(n22637), .B(n22636), .Z(n47918) );
  NANDN U42910 ( .A(x[7142]), .B(y[7142]), .Z(n50840) );
  NAND U42911 ( .A(n50840), .B(n22638), .Z(n47916) );
  XNOR U42912 ( .A(x[7142]), .B(y[7142]), .Z(n22640) );
  AND U42913 ( .A(n22640), .B(n22639), .Z(n47914) );
  ANDN U42914 ( .B(y[7140]), .A(x[7140]), .Z(n59988) );
  NOR U42915 ( .A(n59988), .B(n50839), .Z(n47912) );
  AND U42916 ( .A(n22642), .B(n22641), .Z(n47904) );
  IV U42917 ( .A(n22643), .Z(n59984) );
  ANDN U42918 ( .B(y[7136]), .A(x[7136]), .Z(n59983) );
  NOR U42919 ( .A(n59984), .B(n59983), .Z(n47902) );
  AND U42920 ( .A(n22645), .B(n22644), .Z(n47894) );
  ANDN U42921 ( .B(y[7132]), .A(x[7132]), .Z(n50842) );
  NOR U42922 ( .A(n50842), .B(n59978), .Z(n47892) );
  AND U42923 ( .A(n22647), .B(n22646), .Z(n47884) );
  ANDN U42924 ( .B(y[7128]), .A(x[7128]), .Z(n59971) );
  NOR U42925 ( .A(n59971), .B(n59973), .Z(n47882) );
  AND U42926 ( .A(n22649), .B(n22648), .Z(n47873) );
  AND U42927 ( .A(n22651), .B(n22650), .Z(n47869) );
  AND U42928 ( .A(n22653), .B(n22652), .Z(n47865) );
  NANDN U42929 ( .A(x[7120]), .B(y[7120]), .Z(n59961) );
  ANDN U42930 ( .B(n59961), .A(n59963), .Z(n47863) );
  AND U42931 ( .A(n22655), .B(n22654), .Z(n47855) );
  NANDN U42932 ( .A(x[7116]), .B(y[7116]), .Z(n59955) );
  ANDN U42933 ( .B(n59955), .A(n59957), .Z(n47853) );
  AND U42934 ( .A(n22657), .B(n22656), .Z(n47845) );
  NANDN U42935 ( .A(x[7112]), .B(y[7112]), .Z(n59950) );
  AND U42936 ( .A(n59950), .B(n59953), .Z(n47843) );
  AND U42937 ( .A(n22659), .B(n22658), .Z(n47835) );
  NANDN U42938 ( .A(x[7108]), .B(y[7108]), .Z(n59945) );
  IV U42939 ( .A(n22660), .Z(n50849) );
  ANDN U42940 ( .B(n59945), .A(n50849), .Z(n47833) );
  AND U42941 ( .A(n22662), .B(n22661), .Z(n47825) );
  ANDN U42942 ( .B(y[7104]), .A(x[7104]), .Z(n50851) );
  NOR U42943 ( .A(n50851), .B(n59941), .Z(n47823) );
  AND U42944 ( .A(n22664), .B(n22663), .Z(n47815) );
  ANDN U42945 ( .B(y[7100]), .A(x[7100]), .Z(n50853) );
  NOR U42946 ( .A(n50853), .B(n59936), .Z(n47813) );
  AND U42947 ( .A(n22666), .B(n22665), .Z(n47805) );
  ANDN U42948 ( .B(y[7096]), .A(x[7096]), .Z(n50856) );
  NOR U42949 ( .A(n50856), .B(n59931), .Z(n47803) );
  AND U42950 ( .A(n22667), .B(n50857), .Z(n47797) );
  AND U42951 ( .A(n22669), .B(n22668), .Z(n47795) );
  NANDN U42952 ( .A(x[7092]), .B(y[7092]), .Z(n59926) );
  AND U42953 ( .A(n59926), .B(n22670), .Z(n47793) );
  NAND U42954 ( .A(n22672), .B(n22671), .Z(n47791) );
  AND U42955 ( .A(n22674), .B(n22673), .Z(n47787) );
  NANDN U42956 ( .A(x[7088]), .B(y[7088]), .Z(n59921) );
  ANDN U42957 ( .B(n59921), .A(n59923), .Z(n47785) );
  AND U42958 ( .A(n22676), .B(n22675), .Z(n47777) );
  ANDN U42959 ( .B(y[7084]), .A(x[7084]), .Z(n50860) );
  ANDN U42960 ( .B(n59918), .A(n50860), .Z(n47775) );
  AND U42961 ( .A(n22678), .B(n22677), .Z(n47767) );
  NAND U42962 ( .A(n22680), .B(n22679), .Z(n47763) );
  AND U42963 ( .A(n22682), .B(n22681), .Z(n47759) );
  ANDN U42964 ( .B(y[7076]), .A(x[7076]), .Z(n50863) );
  NOR U42965 ( .A(n50863), .B(n59908), .Z(n47757) );
  AND U42966 ( .A(n22684), .B(n22683), .Z(n47749) );
  ANDN U42967 ( .B(y[7072]), .A(x[7072]), .Z(n50866) );
  NOR U42968 ( .A(n50866), .B(n59903), .Z(n47747) );
  AND U42969 ( .A(n22686), .B(n22685), .Z(n47739) );
  NANDN U42970 ( .A(x[7068]), .B(y[7068]), .Z(n59897) );
  ANDN U42971 ( .B(n59897), .A(n59899), .Z(n47737) );
  AND U42972 ( .A(n22688), .B(n22687), .Z(n47729) );
  NANDN U42973 ( .A(x[7064]), .B(y[7064]), .Z(n59890) );
  ANDN U42974 ( .B(n59890), .A(n59893), .Z(n47727) );
  AND U42975 ( .A(n22690), .B(n22689), .Z(n47719) );
  NANDN U42976 ( .A(x[7060]), .B(y[7060]), .Z(n59886) );
  NAND U42977 ( .A(n59886), .B(n50867), .Z(n47717) );
  AND U42978 ( .A(n22692), .B(n22691), .Z(n47715) );
  NANDN U42979 ( .A(x[7058]), .B(y[7058]), .Z(n22693) );
  NAND U42980 ( .A(n22693), .B(n59885), .Z(n47713) );
  AND U42981 ( .A(n22695), .B(n22694), .Z(n47711) );
  AND U42982 ( .A(n22697), .B(n22696), .Z(n47706) );
  NANDN U42983 ( .A(x[7054]), .B(y[7054]), .Z(n59878) );
  AND U42984 ( .A(n22699), .B(n22698), .Z(n47702) );
  ANDN U42985 ( .B(y[7052]), .A(x[7052]), .Z(n50870) );
  NOR U42986 ( .A(n50870), .B(n59877), .Z(n47700) );
  AND U42987 ( .A(n22701), .B(n22700), .Z(n47692) );
  AND U42988 ( .A(n22703), .B(n22702), .Z(n47688) );
  AND U42989 ( .A(n22705), .B(n22704), .Z(n47684) );
  ANDN U42990 ( .B(y[7044]), .A(x[7044]), .Z(n50872) );
  NOR U42991 ( .A(n50872), .B(n59867), .Z(n47682) );
  AND U42992 ( .A(n22707), .B(n22706), .Z(n47673) );
  NANDN U42993 ( .A(x[7040]), .B(y[7040]), .Z(n59861) );
  ANDN U42994 ( .B(n59861), .A(n22708), .Z(n47671) );
  AND U42995 ( .A(n22710), .B(n22709), .Z(n47662) );
  NANDN U42996 ( .A(x[7036]), .B(y[7036]), .Z(n59855) );
  ANDN U42997 ( .B(n59855), .A(n59857), .Z(n47660) );
  AND U42998 ( .A(n22712), .B(n22711), .Z(n47652) );
  ANDN U42999 ( .B(y[7032]), .A(x[7032]), .Z(n59852) );
  NOR U43000 ( .A(n59852), .B(n50875), .Z(n47650) );
  AND U43001 ( .A(n22714), .B(n22713), .Z(n47642) );
  NANDN U43002 ( .A(x[7028]), .B(y[7028]), .Z(n59847) );
  IV U43003 ( .A(n22715), .Z(n50877) );
  ANDN U43004 ( .B(n59847), .A(n50877), .Z(n47640) );
  AND U43005 ( .A(n22717), .B(n22716), .Z(n47632) );
  ANDN U43006 ( .B(y[7024]), .A(x[7024]), .Z(n50880) );
  NOR U43007 ( .A(n50880), .B(n59843), .Z(n47630) );
  AND U43008 ( .A(n22719), .B(n22718), .Z(n47622) );
  ANDN U43009 ( .B(y[7020]), .A(x[7020]), .Z(n50882) );
  NOR U43010 ( .A(n50882), .B(n59839), .Z(n47620) );
  AND U43011 ( .A(n22721), .B(n22720), .Z(n47612) );
  ANDN U43012 ( .B(y[7016]), .A(x[7016]), .Z(n50885) );
  NOR U43013 ( .A(n50885), .B(n59835), .Z(n47610) );
  AND U43014 ( .A(n22723), .B(n22722), .Z(n47602) );
  NANDN U43015 ( .A(x[7012]), .B(y[7012]), .Z(n59829) );
  ANDN U43016 ( .B(n59829), .A(n59831), .Z(n47600) );
  AND U43017 ( .A(n22725), .B(n22724), .Z(n47592) );
  ANDN U43018 ( .B(y[7008]), .A(x[7008]), .Z(n59822) );
  NOR U43019 ( .A(n59822), .B(n59825), .Z(n47590) );
  AND U43020 ( .A(n22727), .B(n22726), .Z(n47582) );
  NANDN U43021 ( .A(x[7004]), .B(y[7004]), .Z(n59816) );
  AND U43022 ( .A(n59816), .B(n50887), .Z(n47580) );
  NAND U43023 ( .A(n22729), .B(n22728), .Z(n47578) );
  AND U43024 ( .A(n22731), .B(n22730), .Z(n47574) );
  NANDN U43025 ( .A(x[7000]), .B(y[7000]), .Z(n59809) );
  AND U43026 ( .A(n59812), .B(n59809), .Z(n47572) );
  AND U43027 ( .A(n22732), .B(n59810), .Z(n47566) );
  NAND U43028 ( .A(n22734), .B(n22733), .Z(n47564) );
  NANDN U43029 ( .A(x[6996]), .B(y[6996]), .Z(n50890) );
  AND U43030 ( .A(n22735), .B(n50890), .Z(n47562) );
  NAND U43031 ( .A(n22737), .B(n22736), .Z(n47560) );
  AND U43032 ( .A(n22739), .B(n22738), .Z(n47556) );
  ANDN U43033 ( .B(y[6992]), .A(x[6992]), .Z(n59802) );
  NOR U43034 ( .A(n59802), .B(n50891), .Z(n47554) );
  AND U43035 ( .A(n22741), .B(n22740), .Z(n47546) );
  NANDN U43036 ( .A(x[6988]), .B(y[6988]), .Z(n59798) );
  ANDN U43037 ( .B(n59798), .A(n50893), .Z(n47544) );
  AND U43038 ( .A(n22743), .B(n22742), .Z(n47536) );
  ANDN U43039 ( .B(y[6984]), .A(x[6984]), .Z(n50895) );
  NOR U43040 ( .A(n50895), .B(n59794), .Z(n47534) );
  AND U43041 ( .A(n22745), .B(n22744), .Z(n47526) );
  ANDN U43042 ( .B(y[6980]), .A(x[6980]), .Z(n50896) );
  NOR U43043 ( .A(n50896), .B(n59787), .Z(n47524) );
  AND U43044 ( .A(n22747), .B(n22746), .Z(n47516) );
  NAND U43045 ( .A(n22749), .B(n22748), .Z(n47512) );
  NANDN U43046 ( .A(x[6974]), .B(y[6974]), .Z(n59780) );
  AND U43047 ( .A(n22751), .B(n22750), .Z(n47508) );
  NANDN U43048 ( .A(x[6972]), .B(y[6972]), .Z(n59776) );
  ANDN U43049 ( .B(n59776), .A(n59779), .Z(n47506) );
  AND U43050 ( .A(n22753), .B(n22752), .Z(n47498) );
  NANDN U43051 ( .A(x[6968]), .B(y[6968]), .Z(n59770) );
  ANDN U43052 ( .B(n59770), .A(n59772), .Z(n47496) );
  AND U43053 ( .A(n22755), .B(n22754), .Z(n47488) );
  ANDN U43054 ( .B(y[6964]), .A(x[6964]), .Z(n59766) );
  NOR U43055 ( .A(n59766), .B(n50900), .Z(n47486) );
  AND U43056 ( .A(n22757), .B(n22756), .Z(n47478) );
  ANDN U43057 ( .B(y[6960]), .A(x[6960]), .Z(n50905) );
  NOR U43058 ( .A(n50905), .B(n50903), .Z(n47476) );
  AND U43059 ( .A(n22759), .B(n22758), .Z(n47468) );
  ANDN U43060 ( .B(y[6956]), .A(x[6956]), .Z(n22760) );
  NOR U43061 ( .A(n22760), .B(n59760), .Z(n47466) );
  AND U43062 ( .A(n22762), .B(n22761), .Z(n47457) );
  ANDN U43063 ( .B(y[6952]), .A(x[6952]), .Z(n50908) );
  NOR U43064 ( .A(n50908), .B(n59755), .Z(n47455) );
  AND U43065 ( .A(n22764), .B(n22763), .Z(n47447) );
  NANDN U43066 ( .A(x[6948]), .B(y[6948]), .Z(n59748) );
  ANDN U43067 ( .B(n59748), .A(n59751), .Z(n47445) );
  AND U43068 ( .A(n22766), .B(n22765), .Z(n47437) );
  NANDN U43069 ( .A(x[6944]), .B(y[6944]), .Z(n59742) );
  ANDN U43070 ( .B(n59742), .A(n59744), .Z(n47435) );
  AND U43071 ( .A(n22768), .B(n22767), .Z(n47427) );
  ANDN U43072 ( .B(y[6940]), .A(x[6940]), .Z(n22769) );
  ANDN U43073 ( .B(n59739), .A(n22769), .Z(n47425) );
  AND U43074 ( .A(n22771), .B(n22770), .Z(n47416) );
  ANDN U43075 ( .B(y[6936]), .A(x[6936]), .Z(n59732) );
  NOR U43076 ( .A(n59732), .B(n50910), .Z(n47414) );
  AND U43077 ( .A(n22773), .B(n22772), .Z(n47406) );
  ANDN U43078 ( .B(y[6932]), .A(x[6932]), .Z(n50912) );
  NOR U43079 ( .A(n50912), .B(n59727), .Z(n47404) );
  AND U43080 ( .A(n22775), .B(n22774), .Z(n47396) );
  NAND U43081 ( .A(n22777), .B(n22776), .Z(n47392) );
  AND U43082 ( .A(n22779), .B(n22778), .Z(n47388) );
  ANDN U43083 ( .B(y[6924]), .A(x[6924]), .Z(n50916) );
  NOR U43084 ( .A(n50916), .B(n59719), .Z(n47386) );
  AND U43085 ( .A(n22781), .B(n22780), .Z(n47378) );
  NANDN U43086 ( .A(x[6920]), .B(y[6920]), .Z(n59712) );
  ANDN U43087 ( .B(n59712), .A(n59714), .Z(n47376) );
  AND U43088 ( .A(n22783), .B(n22782), .Z(n47368) );
  ANDN U43089 ( .B(y[6916]), .A(x[6916]), .Z(n59706) );
  NOR U43090 ( .A(n59706), .B(n59708), .Z(n47366) );
  AND U43091 ( .A(n22785), .B(n22784), .Z(n47358) );
  ANDN U43092 ( .B(y[6912]), .A(x[6912]), .Z(n59700) );
  NOR U43093 ( .A(n59700), .B(n50918), .Z(n47356) );
  AND U43094 ( .A(n22787), .B(n22786), .Z(n47348) );
  ANDN U43095 ( .B(y[6908]), .A(x[6908]), .Z(n59694) );
  NOR U43096 ( .A(n59694), .B(n59696), .Z(n47346) );
  AND U43097 ( .A(n22789), .B(n22788), .Z(n47337) );
  NANDN U43098 ( .A(x[6904]), .B(y[6904]), .Z(n59691) );
  IV U43099 ( .A(n22790), .Z(n50921) );
  ANDN U43100 ( .B(n59691), .A(n50921), .Z(n47335) );
  AND U43101 ( .A(n22791), .B(n59690), .Z(n47329) );
  AND U43102 ( .A(n22793), .B(n22792), .Z(n47327) );
  ANDN U43103 ( .B(y[6900]), .A(x[6900]), .Z(n59684) );
  NOR U43104 ( .A(n59684), .B(n22794), .Z(n47325) );
  AND U43105 ( .A(n22796), .B(n22795), .Z(n47317) );
  ANDN U43106 ( .B(y[6896]), .A(x[6896]), .Z(n59680) );
  NOR U43107 ( .A(n59680), .B(n50923), .Z(n47315) );
  AND U43108 ( .A(n22798), .B(n22797), .Z(n47307) );
  ANDN U43109 ( .B(y[6892]), .A(x[6892]), .Z(n50925) );
  NOR U43110 ( .A(n50925), .B(n59676), .Z(n47305) );
  AND U43111 ( .A(n22800), .B(n22799), .Z(n47297) );
  NANDN U43112 ( .A(x[6888]), .B(y[6888]), .Z(n50928) );
  ANDN U43113 ( .B(n50928), .A(n59671), .Z(n47295) );
  AND U43114 ( .A(n22802), .B(n22801), .Z(n47286) );
  ANDN U43115 ( .B(y[6884]), .A(x[6884]), .Z(n50929) );
  NOR U43116 ( .A(n50929), .B(n59666), .Z(n47284) );
  AND U43117 ( .A(n22804), .B(n22803), .Z(n47275) );
  NANDN U43118 ( .A(x[6880]), .B(y[6880]), .Z(n59660) );
  ANDN U43119 ( .B(n59660), .A(n59662), .Z(n47273) );
  AND U43120 ( .A(n22806), .B(n22805), .Z(n47265) );
  NANDN U43121 ( .A(x[6876]), .B(y[6876]), .Z(n59653) );
  AND U43122 ( .A(n59653), .B(n59656), .Z(n47263) );
  NAND U43123 ( .A(n22808), .B(n22807), .Z(n47261) );
  AND U43124 ( .A(n22810), .B(n22809), .Z(n47257) );
  NANDN U43125 ( .A(x[6872]), .B(y[6872]), .Z(n59649) );
  AND U43126 ( .A(n59649), .B(n50931), .Z(n47255) );
  ANDN U43127 ( .B(y[6870]), .A(x[6870]), .Z(n50933) );
  AND U43128 ( .A(n22812), .B(n22811), .Z(n47247) );
  ANDN U43129 ( .B(y[6868]), .A(x[6868]), .Z(n59645) );
  ANDN U43130 ( .B(n50934), .A(n59645), .Z(n47245) );
  AND U43131 ( .A(n22814), .B(n22813), .Z(n47237) );
  NANDN U43132 ( .A(x[6864]), .B(y[6864]), .Z(n59638) );
  AND U43133 ( .A(n59638), .B(n59641), .Z(n47235) );
  NAND U43134 ( .A(n22816), .B(n22815), .Z(n47233) );
  AND U43135 ( .A(n22818), .B(n22817), .Z(n47229) );
  ANDN U43136 ( .B(y[6860]), .A(x[6860]), .Z(n50935) );
  NOR U43137 ( .A(n50935), .B(n59634), .Z(n47227) );
  AND U43138 ( .A(n22820), .B(n22819), .Z(n47219) );
  NANDN U43139 ( .A(x[6856]), .B(y[6856]), .Z(n50938) );
  NAND U43140 ( .A(n50938), .B(n59630), .Z(n47217) );
  AND U43141 ( .A(n22822), .B(n22821), .Z(n47215) );
  NANDN U43142 ( .A(x[6854]), .B(y[6854]), .Z(n22823) );
  NAND U43143 ( .A(n22823), .B(n50937), .Z(n47213) );
  AND U43144 ( .A(n22825), .B(n22824), .Z(n47211) );
  NAND U43145 ( .A(n22827), .B(n22826), .Z(n47206) );
  AND U43146 ( .A(n22829), .B(n22828), .Z(n47202) );
  NANDN U43147 ( .A(x[6848]), .B(y[6848]), .Z(n59618) );
  ANDN U43148 ( .B(n59618), .A(n59620), .Z(n47200) );
  AND U43149 ( .A(n22831), .B(n22830), .Z(n47192) );
  NANDN U43150 ( .A(x[6844]), .B(y[6844]), .Z(n59615) );
  AND U43151 ( .A(n59615), .B(n50940), .Z(n47190) );
  NAND U43152 ( .A(n22833), .B(n22832), .Z(n47188) );
  NANDN U43153 ( .A(x[6842]), .B(y[6842]), .Z(n50942) );
  AND U43154 ( .A(n50942), .B(n59614), .Z(n47186) );
  AND U43155 ( .A(n22835), .B(n22834), .Z(n47184) );
  ANDN U43156 ( .B(y[6840]), .A(x[6840]), .Z(n50945) );
  NOR U43157 ( .A(n50945), .B(n50943), .Z(n47182) );
  AND U43158 ( .A(n22837), .B(n22836), .Z(n47173) );
  NANDN U43159 ( .A(x[6836]), .B(y[6836]), .Z(n50948) );
  ANDN U43160 ( .B(n50948), .A(n22838), .Z(n47171) );
  AND U43161 ( .A(n22840), .B(n22839), .Z(n47162) );
  ANDN U43162 ( .B(y[6832]), .A(x[6832]), .Z(n50949) );
  NOR U43163 ( .A(n50949), .B(n59605), .Z(n47160) );
  AND U43164 ( .A(n22842), .B(n22841), .Z(n47151) );
  NANDN U43165 ( .A(x[6828]), .B(y[6828]), .Z(n59599) );
  ANDN U43166 ( .B(n59599), .A(n59601), .Z(n47149) );
  AND U43167 ( .A(n22844), .B(n22843), .Z(n47141) );
  ANDN U43168 ( .B(y[6824]), .A(x[6824]), .Z(n59592) );
  NOR U43169 ( .A(n59592), .B(n59594), .Z(n47139) );
  AND U43170 ( .A(n22846), .B(n22845), .Z(n47131) );
  NANDN U43171 ( .A(x[6820]), .B(y[6820]), .Z(n59588) );
  IV U43172 ( .A(n22847), .Z(n50951) );
  ANDN U43173 ( .B(n59588), .A(n50951), .Z(n47129) );
  AND U43174 ( .A(n22849), .B(n22848), .Z(n47121) );
  NANDN U43175 ( .A(x[6816]), .B(y[6816]), .Z(n59582) );
  AND U43176 ( .A(n59582), .B(n59584), .Z(n47119) );
  NAND U43177 ( .A(n22851), .B(n22850), .Z(n47117) );
  AND U43178 ( .A(n22853), .B(n22852), .Z(n47113) );
  ANDN U43179 ( .B(y[6812]), .A(x[6812]), .Z(n59575) );
  NOR U43180 ( .A(n59575), .B(n59577), .Z(n47111) );
  AND U43181 ( .A(n22855), .B(n22854), .Z(n47103) );
  ANDN U43182 ( .B(n22856), .A(n59571), .Z(n47101) );
  NANDN U43183 ( .A(x[6804]), .B(y[6804]), .Z(n59566) );
  ANDN U43184 ( .B(n59566), .A(n22857), .Z(n47090) );
  AND U43185 ( .A(n22859), .B(n22858), .Z(n47082) );
  NANDN U43186 ( .A(x[6800]), .B(y[6800]), .Z(n59559) );
  ANDN U43187 ( .B(n59559), .A(n59561), .Z(n47080) );
  AND U43188 ( .A(n22861), .B(n22860), .Z(n47072) );
  ANDN U43189 ( .B(y[6796]), .A(x[6796]), .Z(n59555) );
  NOR U43190 ( .A(n59555), .B(n50954), .Z(n47070) );
  AND U43191 ( .A(n22863), .B(n22862), .Z(n47062) );
  AND U43192 ( .A(n22865), .B(n22864), .Z(n47058) );
  AND U43193 ( .A(n22867), .B(n22866), .Z(n47054) );
  ANDN U43194 ( .B(y[6788]), .A(x[6788]), .Z(n50958) );
  NOR U43195 ( .A(n50958), .B(n59545), .Z(n47052) );
  AND U43196 ( .A(n22869), .B(n22868), .Z(n47044) );
  ANDN U43197 ( .B(y[6784]), .A(x[6784]), .Z(n50959) );
  NOR U43198 ( .A(n50959), .B(n59540), .Z(n47042) );
  AND U43199 ( .A(n22871), .B(n22870), .Z(n47034) );
  ANDN U43200 ( .B(y[6780]), .A(x[6780]), .Z(n50961) );
  NOR U43201 ( .A(n50961), .B(n59536), .Z(n47032) );
  AND U43202 ( .A(n22873), .B(n22872), .Z(n47024) );
  NANDN U43203 ( .A(x[6776]), .B(y[6776]), .Z(n59528) );
  ANDN U43204 ( .B(n59528), .A(n59530), .Z(n47022) );
  AND U43205 ( .A(n22875), .B(n22874), .Z(n47014) );
  NAND U43206 ( .A(n22877), .B(n22876), .Z(n47010) );
  NANDN U43207 ( .A(x[6770]), .B(y[6770]), .Z(n50964) );
  AND U43208 ( .A(n22879), .B(n22878), .Z(n47006) );
  ANDN U43209 ( .B(y[6768]), .A(x[6768]), .Z(n59518) );
  NOR U43210 ( .A(n59518), .B(n50963), .Z(n47004) );
  AND U43211 ( .A(n22881), .B(n22880), .Z(n46996) );
  NANDN U43212 ( .A(x[6764]), .B(y[6764]), .Z(n59513) );
  IV U43213 ( .A(n22882), .Z(n50965) );
  ANDN U43214 ( .B(n59513), .A(n50965), .Z(n46994) );
  AND U43215 ( .A(n22884), .B(n22883), .Z(n46986) );
  ANDN U43216 ( .B(y[6760]), .A(x[6760]), .Z(n50967) );
  NOR U43217 ( .A(n50967), .B(n59509), .Z(n46984) );
  AND U43218 ( .A(n22886), .B(n22885), .Z(n46976) );
  ANDN U43219 ( .B(y[6756]), .A(x[6756]), .Z(n50968) );
  NOR U43220 ( .A(n50968), .B(n59504), .Z(n46974) );
  AND U43221 ( .A(n22888), .B(n22887), .Z(n46966) );
  NANDN U43222 ( .A(x[6752]), .B(y[6752]), .Z(n22889) );
  NAND U43223 ( .A(n22889), .B(n59498), .Z(n46964) );
  AND U43224 ( .A(n22891), .B(n22890), .Z(n46962) );
  NANDN U43225 ( .A(x[6750]), .B(y[6750]), .Z(n59494) );
  NAND U43226 ( .A(n59494), .B(n22892), .Z(n46960) );
  AND U43227 ( .A(n22894), .B(n22893), .Z(n46958) );
  NANDN U43228 ( .A(x[6748]), .B(y[6748]), .Z(n59491) );
  ANDN U43229 ( .B(n59491), .A(n59493), .Z(n46956) );
  AND U43230 ( .A(n22896), .B(n22895), .Z(n46948) );
  NANDN U43231 ( .A(x[6744]), .B(y[6744]), .Z(n59484) );
  AND U43232 ( .A(n59484), .B(n59488), .Z(n46946) );
  AND U43233 ( .A(n22898), .B(n22897), .Z(n46938) );
  NANDN U43234 ( .A(x[6740]), .B(y[6740]), .Z(n59480) );
  IV U43235 ( .A(n22899), .Z(n50970) );
  ANDN U43236 ( .B(n59480), .A(n50970), .Z(n46936) );
  AND U43237 ( .A(n22901), .B(n22900), .Z(n46928) );
  NANDN U43238 ( .A(x[6736]), .B(y[6736]), .Z(n22902) );
  AND U43239 ( .A(n22902), .B(n59476), .Z(n46926) );
  NAND U43240 ( .A(n22904), .B(n22903), .Z(n46924) );
  AND U43241 ( .A(n22906), .B(n22905), .Z(n46919) );
  ANDN U43242 ( .B(y[6732]), .A(x[6732]), .Z(n50974) );
  NOR U43243 ( .A(n50974), .B(n59471), .Z(n46917) );
  AND U43244 ( .A(n22908), .B(n22907), .Z(n46909) );
  NANDN U43245 ( .A(x[6728]), .B(y[6728]), .Z(n59465) );
  ANDN U43246 ( .B(n59465), .A(n59467), .Z(n46907) );
  AND U43247 ( .A(n22910), .B(n22909), .Z(n46899) );
  NAND U43248 ( .A(n22912), .B(n22911), .Z(n46895) );
  AND U43249 ( .A(n22914), .B(n22913), .Z(n46891) );
  ANDN U43250 ( .B(y[6720]), .A(x[6720]), .Z(n59455) );
  NOR U43251 ( .A(n59455), .B(n50976), .Z(n46889) );
  IV U43252 ( .A(n22915), .Z(n59454) );
  AND U43253 ( .A(n22916), .B(n59454), .Z(n46883) );
  AND U43254 ( .A(n22918), .B(n22917), .Z(n46881) );
  NANDN U43255 ( .A(x[6716]), .B(y[6716]), .Z(n50979) );
  NAND U43256 ( .A(n50979), .B(n22919), .Z(n46879) );
  AND U43257 ( .A(n22921), .B(n22920), .Z(n46877) );
  NANDN U43258 ( .A(x[6714]), .B(y[6714]), .Z(n59448) );
  NAND U43259 ( .A(n59448), .B(n50978), .Z(n46875) );
  AND U43260 ( .A(n22923), .B(n22922), .Z(n46873) );
  ANDN U43261 ( .B(y[6712]), .A(x[6712]), .Z(n50980) );
  NOR U43262 ( .A(n50980), .B(n59447), .Z(n46871) );
  AND U43263 ( .A(n22925), .B(n22924), .Z(n46863) );
  ANDN U43264 ( .B(y[6708]), .A(x[6708]), .Z(n50983) );
  NOR U43265 ( .A(n50983), .B(n59443), .Z(n46861) );
  AND U43266 ( .A(n22927), .B(n22926), .Z(n46853) );
  NANDN U43267 ( .A(x[6704]), .B(y[6704]), .Z(n59436) );
  ANDN U43268 ( .B(n59436), .A(n59438), .Z(n46851) );
  AND U43269 ( .A(n22929), .B(n22928), .Z(n46843) );
  NANDN U43270 ( .A(x[6700]), .B(y[6700]), .Z(n59430) );
  ANDN U43271 ( .B(n59430), .A(n59432), .Z(n46841) );
  AND U43272 ( .A(n22931), .B(n22930), .Z(n46833) );
  NANDN U43273 ( .A(x[6696]), .B(y[6696]), .Z(n59424) );
  AND U43274 ( .A(n59424), .B(n59428), .Z(n46831) );
  AND U43275 ( .A(n22933), .B(n22932), .Z(n46823) );
  ANDN U43276 ( .B(y[6692]), .A(x[6692]), .Z(n59420) );
  NOR U43277 ( .A(n59420), .B(n50985), .Z(n46821) );
  AND U43278 ( .A(n22935), .B(n22934), .Z(n46813) );
  NANDN U43279 ( .A(x[6688]), .B(y[6688]), .Z(n50990) );
  AND U43280 ( .A(n50990), .B(n50987), .Z(n46811) );
  NAND U43281 ( .A(n22937), .B(n22936), .Z(n46809) );
  AND U43282 ( .A(n22939), .B(n22938), .Z(n46805) );
  ANDN U43283 ( .B(y[6684]), .A(x[6684]), .Z(n50991) );
  NOR U43284 ( .A(n50991), .B(n59414), .Z(n46803) );
  AND U43285 ( .A(n22941), .B(n22940), .Z(n46795) );
  NANDN U43286 ( .A(x[6680]), .B(y[6680]), .Z(n50994) );
  AND U43287 ( .A(n59408), .B(n50994), .Z(n46793) );
  NAND U43288 ( .A(n22943), .B(n22942), .Z(n46791) );
  AND U43289 ( .A(n22945), .B(n22944), .Z(n46787) );
  NANDN U43290 ( .A(x[6676]), .B(y[6676]), .Z(n59402) );
  NAND U43291 ( .A(n59402), .B(n59404), .Z(n46785) );
  AND U43292 ( .A(n22947), .B(n22946), .Z(n46783) );
  NAND U43293 ( .A(n22948), .B(n59401), .Z(n46781) );
  AND U43294 ( .A(n22950), .B(n22949), .Z(n46779) );
  NAND U43295 ( .A(n22952), .B(n22951), .Z(n46777) );
  AND U43296 ( .A(n22954), .B(n22953), .Z(n46775) );
  NANDN U43297 ( .A(x[6670]), .B(y[6670]), .Z(n50996) );
  NAND U43298 ( .A(n50996), .B(n22955), .Z(n46773) );
  AND U43299 ( .A(n22957), .B(n22956), .Z(n46771) );
  ANDN U43300 ( .B(y[6668]), .A(x[6668]), .Z(n50997) );
  NOR U43301 ( .A(n50997), .B(n50995), .Z(n46769) );
  AND U43302 ( .A(n22959), .B(n22958), .Z(n46761) );
  NANDN U43303 ( .A(x[6664]), .B(y[6664]), .Z(n51001) );
  ANDN U43304 ( .B(n51001), .A(n59391), .Z(n46759) );
  AND U43305 ( .A(n22961), .B(n22960), .Z(n46750) );
  ANDN U43306 ( .B(y[6660]), .A(x[6660]), .Z(n51003) );
  NOR U43307 ( .A(n51003), .B(n59388), .Z(n46748) );
  AND U43308 ( .A(n22963), .B(n22962), .Z(n46740) );
  NANDN U43309 ( .A(x[6656]), .B(y[6656]), .Z(n59380) );
  ANDN U43310 ( .B(n59380), .A(n59382), .Z(n46738) );
  AND U43311 ( .A(n22964), .B(n59379), .Z(n46732) );
  AND U43312 ( .A(n22966), .B(n22965), .Z(n46730) );
  NAND U43313 ( .A(n22968), .B(n22967), .Z(n46728) );
  AND U43314 ( .A(n22970), .B(n22969), .Z(n46726) );
  NANDN U43315 ( .A(x[6650]), .B(y[6650]), .Z(n22972) );
  NAND U43316 ( .A(n22972), .B(n22971), .Z(n46724) );
  AND U43317 ( .A(n22974), .B(n22973), .Z(n46722) );
  ANDN U43318 ( .B(y[6648]), .A(x[6648]), .Z(n51006) );
  NOR U43319 ( .A(n51006), .B(n22975), .Z(n46720) );
  AND U43320 ( .A(n22977), .B(n22976), .Z(n46712) );
  ANDN U43321 ( .B(y[6644]), .A(x[6644]), .Z(n51008) );
  NOR U43322 ( .A(n51008), .B(n59370), .Z(n46710) );
  AND U43323 ( .A(n22979), .B(n22978), .Z(n46702) );
  ANDN U43324 ( .B(y[6640]), .A(x[6640]), .Z(n51011) );
  NOR U43325 ( .A(n59365), .B(n51011), .Z(n46700) );
  AND U43326 ( .A(n22981), .B(n22980), .Z(n46692) );
  AND U43327 ( .A(n22983), .B(n22982), .Z(n46688) );
  AND U43328 ( .A(n22985), .B(n22984), .Z(n46683) );
  NAND U43329 ( .A(n22987), .B(n22986), .Z(n46681) );
  AND U43330 ( .A(n22989), .B(n22988), .Z(n46679) );
  NANDN U43331 ( .A(x[6630]), .B(y[6630]), .Z(n51013) );
  NAND U43332 ( .A(n51013), .B(n22990), .Z(n46677) );
  AND U43333 ( .A(n22992), .B(n22991), .Z(n46675) );
  NAND U43334 ( .A(n22993), .B(n51012), .Z(n46673) );
  AND U43335 ( .A(n22995), .B(n22994), .Z(n46671) );
  NANDN U43336 ( .A(x[6626]), .B(y[6626]), .Z(n59348) );
  AND U43337 ( .A(n22997), .B(n22996), .Z(n46666) );
  IV U43338 ( .A(n22998), .Z(n59347) );
  NAND U43339 ( .A(n59347), .B(n22999), .Z(n46664) );
  AND U43340 ( .A(n23001), .B(n23000), .Z(n46662) );
  NAND U43341 ( .A(n23003), .B(n23002), .Z(n46660) );
  AND U43342 ( .A(n23005), .B(n23004), .Z(n46658) );
  NANDN U43343 ( .A(x[6620]), .B(y[6620]), .Z(n59342) );
  NAND U43344 ( .A(n59342), .B(n23006), .Z(n46656) );
  AND U43345 ( .A(n23008), .B(n23007), .Z(n46654) );
  IV U43346 ( .A(n23009), .Z(n59341) );
  NANDN U43347 ( .A(x[6618]), .B(y[6618]), .Z(n59338) );
  NAND U43348 ( .A(n59341), .B(n59338), .Z(n46652) );
  AND U43349 ( .A(n23011), .B(n23010), .Z(n46650) );
  NANDN U43350 ( .A(x[6616]), .B(y[6616]), .Z(n59335) );
  ANDN U43351 ( .B(n59335), .A(n59337), .Z(n46648) );
  AND U43352 ( .A(n23013), .B(n23012), .Z(n46640) );
  ANDN U43353 ( .B(y[6612]), .A(x[6612]), .Z(n59332) );
  NOR U43354 ( .A(n59332), .B(n51016), .Z(n46638) );
  AND U43355 ( .A(n23015), .B(n23014), .Z(n46630) );
  NANDN U43356 ( .A(x[6608]), .B(y[6608]), .Z(n59328) );
  IV U43357 ( .A(n23016), .Z(n51018) );
  ANDN U43358 ( .B(n59328), .A(n51018), .Z(n46628) );
  NANDN U43359 ( .A(x[6606]), .B(y[6606]), .Z(n59324) );
  IV U43360 ( .A(n23017), .Z(n59326) );
  AND U43361 ( .A(n23019), .B(n23018), .Z(n46620) );
  NAND U43362 ( .A(n23021), .B(n23020), .Z(n46616) );
  AND U43363 ( .A(n23023), .B(n23022), .Z(n46612) );
  NAND U43364 ( .A(n23025), .B(n23024), .Z(n46608) );
  AND U43365 ( .A(n23027), .B(n23026), .Z(n46604) );
  NAND U43366 ( .A(n23029), .B(n23028), .Z(n46600) );
  AND U43367 ( .A(n23031), .B(n23030), .Z(n46596) );
  NAND U43368 ( .A(n23033), .B(n23032), .Z(n46592) );
  AND U43369 ( .A(n23035), .B(n23034), .Z(n46588) );
  NAND U43370 ( .A(n23037), .B(n23036), .Z(n46584) );
  AND U43371 ( .A(n23039), .B(n23038), .Z(n46580) );
  NANDN U43372 ( .A(x[6582]), .B(y[6582]), .Z(n59292) );
  AND U43373 ( .A(n59292), .B(n51025), .Z(n46572) );
  NAND U43374 ( .A(n23041), .B(n23040), .Z(n46570) );
  NAND U43375 ( .A(n23043), .B(n23042), .Z(n46566) );
  AND U43376 ( .A(n23045), .B(n23044), .Z(n46562) );
  NAND U43377 ( .A(n23047), .B(n23046), .Z(n46545) );
  NANDN U43378 ( .A(x[6570]), .B(y[6570]), .Z(n59274) );
  AND U43379 ( .A(n23049), .B(n23048), .Z(n46541) );
  NAND U43380 ( .A(n23051), .B(n23050), .Z(n46537) );
  NANDN U43381 ( .A(x[6566]), .B(y[6566]), .Z(n59271) );
  AND U43382 ( .A(n59271), .B(n23052), .Z(n46535) );
  NAND U43383 ( .A(n23054), .B(n23053), .Z(n46533) );
  IV U43384 ( .A(n23055), .Z(n59270) );
  AND U43385 ( .A(n23056), .B(n59270), .Z(n46531) );
  AND U43386 ( .A(n23058), .B(n23057), .Z(n46529) );
  AND U43387 ( .A(n23060), .B(n23059), .Z(n46523) );
  NAND U43388 ( .A(n23062), .B(n23061), .Z(n46518) );
  AND U43389 ( .A(n23064), .B(n23063), .Z(n46514) );
  NANDN U43390 ( .A(x[6554]), .B(y[6554]), .Z(n59257) );
  AND U43391 ( .A(n59257), .B(n51032), .Z(n46506) );
  NAND U43392 ( .A(n23066), .B(n23065), .Z(n46504) );
  NAND U43393 ( .A(n23068), .B(n23067), .Z(n46500) );
  NANDN U43394 ( .A(x[6550]), .B(y[6550]), .Z(n59250) );
  AND U43395 ( .A(n59253), .B(n59250), .Z(n46498) );
  NAND U43396 ( .A(n23070), .B(n23069), .Z(n46496) );
  NAND U43397 ( .A(n23072), .B(n23071), .Z(n46491) );
  NANDN U43398 ( .A(x[6546]), .B(y[6546]), .Z(n51034) );
  AND U43399 ( .A(n23074), .B(n23073), .Z(n46486) );
  NAND U43400 ( .A(n23076), .B(n23075), .Z(n46482) );
  NANDN U43401 ( .A(x[6542]), .B(y[6542]), .Z(n51037) );
  AND U43402 ( .A(n23078), .B(n23077), .Z(n46477) );
  NAND U43403 ( .A(n23080), .B(n23079), .Z(n46473) );
  NANDN U43404 ( .A(x[6538]), .B(y[6538]), .Z(n59237) );
  AND U43405 ( .A(n23082), .B(n23081), .Z(n46469) );
  NAND U43406 ( .A(n23084), .B(n23083), .Z(n46465) );
  NANDN U43407 ( .A(x[6534]), .B(y[6534]), .Z(n51040) );
  AND U43408 ( .A(n23086), .B(n23085), .Z(n46461) );
  AND U43409 ( .A(n23088), .B(n23087), .Z(n46456) );
  NAND U43410 ( .A(n23090), .B(n23089), .Z(n46454) );
  AND U43411 ( .A(n23092), .B(n23091), .Z(n46452) );
  NAND U43412 ( .A(n23094), .B(n23093), .Z(n46447) );
  AND U43413 ( .A(n23096), .B(n23095), .Z(n46443) );
  NAND U43414 ( .A(n23098), .B(n23097), .Z(n46439) );
  NANDN U43415 ( .A(x[6522]), .B(y[6522]), .Z(n59217) );
  AND U43416 ( .A(n23100), .B(n23099), .Z(n46435) );
  NAND U43417 ( .A(n23102), .B(n23101), .Z(n46431) );
  AND U43418 ( .A(n23104), .B(n23103), .Z(n46427) );
  NAND U43419 ( .A(n23106), .B(n23105), .Z(n46423) );
  NANDN U43420 ( .A(x[6514]), .B(y[6514]), .Z(n59207) );
  AND U43421 ( .A(n23108), .B(n23107), .Z(n46419) );
  NAND U43422 ( .A(n23110), .B(n23109), .Z(n46415) );
  AND U43423 ( .A(n23112), .B(n23111), .Z(n46411) );
  NAND U43424 ( .A(n23114), .B(n23113), .Z(n46406) );
  AND U43425 ( .A(n23116), .B(n23115), .Z(n46402) );
  AND U43426 ( .A(n23118), .B(n23117), .Z(n46392) );
  NAND U43427 ( .A(n23120), .B(n23119), .Z(n46388) );
  AND U43428 ( .A(n23122), .B(n23121), .Z(n46384) );
  NAND U43429 ( .A(n23124), .B(n23123), .Z(n46380) );
  AND U43430 ( .A(n23126), .B(n23125), .Z(n46376) );
  NAND U43431 ( .A(n23128), .B(n23127), .Z(n46372) );
  AND U43432 ( .A(n23130), .B(n23129), .Z(n46368) );
  NAND U43433 ( .A(n23132), .B(n23131), .Z(n46364) );
  AND U43434 ( .A(n23134), .B(n23133), .Z(n46360) );
  NAND U43435 ( .A(n23136), .B(n23135), .Z(n46356) );
  AND U43436 ( .A(n23138), .B(n23137), .Z(n46352) );
  NANDN U43437 ( .A(x[6478]), .B(y[6478]), .Z(n59143) );
  AND U43438 ( .A(n59143), .B(n23139), .Z(n46344) );
  NAND U43439 ( .A(n23141), .B(n23140), .Z(n46342) );
  NAND U43440 ( .A(n23143), .B(n23142), .Z(n46338) );
  NANDN U43441 ( .A(x[6474]), .B(y[6474]), .Z(n59132) );
  AND U43442 ( .A(n23145), .B(n23144), .Z(n46334) );
  AND U43443 ( .A(n23147), .B(n23146), .Z(n46323) );
  NAND U43444 ( .A(n23149), .B(n23148), .Z(n46319) );
  NANDN U43445 ( .A(x[6466]), .B(y[6466]), .Z(n59122) );
  AND U43446 ( .A(n23151), .B(n23150), .Z(n46315) );
  NAND U43447 ( .A(n23153), .B(n23152), .Z(n46311) );
  NANDN U43448 ( .A(x[6462]), .B(y[6462]), .Z(n59118) );
  IV U43449 ( .A(n23154), .Z(n51058) );
  AND U43450 ( .A(n23156), .B(n23155), .Z(n46307) );
  NAND U43451 ( .A(n23158), .B(n23157), .Z(n46303) );
  NANDN U43452 ( .A(x[6458]), .B(y[6458]), .Z(n59111) );
  AND U43453 ( .A(n23160), .B(n23159), .Z(n46299) );
  AND U43454 ( .A(n23161), .B(n59112), .Z(n46297) );
  NAND U43455 ( .A(n23163), .B(n23162), .Z(n46295) );
  AND U43456 ( .A(n23165), .B(n23164), .Z(n46293) );
  NAND U43457 ( .A(n23167), .B(n23166), .Z(n46291) );
  NANDN U43458 ( .A(x[6450]), .B(y[6450]), .Z(n51061) );
  AND U43459 ( .A(n23169), .B(n23168), .Z(n46280) );
  NAND U43460 ( .A(n23171), .B(n23170), .Z(n46275) );
  NANDN U43461 ( .A(x[6446]), .B(y[6446]), .Z(n23172) );
  AND U43462 ( .A(n23172), .B(n59097), .Z(n46273) );
  NAND U43463 ( .A(n23174), .B(n23173), .Z(n46271) );
  AND U43464 ( .A(n23176), .B(n23175), .Z(n46269) );
  NAND U43465 ( .A(n23178), .B(n23177), .Z(n46267) );
  NANDN U43466 ( .A(x[6442]), .B(y[6442]), .Z(n59091) );
  AND U43467 ( .A(n23180), .B(n23179), .Z(n46262) );
  NAND U43468 ( .A(n23182), .B(n23181), .Z(n46258) );
  IV U43469 ( .A(n23183), .Z(n59087) );
  AND U43470 ( .A(n23184), .B(n59087), .Z(n46256) );
  AND U43471 ( .A(n59085), .B(n23185), .Z(n46246) );
  AND U43472 ( .A(n23187), .B(n23186), .Z(n46244) );
  AND U43473 ( .A(n23189), .B(n23188), .Z(n46242) );
  NANDN U43474 ( .A(x[6432]), .B(y[6432]), .Z(n51066) );
  AND U43475 ( .A(n51066), .B(n23190), .Z(n46240) );
  NAND U43476 ( .A(n23192), .B(n23191), .Z(n46238) );
  AND U43477 ( .A(n23194), .B(n23193), .Z(n46232) );
  NANDN U43478 ( .A(x[6428]), .B(y[6428]), .Z(n59076) );
  NAND U43479 ( .A(n59076), .B(n23195), .Z(n46230) );
  AND U43480 ( .A(n23197), .B(n23196), .Z(n46228) );
  NANDN U43481 ( .A(x[6426]), .B(y[6426]), .Z(n51068) );
  NAND U43482 ( .A(n59077), .B(n51068), .Z(n46226) );
  AND U43483 ( .A(n23199), .B(n23198), .Z(n46224) );
  NANDN U43484 ( .A(x[6424]), .B(y[6424]), .Z(n59072) );
  AND U43485 ( .A(n59072), .B(n51067), .Z(n46222) );
  NAND U43486 ( .A(n23201), .B(n23200), .Z(n46220) );
  AND U43487 ( .A(n23203), .B(n23202), .Z(n46216) );
  NANDN U43488 ( .A(x[6420]), .B(y[6420]), .Z(n59067) );
  IV U43489 ( .A(n23204), .Z(n59068) );
  AND U43490 ( .A(n59067), .B(n59068), .Z(n46214) );
  NANDN U43491 ( .A(x[6418]), .B(y[6418]), .Z(n51071) );
  AND U43492 ( .A(n23206), .B(n23205), .Z(n46206) );
  ANDN U43493 ( .B(y[6416]), .A(x[6416]), .Z(n59063) );
  NOR U43494 ( .A(n59063), .B(n51070), .Z(n46204) );
  AND U43495 ( .A(n23208), .B(n23207), .Z(n46195) );
  NANDN U43496 ( .A(x[6412]), .B(y[6412]), .Z(n59054) );
  AND U43497 ( .A(n59057), .B(n59054), .Z(n46193) );
  NAND U43498 ( .A(n23210), .B(n23209), .Z(n46191) );
  AND U43499 ( .A(n23212), .B(n23211), .Z(n46187) );
  ANDN U43500 ( .B(y[6408]), .A(x[6408]), .Z(n59051) );
  NOR U43501 ( .A(n59051), .B(n51072), .Z(n46185) );
  AND U43502 ( .A(n23214), .B(n23213), .Z(n46177) );
  ANDN U43503 ( .B(y[6404]), .A(x[6404]), .Z(n59045) );
  NOR U43504 ( .A(n59045), .B(n59048), .Z(n46175) );
  AND U43505 ( .A(n23216), .B(n23215), .Z(n46167) );
  NAND U43506 ( .A(n23218), .B(n23217), .Z(n46163) );
  AND U43507 ( .A(n23220), .B(n23219), .Z(n46158) );
  ANDN U43508 ( .B(y[6396]), .A(x[6396]), .Z(n51079) );
  NOR U43509 ( .A(n51079), .B(n59035), .Z(n46156) );
  AND U43510 ( .A(n23222), .B(n23221), .Z(n46148) );
  ANDN U43511 ( .B(y[6392]), .A(x[6392]), .Z(n59030) );
  NOR U43512 ( .A(n59030), .B(n51080), .Z(n46146) );
  AND U43513 ( .A(n23224), .B(n23223), .Z(n46137) );
  ANDN U43514 ( .B(y[6388]), .A(x[6388]), .Z(n59024) );
  NOR U43515 ( .A(n59024), .B(n59026), .Z(n46135) );
  AND U43516 ( .A(n23226), .B(n23225), .Z(n46127) );
  ANDN U43517 ( .B(y[6384]), .A(x[6384]), .Z(n59020) );
  NOR U43518 ( .A(n59020), .B(n51082), .Z(n46125) );
  AND U43519 ( .A(n23228), .B(n23227), .Z(n46117) );
  ANDN U43520 ( .B(y[6380]), .A(x[6380]), .Z(n59013) );
  NOR U43521 ( .A(n59014), .B(n59013), .Z(n46115) );
  AND U43522 ( .A(n23230), .B(n23229), .Z(n46107) );
  IV U43523 ( .A(n23231), .Z(n51085) );
  AND U43524 ( .A(n23233), .B(n23232), .Z(n46103) );
  IV U43525 ( .A(n23234), .Z(n59008) );
  NAND U43526 ( .A(n59008), .B(n23235), .Z(n46101) );
  AND U43527 ( .A(n23237), .B(n23236), .Z(n46099) );
  NANDN U43528 ( .A(x[6372]), .B(y[6372]), .Z(n51090) );
  AND U43529 ( .A(n51090), .B(n23238), .Z(n46097) );
  NAND U43530 ( .A(n23240), .B(n23239), .Z(n46095) );
  AND U43531 ( .A(n23242), .B(n23241), .Z(n46090) );
  IV U43532 ( .A(n23243), .Z(n59002) );
  AND U43533 ( .A(n23244), .B(n59002), .Z(n46088) );
  NANDN U43534 ( .A(x[6366]), .B(y[6366]), .Z(n51092) );
  AND U43535 ( .A(n23246), .B(n23245), .Z(n46079) );
  AND U43536 ( .A(n23248), .B(n23247), .Z(n46075) );
  NAND U43537 ( .A(n23249), .B(n58996), .Z(n46073) );
  AND U43538 ( .A(n23251), .B(n23250), .Z(n46071) );
  ANDN U43539 ( .B(y[6360]), .A(x[6360]), .Z(n51093) );
  NOR U43540 ( .A(n51093), .B(n23252), .Z(n46069) );
  AND U43541 ( .A(n23254), .B(n23253), .Z(n46061) );
  ANDN U43542 ( .B(y[6356]), .A(x[6356]), .Z(n58987) );
  NOR U43543 ( .A(n58987), .B(n58989), .Z(n46059) );
  AND U43544 ( .A(n23256), .B(n23255), .Z(n46050) );
  ANDN U43545 ( .B(y[6352]), .A(x[6352]), .Z(n51095) );
  NOR U43546 ( .A(n51095), .B(n58984), .Z(n46048) );
  AND U43547 ( .A(n23258), .B(n23257), .Z(n46040) );
  ANDN U43548 ( .B(y[6348]), .A(x[6348]), .Z(n58975) );
  NOR U43549 ( .A(n58975), .B(n58979), .Z(n46038) );
  AND U43550 ( .A(n23259), .B(n58977), .Z(n46032) );
  AND U43551 ( .A(n23261), .B(n23260), .Z(n46030) );
  AND U43552 ( .A(n23263), .B(n23262), .Z(n46024) );
  NAND U43553 ( .A(n23265), .B(n23264), .Z(n46022) );
  AND U43554 ( .A(n23267), .B(n23266), .Z(n46020) );
  AND U43555 ( .A(n23269), .B(n23268), .Z(n46015) );
  NAND U43556 ( .A(n23270), .B(n51098), .Z(n46013) );
  AND U43557 ( .A(n23272), .B(n23271), .Z(n46011) );
  AND U43558 ( .A(n23274), .B(n23273), .Z(n46009) );
  AND U43559 ( .A(n23276), .B(n23275), .Z(n46003) );
  NAND U43560 ( .A(n23278), .B(n23277), .Z(n46001) );
  AND U43561 ( .A(n23280), .B(n23279), .Z(n45995) );
  NAND U43562 ( .A(n23282), .B(n23281), .Z(n45993) );
  AND U43563 ( .A(n23284), .B(n23283), .Z(n45991) );
  AND U43564 ( .A(n23286), .B(n23285), .Z(n45989) );
  NAND U43565 ( .A(n23288), .B(n23287), .Z(n45987) );
  NANDN U43566 ( .A(x[6326]), .B(y[6326]), .Z(n58952) );
  AND U43567 ( .A(n58952), .B(n23289), .Z(n45985) );
  AND U43568 ( .A(n23291), .B(n23290), .Z(n45983) );
  ANDN U43569 ( .B(y[6324]), .A(x[6324]), .Z(n58948) );
  NOR U43570 ( .A(n58948), .B(n58951), .Z(n45981) );
  AND U43571 ( .A(n23293), .B(n23292), .Z(n45973) );
  NANDN U43572 ( .A(x[6320]), .B(y[6320]), .Z(n58945) );
  ANDN U43573 ( .B(n58945), .A(n51100), .Z(n45971) );
  AND U43574 ( .A(n23295), .B(n23294), .Z(n45963) );
  ANDN U43575 ( .B(y[6316]), .A(x[6316]), .Z(n58937) );
  NOR U43576 ( .A(n58937), .B(n58940), .Z(n45961) );
  AND U43577 ( .A(n23297), .B(n23296), .Z(n45953) );
  NANDN U43578 ( .A(x[6312]), .B(y[6312]), .Z(n58934) );
  ANDN U43579 ( .B(n58934), .A(n51102), .Z(n45951) );
  AND U43580 ( .A(n23299), .B(n23298), .Z(n45942) );
  ANDN U43581 ( .B(y[6308]), .A(x[6308]), .Z(n51105) );
  NOR U43582 ( .A(n51105), .B(n58930), .Z(n45940) );
  AND U43583 ( .A(n23301), .B(n23300), .Z(n45932) );
  NANDN U43584 ( .A(x[6304]), .B(y[6304]), .Z(n58925) );
  ANDN U43585 ( .B(n58925), .A(n51107), .Z(n45930) );
  AND U43586 ( .A(n23303), .B(n23302), .Z(n45922) );
  NANDN U43587 ( .A(x[6300]), .B(y[6300]), .Z(n58918) );
  AND U43588 ( .A(n58921), .B(n58918), .Z(n45920) );
  NAND U43589 ( .A(n23305), .B(n23304), .Z(n45918) );
  AND U43590 ( .A(n23307), .B(n23306), .Z(n45914) );
  NANDN U43591 ( .A(x[6296]), .B(y[6296]), .Z(n58915) );
  ANDN U43592 ( .B(n58915), .A(n51109), .Z(n45912) );
  AND U43593 ( .A(n23309), .B(n23308), .Z(n45904) );
  NANDN U43594 ( .A(x[6292]), .B(y[6292]), .Z(n58907) );
  AND U43595 ( .A(n58910), .B(n58907), .Z(n45902) );
  NAND U43596 ( .A(n23311), .B(n23310), .Z(n45900) );
  AND U43597 ( .A(n23313), .B(n23312), .Z(n45896) );
  NANDN U43598 ( .A(x[6288]), .B(y[6288]), .Z(n58904) );
  IV U43599 ( .A(n23314), .Z(n51111) );
  AND U43600 ( .A(n58904), .B(n51111), .Z(n45894) );
  AND U43601 ( .A(n23316), .B(n23315), .Z(n45892) );
  NANDN U43602 ( .A(x[6286]), .B(y[6286]), .Z(n58901) );
  NAND U43603 ( .A(n58901), .B(n58903), .Z(n45890) );
  AND U43604 ( .A(n23318), .B(n23317), .Z(n45888) );
  ANDN U43605 ( .B(y[6284]), .A(x[6284]), .Z(n58897) );
  NOR U43606 ( .A(n58897), .B(n58900), .Z(n45886) );
  AND U43607 ( .A(n23320), .B(n23319), .Z(n45878) );
  NANDN U43608 ( .A(x[6280]), .B(y[6280]), .Z(n58893) );
  IV U43609 ( .A(n23321), .Z(n51113) );
  AND U43610 ( .A(n58893), .B(n51113), .Z(n45876) );
  XNOR U43611 ( .A(y[6280]), .B(x[6280]), .Z(n45872) );
  AND U43612 ( .A(n23323), .B(n23322), .Z(n45868) );
  ANDN U43613 ( .B(y[6276]), .A(x[6276]), .Z(n58886) );
  NOR U43614 ( .A(n58889), .B(n58886), .Z(n45866) );
  AND U43615 ( .A(n23325), .B(n23324), .Z(n45858) );
  NANDN U43616 ( .A(x[6272]), .B(y[6272]), .Z(n58882) );
  ANDN U43617 ( .B(n58882), .A(n51115), .Z(n45856) );
  AND U43618 ( .A(n23327), .B(n23326), .Z(n45848) );
  ANDN U43619 ( .B(y[6268]), .A(x[6268]), .Z(n58876) );
  NOR U43620 ( .A(n58876), .B(n58878), .Z(n45846) );
  AND U43621 ( .A(n23328), .B(n58875), .Z(n45840) );
  AND U43622 ( .A(n23330), .B(n23329), .Z(n45838) );
  NANDN U43623 ( .A(x[6264]), .B(y[6264]), .Z(n51119) );
  NAND U43624 ( .A(n51119), .B(n23331), .Z(n45836) );
  AND U43625 ( .A(n23333), .B(n23332), .Z(n45834) );
  NANDN U43626 ( .A(x[6262]), .B(y[6262]), .Z(n58869) );
  NAND U43627 ( .A(n58869), .B(n58873), .Z(n45832) );
  AND U43628 ( .A(n23335), .B(n23334), .Z(n45830) );
  AND U43629 ( .A(n23337), .B(n23336), .Z(n45826) );
  ANDN U43630 ( .B(y[6258]), .A(x[6258]), .Z(n58864) );
  AND U43631 ( .A(n23339), .B(n23338), .Z(n45821) );
  NANDN U43632 ( .A(x[6256]), .B(y[6256]), .Z(n58861) );
  ANDN U43633 ( .B(n58861), .A(n58863), .Z(n45819) );
  AND U43634 ( .A(n23341), .B(n23340), .Z(n45811) );
  NANDN U43635 ( .A(x[6252]), .B(y[6252]), .Z(n51123) );
  AND U43636 ( .A(n51123), .B(n58858), .Z(n45809) );
  NAND U43637 ( .A(n23343), .B(n23342), .Z(n45807) );
  NANDN U43638 ( .A(x[6250]), .B(y[6250]), .Z(n58853) );
  IV U43639 ( .A(n23344), .Z(n51122) );
  AND U43640 ( .A(n58853), .B(n51122), .Z(n45805) );
  AND U43641 ( .A(n23346), .B(n23345), .Z(n45803) );
  NANDN U43642 ( .A(x[6248]), .B(y[6248]), .Z(n51124) );
  AND U43643 ( .A(n51124), .B(n58852), .Z(n45801) );
  NAND U43644 ( .A(n23348), .B(n23347), .Z(n45799) );
  AND U43645 ( .A(n23350), .B(n23349), .Z(n45794) );
  NAND U43646 ( .A(n23351), .B(n58848), .Z(n45792) );
  AND U43647 ( .A(n23353), .B(n23352), .Z(n45790) );
  NAND U43648 ( .A(n23355), .B(n23354), .Z(n45788) );
  AND U43649 ( .A(n23357), .B(n23356), .Z(n45786) );
  NANDN U43650 ( .A(x[6240]), .B(y[6240]), .Z(n58843) );
  NAND U43651 ( .A(n58843), .B(n23358), .Z(n45784) );
  AND U43652 ( .A(n23360), .B(n23359), .Z(n45782) );
  NANDN U43653 ( .A(x[6238]), .B(y[6238]), .Z(n51129) );
  NAND U43654 ( .A(n58842), .B(n51129), .Z(n45780) );
  AND U43655 ( .A(n23362), .B(n23361), .Z(n45778) );
  ANDN U43656 ( .B(y[6236]), .A(x[6236]), .Z(n58839) );
  NOR U43657 ( .A(n58839), .B(n51128), .Z(n45776) );
  AND U43658 ( .A(n23364), .B(n23363), .Z(n45768) );
  ANDN U43659 ( .B(y[6232]), .A(x[6232]), .Z(n58833) );
  NOR U43660 ( .A(n58833), .B(n58835), .Z(n45766) );
  AND U43661 ( .A(n23366), .B(n23365), .Z(n45758) );
  NANDN U43662 ( .A(x[6228]), .B(y[6228]), .Z(n58828) );
  IV U43663 ( .A(n23367), .Z(n51131) );
  ANDN U43664 ( .B(n58828), .A(n51131), .Z(n45756) );
  AND U43665 ( .A(n23369), .B(n23368), .Z(n45747) );
  NANDN U43666 ( .A(x[6224]), .B(y[6224]), .Z(n51134) );
  AND U43667 ( .A(n51134), .B(n23370), .Z(n45745) );
  NAND U43668 ( .A(n23372), .B(n23371), .Z(n45743) );
  NANDN U43669 ( .A(x[6222]), .B(y[6222]), .Z(n58822) );
  AND U43670 ( .A(n58822), .B(n51133), .Z(n45741) );
  AND U43671 ( .A(n23374), .B(n23373), .Z(n45739) );
  ANDN U43672 ( .B(y[6220]), .A(x[6220]), .Z(n58819) );
  NOR U43673 ( .A(n58819), .B(n58821), .Z(n45737) );
  AND U43674 ( .A(n23376), .B(n23375), .Z(n45728) );
  ANDN U43675 ( .B(y[6216]), .A(x[6216]), .Z(n51136) );
  NOR U43676 ( .A(n51136), .B(n58816), .Z(n45726) );
  AND U43677 ( .A(n23378), .B(n23377), .Z(n45718) );
  NANDN U43678 ( .A(x[6212]), .B(y[6212]), .Z(n58808) );
  ANDN U43679 ( .B(n58808), .A(n58810), .Z(n45716) );
  AND U43680 ( .A(n23380), .B(n23379), .Z(n45707) );
  NANDN U43681 ( .A(x[6208]), .B(y[6208]), .Z(n51140) );
  ANDN U43682 ( .B(n51140), .A(n51139), .Z(n45705) );
  AND U43683 ( .A(n23382), .B(n23381), .Z(n45697) );
  IV U43684 ( .A(n23383), .Z(n58801) );
  ANDN U43685 ( .B(y[6204]), .A(x[6204]), .Z(n58800) );
  NOR U43686 ( .A(n58801), .B(n58800), .Z(n45695) );
  AND U43687 ( .A(n23385), .B(n23384), .Z(n45686) );
  ANDN U43688 ( .B(y[6200]), .A(x[6200]), .Z(n51144) );
  NOR U43689 ( .A(n51144), .B(n58798), .Z(n45684) );
  AND U43690 ( .A(n23387), .B(n23386), .Z(n45676) );
  IV U43691 ( .A(n23388), .Z(n58793) );
  ANDN U43692 ( .B(y[6196]), .A(x[6196]), .Z(n58791) );
  NOR U43693 ( .A(n58793), .B(n58791), .Z(n45674) );
  AND U43694 ( .A(n23390), .B(n23389), .Z(n45665) );
  ANDN U43695 ( .B(y[6192]), .A(x[6192]), .Z(n51148) );
  NOR U43696 ( .A(n51148), .B(n58789), .Z(n45663) );
  AND U43697 ( .A(n23392), .B(n23391), .Z(n45655) );
  ANDN U43698 ( .B(y[6188]), .A(x[6188]), .Z(n58782) );
  NOR U43699 ( .A(n58782), .B(n58784), .Z(n45653) );
  AND U43700 ( .A(n23394), .B(n23393), .Z(n45644) );
  ANDN U43701 ( .B(y[6184]), .A(x[6184]), .Z(n51151) );
  NOR U43702 ( .A(n51151), .B(n58779), .Z(n45642) );
  AND U43703 ( .A(n23396), .B(n23395), .Z(n45634) );
  ANDN U43704 ( .B(y[6180]), .A(x[6180]), .Z(n58772) );
  NOR U43705 ( .A(n58772), .B(n58774), .Z(n45632) );
  AND U43706 ( .A(n23398), .B(n23397), .Z(n45623) );
  ANDN U43707 ( .B(y[6176]), .A(x[6176]), .Z(n51154) );
  ANDN U43708 ( .B(n58770), .A(n51154), .Z(n45621) );
  AND U43709 ( .A(n23400), .B(n23399), .Z(n45613) );
  NANDN U43710 ( .A(x[6172]), .B(y[6172]), .Z(n58759) );
  AND U43711 ( .A(n58759), .B(n58761), .Z(n45611) );
  NAND U43712 ( .A(n23402), .B(n23401), .Z(n45609) );
  IV U43713 ( .A(n23403), .Z(n58758) );
  AND U43714 ( .A(n23405), .B(n23404), .Z(n45605) );
  NAND U43715 ( .A(n23406), .B(n58757), .Z(n45603) );
  AND U43716 ( .A(n23408), .B(n23407), .Z(n45601) );
  NANDN U43717 ( .A(x[6166]), .B(y[6166]), .Z(n58754) );
  NAND U43718 ( .A(n58754), .B(n23409), .Z(n45599) );
  AND U43719 ( .A(n23411), .B(n23410), .Z(n45597) );
  NAND U43720 ( .A(n23412), .B(n58753), .Z(n45595) );
  AND U43721 ( .A(n23414), .B(n23413), .Z(n45593) );
  NANDN U43722 ( .A(x[6162]), .B(y[6162]), .Z(n51160) );
  AND U43723 ( .A(n23416), .B(n23415), .Z(n45588) );
  ANDN U43724 ( .B(y[6160]), .A(x[6160]), .Z(n58747) );
  NOR U43725 ( .A(n58747), .B(n51159), .Z(n45586) );
  AND U43726 ( .A(n23418), .B(n23417), .Z(n45578) );
  ANDN U43727 ( .B(y[6156]), .A(x[6156]), .Z(n58741) );
  NOR U43728 ( .A(n58743), .B(n58741), .Z(n45576) );
  AND U43729 ( .A(n23420), .B(n23419), .Z(n45568) );
  ANDN U43730 ( .B(y[6152]), .A(x[6152]), .Z(n58737) );
  NOR U43731 ( .A(n58737), .B(n51162), .Z(n45566) );
  AND U43732 ( .A(n23422), .B(n23421), .Z(n45558) );
  AND U43733 ( .A(n23424), .B(n23423), .Z(n45554) );
  AND U43734 ( .A(n23425), .B(n58732), .Z(n45552) );
  AND U43735 ( .A(n23427), .B(n23426), .Z(n45550) );
  NANDN U43736 ( .A(x[6144]), .B(y[6144]), .Z(n51166) );
  NAND U43737 ( .A(n51166), .B(n23428), .Z(n45548) );
  AND U43738 ( .A(n23430), .B(n23429), .Z(n45546) );
  AND U43739 ( .A(n23432), .B(n23431), .Z(n45542) );
  AND U43740 ( .A(n23434), .B(n23433), .Z(n45537) );
  NANDN U43741 ( .A(x[6138]), .B(y[6138]), .Z(n58719) );
  NAND U43742 ( .A(n58719), .B(n23435), .Z(n45535) );
  AND U43743 ( .A(n23437), .B(n23436), .Z(n45533) );
  NAND U43744 ( .A(n23439), .B(n23438), .Z(n45528) );
  AND U43745 ( .A(n23441), .B(n23440), .Z(n45523) );
  NAND U43746 ( .A(n23443), .B(n23442), .Z(n45519) );
  AND U43747 ( .A(n23445), .B(n23444), .Z(n45515) );
  NAND U43748 ( .A(n23447), .B(n23446), .Z(n45511) );
  AND U43749 ( .A(n23449), .B(n23448), .Z(n45506) );
  ANDN U43750 ( .B(y[6122]), .A(x[6122]), .Z(n58699) );
  AND U43751 ( .A(n23451), .B(n23450), .Z(n45494) );
  NAND U43752 ( .A(n23453), .B(n23452), .Z(n45490) );
  AND U43753 ( .A(n23455), .B(n23454), .Z(n45486) );
  NAND U43754 ( .A(n23457), .B(n23456), .Z(n45482) );
  AND U43755 ( .A(n23459), .B(n23458), .Z(n45478) );
  NAND U43756 ( .A(n23461), .B(n23460), .Z(n45474) );
  AND U43757 ( .A(n23463), .B(n23462), .Z(n45470) );
  NAND U43758 ( .A(n23465), .B(n23464), .Z(n45465) );
  AND U43759 ( .A(n23467), .B(n23466), .Z(n45461) );
  NAND U43760 ( .A(n23469), .B(n23468), .Z(n45457) );
  AND U43761 ( .A(n23471), .B(n23470), .Z(n45453) );
  NAND U43762 ( .A(n23473), .B(n23472), .Z(n45449) );
  AND U43763 ( .A(n23475), .B(n23474), .Z(n45445) );
  NANDN U43764 ( .A(x[6094]), .B(y[6094]), .Z(n51182) );
  AND U43765 ( .A(n51182), .B(n51179), .Z(n45437) );
  NAND U43766 ( .A(n23477), .B(n23476), .Z(n45435) );
  NAND U43767 ( .A(n23479), .B(n23478), .Z(n45431) );
  NANDN U43768 ( .A(x[6090]), .B(y[6090]), .Z(n58659) );
  AND U43769 ( .A(n23481), .B(n23480), .Z(n45427) );
  NAND U43770 ( .A(n23483), .B(n23482), .Z(n45423) );
  NANDN U43771 ( .A(x[6086]), .B(y[6086]), .Z(n51184) );
  AND U43772 ( .A(n23485), .B(n23484), .Z(n45419) );
  NAND U43773 ( .A(n23487), .B(n23486), .Z(n45415) );
  NANDN U43774 ( .A(x[6082]), .B(y[6082]), .Z(n58649) );
  AND U43775 ( .A(n23489), .B(n23488), .Z(n45411) );
  NAND U43776 ( .A(n23491), .B(n23490), .Z(n45407) );
  AND U43777 ( .A(n23493), .B(n23492), .Z(n45403) );
  NAND U43778 ( .A(n23495), .B(n23494), .Z(n45399) );
  NANDN U43779 ( .A(x[6074]), .B(y[6074]), .Z(n58636) );
  IV U43780 ( .A(n23496), .Z(n58638) );
  AND U43781 ( .A(n58636), .B(n58638), .Z(n45397) );
  NAND U43782 ( .A(n23498), .B(n23497), .Z(n45395) );
  NAND U43783 ( .A(n23500), .B(n23499), .Z(n45391) );
  AND U43784 ( .A(n23502), .B(n23501), .Z(n45387) );
  IV U43785 ( .A(n23503), .Z(n51187) );
  AND U43786 ( .A(n23504), .B(n51187), .Z(n45385) );
  NAND U43787 ( .A(n23506), .B(n23505), .Z(n45383) );
  AND U43788 ( .A(n23508), .B(n23507), .Z(n45381) );
  NAND U43789 ( .A(n23510), .B(n23509), .Z(n45379) );
  NAND U43790 ( .A(n23512), .B(n23511), .Z(n45374) );
  AND U43791 ( .A(n23513), .B(n51189), .Z(n45372) );
  NAND U43792 ( .A(n23515), .B(n23514), .Z(n45370) );
  AND U43793 ( .A(n23517), .B(n23516), .Z(n45368) );
  NAND U43794 ( .A(n23519), .B(n23518), .Z(n45366) );
  NANDN U43795 ( .A(x[6058]), .B(y[6058]), .Z(n51192) );
  AND U43796 ( .A(n23521), .B(n23520), .Z(n45361) );
  NAND U43797 ( .A(n23523), .B(n23522), .Z(n45357) );
  AND U43798 ( .A(n23524), .B(n58617), .Z(n45355) );
  NAND U43799 ( .A(n23526), .B(n23525), .Z(n45353) );
  AND U43800 ( .A(n23528), .B(n23527), .Z(n45351) );
  NAND U43801 ( .A(n23530), .B(n23529), .Z(n45349) );
  AND U43802 ( .A(n23532), .B(n23531), .Z(n45347) );
  NAND U43803 ( .A(n23534), .B(n23533), .Z(n45345) );
  NAND U43804 ( .A(n23536), .B(n23535), .Z(n45340) );
  NANDN U43805 ( .A(x[6046]), .B(y[6046]), .Z(n51194) );
  AND U43806 ( .A(n23538), .B(n23537), .Z(n45336) );
  NAND U43807 ( .A(n23540), .B(n23539), .Z(n45332) );
  NANDN U43808 ( .A(x[6042]), .B(y[6042]), .Z(n58601) );
  AND U43809 ( .A(n23542), .B(n23541), .Z(n45328) );
  NANDN U43810 ( .A(x[6038]), .B(y[6038]), .Z(n23543) );
  NAND U43811 ( .A(n23543), .B(n58598), .Z(n45320) );
  NAND U43812 ( .A(n23545), .B(n23544), .Z(n45311) );
  NANDN U43813 ( .A(x[6034]), .B(y[6034]), .Z(n58589) );
  IV U43814 ( .A(n23546), .Z(n58592) );
  AND U43815 ( .A(n23548), .B(n23547), .Z(n45307) );
  AND U43816 ( .A(n23550), .B(n23549), .Z(n45297) );
  NAND U43817 ( .A(n23552), .B(n23551), .Z(n45293) );
  NANDN U43818 ( .A(x[6026]), .B(y[6026]), .Z(n58578) );
  AND U43819 ( .A(n23554), .B(n23553), .Z(n45289) );
  NAND U43820 ( .A(n23556), .B(n23555), .Z(n45285) );
  NANDN U43821 ( .A(x[6022]), .B(y[6022]), .Z(n23557) );
  AND U43822 ( .A(n23557), .B(n51198), .Z(n45283) );
  NAND U43823 ( .A(n23559), .B(n23558), .Z(n45281) );
  AND U43824 ( .A(n23561), .B(n23560), .Z(n45270) );
  NAND U43825 ( .A(n23563), .B(n23562), .Z(n45266) );
  AND U43826 ( .A(n23565), .B(n23564), .Z(n45261) );
  NAND U43827 ( .A(n23567), .B(n23566), .Z(n45256) );
  AND U43828 ( .A(n23569), .B(n23568), .Z(n45252) );
  NAND U43829 ( .A(n23571), .B(n23570), .Z(n45248) );
  AND U43830 ( .A(n23573), .B(n23572), .Z(n45243) );
  NAND U43831 ( .A(n23575), .B(n23574), .Z(n45238) );
  AND U43832 ( .A(n23577), .B(n23576), .Z(n45234) );
  NAND U43833 ( .A(n23579), .B(n23578), .Z(n45230) );
  AND U43834 ( .A(n23581), .B(n23580), .Z(n45225) );
  NAND U43835 ( .A(n23583), .B(n23582), .Z(n45220) );
  AND U43836 ( .A(n23585), .B(n23584), .Z(n45216) );
  NAND U43837 ( .A(n23587), .B(n23586), .Z(n45212) );
  NANDN U43838 ( .A(x[5990]), .B(y[5990]), .Z(n58533) );
  IV U43839 ( .A(n23588), .Z(n58535) );
  AND U43840 ( .A(n23590), .B(n23589), .Z(n45208) );
  NAND U43841 ( .A(n23592), .B(n23591), .Z(n45203) );
  AND U43842 ( .A(n23594), .B(n23593), .Z(n45199) );
  AND U43843 ( .A(n23596), .B(n23595), .Z(n45195) );
  AND U43844 ( .A(n23598), .B(n23597), .Z(n45191) );
  ANDN U43845 ( .B(y[5980]), .A(x[5980]), .Z(n58518) );
  NAND U43846 ( .A(n23600), .B(n23599), .Z(n45186) );
  NANDN U43847 ( .A(x[5978]), .B(y[5978]), .Z(n51216) );
  AND U43848 ( .A(n23602), .B(n23601), .Z(n45182) );
  NAND U43849 ( .A(n23604), .B(n23603), .Z(n45178) );
  NANDN U43850 ( .A(x[5974]), .B(y[5974]), .Z(n58512) );
  IV U43851 ( .A(n23605), .Z(n58514) );
  AND U43852 ( .A(n23607), .B(n23606), .Z(n45174) );
  NAND U43853 ( .A(n23609), .B(n23608), .Z(n45170) );
  NANDN U43854 ( .A(x[5970]), .B(y[5970]), .Z(n51218) );
  AND U43855 ( .A(n23611), .B(n23610), .Z(n45166) );
  AND U43856 ( .A(n23612), .B(n51217), .Z(n45164) );
  AND U43857 ( .A(n23614), .B(n23613), .Z(n45158) );
  NAND U43858 ( .A(n23616), .B(n23615), .Z(n45156) );
  NAND U43859 ( .A(n23618), .B(n23617), .Z(n45151) );
  NANDN U43860 ( .A(x[5962]), .B(y[5962]), .Z(n58497) );
  AND U43861 ( .A(n23620), .B(n23619), .Z(n45147) );
  IV U43862 ( .A(n23621), .Z(n58496) );
  AND U43863 ( .A(n23622), .B(n58496), .Z(n45145) );
  NAND U43864 ( .A(n23624), .B(n23623), .Z(n45143) );
  NANDN U43865 ( .A(x[5958]), .B(y[5958]), .Z(n51223) );
  AND U43866 ( .A(n23626), .B(n23625), .Z(n45138) );
  AND U43867 ( .A(n23627), .B(n58490), .Z(n45130) );
  NAND U43868 ( .A(n23629), .B(n23628), .Z(n45128) );
  AND U43869 ( .A(n23631), .B(n23630), .Z(n45117) );
  NAND U43870 ( .A(n23633), .B(n23632), .Z(n45112) );
  AND U43871 ( .A(n23635), .B(n23634), .Z(n45107) );
  NAND U43872 ( .A(n23637), .B(n23636), .Z(n45103) );
  AND U43873 ( .A(n23639), .B(n23638), .Z(n45099) );
  NAND U43874 ( .A(n23641), .B(n23640), .Z(n45094) );
  AND U43875 ( .A(n23643), .B(n23642), .Z(n45090) );
  NAND U43876 ( .A(n23645), .B(n23644), .Z(n45085) );
  AND U43877 ( .A(n23647), .B(n23646), .Z(n45080) );
  NANDN U43878 ( .A(x[5930]), .B(y[5930]), .Z(n51232) );
  AND U43879 ( .A(n51232), .B(n58459), .Z(n45072) );
  NAND U43880 ( .A(n23649), .B(n23648), .Z(n45070) );
  NAND U43881 ( .A(n23651), .B(n23650), .Z(n45065) );
  NANDN U43882 ( .A(x[5926]), .B(y[5926]), .Z(n58453) );
  AND U43883 ( .A(n23653), .B(n23652), .Z(n45061) );
  AND U43884 ( .A(n23655), .B(n23654), .Z(n45057) );
  NAND U43885 ( .A(n23656), .B(n58450), .Z(n45055) );
  AND U43886 ( .A(n23658), .B(n23657), .Z(n45053) );
  NAND U43887 ( .A(n23660), .B(n23659), .Z(n45047) );
  AND U43888 ( .A(n23662), .B(n23661), .Z(n45042) );
  NAND U43889 ( .A(n23664), .B(n23663), .Z(n45038) );
  AND U43890 ( .A(n23666), .B(n23665), .Z(n45034) );
  NAND U43891 ( .A(n23668), .B(n23667), .Z(n45029) );
  AND U43892 ( .A(n23670), .B(n23669), .Z(n45025) );
  NAND U43893 ( .A(n23672), .B(n23671), .Z(n45021) );
  AND U43894 ( .A(n23674), .B(n23673), .Z(n45017) );
  NAND U43895 ( .A(n23676), .B(n23675), .Z(n45012) );
  AND U43896 ( .A(n23678), .B(n23677), .Z(n45008) );
  NAND U43897 ( .A(n23680), .B(n23679), .Z(n45004) );
  AND U43898 ( .A(n23682), .B(n23681), .Z(n45000) );
  NAND U43899 ( .A(n23684), .B(n23683), .Z(n44995) );
  AND U43900 ( .A(n23686), .B(n23685), .Z(n44991) );
  NAND U43901 ( .A(n23688), .B(n23687), .Z(n44987) );
  AND U43902 ( .A(n23690), .B(n23689), .Z(n44983) );
  NAND U43903 ( .A(n23692), .B(n23691), .Z(n44978) );
  AND U43904 ( .A(n23694), .B(n23693), .Z(n44974) );
  NAND U43905 ( .A(n23696), .B(n23695), .Z(n44970) );
  AND U43906 ( .A(n23698), .B(n23697), .Z(n44966) );
  NAND U43907 ( .A(n23700), .B(n23699), .Z(n44961) );
  ANDN U43908 ( .B(y[5878]), .A(x[5878]), .Z(n58387) );
  NOR U43909 ( .A(n58387), .B(n58390), .Z(n44959) );
  NAND U43910 ( .A(n23702), .B(n23701), .Z(n44951) );
  NANDN U43911 ( .A(x[5874]), .B(y[5874]), .Z(n58383) );
  AND U43912 ( .A(n23704), .B(n23703), .Z(n44947) );
  IV U43913 ( .A(n23705), .Z(n58382) );
  AND U43914 ( .A(n23706), .B(n58382), .Z(n44945) );
  NAND U43915 ( .A(n23708), .B(n23707), .Z(n44943) );
  NANDN U43916 ( .A(x[5870]), .B(y[5870]), .Z(n51250) );
  AND U43917 ( .A(n23710), .B(n23709), .Z(n44938) );
  NAND U43918 ( .A(n23712), .B(n23711), .Z(n44933) );
  IV U43919 ( .A(n23713), .Z(n58377) );
  AND U43920 ( .A(n23714), .B(n58377), .Z(n44931) );
  NAND U43921 ( .A(n23716), .B(n23715), .Z(n44929) );
  NAND U43922 ( .A(n23718), .B(n23717), .Z(n44924) );
  NANDN U43923 ( .A(x[5862]), .B(y[5862]), .Z(n58372) );
  AND U43924 ( .A(n23720), .B(n23719), .Z(n44920) );
  AND U43925 ( .A(n23721), .B(n58371), .Z(n44918) );
  AND U43926 ( .A(n23723), .B(n23722), .Z(n44916) );
  NAND U43927 ( .A(n23725), .B(n23724), .Z(n44914) );
  AND U43928 ( .A(n23727), .B(n23726), .Z(n44912) );
  NAND U43929 ( .A(n23729), .B(n23728), .Z(n44907) );
  AND U43930 ( .A(n23731), .B(n23730), .Z(n44903) );
  NANDN U43931 ( .A(x[5850]), .B(y[5850]), .Z(n51255) );
  AND U43932 ( .A(n51255), .B(n58359), .Z(n44894) );
  NAND U43933 ( .A(n23733), .B(n23732), .Z(n44892) );
  NAND U43934 ( .A(n23735), .B(n23734), .Z(n44888) );
  NANDN U43935 ( .A(x[5846]), .B(y[5846]), .Z(n58352) );
  AND U43936 ( .A(n23737), .B(n23736), .Z(n44884) );
  NAND U43937 ( .A(n23739), .B(n23738), .Z(n44879) );
  NANDN U43938 ( .A(x[5842]), .B(y[5842]), .Z(n51258) );
  AND U43939 ( .A(n23741), .B(n23740), .Z(n44875) );
  NAND U43940 ( .A(n23743), .B(n23742), .Z(n44871) );
  NANDN U43941 ( .A(x[5838]), .B(y[5838]), .Z(n58342) );
  AND U43942 ( .A(n23745), .B(n23744), .Z(n44867) );
  XNOR U43943 ( .A(x[5836]), .B(y[5836]), .Z(n23747) );
  NAND U43944 ( .A(n23747), .B(n23746), .Z(n44862) );
  NANDN U43945 ( .A(x[5834]), .B(y[5834]), .Z(n23748) );
  AND U43946 ( .A(n23748), .B(n58340), .Z(n44860) );
  NAND U43947 ( .A(n23750), .B(n23749), .Z(n44858) );
  NAND U43948 ( .A(n23752), .B(n23751), .Z(n44853) );
  NANDN U43949 ( .A(x[5830]), .B(y[5830]), .Z(n58331) );
  IV U43950 ( .A(n23753), .Z(n58333) );
  AND U43951 ( .A(n23755), .B(n23754), .Z(n44849) );
  ANDN U43952 ( .B(y[5826]), .A(x[5826]), .Z(n51261) );
  AND U43953 ( .A(n23757), .B(n23756), .Z(n44838) );
  AND U43954 ( .A(n23758), .B(n51262), .Z(n44836) );
  AND U43955 ( .A(n23760), .B(n23759), .Z(n44834) );
  NANDN U43956 ( .A(x[5822]), .B(y[5822]), .Z(n58322) );
  AND U43957 ( .A(n58322), .B(n23761), .Z(n44832) );
  NAND U43958 ( .A(n23763), .B(n23762), .Z(n44830) );
  NAND U43959 ( .A(n23765), .B(n23764), .Z(n44825) );
  NANDN U43960 ( .A(x[5818]), .B(y[5818]), .Z(n23766) );
  AND U43961 ( .A(n23766), .B(n51265), .Z(n44823) );
  NAND U43962 ( .A(n23768), .B(n23767), .Z(n44821) );
  AND U43963 ( .A(n23770), .B(n23769), .Z(n44816) );
  AND U43964 ( .A(n23772), .B(n23771), .Z(n44811) );
  NAND U43965 ( .A(n23774), .B(n23773), .Z(n44806) );
  AND U43966 ( .A(n23776), .B(n23775), .Z(n44802) );
  NAND U43967 ( .A(n23778), .B(n23777), .Z(n44798) );
  AND U43968 ( .A(n23780), .B(n23779), .Z(n44794) );
  NAND U43969 ( .A(n23782), .B(n23781), .Z(n44789) );
  AND U43970 ( .A(n23784), .B(n23783), .Z(n44785) );
  NANDN U43971 ( .A(x[5798]), .B(y[5798]), .Z(n58273) );
  AND U43972 ( .A(n58273), .B(n58276), .Z(n44777) );
  NAND U43973 ( .A(n23786), .B(n23785), .Z(n44775) );
  NAND U43974 ( .A(n23788), .B(n23787), .Z(n44770) );
  NANDN U43975 ( .A(x[5794]), .B(y[5794]), .Z(n58267) );
  AND U43976 ( .A(n23790), .B(n23789), .Z(n44766) );
  NAND U43977 ( .A(n23792), .B(n23791), .Z(n44749) );
  NANDN U43978 ( .A(x[5786]), .B(y[5786]), .Z(n58258) );
  AND U43979 ( .A(n23794), .B(n23793), .Z(n44745) );
  NAND U43980 ( .A(n23796), .B(n23795), .Z(n44741) );
  AND U43981 ( .A(n23798), .B(n23797), .Z(n44737) );
  NAND U43982 ( .A(n23800), .B(n23799), .Z(n44733) );
  AND U43983 ( .A(n23801), .B(n58250), .Z(n44731) );
  NAND U43984 ( .A(n23803), .B(n23802), .Z(n44729) );
  AND U43985 ( .A(n23805), .B(n23804), .Z(n44727) );
  NAND U43986 ( .A(n23807), .B(n23806), .Z(n44725) );
  NANDN U43987 ( .A(x[5774]), .B(y[5774]), .Z(n58243) );
  AND U43988 ( .A(n58243), .B(n23808), .Z(n44723) );
  NAND U43989 ( .A(n23810), .B(n23809), .Z(n44721) );
  AND U43990 ( .A(n23811), .B(n58242), .Z(n44719) );
  NAND U43991 ( .A(n23813), .B(n23812), .Z(n44713) );
  AND U43992 ( .A(n23815), .B(n23814), .Z(n44707) );
  AND U43993 ( .A(n23817), .B(n23816), .Z(n44701) );
  NAND U43994 ( .A(n23819), .B(n23818), .Z(n44699) );
  AND U43995 ( .A(n23821), .B(n23820), .Z(n44697) );
  AND U43996 ( .A(n23823), .B(n23822), .Z(n44695) );
  AND U43997 ( .A(n23825), .B(n23824), .Z(n44693) );
  NAND U43998 ( .A(n23827), .B(n23826), .Z(n44691) );
  NAND U43999 ( .A(n23829), .B(n23828), .Z(n44686) );
  AND U44000 ( .A(n23831), .B(n23830), .Z(n44681) );
  NAND U44001 ( .A(n23833), .B(n23832), .Z(n44676) );
  AND U44002 ( .A(n23835), .B(n23834), .Z(n44672) );
  NAND U44003 ( .A(n23837), .B(n23836), .Z(n44668) );
  AND U44004 ( .A(n23839), .B(n23838), .Z(n44664) );
  NAND U44005 ( .A(n23841), .B(n23840), .Z(n44658) );
  AND U44006 ( .A(n23843), .B(n23842), .Z(n44653) );
  NAND U44007 ( .A(n23845), .B(n23844), .Z(n44649) );
  AND U44008 ( .A(n23847), .B(n23846), .Z(n44645) );
  NAND U44009 ( .A(n23849), .B(n23848), .Z(n44641) );
  AND U44010 ( .A(n23851), .B(n23850), .Z(n44637) );
  NANDN U44011 ( .A(x[5734]), .B(y[5734]), .Z(n58200) );
  ANDN U44012 ( .B(n58200), .A(n58202), .Z(n44629) );
  AND U44013 ( .A(n23853), .B(n23852), .Z(n44612) );
  NAND U44014 ( .A(n23855), .B(n23854), .Z(n44608) );
  AND U44015 ( .A(n23857), .B(n23856), .Z(n44603) );
  NAND U44016 ( .A(n23859), .B(n23858), .Z(n44599) );
  AND U44017 ( .A(n23861), .B(n23860), .Z(n44595) );
  NAND U44018 ( .A(n23863), .B(n23862), .Z(n44591) );
  AND U44019 ( .A(n23865), .B(n23864), .Z(n44587) );
  NAND U44020 ( .A(n23867), .B(n23866), .Z(n44582) );
  AND U44021 ( .A(n23869), .B(n23868), .Z(n44577) );
  NANDN U44022 ( .A(x[5710]), .B(y[5710]), .Z(n51303) );
  AND U44023 ( .A(n51303), .B(n23870), .Z(n44568) );
  NAND U44024 ( .A(n23872), .B(n23871), .Z(n44566) );
  AND U44025 ( .A(n23873), .B(n58170), .Z(n44558) );
  NAND U44026 ( .A(n23875), .B(n23874), .Z(n44556) );
  AND U44027 ( .A(n23877), .B(n23876), .Z(n44554) );
  NAND U44028 ( .A(n23879), .B(n23878), .Z(n44552) );
  NANDN U44029 ( .A(x[5702]), .B(y[5702]), .Z(n58164) );
  AND U44030 ( .A(n23881), .B(n23880), .Z(n44547) );
  NAND U44031 ( .A(n23883), .B(n23882), .Z(n44542) );
  NANDN U44032 ( .A(x[5698]), .B(y[5698]), .Z(n51305) );
  AND U44033 ( .A(n51305), .B(n23884), .Z(n44540) );
  NAND U44034 ( .A(n23886), .B(n23885), .Z(n44538) );
  NAND U44035 ( .A(n23888), .B(n23887), .Z(n44534) );
  NANDN U44036 ( .A(x[5694]), .B(y[5694]), .Z(n51308) );
  IV U44037 ( .A(n23889), .Z(n58156) );
  AND U44038 ( .A(n23891), .B(n23890), .Z(n44530) );
  AND U44039 ( .A(n23892), .B(n51307), .Z(n44528) );
  NAND U44040 ( .A(n23894), .B(n23893), .Z(n44526) );
  NANDN U44041 ( .A(x[5690]), .B(y[5690]), .Z(n58152) );
  AND U44042 ( .A(n23896), .B(n23895), .Z(n44521) );
  NAND U44043 ( .A(n23898), .B(n23897), .Z(n44517) );
  NANDN U44044 ( .A(x[5686]), .B(y[5686]), .Z(n58145) );
  IV U44045 ( .A(n23899), .Z(n58147) );
  AND U44046 ( .A(n23901), .B(n23900), .Z(n44513) );
  IV U44047 ( .A(n23902), .Z(n51310) );
  ANDN U44048 ( .B(y[5682]), .A(x[5682]), .Z(n58142) );
  AND U44049 ( .A(n23904), .B(n23903), .Z(n44503) );
  NAND U44050 ( .A(n23906), .B(n23905), .Z(n44498) );
  NANDN U44051 ( .A(x[5678]), .B(y[5678]), .Z(n58134) );
  AND U44052 ( .A(n23908), .B(n23907), .Z(n44494) );
  NAND U44053 ( .A(n23910), .B(n23909), .Z(n44490) );
  AND U44054 ( .A(n23912), .B(n23911), .Z(n44486) );
  AND U44055 ( .A(n23913), .B(n58127), .Z(n44484) );
  NAND U44056 ( .A(n23915), .B(n23914), .Z(n44482) );
  NANDN U44057 ( .A(x[5670]), .B(y[5670]), .Z(n51316) );
  AND U44058 ( .A(n23917), .B(n23916), .Z(n44477) );
  NAND U44059 ( .A(n23919), .B(n23918), .Z(n44472) );
  AND U44060 ( .A(n23920), .B(n58123), .Z(n44470) );
  NAND U44061 ( .A(n23922), .B(n23921), .Z(n44468) );
  NAND U44062 ( .A(n23924), .B(n23923), .Z(n44463) );
  NANDN U44063 ( .A(x[5662]), .B(y[5662]), .Z(n58117) );
  AND U44064 ( .A(n23926), .B(n23925), .Z(n44459) );
  NAND U44065 ( .A(n23928), .B(n23927), .Z(n44455) );
  NANDN U44066 ( .A(x[5658]), .B(y[5658]), .Z(n58111) );
  IV U44067 ( .A(n23929), .Z(n58113) );
  AND U44068 ( .A(n23931), .B(n23930), .Z(n44451) );
  NANDN U44069 ( .A(x[5654]), .B(y[5654]), .Z(n58106) );
  AND U44070 ( .A(n23933), .B(n23932), .Z(n44441) );
  NAND U44071 ( .A(n23935), .B(n23934), .Z(n44436) );
  NANDN U44072 ( .A(x[5650]), .B(y[5650]), .Z(n51323) );
  AND U44073 ( .A(n51323), .B(n23936), .Z(n44434) );
  NAND U44074 ( .A(n23938), .B(n23937), .Z(n44432) );
  NAND U44075 ( .A(n23940), .B(n23939), .Z(n44428) );
  NANDN U44076 ( .A(x[5646]), .B(y[5646]), .Z(n58097) );
  IV U44077 ( .A(n23941), .Z(n58099) );
  AND U44078 ( .A(n23943), .B(n23942), .Z(n44424) );
  NAND U44079 ( .A(n23945), .B(n23944), .Z(n44420) );
  NANDN U44080 ( .A(x[5642]), .B(y[5642]), .Z(n51325) );
  AND U44081 ( .A(n23947), .B(n23946), .Z(n44416) );
  NAND U44082 ( .A(n23949), .B(n23948), .Z(n44411) );
  NANDN U44083 ( .A(x[5638]), .B(y[5638]), .Z(n58085) );
  AND U44084 ( .A(n23951), .B(n23950), .Z(n44407) );
  NAND U44085 ( .A(n23953), .B(n23952), .Z(n44403) );
  NANDN U44086 ( .A(x[5634]), .B(y[5634]), .Z(n51327) );
  AND U44087 ( .A(n23955), .B(n23954), .Z(n44399) );
  ANDN U44088 ( .B(y[5630]), .A(x[5630]), .Z(n58074) );
  AND U44089 ( .A(n23957), .B(n23956), .Z(n44388) );
  NAND U44090 ( .A(n23959), .B(n23958), .Z(n44384) );
  AND U44091 ( .A(n23961), .B(n23960), .Z(n44380) );
  NAND U44092 ( .A(n23963), .B(n23962), .Z(n44376) );
  AND U44093 ( .A(n23964), .B(n58065), .Z(n44374) );
  NAND U44094 ( .A(n23966), .B(n23965), .Z(n44372) );
  NAND U44095 ( .A(n23968), .B(n23967), .Z(n44367) );
  NANDN U44096 ( .A(x[5618]), .B(y[5618]), .Z(n23969) );
  AND U44097 ( .A(n23969), .B(n51330), .Z(n44365) );
  NAND U44098 ( .A(n23971), .B(n23970), .Z(n44363) );
  NAND U44099 ( .A(n23973), .B(n23972), .Z(n44357) );
  AND U44100 ( .A(n23975), .B(n23974), .Z(n44352) );
  IV U44101 ( .A(n23976), .Z(n58054) );
  AND U44102 ( .A(n23977), .B(n58054), .Z(n44343) );
  NAND U44103 ( .A(n23979), .B(n23978), .Z(n44341) );
  AND U44104 ( .A(n23981), .B(n23980), .Z(n44336) );
  NAND U44105 ( .A(n23982), .B(n51336), .Z(n44334) );
  AND U44106 ( .A(n23984), .B(n23983), .Z(n44332) );
  NAND U44107 ( .A(n23986), .B(n23985), .Z(n44327) );
  NANDN U44108 ( .A(x[5602]), .B(y[5602]), .Z(n51339) );
  AND U44109 ( .A(n51339), .B(n58045), .Z(n44325) );
  NAND U44110 ( .A(n23988), .B(n23987), .Z(n44323) );
  AND U44111 ( .A(n23989), .B(n51338), .Z(n44321) );
  NAND U44112 ( .A(n23991), .B(n23990), .Z(n44319) );
  NANDN U44113 ( .A(x[5598]), .B(y[5598]), .Z(n58038) );
  AND U44114 ( .A(n23992), .B(n58038), .Z(n44317) );
  NAND U44115 ( .A(n23994), .B(n23993), .Z(n44315) );
  NAND U44116 ( .A(n23996), .B(n23995), .Z(n44310) );
  NANDN U44117 ( .A(x[5594]), .B(y[5594]), .Z(n23998) );
  AND U44118 ( .A(n23998), .B(n23997), .Z(n44308) );
  NAND U44119 ( .A(n24000), .B(n23999), .Z(n44306) );
  AND U44120 ( .A(n24002), .B(n24001), .Z(n44304) );
  NAND U44121 ( .A(n24004), .B(n24003), .Z(n44302) );
  NANDN U44122 ( .A(x[5590]), .B(y[5590]), .Z(n51341) );
  AND U44123 ( .A(n24006), .B(n24005), .Z(n44297) );
  AND U44124 ( .A(n24007), .B(n51340), .Z(n44295) );
  NAND U44125 ( .A(n24009), .B(n24008), .Z(n44293) );
  NANDN U44126 ( .A(x[5586]), .B(y[5586]), .Z(n58025) );
  AND U44127 ( .A(n24010), .B(n58025), .Z(n44291) );
  NAND U44128 ( .A(n24012), .B(n24011), .Z(n44289) );
  NAND U44129 ( .A(n24014), .B(n24013), .Z(n44285) );
  NANDN U44130 ( .A(x[5582]), .B(y[5582]), .Z(n44283) );
  AND U44131 ( .A(n24016), .B(n24015), .Z(n44280) );
  AND U44132 ( .A(n24017), .B(n58020), .Z(n44271) );
  AND U44133 ( .A(n58016), .B(n24018), .Z(n44261) );
  AND U44134 ( .A(n24020), .B(n24019), .Z(n44255) );
  AND U44135 ( .A(n24022), .B(n24021), .Z(n44249) );
  NAND U44136 ( .A(n24024), .B(n24023), .Z(n44247) );
  AND U44137 ( .A(n24026), .B(n24025), .Z(n44245) );
  NAND U44138 ( .A(n24028), .B(n24027), .Z(n44243) );
  AND U44139 ( .A(n24030), .B(n24029), .Z(n44241) );
  ANDN U44140 ( .B(y[5566]), .A(x[5566]), .Z(n58004) );
  AND U44141 ( .A(n24032), .B(n24031), .Z(n44236) );
  ANDN U44142 ( .B(y[5564]), .A(x[5564]), .Z(n58001) );
  NOR U44143 ( .A(n58001), .B(n58003), .Z(n44234) );
  AND U44144 ( .A(n24034), .B(n24033), .Z(n44226) );
  NANDN U44145 ( .A(x[5560]), .B(y[5560]), .Z(n51345) );
  ANDN U44146 ( .B(n51345), .A(n57997), .Z(n44224) );
  AND U44147 ( .A(n24036), .B(n24035), .Z(n44215) );
  ANDN U44148 ( .B(y[5556]), .A(x[5556]), .Z(n57989) );
  NOR U44149 ( .A(n57989), .B(n57991), .Z(n44213) );
  AND U44150 ( .A(n24038), .B(n24037), .Z(n44205) );
  NANDN U44151 ( .A(x[5552]), .B(y[5552]), .Z(n51347) );
  ANDN U44152 ( .B(n51347), .A(n57986), .Z(n44203) );
  AND U44153 ( .A(n24040), .B(n24039), .Z(n44194) );
  ANDN U44154 ( .B(y[5548]), .A(x[5548]), .Z(n57978) );
  NOR U44155 ( .A(n57978), .B(n57980), .Z(n44192) );
  AND U44156 ( .A(n24042), .B(n24041), .Z(n44183) );
  NAND U44157 ( .A(n24043), .B(n51350), .Z(n44181) );
  AND U44158 ( .A(n24045), .B(n24044), .Z(n44179) );
  NANDN U44159 ( .A(x[5542]), .B(y[5542]), .Z(n57973) );
  NAND U44160 ( .A(n57973), .B(n24046), .Z(n44177) );
  AND U44161 ( .A(n24048), .B(n24047), .Z(n44175) );
  AND U44162 ( .A(n24050), .B(n24049), .Z(n44170) );
  NAND U44163 ( .A(n24052), .B(n24051), .Z(n44168) );
  AND U44164 ( .A(n24054), .B(n24053), .Z(n44166) );
  ANDN U44165 ( .B(y[5536]), .A(x[5536]), .Z(n57965) );
  NOR U44166 ( .A(n57965), .B(n24055), .Z(n44164) );
  AND U44167 ( .A(n24057), .B(n24056), .Z(n44156) );
  NANDN U44168 ( .A(x[5532]), .B(y[5532]), .Z(n57958) );
  AND U44169 ( .A(n57961), .B(n57958), .Z(n44154) );
  NAND U44170 ( .A(n24059), .B(n24058), .Z(n44152) );
  AND U44171 ( .A(n24061), .B(n24060), .Z(n44148) );
  AND U44172 ( .A(n24062), .B(n51351), .Z(n44146) );
  NAND U44173 ( .A(n24064), .B(n24063), .Z(n44144) );
  AND U44174 ( .A(n24066), .B(n24065), .Z(n44139) );
  NANDN U44175 ( .A(x[5524]), .B(y[5524]), .Z(n51355) );
  ANDN U44176 ( .B(n51355), .A(n57953), .Z(n44137) );
  AND U44177 ( .A(n24068), .B(n24067), .Z(n44128) );
  AND U44178 ( .A(n57948), .B(n57942), .Z(n44126) );
  NAND U44179 ( .A(n57944), .B(n24069), .Z(n44124) );
  AND U44180 ( .A(n24071), .B(n24070), .Z(n57946) );
  AND U44181 ( .A(n24073), .B(n24072), .Z(n44121) );
  NAND U44182 ( .A(n24075), .B(n24074), .Z(n44116) );
  AND U44183 ( .A(n24077), .B(n24076), .Z(n44111) );
  NAND U44184 ( .A(n24079), .B(n24078), .Z(n44107) );
  NANDN U44185 ( .A(x[5510]), .B(y[5510]), .Z(n44105) );
  IV U44186 ( .A(n24080), .Z(n51359) );
  AND U44187 ( .A(n24082), .B(n24081), .Z(n44102) );
  ANDN U44188 ( .B(y[5508]), .A(x[5508]), .Z(n57932) );
  NOR U44189 ( .A(n57932), .B(n24083), .Z(n44100) );
  AND U44190 ( .A(n24085), .B(n24084), .Z(n44092) );
  ANDN U44191 ( .B(y[5504]), .A(x[5504]), .Z(n57925) );
  NOR U44192 ( .A(n57927), .B(n57925), .Z(n44090) );
  AND U44193 ( .A(n24087), .B(n24086), .Z(n44081) );
  NANDN U44194 ( .A(x[5500]), .B(y[5500]), .Z(n51364) );
  NAND U44195 ( .A(n51364), .B(n24088), .Z(n44079) );
  AND U44196 ( .A(n24090), .B(n24089), .Z(n44077) );
  NANDN U44197 ( .A(x[5498]), .B(y[5498]), .Z(n57918) );
  NAND U44198 ( .A(n57918), .B(n57923), .Z(n44075) );
  AND U44199 ( .A(n24092), .B(n24091), .Z(n44073) );
  NAND U44200 ( .A(n57919), .B(n24093), .Z(n44071) );
  AND U44201 ( .A(n24095), .B(n24094), .Z(n44069) );
  ANDN U44202 ( .B(y[5494]), .A(x[5494]), .Z(n57914) );
  AND U44203 ( .A(n24097), .B(n24096), .Z(n44064) );
  ANDN U44204 ( .B(y[5492]), .A(x[5492]), .Z(n57911) );
  NOR U44205 ( .A(n57911), .B(n57913), .Z(n44062) );
  AND U44206 ( .A(n24099), .B(n24098), .Z(n44053) );
  NAND U44207 ( .A(n24101), .B(n24100), .Z(n44048) );
  AND U44208 ( .A(n24103), .B(n24102), .Z(n44043) );
  AND U44209 ( .A(n24104), .B(n57902), .Z(n44041) );
  AND U44210 ( .A(n24106), .B(n24105), .Z(n44039) );
  NAND U44211 ( .A(n24108), .B(n24107), .Z(n44037) );
  AND U44212 ( .A(n24110), .B(n24109), .Z(n44035) );
  NAND U44213 ( .A(n24112), .B(n24111), .Z(n44033) );
  AND U44214 ( .A(n24114), .B(n24113), .Z(n44031) );
  NANDN U44215 ( .A(x[5478]), .B(y[5478]), .Z(n57895) );
  NAND U44216 ( .A(n57895), .B(n24115), .Z(n44029) );
  AND U44217 ( .A(n24117), .B(n24116), .Z(n44027) );
  AND U44218 ( .A(n24119), .B(n24118), .Z(n44022) );
  NAND U44219 ( .A(n24121), .B(n24120), .Z(n44020) );
  AND U44220 ( .A(n24123), .B(n24122), .Z(n44018) );
  ANDN U44221 ( .B(y[5472]), .A(x[5472]), .Z(n57889) );
  NOR U44222 ( .A(n57889), .B(n24124), .Z(n44016) );
  AND U44223 ( .A(n24126), .B(n24125), .Z(n44008) );
  NANDN U44224 ( .A(x[5468]), .B(y[5468]), .Z(n57885) );
  IV U44225 ( .A(n24127), .Z(n51370) );
  ANDN U44226 ( .B(n57885), .A(n51370), .Z(n44006) );
  AND U44227 ( .A(n24129), .B(n24128), .Z(n43996) );
  NANDN U44228 ( .A(x[5464]), .B(y[5464]), .Z(n51374) );
  NAND U44229 ( .A(n51374), .B(n24130), .Z(n43994) );
  AND U44230 ( .A(n24132), .B(n24131), .Z(n43992) );
  NANDN U44231 ( .A(x[5462]), .B(y[5462]), .Z(n24133) );
  NAND U44232 ( .A(n24133), .B(n51373), .Z(n43990) );
  AND U44233 ( .A(n24135), .B(n24134), .Z(n43988) );
  ANDN U44234 ( .B(y[5460]), .A(x[5460]), .Z(n57876) );
  NOR U44235 ( .A(n57876), .B(n24136), .Z(n43986) );
  AND U44236 ( .A(n24138), .B(n24137), .Z(n43978) );
  ANDN U44237 ( .B(y[5456]), .A(x[5456]), .Z(n57873) );
  NOR U44238 ( .A(n57873), .B(n51375), .Z(n43976) );
  AND U44239 ( .A(n24140), .B(n24139), .Z(n43968) );
  NAND U44240 ( .A(n24142), .B(n24141), .Z(n43964) );
  NANDN U44241 ( .A(x[5450]), .B(y[5450]), .Z(n51378) );
  AND U44242 ( .A(n24144), .B(n24143), .Z(n43960) );
  ANDN U44243 ( .B(y[5448]), .A(x[5448]), .Z(n57861) );
  NOR U44244 ( .A(n57861), .B(n51377), .Z(n43958) );
  AND U44245 ( .A(n24146), .B(n24145), .Z(n43950) );
  ANDN U44246 ( .B(y[5444]), .A(x[5444]), .Z(n57854) );
  NOR U44247 ( .A(n57854), .B(n57857), .Z(n43948) );
  AND U44248 ( .A(n24148), .B(n24147), .Z(n43940) );
  ANDN U44249 ( .B(y[5440]), .A(x[5440]), .Z(n57851) );
  NOR U44250 ( .A(n57851), .B(n51379), .Z(n43938) );
  AND U44251 ( .A(n24150), .B(n24149), .Z(n43930) );
  ANDN U44252 ( .B(y[5436]), .A(x[5436]), .Z(n57843) );
  NOR U44253 ( .A(n57843), .B(n57846), .Z(n43928) );
  AND U44254 ( .A(n24152), .B(n24151), .Z(n43920) );
  ANDN U44255 ( .B(y[5432]), .A(x[5432]), .Z(n57840) );
  NOR U44256 ( .A(n57840), .B(n51381), .Z(n43918) );
  AND U44257 ( .A(n24154), .B(n24153), .Z(n43910) );
  NANDN U44258 ( .A(x[5428]), .B(y[5428]), .Z(n57833) );
  AND U44259 ( .A(n57833), .B(n57836), .Z(n43908) );
  NAND U44260 ( .A(n24156), .B(n24155), .Z(n43906) );
  AND U44261 ( .A(n24158), .B(n24157), .Z(n43901) );
  NANDN U44262 ( .A(x[5424]), .B(y[5424]), .Z(n57828) );
  AND U44263 ( .A(n57828), .B(n51383), .Z(n43899) );
  NANDN U44264 ( .A(x[5422]), .B(y[5422]), .Z(n57826) );
  AND U44265 ( .A(n24160), .B(n24159), .Z(n43891) );
  ANDN U44266 ( .B(y[5420]), .A(x[5420]), .Z(n57822) );
  NOR U44267 ( .A(n57822), .B(n57825), .Z(n43889) );
  AND U44268 ( .A(n24162), .B(n24161), .Z(n43881) );
  ANDN U44269 ( .B(y[5416]), .A(x[5416]), .Z(n57819) );
  NOR U44270 ( .A(n57819), .B(n51386), .Z(n43879) );
  AND U44271 ( .A(n24164), .B(n24163), .Z(n43871) );
  ANDN U44272 ( .B(y[5412]), .A(x[5412]), .Z(n57811) );
  NOR U44273 ( .A(n57811), .B(n57813), .Z(n43869) );
  AND U44274 ( .A(n24166), .B(n24165), .Z(n43861) );
  ANDN U44275 ( .B(y[5408]), .A(x[5408]), .Z(n57807) );
  NOR U44276 ( .A(n57807), .B(n51389), .Z(n43859) );
  AND U44277 ( .A(n24168), .B(n24167), .Z(n43850) );
  ANDN U44278 ( .B(y[5404]), .A(x[5404]), .Z(n57800) );
  NOR U44279 ( .A(n57800), .B(n57802), .Z(n43848) );
  AND U44280 ( .A(n24169), .B(n57799), .Z(n43842) );
  AND U44281 ( .A(n24171), .B(n24170), .Z(n43840) );
  NANDN U44282 ( .A(x[5400]), .B(y[5400]), .Z(n57795) );
  NAND U44283 ( .A(n57795), .B(n24172), .Z(n43838) );
  AND U44284 ( .A(n24174), .B(n24173), .Z(n43836) );
  NANDN U44285 ( .A(x[5398]), .B(y[5398]), .Z(n57792) );
  NAND U44286 ( .A(n57792), .B(n57794), .Z(n43834) );
  AND U44287 ( .A(n24176), .B(n24175), .Z(n43832) );
  NANDN U44288 ( .A(x[5396]), .B(y[5396]), .Z(n57788) );
  AND U44289 ( .A(n57791), .B(n57788), .Z(n43830) );
  NAND U44290 ( .A(n24178), .B(n24177), .Z(n43828) );
  NANDN U44291 ( .A(x[5394]), .B(y[5394]), .Z(n51393) );
  AND U44292 ( .A(n51393), .B(n57789), .Z(n43826) );
  AND U44293 ( .A(n24180), .B(n24179), .Z(n43824) );
  NANDN U44294 ( .A(x[5392]), .B(y[5392]), .Z(n57784) );
  ANDN U44295 ( .B(n57784), .A(n51391), .Z(n43822) );
  AND U44296 ( .A(n24182), .B(n24181), .Z(n43813) );
  ANDN U44297 ( .B(y[5388]), .A(x[5388]), .Z(n57777) );
  NOR U44298 ( .A(n57777), .B(n57780), .Z(n43811) );
  AND U44299 ( .A(n24184), .B(n24183), .Z(n43802) );
  ANDN U44300 ( .B(y[5384]), .A(x[5384]), .Z(n57774) );
  NOR U44301 ( .A(n57774), .B(n24185), .Z(n43800) );
  AND U44302 ( .A(n24187), .B(n24186), .Z(n43792) );
  ANDN U44303 ( .B(y[5380]), .A(x[5380]), .Z(n51396) );
  ANDN U44304 ( .B(n57770), .A(n51396), .Z(n43790) );
  AND U44305 ( .A(n24188), .B(n51395), .Z(n43784) );
  AND U44306 ( .A(n24190), .B(n24189), .Z(n43782) );
  NANDN U44307 ( .A(x[5376]), .B(y[5376]), .Z(n57762) );
  NAND U44308 ( .A(n57762), .B(n24191), .Z(n43780) );
  AND U44309 ( .A(n24193), .B(n24192), .Z(n43778) );
  NANDN U44310 ( .A(x[5374]), .B(y[5374]), .Z(n51399) );
  NAND U44311 ( .A(n51399), .B(n57763), .Z(n43776) );
  AND U44312 ( .A(n24195), .B(n24194), .Z(n43774) );
  NANDN U44313 ( .A(x[5372]), .B(y[5372]), .Z(n57759) );
  ANDN U44314 ( .B(n57759), .A(n51398), .Z(n43772) );
  AND U44315 ( .A(n24197), .B(n24196), .Z(n43763) );
  NANDN U44316 ( .A(x[5368]), .B(y[5368]), .Z(n24199) );
  NAND U44317 ( .A(n24199), .B(n24198), .Z(n43761) );
  AND U44318 ( .A(n24201), .B(n24200), .Z(n43759) );
  NANDN U44319 ( .A(x[5366]), .B(y[5366]), .Z(n24203) );
  NAND U44320 ( .A(n24203), .B(n24202), .Z(n43757) );
  AND U44321 ( .A(n24205), .B(n24204), .Z(n43755) );
  ANDN U44322 ( .B(y[5364]), .A(x[5364]), .Z(n57751) );
  NOR U44323 ( .A(n57751), .B(n24206), .Z(n43753) );
  AND U44324 ( .A(n24208), .B(n24207), .Z(n43745) );
  NANDN U44325 ( .A(x[5360]), .B(y[5360]), .Z(n57745) );
  IV U44326 ( .A(n24209), .Z(n51402) );
  ANDN U44327 ( .B(n57745), .A(n51402), .Z(n43743) );
  AND U44328 ( .A(n24211), .B(n24210), .Z(n43734) );
  AND U44329 ( .A(n24213), .B(n24212), .Z(n43729) );
  NAND U44330 ( .A(n24215), .B(n24214), .Z(n43727) );
  AND U44331 ( .A(n24217), .B(n24216), .Z(n43725) );
  ANDN U44332 ( .B(y[5352]), .A(x[5352]), .Z(n57739) );
  NOR U44333 ( .A(n57739), .B(n24218), .Z(n43723) );
  AND U44334 ( .A(n24220), .B(n24219), .Z(n43715) );
  NANDN U44335 ( .A(x[5348]), .B(y[5348]), .Z(n24221) );
  NAND U44336 ( .A(n51408), .B(n24221), .Z(n43713) );
  AND U44337 ( .A(n24223), .B(n24222), .Z(n43711) );
  NANDN U44338 ( .A(x[5346]), .B(y[5346]), .Z(n24225) );
  NAND U44339 ( .A(n24225), .B(n24224), .Z(n43709) );
  AND U44340 ( .A(n24227), .B(n24226), .Z(n43707) );
  NANDN U44341 ( .A(x[5344]), .B(y[5344]), .Z(n24229) );
  NAND U44342 ( .A(n24229), .B(n24228), .Z(n43705) );
  AND U44343 ( .A(n24231), .B(n24230), .Z(n43703) );
  NANDN U44344 ( .A(x[5342]), .B(y[5342]), .Z(n24233) );
  NAND U44345 ( .A(n24233), .B(n24232), .Z(n43701) );
  AND U44346 ( .A(n24235), .B(n24234), .Z(n43699) );
  ANDN U44347 ( .B(y[5340]), .A(x[5340]), .Z(n57726) );
  NOR U44348 ( .A(n57726), .B(n24236), .Z(n43697) );
  AND U44349 ( .A(n24237), .B(n57725), .Z(n43691) );
  AND U44350 ( .A(n24239), .B(n24238), .Z(n43689) );
  NANDN U44351 ( .A(x[5336]), .B(y[5336]), .Z(n51413) );
  NAND U44352 ( .A(n51413), .B(n24240), .Z(n43687) );
  AND U44353 ( .A(n24242), .B(n24241), .Z(n43685) );
  NANDN U44354 ( .A(x[5334]), .B(y[5334]), .Z(n57718) );
  IV U44355 ( .A(n24243), .Z(n57720) );
  NAND U44356 ( .A(n57718), .B(n57720), .Z(n43683) );
  AND U44357 ( .A(n24245), .B(n24244), .Z(n43681) );
  NAND U44358 ( .A(n57719), .B(n24246), .Z(n43679) );
  AND U44359 ( .A(n24248), .B(n24247), .Z(n43677) );
  ANDN U44360 ( .B(y[5330]), .A(x[5330]), .Z(n57714) );
  AND U44361 ( .A(n24250), .B(n24249), .Z(n43672) );
  ANDN U44362 ( .B(y[5328]), .A(x[5328]), .Z(n57709) );
  NOR U44363 ( .A(n57709), .B(n57713), .Z(n43670) );
  AND U44364 ( .A(n24252), .B(n24251), .Z(n43662) );
  ANDN U44365 ( .B(y[5324]), .A(x[5324]), .Z(n51415) );
  NOR U44366 ( .A(n51415), .B(n57706), .Z(n43660) );
  AND U44367 ( .A(n24254), .B(n24253), .Z(n43652) );
  IV U44368 ( .A(n24255), .Z(n57701) );
  NAND U44369 ( .A(n24257), .B(n24256), .Z(n43647) );
  AND U44370 ( .A(n24259), .B(n24258), .Z(n43642) );
  NANDN U44371 ( .A(x[5316]), .B(y[5316]), .Z(n57696) );
  IV U44372 ( .A(n24260), .Z(n51418) );
  AND U44373 ( .A(n57696), .B(n51418), .Z(n43640) );
  NAND U44374 ( .A(n24262), .B(n24261), .Z(n43638) );
  IV U44375 ( .A(n24263), .Z(n57695) );
  AND U44376 ( .A(n24264), .B(n57695), .Z(n43636) );
  AND U44377 ( .A(n24266), .B(n24265), .Z(n43634) );
  NANDN U44378 ( .A(x[5312]), .B(y[5312]), .Z(n51422) );
  AND U44379 ( .A(n51422), .B(n24267), .Z(n43632) );
  AND U44380 ( .A(n24268), .B(n51421), .Z(n43626) );
  NAND U44381 ( .A(n24270), .B(n24269), .Z(n43624) );
  NANDN U44382 ( .A(x[5308]), .B(y[5308]), .Z(n57688) );
  AND U44383 ( .A(n57688), .B(n24271), .Z(n43622) );
  NAND U44384 ( .A(n24273), .B(n24272), .Z(n43620) );
  NANDN U44385 ( .A(x[5306]), .B(y[5306]), .Z(n51425) );
  AND U44386 ( .A(n51425), .B(n57689), .Z(n43618) );
  AND U44387 ( .A(n24275), .B(n24274), .Z(n43616) );
  ANDN U44388 ( .B(y[5304]), .A(x[5304]), .Z(n57686) );
  NOR U44389 ( .A(n57686), .B(n51424), .Z(n43614) );
  IV U44390 ( .A(n24276), .Z(n57684) );
  AND U44391 ( .A(n24277), .B(n57684), .Z(n43608) );
  AND U44392 ( .A(n24279), .B(n24278), .Z(n43606) );
  NANDN U44393 ( .A(x[5300]), .B(y[5300]), .Z(n51428) );
  ANDN U44394 ( .B(n51428), .A(n24280), .Z(n43604) );
  IV U44395 ( .A(n24281), .Z(n51427) );
  AND U44396 ( .A(n24282), .B(n51427), .Z(n43598) );
  AND U44397 ( .A(n24284), .B(n24283), .Z(n43596) );
  NAND U44398 ( .A(n24286), .B(n24285), .Z(n43594) );
  AND U44399 ( .A(n24288), .B(n24287), .Z(n43592) );
  NAND U44400 ( .A(n24290), .B(n24289), .Z(n43590) );
  AND U44401 ( .A(n24292), .B(n24291), .Z(n43588) );
  NANDN U44402 ( .A(x[5292]), .B(y[5292]), .Z(n57674) );
  NAND U44403 ( .A(n57674), .B(n24293), .Z(n43586) );
  XNOR U44404 ( .A(x[5292]), .B(y[5292]), .Z(n24295) );
  AND U44405 ( .A(n24295), .B(n24294), .Z(n43584) );
  NAND U44406 ( .A(n24296), .B(n57673), .Z(n43582) );
  AND U44407 ( .A(n24298), .B(n24297), .Z(n43580) );
  AND U44408 ( .A(n24300), .B(n24299), .Z(n43574) );
  NAND U44409 ( .A(n24302), .B(n24301), .Z(n43572) );
  AND U44410 ( .A(n24304), .B(n24303), .Z(n43570) );
  ANDN U44411 ( .B(y[5284]), .A(x[5284]), .Z(n57663) );
  NOR U44412 ( .A(n57663), .B(n24305), .Z(n43568) );
  AND U44413 ( .A(n24306), .B(n57664), .Z(n43562) );
  AND U44414 ( .A(n24308), .B(n24307), .Z(n43560) );
  NAND U44415 ( .A(n24310), .B(n24309), .Z(n43558) );
  AND U44416 ( .A(n24312), .B(n24311), .Z(n43556) );
  ANDN U44417 ( .B(y[5278]), .A(x[5278]), .Z(n57657) );
  AND U44418 ( .A(n24314), .B(n24313), .Z(n43551) );
  NAND U44419 ( .A(n24315), .B(n57658), .Z(n43549) );
  AND U44420 ( .A(n24317), .B(n24316), .Z(n43547) );
  NAND U44421 ( .A(n24319), .B(n24318), .Z(n43545) );
  AND U44422 ( .A(n24321), .B(n24320), .Z(n43543) );
  NANDN U44423 ( .A(x[5272]), .B(y[5272]), .Z(n57651) );
  AND U44424 ( .A(n57651), .B(n24322), .Z(n43541) );
  ANDN U44425 ( .B(y[5270]), .A(x[5270]), .Z(n43534) );
  AND U44426 ( .A(n24324), .B(n24323), .Z(n43532) );
  NAND U44427 ( .A(n24326), .B(n24325), .Z(n43530) );
  AND U44428 ( .A(n24328), .B(n24327), .Z(n43528) );
  NANDN U44429 ( .A(x[5266]), .B(y[5266]), .Z(n57643) );
  NAND U44430 ( .A(n57643), .B(n24329), .Z(n43526) );
  AND U44431 ( .A(n24331), .B(n24330), .Z(n43524) );
  NANDN U44432 ( .A(x[5264]), .B(y[5264]), .Z(n51438) );
  IV U44433 ( .A(n24332), .Z(n57642) );
  ANDN U44434 ( .B(n51438), .A(n57642), .Z(n43522) );
  AND U44435 ( .A(n24334), .B(n24333), .Z(n43513) );
  NANDN U44436 ( .A(x[5260]), .B(y[5260]), .Z(n57636) );
  ANDN U44437 ( .B(n57636), .A(n57638), .Z(n43511) );
  IV U44438 ( .A(n24335), .Z(n57635) );
  AND U44439 ( .A(n24336), .B(n57635), .Z(n43505) );
  AND U44440 ( .A(n24338), .B(n24337), .Z(n43503) );
  ANDN U44441 ( .B(y[5256]), .A(x[5256]), .Z(n57631) );
  NOR U44442 ( .A(n57631), .B(n24339), .Z(n43501) );
  AND U44443 ( .A(n24341), .B(n24340), .Z(n43492) );
  NANDN U44444 ( .A(x[5252]), .B(y[5252]), .Z(n57624) );
  IV U44445 ( .A(n24342), .Z(n57626) );
  NAND U44446 ( .A(n57624), .B(n57626), .Z(n43490) );
  AND U44447 ( .A(n24344), .B(n24343), .Z(n43488) );
  NAND U44448 ( .A(n57625), .B(n24345), .Z(n43486) );
  AND U44449 ( .A(n24347), .B(n24346), .Z(n43484) );
  NAND U44450 ( .A(n24349), .B(n24348), .Z(n43479) );
  AND U44451 ( .A(n24351), .B(n24350), .Z(n43474) );
  NAND U44452 ( .A(n24352), .B(n57618), .Z(n43472) );
  AND U44453 ( .A(n24354), .B(n24353), .Z(n43470) );
  NANDN U44454 ( .A(x[5242]), .B(y[5242]), .Z(n57612) );
  NAND U44455 ( .A(n57612), .B(n24355), .Z(n43468) );
  AND U44456 ( .A(n24357), .B(n24356), .Z(n43466) );
  ANDN U44457 ( .B(y[5240]), .A(x[5240]), .Z(n57609) );
  NOR U44458 ( .A(n57609), .B(n57611), .Z(n43464) );
  AND U44459 ( .A(n24359), .B(n24358), .Z(n43456) );
  ANDN U44460 ( .B(y[5236]), .A(x[5236]), .Z(n57602) );
  NOR U44461 ( .A(n57602), .B(n57606), .Z(n43454) );
  AND U44462 ( .A(n24360), .B(n57603), .Z(n43448) );
  AND U44463 ( .A(n24362), .B(n24361), .Z(n43446) );
  ANDN U44464 ( .B(y[5232]), .A(x[5232]), .Z(n57597) );
  NOR U44465 ( .A(n57597), .B(n24363), .Z(n43444) );
  AND U44466 ( .A(n24365), .B(n24364), .Z(n43436) );
  NAND U44467 ( .A(n51441), .B(n24366), .Z(n43434) );
  AND U44468 ( .A(n24368), .B(n24367), .Z(n43432) );
  NANDN U44469 ( .A(x[5226]), .B(y[5226]), .Z(n57590) );
  NAND U44470 ( .A(n57590), .B(n24369), .Z(n43430) );
  AND U44471 ( .A(n24371), .B(n24370), .Z(n43428) );
  ANDN U44472 ( .B(y[5224]), .A(x[5224]), .Z(n51445) );
  NOR U44473 ( .A(n51445), .B(n57591), .Z(n43426) );
  AND U44474 ( .A(n24373), .B(n24372), .Z(n43417) );
  ANDN U44475 ( .B(y[5220]), .A(x[5220]), .Z(n57585) );
  NOR U44476 ( .A(n57585), .B(n24374), .Z(n43415) );
  AND U44477 ( .A(n24376), .B(n24375), .Z(n43406) );
  NANDN U44478 ( .A(x[5216]), .B(y[5216]), .Z(n51449) );
  NAND U44479 ( .A(n51449), .B(n24377), .Z(n43404) );
  AND U44480 ( .A(n24379), .B(n24378), .Z(n43402) );
  NANDN U44481 ( .A(x[5214]), .B(y[5214]), .Z(n57578) );
  NAND U44482 ( .A(n57578), .B(n57581), .Z(n43400) );
  AND U44483 ( .A(n24381), .B(n24380), .Z(n43398) );
  ANDN U44484 ( .B(y[5212]), .A(x[5212]), .Z(n51451) );
  ANDN U44485 ( .B(n57579), .A(n51451), .Z(n43396) );
  AND U44486 ( .A(n24383), .B(n24382), .Z(n43388) );
  ANDN U44487 ( .B(y[5208]), .A(x[5208]), .Z(n57571) );
  NOR U44488 ( .A(n57572), .B(n57571), .Z(n43386) );
  AND U44489 ( .A(n24384), .B(n57570), .Z(n43380) );
  AND U44490 ( .A(n24386), .B(n24385), .Z(n43378) );
  NAND U44491 ( .A(n24388), .B(n24387), .Z(n43376) );
  AND U44492 ( .A(n24390), .B(n24389), .Z(n43374) );
  NANDN U44493 ( .A(x[5202]), .B(y[5202]), .Z(n51455) );
  NAND U44494 ( .A(n51455), .B(n24391), .Z(n43372) );
  AND U44495 ( .A(n24393), .B(n24392), .Z(n43370) );
  NANDN U44496 ( .A(x[5200]), .B(y[5200]), .Z(n51458) );
  ANDN U44497 ( .B(n51458), .A(n51456), .Z(n43368) );
  AND U44498 ( .A(n24395), .B(n24394), .Z(n43359) );
  ANDN U44499 ( .B(y[5196]), .A(x[5196]), .Z(n57559) );
  NOR U44500 ( .A(n57559), .B(n57561), .Z(n43357) );
  AND U44501 ( .A(n24397), .B(n24396), .Z(n43348) );
  NANDN U44502 ( .A(x[5192]), .B(y[5192]), .Z(n51461) );
  AND U44503 ( .A(n24399), .B(n24398), .Z(n43344) );
  NAND U44504 ( .A(n51460), .B(n24400), .Z(n43342) );
  AND U44505 ( .A(n24402), .B(n24401), .Z(n43340) );
  NANDN U44506 ( .A(x[5188]), .B(y[5188]), .Z(n51464) );
  ANDN U44507 ( .B(n51464), .A(n24403), .Z(n43338) );
  IV U44508 ( .A(n24404), .Z(n51463) );
  AND U44509 ( .A(n24405), .B(n51463), .Z(n43332) );
  AND U44510 ( .A(n24407), .B(n24406), .Z(n43330) );
  NANDN U44511 ( .A(x[5184]), .B(y[5184]), .Z(n57547) );
  AND U44512 ( .A(n57547), .B(n24408), .Z(n43328) );
  IV U44513 ( .A(n24409), .Z(n57546) );
  ANDN U44514 ( .B(y[5182]), .A(x[5182]), .Z(n57544) );
  AND U44515 ( .A(n24411), .B(n24410), .Z(n43320) );
  ANDN U44516 ( .B(y[5180]), .A(x[5180]), .Z(n57540) );
  NOR U44517 ( .A(n57543), .B(n57540), .Z(n43318) );
  AND U44518 ( .A(n24412), .B(n57539), .Z(n43312) );
  AND U44519 ( .A(n24414), .B(n24413), .Z(n43310) );
  ANDN U44520 ( .B(y[5176]), .A(x[5176]), .Z(n57535) );
  NOR U44521 ( .A(n57535), .B(n24415), .Z(n43308) );
  AND U44522 ( .A(n24417), .B(n24416), .Z(n43299) );
  ANDN U44523 ( .B(y[5172]), .A(x[5172]), .Z(n51467) );
  NOR U44524 ( .A(n51467), .B(n57532), .Z(n43297) );
  AND U44525 ( .A(n24419), .B(n24418), .Z(n43289) );
  NAND U44526 ( .A(n24420), .B(n57527), .Z(n43287) );
  AND U44527 ( .A(n24422), .B(n24421), .Z(n43285) );
  NANDN U44528 ( .A(x[5166]), .B(y[5166]), .Z(n51469) );
  AND U44529 ( .A(n24424), .B(n24423), .Z(n43280) );
  IV U44530 ( .A(n24425), .Z(n51468) );
  NANDN U44531 ( .A(x[5164]), .B(y[5164]), .Z(n57521) );
  NAND U44532 ( .A(n51468), .B(n57521), .Z(n43278) );
  AND U44533 ( .A(n24427), .B(n24426), .Z(n43276) );
  NAND U44534 ( .A(n24428), .B(n57520), .Z(n43274) );
  AND U44535 ( .A(n24430), .B(n24429), .Z(n43272) );
  NAND U44536 ( .A(n24432), .B(n24431), .Z(n43266) );
  AND U44537 ( .A(n24434), .B(n24433), .Z(n43261) );
  NAND U44538 ( .A(n24436), .B(n24435), .Z(n43257) );
  AND U44539 ( .A(n24437), .B(n57510), .Z(n43255) );
  NAND U44540 ( .A(n24439), .B(n24438), .Z(n43253) );
  NANDN U44541 ( .A(x[5152]), .B(y[5152]), .Z(n57506) );
  AND U44542 ( .A(n24440), .B(n57506), .Z(n43251) );
  AND U44543 ( .A(n24442), .B(n24441), .Z(n43242) );
  NANDN U44544 ( .A(x[5148]), .B(y[5148]), .Z(n51474) );
  ANDN U44545 ( .B(n51474), .A(n24443), .Z(n43240) );
  XNOR U44546 ( .A(x[5146]), .B(y[5146]), .Z(n24445) );
  AND U44547 ( .A(n24445), .B(n24444), .Z(n43231) );
  NAND U44548 ( .A(n24446), .B(n57500), .Z(n43229) );
  AND U44549 ( .A(n24448), .B(n24447), .Z(n43227) );
  NANDN U44550 ( .A(x[5142]), .B(y[5142]), .Z(n24450) );
  NAND U44551 ( .A(n24450), .B(n24449), .Z(n43225) );
  AND U44552 ( .A(n24452), .B(n24451), .Z(n43223) );
  NAND U44553 ( .A(n24454), .B(n24453), .Z(n43221) );
  AND U44554 ( .A(n24456), .B(n24455), .Z(n43219) );
  NANDN U44555 ( .A(x[5138]), .B(y[5138]), .Z(n57492) );
  NAND U44556 ( .A(n57492), .B(n24457), .Z(n43217) );
  AND U44557 ( .A(n24459), .B(n24458), .Z(n43215) );
  NANDN U44558 ( .A(x[5136]), .B(y[5136]), .Z(n51478) );
  IV U44559 ( .A(n24460), .Z(n57491) );
  ANDN U44560 ( .B(n51478), .A(n57491), .Z(n43213) );
  AND U44561 ( .A(n24462), .B(n24461), .Z(n43204) );
  ANDN U44562 ( .B(y[5132]), .A(x[5132]), .Z(n57485) );
  NOR U44563 ( .A(n57485), .B(n57487), .Z(n43202) );
  AND U44564 ( .A(n24464), .B(n24463), .Z(n43193) );
  ANDN U44565 ( .B(y[5128]), .A(x[5128]), .Z(n51481) );
  NOR U44566 ( .A(n51481), .B(n57481), .Z(n43191) );
  AND U44567 ( .A(n24466), .B(n24465), .Z(n43182) );
  NANDN U44568 ( .A(x[5124]), .B(y[5124]), .Z(n24468) );
  NAND U44569 ( .A(n24468), .B(n24467), .Z(n43180) );
  AND U44570 ( .A(n24470), .B(n24469), .Z(n43178) );
  NANDN U44571 ( .A(x[5122]), .B(y[5122]), .Z(n24472) );
  NAND U44572 ( .A(n24472), .B(n24471), .Z(n43176) );
  AND U44573 ( .A(n24474), .B(n24473), .Z(n43174) );
  NAND U44574 ( .A(n24476), .B(n24475), .Z(n43172) );
  AND U44575 ( .A(n24478), .B(n24477), .Z(n43170) );
  NANDN U44576 ( .A(x[5118]), .B(y[5118]), .Z(n57467) );
  NAND U44577 ( .A(n57467), .B(n24479), .Z(n43168) );
  AND U44578 ( .A(n24481), .B(n24480), .Z(n43166) );
  NANDN U44579 ( .A(x[5116]), .B(y[5116]), .Z(n51483) );
  AND U44580 ( .A(n51483), .B(n57469), .Z(n43164) );
  NAND U44581 ( .A(n24483), .B(n24482), .Z(n43162) );
  AND U44582 ( .A(n24485), .B(n24484), .Z(n43158) );
  ANDN U44583 ( .B(y[5112]), .A(x[5112]), .Z(n57460) );
  NOR U44584 ( .A(n57460), .B(n57462), .Z(n43156) );
  AND U44585 ( .A(n24487), .B(n24486), .Z(n43147) );
  NANDN U44586 ( .A(x[5108]), .B(y[5108]), .Z(n51487) );
  AND U44587 ( .A(n51487), .B(n51484), .Z(n43145) );
  NAND U44588 ( .A(n24489), .B(n24488), .Z(n43143) );
  AND U44589 ( .A(n24491), .B(n24490), .Z(n43139) );
  NANDN U44590 ( .A(x[5104]), .B(y[5104]), .Z(n24492) );
  NAND U44591 ( .A(n24492), .B(n57454), .Z(n43137) );
  AND U44592 ( .A(n24494), .B(n24493), .Z(n43135) );
  NANDN U44593 ( .A(x[5102]), .B(y[5102]), .Z(n24496) );
  NAND U44594 ( .A(n24496), .B(n24495), .Z(n43133) );
  AND U44595 ( .A(n24498), .B(n24497), .Z(n43131) );
  NAND U44596 ( .A(n24500), .B(n24499), .Z(n43125) );
  AND U44597 ( .A(n24502), .B(n24501), .Z(n43119) );
  NANDN U44598 ( .A(x[5096]), .B(y[5096]), .Z(n51489) );
  ANDN U44599 ( .B(n51489), .A(n24503), .Z(n43117) );
  AND U44600 ( .A(n24505), .B(n24504), .Z(n43108) );
  NAND U44601 ( .A(n24506), .B(n57441), .Z(n43106) );
  AND U44602 ( .A(n24508), .B(n24507), .Z(n43104) );
  NAND U44603 ( .A(n24510), .B(n24509), .Z(n43102) );
  AND U44604 ( .A(n24512), .B(n24511), .Z(n43100) );
  NANDN U44605 ( .A(x[5088]), .B(y[5088]), .Z(n57433) );
  NAND U44606 ( .A(n57433), .B(n24513), .Z(n43098) );
  AND U44607 ( .A(n24515), .B(n24514), .Z(n43096) );
  NANDN U44608 ( .A(x[5086]), .B(y[5086]), .Z(n57430) );
  NAND U44609 ( .A(n57430), .B(n57432), .Z(n43094) );
  AND U44610 ( .A(n24517), .B(n24516), .Z(n43092) );
  ANDN U44611 ( .B(y[5084]), .A(x[5084]), .Z(n57428) );
  NOR U44612 ( .A(n57429), .B(n57428), .Z(n43090) );
  AND U44613 ( .A(n24519), .B(n24518), .Z(n43082) );
  ANDN U44614 ( .B(y[5080]), .A(x[5080]), .Z(n57424) );
  NOR U44615 ( .A(n57424), .B(n51492), .Z(n43080) );
  AND U44616 ( .A(n24520), .B(n57423), .Z(n43074) );
  AND U44617 ( .A(n24522), .B(n24521), .Z(n43072) );
  ANDN U44618 ( .B(y[5076]), .A(x[5076]), .Z(n51493) );
  NOR U44619 ( .A(n51493), .B(n24523), .Z(n43070) );
  AND U44620 ( .A(n24524), .B(n51494), .Z(n43064) );
  AND U44621 ( .A(n24526), .B(n24525), .Z(n43062) );
  NANDN U44622 ( .A(x[5072]), .B(y[5072]), .Z(n57414) );
  NAND U44623 ( .A(n57414), .B(n24527), .Z(n43060) );
  AND U44624 ( .A(n24529), .B(n24528), .Z(n43058) );
  NAND U44625 ( .A(n57415), .B(n24530), .Z(n43056) );
  AND U44626 ( .A(n24532), .B(n24531), .Z(n43054) );
  ANDN U44627 ( .B(y[5068]), .A(x[5068]), .Z(n57410) );
  NOR U44628 ( .A(n57410), .B(n24533), .Z(n43052) );
  AND U44629 ( .A(n24535), .B(n24534), .Z(n43044) );
  ANDN U44630 ( .B(y[5064]), .A(x[5064]), .Z(n57402) );
  NOR U44631 ( .A(n57402), .B(n57405), .Z(n43042) );
  AND U44632 ( .A(n24537), .B(n24536), .Z(n43034) );
  ANDN U44633 ( .B(y[5060]), .A(x[5060]), .Z(n57399) );
  NOR U44634 ( .A(n57399), .B(n51496), .Z(n43032) );
  AND U44635 ( .A(n24538), .B(n57398), .Z(n43026) );
  AND U44636 ( .A(n24540), .B(n24539), .Z(n43024) );
  NAND U44637 ( .A(n24542), .B(n24541), .Z(n43022) );
  AND U44638 ( .A(n24544), .B(n24543), .Z(n43020) );
  NANDN U44639 ( .A(x[5054]), .B(y[5054]), .Z(n57392) );
  NAND U44640 ( .A(n57392), .B(n24545), .Z(n43018) );
  AND U44641 ( .A(n24547), .B(n24546), .Z(n43016) );
  ANDN U44642 ( .B(y[5052]), .A(x[5052]), .Z(n57388) );
  NOR U44643 ( .A(n57388), .B(n57390), .Z(n43014) );
  AND U44644 ( .A(n24549), .B(n24548), .Z(n43006) );
  NAND U44645 ( .A(n51497), .B(n24550), .Z(n43004) );
  AND U44646 ( .A(n24552), .B(n24551), .Z(n43002) );
  NANDN U44647 ( .A(x[5046]), .B(y[5046]), .Z(n57381) );
  NAND U44648 ( .A(n57381), .B(n24553), .Z(n43000) );
  AND U44649 ( .A(n24555), .B(n24554), .Z(n42998) );
  NAND U44650 ( .A(n57382), .B(n24556), .Z(n42996) );
  AND U44651 ( .A(n24558), .B(n24557), .Z(n42994) );
  ANDN U44652 ( .B(y[5042]), .A(x[5042]), .Z(n57378) );
  AND U44653 ( .A(n24560), .B(n24559), .Z(n42989) );
  NAND U44654 ( .A(n24561), .B(n57377), .Z(n42987) );
  AND U44655 ( .A(n24563), .B(n24562), .Z(n42985) );
  NANDN U44656 ( .A(x[5038]), .B(y[5038]), .Z(n51502) );
  NAND U44657 ( .A(n51502), .B(n24564), .Z(n42983) );
  AND U44658 ( .A(n24566), .B(n24565), .Z(n42981) );
  AND U44659 ( .A(n24568), .B(n24567), .Z(n42976) );
  NAND U44660 ( .A(n24570), .B(n24569), .Z(n42974) );
  AND U44661 ( .A(n24572), .B(n24571), .Z(n42972) );
  NAND U44662 ( .A(n24574), .B(n24573), .Z(n42970) );
  AND U44663 ( .A(n24576), .B(n24575), .Z(n42968) );
  NANDN U44664 ( .A(x[5030]), .B(y[5030]), .Z(n57366) );
  NAND U44665 ( .A(n57366), .B(n24577), .Z(n42966) );
  AND U44666 ( .A(n24579), .B(n24578), .Z(n42964) );
  ANDN U44667 ( .B(y[5028]), .A(x[5028]), .Z(n57361) );
  NOR U44668 ( .A(n57361), .B(n57365), .Z(n42962) );
  AND U44669 ( .A(n24581), .B(n24580), .Z(n42953) );
  AND U44670 ( .A(n24583), .B(n24582), .Z(n42948) );
  AND U44671 ( .A(n24585), .B(n24584), .Z(n42944) );
  NAND U44672 ( .A(n57354), .B(n24586), .Z(n42942) );
  AND U44673 ( .A(n24588), .B(n24587), .Z(n42940) );
  ANDN U44674 ( .B(y[5018]), .A(x[5018]), .Z(n57351) );
  AND U44675 ( .A(n24590), .B(n24589), .Z(n42935) );
  ANDN U44676 ( .B(y[5016]), .A(x[5016]), .Z(n57345) );
  NOR U44677 ( .A(n57349), .B(n57345), .Z(n42933) );
  AND U44678 ( .A(n24591), .B(n57346), .Z(n42927) );
  AND U44679 ( .A(n24593), .B(n24592), .Z(n42925) );
  NANDN U44680 ( .A(x[5012]), .B(y[5012]), .Z(n57341) );
  NAND U44681 ( .A(n57341), .B(n24594), .Z(n42923) );
  AND U44682 ( .A(n24596), .B(n24595), .Z(n42921) );
  IV U44683 ( .A(n24597), .Z(n57340) );
  NANDN U44684 ( .A(x[5010]), .B(y[5010]), .Z(n57338) );
  NAND U44685 ( .A(n57340), .B(n57338), .Z(n42919) );
  AND U44686 ( .A(n24599), .B(n24598), .Z(n42917) );
  ANDN U44687 ( .B(y[5008]), .A(x[5008]), .Z(n57335) );
  NOR U44688 ( .A(n57335), .B(n57337), .Z(n42915) );
  AND U44689 ( .A(n24600), .B(n57336), .Z(n42909) );
  AND U44690 ( .A(n24602), .B(n24601), .Z(n42907) );
  ANDN U44691 ( .B(y[5004]), .A(x[5004]), .Z(n57332) );
  NOR U44692 ( .A(n57332), .B(n24603), .Z(n42905) );
  AND U44693 ( .A(n24605), .B(n24604), .Z(n42896) );
  AND U44694 ( .A(n24606), .B(n57329), .Z(n42894) );
  NAND U44695 ( .A(n24608), .B(n24607), .Z(n42892) );
  NANDN U44696 ( .A(x[4998]), .B(y[4998]), .Z(n57324) );
  AND U44697 ( .A(n24610), .B(n24609), .Z(n42887) );
  NANDN U44698 ( .A(x[4996]), .B(y[4996]), .Z(n57321) );
  AND U44699 ( .A(n57321), .B(n57323), .Z(n42885) );
  AND U44700 ( .A(n24612), .B(n24611), .Z(n42875) );
  ANDN U44701 ( .B(y[4992]), .A(x[4992]), .Z(n57316) );
  NOR U44702 ( .A(n57316), .B(n24613), .Z(n42873) );
  AND U44703 ( .A(n24615), .B(n24614), .Z(n42864) );
  ANDN U44704 ( .B(y[4988]), .A(x[4988]), .Z(n57309) );
  NOR U44705 ( .A(n57311), .B(n57309), .Z(n42862) );
  AND U44706 ( .A(n24617), .B(n24616), .Z(n42854) );
  ANDN U44707 ( .B(y[4984]), .A(x[4984]), .Z(n57304) );
  NOR U44708 ( .A(n57304), .B(n57306), .Z(n42852) );
  AND U44709 ( .A(n24619), .B(n24618), .Z(n42844) );
  ANDN U44710 ( .B(y[4980]), .A(x[4980]), .Z(n51512) );
  NOR U44711 ( .A(n57299), .B(n51512), .Z(n42842) );
  AND U44712 ( .A(n24621), .B(n24620), .Z(n42833) );
  NAND U44713 ( .A(n24623), .B(n24622), .Z(n42831) );
  AND U44714 ( .A(n24625), .B(n24624), .Z(n42829) );
  NANDN U44715 ( .A(x[4974]), .B(y[4974]), .Z(n24627) );
  NAND U44716 ( .A(n24627), .B(n24626), .Z(n42827) );
  AND U44717 ( .A(n24629), .B(n24628), .Z(n42825) );
  NAND U44718 ( .A(n24631), .B(n24630), .Z(n42823) );
  AND U44719 ( .A(n24633), .B(n24632), .Z(n42821) );
  NANDN U44720 ( .A(x[4970]), .B(y[4970]), .Z(n57287) );
  NAND U44721 ( .A(n57287), .B(n24634), .Z(n42819) );
  AND U44722 ( .A(n24636), .B(n24635), .Z(n42817) );
  NAND U44723 ( .A(n24637), .B(n57288), .Z(n42815) );
  AND U44724 ( .A(n24639), .B(n24638), .Z(n42813) );
  ANDN U44725 ( .B(y[4966]), .A(x[4966]), .Z(n57281) );
  AND U44726 ( .A(n24641), .B(n24640), .Z(n42808) );
  NANDN U44727 ( .A(x[4964]), .B(y[4964]), .Z(n57278) );
  ANDN U44728 ( .B(n57278), .A(n57280), .Z(n42806) );
  AND U44729 ( .A(n24643), .B(n24642), .Z(n42797) );
  NANDN U44730 ( .A(x[4960]), .B(y[4960]), .Z(n51518) );
  AND U44731 ( .A(n51518), .B(n51516), .Z(n42795) );
  NAND U44732 ( .A(n24645), .B(n24644), .Z(n42793) );
  AND U44733 ( .A(n24647), .B(n24646), .Z(n42789) );
  ANDN U44734 ( .B(y[4956]), .A(x[4956]), .Z(n57270) );
  NOR U44735 ( .A(n57270), .B(n57272), .Z(n42787) );
  XNOR U44736 ( .A(x[4954]), .B(y[4954]), .Z(n24649) );
  AND U44737 ( .A(n24649), .B(n24648), .Z(n42778) );
  NAND U44738 ( .A(n24650), .B(n57266), .Z(n42776) );
  AND U44739 ( .A(n24652), .B(n24651), .Z(n42774) );
  NANDN U44740 ( .A(x[4950]), .B(y[4950]), .Z(n51520) );
  NAND U44741 ( .A(n51520), .B(n24653), .Z(n42772) );
  AND U44742 ( .A(n24655), .B(n24654), .Z(n42770) );
  ANDN U44743 ( .B(y[4948]), .A(x[4948]), .Z(n57258) );
  NOR U44744 ( .A(n57261), .B(n57258), .Z(n42768) );
  AND U44745 ( .A(n24657), .B(n24656), .Z(n42760) );
  ANDN U44746 ( .B(y[4944]), .A(x[4944]), .Z(n57255) );
  NOR U44747 ( .A(n57255), .B(n51521), .Z(n42758) );
  AND U44748 ( .A(n24659), .B(n24658), .Z(n42750) );
  NANDN U44749 ( .A(x[4940]), .B(y[4940]), .Z(n57247) );
  AND U44750 ( .A(n57250), .B(n57247), .Z(n42748) );
  AND U44751 ( .A(n24660), .B(n57248), .Z(n42742) );
  NAND U44752 ( .A(n24662), .B(n24661), .Z(n42740) );
  NAND U44753 ( .A(n24664), .B(n24663), .Z(n42735) );
  NANDN U44754 ( .A(x[4934]), .B(y[4934]), .Z(n57241) );
  IV U44755 ( .A(n24665), .Z(n57243) );
  AND U44756 ( .A(n57241), .B(n57243), .Z(n42733) );
  NAND U44757 ( .A(n24667), .B(n24666), .Z(n42731) );
  AND U44758 ( .A(n24668), .B(n57240), .Z(n42729) );
  AND U44759 ( .A(n24670), .B(n24669), .Z(n42727) );
  AND U44760 ( .A(n24672), .B(n24671), .Z(n42722) );
  ANDN U44761 ( .B(y[4928]), .A(x[4928]), .Z(n57233) );
  NAND U44762 ( .A(n24674), .B(n24673), .Z(n42718) );
  NANDN U44763 ( .A(x[4926]), .B(y[4926]), .Z(n51526) );
  AND U44764 ( .A(n24676), .B(n24675), .Z(n42714) );
  AND U44765 ( .A(n24677), .B(n57228), .Z(n42705) );
  NAND U44766 ( .A(n24679), .B(n24678), .Z(n42703) );
  AND U44767 ( .A(n24681), .B(n24680), .Z(n42701) );
  NAND U44768 ( .A(n24683), .B(n24682), .Z(n42699) );
  NANDN U44769 ( .A(x[4918]), .B(y[4918]), .Z(n51530) );
  AND U44770 ( .A(n24685), .B(n24684), .Z(n42694) );
  NAND U44771 ( .A(n24687), .B(n24686), .Z(n42690) );
  NANDN U44772 ( .A(x[4914]), .B(y[4914]), .Z(n57217) );
  AND U44773 ( .A(n24689), .B(n24688), .Z(n42686) );
  AND U44774 ( .A(n24690), .B(n57218), .Z(n42684) );
  AND U44775 ( .A(n24692), .B(n24691), .Z(n42678) );
  NAND U44776 ( .A(n24694), .B(n24693), .Z(n42676) );
  AND U44777 ( .A(n24696), .B(n24695), .Z(n42674) );
  NAND U44778 ( .A(n24698), .B(n24697), .Z(n42672) );
  NANDN U44779 ( .A(x[4906]), .B(y[4906]), .Z(n51534) );
  AND U44780 ( .A(n51534), .B(n24699), .Z(n42670) );
  NAND U44781 ( .A(n24701), .B(n24700), .Z(n42668) );
  IV U44782 ( .A(n24702), .Z(n51533) );
  AND U44783 ( .A(n24703), .B(n51533), .Z(n42666) );
  AND U44784 ( .A(n24705), .B(n24704), .Z(n42660) );
  NAND U44785 ( .A(n24707), .B(n24706), .Z(n42658) );
  AND U44786 ( .A(n24709), .B(n24708), .Z(n42656) );
  AND U44787 ( .A(n24711), .B(n24710), .Z(n42650) );
  NAND U44788 ( .A(n24713), .B(n24712), .Z(n42648) );
  AND U44789 ( .A(n24715), .B(n24714), .Z(n42646) );
  AND U44790 ( .A(n24717), .B(n24716), .Z(n42640) );
  NAND U44791 ( .A(n24719), .B(n24718), .Z(n42638) );
  AND U44792 ( .A(n24721), .B(n24720), .Z(n42636) );
  AND U44793 ( .A(n24723), .B(n24722), .Z(n42630) );
  NAND U44794 ( .A(n24725), .B(n24724), .Z(n42628) );
  AND U44795 ( .A(n24727), .B(n24726), .Z(n42626) );
  NAND U44796 ( .A(n24729), .B(n24728), .Z(n42624) );
  NANDN U44797 ( .A(x[4886]), .B(y[4886]), .Z(n57190) );
  AND U44798 ( .A(n24731), .B(n24730), .Z(n42619) );
  AND U44799 ( .A(n24732), .B(n57189), .Z(n42617) );
  NAND U44800 ( .A(n24734), .B(n24733), .Z(n42615) );
  NANDN U44801 ( .A(x[4882]), .B(y[4882]), .Z(n24736) );
  AND U44802 ( .A(n24736), .B(n24735), .Z(n42613) );
  NAND U44803 ( .A(n24738), .B(n24737), .Z(n42611) );
  NAND U44804 ( .A(n24740), .B(n24739), .Z(n42605) );
  NANDN U44805 ( .A(x[4878]), .B(y[4878]), .Z(n24742) );
  AND U44806 ( .A(n24742), .B(n24741), .Z(n42603) );
  NAND U44807 ( .A(n24744), .B(n24743), .Z(n42601) );
  NAND U44808 ( .A(n24746), .B(n24745), .Z(n42596) );
  NANDN U44809 ( .A(x[4874]), .B(y[4874]), .Z(n57176) );
  IV U44810 ( .A(n24747), .Z(n57178) );
  AND U44811 ( .A(n24749), .B(n24748), .Z(n42592) );
  NAND U44812 ( .A(n24751), .B(n24750), .Z(n42588) );
  NANDN U44813 ( .A(x[4870]), .B(y[4870]), .Z(n51538) );
  AND U44814 ( .A(n24753), .B(n24752), .Z(n42584) );
  IV U44815 ( .A(n24754), .Z(n57165) );
  ANDN U44816 ( .B(y[4866]), .A(x[4866]), .Z(n57163) );
  AND U44817 ( .A(n24756), .B(n24755), .Z(n42574) );
  NAND U44818 ( .A(n24758), .B(n24757), .Z(n42569) );
  NANDN U44819 ( .A(x[4862]), .B(y[4862]), .Z(n51541) );
  AND U44820 ( .A(n24760), .B(n24759), .Z(n42565) );
  NAND U44821 ( .A(n24762), .B(n24761), .Z(n42561) );
  AND U44822 ( .A(n24764), .B(n24763), .Z(n42556) );
  NAND U44823 ( .A(n24766), .B(n24765), .Z(n42552) );
  NANDN U44824 ( .A(x[4854]), .B(y[4854]), .Z(n51543) );
  AND U44825 ( .A(n24768), .B(n24767), .Z(n42548) );
  AND U44826 ( .A(n24769), .B(n51542), .Z(n42546) );
  NAND U44827 ( .A(n24771), .B(n24770), .Z(n42544) );
  NANDN U44828 ( .A(x[4850]), .B(y[4850]), .Z(n57142) );
  AND U44829 ( .A(n24773), .B(n24772), .Z(n42539) );
  AND U44830 ( .A(n24774), .B(n57143), .Z(n42537) );
  NAND U44831 ( .A(n24776), .B(n24775), .Z(n42535) );
  AND U44832 ( .A(n24778), .B(n24777), .Z(n42530) );
  NAND U44833 ( .A(n24780), .B(n24779), .Z(n42525) );
  AND U44834 ( .A(n24782), .B(n24781), .Z(n42521) );
  NANDN U44835 ( .A(x[4838]), .B(y[4838]), .Z(n24783) );
  AND U44836 ( .A(n24783), .B(n51544), .Z(n42513) );
  NAND U44837 ( .A(n24785), .B(n24784), .Z(n42511) );
  NAND U44838 ( .A(n24787), .B(n24786), .Z(n42506) );
  NANDN U44839 ( .A(x[4834]), .B(y[4834]), .Z(n24788) );
  AND U44840 ( .A(n24788), .B(n57123), .Z(n42504) );
  NAND U44841 ( .A(n24790), .B(n24789), .Z(n42502) );
  NAND U44842 ( .A(n24792), .B(n24791), .Z(n42496) );
  NANDN U44843 ( .A(x[4830]), .B(y[4830]), .Z(n24794) );
  AND U44844 ( .A(n24794), .B(n24793), .Z(n42494) );
  NAND U44845 ( .A(n24796), .B(n24795), .Z(n42492) );
  NAND U44846 ( .A(n24798), .B(n24797), .Z(n42487) );
  NANDN U44847 ( .A(x[4826]), .B(y[4826]), .Z(n24799) );
  AND U44848 ( .A(n24799), .B(n51546), .Z(n42485) );
  NAND U44849 ( .A(n24801), .B(n24800), .Z(n42483) );
  AND U44850 ( .A(n24803), .B(n24802), .Z(n42481) );
  NAND U44851 ( .A(n24805), .B(n24804), .Z(n42479) );
  NANDN U44852 ( .A(x[4822]), .B(y[4822]), .Z(n51549) );
  AND U44853 ( .A(n24807), .B(n24806), .Z(n42474) );
  AND U44854 ( .A(n24808), .B(n51548), .Z(n42472) );
  NANDN U44855 ( .A(x[4818]), .B(y[4818]), .Z(n24810) );
  AND U44856 ( .A(n24810), .B(n24809), .Z(n42466) );
  NAND U44857 ( .A(n24812), .B(n24811), .Z(n42464) );
  NANDN U44858 ( .A(x[4816]), .B(y[4816]), .Z(n24814) );
  AND U44859 ( .A(n24814), .B(n24813), .Z(n42462) );
  AND U44860 ( .A(n24816), .B(n24815), .Z(n42456) );
  NAND U44861 ( .A(n24818), .B(n24817), .Z(n42454) );
  AND U44862 ( .A(n24820), .B(n24819), .Z(n42452) );
  AND U44863 ( .A(n24822), .B(n24821), .Z(n42450) );
  NAND U44864 ( .A(n51555), .B(n24823), .Z(n42439) );
  NAND U44865 ( .A(n24827), .B(n24826), .Z(n57094) );
  IV U44866 ( .A(n24828), .Z(n57093) );
  AND U44867 ( .A(n24829), .B(n57093), .Z(n42435) );
  AND U44868 ( .A(n57092), .B(n24830), .Z(n42433) );
  AND U44869 ( .A(n24832), .B(n24831), .Z(n42431) );
  NAND U44870 ( .A(n24834), .B(n24833), .Z(n42429) );
  AND U44871 ( .A(n24836), .B(n24835), .Z(n42427) );
  AND U44872 ( .A(n24838), .B(n24837), .Z(n42421) );
  AND U44873 ( .A(n51557), .B(n24839), .Z(n42415) );
  AND U44874 ( .A(n24841), .B(n24840), .Z(n42410) );
  NANDN U44875 ( .A(x[4792]), .B(y[4792]), .Z(n24843) );
  AND U44876 ( .A(n24843), .B(n24842), .Z(n42405) );
  NANDN U44877 ( .A(x[4790]), .B(y[4790]), .Z(n24845) );
  AND U44878 ( .A(n24845), .B(n24844), .Z(n42399) );
  NANDN U44879 ( .A(x[4788]), .B(y[4788]), .Z(n24847) );
  AND U44880 ( .A(n24847), .B(n24846), .Z(n42393) );
  NANDN U44881 ( .A(x[4786]), .B(y[4786]), .Z(n24849) );
  AND U44882 ( .A(n24849), .B(n24848), .Z(n42387) );
  NANDN U44883 ( .A(x[4784]), .B(y[4784]), .Z(n24851) );
  AND U44884 ( .A(n24851), .B(n24850), .Z(n42381) );
  NANDN U44885 ( .A(x[4782]), .B(y[4782]), .Z(n24853) );
  AND U44886 ( .A(n24853), .B(n24852), .Z(n42375) );
  AND U44887 ( .A(n24855), .B(n24854), .Z(n42365) );
  NANDN U44888 ( .A(x[4778]), .B(y[4778]), .Z(n57064) );
  AND U44889 ( .A(n57064), .B(n24856), .Z(n42363) );
  NAND U44890 ( .A(n24858), .B(n24857), .Z(n42361) );
  NANDN U44891 ( .A(x[4776]), .B(y[4776]), .Z(n57061) );
  AND U44892 ( .A(n57063), .B(n57061), .Z(n42359) );
  NANDN U44893 ( .A(x[4774]), .B(y[4774]), .Z(n24859) );
  AND U44894 ( .A(n24859), .B(n57062), .Z(n42353) );
  NANDN U44895 ( .A(x[4772]), .B(y[4772]), .Z(n24861) );
  AND U44896 ( .A(n24861), .B(n24860), .Z(n42347) );
  AND U44897 ( .A(n24863), .B(n24862), .Z(n42345) );
  NANDN U44898 ( .A(x[4770]), .B(y[4770]), .Z(n57053) );
  AND U44899 ( .A(n24864), .B(n57053), .Z(n42343) );
  NAND U44900 ( .A(n24866), .B(n24865), .Z(n42341) );
  NANDN U44901 ( .A(x[4768]), .B(y[4768]), .Z(n24867) );
  AND U44902 ( .A(n24867), .B(n57055), .Z(n42339) );
  NANDN U44903 ( .A(x[4764]), .B(y[4764]), .Z(n24868) );
  AND U44904 ( .A(n24868), .B(n57048), .Z(n42326) );
  ANDN U44905 ( .B(y[4762]), .A(x[4762]), .Z(n24870) );
  NOR U44906 ( .A(n24870), .B(n24869), .Z(n42320) );
  NANDN U44907 ( .A(x[4760]), .B(y[4760]), .Z(n24872) );
  AND U44908 ( .A(n24872), .B(n24871), .Z(n42314) );
  NANDN U44909 ( .A(x[4758]), .B(y[4758]), .Z(n24874) );
  AND U44910 ( .A(n24874), .B(n24873), .Z(n42308) );
  NANDN U44911 ( .A(x[4756]), .B(y[4756]), .Z(n24876) );
  AND U44912 ( .A(n24876), .B(n24875), .Z(n42302) );
  NANDN U44913 ( .A(x[4754]), .B(y[4754]), .Z(n24878) );
  AND U44914 ( .A(n24878), .B(n24877), .Z(n42296) );
  NANDN U44915 ( .A(x[4752]), .B(y[4752]), .Z(n24880) );
  AND U44916 ( .A(n24880), .B(n24879), .Z(n42290) );
  NANDN U44917 ( .A(x[4750]), .B(y[4750]), .Z(n24882) );
  AND U44918 ( .A(n24882), .B(n24881), .Z(n42284) );
  NAND U44919 ( .A(n24884), .B(n24883), .Z(n42282) );
  NAND U44920 ( .A(n24886), .B(n24885), .Z(n42277) );
  NAND U44921 ( .A(n24888), .B(n24887), .Z(n42272) );
  AND U44922 ( .A(n24890), .B(n24889), .Z(n42252) );
  NAND U44923 ( .A(n24892), .B(n24891), .Z(n42223) );
  NANDN U44924 ( .A(x[4730]), .B(y[4730]), .Z(n57013) );
  AND U44925 ( .A(n57013), .B(n57015), .Z(n42221) );
  IV U44926 ( .A(n24893), .Z(n57014) );
  NANDN U44927 ( .A(x[4728]), .B(y[4728]), .Z(n51572) );
  AND U44928 ( .A(n24895), .B(n24894), .Z(n42213) );
  NANDN U44929 ( .A(x[4726]), .B(y[4726]), .Z(n57008) );
  IV U44930 ( .A(n24896), .Z(n51571) );
  AND U44931 ( .A(n57008), .B(n51571), .Z(n42211) );
  NAND U44932 ( .A(n24898), .B(n24897), .Z(n42209) );
  NANDN U44933 ( .A(x[4724]), .B(y[4724]), .Z(n57006) );
  IV U44934 ( .A(n24899), .Z(n57007) );
  AND U44935 ( .A(n57006), .B(n57007), .Z(n42207) );
  NAND U44936 ( .A(n24901), .B(n24900), .Z(n42205) );
  NAND U44937 ( .A(n24903), .B(n24902), .Z(n42200) );
  NAND U44938 ( .A(n24905), .B(n24904), .Z(n42194) );
  AND U44939 ( .A(n24907), .B(n24906), .Z(n42192) );
  NAND U44940 ( .A(n24909), .B(n24908), .Z(n42190) );
  NAND U44941 ( .A(n24911), .B(n24910), .Z(n42176) );
  NANDN U44942 ( .A(x[4712]), .B(y[4712]), .Z(n24913) );
  AND U44943 ( .A(n24913), .B(n24912), .Z(n42174) );
  NANDN U44944 ( .A(x[4710]), .B(y[4710]), .Z(n56990) );
  NAND U44945 ( .A(n56990), .B(n24914), .Z(n42168) );
  ANDN U44946 ( .B(y[4708]), .A(x[4708]), .Z(n56987) );
  AND U44947 ( .A(n24916), .B(n24915), .Z(n42160) );
  AND U44948 ( .A(n56988), .B(n24917), .Z(n42158) );
  NAND U44949 ( .A(n24919), .B(n24918), .Z(n42156) );
  NANDN U44950 ( .A(x[4704]), .B(y[4704]), .Z(n24921) );
  AND U44951 ( .A(n24921), .B(n24920), .Z(n42154) );
  NANDN U44952 ( .A(x[4702]), .B(y[4702]), .Z(n24923) );
  AND U44953 ( .A(n24923), .B(n24922), .Z(n42148) );
  NANDN U44954 ( .A(x[4700]), .B(y[4700]), .Z(n24925) );
  AND U44955 ( .A(n24925), .B(n24924), .Z(n42142) );
  AND U44956 ( .A(n24927), .B(n24926), .Z(n42132) );
  NANDN U44957 ( .A(x[4696]), .B(y[4696]), .Z(n56973) );
  NAND U44958 ( .A(n56973), .B(n24928), .Z(n42130) );
  AND U44959 ( .A(n24930), .B(n24929), .Z(n42128) );
  AND U44960 ( .A(n24932), .B(n24931), .Z(n42123) );
  AND U44961 ( .A(n24934), .B(n24933), .Z(n42118) );
  ANDN U44962 ( .B(y[4690]), .A(x[4690]), .Z(n56964) );
  AND U44963 ( .A(n24936), .B(n24935), .Z(n42107) );
  ANDN U44964 ( .B(y[4686]), .A(x[4686]), .Z(n42105) );
  NAND U44965 ( .A(n24938), .B(n24937), .Z(n42101) );
  NANDN U44966 ( .A(x[4684]), .B(y[4684]), .Z(n24940) );
  AND U44967 ( .A(n24940), .B(n24939), .Z(n42099) );
  NANDN U44968 ( .A(x[4682]), .B(y[4682]), .Z(n51578) );
  NAND U44969 ( .A(n51578), .B(n24941), .Z(n42093) );
  AND U44970 ( .A(n24943), .B(n24942), .Z(n42085) );
  ANDN U44971 ( .B(y[4678]), .A(x[4678]), .Z(n24944) );
  NOR U44972 ( .A(n56953), .B(n24944), .Z(n42083) );
  NANDN U44973 ( .A(x[4676]), .B(y[4676]), .Z(n51580) );
  AND U44974 ( .A(n51580), .B(n24945), .Z(n42077) );
  NANDN U44975 ( .A(x[4674]), .B(y[4674]), .Z(n24946) );
  AND U44976 ( .A(n24946), .B(n51579), .Z(n42071) );
  NANDN U44977 ( .A(x[4672]), .B(y[4672]), .Z(n24948) );
  AND U44978 ( .A(n24948), .B(n24947), .Z(n42065) );
  NANDN U44979 ( .A(x[4670]), .B(y[4670]), .Z(n24950) );
  AND U44980 ( .A(n24950), .B(n24949), .Z(n42059) );
  NANDN U44981 ( .A(x[4668]), .B(y[4668]), .Z(n24952) );
  AND U44982 ( .A(n24952), .B(n24951), .Z(n42053) );
  AND U44983 ( .A(n24954), .B(n24953), .Z(n42043) );
  AND U44984 ( .A(n24956), .B(n24955), .Z(n42037) );
  AND U44985 ( .A(n24958), .B(n24957), .Z(n42032) );
  AND U44986 ( .A(n24960), .B(n24959), .Z(n42027) );
  ANDN U44987 ( .B(y[4658]), .A(x[4658]), .Z(n42025) );
  NAND U44988 ( .A(n24962), .B(n24961), .Z(n41998) );
  NANDN U44989 ( .A(x[4650]), .B(y[4650]), .Z(n24963) );
  AND U44990 ( .A(n24963), .B(n56924), .Z(n41996) );
  NANDN U44991 ( .A(x[4646]), .B(y[4646]), .Z(n51585) );
  AND U44992 ( .A(n51585), .B(n56918), .Z(n41987) );
  NAND U44993 ( .A(n24967), .B(n24966), .Z(n41985) );
  NANDN U44994 ( .A(x[4644]), .B(y[4644]), .Z(n56915) );
  AND U44995 ( .A(n56915), .B(n51584), .Z(n41983) );
  ANDN U44996 ( .B(y[4642]), .A(x[4642]), .Z(n24968) );
  NOR U44997 ( .A(n56914), .B(n24968), .Z(n41977) );
  NANDN U44998 ( .A(x[4640]), .B(y[4640]), .Z(n24970) );
  AND U44999 ( .A(n24970), .B(n24969), .Z(n41971) );
  NAND U45000 ( .A(n51587), .B(n24971), .Z(n41969) );
  AND U45001 ( .A(n56906), .B(n24972), .Z(n41961) );
  NAND U45002 ( .A(n56905), .B(n24973), .Z(n41959) );
  AND U45003 ( .A(n24975), .B(n24974), .Z(n41913) );
  ANDN U45004 ( .B(y[4622]), .A(x[4622]), .Z(n41911) );
  NAND U45005 ( .A(n24977), .B(n24976), .Z(n41894) );
  NANDN U45006 ( .A(x[4616]), .B(y[4616]), .Z(n24978) );
  AND U45007 ( .A(n24978), .B(n51592), .Z(n41892) );
  NAND U45008 ( .A(n24980), .B(n24979), .Z(n41886) );
  ANDN U45009 ( .B(y[4612]), .A(x[4612]), .Z(n51595) );
  AND U45010 ( .A(n24982), .B(n24981), .Z(n41877) );
  NANDN U45011 ( .A(x[4610]), .B(y[4610]), .Z(n24983) );
  AND U45012 ( .A(n24983), .B(n51594), .Z(n41875) );
  NAND U45013 ( .A(n24985), .B(n24984), .Z(n41873) );
  NANDN U45014 ( .A(x[4608]), .B(y[4608]), .Z(n56876) );
  AND U45015 ( .A(n56876), .B(n24986), .Z(n41871) );
  NANDN U45016 ( .A(x[4606]), .B(y[4606]), .Z(n24987) );
  AND U45017 ( .A(n24987), .B(n56877), .Z(n41865) );
  NANDN U45018 ( .A(x[4604]), .B(y[4604]), .Z(n24989) );
  AND U45019 ( .A(n24989), .B(n24988), .Z(n41859) );
  NANDN U45020 ( .A(x[4602]), .B(y[4602]), .Z(n24991) );
  AND U45021 ( .A(n24991), .B(n24990), .Z(n41853) );
  NAND U45022 ( .A(n24993), .B(n24992), .Z(n41843) );
  AND U45023 ( .A(n24995), .B(n24994), .Z(n41837) );
  NANDN U45024 ( .A(x[4596]), .B(y[4596]), .Z(n24997) );
  AND U45025 ( .A(n24997), .B(n24996), .Z(n41835) );
  NAND U45026 ( .A(n24999), .B(n24998), .Z(n41833) );
  NANDN U45027 ( .A(x[4594]), .B(y[4594]), .Z(n25001) );
  AND U45028 ( .A(n25001), .B(n25000), .Z(n41831) );
  NANDN U45029 ( .A(x[4592]), .B(y[4592]), .Z(n25003) );
  AND U45030 ( .A(n25003), .B(n25002), .Z(n41825) );
  AND U45031 ( .A(n25005), .B(n25004), .Z(n41815) );
  AND U45032 ( .A(n25007), .B(n25006), .Z(n41810) );
  XNOR U45033 ( .A(x[4586]), .B(y[4586]), .Z(n25009) );
  AND U45034 ( .A(n25009), .B(n25008), .Z(n41806) );
  ANDN U45035 ( .B(y[4584]), .A(x[4584]), .Z(n41804) );
  NAND U45036 ( .A(n56838), .B(n25010), .Z(n41758) );
  NANDN U45037 ( .A(x[4570]), .B(y[4570]), .Z(n56834) );
  NAND U45038 ( .A(n56834), .B(n25011), .Z(n41752) );
  AND U45039 ( .A(n25013), .B(n25012), .Z(n41744) );
  NANDN U45040 ( .A(x[4566]), .B(y[4566]), .Z(n56827) );
  NAND U45041 ( .A(n56827), .B(n56830), .Z(n41742) );
  AND U45042 ( .A(n25015), .B(n25014), .Z(n41740) );
  NANDN U45043 ( .A(x[4564]), .B(y[4564]), .Z(n51602) );
  AND U45044 ( .A(n25017), .B(n25016), .Z(n41736) );
  AND U45045 ( .A(n25019), .B(n25018), .Z(n41731) );
  NANDN U45046 ( .A(x[4558]), .B(y[4558]), .Z(n25021) );
  NAND U45047 ( .A(n25021), .B(n25020), .Z(n41721) );
  AND U45048 ( .A(n25023), .B(n25022), .Z(n41719) );
  NANDN U45049 ( .A(x[4556]), .B(y[4556]), .Z(n25025) );
  NAND U45050 ( .A(n25025), .B(n25024), .Z(n41717) );
  NANDN U45051 ( .A(x[4552]), .B(y[4552]), .Z(n51604) );
  NAND U45052 ( .A(n51604), .B(n25026), .Z(n41703) );
  ANDN U45053 ( .B(y[4550]), .A(x[4550]), .Z(n56812) );
  AND U45054 ( .A(n25028), .B(n25027), .Z(n41695) );
  NANDN U45055 ( .A(x[4548]), .B(y[4548]), .Z(n56809) );
  AND U45056 ( .A(n56809), .B(n56811), .Z(n41693) );
  NAND U45057 ( .A(n25030), .B(n25029), .Z(n41691) );
  NANDN U45058 ( .A(x[4546]), .B(y[4546]), .Z(n25031) );
  AND U45059 ( .A(n25031), .B(n56808), .Z(n41689) );
  NANDN U45060 ( .A(x[4544]), .B(y[4544]), .Z(n25033) );
  AND U45061 ( .A(n25033), .B(n25032), .Z(n41683) );
  AND U45062 ( .A(n25035), .B(n25034), .Z(n41677) );
  NANDN U45063 ( .A(x[4540]), .B(y[4540]), .Z(n25037) );
  AND U45064 ( .A(n25037), .B(n25036), .Z(n41671) );
  NANDN U45065 ( .A(x[4538]), .B(y[4538]), .Z(n56789) );
  AND U45066 ( .A(n56789), .B(n25038), .Z(n41665) );
  NAND U45067 ( .A(n25040), .B(n25039), .Z(n41663) );
  NAND U45068 ( .A(n25042), .B(n25041), .Z(n41658) );
  NAND U45069 ( .A(n25044), .B(n25043), .Z(n41652) );
  IV U45070 ( .A(n25045), .Z(n56767) );
  NANDN U45071 ( .A(x[4528]), .B(y[4528]), .Z(n25046) );
  NAND U45072 ( .A(n56767), .B(n25046), .Z(n41637) );
  NANDN U45073 ( .A(x[4526]), .B(y[4526]), .Z(n25048) );
  NAND U45074 ( .A(n25048), .B(n25047), .Z(n41631) );
  AND U45075 ( .A(n25050), .B(n25049), .Z(n41617) );
  NANDN U45076 ( .A(x[4520]), .B(y[4520]), .Z(n25052) );
  AND U45077 ( .A(n25052), .B(n25051), .Z(n41611) );
  AND U45078 ( .A(n25054), .B(n25053), .Z(n41602) );
  NANDN U45079 ( .A(x[4516]), .B(y[4516]), .Z(n25055) );
  AND U45080 ( .A(n25055), .B(n56755), .Z(n41600) );
  NAND U45081 ( .A(n25057), .B(n25056), .Z(n41598) );
  NANDN U45082 ( .A(x[4514]), .B(y[4514]), .Z(n25059) );
  AND U45083 ( .A(n25059), .B(n25058), .Z(n41596) );
  NANDN U45084 ( .A(x[4512]), .B(y[4512]), .Z(n25061) );
  AND U45085 ( .A(n25061), .B(n25060), .Z(n41590) );
  NAND U45086 ( .A(n25063), .B(n25062), .Z(n41580) );
  NAND U45087 ( .A(n25065), .B(n25064), .Z(n41574) );
  NAND U45088 ( .A(n25067), .B(n25066), .Z(n41568) );
  AND U45089 ( .A(n25069), .B(n25068), .Z(n41566) );
  NAND U45090 ( .A(n25071), .B(n25070), .Z(n41564) );
  AND U45091 ( .A(n25073), .B(n25072), .Z(n41530) );
  AND U45092 ( .A(n25075), .B(n25074), .Z(n41528) );
  NAND U45093 ( .A(n25077), .B(n25076), .Z(n41526) );
  AND U45094 ( .A(n56731), .B(n25078), .Z(n41524) );
  NAND U45095 ( .A(n25080), .B(n25079), .Z(n56730) );
  AND U45096 ( .A(n25083), .B(n56728), .Z(n41520) );
  NAND U45097 ( .A(n56727), .B(n25084), .Z(n41518) );
  NANDN U45098 ( .A(x[4486]), .B(y[4486]), .Z(n56722) );
  AND U45099 ( .A(n25086), .B(n25085), .Z(n41513) );
  AND U45100 ( .A(n25088), .B(n25087), .Z(n41508) );
  AND U45101 ( .A(n25090), .B(n25089), .Z(n41502) );
  AND U45102 ( .A(n25092), .B(n25091), .Z(n41500) );
  NAND U45103 ( .A(n25094), .B(n25093), .Z(n41498) );
  NANDN U45104 ( .A(x[4476]), .B(y[4476]), .Z(n25095) );
  NAND U45105 ( .A(n25095), .B(n51612), .Z(n41489) );
  NANDN U45106 ( .A(x[4474]), .B(y[4474]), .Z(n25097) );
  NAND U45107 ( .A(n25097), .B(n25096), .Z(n41483) );
  ANDN U45108 ( .B(y[4472]), .A(x[4472]), .Z(n41477) );
  NANDN U45109 ( .A(x[4470]), .B(y[4470]), .Z(n25099) );
  AND U45110 ( .A(n25099), .B(n25098), .Z(n41469) );
  NANDN U45111 ( .A(x[4468]), .B(y[4468]), .Z(n25101) );
  AND U45112 ( .A(n25101), .B(n25100), .Z(n41463) );
  NANDN U45113 ( .A(x[4466]), .B(y[4466]), .Z(n25103) );
  AND U45114 ( .A(n25103), .B(n25102), .Z(n41457) );
  NAND U45115 ( .A(n25105), .B(n25104), .Z(n41455) );
  ANDN U45116 ( .B(y[4464]), .A(x[4464]), .Z(n41451) );
  AND U45117 ( .A(n25107), .B(n25106), .Z(n41449) );
  NANDN U45118 ( .A(x[4460]), .B(y[4460]), .Z(n51619) );
  NAND U45119 ( .A(n56699), .B(n51619), .Z(n41440) );
  AND U45120 ( .A(n25109), .B(n25108), .Z(n41438) );
  NANDN U45121 ( .A(x[4458]), .B(y[4458]), .Z(n25110) );
  NAND U45122 ( .A(n51617), .B(n25110), .Z(n41436) );
  AND U45123 ( .A(n25112), .B(n25111), .Z(n41434) );
  ANDN U45124 ( .B(y[4456]), .A(x[4456]), .Z(n41432) );
  AND U45125 ( .A(n25114), .B(n25113), .Z(n41424) );
  NAND U45126 ( .A(n25116), .B(n25115), .Z(n41422) );
  AND U45127 ( .A(n25118), .B(n25117), .Z(n41409) );
  ANDN U45128 ( .B(y[4448]), .A(x[4448]), .Z(n41407) );
  AND U45129 ( .A(n25120), .B(n25119), .Z(n41396) );
  ANDN U45130 ( .B(y[4444]), .A(x[4444]), .Z(n41394) );
  NAND U45131 ( .A(n25122), .B(n25121), .Z(n41346) );
  NANDN U45132 ( .A(x[4430]), .B(y[4430]), .Z(n56669) );
  NAND U45133 ( .A(n56669), .B(n25123), .Z(n41340) );
  ANDN U45134 ( .B(y[4428]), .A(x[4428]), .Z(n56666) );
  AND U45135 ( .A(n25125), .B(n25124), .Z(n41332) );
  NANDN U45136 ( .A(x[4426]), .B(y[4426]), .Z(n25127) );
  IV U45137 ( .A(n25126), .Z(n56665) );
  AND U45138 ( .A(n25127), .B(n56665), .Z(n41330) );
  NAND U45139 ( .A(n25129), .B(n25128), .Z(n41328) );
  NANDN U45140 ( .A(x[4424]), .B(y[4424]), .Z(n25131) );
  AND U45141 ( .A(n25131), .B(n25130), .Z(n41326) );
  NAND U45142 ( .A(n25133), .B(n25132), .Z(n41324) );
  NAND U45143 ( .A(n25135), .B(n25134), .Z(n41318) );
  NAND U45144 ( .A(n25137), .B(n25136), .Z(n41312) );
  NAND U45145 ( .A(n25139), .B(n25138), .Z(n41306) );
  AND U45146 ( .A(n25141), .B(n25140), .Z(n41304) );
  NAND U45147 ( .A(n25143), .B(n25142), .Z(n41302) );
  XNOR U45148 ( .A(x[4412]), .B(y[4412]), .Z(n41289) );
  IV U45149 ( .A(n25144), .Z(n56652) );
  NAND U45150 ( .A(n56652), .B(n25145), .Z(n41287) );
  NANDN U45151 ( .A(x[4408]), .B(y[4408]), .Z(n51635) );
  NAND U45152 ( .A(n51635), .B(n25146), .Z(n41281) );
  ANDN U45153 ( .B(y[4406]), .A(x[4406]), .Z(n56647) );
  AND U45154 ( .A(n25148), .B(n25147), .Z(n41273) );
  NANDN U45155 ( .A(x[4404]), .B(y[4404]), .Z(n25150) );
  IV U45156 ( .A(n25149), .Z(n56646) );
  AND U45157 ( .A(n25150), .B(n56646), .Z(n41271) );
  NAND U45158 ( .A(n25152), .B(n25151), .Z(n41269) );
  NANDN U45159 ( .A(x[4402]), .B(y[4402]), .Z(n25154) );
  AND U45160 ( .A(n25154), .B(n25153), .Z(n41267) );
  NANDN U45161 ( .A(x[4400]), .B(y[4400]), .Z(n25156) );
  AND U45162 ( .A(n25156), .B(n25155), .Z(n41261) );
  ANDN U45163 ( .B(y[4398]), .A(x[4398]), .Z(n41255) );
  AND U45164 ( .A(n25158), .B(n25157), .Z(n41251) );
  AND U45165 ( .A(n25160), .B(n25159), .Z(n41245) );
  NAND U45166 ( .A(n25162), .B(n25161), .Z(n41240) );
  AND U45167 ( .A(n25164), .B(n25163), .Z(n41235) );
  NANDN U45168 ( .A(x[4388]), .B(y[4388]), .Z(n25166) );
  NAND U45169 ( .A(n25166), .B(n25165), .Z(n41225) );
  NANDN U45170 ( .A(x[4386]), .B(y[4386]), .Z(n25168) );
  NAND U45171 ( .A(n25168), .B(n25167), .Z(n41219) );
  ANDN U45172 ( .B(y[4384]), .A(x[4384]), .Z(n41211) );
  AND U45173 ( .A(n25170), .B(n25169), .Z(n41209) );
  ANDN U45174 ( .B(y[4382]), .A(x[4382]), .Z(n41207) );
  NAND U45175 ( .A(n25172), .B(n25171), .Z(n41195) );
  NAND U45176 ( .A(n25174), .B(n25173), .Z(n41189) );
  AND U45177 ( .A(n25176), .B(n25175), .Z(n41187) );
  NAND U45178 ( .A(n25178), .B(n25177), .Z(n41185) );
  AND U45179 ( .A(n25179), .B(n51643), .Z(n41176) );
  NAND U45180 ( .A(n25181), .B(n25180), .Z(n41174) );
  AND U45181 ( .A(n25183), .B(n25182), .Z(n41172) );
  NANDN U45182 ( .A(x[4368]), .B(y[4368]), .Z(n25185) );
  AND U45183 ( .A(n25185), .B(n25184), .Z(n41166) );
  ANDN U45184 ( .B(y[4366]), .A(x[4366]), .Z(n51646) );
  AND U45185 ( .A(n25187), .B(n25186), .Z(n41157) );
  NANDN U45186 ( .A(x[4364]), .B(y[4364]), .Z(n56608) );
  IV U45187 ( .A(n25188), .Z(n56609) );
  AND U45188 ( .A(n56608), .B(n56609), .Z(n41155) );
  NAND U45189 ( .A(n25190), .B(n25189), .Z(n41153) );
  NANDN U45190 ( .A(x[4362]), .B(y[4362]), .Z(n25191) );
  AND U45191 ( .A(n25191), .B(n56606), .Z(n41151) );
  NANDN U45192 ( .A(x[4360]), .B(y[4360]), .Z(n56601) );
  AND U45193 ( .A(n56601), .B(n25192), .Z(n41145) );
  NAND U45194 ( .A(n25194), .B(n25193), .Z(n41143) );
  NAND U45195 ( .A(n25196), .B(n25195), .Z(n41138) );
  AND U45196 ( .A(n25198), .B(n25197), .Z(n41128) );
  NAND U45197 ( .A(n25200), .B(n25199), .Z(n41116) );
  AND U45198 ( .A(n25202), .B(n25201), .Z(n41114) );
  AND U45199 ( .A(n25204), .B(n25203), .Z(n41108) );
  AND U45200 ( .A(n25206), .B(n25205), .Z(n41102) );
  AND U45201 ( .A(n25208), .B(n25207), .Z(n41096) );
  NANDN U45202 ( .A(x[4340]), .B(y[4340]), .Z(n25210) );
  AND U45203 ( .A(n25210), .B(n25209), .Z(n41090) );
  AND U45204 ( .A(n25212), .B(n25211), .Z(n41084) );
  NANDN U45205 ( .A(x[4336]), .B(y[4336]), .Z(n56579) );
  AND U45206 ( .A(n25213), .B(n56579), .Z(n41078) );
  NAND U45207 ( .A(n25215), .B(n25214), .Z(n41069) );
  NAND U45208 ( .A(n25217), .B(n25216), .Z(n41063) );
  NAND U45209 ( .A(n25219), .B(n25218), .Z(n41057) );
  AND U45210 ( .A(n25221), .B(n25220), .Z(n41055) );
  NAND U45211 ( .A(n25223), .B(n25222), .Z(n41053) );
  AND U45212 ( .A(n25225), .B(n25224), .Z(n41025) );
  ANDN U45213 ( .B(y[4316]), .A(x[4316]), .Z(n41013) );
  AND U45214 ( .A(n25227), .B(n25226), .Z(n41011) );
  AND U45215 ( .A(n25229), .B(n25228), .Z(n41005) );
  AND U45216 ( .A(n25231), .B(n25230), .Z(n40999) );
  AND U45217 ( .A(n25233), .B(n25232), .Z(n40993) );
  AND U45218 ( .A(n25235), .B(n25234), .Z(n40983) );
  NAND U45219 ( .A(n25237), .B(n25236), .Z(n40981) );
  NAND U45220 ( .A(n25239), .B(n25238), .Z(n40970) );
  NANDN U45221 ( .A(x[4300]), .B(y[4300]), .Z(n25240) );
  AND U45222 ( .A(n25240), .B(n56545), .Z(n40968) );
  NANDN U45223 ( .A(x[4298]), .B(y[4298]), .Z(n25242) );
  AND U45224 ( .A(n25242), .B(n25241), .Z(n40962) );
  AND U45225 ( .A(n25244), .B(n25243), .Z(n40956) );
  AND U45226 ( .A(n25246), .B(n25245), .Z(n40954) );
  ANDN U45227 ( .B(y[4294]), .A(x[4294]), .Z(n25248) );
  NOR U45228 ( .A(n25248), .B(n25247), .Z(n40952) );
  AND U45229 ( .A(n25250), .B(n25249), .Z(n40946) );
  AND U45230 ( .A(n25252), .B(n25251), .Z(n40936) );
  AND U45231 ( .A(n25254), .B(n25253), .Z(n40930) );
  NAND U45232 ( .A(n25256), .B(n25255), .Z(n40924) );
  NAND U45233 ( .A(n25258), .B(n25257), .Z(n40918) );
  NANDN U45234 ( .A(x[4282]), .B(y[4282]), .Z(n25260) );
  AND U45235 ( .A(n25260), .B(n25259), .Z(n40916) );
  NAND U45236 ( .A(n25262), .B(n25261), .Z(n40914) );
  NANDN U45237 ( .A(x[4278]), .B(y[4278]), .Z(n25264) );
  AND U45238 ( .A(n25264), .B(n25263), .Z(n40904) );
  NAND U45239 ( .A(n25266), .B(n25265), .Z(n40898) );
  NANDN U45240 ( .A(x[4274]), .B(y[4274]), .Z(n56518) );
  NAND U45241 ( .A(n56518), .B(n25267), .Z(n40892) );
  IV U45242 ( .A(n25268), .Z(n56517) );
  NAND U45243 ( .A(n56517), .B(n25269), .Z(n40886) );
  AND U45244 ( .A(n25271), .B(n25270), .Z(n40884) );
  NANDN U45245 ( .A(x[4270]), .B(y[4270]), .Z(n51669) );
  NAND U45246 ( .A(n51669), .B(n25272), .Z(n40882) );
  AND U45247 ( .A(n25274), .B(n25273), .Z(n40880) );
  IV U45248 ( .A(n25275), .Z(n51668) );
  NAND U45249 ( .A(n51668), .B(n25276), .Z(n40878) );
  AND U45250 ( .A(n25278), .B(n25277), .Z(n40876) );
  NAND U45251 ( .A(n25280), .B(n25279), .Z(n40870) );
  AND U45252 ( .A(n25282), .B(n25281), .Z(n40864) );
  NANDN U45253 ( .A(x[4262]), .B(y[4262]), .Z(n25284) );
  NAND U45254 ( .A(n25284), .B(n25283), .Z(n40862) );
  AND U45255 ( .A(n25286), .B(n25285), .Z(n40860) );
  AND U45256 ( .A(n25288), .B(n25287), .Z(n40840) );
  AND U45257 ( .A(n25290), .B(n25289), .Z(n40834) );
  AND U45258 ( .A(n25292), .B(n25291), .Z(n40824) );
  NAND U45259 ( .A(n25294), .B(n25293), .Z(n40822) );
  AND U45260 ( .A(n25296), .B(n25295), .Z(n40806) );
  AND U45261 ( .A(n25298), .B(n25297), .Z(n40804) );
  NAND U45262 ( .A(n25300), .B(n25299), .Z(n40802) );
  NAND U45263 ( .A(n25302), .B(n25301), .Z(n40792) );
  NANDN U45264 ( .A(x[4238]), .B(y[4238]), .Z(n25304) );
  AND U45265 ( .A(n25304), .B(n25303), .Z(n40790) );
  NANDN U45266 ( .A(x[4236]), .B(y[4236]), .Z(n51677) );
  NAND U45267 ( .A(n51677), .B(n25305), .Z(n40784) );
  NAND U45268 ( .A(n25306), .B(n51676), .Z(n40778) );
  AND U45269 ( .A(n25308), .B(n25307), .Z(n40776) );
  NANDN U45270 ( .A(x[4232]), .B(y[4232]), .Z(n56467) );
  AND U45271 ( .A(n56467), .B(n25309), .Z(n40774) );
  NAND U45272 ( .A(n25311), .B(n25310), .Z(n40772) );
  NANDN U45273 ( .A(x[4230]), .B(y[4230]), .Z(n25312) );
  AND U45274 ( .A(n25312), .B(n56470), .Z(n40770) );
  NAND U45275 ( .A(n25314), .B(n25313), .Z(n40760) );
  NAND U45276 ( .A(n25316), .B(n25315), .Z(n40754) );
  NAND U45277 ( .A(n25318), .B(n25317), .Z(n40748) );
  AND U45278 ( .A(n25320), .B(n25319), .Z(n40746) );
  NAND U45279 ( .A(n25322), .B(n25321), .Z(n40732) );
  NAND U45280 ( .A(n25324), .B(n25323), .Z(n40726) );
  ANDN U45281 ( .B(y[4214]), .A(x[4214]), .Z(n51678) );
  AND U45282 ( .A(n25326), .B(n25325), .Z(n40717) );
  AND U45283 ( .A(n51679), .B(n25327), .Z(n40715) );
  NAND U45284 ( .A(n25329), .B(n25328), .Z(n40713) );
  AND U45285 ( .A(n25331), .B(n25330), .Z(n40711) );
  AND U45286 ( .A(n25333), .B(n25332), .Z(n40705) );
  AND U45287 ( .A(n25335), .B(n25334), .Z(n40699) );
  NANDN U45288 ( .A(x[4204]), .B(y[4204]), .Z(n56428) );
  AND U45289 ( .A(n25336), .B(n56428), .Z(n40693) );
  NANDN U45290 ( .A(x[4202]), .B(y[4202]), .Z(n51681) );
  AND U45291 ( .A(n51681), .B(n56427), .Z(n40687) );
  IV U45292 ( .A(n25337), .Z(n51680) );
  AND U45293 ( .A(n25339), .B(n25338), .Z(n40678) );
  ANDN U45294 ( .B(y[4198]), .A(x[4198]), .Z(n40676) );
  NAND U45295 ( .A(n25341), .B(n25340), .Z(n40672) );
  AND U45296 ( .A(n25343), .B(n25342), .Z(n40666) );
  NAND U45297 ( .A(n25345), .B(n25344), .Z(n40652) );
  AND U45298 ( .A(n25347), .B(n25346), .Z(n40638) );
  AND U45299 ( .A(n25349), .B(n25348), .Z(n40632) );
  AND U45300 ( .A(n25351), .B(n25350), .Z(n40626) );
  AND U45301 ( .A(n25353), .B(n25352), .Z(n40620) );
  NAND U45302 ( .A(n25355), .B(n25354), .Z(n40610) );
  NAND U45303 ( .A(n25357), .B(n25356), .Z(n40604) );
  AND U45304 ( .A(n25359), .B(n25358), .Z(n40590) );
  AND U45305 ( .A(n25361), .B(n25360), .Z(n40584) );
  AND U45306 ( .A(n25363), .B(n25362), .Z(n40578) );
  AND U45307 ( .A(n25365), .B(n25364), .Z(n40568) );
  AND U45308 ( .A(n25367), .B(n25366), .Z(n40566) );
  NAND U45309 ( .A(n25369), .B(n25368), .Z(n40564) );
  AND U45310 ( .A(n25371), .B(n25370), .Z(n40562) );
  NANDN U45311 ( .A(x[4160]), .B(y[4160]), .Z(n25373) );
  AND U45312 ( .A(n25373), .B(n25372), .Z(n40556) );
  NANDN U45313 ( .A(x[4158]), .B(y[4158]), .Z(n25375) );
  AND U45314 ( .A(n25375), .B(n25374), .Z(n40550) );
  NANDN U45315 ( .A(x[4156]), .B(y[4156]), .Z(n25377) );
  AND U45316 ( .A(n25377), .B(n25376), .Z(n40544) );
  NANDN U45317 ( .A(x[4154]), .B(y[4154]), .Z(n51693) );
  AND U45318 ( .A(n51693), .B(n25378), .Z(n40538) );
  NANDN U45319 ( .A(x[4152]), .B(y[4152]), .Z(n56381) );
  AND U45320 ( .A(n56381), .B(n51692), .Z(n40532) );
  NAND U45321 ( .A(n25380), .B(n25379), .Z(n40530) );
  NAND U45322 ( .A(n25382), .B(n25381), .Z(n40524) );
  NAND U45323 ( .A(n25384), .B(n25383), .Z(n40519) );
  AND U45324 ( .A(n25386), .B(n25385), .Z(n40514) );
  AND U45325 ( .A(n25388), .B(n25387), .Z(n40508) );
  NAND U45326 ( .A(n25390), .B(n25389), .Z(n40498) );
  NAND U45327 ( .A(n25392), .B(n25391), .Z(n40492) );
  NAND U45328 ( .A(n25394), .B(n25393), .Z(n40486) );
  AND U45329 ( .A(n25396), .B(n25395), .Z(n40484) );
  ANDN U45330 ( .B(y[4134]), .A(x[4134]), .Z(n56365) );
  NOR U45331 ( .A(n56365), .B(n25397), .Z(n40482) );
  AND U45332 ( .A(n25398), .B(n56364), .Z(n40476) );
  NANDN U45333 ( .A(x[4128]), .B(y[4128]), .Z(n56359) );
  AND U45334 ( .A(n56359), .B(n25399), .Z(n40462) );
  AND U45335 ( .A(n25400), .B(n56358), .Z(n40456) );
  AND U45336 ( .A(n25402), .B(n25401), .Z(n40454) );
  NAND U45337 ( .A(n25404), .B(n25403), .Z(n40448) );
  NAND U45338 ( .A(n25406), .B(n25405), .Z(n40442) );
  NAND U45339 ( .A(n25408), .B(n25407), .Z(n40436) );
  AND U45340 ( .A(n25410), .B(n25409), .Z(n40422) );
  AND U45341 ( .A(n25412), .B(n25411), .Z(n40416) );
  AND U45342 ( .A(n25414), .B(n25413), .Z(n40410) );
  AND U45343 ( .A(n25416), .B(n25415), .Z(n40404) );
  AND U45344 ( .A(n25418), .B(n25417), .Z(n40398) );
  AND U45345 ( .A(n25420), .B(n25419), .Z(n40392) );
  AND U45346 ( .A(n25422), .B(n25421), .Z(n40386) );
  AND U45347 ( .A(n25424), .B(n25423), .Z(n40380) );
  NAND U45348 ( .A(n25426), .B(n25425), .Z(n40370) );
  NANDN U45349 ( .A(x[4096]), .B(y[4096]), .Z(n56330) );
  NAND U45350 ( .A(n56330), .B(n25427), .Z(n40364) );
  NAND U45351 ( .A(n25428), .B(n56329), .Z(n40358) );
  AND U45352 ( .A(n25430), .B(n25429), .Z(n40356) );
  NANDN U45353 ( .A(x[4092]), .B(y[4092]), .Z(n51712) );
  AND U45354 ( .A(n51712), .B(n25431), .Z(n40354) );
  NAND U45355 ( .A(n25433), .B(n25432), .Z(n40352) );
  AND U45356 ( .A(n25434), .B(n51711), .Z(n40350) );
  NANDN U45357 ( .A(x[4088]), .B(y[4088]), .Z(n25436) );
  AND U45358 ( .A(n25436), .B(n25435), .Z(n40344) );
  AND U45359 ( .A(n25438), .B(n25437), .Z(n40334) );
  AND U45360 ( .A(n25440), .B(n25439), .Z(n40329) );
  AND U45361 ( .A(n25442), .B(n25441), .Z(n40325) );
  ANDN U45362 ( .B(y[4080]), .A(x[4080]), .Z(n40323) );
  AND U45363 ( .A(n25444), .B(n25443), .Z(n40316) );
  AND U45364 ( .A(n25446), .B(n25445), .Z(n40314) );
  NAND U45365 ( .A(n25448), .B(n25447), .Z(n40312) );
  AND U45366 ( .A(n25450), .B(n25449), .Z(n40310) );
  NAND U45367 ( .A(n25452), .B(n25451), .Z(n40300) );
  NAND U45368 ( .A(n25454), .B(n25453), .Z(n40294) );
  NANDN U45369 ( .A(x[4068]), .B(y[4068]), .Z(n25456) );
  NAND U45370 ( .A(n25456), .B(n25455), .Z(n40288) );
  NAND U45371 ( .A(n25458), .B(n25457), .Z(n40282) );
  AND U45372 ( .A(n25460), .B(n25459), .Z(n40280) );
  NAND U45373 ( .A(n25462), .B(n25461), .Z(n40278) );
  AND U45374 ( .A(n25464), .B(n25463), .Z(n40272) );
  NANDN U45375 ( .A(x[4060]), .B(y[4060]), .Z(n25466) );
  AND U45376 ( .A(n25466), .B(n25465), .Z(n40266) );
  AND U45377 ( .A(n25468), .B(n25467), .Z(n40252) );
  NAND U45378 ( .A(n25470), .B(n25469), .Z(n40242) );
  NAND U45379 ( .A(n25472), .B(n25471), .Z(n40236) );
  NAND U45380 ( .A(n25474), .B(n25473), .Z(n40230) );
  NANDN U45381 ( .A(x[4048]), .B(y[4048]), .Z(n25476) );
  AND U45382 ( .A(n25476), .B(n25475), .Z(n40228) );
  NAND U45383 ( .A(n25478), .B(n25477), .Z(n40226) );
  NAND U45384 ( .A(n25480), .B(n25479), .Z(n40216) );
  NAND U45385 ( .A(n25482), .B(n25481), .Z(n40210) );
  NAND U45386 ( .A(n25484), .B(n25483), .Z(n40204) );
  AND U45387 ( .A(n25486), .B(n25485), .Z(n40202) );
  NAND U45388 ( .A(n25488), .B(n25487), .Z(n40200) );
  AND U45389 ( .A(n25490), .B(n25489), .Z(n40194) );
  NANDN U45390 ( .A(x[4034]), .B(y[4034]), .Z(n56279) );
  AND U45391 ( .A(n25491), .B(n56279), .Z(n40188) );
  NANDN U45392 ( .A(x[4032]), .B(y[4032]), .Z(n56276) );
  AND U45393 ( .A(n56276), .B(n56278), .Z(n40182) );
  AND U45394 ( .A(n25492), .B(n51731), .Z(n40176) );
  AND U45395 ( .A(n25494), .B(n25493), .Z(n40174) );
  NANDN U45396 ( .A(x[4028]), .B(y[4028]), .Z(n56271) );
  AND U45397 ( .A(n25495), .B(n56271), .Z(n40172) );
  NAND U45398 ( .A(n25497), .B(n25496), .Z(n40170) );
  AND U45399 ( .A(n25498), .B(n56273), .Z(n40168) );
  AND U45400 ( .A(n25500), .B(n25499), .Z(n40162) );
  AND U45401 ( .A(n25502), .B(n25501), .Z(n40156) );
  AND U45402 ( .A(n25504), .B(n25503), .Z(n40150) );
  AND U45403 ( .A(n25506), .B(n25505), .Z(n40144) );
  AND U45404 ( .A(n25508), .B(n25507), .Z(n40138) );
  NANDN U45405 ( .A(x[4014]), .B(y[4014]), .Z(n25510) );
  AND U45406 ( .A(n25510), .B(n25509), .Z(n40132) );
  AND U45407 ( .A(n25512), .B(n25511), .Z(n40122) );
  AND U45408 ( .A(n25514), .B(n25513), .Z(n40116) );
  ANDN U45409 ( .B(y[4008]), .A(x[4008]), .Z(n40114) );
  NAND U45410 ( .A(n25516), .B(n25515), .Z(n40110) );
  NAND U45411 ( .A(n25518), .B(n25517), .Z(n40104) );
  AND U45412 ( .A(n25520), .B(n25519), .Z(n40102) );
  NAND U45413 ( .A(n25522), .B(n25521), .Z(n40100) );
  NAND U45414 ( .A(n25524), .B(n25523), .Z(n40095) );
  NANDN U45415 ( .A(x[4000]), .B(y[4000]), .Z(n51742) );
  AND U45416 ( .A(n51742), .B(n56245), .Z(n40093) );
  NANDN U45417 ( .A(x[3998]), .B(y[3998]), .Z(n56242) );
  AND U45418 ( .A(n25526), .B(n25525), .Z(n40085) );
  AND U45419 ( .A(n56241), .B(n25527), .Z(n40083) );
  NAND U45420 ( .A(n25529), .B(n25528), .Z(n40081) );
  NANDN U45421 ( .A(x[3994]), .B(y[3994]), .Z(n51744) );
  AND U45422 ( .A(n51744), .B(n25530), .Z(n40079) );
  NAND U45423 ( .A(n25532), .B(n25531), .Z(n40071) );
  AND U45424 ( .A(n25534), .B(n25533), .Z(n40066) );
  NANDN U45425 ( .A(x[3988]), .B(y[3988]), .Z(n51746) );
  NAND U45426 ( .A(n51746), .B(n25535), .Z(n40064) );
  AND U45427 ( .A(n25537), .B(n25536), .Z(n40062) );
  NAND U45428 ( .A(n25539), .B(n25538), .Z(n40057) );
  NAND U45429 ( .A(n25541), .B(n25540), .Z(n40052) );
  AND U45430 ( .A(n25542), .B(n56227), .Z(n40050) );
  NANDN U45431 ( .A(x[3980]), .B(y[3980]), .Z(n25544) );
  NAND U45432 ( .A(n25544), .B(n25543), .Z(n40044) );
  NAND U45433 ( .A(n25546), .B(n25545), .Z(n40038) );
  NANDN U45434 ( .A(x[3976]), .B(y[3976]), .Z(n25548) );
  NAND U45435 ( .A(n25548), .B(n25547), .Z(n40032) );
  ANDN U45436 ( .B(y[3974]), .A(x[3974]), .Z(n40024) );
  AND U45437 ( .A(n25550), .B(n25549), .Z(n40022) );
  NANDN U45438 ( .A(x[3972]), .B(y[3972]), .Z(n25551) );
  AND U45439 ( .A(n25552), .B(n25551), .Z(n40020) );
  NAND U45440 ( .A(n25554), .B(n25553), .Z(n40018) );
  NANDN U45441 ( .A(x[3970]), .B(y[3970]), .Z(n25556) );
  AND U45442 ( .A(n25556), .B(n25555), .Z(n40016) );
  NAND U45443 ( .A(n25558), .B(n25557), .Z(n40002) );
  AND U45444 ( .A(n25560), .B(n25559), .Z(n40000) );
  ANDN U45445 ( .B(y[3964]), .A(x[3964]), .Z(n56207) );
  NAND U45446 ( .A(n25562), .B(n25561), .Z(n39995) );
  NAND U45447 ( .A(n25564), .B(n25563), .Z(n39990) );
  AND U45448 ( .A(n25566), .B(n25565), .Z(n39988) );
  NAND U45449 ( .A(n25568), .B(n25567), .Z(n39986) );
  AND U45450 ( .A(n25569), .B(n56199), .Z(n39977) );
  NAND U45451 ( .A(n51754), .B(n25570), .Z(n39971) );
  XNOR U45452 ( .A(y[3952]), .B(x[3952]), .Z(n25573) );
  AND U45453 ( .A(n25573), .B(n25572), .Z(n39965) );
  IV U45454 ( .A(n25574), .Z(n56194) );
  AND U45455 ( .A(n25575), .B(n56194), .Z(n39963) );
  NAND U45456 ( .A(n25577), .B(n25576), .Z(n39961) );
  NANDN U45457 ( .A(x[3948]), .B(y[3948]), .Z(n25579) );
  AND U45458 ( .A(n25579), .B(n25578), .Z(n39959) );
  NAND U45459 ( .A(n25581), .B(n25580), .Z(n39957) );
  AND U45460 ( .A(n25583), .B(n25582), .Z(n39951) );
  AND U45461 ( .A(n25585), .B(n25584), .Z(n39945) );
  NAND U45462 ( .A(n25587), .B(n25586), .Z(n39943) );
  AND U45463 ( .A(n25589), .B(n25588), .Z(n39941) );
  NAND U45464 ( .A(n25591), .B(n25590), .Z(n39935) );
  NAND U45465 ( .A(n25593), .B(n25592), .Z(n39929) );
  AND U45466 ( .A(n25595), .B(n25594), .Z(n39927) );
  NAND U45467 ( .A(n25597), .B(n25596), .Z(n39925) );
  AND U45468 ( .A(n25598), .B(n51761), .Z(n39910) );
  AND U45469 ( .A(n25600), .B(n25599), .Z(n39908) );
  NAND U45470 ( .A(n25602), .B(n25601), .Z(n39906) );
  AND U45471 ( .A(n25604), .B(n25603), .Z(n39904) );
  AND U45472 ( .A(n25606), .B(n25605), .Z(n39898) );
  AND U45473 ( .A(n25608), .B(n25607), .Z(n39892) );
  AND U45474 ( .A(n25610), .B(n25609), .Z(n39886) );
  NAND U45475 ( .A(n25612), .B(n25611), .Z(n39876) );
  NAND U45476 ( .A(n25614), .B(n25613), .Z(n39870) );
  NAND U45477 ( .A(n25616), .B(n25615), .Z(n39864) );
  AND U45478 ( .A(n25618), .B(n25617), .Z(n39862) );
  NAND U45479 ( .A(n25620), .B(n25619), .Z(n39860) );
  NANDN U45480 ( .A(x[3910]), .B(y[3910]), .Z(n25622) );
  AND U45481 ( .A(n25622), .B(n25621), .Z(n39854) );
  NANDN U45482 ( .A(x[3908]), .B(y[3908]), .Z(n25624) );
  AND U45483 ( .A(n25624), .B(n25623), .Z(n39848) );
  AND U45484 ( .A(n25626), .B(n25625), .Z(n39842) );
  NANDN U45485 ( .A(x[3904]), .B(y[3904]), .Z(n25628) );
  AND U45486 ( .A(n25628), .B(n25627), .Z(n39836) );
  NANDN U45487 ( .A(x[3902]), .B(y[3902]), .Z(n25630) );
  AND U45488 ( .A(n25630), .B(n25629), .Z(n39830) );
  NANDN U45489 ( .A(x[3898]), .B(y[3898]), .Z(n25632) );
  NAND U45490 ( .A(n25632), .B(n25631), .Z(n39816) );
  AND U45491 ( .A(n25634), .B(n25633), .Z(n39814) );
  NAND U45492 ( .A(n25636), .B(n25635), .Z(n39808) );
  AND U45493 ( .A(n25638), .B(n25637), .Z(n39802) );
  AND U45494 ( .A(n25640), .B(n25639), .Z(n39796) );
  AND U45495 ( .A(n25642), .B(n25641), .Z(n39794) );
  NAND U45496 ( .A(n25644), .B(n25643), .Z(n39792) );
  AND U45497 ( .A(n25645), .B(n56136), .Z(n39783) );
  AND U45498 ( .A(n25647), .B(n25646), .Z(n39781) );
  NAND U45499 ( .A(n25649), .B(n25648), .Z(n39779) );
  AND U45500 ( .A(n25651), .B(n25650), .Z(n39777) );
  NANDN U45501 ( .A(x[3882]), .B(y[3882]), .Z(n56129) );
  NAND U45502 ( .A(n56129), .B(n25652), .Z(n39775) );
  NANDN U45503 ( .A(x[3880]), .B(y[3880]), .Z(n56126) );
  NAND U45504 ( .A(n56126), .B(n56128), .Z(n39769) );
  NANDN U45505 ( .A(x[3878]), .B(y[3878]), .Z(n51775) );
  AND U45506 ( .A(n25654), .B(n25653), .Z(n39761) );
  IV U45507 ( .A(n25655), .Z(n51774) );
  AND U45508 ( .A(n25656), .B(n51774), .Z(n39759) );
  NAND U45509 ( .A(n25658), .B(n25657), .Z(n39757) );
  NANDN U45510 ( .A(x[3874]), .B(y[3874]), .Z(n56120) );
  AND U45511 ( .A(n56120), .B(n25659), .Z(n39755) );
  NAND U45512 ( .A(n25661), .B(n25660), .Z(n39742) );
  AND U45513 ( .A(n25663), .B(n25662), .Z(n39740) );
  NAND U45514 ( .A(n25665), .B(n25664), .Z(n39734) );
  NAND U45515 ( .A(n25667), .B(n25666), .Z(n39728) );
  AND U45516 ( .A(n25669), .B(n25668), .Z(n39726) );
  NAND U45517 ( .A(n25671), .B(n25670), .Z(n39724) );
  NAND U45518 ( .A(n25673), .B(n25672), .Z(n39714) );
  NAND U45519 ( .A(n25675), .B(n25674), .Z(n39708) );
  NAND U45520 ( .A(n25677), .B(n25676), .Z(n39702) );
  ANDN U45521 ( .B(y[3854]), .A(x[3854]), .Z(n56102) );
  AND U45522 ( .A(n25679), .B(n25678), .Z(n39693) );
  IV U45523 ( .A(n25680), .Z(n56101) );
  AND U45524 ( .A(n25681), .B(n56101), .Z(n39691) );
  NAND U45525 ( .A(n25683), .B(n25682), .Z(n39689) );
  AND U45526 ( .A(n25685), .B(n25684), .Z(n39687) );
  NAND U45527 ( .A(n25687), .B(n25686), .Z(n39677) );
  NAND U45528 ( .A(n25689), .B(n25688), .Z(n39671) );
  AND U45529 ( .A(n25691), .B(n25690), .Z(n39669) );
  NAND U45530 ( .A(n25693), .B(n25692), .Z(n39667) );
  NAND U45531 ( .A(n56088), .B(n25694), .Z(n39652) );
  NANDN U45532 ( .A(x[3836]), .B(y[3836]), .Z(n56081) );
  NAND U45533 ( .A(n56081), .B(n25695), .Z(n39646) );
  ANDN U45534 ( .B(y[3834]), .A(x[3834]), .Z(n51785) );
  AND U45535 ( .A(n25697), .B(n25696), .Z(n39638) );
  NANDN U45536 ( .A(x[3832]), .B(y[3832]), .Z(n51788) );
  AND U45537 ( .A(n51788), .B(n51786), .Z(n39636) );
  NAND U45538 ( .A(n25699), .B(n25698), .Z(n39634) );
  AND U45539 ( .A(n25700), .B(n51787), .Z(n39632) );
  NANDN U45540 ( .A(x[3828]), .B(y[3828]), .Z(n25702) );
  AND U45541 ( .A(n25702), .B(n25701), .Z(n39626) );
  NANDN U45542 ( .A(x[3826]), .B(y[3826]), .Z(n25704) );
  AND U45543 ( .A(n25704), .B(n25703), .Z(n39620) );
  NANDN U45544 ( .A(x[3824]), .B(y[3824]), .Z(n25706) );
  AND U45545 ( .A(n25706), .B(n25705), .Z(n39614) );
  NANDN U45546 ( .A(x[3822]), .B(y[3822]), .Z(n25708) );
  AND U45547 ( .A(n25708), .B(n25707), .Z(n39608) );
  NANDN U45548 ( .A(x[3820]), .B(y[3820]), .Z(n25710) );
  AND U45549 ( .A(n25710), .B(n25709), .Z(n39602) );
  NAND U45550 ( .A(n25712), .B(n25711), .Z(n39600) );
  NAND U45551 ( .A(n25714), .B(n25713), .Z(n39594) );
  AND U45552 ( .A(n25716), .B(n25715), .Z(n39580) );
  AND U45553 ( .A(n25718), .B(n25717), .Z(n39574) );
  AND U45554 ( .A(n25720), .B(n25719), .Z(n39568) );
  AND U45555 ( .A(n25722), .B(n25721), .Z(n39562) );
  NAND U45556 ( .A(n25724), .B(n25723), .Z(n39548) );
  AND U45557 ( .A(n56049), .B(n25725), .Z(n39546) );
  NAND U45558 ( .A(n25729), .B(n25728), .Z(n39540) );
  NANDN U45559 ( .A(x[3798]), .B(y[3798]), .Z(n51797) );
  AND U45560 ( .A(n56047), .B(n51797), .Z(n39538) );
  NAND U45561 ( .A(n25731), .B(n25730), .Z(n39536) );
  NANDN U45562 ( .A(x[3796]), .B(y[3796]), .Z(n39533) );
  NAND U45563 ( .A(n25733), .B(n25732), .Z(n39531) );
  NAND U45564 ( .A(n25735), .B(n25734), .Z(n39525) );
  AND U45565 ( .A(n25737), .B(n25736), .Z(n39523) );
  NAND U45566 ( .A(n25739), .B(n25738), .Z(n39521) );
  AND U45567 ( .A(n25741), .B(n25740), .Z(n39511) );
  AND U45568 ( .A(n25743), .B(n25742), .Z(n39509) );
  NAND U45569 ( .A(n25745), .B(n25744), .Z(n39507) );
  AND U45570 ( .A(n25747), .B(n25746), .Z(n39505) );
  NAND U45571 ( .A(n25749), .B(n25748), .Z(n39495) );
  NANDN U45572 ( .A(x[3780]), .B(y[3780]), .Z(n56027) );
  NAND U45573 ( .A(n56027), .B(n25750), .Z(n39489) );
  ANDN U45574 ( .B(y[3778]), .A(x[3778]), .Z(n56024) );
  AND U45575 ( .A(n25752), .B(n25751), .Z(n39481) );
  NANDN U45576 ( .A(x[3776]), .B(y[3776]), .Z(n56020) );
  AND U45577 ( .A(n56023), .B(n56020), .Z(n39479) );
  NAND U45578 ( .A(n25754), .B(n25753), .Z(n39477) );
  AND U45579 ( .A(n25755), .B(n56021), .Z(n39475) );
  NANDN U45580 ( .A(x[3772]), .B(y[3772]), .Z(n56017) );
  AND U45581 ( .A(n25756), .B(n56017), .Z(n39469) );
  AND U45582 ( .A(n25758), .B(n25757), .Z(n39460) );
  NAND U45583 ( .A(n25760), .B(n25759), .Z(n39458) );
  AND U45584 ( .A(n25762), .B(n25761), .Z(n39456) );
  NAND U45585 ( .A(n25764), .B(n25763), .Z(n39454) );
  AND U45586 ( .A(n25766), .B(n25765), .Z(n39448) );
  AND U45587 ( .A(n25768), .B(n25767), .Z(n39442) );
  AND U45588 ( .A(n25770), .B(n25769), .Z(n39432) );
  AND U45589 ( .A(n25772), .B(n25771), .Z(n39426) );
  AND U45590 ( .A(n25774), .B(n25773), .Z(n39420) );
  AND U45591 ( .A(n25776), .B(n25775), .Z(n39414) );
  AND U45592 ( .A(n25778), .B(n25777), .Z(n39412) );
  NAND U45593 ( .A(n25780), .B(n25779), .Z(n39410) );
  AND U45594 ( .A(n25782), .B(n25781), .Z(n39400) );
  AND U45595 ( .A(n25784), .B(n25783), .Z(n39398) );
  NAND U45596 ( .A(n25786), .B(n25785), .Z(n39396) );
  NAND U45597 ( .A(n25788), .B(n25787), .Z(n39390) );
  NAND U45598 ( .A(n25790), .B(n25789), .Z(n39384) );
  NAND U45599 ( .A(n25792), .B(n25791), .Z(n39378) );
  AND U45600 ( .A(n25794), .B(n25793), .Z(n39376) );
  NAND U45601 ( .A(n25796), .B(n25795), .Z(n39374) );
  AND U45602 ( .A(n25798), .B(n25797), .Z(n39368) );
  AND U45603 ( .A(n25800), .B(n25799), .Z(n39362) );
  NANDN U45604 ( .A(x[3732]), .B(y[3732]), .Z(n51814) );
  AND U45605 ( .A(n51814), .B(n25801), .Z(n39356) );
  NANDN U45606 ( .A(x[3730]), .B(y[3730]), .Z(n55984) );
  IV U45607 ( .A(n25802), .Z(n51813) );
  AND U45608 ( .A(n55984), .B(n51813), .Z(n39350) );
  AND U45609 ( .A(n25803), .B(n55983), .Z(n39344) );
  NAND U45610 ( .A(n25805), .B(n25804), .Z(n39342) );
  NAND U45611 ( .A(n25807), .B(n25806), .Z(n39336) );
  NANDN U45612 ( .A(x[3724]), .B(y[3724]), .Z(n55975) );
  NANDN U45613 ( .A(x[3722]), .B(y[3722]), .Z(n55971) );
  AND U45614 ( .A(n55971), .B(n55974), .Z(n39327) );
  NAND U45615 ( .A(n25809), .B(n25808), .Z(n39325) );
  IV U45616 ( .A(n25810), .Z(n55972) );
  AND U45617 ( .A(n25811), .B(n55972), .Z(n39323) );
  AND U45618 ( .A(n25813), .B(n25812), .Z(n39321) );
  AND U45619 ( .A(n25815), .B(n25814), .Z(n39315) );
  AND U45620 ( .A(n25817), .B(n25816), .Z(n39309) );
  AND U45621 ( .A(n25819), .B(n25818), .Z(n39303) );
  NAND U45622 ( .A(n25821), .B(n25820), .Z(n39293) );
  NAND U45623 ( .A(n25823), .B(n25822), .Z(n39287) );
  NAND U45624 ( .A(n25825), .B(n25824), .Z(n39278) );
  AND U45625 ( .A(n25826), .B(n55957), .Z(n39276) );
  AND U45626 ( .A(n25828), .B(n25827), .Z(n39274) );
  NAND U45627 ( .A(n25830), .B(n25829), .Z(n39272) );
  AND U45628 ( .A(n25832), .B(n25831), .Z(n39270) );
  NAND U45629 ( .A(n25834), .B(n25833), .Z(n39264) );
  NAND U45630 ( .A(n25836), .B(n25835), .Z(n39258) );
  AND U45631 ( .A(n25838), .B(n25837), .Z(n39256) );
  NAND U45632 ( .A(n25840), .B(n25839), .Z(n39254) );
  AND U45633 ( .A(n25841), .B(n55946), .Z(n39245) );
  AND U45634 ( .A(n25843), .B(n25842), .Z(n39243) );
  NAND U45635 ( .A(n25845), .B(n25844), .Z(n39241) );
  AND U45636 ( .A(n25847), .B(n25846), .Z(n39239) );
  AND U45637 ( .A(n25849), .B(n25848), .Z(n39233) );
  AND U45638 ( .A(n25851), .B(n25850), .Z(n39227) );
  AND U45639 ( .A(n25853), .B(n25852), .Z(n39221) );
  AND U45640 ( .A(n25855), .B(n25854), .Z(n39211) );
  NAND U45641 ( .A(n25857), .B(n25856), .Z(n39209) );
  AND U45642 ( .A(n25859), .B(n25858), .Z(n39207) );
  NAND U45643 ( .A(n25861), .B(n25860), .Z(n39205) );
  AND U45644 ( .A(n25863), .B(n25862), .Z(n39199) );
  NAND U45645 ( .A(n25865), .B(n25864), .Z(n39197) );
  AND U45646 ( .A(n25867), .B(n25866), .Z(n39195) );
  AND U45647 ( .A(n25869), .B(n25868), .Z(n39193) );
  NAND U45648 ( .A(n25871), .B(n25870), .Z(n39191) );
  NAND U45649 ( .A(n25873), .B(n25872), .Z(n39181) );
  NAND U45650 ( .A(n25875), .B(n25874), .Z(n39175) );
  NAND U45651 ( .A(n25877), .B(n25876), .Z(n39169) );
  AND U45652 ( .A(n25879), .B(n25878), .Z(n39167) );
  AND U45653 ( .A(n25881), .B(n25880), .Z(n39162) );
  AND U45654 ( .A(n55920), .B(n25882), .Z(n39160) );
  NAND U45655 ( .A(n25884), .B(n25883), .Z(n39158) );
  AND U45656 ( .A(n25886), .B(n25885), .Z(n39156) );
  AND U45657 ( .A(n25888), .B(n25887), .Z(n39154) );
  NANDN U45658 ( .A(x[3656]), .B(y[3656]), .Z(n55915) );
  AND U45659 ( .A(n55915), .B(n25889), .Z(n39152) );
  NAND U45660 ( .A(n25891), .B(n25890), .Z(n39150) );
  AND U45661 ( .A(n25892), .B(n55914), .Z(n39148) );
  NAND U45662 ( .A(n25894), .B(n25893), .Z(n39146) );
  ANDN U45663 ( .B(y[3652]), .A(x[3652]), .Z(n39142) );
  AND U45664 ( .A(n25896), .B(n25895), .Z(n39140) );
  AND U45665 ( .A(n25897), .B(n55907), .Z(n39134) );
  AND U45666 ( .A(n25898), .B(n55906), .Z(n39132) );
  NAND U45667 ( .A(n25900), .B(n25899), .Z(n39130) );
  NANDN U45668 ( .A(x[3644]), .B(y[3644]), .Z(n25901) );
  NAND U45669 ( .A(n25901), .B(n51837), .Z(n39122) );
  NAND U45670 ( .A(n25903), .B(n25902), .Z(n39116) );
  AND U45671 ( .A(n25905), .B(n25904), .Z(n39102) );
  NANDN U45672 ( .A(x[3636]), .B(y[3636]), .Z(n25907) );
  AND U45673 ( .A(n25907), .B(n25906), .Z(n39096) );
  AND U45674 ( .A(n25909), .B(n25908), .Z(n39090) );
  AND U45675 ( .A(n25911), .B(n25910), .Z(n39084) );
  NANDN U45676 ( .A(x[3630]), .B(y[3630]), .Z(n51845) );
  AND U45677 ( .A(n51845), .B(n25912), .Z(n39078) );
  NAND U45678 ( .A(n25914), .B(n25913), .Z(n39068) );
  NAND U45679 ( .A(n25916), .B(n25915), .Z(n39062) );
  NAND U45680 ( .A(n25918), .B(n25917), .Z(n39056) );
  AND U45681 ( .A(n25920), .B(n25919), .Z(n39050) );
  AND U45682 ( .A(n25922), .B(n25921), .Z(n39044) );
  AND U45683 ( .A(n25924), .B(n25923), .Z(n39034) );
  NAND U45684 ( .A(n25926), .B(n25925), .Z(n39032) );
  NAND U45685 ( .A(n25928), .B(n25927), .Z(n39027) );
  AND U45686 ( .A(n25930), .B(n25929), .Z(n39022) );
  AND U45687 ( .A(n25932), .B(n25931), .Z(n39016) );
  AND U45688 ( .A(n25934), .B(n25933), .Z(n39010) );
  AND U45689 ( .A(n25936), .B(n25935), .Z(n39004) );
  NAND U45690 ( .A(n25938), .B(n25937), .Z(n38994) );
  NAND U45691 ( .A(n25940), .B(n25939), .Z(n38988) );
  NANDN U45692 ( .A(x[3598]), .B(y[3598]), .Z(n25942) );
  NAND U45693 ( .A(n25942), .B(n25941), .Z(n38982) );
  AND U45694 ( .A(n25944), .B(n25943), .Z(n38972) );
  ANDN U45695 ( .B(y[3594]), .A(x[3594]), .Z(n25946) );
  NOR U45696 ( .A(n25946), .B(n25945), .Z(n38970) );
  AND U45697 ( .A(n25948), .B(n25947), .Z(n38964) );
  AND U45698 ( .A(n25950), .B(n25949), .Z(n38954) );
  NANDN U45699 ( .A(x[3586]), .B(y[3586]), .Z(n25952) );
  AND U45700 ( .A(n25952), .B(n25951), .Z(n38944) );
  NANDN U45701 ( .A(x[3584]), .B(y[3584]), .Z(n55849) );
  AND U45702 ( .A(n55849), .B(n25953), .Z(n38938) );
  AND U45703 ( .A(n25954), .B(n55848), .Z(n38932) );
  NAND U45704 ( .A(n25956), .B(n25955), .Z(n38930) );
  AND U45705 ( .A(n25958), .B(n25957), .Z(n38916) );
  AND U45706 ( .A(n25960), .B(n25959), .Z(n38910) );
  AND U45707 ( .A(n25962), .B(n25961), .Z(n38904) );
  NAND U45708 ( .A(n25964), .B(n25963), .Z(n38899) );
  IV U45709 ( .A(n25965), .Z(n55836) );
  AND U45710 ( .A(n25966), .B(n55836), .Z(n38897) );
  NAND U45711 ( .A(n25968), .B(n25967), .Z(n38895) );
  AND U45712 ( .A(n25969), .B(n55831), .Z(n38886) );
  AND U45713 ( .A(n25971), .B(n25970), .Z(n38884) );
  NAND U45714 ( .A(n25973), .B(n25972), .Z(n38882) );
  AND U45715 ( .A(n25975), .B(n25974), .Z(n38880) );
  AND U45716 ( .A(n25977), .B(n25976), .Z(n38874) );
  AND U45717 ( .A(n25979), .B(n25978), .Z(n38868) );
  AND U45718 ( .A(n25981), .B(n25980), .Z(n38862) );
  NAND U45719 ( .A(n25983), .B(n25982), .Z(n38848) );
  AND U45720 ( .A(n25985), .B(n25984), .Z(n38846) );
  NANDN U45721 ( .A(x[3550]), .B(y[3550]), .Z(n55815) );
  AND U45722 ( .A(n25986), .B(n55815), .Z(n38840) );
  XNOR U45723 ( .A(y[3550]), .B(x[3550]), .Z(n38836) );
  AND U45724 ( .A(n25988), .B(n25987), .Z(n38831) );
  NAND U45725 ( .A(n25990), .B(n25989), .Z(n38829) );
  AND U45726 ( .A(n25992), .B(n25991), .Z(n38823) );
  NANDN U45727 ( .A(x[3542]), .B(y[3542]), .Z(n51866) );
  AND U45728 ( .A(n51866), .B(n25993), .Z(n38817) );
  AND U45729 ( .A(n25994), .B(n51865), .Z(n38811) );
  NAND U45730 ( .A(n25996), .B(n25995), .Z(n38809) );
  AND U45731 ( .A(n25998), .B(n25997), .Z(n38803) );
  AND U45732 ( .A(n26000), .B(n25999), .Z(n38798) );
  IV U45733 ( .A(n26001), .Z(n55800) );
  AND U45734 ( .A(n26002), .B(n55800), .Z(n38796) );
  NAND U45735 ( .A(n26004), .B(n26003), .Z(n38794) );
  IV U45736 ( .A(n26005), .Z(n51869) );
  NAND U45737 ( .A(n51869), .B(n26006), .Z(n38785) );
  NAND U45738 ( .A(n26008), .B(n26007), .Z(n38779) );
  ANDN U45739 ( .B(y[3526]), .A(x[3526]), .Z(n55794) );
  AND U45740 ( .A(n26010), .B(n26009), .Z(n38770) );
  AND U45741 ( .A(n55795), .B(n26011), .Z(n38768) );
  NAND U45742 ( .A(n26013), .B(n26012), .Z(n38766) );
  AND U45743 ( .A(n26015), .B(n26014), .Z(n38764) );
  NANDN U45744 ( .A(x[3518]), .B(y[3518]), .Z(n26017) );
  AND U45745 ( .A(n26017), .B(n26016), .Z(n38750) );
  NAND U45746 ( .A(n26019), .B(n26018), .Z(n38740) );
  NAND U45747 ( .A(n26021), .B(n26020), .Z(n38734) );
  NAND U45748 ( .A(n26023), .B(n26022), .Z(n38728) );
  NAND U45749 ( .A(n26025), .B(n26024), .Z(n38722) );
  AND U45750 ( .A(n26027), .B(n26026), .Z(n38720) );
  NAND U45751 ( .A(n26029), .B(n26028), .Z(n38718) );
  NAND U45752 ( .A(n26030), .B(n55774), .Z(n38709) );
  NAND U45753 ( .A(n26032), .B(n26031), .Z(n38703) );
  NAND U45754 ( .A(n26034), .B(n26033), .Z(n38697) );
  AND U45755 ( .A(n26036), .B(n26035), .Z(n38695) );
  AND U45756 ( .A(n26037), .B(n55766), .Z(n38693) );
  NAND U45757 ( .A(n51878), .B(n26038), .Z(n38691) );
  AND U45758 ( .A(n26041), .B(n26040), .Z(n38688) );
  AND U45759 ( .A(n26042), .B(n55764), .Z(n38686) );
  NAND U45760 ( .A(n26044), .B(n26043), .Z(n38684) );
  AND U45761 ( .A(n26046), .B(n26045), .Z(n38682) );
  AND U45762 ( .A(n26048), .B(n26047), .Z(n38676) );
  NANDN U45763 ( .A(x[3488]), .B(y[3488]), .Z(n26050) );
  AND U45764 ( .A(n26050), .B(n26049), .Z(n38670) );
  NAND U45765 ( .A(n26052), .B(n26051), .Z(n38668) );
  NAND U45766 ( .A(n26054), .B(n26053), .Z(n38654) );
  NAND U45767 ( .A(n26056), .B(n26055), .Z(n38648) );
  AND U45768 ( .A(n26058), .B(n26057), .Z(n38646) );
  NAND U45769 ( .A(n26060), .B(n26059), .Z(n38644) );
  AND U45770 ( .A(n26061), .B(n51881), .Z(n38635) );
  AND U45771 ( .A(n26063), .B(n26062), .Z(n38633) );
  NAND U45772 ( .A(n26065), .B(n26064), .Z(n38631) );
  AND U45773 ( .A(n26067), .B(n26066), .Z(n38629) );
  NAND U45774 ( .A(n26069), .B(n26068), .Z(n38619) );
  NAND U45775 ( .A(n26071), .B(n26070), .Z(n38613) );
  NAND U45776 ( .A(n26073), .B(n26072), .Z(n38607) );
  NAND U45777 ( .A(n26075), .B(n26074), .Z(n38601) );
  NANDN U45778 ( .A(x[3462]), .B(y[3462]), .Z(n55716) );
  NAND U45779 ( .A(n55716), .B(n26076), .Z(n38595) );
  AND U45780 ( .A(n26077), .B(n55715), .Z(n38589) );
  AND U45781 ( .A(n26079), .B(n26078), .Z(n38587) );
  NAND U45782 ( .A(n26081), .B(n26080), .Z(n38585) );
  AND U45783 ( .A(n26083), .B(n26082), .Z(n38583) );
  NAND U45784 ( .A(n26085), .B(n26084), .Z(n38581) );
  AND U45785 ( .A(n26087), .B(n26086), .Z(n38579) );
  AND U45786 ( .A(n26089), .B(n26088), .Z(n38577) );
  NAND U45787 ( .A(n26091), .B(n26090), .Z(n38575) );
  AND U45788 ( .A(n26093), .B(n26092), .Z(n38573) );
  NAND U45789 ( .A(n26095), .B(n26094), .Z(n38571) );
  NAND U45790 ( .A(n26097), .B(n26096), .Z(n38565) );
  NAND U45791 ( .A(n26099), .B(n26098), .Z(n38559) );
  NAND U45792 ( .A(n26101), .B(n26100), .Z(n38553) );
  AND U45793 ( .A(n26103), .B(n26102), .Z(n38551) );
  NAND U45794 ( .A(n26105), .B(n26104), .Z(n38549) );
  AND U45795 ( .A(n26107), .B(n26106), .Z(n38543) );
  AND U45796 ( .A(n26109), .B(n26108), .Z(n38537) );
  NANDN U45797 ( .A(x[3438]), .B(y[3438]), .Z(n26111) );
  NAND U45798 ( .A(n26111), .B(n26110), .Z(n38535) );
  AND U45799 ( .A(n26113), .B(n26112), .Z(n38525) );
  AND U45800 ( .A(n26115), .B(n26114), .Z(n38519) );
  AND U45801 ( .A(n26116), .B(n55658), .Z(n38510) );
  AND U45802 ( .A(n26118), .B(n26117), .Z(n38508) );
  NAND U45803 ( .A(n26120), .B(n26119), .Z(n38506) );
  AND U45804 ( .A(n26122), .B(n26121), .Z(n38504) );
  NAND U45805 ( .A(n26123), .B(n55649), .Z(n38487) );
  NAND U45806 ( .A(n26125), .B(n26124), .Z(n38481) );
  ANDN U45807 ( .B(y[3418]), .A(x[3418]), .Z(n55642) );
  AND U45808 ( .A(n26127), .B(n26126), .Z(n38472) );
  AND U45809 ( .A(n55641), .B(n26128), .Z(n38470) );
  NAND U45810 ( .A(n26130), .B(n26129), .Z(n38468) );
  AND U45811 ( .A(n26132), .B(n26131), .Z(n38466) );
  AND U45812 ( .A(n26134), .B(n26133), .Z(n38460) );
  AND U45813 ( .A(n26136), .B(n26135), .Z(n38454) );
  NANDN U45814 ( .A(x[3408]), .B(y[3408]), .Z(n55631) );
  AND U45815 ( .A(n26137), .B(n55631), .Z(n38448) );
  AND U45816 ( .A(n26138), .B(n51883), .Z(n38442) );
  AND U45817 ( .A(n26140), .B(n26139), .Z(n38436) );
  AND U45818 ( .A(n26142), .B(n26141), .Z(n38430) );
  NANDN U45819 ( .A(x[3400]), .B(y[3400]), .Z(n26144) );
  AND U45820 ( .A(n26144), .B(n26143), .Z(n38424) );
  NANDN U45821 ( .A(x[3398]), .B(y[3398]), .Z(n55621) );
  AND U45822 ( .A(n55621), .B(n26145), .Z(n38418) );
  NANDN U45823 ( .A(x[3396]), .B(y[3396]), .Z(n55617) );
  AND U45824 ( .A(n55617), .B(n55620), .Z(n38412) );
  NAND U45825 ( .A(n26147), .B(n26146), .Z(n38410) );
  NAND U45826 ( .A(n26149), .B(n26148), .Z(n38405) );
  AND U45827 ( .A(n26151), .B(n26150), .Z(n38403) );
  NAND U45828 ( .A(n26153), .B(n26152), .Z(n38401) );
  AND U45829 ( .A(n26155), .B(n26154), .Z(n38396) );
  IV U45830 ( .A(n26156), .Z(n55610) );
  NAND U45831 ( .A(n55610), .B(n26157), .Z(n38394) );
  AND U45832 ( .A(n26159), .B(n26158), .Z(n38392) );
  NAND U45833 ( .A(n26161), .B(n26160), .Z(n38390) );
  NAND U45834 ( .A(n26163), .B(n26162), .Z(n38384) );
  ANDN U45835 ( .B(y[3382]), .A(x[3382]), .Z(n55605) );
  AND U45836 ( .A(n26164), .B(n55604), .Z(n38371) );
  AND U45837 ( .A(n26166), .B(n26165), .Z(n38365) );
  AND U45838 ( .A(n26168), .B(n26167), .Z(n38351) );
  AND U45839 ( .A(n26170), .B(n26169), .Z(n38345) );
  AND U45840 ( .A(n26172), .B(n26171), .Z(n38339) );
  NANDN U45841 ( .A(x[3368]), .B(y[3368]), .Z(n26174) );
  AND U45842 ( .A(n26174), .B(n26173), .Z(n38333) );
  AND U45843 ( .A(n26176), .B(n26175), .Z(n38327) );
  AND U45844 ( .A(n26178), .B(n26177), .Z(n38321) );
  AND U45845 ( .A(n26180), .B(n26179), .Z(n38315) );
  AND U45846 ( .A(n26182), .B(n26181), .Z(n38309) );
  AND U45847 ( .A(n26184), .B(n26183), .Z(n38303) );
  AND U45848 ( .A(n26186), .B(n26185), .Z(n38297) );
  NAND U45849 ( .A(n26188), .B(n26187), .Z(n38295) );
  NAND U45850 ( .A(n26190), .B(n26189), .Z(n38290) );
  NAND U45851 ( .A(n26192), .B(n26191), .Z(n38285) );
  AND U45852 ( .A(n26194), .B(n26193), .Z(n38283) );
  NAND U45853 ( .A(n26196), .B(n26195), .Z(n38281) );
  NAND U45854 ( .A(n26198), .B(n26197), .Z(n38275) );
  NANDN U45855 ( .A(x[3346]), .B(y[3346]), .Z(n26200) );
  AND U45856 ( .A(n26200), .B(n26199), .Z(n38273) );
  NAND U45857 ( .A(n51905), .B(n26201), .Z(n38268) );
  NAND U45858 ( .A(n51906), .B(n26202), .Z(n38263) );
  AND U45859 ( .A(n26204), .B(n26203), .Z(n38261) );
  NANDN U45860 ( .A(x[3340]), .B(y[3340]), .Z(n26205) );
  AND U45861 ( .A(n26206), .B(n26205), .Z(n38259) );
  NAND U45862 ( .A(n26208), .B(n26207), .Z(n38257) );
  AND U45863 ( .A(n26210), .B(n26209), .Z(n38255) );
  AND U45864 ( .A(n26212), .B(n26211), .Z(n38249) );
  NANDN U45865 ( .A(x[3334]), .B(y[3334]), .Z(n26214) );
  AND U45866 ( .A(n26214), .B(n26213), .Z(n38243) );
  NANDN U45867 ( .A(x[3332]), .B(y[3332]), .Z(n26216) );
  AND U45868 ( .A(n26216), .B(n26215), .Z(n38237) );
  AND U45869 ( .A(n26218), .B(n26217), .Z(n38231) );
  NANDN U45870 ( .A(x[3328]), .B(y[3328]), .Z(n26220) );
  AND U45871 ( .A(n26220), .B(n26219), .Z(n38225) );
  AND U45872 ( .A(n26222), .B(n26221), .Z(n38211) );
  AND U45873 ( .A(n26224), .B(n26223), .Z(n38205) );
  AND U45874 ( .A(n26226), .B(n26225), .Z(n38199) );
  AND U45875 ( .A(n26228), .B(n26227), .Z(n38193) );
  AND U45876 ( .A(n26230), .B(n26229), .Z(n38187) );
  AND U45877 ( .A(n26232), .B(n26231), .Z(n38181) );
  AND U45878 ( .A(n26234), .B(n26233), .Z(n38175) );
  AND U45879 ( .A(n26236), .B(n26235), .Z(n38169) );
  AND U45880 ( .A(n26238), .B(n26237), .Z(n38163) );
  AND U45881 ( .A(n26240), .B(n26239), .Z(n38157) );
  NANDN U45882 ( .A(x[3304]), .B(y[3304]), .Z(n55541) );
  AND U45883 ( .A(n55541), .B(n26241), .Z(n38151) );
  AND U45884 ( .A(n26242), .B(n55540), .Z(n38145) );
  NANDN U45885 ( .A(x[3300]), .B(y[3300]), .Z(n26244) );
  AND U45886 ( .A(n26244), .B(n26243), .Z(n38139) );
  AND U45887 ( .A(n26246), .B(n26245), .Z(n38133) );
  AND U45888 ( .A(n26248), .B(n26247), .Z(n38127) );
  AND U45889 ( .A(n26250), .B(n26249), .Z(n38121) );
  AND U45890 ( .A(n26252), .B(n26251), .Z(n38115) );
  AND U45891 ( .A(n26254), .B(n26253), .Z(n38109) );
  NANDN U45892 ( .A(x[3288]), .B(y[3288]), .Z(n26256) );
  AND U45893 ( .A(n26256), .B(n26255), .Z(n38103) );
  AND U45894 ( .A(n26258), .B(n26257), .Z(n38097) );
  NANDN U45895 ( .A(x[3284]), .B(y[3284]), .Z(n26260) );
  AND U45896 ( .A(n26260), .B(n26259), .Z(n38091) );
  NANDN U45897 ( .A(x[3282]), .B(y[3282]), .Z(n26262) );
  AND U45898 ( .A(n26262), .B(n26261), .Z(n38085) );
  AND U45899 ( .A(n26264), .B(n26263), .Z(n38079) );
  AND U45900 ( .A(n26266), .B(n26265), .Z(n38073) );
  AND U45901 ( .A(n26268), .B(n26267), .Z(n38067) );
  AND U45902 ( .A(n26270), .B(n26269), .Z(n38061) );
  AND U45903 ( .A(n26272), .B(n26271), .Z(n38051) );
  NAND U45904 ( .A(n26274), .B(n26273), .Z(n38049) );
  AND U45905 ( .A(n26276), .B(n26275), .Z(n38047) );
  NANDN U45906 ( .A(x[3268]), .B(y[3268]), .Z(n51929) );
  AND U45907 ( .A(n51929), .B(n26277), .Z(n38045) );
  NAND U45908 ( .A(n26279), .B(n26278), .Z(n38043) );
  AND U45909 ( .A(n26280), .B(n51928), .Z(n38041) );
  AND U45910 ( .A(n26282), .B(n26281), .Z(n38035) );
  AND U45911 ( .A(n26284), .B(n26283), .Z(n38029) );
  AND U45912 ( .A(n26286), .B(n26285), .Z(n38023) );
  AND U45913 ( .A(n26288), .B(n26287), .Z(n38017) );
  AND U45914 ( .A(n26290), .B(n26289), .Z(n38011) );
  NANDN U45915 ( .A(x[3254]), .B(y[3254]), .Z(n26292) );
  AND U45916 ( .A(n26292), .B(n26291), .Z(n38005) );
  NAND U45917 ( .A(n26294), .B(n26293), .Z(n37995) );
  NAND U45918 ( .A(n26296), .B(n26295), .Z(n37989) );
  NAND U45919 ( .A(n26298), .B(n26297), .Z(n37983) );
  AND U45920 ( .A(n26300), .B(n26299), .Z(n37981) );
  NAND U45921 ( .A(n26302), .B(n26301), .Z(n37979) );
  AND U45922 ( .A(n26304), .B(n26303), .Z(n37973) );
  AND U45923 ( .A(n26306), .B(n26305), .Z(n37967) );
  NAND U45924 ( .A(n26308), .B(n26307), .Z(n37957) );
  NAND U45925 ( .A(n26310), .B(n26309), .Z(n37951) );
  NAND U45926 ( .A(n26312), .B(n26311), .Z(n37945) );
  ANDN U45927 ( .B(y[3232]), .A(x[3232]), .Z(n55480) );
  AND U45928 ( .A(n26314), .B(n26313), .Z(n37936) );
  AND U45929 ( .A(n55479), .B(n26315), .Z(n37934) );
  NAND U45930 ( .A(n26317), .B(n26316), .Z(n37932) );
  NANDN U45931 ( .A(x[3228]), .B(y[3228]), .Z(n55473) );
  AND U45932 ( .A(n26318), .B(n55473), .Z(n37930) );
  AND U45933 ( .A(n26319), .B(n55472), .Z(n37924) );
  AND U45934 ( .A(n26321), .B(n26320), .Z(n37918) );
  AND U45935 ( .A(n26323), .B(n26322), .Z(n37912) );
  ANDN U45936 ( .B(y[3220]), .A(x[3220]), .Z(n26325) );
  NOR U45937 ( .A(n26325), .B(n26324), .Z(n37906) );
  AND U45938 ( .A(n26327), .B(n26326), .Z(n37900) );
  NANDN U45939 ( .A(x[3216]), .B(y[3216]), .Z(n26329) );
  AND U45940 ( .A(n26329), .B(n26328), .Z(n37894) );
  NANDN U45941 ( .A(x[3214]), .B(y[3214]), .Z(n26331) );
  AND U45942 ( .A(n26331), .B(n26330), .Z(n37888) );
  NANDN U45943 ( .A(x[3212]), .B(y[3212]), .Z(n26333) );
  AND U45944 ( .A(n26333), .B(n26332), .Z(n37882) );
  AND U45945 ( .A(n26335), .B(n26334), .Z(n37876) );
  AND U45946 ( .A(n26337), .B(n26336), .Z(n37870) );
  AND U45947 ( .A(n26339), .B(n26338), .Z(n37864) );
  AND U45948 ( .A(n26341), .B(n26340), .Z(n37858) );
  AND U45949 ( .A(n26343), .B(n26342), .Z(n37852) );
  NANDN U45950 ( .A(x[3200]), .B(y[3200]), .Z(n51951) );
  AND U45951 ( .A(n51951), .B(n26344), .Z(n37846) );
  IV U45952 ( .A(n26345), .Z(n51950) );
  AND U45953 ( .A(n26346), .B(n51950), .Z(n37840) );
  NAND U45954 ( .A(n26348), .B(n26347), .Z(n37838) );
  NAND U45955 ( .A(n26350), .B(n26349), .Z(n37832) );
  AND U45956 ( .A(n26352), .B(n26351), .Z(n37823) );
  NAND U45957 ( .A(n26353), .B(n51955), .Z(n37821) );
  AND U45958 ( .A(n26355), .B(n26354), .Z(n37816) );
  IV U45959 ( .A(n26356), .Z(n51956) );
  NAND U45960 ( .A(n51956), .B(n26357), .Z(n37814) );
  AND U45961 ( .A(n26359), .B(n26358), .Z(n37812) );
  AND U45962 ( .A(n26361), .B(n26360), .Z(n37806) );
  AND U45963 ( .A(n26363), .B(n26362), .Z(n37796) );
  NAND U45964 ( .A(n26365), .B(n26364), .Z(n37794) );
  AND U45965 ( .A(n26367), .B(n26366), .Z(n37792) );
  AND U45966 ( .A(n26369), .B(n26368), .Z(n37790) );
  AND U45967 ( .A(n26371), .B(n26370), .Z(n37784) );
  NANDN U45968 ( .A(x[3176]), .B(y[3176]), .Z(n26373) );
  NAND U45969 ( .A(n26373), .B(n26372), .Z(n37782) );
  AND U45970 ( .A(n26375), .B(n26374), .Z(n37780) );
  AND U45971 ( .A(n26377), .B(n26376), .Z(n37774) );
  AND U45972 ( .A(n26379), .B(n26378), .Z(n37768) );
  NAND U45973 ( .A(n26381), .B(n26380), .Z(n37758) );
  NAND U45974 ( .A(n26383), .B(n26382), .Z(n37752) );
  ANDN U45975 ( .B(y[3164]), .A(x[3164]), .Z(n55420) );
  AND U45976 ( .A(n26385), .B(n26384), .Z(n37743) );
  NANDN U45977 ( .A(x[3162]), .B(y[3162]), .Z(n51961) );
  AND U45978 ( .A(n55419), .B(n51961), .Z(n37741) );
  NAND U45979 ( .A(n26387), .B(n26386), .Z(n37739) );
  IV U45980 ( .A(n26388), .Z(n55416) );
  AND U45981 ( .A(n26389), .B(n55416), .Z(n37737) );
  NANDN U45982 ( .A(x[3158]), .B(y[3158]), .Z(n51963) );
  AND U45983 ( .A(n51963), .B(n26390), .Z(n37731) );
  AND U45984 ( .A(n26391), .B(n51962), .Z(n37725) );
  AND U45985 ( .A(n26393), .B(n26392), .Z(n37719) );
  AND U45986 ( .A(n26395), .B(n26394), .Z(n37705) );
  NANDN U45987 ( .A(x[3148]), .B(y[3148]), .Z(n26397) );
  AND U45988 ( .A(n26397), .B(n26396), .Z(n37699) );
  AND U45989 ( .A(n26399), .B(n26398), .Z(n37693) );
  AND U45990 ( .A(n26401), .B(n26400), .Z(n37687) );
  NANDN U45991 ( .A(x[3142]), .B(y[3142]), .Z(n26403) );
  AND U45992 ( .A(n26403), .B(n26402), .Z(n37681) );
  AND U45993 ( .A(n26405), .B(n26404), .Z(n37679) );
  NANDN U45994 ( .A(x[3140]), .B(y[3140]), .Z(n55394) );
  AND U45995 ( .A(n55394), .B(n26406), .Z(n37677) );
  NAND U45996 ( .A(n26408), .B(n26407), .Z(n37675) );
  AND U45997 ( .A(n26409), .B(n55393), .Z(n37673) );
  NANDN U45998 ( .A(x[3136]), .B(y[3136]), .Z(n26411) );
  AND U45999 ( .A(n26411), .B(n26410), .Z(n37667) );
  NANDN U46000 ( .A(x[3134]), .B(y[3134]), .Z(n26413) );
  AND U46001 ( .A(n26413), .B(n26412), .Z(n37661) );
  AND U46002 ( .A(n26415), .B(n26414), .Z(n37655) );
  AND U46003 ( .A(n26417), .B(n26416), .Z(n37649) );
  NAND U46004 ( .A(n26419), .B(n26418), .Z(n37639) );
  NAND U46005 ( .A(n26421), .B(n26420), .Z(n37633) );
  NAND U46006 ( .A(n26423), .B(n26422), .Z(n37627) );
  AND U46007 ( .A(n26425), .B(n26424), .Z(n37625) );
  AND U46008 ( .A(n26427), .B(n26426), .Z(n37623) );
  NAND U46009 ( .A(n26429), .B(n26428), .Z(n37621) );
  ANDN U46010 ( .B(n26431), .A(n26430), .Z(n37619) );
  NAND U46011 ( .A(n26433), .B(n26432), .Z(n37605) );
  AND U46012 ( .A(n26435), .B(n26434), .Z(n37603) );
  NAND U46013 ( .A(n26437), .B(n26436), .Z(n37601) );
  AND U46014 ( .A(n26439), .B(n26438), .Z(n37599) );
  NAND U46015 ( .A(n26441), .B(n26440), .Z(n37593) );
  NAND U46016 ( .A(n26443), .B(n26442), .Z(n37587) );
  NAND U46017 ( .A(n26445), .B(n26444), .Z(n37581) );
  AND U46018 ( .A(n26447), .B(n26446), .Z(n37579) );
  NAND U46019 ( .A(n26449), .B(n26448), .Z(n37577) );
  AND U46020 ( .A(n26451), .B(n26450), .Z(n37567) );
  AND U46021 ( .A(n26453), .B(n26452), .Z(n37565) );
  NAND U46022 ( .A(n26455), .B(n26454), .Z(n37563) );
  AND U46023 ( .A(n26457), .B(n26456), .Z(n37561) );
  NAND U46024 ( .A(n26459), .B(n26458), .Z(n37551) );
  NAND U46025 ( .A(n26461), .B(n26460), .Z(n37545) );
  NAND U46026 ( .A(n26463), .B(n26462), .Z(n37539) );
  NANDN U46027 ( .A(x[3088]), .B(y[3088]), .Z(n55320) );
  NAND U46028 ( .A(n55320), .B(n26464), .Z(n37533) );
  AND U46029 ( .A(n26465), .B(n55319), .Z(n37527) );
  AND U46030 ( .A(n26467), .B(n26466), .Z(n37521) );
  AND U46031 ( .A(n26469), .B(n26468), .Z(n37515) );
  NANDN U46032 ( .A(x[3080]), .B(y[3080]), .Z(n51967) );
  AND U46033 ( .A(n26470), .B(n51967), .Z(n37509) );
  NAND U46034 ( .A(n26472), .B(n26471), .Z(n37507) );
  AND U46035 ( .A(n26474), .B(n26473), .Z(n37502) );
  NAND U46036 ( .A(n26475), .B(n55306), .Z(n37493) );
  NAND U46037 ( .A(n26477), .B(n26476), .Z(n37487) );
  NAND U46038 ( .A(n26479), .B(n26478), .Z(n37481) );
  NANDN U46039 ( .A(x[3068]), .B(y[3068]), .Z(n26481) );
  NAND U46040 ( .A(n26481), .B(n26480), .Z(n37475) );
  AND U46041 ( .A(n26483), .B(n26482), .Z(n37473) );
  NANDN U46042 ( .A(x[3066]), .B(y[3066]), .Z(n26484) );
  AND U46043 ( .A(n26485), .B(n26484), .Z(n37471) );
  NAND U46044 ( .A(n26487), .B(n26486), .Z(n37469) );
  NANDN U46045 ( .A(x[3064]), .B(y[3064]), .Z(n26489) );
  AND U46046 ( .A(n26489), .B(n26488), .Z(n37467) );
  NANDN U46047 ( .A(x[3062]), .B(y[3062]), .Z(n26491) );
  AND U46048 ( .A(n26491), .B(n26490), .Z(n37461) );
  NANDN U46049 ( .A(x[3060]), .B(y[3060]), .Z(n26493) );
  AND U46050 ( .A(n26493), .B(n26492), .Z(n37455) );
  AND U46051 ( .A(n26495), .B(n26494), .Z(n37449) );
  AND U46052 ( .A(n26497), .B(n26496), .Z(n37443) );
  AND U46053 ( .A(n26499), .B(n26498), .Z(n37437) );
  NAND U46054 ( .A(n26501), .B(n26500), .Z(n37435) );
  AND U46055 ( .A(n26503), .B(n26502), .Z(n37429) );
  NAND U46056 ( .A(n26505), .B(n26504), .Z(n37424) );
  AND U46057 ( .A(n26506), .B(n55284), .Z(n37422) );
  NAND U46058 ( .A(n26508), .B(n26507), .Z(n37420) );
  XOR U46059 ( .A(x[3046]), .B(y[3046]), .Z(n37413) );
  AND U46060 ( .A(n26509), .B(n55272), .Z(n37403) );
  AND U46061 ( .A(n55273), .B(n26510), .Z(n37401) );
  NAND U46062 ( .A(n26512), .B(n26511), .Z(n37399) );
  AND U46063 ( .A(n26514), .B(n26513), .Z(n37390) );
  AND U46064 ( .A(n26516), .B(n26515), .Z(n37384) );
  AND U46065 ( .A(n26518), .B(n26517), .Z(n37378) );
  NANDN U46066 ( .A(x[3028]), .B(y[3028]), .Z(n26520) );
  AND U46067 ( .A(n26520), .B(n26519), .Z(n37364) );
  AND U46068 ( .A(n26522), .B(n26521), .Z(n37358) );
  AND U46069 ( .A(n26524), .B(n26523), .Z(n37352) );
  NAND U46070 ( .A(n26526), .B(n26525), .Z(n37342) );
  NAND U46071 ( .A(n26528), .B(n26527), .Z(n37336) );
  NANDN U46072 ( .A(x[3014]), .B(y[3014]), .Z(n51978) );
  NAND U46073 ( .A(n51978), .B(n26529), .Z(n37318) );
  AND U46074 ( .A(n26531), .B(n26530), .Z(n37305) );
  NANDN U46075 ( .A(x[3008]), .B(y[3008]), .Z(n55217) );
  AND U46076 ( .A(n26532), .B(n55217), .Z(n37299) );
  AND U46077 ( .A(n26533), .B(n55216), .Z(n37293) );
  AND U46078 ( .A(n26535), .B(n26534), .Z(n37287) );
  AND U46079 ( .A(n26537), .B(n26536), .Z(n37281) );
  AND U46080 ( .A(n26539), .B(n26538), .Z(n37275) );
  AND U46081 ( .A(n26541), .B(n26540), .Z(n37269) );
  NANDN U46082 ( .A(x[2996]), .B(y[2996]), .Z(n26543) );
  AND U46083 ( .A(n26543), .B(n26542), .Z(n37263) );
  NANDN U46084 ( .A(x[2994]), .B(y[2994]), .Z(n26545) );
  AND U46085 ( .A(n26545), .B(n26544), .Z(n37257) );
  AND U46086 ( .A(n26547), .B(n26546), .Z(n37251) );
  AND U46087 ( .A(n26549), .B(n26548), .Z(n37245) );
  AND U46088 ( .A(n26551), .B(n26550), .Z(n37235) );
  AND U46089 ( .A(n26553), .B(n26552), .Z(n37229) );
  NAND U46090 ( .A(n26555), .B(n26554), .Z(n37227) );
  AND U46091 ( .A(n26557), .B(n26556), .Z(n37225) );
  AND U46092 ( .A(n26559), .B(n26558), .Z(n37223) );
  NAND U46093 ( .A(n26561), .B(n26560), .Z(n37221) );
  NANDN U46094 ( .A(x[2980]), .B(y[2980]), .Z(n26563) );
  AND U46095 ( .A(n26563), .B(n26562), .Z(n37219) );
  AND U46096 ( .A(n26565), .B(n26564), .Z(n37217) );
  NANDN U46097 ( .A(x[2978]), .B(y[2978]), .Z(n26567) );
  AND U46098 ( .A(n26567), .B(n26566), .Z(n37215) );
  NAND U46099 ( .A(n26569), .B(n26568), .Z(n37213) );
  AND U46100 ( .A(n26571), .B(n26570), .Z(n37211) );
  AND U46101 ( .A(n26573), .B(n26572), .Z(n37205) );
  AND U46102 ( .A(n26575), .B(n26574), .Z(n37199) );
  NANDN U46103 ( .A(x[2970]), .B(y[2970]), .Z(n55176) );
  AND U46104 ( .A(n55176), .B(n26576), .Z(n37193) );
  IV U46105 ( .A(n26577), .Z(n55175) );
  AND U46106 ( .A(n26578), .B(n55175), .Z(n37187) );
  AND U46107 ( .A(n26580), .B(n26579), .Z(n37181) );
  NANDN U46108 ( .A(x[2964]), .B(y[2964]), .Z(n55172) );
  AND U46109 ( .A(n55172), .B(n26581), .Z(n37175) );
  NAND U46110 ( .A(n26583), .B(n26582), .Z(n37166) );
  NAND U46111 ( .A(n26585), .B(n26584), .Z(n37160) );
  NAND U46112 ( .A(n26587), .B(n26586), .Z(n37154) );
  AND U46113 ( .A(n26589), .B(n26588), .Z(n37152) );
  AND U46114 ( .A(n26591), .B(n26590), .Z(n37150) );
  NAND U46115 ( .A(n55161), .B(n26592), .Z(n37148) );
  AND U46116 ( .A(n26594), .B(n26593), .Z(n37146) );
  AND U46117 ( .A(n26596), .B(n26595), .Z(n37142) );
  NAND U46118 ( .A(n26598), .B(n26597), .Z(n37140) );
  NANDN U46119 ( .A(x[2948]), .B(y[2948]), .Z(n26600) );
  NAND U46120 ( .A(n26600), .B(n26599), .Z(n37134) );
  NAND U46121 ( .A(n26602), .B(n26601), .Z(n37128) );
  NAND U46122 ( .A(n26604), .B(n26603), .Z(n37122) );
  AND U46123 ( .A(n26606), .B(n26605), .Z(n37120) );
  NAND U46124 ( .A(n26608), .B(n26607), .Z(n37118) );
  AND U46125 ( .A(n26610), .B(n26609), .Z(n37112) );
  NANDN U46126 ( .A(x[2938]), .B(y[2938]), .Z(n55146) );
  AND U46127 ( .A(n26611), .B(n55146), .Z(n37106) );
  AND U46128 ( .A(n26612), .B(n55145), .Z(n37100) );
  AND U46129 ( .A(n26614), .B(n26613), .Z(n37094) );
  AND U46130 ( .A(n26616), .B(n26615), .Z(n37088) );
  AND U46131 ( .A(n26618), .B(n26617), .Z(n37082) );
  AND U46132 ( .A(n26620), .B(n26619), .Z(n37076) );
  AND U46133 ( .A(n26622), .B(n26621), .Z(n37070) );
  AND U46134 ( .A(n26624), .B(n26623), .Z(n37064) );
  AND U46135 ( .A(n26626), .B(n26625), .Z(n37058) );
  AND U46136 ( .A(n26628), .B(n26627), .Z(n37052) );
  AND U46137 ( .A(n26630), .B(n26629), .Z(n37046) );
  AND U46138 ( .A(n26632), .B(n26631), .Z(n37040) );
  NANDN U46139 ( .A(x[2914]), .B(y[2914]), .Z(n26634) );
  AND U46140 ( .A(n26634), .B(n26633), .Z(n37034) );
  NAND U46141 ( .A(n26636), .B(n26635), .Z(n37032) );
  AND U46142 ( .A(n26638), .B(n26637), .Z(n37026) );
  AND U46143 ( .A(n26640), .B(n26639), .Z(n37020) );
  NANDN U46144 ( .A(x[2908]), .B(y[2908]), .Z(n26642) );
  AND U46145 ( .A(n26642), .B(n26641), .Z(n37018) );
  NAND U46146 ( .A(n26644), .B(n26643), .Z(n37016) );
  AND U46147 ( .A(n26646), .B(n26645), .Z(n37006) );
  AND U46148 ( .A(n26648), .B(n26647), .Z(n37004) );
  NAND U46149 ( .A(n26650), .B(n26649), .Z(n37002) );
  AND U46150 ( .A(n26652), .B(n26651), .Z(n37000) );
  AND U46151 ( .A(n26654), .B(n26653), .Z(n36994) );
  AND U46152 ( .A(n26656), .B(n26655), .Z(n36988) );
  AND U46153 ( .A(n26658), .B(n26657), .Z(n36982) );
  AND U46154 ( .A(n26660), .B(n26659), .Z(n36976) );
  AND U46155 ( .A(n26662), .B(n26661), .Z(n36970) );
  NAND U46156 ( .A(n55096), .B(n26663), .Z(n36968) );
  NAND U46157 ( .A(n26664), .B(n55094), .Z(n36962) );
  AND U46158 ( .A(n26665), .B(n51994), .Z(n36960) );
  AND U46159 ( .A(n26667), .B(n26666), .Z(n36958) );
  NAND U46160 ( .A(n26669), .B(n26668), .Z(n36952) );
  NAND U46161 ( .A(n26671), .B(n26670), .Z(n36946) );
  NAND U46162 ( .A(n26673), .B(n26672), .Z(n36940) );
  NAND U46163 ( .A(n26675), .B(n26674), .Z(n36934) );
  AND U46164 ( .A(n26677), .B(n26676), .Z(n36932) );
  NAND U46165 ( .A(n26679), .B(n26678), .Z(n36930) );
  AND U46166 ( .A(n26681), .B(n26680), .Z(n36924) );
  NAND U46167 ( .A(n26683), .B(n26682), .Z(n36922) );
  AND U46168 ( .A(n26685), .B(n26684), .Z(n36920) );
  AND U46169 ( .A(n26687), .B(n26686), .Z(n36914) );
  AND U46170 ( .A(n26689), .B(n26688), .Z(n36908) );
  AND U46171 ( .A(n26691), .B(n26690), .Z(n36902) );
  AND U46172 ( .A(n26693), .B(n26692), .Z(n36896) );
  NAND U46173 ( .A(n26695), .B(n26694), .Z(n36886) );
  NAND U46174 ( .A(n26697), .B(n26696), .Z(n36880) );
  AND U46175 ( .A(n26699), .B(n26698), .Z(n36866) );
  AND U46176 ( .A(n26701), .B(n26700), .Z(n36860) );
  AND U46177 ( .A(n26703), .B(n26702), .Z(n36854) );
  NANDN U46178 ( .A(x[2846]), .B(y[2846]), .Z(n26705) );
  NAND U46179 ( .A(n26705), .B(n26704), .Z(n36840) );
  AND U46180 ( .A(n26707), .B(n26706), .Z(n36838) );
  AND U46181 ( .A(n26709), .B(n26708), .Z(n36832) );
  AND U46182 ( .A(n26711), .B(n26710), .Z(n36826) );
  AND U46183 ( .A(n26713), .B(n26712), .Z(n36824) );
  NAND U46184 ( .A(n26715), .B(n26714), .Z(n36822) );
  AND U46185 ( .A(n26717), .B(n26716), .Z(n36816) );
  NANDN U46186 ( .A(x[2836]), .B(y[2836]), .Z(n55053) );
  NAND U46187 ( .A(n55053), .B(n26718), .Z(n36814) );
  AND U46188 ( .A(n26720), .B(n26719), .Z(n36812) );
  AND U46189 ( .A(n26722), .B(n26721), .Z(n36807) );
  AND U46190 ( .A(n26724), .B(n26723), .Z(n36801) );
  AND U46191 ( .A(n26726), .B(n26725), .Z(n36795) );
  NAND U46192 ( .A(n26728), .B(n26727), .Z(n36781) );
  AND U46193 ( .A(n26730), .B(n26729), .Z(n36779) );
  NANDN U46194 ( .A(x[2822]), .B(y[2822]), .Z(n52012) );
  NAND U46195 ( .A(n52012), .B(n26731), .Z(n36773) );
  IV U46196 ( .A(n26732), .Z(n55037) );
  NAND U46197 ( .A(n55037), .B(n26733), .Z(n36767) );
  AND U46198 ( .A(n26735), .B(n26734), .Z(n36765) );
  NANDN U46199 ( .A(x[2818]), .B(y[2818]), .Z(n55034) );
  AND U46200 ( .A(n55034), .B(n26736), .Z(n36763) );
  NAND U46201 ( .A(n26738), .B(n26737), .Z(n36761) );
  NANDN U46202 ( .A(x[2816]), .B(y[2816]), .Z(n55029) );
  IV U46203 ( .A(n26739), .Z(n55033) );
  AND U46204 ( .A(n55029), .B(n55033), .Z(n36759) );
  AND U46205 ( .A(n26740), .B(n55030), .Z(n36753) );
  AND U46206 ( .A(n26742), .B(n26741), .Z(n36747) );
  AND U46207 ( .A(n26744), .B(n26743), .Z(n36741) );
  AND U46208 ( .A(n26746), .B(n26745), .Z(n36735) );
  AND U46209 ( .A(n26748), .B(n26747), .Z(n36729) );
  NAND U46210 ( .A(n26750), .B(n26749), .Z(n36719) );
  NAND U46211 ( .A(n26752), .B(n26751), .Z(n36713) );
  NAND U46212 ( .A(n26754), .B(n26753), .Z(n36707) );
  AND U46213 ( .A(n26756), .B(n26755), .Z(n36705) );
  NAND U46214 ( .A(n26758), .B(n26757), .Z(n36694) );
  ANDN U46215 ( .B(y[2792]), .A(x[2792]), .Z(n36686) );
  AND U46216 ( .A(n26760), .B(n26759), .Z(n36684) );
  ANDN U46217 ( .B(y[2790]), .A(x[2790]), .Z(n52015) );
  NOR U46218 ( .A(n52015), .B(n26761), .Z(n36682) );
  IV U46219 ( .A(n26762), .Z(n55003) );
  AND U46220 ( .A(n26763), .B(n55003), .Z(n36676) );
  AND U46221 ( .A(n26765), .B(n26764), .Z(n36662) );
  AND U46222 ( .A(n26767), .B(n26766), .Z(n36652) );
  AND U46223 ( .A(n26769), .B(n26768), .Z(n36646) );
  AND U46224 ( .A(n26771), .B(n26770), .Z(n36641) );
  AND U46225 ( .A(n26773), .B(n26772), .Z(n36637) );
  NAND U46226 ( .A(n26774), .B(n54978), .Z(n36635) );
  AND U46227 ( .A(n26776), .B(n26775), .Z(n36633) );
  AND U46228 ( .A(n26778), .B(n26777), .Z(n36627) );
  NANDN U46229 ( .A(x[2768]), .B(y[2768]), .Z(n54960) );
  NAND U46230 ( .A(n54960), .B(n26779), .Z(n36617) );
  NAND U46231 ( .A(n26780), .B(n54959), .Z(n36611) );
  ANDN U46232 ( .B(y[2764]), .A(x[2764]), .Z(n36605) );
  AND U46233 ( .A(n26782), .B(n26781), .Z(n36597) );
  NANDN U46234 ( .A(x[2760]), .B(y[2760]), .Z(n26784) );
  AND U46235 ( .A(n26784), .B(n26783), .Z(n36591) );
  NAND U46236 ( .A(n26786), .B(n26785), .Z(n36581) );
  NAND U46237 ( .A(n26788), .B(n26787), .Z(n36575) );
  NAND U46238 ( .A(n26790), .B(n26789), .Z(n36569) );
  NAND U46239 ( .A(n26792), .B(n26791), .Z(n36563) );
  AND U46240 ( .A(n26793), .B(n52019), .Z(n36554) );
  NAND U46241 ( .A(n26795), .B(n26794), .Z(n36552) );
  AND U46242 ( .A(n26797), .B(n26796), .Z(n36550) );
  AND U46243 ( .A(n26799), .B(n26798), .Z(n36544) );
  AND U46244 ( .A(n54933), .B(n26800), .Z(n36533) );
  NAND U46245 ( .A(n26802), .B(n26801), .Z(n36531) );
  IV U46246 ( .A(n26803), .Z(n54929) );
  AND U46247 ( .A(n26804), .B(n54929), .Z(n36525) );
  NAND U46248 ( .A(n26806), .B(n26805), .Z(n54928) );
  IV U46249 ( .A(n26807), .Z(n54927) );
  AND U46250 ( .A(n26808), .B(n54927), .Z(n36522) );
  AND U46251 ( .A(n26810), .B(n26809), .Z(n36517) );
  AND U46252 ( .A(n26812), .B(n26811), .Z(n36511) );
  AND U46253 ( .A(n26814), .B(n26813), .Z(n36505) );
  AND U46254 ( .A(n26816), .B(n26815), .Z(n36499) );
  AND U46255 ( .A(n26818), .B(n26817), .Z(n36493) );
  AND U46256 ( .A(n26820), .B(n26819), .Z(n36487) );
  AND U46257 ( .A(n26822), .B(n26821), .Z(n36481) );
  NAND U46258 ( .A(n26824), .B(n26823), .Z(n36471) );
  NANDN U46259 ( .A(x[2716]), .B(y[2716]), .Z(n54884) );
  NAND U46260 ( .A(n54884), .B(n26825), .Z(n36465) );
  ANDN U46261 ( .B(y[2714]), .A(x[2714]), .Z(n54881) );
  AND U46262 ( .A(n26827), .B(n26826), .Z(n36457) );
  IV U46263 ( .A(n26828), .Z(n54880) );
  AND U46264 ( .A(n26829), .B(n54880), .Z(n36455) );
  NAND U46265 ( .A(n26831), .B(n26830), .Z(n36453) );
  NAND U46266 ( .A(n26833), .B(n26832), .Z(n36441) );
  AND U46267 ( .A(n26835), .B(n26834), .Z(n36431) );
  NAND U46268 ( .A(n26837), .B(n26836), .Z(n36429) );
  AND U46269 ( .A(n26839), .B(n26838), .Z(n36424) );
  AND U46270 ( .A(n26841), .B(n26840), .Z(n36419) );
  AND U46271 ( .A(n26843), .B(n26842), .Z(n36413) );
  AND U46272 ( .A(n26845), .B(n26844), .Z(n36403) );
  NAND U46273 ( .A(n26847), .B(n26846), .Z(n36401) );
  NANDN U46274 ( .A(x[2692]), .B(y[2692]), .Z(n26849) );
  AND U46275 ( .A(n26849), .B(n26848), .Z(n36399) );
  AND U46276 ( .A(n26851), .B(n26850), .Z(n36397) );
  NAND U46277 ( .A(n26853), .B(n26852), .Z(n36395) );
  AND U46278 ( .A(n26855), .B(n26854), .Z(n36393) );
  AND U46279 ( .A(n26857), .B(n26856), .Z(n36387) );
  AND U46280 ( .A(n26859), .B(n26858), .Z(n36381) );
  AND U46281 ( .A(n26861), .B(n26860), .Z(n36375) );
  AND U46282 ( .A(n26863), .B(n26862), .Z(n36369) );
  AND U46283 ( .A(n26865), .B(n26864), .Z(n36363) );
  AND U46284 ( .A(n26867), .B(n26866), .Z(n36357) );
  NAND U46285 ( .A(n26869), .B(n26868), .Z(n36347) );
  NANDN U46286 ( .A(x[2672]), .B(y[2672]), .Z(n54838) );
  NAND U46287 ( .A(n54838), .B(n26870), .Z(n36341) );
  NANDN U46288 ( .A(x[2668]), .B(y[2668]), .Z(n52031) );
  AND U46289 ( .A(n52031), .B(n26871), .Z(n36328) );
  IV U46290 ( .A(n26872), .Z(n52030) );
  AND U46291 ( .A(n26873), .B(n52030), .Z(n36322) );
  AND U46292 ( .A(n26875), .B(n26874), .Z(n36316) );
  NANDN U46293 ( .A(x[2662]), .B(y[2662]), .Z(n26877) );
  AND U46294 ( .A(n26877), .B(n26876), .Z(n36310) );
  AND U46295 ( .A(n26879), .B(n26878), .Z(n36304) );
  AND U46296 ( .A(n26881), .B(n26880), .Z(n36298) );
  AND U46297 ( .A(n26883), .B(n26882), .Z(n36288) );
  NAND U46298 ( .A(n26885), .B(n26884), .Z(n36286) );
  AND U46299 ( .A(n26887), .B(n26886), .Z(n36284) );
  NANDN U46300 ( .A(x[2652]), .B(y[2652]), .Z(n26888) );
  AND U46301 ( .A(n26889), .B(n26888), .Z(n36282) );
  NAND U46302 ( .A(n26891), .B(n26890), .Z(n36280) );
  NANDN U46303 ( .A(x[2650]), .B(y[2650]), .Z(n26893) );
  AND U46304 ( .A(n26893), .B(n26892), .Z(n36278) );
  AND U46305 ( .A(n26895), .B(n26894), .Z(n36272) );
  NAND U46306 ( .A(n26897), .B(n26896), .Z(n36270) );
  AND U46307 ( .A(n26899), .B(n26898), .Z(n36264) );
  ANDN U46308 ( .B(y[2644]), .A(x[2644]), .Z(n36262) );
  NAND U46309 ( .A(n26901), .B(n26900), .Z(n36258) );
  NAND U46310 ( .A(n26903), .B(n26902), .Z(n36252) );
  AND U46311 ( .A(n26905), .B(n26904), .Z(n36250) );
  ANDN U46312 ( .B(y[2638]), .A(x[2638]), .Z(n36244) );
  AND U46313 ( .A(n26907), .B(n26906), .Z(n36236) );
  NAND U46314 ( .A(n26909), .B(n26908), .Z(n36234) );
  AND U46315 ( .A(n26911), .B(n26910), .Z(n36232) );
  NANDN U46316 ( .A(x[2632]), .B(y[2632]), .Z(n52047) );
  XOR U46317 ( .A(x[2630]), .B(y[2630]), .Z(n26912) );
  NOR U46318 ( .A(n26913), .B(n26912), .Z(n36217) );
  AND U46319 ( .A(n26915), .B(n26914), .Z(n36212) );
  NAND U46320 ( .A(n26917), .B(n26916), .Z(n36202) );
  AND U46321 ( .A(n26919), .B(n26918), .Z(n36200) );
  NAND U46322 ( .A(n26921), .B(n26920), .Z(n36198) );
  AND U46323 ( .A(n26923), .B(n26922), .Z(n36196) );
  ANDN U46324 ( .B(y[2620]), .A(x[2620]), .Z(n36192) );
  AND U46325 ( .A(n26925), .B(n26924), .Z(n36190) );
  ANDN U46326 ( .B(y[2618]), .A(x[2618]), .Z(n52050) );
  NANDN U46327 ( .A(x[2616]), .B(y[2616]), .Z(n54789) );
  AND U46328 ( .A(n54792), .B(n54789), .Z(n36181) );
  NANDN U46329 ( .A(x[2612]), .B(y[2612]), .Z(n26927) );
  AND U46330 ( .A(n26927), .B(n26926), .Z(n36168) );
  NANDN U46331 ( .A(x[2610]), .B(y[2610]), .Z(n26929) );
  AND U46332 ( .A(n26929), .B(n26928), .Z(n36162) );
  NANDN U46333 ( .A(x[2608]), .B(y[2608]), .Z(n26931) );
  AND U46334 ( .A(n26931), .B(n26930), .Z(n36156) );
  AND U46335 ( .A(n26933), .B(n26932), .Z(n36142) );
  AND U46336 ( .A(n26935), .B(n26934), .Z(n36136) );
  AND U46337 ( .A(n26937), .B(n26936), .Z(n36130) );
  AND U46338 ( .A(n26939), .B(n26938), .Z(n36124) );
  NANDN U46339 ( .A(x[2594]), .B(y[2594]), .Z(n26941) );
  AND U46340 ( .A(n26941), .B(n26940), .Z(n36110) );
  NANDN U46341 ( .A(x[2592]), .B(y[2592]), .Z(n36104) );
  AND U46342 ( .A(n26943), .B(n26942), .Z(n36100) );
  ANDN U46343 ( .B(y[2590]), .A(x[2590]), .Z(n26944) );
  NOR U46344 ( .A(n26945), .B(n26944), .Z(n36098) );
  NANDN U46345 ( .A(x[2588]), .B(y[2588]), .Z(n26947) );
  AND U46346 ( .A(n26947), .B(n26946), .Z(n36092) );
  NANDN U46347 ( .A(x[2586]), .B(y[2586]), .Z(n36086) );
  NAND U46348 ( .A(n26951), .B(n26950), .Z(n54754) );
  IV U46349 ( .A(n26954), .Z(n26956) );
  NAND U46350 ( .A(n26956), .B(n26955), .Z(n54752) );
  AND U46351 ( .A(n26958), .B(n26957), .Z(n54751) );
  ANDN U46352 ( .B(y[2574]), .A(x[2574]), .Z(n36054) );
  AND U46353 ( .A(n26960), .B(n26959), .Z(n36048) );
  NAND U46354 ( .A(n26962), .B(n26961), .Z(n36046) );
  AND U46355 ( .A(n26964), .B(n26963), .Z(n36044) );
  AND U46356 ( .A(n26966), .B(n26965), .Z(n36038) );
  NAND U46357 ( .A(n54739), .B(n26967), .Z(n36029) );
  AND U46358 ( .A(n26970), .B(n54730), .Z(n36009) );
  NANDN U46359 ( .A(x[2556]), .B(y[2556]), .Z(n26971) );
  AND U46360 ( .A(n26971), .B(n54728), .Z(n36004) );
  NANDN U46361 ( .A(x[2552]), .B(y[2552]), .Z(n26973) );
  AND U46362 ( .A(n26973), .B(n26972), .Z(n35990) );
  NAND U46363 ( .A(n26975), .B(n26974), .Z(n35988) );
  NOR U46364 ( .A(n26977), .B(n26976), .Z(n35960) );
  AND U46365 ( .A(n26979), .B(n26978), .Z(n35954) );
  ANDN U46366 ( .B(y[2538]), .A(x[2538]), .Z(n26980) );
  NOR U46367 ( .A(n26981), .B(n26980), .Z(n35944) );
  IV U46368 ( .A(n26982), .Z(n52061) );
  NAND U46369 ( .A(n26986), .B(n26985), .Z(n35939) );
  AND U46370 ( .A(n26987), .B(n54707), .Z(n35937) );
  AND U46371 ( .A(n26989), .B(n26988), .Z(n35931) );
  IV U46372 ( .A(n26990), .Z(n54701) );
  NAND U46373 ( .A(n54701), .B(n26991), .Z(n35922) );
  AND U46374 ( .A(n26993), .B(n26992), .Z(n52065) );
  NAND U46375 ( .A(n26995), .B(n26994), .Z(n35897) );
  NOR U46376 ( .A(n26997), .B(n26996), .Z(n35891) );
  IV U46377 ( .A(n26998), .Z(n26999) );
  AND U46378 ( .A(n27000), .B(n26999), .Z(n54690) );
  IV U46379 ( .A(n27003), .Z(n27004) );
  AND U46380 ( .A(n27005), .B(n27004), .Z(n54686) );
  IV U46381 ( .A(n27006), .Z(n27007) );
  AND U46382 ( .A(n27008), .B(n27007), .Z(n54685) );
  AND U46383 ( .A(n27009), .B(n54684), .Z(n35876) );
  ANDN U46384 ( .B(y[2510]), .A(x[2510]), .Z(n27010) );
  NOR U46385 ( .A(n54683), .B(n27010), .Z(n35874) );
  NANDN U46386 ( .A(x[2508]), .B(y[2508]), .Z(n27012) );
  AND U46387 ( .A(n27012), .B(n27011), .Z(n35868) );
  NOR U46388 ( .A(n27014), .B(n27013), .Z(n35858) );
  AND U46389 ( .A(n27016), .B(n27015), .Z(n35852) );
  AND U46390 ( .A(n27018), .B(n27017), .Z(n35846) );
  ANDN U46391 ( .B(y[2500]), .A(x[2500]), .Z(n35844) );
  NANDN U46392 ( .A(x[2498]), .B(y[2498]), .Z(n52071) );
  AND U46393 ( .A(n52071), .B(n27019), .Z(n35836) );
  NANDN U46394 ( .A(x[2496]), .B(y[2496]), .Z(n27021) );
  IV U46395 ( .A(n27020), .Z(n52070) );
  AND U46396 ( .A(n27021), .B(n52070), .Z(n35830) );
  AND U46397 ( .A(n27023), .B(n27022), .Z(n35816) );
  AND U46398 ( .A(n27025), .B(n27024), .Z(n35806) );
  AND U46399 ( .A(n27027), .B(n27026), .Z(n35796) );
  NAND U46400 ( .A(n27029), .B(n27028), .Z(n35794) );
  AND U46401 ( .A(n27031), .B(n27030), .Z(n35788) );
  NOR U46402 ( .A(n27033), .B(n27032), .Z(n35786) );
  AND U46403 ( .A(n27035), .B(n27034), .Z(n35780) );
  NAND U46404 ( .A(n52078), .B(n27036), .Z(n35770) );
  IV U46405 ( .A(n27037), .Z(n54651) );
  NANDN U46406 ( .A(x[2474]), .B(y[2474]), .Z(n35763) );
  AND U46407 ( .A(n27039), .B(n27038), .Z(n35760) );
  NAND U46408 ( .A(n27041), .B(n27040), .Z(n35758) );
  AND U46409 ( .A(n27043), .B(n27042), .Z(n35748) );
  NAND U46410 ( .A(n27045), .B(n27044), .Z(n35746) );
  NAND U46411 ( .A(n27047), .B(n27046), .Z(n35724) );
  AND U46412 ( .A(n27049), .B(n27048), .Z(n35722) );
  IV U46413 ( .A(n27050), .Z(n54633) );
  NAND U46414 ( .A(n54633), .B(n27051), .Z(n35720) );
  AND U46415 ( .A(n27052), .B(n54632), .Z(n35718) );
  NAND U46416 ( .A(n27056), .B(n27055), .Z(n54630) );
  IV U46417 ( .A(n27059), .Z(n27060) );
  AND U46418 ( .A(n27061), .B(n27060), .Z(n54627) );
  NAND U46419 ( .A(n27063), .B(n27062), .Z(n35703) );
  XOR U46420 ( .A(x[2448]), .B(y[2448]), .Z(n35688) );
  AND U46421 ( .A(n27065), .B(n27064), .Z(n35682) );
  IV U46422 ( .A(n27066), .Z(n54615) );
  NAND U46423 ( .A(n54615), .B(n27067), .Z(n35680) );
  AND U46424 ( .A(n27069), .B(n27068), .Z(n35678) );
  AND U46425 ( .A(n27071), .B(n27070), .Z(n35666) );
  AND U46426 ( .A(n54609), .B(n27072), .Z(n35661) );
  AND U46427 ( .A(n27074), .B(n27073), .Z(n54607) );
  IV U46428 ( .A(n27075), .Z(n54605) );
  AND U46429 ( .A(n27077), .B(n27076), .Z(n35647) );
  ANDN U46430 ( .B(y[2430]), .A(x[2430]), .Z(n35645) );
  AND U46431 ( .A(n54583), .B(n27078), .Z(n35602) );
  IV U46432 ( .A(n27079), .Z(n54582) );
  NOR U46433 ( .A(n54582), .B(n27080), .Z(n35600) );
  AND U46434 ( .A(n27082), .B(n27081), .Z(n35594) );
  ANDN U46435 ( .B(n27086), .A(n27085), .Z(n54574) );
  AND U46436 ( .A(n27088), .B(n27087), .Z(n54573) );
  AND U46437 ( .A(n54560), .B(n27089), .Z(n35551) );
  NANDN U46438 ( .A(y[2389]), .B(x[2389]), .Z(n27094) );
  IV U46439 ( .A(n27092), .Z(n27093) );
  AND U46440 ( .A(n27094), .B(n27093), .Z(n54554) );
  IV U46441 ( .A(n27095), .Z(n27096) );
  AND U46442 ( .A(n27097), .B(n27096), .Z(n54553) );
  NAND U46443 ( .A(n27099), .B(n27098), .Z(n54552) );
  AND U46444 ( .A(n27100), .B(n54548), .Z(n35531) );
  AND U46445 ( .A(n27102), .B(n27101), .Z(n35514) );
  AND U46446 ( .A(n27104), .B(n27103), .Z(n35508) );
  AND U46447 ( .A(n27106), .B(n27105), .Z(n35502) );
  AND U46448 ( .A(n27108), .B(n27107), .Z(n35496) );
  AND U46449 ( .A(n27110), .B(n27109), .Z(n35490) );
  AND U46450 ( .A(n27112), .B(n27111), .Z(n35484) );
  IV U46451 ( .A(n27113), .Z(n54527) );
  NANDN U46452 ( .A(x[2358]), .B(y[2358]), .Z(n27114) );
  OR U46453 ( .A(n27115), .B(n27114), .Z(n27116) );
  AND U46454 ( .A(n54523), .B(n27116), .Z(n35464) );
  AND U46455 ( .A(n27117), .B(n54522), .Z(n35462) );
  NAND U46456 ( .A(n27119), .B(n27118), .Z(n35460) );
  AND U46457 ( .A(n27121), .B(n27120), .Z(n35458) );
  AND U46458 ( .A(n27123), .B(n27122), .Z(n35452) );
  NAND U46459 ( .A(n27125), .B(n27124), .Z(n35438) );
  AND U46460 ( .A(n27127), .B(n27126), .Z(n35436) );
  NAND U46461 ( .A(n27129), .B(n27128), .Z(n35434) );
  AND U46462 ( .A(n27131), .B(n27130), .Z(n35432) );
  AND U46463 ( .A(n27133), .B(n27132), .Z(n35430) );
  NAND U46464 ( .A(n27135), .B(n27134), .Z(n35428) );
  AND U46465 ( .A(n27137), .B(n27136), .Z(n35418) );
  AND U46466 ( .A(n27139), .B(n27138), .Z(n54504) );
  AND U46467 ( .A(n27143), .B(n27142), .Z(n52099) );
  IV U46468 ( .A(n27144), .Z(n54498) );
  AND U46469 ( .A(n27146), .B(n27145), .Z(n35383) );
  AND U46470 ( .A(n27148), .B(n27147), .Z(n35377) );
  AND U46471 ( .A(n27150), .B(n27149), .Z(n35371) );
  OR U46472 ( .A(n27152), .B(n27151), .Z(n27153) );
  NAND U46473 ( .A(n27154), .B(n27153), .Z(n27155) );
  NANDN U46474 ( .A(n27156), .B(n27155), .Z(n54488) );
  AND U46475 ( .A(n27157), .B(n54486), .Z(n54484) );
  NAND U46476 ( .A(n54482), .B(n27158), .Z(n35352) );
  NOR U46477 ( .A(n27162), .B(n27161), .Z(n35338) );
  AND U46478 ( .A(n27164), .B(n27163), .Z(n35332) );
  ANDN U46479 ( .B(y[2306]), .A(x[2306]), .Z(n52105) );
  AND U46480 ( .A(n27166), .B(n27165), .Z(n35316) );
  AND U46481 ( .A(n27168), .B(n27167), .Z(n35310) );
  XNOR U46482 ( .A(y[2300]), .B(x[2300]), .Z(n54469) );
  AND U46483 ( .A(n27170), .B(n27169), .Z(n35298) );
  IV U46484 ( .A(n27171), .Z(n54461) );
  AND U46485 ( .A(n27172), .B(n54461), .Z(n35288) );
  NAND U46486 ( .A(n27174), .B(n27173), .Z(n54460) );
  IV U46487 ( .A(n27175), .Z(n54459) );
  AND U46488 ( .A(n27176), .B(n54459), .Z(n35285) );
  IV U46489 ( .A(n27177), .Z(n54458) );
  AND U46490 ( .A(n27179), .B(n27178), .Z(n35280) );
  NANDN U46491 ( .A(x[2288]), .B(y[2288]), .Z(n27181) );
  NAND U46492 ( .A(n27181), .B(n27180), .Z(n35278) );
  AND U46493 ( .A(n27182), .B(n52111), .Z(n35269) );
  NAND U46494 ( .A(n27184), .B(n27183), .Z(n52112) );
  XNOR U46495 ( .A(x[2284]), .B(y[2284]), .Z(n27187) );
  IV U46496 ( .A(n27185), .Z(n27186) );
  AND U46497 ( .A(n27187), .B(n27186), .Z(n54450) );
  IV U46498 ( .A(n27188), .Z(n27189) );
  AND U46499 ( .A(n27190), .B(n27189), .Z(n54448) );
  AND U46500 ( .A(n27192), .B(n27191), .Z(n35251) );
  NAND U46501 ( .A(n27194), .B(n27193), .Z(n35249) );
  AND U46502 ( .A(n27196), .B(n27195), .Z(n35247) );
  IV U46503 ( .A(n27197), .Z(n27199) );
  NAND U46504 ( .A(n27199), .B(n27198), .Z(n54439) );
  IV U46505 ( .A(n27203), .Z(n27204) );
  AND U46506 ( .A(n27205), .B(n27204), .Z(n54435) );
  IV U46507 ( .A(n27206), .Z(n54434) );
  AND U46508 ( .A(n27208), .B(n27207), .Z(n35223) );
  AND U46509 ( .A(n27210), .B(n27209), .Z(n35205) );
  IV U46510 ( .A(n27211), .Z(n54419) );
  AND U46511 ( .A(n27212), .B(n54419), .Z(n35187) );
  NAND U46512 ( .A(n27214), .B(n27213), .Z(n54418) );
  AND U46513 ( .A(n27220), .B(n27219), .Z(n35171) );
  NAND U46514 ( .A(n27222), .B(n27221), .Z(n35169) );
  AND U46515 ( .A(n27223), .B(n52118), .Z(n35167) );
  IV U46516 ( .A(n27224), .Z(n54404) );
  NAND U46517 ( .A(n27226), .B(n27225), .Z(n35129) );
  IV U46518 ( .A(n27227), .Z(n54393) );
  IV U46519 ( .A(n27228), .Z(n54392) );
  IV U46520 ( .A(n27229), .Z(n54391) );
  NANDN U46521 ( .A(x[2226]), .B(y[2226]), .Z(n27231) );
  AND U46522 ( .A(n27231), .B(n27230), .Z(n35112) );
  NAND U46523 ( .A(n27233), .B(n27232), .Z(n35110) );
  AND U46524 ( .A(n27235), .B(n27234), .Z(n35108) );
  AND U46525 ( .A(n27237), .B(n27236), .Z(n35102) );
  IV U46526 ( .A(n27238), .Z(n54384) );
  IV U46527 ( .A(n27239), .Z(n54379) );
  ANDN U46528 ( .B(y[2208]), .A(x[2208]), .Z(n35076) );
  AND U46529 ( .A(n27245), .B(n27244), .Z(n35069) );
  AND U46530 ( .A(n27247), .B(n27246), .Z(n35063) );
  NAND U46531 ( .A(n27249), .B(n27248), .Z(n54356) );
  AND U46532 ( .A(n27251), .B(n27250), .Z(n35003) );
  NAND U46533 ( .A(n54346), .B(n27252), .Z(n34993) );
  NOR U46534 ( .A(n27254), .B(n27253), .Z(n34983) );
  AND U46535 ( .A(n27256), .B(n27255), .Z(n34977) );
  AND U46536 ( .A(n27258), .B(n27257), .Z(n54339) );
  AND U46537 ( .A(n27260), .B(n27259), .Z(n34957) );
  IV U46538 ( .A(n27261), .Z(n54328) );
  AND U46539 ( .A(n27262), .B(n54328), .Z(n34951) );
  IV U46540 ( .A(n27263), .Z(n54326) );
  IV U46541 ( .A(n27265), .Z(n27266) );
  AND U46542 ( .A(n27267), .B(n27266), .Z(n54308) );
  AND U46543 ( .A(n27268), .B(n54307), .Z(n34910) );
  NANDN U46544 ( .A(x[2144]), .B(y[2144]), .Z(n34905) );
  AND U46545 ( .A(n27270), .B(n27269), .Z(n34901) );
  AND U46546 ( .A(n27272), .B(n27271), .Z(n34895) );
  ANDN U46547 ( .B(y[2140]), .A(x[2140]), .Z(n34891) );
  AND U46548 ( .A(n27274), .B(n27273), .Z(n34889) );
  AND U46549 ( .A(n27276), .B(n27275), .Z(n34867) );
  AND U46550 ( .A(n27278), .B(n27277), .Z(n34861) );
  XNOR U46551 ( .A(x[2130]), .B(y[2130]), .Z(n34855) );
  AND U46552 ( .A(n27280), .B(n27279), .Z(n34834) );
  AND U46553 ( .A(n27282), .B(n27281), .Z(n34812) );
  IV U46554 ( .A(n27283), .Z(n54273) );
  IV U46555 ( .A(n27284), .Z(n54272) );
  IV U46556 ( .A(n27285), .Z(n54271) );
  AND U46557 ( .A(n27287), .B(n27286), .Z(n34774) );
  AND U46558 ( .A(n27289), .B(n27288), .Z(n34752) );
  IV U46559 ( .A(n27290), .Z(n54254) );
  XNOR U46560 ( .A(x[2092]), .B(y[2092]), .Z(n27291) );
  AND U46561 ( .A(n27292), .B(n27291), .Z(n54251) );
  AND U46562 ( .A(n27296), .B(n27295), .Z(n54248) );
  NAND U46563 ( .A(n54245), .B(n27297), .Z(n34730) );
  IV U46564 ( .A(n27298), .Z(n54239) );
  AND U46565 ( .A(n54244), .B(n54239), .Z(n34728) );
  IV U46566 ( .A(n27303), .Z(n54223) );
  AND U46567 ( .A(n27304), .B(n54223), .Z(n34709) );
  AND U46568 ( .A(n27306), .B(n27305), .Z(n34704) );
  NAND U46569 ( .A(n27308), .B(n27307), .Z(n34694) );
  AND U46570 ( .A(n27310), .B(n27309), .Z(n34692) );
  NAND U46571 ( .A(n27312), .B(n27311), .Z(n34690) );
  AND U46572 ( .A(n27314), .B(n27313), .Z(n34688) );
  ANDN U46573 ( .B(y[2068]), .A(x[2068]), .Z(n34684) );
  AND U46574 ( .A(n27316), .B(n27315), .Z(n34682) );
  NOR U46575 ( .A(n27318), .B(n27317), .Z(n34672) );
  IV U46576 ( .A(n27319), .Z(n54202) );
  AND U46577 ( .A(n27320), .B(n54202), .Z(n34666) );
  AND U46578 ( .A(n27321), .B(n54196), .Z(n34650) );
  AND U46579 ( .A(n27323), .B(n27322), .Z(n34645) );
  NAND U46580 ( .A(n27325), .B(n27324), .Z(n54189) );
  AND U46581 ( .A(n54188), .B(n27326), .Z(n34636) );
  NANDN U46582 ( .A(x[2048]), .B(y[2048]), .Z(n34631) );
  AND U46583 ( .A(n27328), .B(n27327), .Z(n34615) );
  AND U46584 ( .A(n27330), .B(n27329), .Z(n34605) );
  AND U46585 ( .A(n27332), .B(n27331), .Z(n34599) );
  AND U46586 ( .A(n27334), .B(n27333), .Z(n34585) );
  NAND U46587 ( .A(n27336), .B(n27335), .Z(n34583) );
  AND U46588 ( .A(n27338), .B(n27337), .Z(n34581) );
  NAND U46589 ( .A(n27340), .B(n27339), .Z(n34579) );
  AND U46590 ( .A(n27342), .B(n27341), .Z(n34577) );
  AND U46591 ( .A(n27344), .B(n27343), .Z(n54166) );
  AND U46592 ( .A(n54161), .B(n27345), .Z(n34560) );
  IV U46593 ( .A(n27350), .Z(n27351) );
  AND U46594 ( .A(n27352), .B(n27351), .Z(n54153) );
  IV U46595 ( .A(n27353), .Z(n27355) );
  NAND U46596 ( .A(n27355), .B(n27354), .Z(n54152) );
  IV U46597 ( .A(n27356), .Z(n54151) );
  AND U46598 ( .A(n27357), .B(n54151), .Z(n34543) );
  AND U46599 ( .A(n27359), .B(n27358), .Z(n34538) );
  IV U46600 ( .A(n27360), .Z(n54144) );
  IV U46601 ( .A(n27363), .Z(n54140) );
  NAND U46602 ( .A(n54135), .B(n27364), .Z(n34505) );
  AND U46603 ( .A(n27366), .B(n27365), .Z(n54134) );
  IV U46604 ( .A(n27367), .Z(n54133) );
  AND U46605 ( .A(n27369), .B(n27368), .Z(n34495) );
  AND U46606 ( .A(n27371), .B(n27370), .Z(n34485) );
  NAND U46607 ( .A(n27373), .B(n27372), .Z(n34483) );
  AND U46608 ( .A(n27375), .B(n27374), .Z(n34481) );
  NAND U46609 ( .A(n27377), .B(n27376), .Z(n34479) );
  AND U46610 ( .A(n27379), .B(n27378), .Z(n34477) );
  NOR U46611 ( .A(n27381), .B(n27380), .Z(n34475) );
  AND U46612 ( .A(n27383), .B(n27382), .Z(n34469) );
  NAND U46613 ( .A(n54119), .B(n27384), .Z(n34460) );
  AND U46614 ( .A(n27386), .B(n27385), .Z(n54118) );
  AND U46615 ( .A(n27388), .B(n27387), .Z(n34451) );
  NAND U46616 ( .A(n27390), .B(n27389), .Z(n34449) );
  AND U46617 ( .A(n27392), .B(n27391), .Z(n34447) );
  AND U46618 ( .A(n27394), .B(n27393), .Z(n34441) );
  AND U46619 ( .A(n54108), .B(n27395), .Z(n34436) );
  AND U46620 ( .A(n27396), .B(n54106), .Z(n34432) );
  IV U46621 ( .A(n27397), .Z(n54103) );
  AND U46622 ( .A(n27398), .B(n54103), .Z(n34428) );
  NANDN U46623 ( .A(x[1972]), .B(y[1972]), .Z(n27399) );
  AND U46624 ( .A(n27399), .B(n54102), .Z(n34426) );
  NAND U46625 ( .A(n27401), .B(n27400), .Z(n34424) );
  NANDN U46626 ( .A(x[1970]), .B(y[1970]), .Z(n27403) );
  AND U46627 ( .A(n27403), .B(n27402), .Z(n34422) );
  IV U46628 ( .A(n27404), .Z(n52169) );
  NANDN U46629 ( .A(x[1958]), .B(y[1958]), .Z(n27410) );
  AND U46630 ( .A(n27410), .B(n27409), .Z(n34401) );
  AND U46631 ( .A(n27412), .B(n27411), .Z(n34391) );
  NAND U46632 ( .A(n27414), .B(n27413), .Z(n34389) );
  AND U46633 ( .A(n27416), .B(n27415), .Z(n34387) );
  AND U46634 ( .A(n27418), .B(n27417), .Z(n34381) );
  AND U46635 ( .A(n27420), .B(n27419), .Z(n34375) );
  AND U46636 ( .A(n27422), .B(n27421), .Z(n34369) );
  AND U46637 ( .A(n27424), .B(n27423), .Z(n34363) );
  AND U46638 ( .A(n27426), .B(n27425), .Z(n34357) );
  AND U46639 ( .A(n27428), .B(n27427), .Z(n34347) );
  IV U46640 ( .A(n27429), .Z(n54074) );
  IV U46641 ( .A(n27432), .Z(n27433) );
  AND U46642 ( .A(n27434), .B(n27433), .Z(n54069) );
  AND U46643 ( .A(n27436), .B(n27435), .Z(n54068) );
  AND U46644 ( .A(n54067), .B(n27437), .Z(n34333) );
  ANDN U46645 ( .B(y[1932]), .A(x[1932]), .Z(n27438) );
  NOR U46646 ( .A(n54066), .B(n27438), .Z(n34331) );
  OR U46647 ( .A(n27440), .B(n27439), .Z(n27441) );
  AND U46648 ( .A(n54062), .B(n27441), .Z(n34324) );
  IV U46649 ( .A(n27442), .Z(n54061) );
  AND U46650 ( .A(n27444), .B(n27443), .Z(n34319) );
  AND U46651 ( .A(n27446), .B(n27445), .Z(n34313) );
  AND U46652 ( .A(n54056), .B(n27447), .Z(n34308) );
  AND U46653 ( .A(n54053), .B(n27448), .Z(n34299) );
  AND U46654 ( .A(n27450), .B(n27449), .Z(n34274) );
  AND U46655 ( .A(n27456), .B(n27455), .Z(n34253) );
  NAND U46656 ( .A(n27458), .B(n27457), .Z(n34239) );
  NAND U46657 ( .A(n27459), .B(n54029), .Z(n34234) );
  NANDN U46658 ( .A(x[1892]), .B(y[1892]), .Z(n27461) );
  AND U46659 ( .A(n27461), .B(n27460), .Z(n54028) );
  AND U46660 ( .A(n27465), .B(n27464), .Z(n54026) );
  AND U46661 ( .A(n27469), .B(n27468), .Z(n34225) );
  NAND U46662 ( .A(n27471), .B(n27470), .Z(n34223) );
  AND U46663 ( .A(n27472), .B(n54019), .Z(n34221) );
  AND U46664 ( .A(n27474), .B(n27473), .Z(n54017) );
  NAND U46665 ( .A(n54016), .B(n27475), .Z(n34215) );
  IV U46666 ( .A(n27476), .Z(n54015) );
  AND U46667 ( .A(n27477), .B(n54015), .Z(n34213) );
  AND U46668 ( .A(n27479), .B(n27478), .Z(n34207) );
  AND U46669 ( .A(n27481), .B(n27480), .Z(n34197) );
  AND U46670 ( .A(n27483), .B(n27482), .Z(n34191) );
  AND U46671 ( .A(n27485), .B(n27484), .Z(n34185) );
  NAND U46672 ( .A(n27487), .B(n27486), .Z(n34171) );
  AND U46673 ( .A(n27489), .B(n27488), .Z(n34169) );
  NAND U46674 ( .A(n27491), .B(n27490), .Z(n34167) );
  AND U46675 ( .A(n27493), .B(n27492), .Z(n34165) );
  AND U46676 ( .A(n27495), .B(n27494), .Z(n34163) );
  NAND U46677 ( .A(n27497), .B(n27496), .Z(n34161) );
  AND U46678 ( .A(n27498), .B(n53998), .Z(n34159) );
  NANDN U46679 ( .A(x[1860]), .B(y[1860]), .Z(n27500) );
  NAND U46680 ( .A(n27500), .B(n27499), .Z(n52197) );
  AND U46681 ( .A(n27504), .B(n27503), .Z(n53995) );
  ANDN U46682 ( .B(y[1846]), .A(x[1846]), .Z(n27509) );
  NOR U46683 ( .A(n27510), .B(n27509), .Z(n34129) );
  AND U46684 ( .A(n27512), .B(n27511), .Z(n34123) );
  ANDN U46685 ( .B(y[1842]), .A(x[1842]), .Z(n53977) );
  AND U46686 ( .A(n27514), .B(n27513), .Z(n53976) );
  NAND U46687 ( .A(n53966), .B(n27517), .Z(n34096) );
  AND U46688 ( .A(n27518), .B(n53965), .Z(n34094) );
  ANDN U46689 ( .B(y[1832]), .A(x[1832]), .Z(n34092) );
  AND U46690 ( .A(n27520), .B(n27519), .Z(n34068) );
  NAND U46691 ( .A(n52199), .B(n27521), .Z(n34059) );
  IV U46692 ( .A(n27526), .Z(n27527) );
  AND U46693 ( .A(n27528), .B(n27527), .Z(n53950) );
  IV U46694 ( .A(n27529), .Z(n27531) );
  NAND U46695 ( .A(n27531), .B(n27530), .Z(n53949) );
  AND U46696 ( .A(n53947), .B(n27532), .Z(n34050) );
  NAND U46697 ( .A(n27534), .B(n27533), .Z(n34033) );
  AND U46698 ( .A(n27536), .B(n27535), .Z(n34031) );
  NAND U46699 ( .A(n53940), .B(n27537), .Z(n34029) );
  AND U46700 ( .A(n27538), .B(n53939), .Z(n34027) );
  NANDN U46701 ( .A(x[1806]), .B(y[1806]), .Z(n27544) );
  IV U46702 ( .A(n27542), .Z(n27543) );
  AND U46703 ( .A(n27544), .B(n27543), .Z(n53936) );
  IV U46704 ( .A(n27545), .Z(n27547) );
  NAND U46705 ( .A(n27547), .B(n27546), .Z(n53935) );
  IV U46706 ( .A(n27548), .Z(n53934) );
  AND U46707 ( .A(n27549), .B(n53934), .Z(n34021) );
  OR U46708 ( .A(n27551), .B(n27550), .Z(n27552) );
  AND U46709 ( .A(n53923), .B(n27552), .Z(n34003) );
  NAND U46710 ( .A(n53922), .B(n27553), .Z(n34001) );
  AND U46711 ( .A(n27555), .B(n27554), .Z(n33999) );
  XNOR U46712 ( .A(y[1791]), .B(x[1791]), .Z(n33991) );
  NAND U46713 ( .A(n27557), .B(n27556), .Z(n33979) );
  AND U46714 ( .A(n27559), .B(n27558), .Z(n33977) );
  IV U46715 ( .A(n27562), .Z(n53904) );
  AND U46716 ( .A(n27568), .B(n53895), .Z(n33958) );
  NAND U46717 ( .A(n27570), .B(n27569), .Z(n33941) );
  AND U46718 ( .A(n27572), .B(n27571), .Z(n33939) );
  NAND U46719 ( .A(n27574), .B(n27573), .Z(n33937) );
  AND U46720 ( .A(n27576), .B(n27575), .Z(n33935) );
  AND U46721 ( .A(n53883), .B(n27577), .Z(n33929) );
  AND U46722 ( .A(n27581), .B(n27580), .Z(n33923) );
  AND U46723 ( .A(n27583), .B(n27582), .Z(n33921) );
  IV U46724 ( .A(n27584), .Z(n53875) );
  AND U46725 ( .A(n27585), .B(n53875), .Z(n33919) );
  NAND U46726 ( .A(n52213), .B(n27586), .Z(n33917) );
  AND U46727 ( .A(n53863), .B(n27587), .Z(n33892) );
  NAND U46728 ( .A(n27591), .B(n27590), .Z(n53860) );
  IV U46729 ( .A(n27592), .Z(n53859) );
  AND U46730 ( .A(n27593), .B(n53859), .Z(n33885) );
  IV U46731 ( .A(n27594), .Z(n53857) );
  NOR U46732 ( .A(n53857), .B(n27595), .Z(n33883) );
  AND U46733 ( .A(n27597), .B(n27596), .Z(n33877) );
  NANDN U46734 ( .A(x[1728]), .B(y[1728]), .Z(n53851) );
  NOR U46735 ( .A(n27599), .B(n27598), .Z(n33868) );
  IV U46736 ( .A(n27604), .Z(n53844) );
  IV U46737 ( .A(n27605), .Z(n53843) );
  AND U46738 ( .A(n27606), .B(n53843), .Z(n33856) );
  NAND U46739 ( .A(n52221), .B(n27607), .Z(n33847) );
  IV U46740 ( .A(n27610), .Z(n53837) );
  AND U46741 ( .A(n27612), .B(n27611), .Z(n33838) );
  AND U46742 ( .A(n27614), .B(n27613), .Z(n33832) );
  NAND U46743 ( .A(n27616), .B(n27615), .Z(n33818) );
  AND U46744 ( .A(n27618), .B(n27617), .Z(n33812) );
  AND U46745 ( .A(n27620), .B(n27619), .Z(n33806) );
  AND U46746 ( .A(n27622), .B(n27621), .Z(n33800) );
  AND U46747 ( .A(n27624), .B(n27623), .Z(n33794) );
  AND U46748 ( .A(n27626), .B(n27625), .Z(n33788) );
  AND U46749 ( .A(n27628), .B(n27627), .Z(n33782) );
  AND U46750 ( .A(n53819), .B(n27629), .Z(n33777) );
  AND U46751 ( .A(n27633), .B(n27632), .Z(n53817) );
  AND U46752 ( .A(n52234), .B(n27636), .Z(n33772) );
  AND U46753 ( .A(n53814), .B(n27637), .Z(n33768) );
  IV U46754 ( .A(n27638), .Z(n27640) );
  NAND U46755 ( .A(n27640), .B(n27639), .Z(n53813) );
  IV U46756 ( .A(n27641), .Z(n53812) );
  AND U46757 ( .A(n27643), .B(n27642), .Z(n33759) );
  AND U46758 ( .A(n27645), .B(n27644), .Z(n33749) );
  AND U46759 ( .A(n53800), .B(n27646), .Z(n33736) );
  OR U46760 ( .A(n27650), .B(n27649), .Z(n27651) );
  AND U46761 ( .A(n53797), .B(n27651), .Z(n33729) );
  AND U46762 ( .A(n27653), .B(n27652), .Z(n33723) );
  AND U46763 ( .A(n27655), .B(n27654), .Z(n33717) );
  AND U46764 ( .A(n27657), .B(n27656), .Z(n33711) );
  AND U46765 ( .A(n27658), .B(n53780), .Z(n33701) );
  AND U46766 ( .A(n27660), .B(n27659), .Z(n33692) );
  NAND U46767 ( .A(n27662), .B(n27661), .Z(n33690) );
  AND U46768 ( .A(n27664), .B(n27663), .Z(n33688) );
  NAND U46769 ( .A(n27666), .B(n27665), .Z(n33686) );
  NANDN U46770 ( .A(x[1654]), .B(y[1654]), .Z(n27668) );
  AND U46771 ( .A(n27668), .B(n27667), .Z(n33684) );
  NAND U46772 ( .A(n27670), .B(n27669), .Z(n33682) );
  AND U46773 ( .A(n27672), .B(n27671), .Z(n33680) );
  AND U46774 ( .A(n27673), .B(n53754), .Z(n33674) );
  XNOR U46775 ( .A(y[1646]), .B(x[1646]), .Z(n33664) );
  AND U46776 ( .A(n27675), .B(n27674), .Z(n33660) );
  AND U46777 ( .A(n27677), .B(n27676), .Z(n33658) );
  NAND U46778 ( .A(n52241), .B(n27678), .Z(n33656) );
  IV U46779 ( .A(n27679), .Z(n53747) );
  AND U46780 ( .A(n27680), .B(n53747), .Z(n33654) );
  AND U46781 ( .A(n27682), .B(n27681), .Z(n52242) );
  AND U46782 ( .A(n27686), .B(n27685), .Z(n53745) );
  AND U46783 ( .A(n27687), .B(n52243), .Z(n33646) );
  ANDN U46784 ( .B(y[1634]), .A(x[1634]), .Z(n33641) );
  NAND U46785 ( .A(n27689), .B(n27688), .Z(n33634) );
  AND U46786 ( .A(n27693), .B(n27692), .Z(n33612) );
  AND U46787 ( .A(n27695), .B(n27694), .Z(n33590) );
  AND U46788 ( .A(n27697), .B(n27696), .Z(n33568) );
  IV U46789 ( .A(n27704), .Z(n27705) );
  AND U46790 ( .A(n27706), .B(n27705), .Z(n53700) );
  AND U46791 ( .A(n27707), .B(n53699), .Z(n33526) );
  AND U46792 ( .A(n27709), .B(n27708), .Z(n33521) );
  NAND U46793 ( .A(n27710), .B(n53683), .Z(n27712) );
  ANDN U46794 ( .B(n27712), .A(n27711), .Z(n27713) );
  NANDN U46795 ( .A(n27714), .B(n27713), .Z(n33493) );
  NOR U46796 ( .A(n27716), .B(n27715), .Z(n33487) );
  AND U46797 ( .A(n27718), .B(n27717), .Z(n33481) );
  NANDN U46798 ( .A(x[1576]), .B(y[1576]), .Z(n33475) );
  NAND U46799 ( .A(n27720), .B(n27719), .Z(n33471) );
  AND U46800 ( .A(n27722), .B(n27721), .Z(n33469) );
  NAND U46801 ( .A(n27724), .B(n27723), .Z(n33467) );
  AND U46802 ( .A(n27726), .B(n27725), .Z(n33465) );
  AND U46803 ( .A(n27728), .B(n27727), .Z(n33459) );
  NAND U46804 ( .A(n53650), .B(n27729), .Z(n33450) );
  AND U46805 ( .A(n27731), .B(n27730), .Z(n53649) );
  NANDN U46806 ( .A(x[1564]), .B(y[1564]), .Z(n33444) );
  NOR U46807 ( .A(n27733), .B(n27732), .Z(n33441) );
  AND U46808 ( .A(n27735), .B(n27734), .Z(n33435) );
  NAND U46809 ( .A(n27741), .B(n27740), .Z(n33409) );
  AND U46810 ( .A(n27743), .B(n27742), .Z(n33407) );
  NAND U46811 ( .A(n53621), .B(n27744), .Z(n33405) );
  AND U46812 ( .A(n27745), .B(n53622), .Z(n33403) );
  AND U46813 ( .A(n27747), .B(n27746), .Z(n33390) );
  NAND U46814 ( .A(n27749), .B(n27748), .Z(n33388) );
  NAND U46815 ( .A(n27751), .B(n27750), .Z(n33378) );
  AND U46816 ( .A(n27753), .B(n27752), .Z(n33376) );
  NAND U46817 ( .A(n27755), .B(n27754), .Z(n33374) );
  NANDN U46818 ( .A(x[1536]), .B(y[1536]), .Z(n27756) );
  AND U46819 ( .A(n27757), .B(n27756), .Z(n33372) );
  NANDN U46820 ( .A(x[1530]), .B(y[1530]), .Z(n27759) );
  AND U46821 ( .A(n27759), .B(n27758), .Z(n33356) );
  AND U46822 ( .A(n27761), .B(n27760), .Z(n33350) );
  AND U46823 ( .A(n27763), .B(n27762), .Z(n53597) );
  NOR U46824 ( .A(n27767), .B(n27766), .Z(n33331) );
  NAND U46825 ( .A(n27769), .B(n27768), .Z(n53588) );
  ANDN U46826 ( .B(y[1512]), .A(x[1512]), .Z(n33314) );
  AND U46827 ( .A(n27775), .B(n27774), .Z(n33307) );
  NAND U46828 ( .A(n27777), .B(n27776), .Z(n33305) );
  AND U46829 ( .A(n27779), .B(n27778), .Z(n33303) );
  IV U46830 ( .A(n27780), .Z(n53577) );
  AND U46831 ( .A(n27781), .B(n53577), .Z(n33297) );
  NAND U46832 ( .A(n27783), .B(n27782), .Z(n53576) );
  AND U46833 ( .A(n27784), .B(n53575), .Z(n33294) );
  IV U46834 ( .A(n27785), .Z(n53574) );
  NAND U46835 ( .A(n53569), .B(n27786), .Z(n33282) );
  AND U46836 ( .A(n27790), .B(n27789), .Z(n33273) );
  AND U46837 ( .A(n27792), .B(n27791), .Z(n33267) );
  AND U46838 ( .A(n27794), .B(n27793), .Z(n33261) );
  NANDN U46839 ( .A(x[1490]), .B(y[1490]), .Z(n27795) );
  AND U46840 ( .A(n27796), .B(n27795), .Z(n33255) );
  AND U46841 ( .A(n27798), .B(n27797), .Z(n33249) );
  NOR U46842 ( .A(n27800), .B(n27799), .Z(n33239) );
  AND U46843 ( .A(n27801), .B(n52266), .Z(n33234) );
  NAND U46844 ( .A(n27803), .B(n27802), .Z(n33227) );
  OR U46845 ( .A(n27805), .B(n27804), .Z(n27806) );
  NAND U46846 ( .A(n27807), .B(n27806), .Z(n27808) );
  NANDN U46847 ( .A(n27809), .B(n27808), .Z(n53539) );
  AND U46848 ( .A(n27810), .B(n53538), .Z(n33198) );
  IV U46849 ( .A(n27811), .Z(n53537) );
  NAND U46850 ( .A(n53533), .B(n27812), .Z(n33186) );
  IV U46851 ( .A(n27815), .Z(n53531) );
  AND U46852 ( .A(n27817), .B(n27816), .Z(n33164) );
  NAND U46853 ( .A(n27819), .B(n27818), .Z(n33154) );
  AND U46854 ( .A(n27821), .B(n27820), .Z(n33152) );
  NAND U46855 ( .A(n27823), .B(n27822), .Z(n33150) );
  AND U46856 ( .A(n27825), .B(n27824), .Z(n33148) );
  OR U46857 ( .A(n27827), .B(n27826), .Z(n27828) );
  AND U46858 ( .A(n27829), .B(n27828), .Z(n33124) );
  IV U46859 ( .A(n27830), .Z(n53515) );
  AND U46860 ( .A(n27831), .B(n53515), .Z(n33121) );
  IV U46861 ( .A(n27834), .Z(n27835) );
  AND U46862 ( .A(n27836), .B(n27835), .Z(n53506) );
  AND U46863 ( .A(n27838), .B(n27837), .Z(n53505) );
  IV U46864 ( .A(n27839), .Z(n27840) );
  AND U46865 ( .A(n27841), .B(n27840), .Z(n53504) );
  AND U46866 ( .A(n27845), .B(n27844), .Z(n52279) );
  IV U46867 ( .A(n27846), .Z(n27847) );
  AND U46868 ( .A(n27848), .B(n27847), .Z(n53494) );
  NOR U46869 ( .A(n27850), .B(n27849), .Z(n33067) );
  AND U46870 ( .A(n53488), .B(n27851), .Z(n33061) );
  NAND U46871 ( .A(n27853), .B(n27852), .Z(n53487) );
  AND U46872 ( .A(n27854), .B(n53486), .Z(n33058) );
  IV U46873 ( .A(n27855), .Z(n53485) );
  AND U46874 ( .A(n27857), .B(n27856), .Z(n33049) );
  NAND U46875 ( .A(n27859), .B(n27858), .Z(n27860) );
  NANDN U46876 ( .A(n27861), .B(n27860), .Z(n33045) );
  IV U46877 ( .A(n27862), .Z(n53476) );
  AND U46878 ( .A(n27863), .B(n53476), .Z(n33036) );
  AND U46879 ( .A(n27865), .B(n27864), .Z(n33026) );
  NAND U46880 ( .A(n27869), .B(n27868), .Z(n53468) );
  AND U46881 ( .A(n27871), .B(n27870), .Z(n53467) );
  AND U46882 ( .A(n27873), .B(n27872), .Z(n33006) );
  NAND U46883 ( .A(n27875), .B(n27874), .Z(n33004) );
  AND U46884 ( .A(n27877), .B(n27876), .Z(n32994) );
  AND U46885 ( .A(n27878), .B(n53456), .Z(n32989) );
  IV U46886 ( .A(n27883), .Z(n27885) );
  ANDN U46887 ( .B(n27885), .A(n27884), .Z(n53453) );
  AND U46888 ( .A(n27887), .B(n27886), .Z(n52284) );
  IV U46889 ( .A(n27888), .Z(n27889) );
  OR U46890 ( .A(n27890), .B(n27889), .Z(n27891) );
  AND U46891 ( .A(n27892), .B(n27891), .Z(n53446) );
  NANDN U46892 ( .A(x[1372]), .B(y[1372]), .Z(n27894) );
  AND U46893 ( .A(n27894), .B(n27893), .Z(n32954) );
  AND U46894 ( .A(n27896), .B(n27895), .Z(n32944) );
  NAND U46895 ( .A(n27898), .B(n27897), .Z(n32942) );
  AND U46896 ( .A(n27900), .B(n27899), .Z(n32940) );
  AND U46897 ( .A(n27902), .B(n27901), .Z(n32930) );
  AND U46898 ( .A(n27904), .B(n27903), .Z(n32920) );
  AND U46899 ( .A(n27906), .B(n27905), .Z(n32914) );
  AND U46900 ( .A(n27908), .B(n27907), .Z(n32908) );
  AND U46901 ( .A(n27910), .B(n27909), .Z(n32902) );
  AND U46902 ( .A(n27912), .B(n27911), .Z(n32896) );
  IV U46903 ( .A(n27913), .Z(n52301) );
  AND U46904 ( .A(n27914), .B(n52301), .Z(n32886) );
  AND U46905 ( .A(n27916), .B(n27915), .Z(n32865) );
  NOR U46906 ( .A(n27918), .B(n27917), .Z(n32855) );
  AND U46907 ( .A(n27919), .B(n53412), .Z(n32850) );
  AND U46908 ( .A(n27921), .B(n27920), .Z(n32845) );
  NANDN U46909 ( .A(x[1334]), .B(y[1334]), .Z(n27923) );
  AND U46910 ( .A(n27923), .B(n27922), .Z(n32840) );
  NAND U46911 ( .A(n27925), .B(n27924), .Z(n32830) );
  AND U46912 ( .A(n27927), .B(n27926), .Z(n32828) );
  NAND U46913 ( .A(n27929), .B(n27928), .Z(n32826) );
  AND U46914 ( .A(n27931), .B(n27930), .Z(n32824) );
  AND U46915 ( .A(n27933), .B(n27932), .Z(n32818) );
  NOR U46916 ( .A(n27935), .B(n27934), .Z(n32808) );
  ANDN U46917 ( .B(y[1322]), .A(x[1322]), .Z(n32804) );
  AND U46918 ( .A(n27937), .B(n27936), .Z(n32786) );
  OR U46919 ( .A(n27939), .B(n27938), .Z(n27940) );
  AND U46920 ( .A(n27941), .B(n27940), .Z(n32763) );
  NAND U46921 ( .A(n27945), .B(n27944), .Z(n52309) );
  AND U46922 ( .A(n27947), .B(n27946), .Z(n32716) );
  NAND U46923 ( .A(n27949), .B(n27948), .Z(n32702) );
  AND U46924 ( .A(n27951), .B(n27950), .Z(n32700) );
  NAND U46925 ( .A(n27953), .B(n27952), .Z(n32690) );
  AND U46926 ( .A(n27955), .B(n27954), .Z(n32688) );
  NOR U46927 ( .A(n27957), .B(n27956), .Z(n32678) );
  AND U46928 ( .A(n27959), .B(n27958), .Z(n53328) );
  XNOR U46929 ( .A(x[1273]), .B(y[1273]), .Z(n32658) );
  NANDN U46930 ( .A(y[1267]), .B(x[1267]), .Z(n27964) );
  AND U46931 ( .A(n27965), .B(n27964), .Z(n53317) );
  AND U46932 ( .A(n27969), .B(n27968), .Z(n53315) );
  AND U46933 ( .A(n27970), .B(n53313), .Z(n32637) );
  NAND U46934 ( .A(n27972), .B(n27971), .Z(n32623) );
  AND U46935 ( .A(n27974), .B(n27973), .Z(n32621) );
  NOR U46936 ( .A(n27976), .B(n27975), .Z(n32611) );
  IV U46937 ( .A(n27977), .Z(n53301) );
  NAND U46938 ( .A(n27979), .B(n27978), .Z(n53299) );
  NAND U46939 ( .A(n53291), .B(n27980), .Z(n32576) );
  ANDN U46940 ( .B(y[1236]), .A(x[1236]), .Z(n32561) );
  NAND U46941 ( .A(n27986), .B(n27985), .Z(n32545) );
  AND U46942 ( .A(n27988), .B(n27987), .Z(n32543) );
  AND U46943 ( .A(n27990), .B(n27989), .Z(n32533) );
  NAND U46944 ( .A(n27992), .B(n27991), .Z(n52317) );
  AND U46945 ( .A(n27993), .B(n53272), .Z(n32520) );
  AND U46946 ( .A(n27995), .B(n27994), .Z(n53262) );
  IV U46947 ( .A(n28000), .Z(n28002) );
  NAND U46948 ( .A(n28002), .B(n28001), .Z(n53259) );
  IV U46949 ( .A(n28003), .Z(n53258) );
  NOR U46950 ( .A(n28005), .B(n28004), .Z(n32466) );
  AND U46951 ( .A(n28007), .B(n28006), .Z(n52320) );
  AND U46952 ( .A(n28008), .B(n52321), .Z(n32441) );
  NOR U46953 ( .A(n28010), .B(n28009), .Z(n32432) );
  NAND U46954 ( .A(n28014), .B(n28013), .Z(n53233) );
  AND U46955 ( .A(n28016), .B(n28015), .Z(n32400) );
  NANDN U46956 ( .A(x[1180]), .B(y[1180]), .Z(n32390) );
  NAND U46957 ( .A(n28018), .B(n28017), .Z(n32386) );
  AND U46958 ( .A(n28020), .B(n28019), .Z(n32384) );
  AND U46959 ( .A(n28022), .B(n28021), .Z(n32374) );
  NAND U46960 ( .A(n28024), .B(n28023), .Z(n53216) );
  AND U46961 ( .A(n53215), .B(n28025), .Z(n32365) );
  ANDN U46962 ( .B(y[1170]), .A(x[1170]), .Z(n32362) );
  NOR U46963 ( .A(n28027), .B(n28026), .Z(n32356) );
  IV U46964 ( .A(n28028), .Z(n53207) );
  IV U46965 ( .A(n28033), .Z(n53202) );
  NAND U46966 ( .A(n28035), .B(n28034), .Z(n32324) );
  AND U46967 ( .A(n28037), .B(n28036), .Z(n32322) );
  NAND U46968 ( .A(n28039), .B(n28038), .Z(n32312) );
  AND U46969 ( .A(n28041), .B(n28040), .Z(n32310) );
  AND U46970 ( .A(n28043), .B(n28042), .Z(n32300) );
  NAND U46971 ( .A(n28045), .B(n28044), .Z(n53186) );
  ANDN U46972 ( .B(y[1142]), .A(x[1142]), .Z(n32281) );
  ANDN U46973 ( .B(y[1140]), .A(x[1140]), .Z(n28047) );
  NOR U46974 ( .A(n28047), .B(n28046), .Z(n32273) );
  AND U46975 ( .A(n28049), .B(n28048), .Z(n32259) );
  NAND U46976 ( .A(n28051), .B(n28050), .Z(n32245) );
  AND U46977 ( .A(n28053), .B(n28052), .Z(n32243) );
  NAND U46978 ( .A(n28055), .B(n28054), .Z(n32233) );
  AND U46979 ( .A(n28057), .B(n28056), .Z(n32231) );
  AND U46980 ( .A(n28059), .B(n28058), .Z(n32221) );
  AND U46981 ( .A(n28062), .B(n53164), .Z(n32207) );
  ANDN U46982 ( .B(y[1116]), .A(x[1116]), .Z(n32198) );
  AND U46983 ( .A(n53147), .B(n28067), .Z(n32178) );
  AND U46984 ( .A(n28069), .B(n28068), .Z(n32157) );
  NAND U46985 ( .A(n28071), .B(n28070), .Z(n32115) );
  AND U46986 ( .A(n28073), .B(n28072), .Z(n32113) );
  NAND U46987 ( .A(n28075), .B(n28074), .Z(n32103) );
  AND U46988 ( .A(n28077), .B(n28076), .Z(n32101) );
  NAND U46989 ( .A(n28079), .B(n28078), .Z(n32091) );
  AND U46990 ( .A(n28081), .B(n28080), .Z(n32089) );
  NAND U46991 ( .A(n28083), .B(n28082), .Z(n32079) );
  AND U46992 ( .A(n28085), .B(n28084), .Z(n32077) );
  NOR U46993 ( .A(n28087), .B(n28086), .Z(n32067) );
  NAND U46994 ( .A(n28091), .B(n28090), .Z(n53089) );
  IV U46995 ( .A(n28092), .Z(n53088) );
  IV U46996 ( .A(n28093), .Z(n53084) );
  NAND U46997 ( .A(n28095), .B(n28094), .Z(n53082) );
  AND U46998 ( .A(n28096), .B(n53081), .Z(n32036) );
  AND U46999 ( .A(n28098), .B(n28097), .Z(n32011) );
  ANDN U47000 ( .B(y[1050]), .A(x[1050]), .Z(n31989) );
  ANDN U47001 ( .B(y[1048]), .A(x[1048]), .Z(n31981) );
  ANDN U47002 ( .B(y[1046]), .A(x[1046]), .Z(n31973) );
  NOR U47003 ( .A(n28100), .B(n28099), .Z(n31948) );
  AND U47004 ( .A(n53049), .B(n28101), .Z(n31929) );
  ANDN U47005 ( .B(y[1032]), .A(x[1032]), .Z(n31926) );
  AND U47006 ( .A(n28103), .B(n28102), .Z(n31924) );
  AND U47007 ( .A(n28105), .B(n28104), .Z(n31914) );
  NAND U47008 ( .A(n28107), .B(n28106), .Z(n53038) );
  AND U47009 ( .A(n53037), .B(n28108), .Z(n31901) );
  NOR U47010 ( .A(n28110), .B(n28109), .Z(n31892) );
  IV U47011 ( .A(n28111), .Z(n53028) );
  IV U47012 ( .A(n28112), .Z(n53027) );
  IV U47013 ( .A(n28115), .Z(n53024) );
  XNOR U47014 ( .A(x[1007]), .B(y[1007]), .Z(n31856) );
  NAND U47015 ( .A(n28117), .B(n28116), .Z(n31844) );
  AND U47016 ( .A(n28119), .B(n28118), .Z(n31842) );
  NOR U47017 ( .A(n28121), .B(n28120), .Z(n31832) );
  AND U47018 ( .A(n28122), .B(n53004), .Z(n31813) );
  ANDN U47019 ( .B(y[982]), .A(x[982]), .Z(n31774) );
  NOR U47020 ( .A(n28124), .B(n28123), .Z(n31768) );
  AND U47021 ( .A(n28126), .B(n28125), .Z(n52980) );
  NAND U47022 ( .A(n52978), .B(n28127), .Z(n31747) );
  NANDN U47023 ( .A(x[972]), .B(y[972]), .Z(n31744) );
  NANDN U47024 ( .A(x[970]), .B(y[970]), .Z(n28128) );
  AND U47025 ( .A(n28129), .B(n28128), .Z(n31738) );
  NAND U47026 ( .A(n28131), .B(n28130), .Z(n31709) );
  AND U47027 ( .A(n28133), .B(n28132), .Z(n31707) );
  NAND U47028 ( .A(n28135), .B(n28134), .Z(n31697) );
  AND U47029 ( .A(n28137), .B(n28136), .Z(n31695) );
  NAND U47030 ( .A(n28139), .B(n28138), .Z(n31685) );
  AND U47031 ( .A(n28141), .B(n28140), .Z(n31683) );
  NOR U47032 ( .A(n28143), .B(n28142), .Z(n31673) );
  AND U47033 ( .A(n28144), .B(n52945), .Z(n31654) );
  AND U47034 ( .A(n28146), .B(n28145), .Z(n31633) );
  ANDN U47035 ( .B(n28148), .A(n28147), .Z(n52935) );
  IV U47036 ( .A(n28149), .Z(n52931) );
  IV U47037 ( .A(n28150), .Z(n52930) );
  IV U47038 ( .A(n28151), .Z(n52924) );
  NOR U47039 ( .A(n28155), .B(n28154), .Z(n31591) );
  IV U47040 ( .A(n28156), .Z(n52914) );
  NANDN U47041 ( .A(x[914]), .B(y[914]), .Z(n28158) );
  AND U47042 ( .A(n28158), .B(n28157), .Z(n52912) );
  ANDN U47043 ( .B(y[912]), .A(x[912]), .Z(n28159) );
  NOR U47044 ( .A(n52910), .B(n28159), .Z(n31565) );
  AND U47045 ( .A(n28161), .B(n28160), .Z(n31559) );
  AND U47046 ( .A(n28163), .B(n28162), .Z(n31549) );
  NAND U47047 ( .A(n28165), .B(n28164), .Z(n31535) );
  AND U47048 ( .A(n28167), .B(n28166), .Z(n31533) );
  AND U47049 ( .A(n28169), .B(n28168), .Z(n31523) );
  NANDN U47050 ( .A(x[896]), .B(y[896]), .Z(n31513) );
  NAND U47051 ( .A(n28171), .B(n28170), .Z(n31509) );
  AND U47052 ( .A(n28173), .B(n28172), .Z(n31507) );
  NANDN U47053 ( .A(x[892]), .B(y[892]), .Z(n31501) );
  NANDN U47054 ( .A(n52375), .B(n28174), .Z(n28176) );
  ANDN U47055 ( .B(n28176), .A(n28175), .Z(n31477) );
  AND U47056 ( .A(n28178), .B(n28177), .Z(n31468) );
  ANDN U47057 ( .B(n28182), .A(n28181), .Z(n52872) );
  AND U47058 ( .A(n28184), .B(n28183), .Z(n31395) );
  ANDN U47059 ( .B(y[852]), .A(x[852]), .Z(n31377) );
  NAND U47060 ( .A(n28186), .B(n28185), .Z(n31369) );
  AND U47061 ( .A(n28188), .B(n28187), .Z(n31367) );
  AND U47062 ( .A(n28190), .B(n28189), .Z(n31357) );
  IV U47063 ( .A(n28191), .Z(n52861) );
  AND U47064 ( .A(n28192), .B(n52859), .Z(n31349) );
  ANDN U47065 ( .B(y[842]), .A(x[842]), .Z(n31346) );
  NAND U47066 ( .A(n28194), .B(n28193), .Z(n31340) );
  AND U47067 ( .A(n28196), .B(n28195), .Z(n31338) );
  NAND U47068 ( .A(n28198), .B(n28197), .Z(n52397) );
  NANDN U47069 ( .A(x[828]), .B(y[828]), .Z(n28199) );
  AND U47070 ( .A(n28200), .B(n28199), .Z(n31306) );
  NANDN U47071 ( .A(x[826]), .B(y[826]), .Z(n31296) );
  NAND U47072 ( .A(n28202), .B(n28201), .Z(n31280) );
  AND U47073 ( .A(n28204), .B(n28203), .Z(n31278) );
  AND U47074 ( .A(n28206), .B(n28205), .Z(n31268) );
  NAND U47075 ( .A(n28208), .B(n28207), .Z(n52805) );
  AND U47076 ( .A(n52804), .B(n28209), .Z(n31259) );
  NAND U47077 ( .A(n28211), .B(n28210), .Z(n31250) );
  AND U47078 ( .A(n28213), .B(n28212), .Z(n31248) );
  ANDN U47079 ( .B(y[806]), .A(x[806]), .Z(n28215) );
  NOR U47080 ( .A(n28215), .B(n28214), .Z(n31238) );
  AND U47081 ( .A(n28217), .B(n28216), .Z(n31224) );
  AND U47082 ( .A(n28219), .B(n28218), .Z(n31210) );
  NAND U47083 ( .A(n28221), .B(n28220), .Z(n52399) );
  AND U47084 ( .A(n28222), .B(n52764), .Z(n31197) );
  NOR U47085 ( .A(n28224), .B(n28223), .Z(n31188) );
  AND U47086 ( .A(n28226), .B(n28225), .Z(n52754) );
  AND U47087 ( .A(n28228), .B(n28227), .Z(n31154) );
  NOR U47088 ( .A(n28230), .B(n28229), .Z(n31132) );
  NAND U47089 ( .A(n28232), .B(n28231), .Z(n52736) );
  AND U47090 ( .A(n28233), .B(n52735), .Z(n31106) );
  NAND U47091 ( .A(n28235), .B(n28234), .Z(n31097) );
  AND U47092 ( .A(n28237), .B(n28236), .Z(n31095) );
  NAND U47093 ( .A(n28239), .B(n28238), .Z(n31085) );
  AND U47094 ( .A(n28241), .B(n28240), .Z(n31083) );
  NAND U47095 ( .A(n28243), .B(n28242), .Z(n31073) );
  AND U47096 ( .A(n28245), .B(n28244), .Z(n31071) );
  NOR U47097 ( .A(n28247), .B(n28246), .Z(n31061) );
  IV U47098 ( .A(n28248), .Z(n52702) );
  NOR U47099 ( .A(n28250), .B(n28249), .Z(n31039) );
  NOR U47100 ( .A(n28252), .B(n28251), .Z(n30996) );
  AND U47101 ( .A(n28254), .B(n28253), .Z(n30990) );
  NAND U47102 ( .A(n28256), .B(n28255), .Z(n52411) );
  AND U47103 ( .A(n28257), .B(n52669), .Z(n30981) );
  NOR U47104 ( .A(n28259), .B(n28258), .Z(n30972) );
  AND U47105 ( .A(n28261), .B(n28260), .Z(n52658) );
  IV U47106 ( .A(n28262), .Z(n52657) );
  XNOR U47107 ( .A(x[705]), .B(y[705]), .Z(n30932) );
  ANDN U47108 ( .B(y[696]), .A(x[696]), .Z(n28263) );
  NOR U47109 ( .A(n28264), .B(n28263), .Z(n30900) );
  AND U47110 ( .A(n28266), .B(n28265), .Z(n30878) );
  NOR U47111 ( .A(n28270), .B(n28269), .Z(n30850) );
  AND U47112 ( .A(n28274), .B(n28273), .Z(n30810) );
  ANDN U47113 ( .B(n28276), .A(n28275), .Z(n52591) );
  ANDN U47114 ( .B(y[652]), .A(x[652]), .Z(n30766) );
  AND U47115 ( .A(n28278), .B(n28277), .Z(n30746) );
  NAND U47116 ( .A(n28280), .B(n28279), .Z(n52428) );
  AND U47117 ( .A(n28282), .B(n28281), .Z(n30723) );
  AND U47118 ( .A(n28284), .B(n28283), .Z(n30701) );
  ANDN U47119 ( .B(y[630]), .A(x[630]), .Z(n30691) );
  AND U47120 ( .A(n28286), .B(n28285), .Z(n30679) );
  AND U47121 ( .A(n28288), .B(n28287), .Z(n30657) );
  ANDN U47122 ( .B(y[620]), .A(x[620]), .Z(n30655) );
  NAND U47123 ( .A(n28292), .B(n28291), .Z(n52522) );
  NANDN U47124 ( .A(x[610]), .B(y[610]), .Z(n28298) );
  NAND U47125 ( .A(n28298), .B(n28297), .Z(n52429) );
  IV U47126 ( .A(n28299), .Z(n28300) );
  AND U47127 ( .A(n28301), .B(n28300), .Z(n52514) );
  IV U47128 ( .A(n28302), .Z(n28303) );
  AND U47129 ( .A(n28304), .B(n28303), .Z(n52507) );
  NAND U47130 ( .A(n28306), .B(n28305), .Z(n52430) );
  IV U47131 ( .A(n28307), .Z(n28308) );
  AND U47132 ( .A(n28309), .B(n28308), .Z(n52506) );
  ANDN U47133 ( .B(y[602]), .A(x[602]), .Z(n30618) );
  NAND U47134 ( .A(n28313), .B(n28312), .Z(n52499) );
  IV U47135 ( .A(n28314), .Z(n28315) );
  AND U47136 ( .A(n28316), .B(n28315), .Z(n52498) );
  AND U47137 ( .A(n52494), .B(n52496), .Z(n30605) );
  IV U47138 ( .A(n28319), .Z(n28320) );
  AND U47139 ( .A(n28321), .B(n28320), .Z(n52490) );
  ANDN U47140 ( .B(n52488), .A(n52486), .Z(n30592) );
  IV U47141 ( .A(n28322), .Z(n28324) );
  NAND U47142 ( .A(n28324), .B(n28323), .Z(n52484) );
  AND U47143 ( .A(n28326), .B(n28325), .Z(n52483) );
  AND U47144 ( .A(n52478), .B(n52480), .Z(n30581) );
  IV U47145 ( .A(n28329), .Z(n28330) );
  AND U47146 ( .A(n28331), .B(n28330), .Z(n52476) );
  NAND U47147 ( .A(n28333), .B(n28332), .Z(n52432) );
  IV U47148 ( .A(n28336), .Z(n28337) );
  AND U47149 ( .A(n28338), .B(n28337), .Z(n52468) );
  NAND U47150 ( .A(n28340), .B(n28339), .Z(n52433) );
  NAND U47151 ( .A(n28344), .B(n28343), .Z(n52434) );
  IV U47152 ( .A(n28347), .Z(n28348) );
  AND U47153 ( .A(n28349), .B(n28348), .Z(n52463) );
  ANDN U47154 ( .B(y[566]), .A(x[566]), .Z(n30551) );
  AND U47155 ( .A(n52458), .B(n52460), .Z(n30548) );
  IV U47156 ( .A(n28350), .Z(n28351) );
  AND U47157 ( .A(n28352), .B(n28351), .Z(n52456) );
  IV U47158 ( .A(n28353), .Z(n28354) );
  AND U47159 ( .A(n28355), .B(n28354), .Z(n52455) );
  ANDN U47160 ( .B(y[560]), .A(x[560]), .Z(n30538) );
  AND U47161 ( .A(n52451), .B(n52453), .Z(n30535) );
  AND U47162 ( .A(n52445), .B(n52442), .Z(n30522) );
  NAND U47163 ( .A(n28363), .B(n28362), .Z(n52438) );
  NANDN U47164 ( .A(x[548]), .B(y[548]), .Z(n28364) );
  AND U47165 ( .A(n28365), .B(n28364), .Z(n30513) );
  ANDN U47166 ( .B(x[548]), .A(y[548]), .Z(n30511) );
  AND U47167 ( .A(n28367), .B(n28366), .Z(n30507) );
  AND U47168 ( .A(n28369), .B(n28368), .Z(n30485) );
  AND U47169 ( .A(n28371), .B(n28370), .Z(n30427) );
  AND U47170 ( .A(n28373), .B(n28372), .Z(n30405) );
  AND U47171 ( .A(n28375), .B(n28374), .Z(n30383) );
  AND U47172 ( .A(n28377), .B(n28376), .Z(n30361) );
  AND U47173 ( .A(n28379), .B(n28378), .Z(n30339) );
  AND U47174 ( .A(n28381), .B(n28380), .Z(n30317) );
  AND U47175 ( .A(n28383), .B(n28382), .Z(n30295) );
  AND U47176 ( .A(n28385), .B(n28384), .Z(n30273) );
  AND U47177 ( .A(n28387), .B(n28386), .Z(n30251) );
  AND U47178 ( .A(n28389), .B(n28388), .Z(n30229) );
  AND U47179 ( .A(n28391), .B(n28390), .Z(n30207) );
  AND U47180 ( .A(n28393), .B(n28392), .Z(n30185) );
  AND U47181 ( .A(n28395), .B(n28394), .Z(n30163) );
  AND U47182 ( .A(n28397), .B(n28396), .Z(n30141) );
  AND U47183 ( .A(n28399), .B(n28398), .Z(n30119) );
  AND U47184 ( .A(n28401), .B(n28400), .Z(n30097) );
  AND U47185 ( .A(n28403), .B(n28402), .Z(n30075) );
  AND U47186 ( .A(n28405), .B(n28404), .Z(n30053) );
  AND U47187 ( .A(n28407), .B(n28406), .Z(n30031) );
  AND U47188 ( .A(n28409), .B(n28408), .Z(n30009) );
  AND U47189 ( .A(n28411), .B(n28410), .Z(n29987) );
  AND U47190 ( .A(n28413), .B(n28412), .Z(n29965) );
  AND U47191 ( .A(n28415), .B(n28414), .Z(n29943) );
  AND U47192 ( .A(n28417), .B(n28416), .Z(n29921) );
  AND U47193 ( .A(n28419), .B(n28418), .Z(n29899) );
  AND U47194 ( .A(n28421), .B(n28420), .Z(n29877) );
  NANDN U47195 ( .A(x[364]), .B(y[364]), .Z(n28423) );
  AND U47196 ( .A(n28423), .B(n28422), .Z(n29855) );
  AND U47197 ( .A(n28425), .B(n28424), .Z(n29833) );
  AND U47198 ( .A(n28427), .B(n28426), .Z(n29811) );
  NANDN U47199 ( .A(x[350]), .B(y[350]), .Z(n29805) );
  AND U47200 ( .A(n28429), .B(n28428), .Z(n29789) );
  AND U47201 ( .A(n28431), .B(n28430), .Z(n29767) );
  NANDN U47202 ( .A(x[338]), .B(y[338]), .Z(n29761) );
  AND U47203 ( .A(n28433), .B(n28432), .Z(n29745) );
  AND U47204 ( .A(n28435), .B(n28434), .Z(n29723) );
  AND U47205 ( .A(n28437), .B(n28436), .Z(n29701) );
  AND U47206 ( .A(n28439), .B(n28438), .Z(n29679) );
  AND U47207 ( .A(n28441), .B(n28440), .Z(n29657) );
  AND U47208 ( .A(n28443), .B(n28442), .Z(n29635) );
  AND U47209 ( .A(n28445), .B(n28444), .Z(n29613) );
  AND U47210 ( .A(n28447), .B(n28446), .Z(n29591) );
  AND U47211 ( .A(n28449), .B(n28448), .Z(n29569) );
  AND U47212 ( .A(n28451), .B(n28450), .Z(n29547) );
  NANDN U47213 ( .A(x[274]), .B(y[274]), .Z(n28452) );
  AND U47214 ( .A(n28453), .B(n28452), .Z(n29527) );
  AND U47215 ( .A(n28455), .B(n28454), .Z(n29477) );
  AND U47216 ( .A(n28457), .B(n28456), .Z(n29455) );
  AND U47217 ( .A(n28459), .B(n28458), .Z(n29433) );
  AND U47218 ( .A(n28461), .B(n28460), .Z(n29411) );
  AND U47219 ( .A(n28463), .B(n28462), .Z(n29389) );
  NANDN U47220 ( .A(x[228]), .B(y[228]), .Z(n28465) );
  AND U47221 ( .A(n28465), .B(n28464), .Z(n29367) );
  AND U47222 ( .A(n28467), .B(n28466), .Z(n29345) );
  AND U47223 ( .A(n28469), .B(n28468), .Z(n29323) );
  AND U47224 ( .A(n28471), .B(n28470), .Z(n29301) );
  AND U47225 ( .A(n28473), .B(n28472), .Z(n29279) );
  AND U47226 ( .A(n28475), .B(n28474), .Z(n29257) );
  XNOR U47227 ( .A(x[189]), .B(y[189]), .Z(n29225) );
  AND U47228 ( .A(n28477), .B(n28476), .Z(n29217) );
  AND U47229 ( .A(n28479), .B(n28478), .Z(n29195) );
  AND U47230 ( .A(n28481), .B(n28480), .Z(n29173) );
  NANDN U47231 ( .A(x[172]), .B(y[172]), .Z(n29167) );
  AND U47232 ( .A(n28483), .B(n28482), .Z(n29151) );
  AND U47233 ( .A(n28485), .B(n28484), .Z(n29129) );
  AND U47234 ( .A(n28487), .B(n28486), .Z(n29107) );
  AND U47235 ( .A(n28489), .B(n28488), .Z(n29085) );
  AND U47236 ( .A(n28491), .B(n28490), .Z(n29057) );
  AND U47237 ( .A(n28493), .B(n28492), .Z(n29035) );
  AND U47238 ( .A(n28495), .B(n28494), .Z(n29013) );
  AND U47239 ( .A(n28497), .B(n28496), .Z(n28991) );
  AND U47240 ( .A(n28499), .B(n28498), .Z(n28969) );
  AND U47241 ( .A(n28501), .B(n28500), .Z(n28947) );
  AND U47242 ( .A(n28503), .B(n28502), .Z(n28925) );
  AND U47243 ( .A(n28505), .B(n28504), .Z(n28903) );
  AND U47244 ( .A(n28507), .B(n28506), .Z(n28881) );
  AND U47245 ( .A(n28509), .B(n28508), .Z(n28859) );
  AND U47246 ( .A(n28511), .B(n28510), .Z(n28837) );
  AND U47247 ( .A(n28513), .B(n28512), .Z(n28815) );
  AND U47248 ( .A(n28515), .B(n28514), .Z(n28793) );
  AND U47249 ( .A(n28517), .B(n28516), .Z(n28771) );
  AND U47250 ( .A(n28519), .B(n28518), .Z(n28749) );
  AND U47251 ( .A(n28521), .B(n28520), .Z(n28727) );
  AND U47252 ( .A(n28523), .B(n28522), .Z(n28705) );
  AND U47253 ( .A(n28525), .B(n28524), .Z(n28683) );
  AND U47254 ( .A(n28527), .B(n28526), .Z(n28655) );
  AND U47255 ( .A(n28529), .B(n28528), .Z(n28633) );
  NANDN U47256 ( .A(x[20]), .B(y[20]), .Z(n28531) );
  AND U47257 ( .A(n28531), .B(n28530), .Z(n28611) );
  AND U47258 ( .A(n28533), .B(n28532), .Z(n28589) );
  AND U47259 ( .A(n28535), .B(n28534), .Z(n28567) );
  AND U47260 ( .A(n28537), .B(n28536), .Z(n28545) );
  NANDN U47261 ( .A(x[0]), .B(y[0]), .Z(n28538) );
  NAND U47262 ( .A(n28539), .B(n28538), .Z(n28540) );
  NANDN U47263 ( .A(n28541), .B(n28540), .Z(n28543) );
  OR U47264 ( .A(n28543), .B(n28542), .Z(n28544) );
  AND U47265 ( .A(n28545), .B(n28544), .Z(n28547) );
  NOR U47266 ( .A(n28547), .B(n28546), .Z(n28548) );
  NANDN U47267 ( .A(n28549), .B(n28548), .Z(n28550) );
  AND U47268 ( .A(n28551), .B(n28550), .Z(n28553) );
  NAND U47269 ( .A(n28553), .B(n28552), .Z(n28555) );
  ANDN U47270 ( .B(n28555), .A(n28554), .Z(n28556) );
  NANDN U47271 ( .A(n28557), .B(n28556), .Z(n28561) );
  AND U47272 ( .A(n28559), .B(n28558), .Z(n28560) );
  NAND U47273 ( .A(n28561), .B(n28560), .Z(n28562) );
  NANDN U47274 ( .A(n28563), .B(n28562), .Z(n28565) );
  OR U47275 ( .A(n28565), .B(n28564), .Z(n28566) );
  AND U47276 ( .A(n28567), .B(n28566), .Z(n28569) );
  NOR U47277 ( .A(n28569), .B(n28568), .Z(n28570) );
  NANDN U47278 ( .A(n28571), .B(n28570), .Z(n28572) );
  AND U47279 ( .A(n28573), .B(n28572), .Z(n28575) );
  NAND U47280 ( .A(n28575), .B(n28574), .Z(n28577) );
  ANDN U47281 ( .B(n28577), .A(n28576), .Z(n28578) );
  NANDN U47282 ( .A(n28579), .B(n28578), .Z(n28583) );
  AND U47283 ( .A(n28581), .B(n28580), .Z(n28582) );
  NAND U47284 ( .A(n28583), .B(n28582), .Z(n28584) );
  NANDN U47285 ( .A(n28585), .B(n28584), .Z(n28587) );
  OR U47286 ( .A(n28587), .B(n28586), .Z(n28588) );
  AND U47287 ( .A(n28589), .B(n28588), .Z(n28591) );
  NOR U47288 ( .A(n28591), .B(n28590), .Z(n28592) );
  NANDN U47289 ( .A(n28593), .B(n28592), .Z(n28594) );
  AND U47290 ( .A(n28595), .B(n28594), .Z(n28597) );
  NAND U47291 ( .A(n28597), .B(n28596), .Z(n28599) );
  ANDN U47292 ( .B(n28599), .A(n28598), .Z(n28600) );
  NANDN U47293 ( .A(n28601), .B(n28600), .Z(n28602) );
  AND U47294 ( .A(n28603), .B(n28602), .Z(n28604) );
  NAND U47295 ( .A(n28605), .B(n28604), .Z(n28606) );
  NANDN U47296 ( .A(n28607), .B(n28606), .Z(n28609) );
  OR U47297 ( .A(n28609), .B(n28608), .Z(n28610) );
  AND U47298 ( .A(n28611), .B(n28610), .Z(n28613) );
  NOR U47299 ( .A(n28613), .B(n28612), .Z(n28614) );
  NANDN U47300 ( .A(n28615), .B(n28614), .Z(n28616) );
  AND U47301 ( .A(n28617), .B(n28616), .Z(n28619) );
  NAND U47302 ( .A(n28619), .B(n28618), .Z(n28621) );
  ANDN U47303 ( .B(n28621), .A(n28620), .Z(n28622) );
  NANDN U47304 ( .A(n28623), .B(n28622), .Z(n28627) );
  AND U47305 ( .A(n28625), .B(n28624), .Z(n28626) );
  NAND U47306 ( .A(n28627), .B(n28626), .Z(n28628) );
  NANDN U47307 ( .A(n28629), .B(n28628), .Z(n28631) );
  OR U47308 ( .A(n28631), .B(n28630), .Z(n28632) );
  AND U47309 ( .A(n28633), .B(n28632), .Z(n28635) );
  NOR U47310 ( .A(n28635), .B(n28634), .Z(n28636) );
  NANDN U47311 ( .A(n28637), .B(n28636), .Z(n28638) );
  AND U47312 ( .A(n28639), .B(n28638), .Z(n28641) );
  NAND U47313 ( .A(n28641), .B(n28640), .Z(n28643) );
  ANDN U47314 ( .B(n28643), .A(n28642), .Z(n28644) );
  NANDN U47315 ( .A(n28645), .B(n28644), .Z(n28649) );
  AND U47316 ( .A(n28647), .B(n28646), .Z(n28648) );
  NAND U47317 ( .A(n28649), .B(n28648), .Z(n28650) );
  NANDN U47318 ( .A(n28651), .B(n28650), .Z(n28653) );
  OR U47319 ( .A(n28653), .B(n28652), .Z(n28654) );
  AND U47320 ( .A(n28655), .B(n28654), .Z(n28657) );
  NOR U47321 ( .A(n28657), .B(n28656), .Z(n28658) );
  NANDN U47322 ( .A(n28659), .B(n28658), .Z(n28660) );
  AND U47323 ( .A(n28661), .B(n28660), .Z(n28663) );
  NAND U47324 ( .A(n28663), .B(n28662), .Z(n28665) );
  ANDN U47325 ( .B(n28665), .A(n28664), .Z(n28666) );
  NANDN U47326 ( .A(n28667), .B(n28666), .Z(n28671) );
  AND U47327 ( .A(n28669), .B(n28668), .Z(n28670) );
  NAND U47328 ( .A(n28671), .B(n28670), .Z(n28672) );
  NANDN U47329 ( .A(n28673), .B(n28672), .Z(n28675) );
  OR U47330 ( .A(n28675), .B(n28674), .Z(n28676) );
  NAND U47331 ( .A(n28677), .B(n28676), .Z(n28678) );
  NANDN U47332 ( .A(n28679), .B(n28678), .Z(n28681) );
  OR U47333 ( .A(n28681), .B(n28680), .Z(n28682) );
  AND U47334 ( .A(n28683), .B(n28682), .Z(n28685) );
  NOR U47335 ( .A(n28685), .B(n28684), .Z(n28686) );
  NANDN U47336 ( .A(n28687), .B(n28686), .Z(n28688) );
  AND U47337 ( .A(n28689), .B(n28688), .Z(n28691) );
  NAND U47338 ( .A(n28691), .B(n28690), .Z(n28693) );
  ANDN U47339 ( .B(n28693), .A(n28692), .Z(n28694) );
  NANDN U47340 ( .A(n28695), .B(n28694), .Z(n28699) );
  AND U47341 ( .A(n28697), .B(n28696), .Z(n28698) );
  NAND U47342 ( .A(n28699), .B(n28698), .Z(n28700) );
  NANDN U47343 ( .A(n28701), .B(n28700), .Z(n28703) );
  OR U47344 ( .A(n28703), .B(n28702), .Z(n28704) );
  AND U47345 ( .A(n28705), .B(n28704), .Z(n28707) );
  NOR U47346 ( .A(n28707), .B(n28706), .Z(n28708) );
  NANDN U47347 ( .A(n28709), .B(n28708), .Z(n28710) );
  AND U47348 ( .A(n28711), .B(n28710), .Z(n28713) );
  NAND U47349 ( .A(n28713), .B(n28712), .Z(n28715) );
  ANDN U47350 ( .B(n28715), .A(n28714), .Z(n28716) );
  NANDN U47351 ( .A(n28717), .B(n28716), .Z(n28721) );
  AND U47352 ( .A(n28719), .B(n28718), .Z(n28720) );
  NAND U47353 ( .A(n28721), .B(n28720), .Z(n28722) );
  NANDN U47354 ( .A(n28723), .B(n28722), .Z(n28725) );
  OR U47355 ( .A(n28725), .B(n28724), .Z(n28726) );
  AND U47356 ( .A(n28727), .B(n28726), .Z(n28729) );
  NOR U47357 ( .A(n28729), .B(n28728), .Z(n28730) );
  NANDN U47358 ( .A(n28731), .B(n28730), .Z(n28732) );
  AND U47359 ( .A(n28733), .B(n28732), .Z(n28735) );
  NAND U47360 ( .A(n28735), .B(n28734), .Z(n28737) );
  ANDN U47361 ( .B(n28737), .A(n28736), .Z(n28738) );
  NANDN U47362 ( .A(n28739), .B(n28738), .Z(n28743) );
  AND U47363 ( .A(n28741), .B(n28740), .Z(n28742) );
  NAND U47364 ( .A(n28743), .B(n28742), .Z(n28744) );
  NANDN U47365 ( .A(n28745), .B(n28744), .Z(n28747) );
  OR U47366 ( .A(n28747), .B(n28746), .Z(n28748) );
  AND U47367 ( .A(n28749), .B(n28748), .Z(n28751) );
  NOR U47368 ( .A(n28751), .B(n28750), .Z(n28752) );
  NANDN U47369 ( .A(n28753), .B(n28752), .Z(n28754) );
  AND U47370 ( .A(n28755), .B(n28754), .Z(n28757) );
  NAND U47371 ( .A(n28757), .B(n28756), .Z(n28759) );
  ANDN U47372 ( .B(n28759), .A(n28758), .Z(n28760) );
  NANDN U47373 ( .A(n28761), .B(n28760), .Z(n28765) );
  AND U47374 ( .A(n28763), .B(n28762), .Z(n28764) );
  NAND U47375 ( .A(n28765), .B(n28764), .Z(n28766) );
  NANDN U47376 ( .A(n28767), .B(n28766), .Z(n28769) );
  OR U47377 ( .A(n28769), .B(n28768), .Z(n28770) );
  AND U47378 ( .A(n28771), .B(n28770), .Z(n28773) );
  NOR U47379 ( .A(n28773), .B(n28772), .Z(n28774) );
  NANDN U47380 ( .A(n28775), .B(n28774), .Z(n28776) );
  AND U47381 ( .A(n28777), .B(n28776), .Z(n28779) );
  NAND U47382 ( .A(n28779), .B(n28778), .Z(n28781) );
  ANDN U47383 ( .B(n28781), .A(n28780), .Z(n28782) );
  NANDN U47384 ( .A(n28783), .B(n28782), .Z(n28787) );
  AND U47385 ( .A(n28785), .B(n28784), .Z(n28786) );
  NAND U47386 ( .A(n28787), .B(n28786), .Z(n28788) );
  NANDN U47387 ( .A(n28789), .B(n28788), .Z(n28791) );
  OR U47388 ( .A(n28791), .B(n28790), .Z(n28792) );
  AND U47389 ( .A(n28793), .B(n28792), .Z(n28795) );
  NOR U47390 ( .A(n28795), .B(n28794), .Z(n28796) );
  NANDN U47391 ( .A(n28797), .B(n28796), .Z(n28798) );
  AND U47392 ( .A(n28799), .B(n28798), .Z(n28801) );
  NAND U47393 ( .A(n28801), .B(n28800), .Z(n28803) );
  ANDN U47394 ( .B(n28803), .A(n28802), .Z(n28804) );
  NANDN U47395 ( .A(n28805), .B(n28804), .Z(n28809) );
  AND U47396 ( .A(n28807), .B(n28806), .Z(n28808) );
  NAND U47397 ( .A(n28809), .B(n28808), .Z(n28810) );
  NANDN U47398 ( .A(n28811), .B(n28810), .Z(n28813) );
  OR U47399 ( .A(n28813), .B(n28812), .Z(n28814) );
  AND U47400 ( .A(n28815), .B(n28814), .Z(n28817) );
  NOR U47401 ( .A(n28817), .B(n28816), .Z(n28818) );
  NANDN U47402 ( .A(n28819), .B(n28818), .Z(n28820) );
  AND U47403 ( .A(n28821), .B(n28820), .Z(n28823) );
  NAND U47404 ( .A(n28823), .B(n28822), .Z(n28825) );
  ANDN U47405 ( .B(n28825), .A(n28824), .Z(n28826) );
  NANDN U47406 ( .A(n28827), .B(n28826), .Z(n28831) );
  AND U47407 ( .A(n28829), .B(n28828), .Z(n28830) );
  NAND U47408 ( .A(n28831), .B(n28830), .Z(n28832) );
  NANDN U47409 ( .A(n28833), .B(n28832), .Z(n28835) );
  OR U47410 ( .A(n28835), .B(n28834), .Z(n28836) );
  AND U47411 ( .A(n28837), .B(n28836), .Z(n28839) );
  NOR U47412 ( .A(n28839), .B(n28838), .Z(n28840) );
  NANDN U47413 ( .A(n28841), .B(n28840), .Z(n28842) );
  AND U47414 ( .A(n28843), .B(n28842), .Z(n28845) );
  NAND U47415 ( .A(n28845), .B(n28844), .Z(n28847) );
  ANDN U47416 ( .B(n28847), .A(n28846), .Z(n28848) );
  NANDN U47417 ( .A(n28849), .B(n28848), .Z(n28853) );
  AND U47418 ( .A(n28851), .B(n28850), .Z(n28852) );
  NAND U47419 ( .A(n28853), .B(n28852), .Z(n28854) );
  NANDN U47420 ( .A(n28855), .B(n28854), .Z(n28857) );
  OR U47421 ( .A(n28857), .B(n28856), .Z(n28858) );
  AND U47422 ( .A(n28859), .B(n28858), .Z(n28861) );
  NOR U47423 ( .A(n28861), .B(n28860), .Z(n28862) );
  NANDN U47424 ( .A(n28863), .B(n28862), .Z(n28864) );
  AND U47425 ( .A(n28865), .B(n28864), .Z(n28867) );
  NAND U47426 ( .A(n28867), .B(n28866), .Z(n28869) );
  ANDN U47427 ( .B(n28869), .A(n28868), .Z(n28870) );
  NANDN U47428 ( .A(n28871), .B(n28870), .Z(n28875) );
  AND U47429 ( .A(n28873), .B(n28872), .Z(n28874) );
  NAND U47430 ( .A(n28875), .B(n28874), .Z(n28876) );
  NANDN U47431 ( .A(n28877), .B(n28876), .Z(n28879) );
  OR U47432 ( .A(n28879), .B(n28878), .Z(n28880) );
  AND U47433 ( .A(n28881), .B(n28880), .Z(n28883) );
  NOR U47434 ( .A(n28883), .B(n28882), .Z(n28884) );
  NANDN U47435 ( .A(n28885), .B(n28884), .Z(n28886) );
  AND U47436 ( .A(n28887), .B(n28886), .Z(n28889) );
  NAND U47437 ( .A(n28889), .B(n28888), .Z(n28891) );
  ANDN U47438 ( .B(n28891), .A(n28890), .Z(n28892) );
  NANDN U47439 ( .A(n28893), .B(n28892), .Z(n28897) );
  AND U47440 ( .A(n28895), .B(n28894), .Z(n28896) );
  NAND U47441 ( .A(n28897), .B(n28896), .Z(n28898) );
  NANDN U47442 ( .A(n28899), .B(n28898), .Z(n28901) );
  OR U47443 ( .A(n28901), .B(n28900), .Z(n28902) );
  AND U47444 ( .A(n28903), .B(n28902), .Z(n28905) );
  NOR U47445 ( .A(n28905), .B(n28904), .Z(n28906) );
  NANDN U47446 ( .A(n28907), .B(n28906), .Z(n28908) );
  AND U47447 ( .A(n28909), .B(n28908), .Z(n28911) );
  NAND U47448 ( .A(n28911), .B(n28910), .Z(n28913) );
  ANDN U47449 ( .B(n28913), .A(n28912), .Z(n28914) );
  NANDN U47450 ( .A(n28915), .B(n28914), .Z(n28919) );
  AND U47451 ( .A(n28917), .B(n28916), .Z(n28918) );
  NAND U47452 ( .A(n28919), .B(n28918), .Z(n28920) );
  NANDN U47453 ( .A(n28921), .B(n28920), .Z(n28923) );
  OR U47454 ( .A(n28923), .B(n28922), .Z(n28924) );
  AND U47455 ( .A(n28925), .B(n28924), .Z(n28927) );
  NOR U47456 ( .A(n28927), .B(n28926), .Z(n28928) );
  NANDN U47457 ( .A(n28929), .B(n28928), .Z(n28930) );
  AND U47458 ( .A(n28931), .B(n28930), .Z(n28933) );
  NAND U47459 ( .A(n28933), .B(n28932), .Z(n28935) );
  ANDN U47460 ( .B(n28935), .A(n28934), .Z(n28936) );
  NANDN U47461 ( .A(n28937), .B(n28936), .Z(n28941) );
  AND U47462 ( .A(n28939), .B(n28938), .Z(n28940) );
  NAND U47463 ( .A(n28941), .B(n28940), .Z(n28942) );
  NANDN U47464 ( .A(n28943), .B(n28942), .Z(n28945) );
  OR U47465 ( .A(n28945), .B(n28944), .Z(n28946) );
  AND U47466 ( .A(n28947), .B(n28946), .Z(n28949) );
  NOR U47467 ( .A(n28949), .B(n28948), .Z(n28950) );
  NANDN U47468 ( .A(n28951), .B(n28950), .Z(n28952) );
  AND U47469 ( .A(n28953), .B(n28952), .Z(n28955) );
  NAND U47470 ( .A(n28955), .B(n28954), .Z(n28957) );
  ANDN U47471 ( .B(n28957), .A(n28956), .Z(n28958) );
  NANDN U47472 ( .A(n28959), .B(n28958), .Z(n28963) );
  AND U47473 ( .A(n28961), .B(n28960), .Z(n28962) );
  NAND U47474 ( .A(n28963), .B(n28962), .Z(n28964) );
  NANDN U47475 ( .A(n28965), .B(n28964), .Z(n28967) );
  OR U47476 ( .A(n28967), .B(n28966), .Z(n28968) );
  AND U47477 ( .A(n28969), .B(n28968), .Z(n28971) );
  NOR U47478 ( .A(n28971), .B(n28970), .Z(n28972) );
  NANDN U47479 ( .A(n28973), .B(n28972), .Z(n28974) );
  AND U47480 ( .A(n28975), .B(n28974), .Z(n28977) );
  NAND U47481 ( .A(n28977), .B(n28976), .Z(n28979) );
  ANDN U47482 ( .B(n28979), .A(n28978), .Z(n28980) );
  NANDN U47483 ( .A(n28981), .B(n28980), .Z(n28985) );
  AND U47484 ( .A(n28983), .B(n28982), .Z(n28984) );
  NAND U47485 ( .A(n28985), .B(n28984), .Z(n28986) );
  NANDN U47486 ( .A(n28987), .B(n28986), .Z(n28989) );
  OR U47487 ( .A(n28989), .B(n28988), .Z(n28990) );
  AND U47488 ( .A(n28991), .B(n28990), .Z(n28993) );
  NOR U47489 ( .A(n28993), .B(n28992), .Z(n28994) );
  NANDN U47490 ( .A(n28995), .B(n28994), .Z(n28996) );
  AND U47491 ( .A(n28997), .B(n28996), .Z(n28999) );
  NAND U47492 ( .A(n28999), .B(n28998), .Z(n29001) );
  ANDN U47493 ( .B(n29001), .A(n29000), .Z(n29002) );
  NANDN U47494 ( .A(n29003), .B(n29002), .Z(n29007) );
  AND U47495 ( .A(n29005), .B(n29004), .Z(n29006) );
  NAND U47496 ( .A(n29007), .B(n29006), .Z(n29008) );
  NANDN U47497 ( .A(n29009), .B(n29008), .Z(n29011) );
  OR U47498 ( .A(n29011), .B(n29010), .Z(n29012) );
  AND U47499 ( .A(n29013), .B(n29012), .Z(n29015) );
  NOR U47500 ( .A(n29015), .B(n29014), .Z(n29016) );
  NANDN U47501 ( .A(n29017), .B(n29016), .Z(n29018) );
  AND U47502 ( .A(n29019), .B(n29018), .Z(n29021) );
  NAND U47503 ( .A(n29021), .B(n29020), .Z(n29023) );
  ANDN U47504 ( .B(n29023), .A(n29022), .Z(n29024) );
  NANDN U47505 ( .A(n29025), .B(n29024), .Z(n29029) );
  AND U47506 ( .A(n29027), .B(n29026), .Z(n29028) );
  NAND U47507 ( .A(n29029), .B(n29028), .Z(n29030) );
  NANDN U47508 ( .A(n29031), .B(n29030), .Z(n29033) );
  OR U47509 ( .A(n29033), .B(n29032), .Z(n29034) );
  AND U47510 ( .A(n29035), .B(n29034), .Z(n29037) );
  NOR U47511 ( .A(n29037), .B(n29036), .Z(n29038) );
  NANDN U47512 ( .A(n29039), .B(n29038), .Z(n29040) );
  AND U47513 ( .A(n29041), .B(n29040), .Z(n29043) );
  NAND U47514 ( .A(n29043), .B(n29042), .Z(n29045) );
  ANDN U47515 ( .B(n29045), .A(n29044), .Z(n29046) );
  NANDN U47516 ( .A(n29047), .B(n29046), .Z(n29051) );
  AND U47517 ( .A(n29049), .B(n29048), .Z(n29050) );
  NAND U47518 ( .A(n29051), .B(n29050), .Z(n29052) );
  NANDN U47519 ( .A(n29053), .B(n29052), .Z(n29055) );
  OR U47520 ( .A(n29055), .B(n29054), .Z(n29056) );
  AND U47521 ( .A(n29057), .B(n29056), .Z(n29059) );
  NOR U47522 ( .A(n29059), .B(n29058), .Z(n29060) );
  NANDN U47523 ( .A(n29061), .B(n29060), .Z(n29062) );
  AND U47524 ( .A(n29063), .B(n29062), .Z(n29065) );
  NAND U47525 ( .A(n29065), .B(n29064), .Z(n29067) );
  ANDN U47526 ( .B(n29067), .A(n29066), .Z(n29068) );
  NANDN U47527 ( .A(n29069), .B(n29068), .Z(n29073) );
  AND U47528 ( .A(n29071), .B(n29070), .Z(n29072) );
  NAND U47529 ( .A(n29073), .B(n29072), .Z(n29074) );
  NANDN U47530 ( .A(n29075), .B(n29074), .Z(n29077) );
  NAND U47531 ( .A(n29077), .B(n29076), .Z(n29078) );
  NANDN U47532 ( .A(n29079), .B(n29078), .Z(n29080) );
  AND U47533 ( .A(n29081), .B(n29080), .Z(n29082) );
  OR U47534 ( .A(n29083), .B(n29082), .Z(n29084) );
  AND U47535 ( .A(n29085), .B(n29084), .Z(n29087) );
  NOR U47536 ( .A(n29087), .B(n29086), .Z(n29088) );
  NANDN U47537 ( .A(n29089), .B(n29088), .Z(n29090) );
  AND U47538 ( .A(n29091), .B(n29090), .Z(n29093) );
  NAND U47539 ( .A(n29093), .B(n29092), .Z(n29095) );
  ANDN U47540 ( .B(n29095), .A(n29094), .Z(n29096) );
  NANDN U47541 ( .A(n29097), .B(n29096), .Z(n29101) );
  AND U47542 ( .A(n29099), .B(n29098), .Z(n29100) );
  NAND U47543 ( .A(n29101), .B(n29100), .Z(n29102) );
  NANDN U47544 ( .A(n29103), .B(n29102), .Z(n29105) );
  OR U47545 ( .A(n29105), .B(n29104), .Z(n29106) );
  AND U47546 ( .A(n29107), .B(n29106), .Z(n29109) );
  NOR U47547 ( .A(n29109), .B(n29108), .Z(n29110) );
  NANDN U47548 ( .A(n29111), .B(n29110), .Z(n29112) );
  AND U47549 ( .A(n29113), .B(n29112), .Z(n29115) );
  NAND U47550 ( .A(n29115), .B(n29114), .Z(n29117) );
  ANDN U47551 ( .B(n29117), .A(n29116), .Z(n29118) );
  NANDN U47552 ( .A(n29119), .B(n29118), .Z(n29123) );
  AND U47553 ( .A(n29121), .B(n29120), .Z(n29122) );
  NAND U47554 ( .A(n29123), .B(n29122), .Z(n29124) );
  NANDN U47555 ( .A(n29125), .B(n29124), .Z(n29127) );
  OR U47556 ( .A(n29127), .B(n29126), .Z(n29128) );
  AND U47557 ( .A(n29129), .B(n29128), .Z(n29131) );
  NOR U47558 ( .A(n29131), .B(n29130), .Z(n29132) );
  NANDN U47559 ( .A(n29133), .B(n29132), .Z(n29134) );
  AND U47560 ( .A(n29135), .B(n29134), .Z(n29137) );
  NAND U47561 ( .A(n29137), .B(n29136), .Z(n29139) );
  ANDN U47562 ( .B(n29139), .A(n29138), .Z(n29140) );
  NANDN U47563 ( .A(n29141), .B(n29140), .Z(n29145) );
  AND U47564 ( .A(n29143), .B(n29142), .Z(n29144) );
  NAND U47565 ( .A(n29145), .B(n29144), .Z(n29146) );
  NANDN U47566 ( .A(n29147), .B(n29146), .Z(n29149) );
  OR U47567 ( .A(n29149), .B(n29148), .Z(n29150) );
  AND U47568 ( .A(n29151), .B(n29150), .Z(n29153) );
  NOR U47569 ( .A(n29153), .B(n29152), .Z(n29154) );
  NANDN U47570 ( .A(n29155), .B(n29154), .Z(n29156) );
  AND U47571 ( .A(n29157), .B(n29156), .Z(n29159) );
  NAND U47572 ( .A(n29159), .B(n29158), .Z(n29161) );
  ANDN U47573 ( .B(n29161), .A(n29160), .Z(n29162) );
  NANDN U47574 ( .A(n29163), .B(n29162), .Z(n29164) );
  AND U47575 ( .A(n29165), .B(n29164), .Z(n29166) );
  NAND U47576 ( .A(n29167), .B(n29166), .Z(n29168) );
  NANDN U47577 ( .A(n29169), .B(n29168), .Z(n29171) );
  OR U47578 ( .A(n29171), .B(n29170), .Z(n29172) );
  AND U47579 ( .A(n29173), .B(n29172), .Z(n29175) );
  NOR U47580 ( .A(n29175), .B(n29174), .Z(n29176) );
  NANDN U47581 ( .A(n29177), .B(n29176), .Z(n29178) );
  AND U47582 ( .A(n29179), .B(n29178), .Z(n29181) );
  NAND U47583 ( .A(n29181), .B(n29180), .Z(n29183) );
  ANDN U47584 ( .B(n29183), .A(n29182), .Z(n29184) );
  NANDN U47585 ( .A(n29185), .B(n29184), .Z(n29189) );
  AND U47586 ( .A(n29187), .B(n29186), .Z(n29188) );
  NAND U47587 ( .A(n29189), .B(n29188), .Z(n29190) );
  NANDN U47588 ( .A(n29191), .B(n29190), .Z(n29193) );
  OR U47589 ( .A(n29193), .B(n29192), .Z(n29194) );
  AND U47590 ( .A(n29195), .B(n29194), .Z(n29197) );
  NOR U47591 ( .A(n29197), .B(n29196), .Z(n29198) );
  NANDN U47592 ( .A(n29199), .B(n29198), .Z(n29200) );
  AND U47593 ( .A(n29201), .B(n29200), .Z(n29203) );
  NAND U47594 ( .A(n29203), .B(n29202), .Z(n29205) );
  ANDN U47595 ( .B(n29205), .A(n29204), .Z(n29206) );
  NANDN U47596 ( .A(n29207), .B(n29206), .Z(n29211) );
  AND U47597 ( .A(n29209), .B(n29208), .Z(n29210) );
  NAND U47598 ( .A(n29211), .B(n29210), .Z(n29212) );
  NANDN U47599 ( .A(n29213), .B(n29212), .Z(n29215) );
  OR U47600 ( .A(n29215), .B(n29214), .Z(n29216) );
  AND U47601 ( .A(n29217), .B(n29216), .Z(n29219) );
  NOR U47602 ( .A(n29219), .B(n29218), .Z(n29220) );
  NANDN U47603 ( .A(n29221), .B(n29220), .Z(n29222) );
  AND U47604 ( .A(n29223), .B(n29222), .Z(n29224) );
  NAND U47605 ( .A(n29225), .B(n29224), .Z(n29226) );
  NAND U47606 ( .A(n29227), .B(n29226), .Z(n29228) );
  AND U47607 ( .A(n29229), .B(n29228), .Z(n29231) );
  OR U47608 ( .A(n29231), .B(n29230), .Z(n29232) );
  NAND U47609 ( .A(n29233), .B(n29232), .Z(n29234) );
  NANDN U47610 ( .A(n29235), .B(n29234), .Z(n29237) );
  NAND U47611 ( .A(n29237), .B(n29236), .Z(n29238) );
  NANDN U47612 ( .A(n29239), .B(n29238), .Z(n29240) );
  AND U47613 ( .A(n29241), .B(n29240), .Z(n29243) );
  NAND U47614 ( .A(n29243), .B(n29242), .Z(n29245) );
  ANDN U47615 ( .B(n29245), .A(n29244), .Z(n29246) );
  NANDN U47616 ( .A(n29247), .B(n29246), .Z(n29251) );
  AND U47617 ( .A(n29249), .B(n29248), .Z(n29250) );
  NAND U47618 ( .A(n29251), .B(n29250), .Z(n29252) );
  NANDN U47619 ( .A(n29253), .B(n29252), .Z(n29255) );
  OR U47620 ( .A(n29255), .B(n29254), .Z(n29256) );
  AND U47621 ( .A(n29257), .B(n29256), .Z(n29259) );
  NOR U47622 ( .A(n29259), .B(n29258), .Z(n29260) );
  NANDN U47623 ( .A(n29261), .B(n29260), .Z(n29262) );
  AND U47624 ( .A(n29263), .B(n29262), .Z(n29265) );
  NAND U47625 ( .A(n29265), .B(n29264), .Z(n29267) );
  ANDN U47626 ( .B(n29267), .A(n29266), .Z(n29268) );
  NANDN U47627 ( .A(n29269), .B(n29268), .Z(n29273) );
  AND U47628 ( .A(n29271), .B(n29270), .Z(n29272) );
  NAND U47629 ( .A(n29273), .B(n29272), .Z(n29274) );
  NANDN U47630 ( .A(n29275), .B(n29274), .Z(n29277) );
  OR U47631 ( .A(n29277), .B(n29276), .Z(n29278) );
  AND U47632 ( .A(n29279), .B(n29278), .Z(n29281) );
  NOR U47633 ( .A(n29281), .B(n29280), .Z(n29282) );
  NANDN U47634 ( .A(n29283), .B(n29282), .Z(n29284) );
  AND U47635 ( .A(n29285), .B(n29284), .Z(n29287) );
  NAND U47636 ( .A(n29287), .B(n29286), .Z(n29289) );
  ANDN U47637 ( .B(n29289), .A(n29288), .Z(n29290) );
  NANDN U47638 ( .A(n29291), .B(n29290), .Z(n29295) );
  AND U47639 ( .A(n29293), .B(n29292), .Z(n29294) );
  NAND U47640 ( .A(n29295), .B(n29294), .Z(n29296) );
  NANDN U47641 ( .A(n29297), .B(n29296), .Z(n29299) );
  OR U47642 ( .A(n29299), .B(n29298), .Z(n29300) );
  AND U47643 ( .A(n29301), .B(n29300), .Z(n29303) );
  NOR U47644 ( .A(n29303), .B(n29302), .Z(n29304) );
  NANDN U47645 ( .A(n29305), .B(n29304), .Z(n29306) );
  AND U47646 ( .A(n29307), .B(n29306), .Z(n29309) );
  NAND U47647 ( .A(n29309), .B(n29308), .Z(n29311) );
  ANDN U47648 ( .B(n29311), .A(n29310), .Z(n29312) );
  NANDN U47649 ( .A(n29313), .B(n29312), .Z(n29317) );
  AND U47650 ( .A(n29315), .B(n29314), .Z(n29316) );
  NAND U47651 ( .A(n29317), .B(n29316), .Z(n29318) );
  NANDN U47652 ( .A(n29319), .B(n29318), .Z(n29321) );
  OR U47653 ( .A(n29321), .B(n29320), .Z(n29322) );
  AND U47654 ( .A(n29323), .B(n29322), .Z(n29325) );
  NOR U47655 ( .A(n29325), .B(n29324), .Z(n29326) );
  NANDN U47656 ( .A(n29327), .B(n29326), .Z(n29328) );
  AND U47657 ( .A(n29329), .B(n29328), .Z(n29331) );
  NAND U47658 ( .A(n29331), .B(n29330), .Z(n29333) );
  ANDN U47659 ( .B(n29333), .A(n29332), .Z(n29334) );
  NANDN U47660 ( .A(n29335), .B(n29334), .Z(n29339) );
  AND U47661 ( .A(n29337), .B(n29336), .Z(n29338) );
  NAND U47662 ( .A(n29339), .B(n29338), .Z(n29340) );
  NANDN U47663 ( .A(n29341), .B(n29340), .Z(n29343) );
  OR U47664 ( .A(n29343), .B(n29342), .Z(n29344) );
  AND U47665 ( .A(n29345), .B(n29344), .Z(n29347) );
  NOR U47666 ( .A(n29347), .B(n29346), .Z(n29348) );
  NANDN U47667 ( .A(n29349), .B(n29348), .Z(n29350) );
  AND U47668 ( .A(n29351), .B(n29350), .Z(n29353) );
  NAND U47669 ( .A(n29353), .B(n29352), .Z(n29355) );
  ANDN U47670 ( .B(n29355), .A(n29354), .Z(n29356) );
  NANDN U47671 ( .A(n29357), .B(n29356), .Z(n29358) );
  AND U47672 ( .A(n29359), .B(n29358), .Z(n29360) );
  NAND U47673 ( .A(n29361), .B(n29360), .Z(n29362) );
  NANDN U47674 ( .A(n29363), .B(n29362), .Z(n29365) );
  OR U47675 ( .A(n29365), .B(n29364), .Z(n29366) );
  AND U47676 ( .A(n29367), .B(n29366), .Z(n29369) );
  NOR U47677 ( .A(n29369), .B(n29368), .Z(n29370) );
  NANDN U47678 ( .A(n29371), .B(n29370), .Z(n29372) );
  AND U47679 ( .A(n29373), .B(n29372), .Z(n29375) );
  NAND U47680 ( .A(n29375), .B(n29374), .Z(n29377) );
  ANDN U47681 ( .B(n29377), .A(n29376), .Z(n29378) );
  NANDN U47682 ( .A(n29379), .B(n29378), .Z(n29383) );
  AND U47683 ( .A(n29381), .B(n29380), .Z(n29382) );
  NAND U47684 ( .A(n29383), .B(n29382), .Z(n29384) );
  NANDN U47685 ( .A(n29385), .B(n29384), .Z(n29387) );
  OR U47686 ( .A(n29387), .B(n29386), .Z(n29388) );
  AND U47687 ( .A(n29389), .B(n29388), .Z(n29391) );
  NOR U47688 ( .A(n29391), .B(n29390), .Z(n29392) );
  NANDN U47689 ( .A(n29393), .B(n29392), .Z(n29394) );
  AND U47690 ( .A(n29395), .B(n29394), .Z(n29397) );
  NAND U47691 ( .A(n29397), .B(n29396), .Z(n29399) );
  ANDN U47692 ( .B(n29399), .A(n29398), .Z(n29400) );
  NANDN U47693 ( .A(n29401), .B(n29400), .Z(n29405) );
  AND U47694 ( .A(n29403), .B(n29402), .Z(n29404) );
  NAND U47695 ( .A(n29405), .B(n29404), .Z(n29406) );
  NANDN U47696 ( .A(n29407), .B(n29406), .Z(n29409) );
  OR U47697 ( .A(n29409), .B(n29408), .Z(n29410) );
  AND U47698 ( .A(n29411), .B(n29410), .Z(n29413) );
  NOR U47699 ( .A(n29413), .B(n29412), .Z(n29414) );
  NANDN U47700 ( .A(n29415), .B(n29414), .Z(n29416) );
  AND U47701 ( .A(n29417), .B(n29416), .Z(n29419) );
  NAND U47702 ( .A(n29419), .B(n29418), .Z(n29421) );
  ANDN U47703 ( .B(n29421), .A(n29420), .Z(n29422) );
  NANDN U47704 ( .A(n29423), .B(n29422), .Z(n29427) );
  AND U47705 ( .A(n29425), .B(n29424), .Z(n29426) );
  NAND U47706 ( .A(n29427), .B(n29426), .Z(n29428) );
  NANDN U47707 ( .A(n29429), .B(n29428), .Z(n29431) );
  OR U47708 ( .A(n29431), .B(n29430), .Z(n29432) );
  AND U47709 ( .A(n29433), .B(n29432), .Z(n29435) );
  NOR U47710 ( .A(n29435), .B(n29434), .Z(n29436) );
  NANDN U47711 ( .A(n29437), .B(n29436), .Z(n29438) );
  AND U47712 ( .A(n29439), .B(n29438), .Z(n29441) );
  NAND U47713 ( .A(n29441), .B(n29440), .Z(n29443) );
  ANDN U47714 ( .B(n29443), .A(n29442), .Z(n29444) );
  NANDN U47715 ( .A(n29445), .B(n29444), .Z(n29449) );
  AND U47716 ( .A(n29447), .B(n29446), .Z(n29448) );
  NAND U47717 ( .A(n29449), .B(n29448), .Z(n29450) );
  NANDN U47718 ( .A(n29451), .B(n29450), .Z(n29453) );
  OR U47719 ( .A(n29453), .B(n29452), .Z(n29454) );
  AND U47720 ( .A(n29455), .B(n29454), .Z(n29457) );
  NOR U47721 ( .A(n29457), .B(n29456), .Z(n29458) );
  NANDN U47722 ( .A(n29459), .B(n29458), .Z(n29460) );
  AND U47723 ( .A(n29461), .B(n29460), .Z(n29463) );
  NAND U47724 ( .A(n29463), .B(n29462), .Z(n29465) );
  ANDN U47725 ( .B(n29465), .A(n29464), .Z(n29466) );
  NANDN U47726 ( .A(n29467), .B(n29466), .Z(n29471) );
  AND U47727 ( .A(n29469), .B(n29468), .Z(n29470) );
  NAND U47728 ( .A(n29471), .B(n29470), .Z(n29472) );
  NANDN U47729 ( .A(n29473), .B(n29472), .Z(n29475) );
  OR U47730 ( .A(n29475), .B(n29474), .Z(n29476) );
  AND U47731 ( .A(n29477), .B(n29476), .Z(n29479) );
  NOR U47732 ( .A(n29479), .B(n29478), .Z(n29480) );
  NANDN U47733 ( .A(n29481), .B(n29480), .Z(n29482) );
  AND U47734 ( .A(n29483), .B(n29482), .Z(n29485) );
  NAND U47735 ( .A(n29485), .B(n29484), .Z(n29487) );
  ANDN U47736 ( .B(n29487), .A(n29486), .Z(n29488) );
  NANDN U47737 ( .A(n29489), .B(n29488), .Z(n29493) );
  AND U47738 ( .A(n29491), .B(n29490), .Z(n29492) );
  NAND U47739 ( .A(n29493), .B(n29492), .Z(n29494) );
  NANDN U47740 ( .A(n29495), .B(n29494), .Z(n29498) );
  NANDN U47741 ( .A(y[264]), .B(n29498), .Z(n29497) );
  ANDN U47742 ( .B(n29497), .A(n29496), .Z(n29501) );
  XNOR U47743 ( .A(n29498), .B(y[264]), .Z(n29499) );
  NAND U47744 ( .A(n29499), .B(x[264]), .Z(n29500) );
  NAND U47745 ( .A(n29501), .B(n29500), .Z(n29502) );
  NAND U47746 ( .A(n29503), .B(n29502), .Z(n29504) );
  NANDN U47747 ( .A(n29505), .B(n29504), .Z(n29506) );
  AND U47748 ( .A(n29507), .B(n29506), .Z(n29508) );
  OR U47749 ( .A(n29509), .B(n29508), .Z(n29510) );
  NAND U47750 ( .A(n29511), .B(n29510), .Z(n29512) );
  NANDN U47751 ( .A(n29513), .B(n29512), .Z(n29515) );
  NAND U47752 ( .A(n29515), .B(n29514), .Z(n29516) );
  NANDN U47753 ( .A(n29517), .B(n29516), .Z(n29518) );
  AND U47754 ( .A(n29519), .B(n29518), .Z(n29521) );
  NAND U47755 ( .A(n29521), .B(n29520), .Z(n29523) );
  ANDN U47756 ( .B(x[274]), .A(y[274]), .Z(n29522) );
  ANDN U47757 ( .B(n29523), .A(n29522), .Z(n29524) );
  NANDN U47758 ( .A(n29525), .B(n29524), .Z(n29526) );
  NAND U47759 ( .A(n29527), .B(n29526), .Z(n29528) );
  NANDN U47760 ( .A(n29529), .B(n29528), .Z(n29530) );
  AND U47761 ( .A(n29531), .B(n29530), .Z(n29533) );
  NAND U47762 ( .A(n29533), .B(n29532), .Z(n29535) );
  ANDN U47763 ( .B(n29535), .A(n29534), .Z(n29536) );
  NANDN U47764 ( .A(n29537), .B(n29536), .Z(n29541) );
  AND U47765 ( .A(n29539), .B(n29538), .Z(n29540) );
  NAND U47766 ( .A(n29541), .B(n29540), .Z(n29542) );
  NANDN U47767 ( .A(n29543), .B(n29542), .Z(n29545) );
  OR U47768 ( .A(n29545), .B(n29544), .Z(n29546) );
  AND U47769 ( .A(n29547), .B(n29546), .Z(n29549) );
  NOR U47770 ( .A(n29549), .B(n29548), .Z(n29550) );
  NANDN U47771 ( .A(n29551), .B(n29550), .Z(n29552) );
  AND U47772 ( .A(n29553), .B(n29552), .Z(n29555) );
  NAND U47773 ( .A(n29555), .B(n29554), .Z(n29557) );
  ANDN U47774 ( .B(n29557), .A(n29556), .Z(n29558) );
  NANDN U47775 ( .A(n29559), .B(n29558), .Z(n29563) );
  AND U47776 ( .A(n29561), .B(n29560), .Z(n29562) );
  NAND U47777 ( .A(n29563), .B(n29562), .Z(n29564) );
  NANDN U47778 ( .A(n29565), .B(n29564), .Z(n29567) );
  OR U47779 ( .A(n29567), .B(n29566), .Z(n29568) );
  AND U47780 ( .A(n29569), .B(n29568), .Z(n29571) );
  NOR U47781 ( .A(n29571), .B(n29570), .Z(n29572) );
  NANDN U47782 ( .A(n29573), .B(n29572), .Z(n29574) );
  AND U47783 ( .A(n29575), .B(n29574), .Z(n29577) );
  NAND U47784 ( .A(n29577), .B(n29576), .Z(n29579) );
  ANDN U47785 ( .B(n29579), .A(n29578), .Z(n29580) );
  NANDN U47786 ( .A(n29581), .B(n29580), .Z(n29585) );
  AND U47787 ( .A(n29583), .B(n29582), .Z(n29584) );
  NAND U47788 ( .A(n29585), .B(n29584), .Z(n29586) );
  NANDN U47789 ( .A(n29587), .B(n29586), .Z(n29589) );
  OR U47790 ( .A(n29589), .B(n29588), .Z(n29590) );
  AND U47791 ( .A(n29591), .B(n29590), .Z(n29593) );
  NOR U47792 ( .A(n29593), .B(n29592), .Z(n29594) );
  NANDN U47793 ( .A(n29595), .B(n29594), .Z(n29596) );
  AND U47794 ( .A(n29597), .B(n29596), .Z(n29599) );
  NAND U47795 ( .A(n29599), .B(n29598), .Z(n29601) );
  ANDN U47796 ( .B(n29601), .A(n29600), .Z(n29602) );
  NANDN U47797 ( .A(n29603), .B(n29602), .Z(n29607) );
  AND U47798 ( .A(n29605), .B(n29604), .Z(n29606) );
  NAND U47799 ( .A(n29607), .B(n29606), .Z(n29608) );
  NANDN U47800 ( .A(n29609), .B(n29608), .Z(n29611) );
  OR U47801 ( .A(n29611), .B(n29610), .Z(n29612) );
  AND U47802 ( .A(n29613), .B(n29612), .Z(n29615) );
  NOR U47803 ( .A(n29615), .B(n29614), .Z(n29616) );
  NANDN U47804 ( .A(n29617), .B(n29616), .Z(n29618) );
  AND U47805 ( .A(n29619), .B(n29618), .Z(n29621) );
  NAND U47806 ( .A(n29621), .B(n29620), .Z(n29623) );
  ANDN U47807 ( .B(n29623), .A(n29622), .Z(n29624) );
  NANDN U47808 ( .A(n29625), .B(n29624), .Z(n29629) );
  AND U47809 ( .A(n29627), .B(n29626), .Z(n29628) );
  NAND U47810 ( .A(n29629), .B(n29628), .Z(n29630) );
  NANDN U47811 ( .A(n29631), .B(n29630), .Z(n29633) );
  OR U47812 ( .A(n29633), .B(n29632), .Z(n29634) );
  AND U47813 ( .A(n29635), .B(n29634), .Z(n29637) );
  NOR U47814 ( .A(n29637), .B(n29636), .Z(n29638) );
  NANDN U47815 ( .A(n29639), .B(n29638), .Z(n29640) );
  AND U47816 ( .A(n29641), .B(n29640), .Z(n29643) );
  NAND U47817 ( .A(n29643), .B(n29642), .Z(n29645) );
  ANDN U47818 ( .B(n29645), .A(n29644), .Z(n29646) );
  NANDN U47819 ( .A(n29647), .B(n29646), .Z(n29651) );
  AND U47820 ( .A(n29649), .B(n29648), .Z(n29650) );
  NAND U47821 ( .A(n29651), .B(n29650), .Z(n29652) );
  NANDN U47822 ( .A(n29653), .B(n29652), .Z(n29655) );
  OR U47823 ( .A(n29655), .B(n29654), .Z(n29656) );
  AND U47824 ( .A(n29657), .B(n29656), .Z(n29659) );
  NOR U47825 ( .A(n29659), .B(n29658), .Z(n29660) );
  NANDN U47826 ( .A(n29661), .B(n29660), .Z(n29662) );
  AND U47827 ( .A(n29663), .B(n29662), .Z(n29665) );
  NAND U47828 ( .A(n29665), .B(n29664), .Z(n29667) );
  ANDN U47829 ( .B(n29667), .A(n29666), .Z(n29668) );
  NANDN U47830 ( .A(n29669), .B(n29668), .Z(n29673) );
  AND U47831 ( .A(n29671), .B(n29670), .Z(n29672) );
  NAND U47832 ( .A(n29673), .B(n29672), .Z(n29674) );
  NANDN U47833 ( .A(n29675), .B(n29674), .Z(n29677) );
  OR U47834 ( .A(n29677), .B(n29676), .Z(n29678) );
  AND U47835 ( .A(n29679), .B(n29678), .Z(n29681) );
  NOR U47836 ( .A(n29681), .B(n29680), .Z(n29682) );
  NANDN U47837 ( .A(n29683), .B(n29682), .Z(n29684) );
  AND U47838 ( .A(n29685), .B(n29684), .Z(n29687) );
  NAND U47839 ( .A(n29687), .B(n29686), .Z(n29689) );
  ANDN U47840 ( .B(n29689), .A(n29688), .Z(n29690) );
  NANDN U47841 ( .A(n29691), .B(n29690), .Z(n29695) );
  AND U47842 ( .A(n29693), .B(n29692), .Z(n29694) );
  NAND U47843 ( .A(n29695), .B(n29694), .Z(n29696) );
  NANDN U47844 ( .A(n29697), .B(n29696), .Z(n29699) );
  OR U47845 ( .A(n29699), .B(n29698), .Z(n29700) );
  AND U47846 ( .A(n29701), .B(n29700), .Z(n29703) );
  NOR U47847 ( .A(n29703), .B(n29702), .Z(n29704) );
  NANDN U47848 ( .A(n29705), .B(n29704), .Z(n29706) );
  AND U47849 ( .A(n29707), .B(n29706), .Z(n29709) );
  NAND U47850 ( .A(n29709), .B(n29708), .Z(n29711) );
  ANDN U47851 ( .B(n29711), .A(n29710), .Z(n29712) );
  NANDN U47852 ( .A(n29713), .B(n29712), .Z(n29717) );
  AND U47853 ( .A(n29715), .B(n29714), .Z(n29716) );
  NAND U47854 ( .A(n29717), .B(n29716), .Z(n29718) );
  NANDN U47855 ( .A(n29719), .B(n29718), .Z(n29721) );
  OR U47856 ( .A(n29721), .B(n29720), .Z(n29722) );
  AND U47857 ( .A(n29723), .B(n29722), .Z(n29725) );
  NOR U47858 ( .A(n29725), .B(n29724), .Z(n29726) );
  NANDN U47859 ( .A(n29727), .B(n29726), .Z(n29728) );
  AND U47860 ( .A(n29729), .B(n29728), .Z(n29731) );
  NAND U47861 ( .A(n29731), .B(n29730), .Z(n29733) );
  ANDN U47862 ( .B(n29733), .A(n29732), .Z(n29734) );
  NANDN U47863 ( .A(n29735), .B(n29734), .Z(n29739) );
  AND U47864 ( .A(n29737), .B(n29736), .Z(n29738) );
  NAND U47865 ( .A(n29739), .B(n29738), .Z(n29740) );
  NANDN U47866 ( .A(n29741), .B(n29740), .Z(n29743) );
  OR U47867 ( .A(n29743), .B(n29742), .Z(n29744) );
  AND U47868 ( .A(n29745), .B(n29744), .Z(n29747) );
  NOR U47869 ( .A(n29747), .B(n29746), .Z(n29748) );
  NANDN U47870 ( .A(n29749), .B(n29748), .Z(n29750) );
  AND U47871 ( .A(n29751), .B(n29750), .Z(n29753) );
  NAND U47872 ( .A(n29753), .B(n29752), .Z(n29755) );
  ANDN U47873 ( .B(n29755), .A(n29754), .Z(n29756) );
  NANDN U47874 ( .A(n29757), .B(n29756), .Z(n29758) );
  AND U47875 ( .A(n29759), .B(n29758), .Z(n29760) );
  NAND U47876 ( .A(n29761), .B(n29760), .Z(n29762) );
  NANDN U47877 ( .A(n29763), .B(n29762), .Z(n29765) );
  OR U47878 ( .A(n29765), .B(n29764), .Z(n29766) );
  AND U47879 ( .A(n29767), .B(n29766), .Z(n29769) );
  NOR U47880 ( .A(n29769), .B(n29768), .Z(n29770) );
  NANDN U47881 ( .A(n29771), .B(n29770), .Z(n29772) );
  AND U47882 ( .A(n29773), .B(n29772), .Z(n29775) );
  NAND U47883 ( .A(n29775), .B(n29774), .Z(n29777) );
  ANDN U47884 ( .B(n29777), .A(n29776), .Z(n29778) );
  NANDN U47885 ( .A(n29779), .B(n29778), .Z(n29783) );
  AND U47886 ( .A(n29781), .B(n29780), .Z(n29782) );
  NAND U47887 ( .A(n29783), .B(n29782), .Z(n29784) );
  NANDN U47888 ( .A(n29785), .B(n29784), .Z(n29787) );
  OR U47889 ( .A(n29787), .B(n29786), .Z(n29788) );
  AND U47890 ( .A(n29789), .B(n29788), .Z(n29791) );
  NOR U47891 ( .A(n29791), .B(n29790), .Z(n29792) );
  NANDN U47892 ( .A(n29793), .B(n29792), .Z(n29794) );
  AND U47893 ( .A(n29795), .B(n29794), .Z(n29797) );
  NAND U47894 ( .A(n29797), .B(n29796), .Z(n29799) );
  ANDN U47895 ( .B(n29799), .A(n29798), .Z(n29800) );
  NANDN U47896 ( .A(n29801), .B(n29800), .Z(n29802) );
  AND U47897 ( .A(n29803), .B(n29802), .Z(n29804) );
  NAND U47898 ( .A(n29805), .B(n29804), .Z(n29806) );
  NANDN U47899 ( .A(n29807), .B(n29806), .Z(n29809) );
  OR U47900 ( .A(n29809), .B(n29808), .Z(n29810) );
  AND U47901 ( .A(n29811), .B(n29810), .Z(n29813) );
  NOR U47902 ( .A(n29813), .B(n29812), .Z(n29814) );
  NANDN U47903 ( .A(n29815), .B(n29814), .Z(n29816) );
  AND U47904 ( .A(n29817), .B(n29816), .Z(n29819) );
  NAND U47905 ( .A(n29819), .B(n29818), .Z(n29821) );
  ANDN U47906 ( .B(n29821), .A(n29820), .Z(n29822) );
  NANDN U47907 ( .A(n29823), .B(n29822), .Z(n29827) );
  AND U47908 ( .A(n29825), .B(n29824), .Z(n29826) );
  NAND U47909 ( .A(n29827), .B(n29826), .Z(n29828) );
  NANDN U47910 ( .A(n29829), .B(n29828), .Z(n29831) );
  OR U47911 ( .A(n29831), .B(n29830), .Z(n29832) );
  AND U47912 ( .A(n29833), .B(n29832), .Z(n29835) );
  NOR U47913 ( .A(n29835), .B(n29834), .Z(n29836) );
  NANDN U47914 ( .A(n29837), .B(n29836), .Z(n29838) );
  AND U47915 ( .A(n29839), .B(n29838), .Z(n29841) );
  NAND U47916 ( .A(n29841), .B(n29840), .Z(n29843) );
  ANDN U47917 ( .B(n29843), .A(n29842), .Z(n29844) );
  NANDN U47918 ( .A(n29845), .B(n29844), .Z(n29846) );
  AND U47919 ( .A(n29847), .B(n29846), .Z(n29848) );
  NAND U47920 ( .A(n29849), .B(n29848), .Z(n29850) );
  NANDN U47921 ( .A(n29851), .B(n29850), .Z(n29853) );
  OR U47922 ( .A(n29853), .B(n29852), .Z(n29854) );
  AND U47923 ( .A(n29855), .B(n29854), .Z(n29857) );
  NOR U47924 ( .A(n29857), .B(n29856), .Z(n29858) );
  NANDN U47925 ( .A(n29859), .B(n29858), .Z(n29860) );
  AND U47926 ( .A(n29861), .B(n29860), .Z(n29863) );
  NAND U47927 ( .A(n29863), .B(n29862), .Z(n29865) );
  ANDN U47928 ( .B(n29865), .A(n29864), .Z(n29866) );
  NANDN U47929 ( .A(n29867), .B(n29866), .Z(n29871) );
  AND U47930 ( .A(n29869), .B(n29868), .Z(n29870) );
  NAND U47931 ( .A(n29871), .B(n29870), .Z(n29872) );
  NANDN U47932 ( .A(n29873), .B(n29872), .Z(n29875) );
  OR U47933 ( .A(n29875), .B(n29874), .Z(n29876) );
  AND U47934 ( .A(n29877), .B(n29876), .Z(n29879) );
  NOR U47935 ( .A(n29879), .B(n29878), .Z(n29880) );
  NANDN U47936 ( .A(n29881), .B(n29880), .Z(n29882) );
  AND U47937 ( .A(n29883), .B(n29882), .Z(n29885) );
  NAND U47938 ( .A(n29885), .B(n29884), .Z(n29887) );
  ANDN U47939 ( .B(n29887), .A(n29886), .Z(n29888) );
  NANDN U47940 ( .A(n29889), .B(n29888), .Z(n29893) );
  AND U47941 ( .A(n29891), .B(n29890), .Z(n29892) );
  NAND U47942 ( .A(n29893), .B(n29892), .Z(n29894) );
  NANDN U47943 ( .A(n29895), .B(n29894), .Z(n29897) );
  OR U47944 ( .A(n29897), .B(n29896), .Z(n29898) );
  AND U47945 ( .A(n29899), .B(n29898), .Z(n29901) );
  NOR U47946 ( .A(n29901), .B(n29900), .Z(n29902) );
  NANDN U47947 ( .A(n29903), .B(n29902), .Z(n29904) );
  AND U47948 ( .A(n29905), .B(n29904), .Z(n29907) );
  NAND U47949 ( .A(n29907), .B(n29906), .Z(n29909) );
  ANDN U47950 ( .B(n29909), .A(n29908), .Z(n29910) );
  NANDN U47951 ( .A(n29911), .B(n29910), .Z(n29915) );
  AND U47952 ( .A(n29913), .B(n29912), .Z(n29914) );
  NAND U47953 ( .A(n29915), .B(n29914), .Z(n29916) );
  NANDN U47954 ( .A(n29917), .B(n29916), .Z(n29919) );
  OR U47955 ( .A(n29919), .B(n29918), .Z(n29920) );
  AND U47956 ( .A(n29921), .B(n29920), .Z(n29923) );
  NOR U47957 ( .A(n29923), .B(n29922), .Z(n29924) );
  NANDN U47958 ( .A(n29925), .B(n29924), .Z(n29926) );
  AND U47959 ( .A(n29927), .B(n29926), .Z(n29929) );
  NAND U47960 ( .A(n29929), .B(n29928), .Z(n29931) );
  ANDN U47961 ( .B(n29931), .A(n29930), .Z(n29932) );
  NANDN U47962 ( .A(n29933), .B(n29932), .Z(n29937) );
  AND U47963 ( .A(n29935), .B(n29934), .Z(n29936) );
  NAND U47964 ( .A(n29937), .B(n29936), .Z(n29938) );
  NANDN U47965 ( .A(n29939), .B(n29938), .Z(n29941) );
  OR U47966 ( .A(n29941), .B(n29940), .Z(n29942) );
  AND U47967 ( .A(n29943), .B(n29942), .Z(n29945) );
  NOR U47968 ( .A(n29945), .B(n29944), .Z(n29946) );
  NANDN U47969 ( .A(n29947), .B(n29946), .Z(n29948) );
  AND U47970 ( .A(n29949), .B(n29948), .Z(n29951) );
  NAND U47971 ( .A(n29951), .B(n29950), .Z(n29953) );
  ANDN U47972 ( .B(n29953), .A(n29952), .Z(n29954) );
  NANDN U47973 ( .A(n29955), .B(n29954), .Z(n29959) );
  AND U47974 ( .A(n29957), .B(n29956), .Z(n29958) );
  NAND U47975 ( .A(n29959), .B(n29958), .Z(n29960) );
  NANDN U47976 ( .A(n29961), .B(n29960), .Z(n29963) );
  OR U47977 ( .A(n29963), .B(n29962), .Z(n29964) );
  AND U47978 ( .A(n29965), .B(n29964), .Z(n29967) );
  NOR U47979 ( .A(n29967), .B(n29966), .Z(n29968) );
  NANDN U47980 ( .A(n29969), .B(n29968), .Z(n29970) );
  AND U47981 ( .A(n29971), .B(n29970), .Z(n29973) );
  NAND U47982 ( .A(n29973), .B(n29972), .Z(n29975) );
  ANDN U47983 ( .B(n29975), .A(n29974), .Z(n29976) );
  NANDN U47984 ( .A(n29977), .B(n29976), .Z(n29981) );
  AND U47985 ( .A(n29979), .B(n29978), .Z(n29980) );
  NAND U47986 ( .A(n29981), .B(n29980), .Z(n29982) );
  NANDN U47987 ( .A(n29983), .B(n29982), .Z(n29985) );
  OR U47988 ( .A(n29985), .B(n29984), .Z(n29986) );
  AND U47989 ( .A(n29987), .B(n29986), .Z(n29989) );
  NOR U47990 ( .A(n29989), .B(n29988), .Z(n29990) );
  NANDN U47991 ( .A(n29991), .B(n29990), .Z(n29992) );
  AND U47992 ( .A(n29993), .B(n29992), .Z(n29995) );
  NAND U47993 ( .A(n29995), .B(n29994), .Z(n29997) );
  ANDN U47994 ( .B(n29997), .A(n29996), .Z(n29998) );
  NANDN U47995 ( .A(n29999), .B(n29998), .Z(n30003) );
  AND U47996 ( .A(n30001), .B(n30000), .Z(n30002) );
  NAND U47997 ( .A(n30003), .B(n30002), .Z(n30004) );
  NANDN U47998 ( .A(n30005), .B(n30004), .Z(n30007) );
  OR U47999 ( .A(n30007), .B(n30006), .Z(n30008) );
  AND U48000 ( .A(n30009), .B(n30008), .Z(n30011) );
  NOR U48001 ( .A(n30011), .B(n30010), .Z(n30012) );
  NANDN U48002 ( .A(n30013), .B(n30012), .Z(n30014) );
  AND U48003 ( .A(n30015), .B(n30014), .Z(n30017) );
  NAND U48004 ( .A(n30017), .B(n30016), .Z(n30019) );
  ANDN U48005 ( .B(n30019), .A(n30018), .Z(n30020) );
  NANDN U48006 ( .A(n30021), .B(n30020), .Z(n30025) );
  AND U48007 ( .A(n30023), .B(n30022), .Z(n30024) );
  NAND U48008 ( .A(n30025), .B(n30024), .Z(n30026) );
  NANDN U48009 ( .A(n30027), .B(n30026), .Z(n30029) );
  OR U48010 ( .A(n30029), .B(n30028), .Z(n30030) );
  AND U48011 ( .A(n30031), .B(n30030), .Z(n30033) );
  NOR U48012 ( .A(n30033), .B(n30032), .Z(n30034) );
  NANDN U48013 ( .A(n30035), .B(n30034), .Z(n30036) );
  AND U48014 ( .A(n30037), .B(n30036), .Z(n30039) );
  NAND U48015 ( .A(n30039), .B(n30038), .Z(n30041) );
  ANDN U48016 ( .B(n30041), .A(n30040), .Z(n30042) );
  NANDN U48017 ( .A(n30043), .B(n30042), .Z(n30047) );
  AND U48018 ( .A(n30045), .B(n30044), .Z(n30046) );
  NAND U48019 ( .A(n30047), .B(n30046), .Z(n30048) );
  NANDN U48020 ( .A(n30049), .B(n30048), .Z(n30051) );
  OR U48021 ( .A(n30051), .B(n30050), .Z(n30052) );
  AND U48022 ( .A(n30053), .B(n30052), .Z(n30055) );
  NOR U48023 ( .A(n30055), .B(n30054), .Z(n30056) );
  NANDN U48024 ( .A(n30057), .B(n30056), .Z(n30058) );
  AND U48025 ( .A(n30059), .B(n30058), .Z(n30061) );
  NAND U48026 ( .A(n30061), .B(n30060), .Z(n30063) );
  ANDN U48027 ( .B(n30063), .A(n30062), .Z(n30064) );
  NANDN U48028 ( .A(n30065), .B(n30064), .Z(n30069) );
  AND U48029 ( .A(n30067), .B(n30066), .Z(n30068) );
  NAND U48030 ( .A(n30069), .B(n30068), .Z(n30070) );
  NANDN U48031 ( .A(n30071), .B(n30070), .Z(n30073) );
  OR U48032 ( .A(n30073), .B(n30072), .Z(n30074) );
  AND U48033 ( .A(n30075), .B(n30074), .Z(n30077) );
  NOR U48034 ( .A(n30077), .B(n30076), .Z(n30078) );
  NANDN U48035 ( .A(n30079), .B(n30078), .Z(n30080) );
  AND U48036 ( .A(n30081), .B(n30080), .Z(n30083) );
  NAND U48037 ( .A(n30083), .B(n30082), .Z(n30085) );
  ANDN U48038 ( .B(n30085), .A(n30084), .Z(n30086) );
  NANDN U48039 ( .A(n30087), .B(n30086), .Z(n30091) );
  AND U48040 ( .A(n30089), .B(n30088), .Z(n30090) );
  NAND U48041 ( .A(n30091), .B(n30090), .Z(n30092) );
  NANDN U48042 ( .A(n30093), .B(n30092), .Z(n30095) );
  OR U48043 ( .A(n30095), .B(n30094), .Z(n30096) );
  AND U48044 ( .A(n30097), .B(n30096), .Z(n30098) );
  NOR U48045 ( .A(n30099), .B(n30098), .Z(n30100) );
  NANDN U48046 ( .A(n30101), .B(n30100), .Z(n30102) );
  AND U48047 ( .A(n30103), .B(n30102), .Z(n30105) );
  NANDN U48048 ( .A(x[432]), .B(y[432]), .Z(n30104) );
  NAND U48049 ( .A(n30105), .B(n30104), .Z(n30107) );
  ANDN U48050 ( .B(n30107), .A(n30106), .Z(n30108) );
  NANDN U48051 ( .A(n30109), .B(n30108), .Z(n30113) );
  AND U48052 ( .A(n30111), .B(n30110), .Z(n30112) );
  NAND U48053 ( .A(n30113), .B(n30112), .Z(n30114) );
  NANDN U48054 ( .A(n30115), .B(n30114), .Z(n30117) );
  OR U48055 ( .A(n30117), .B(n30116), .Z(n30118) );
  AND U48056 ( .A(n30119), .B(n30118), .Z(n30121) );
  NOR U48057 ( .A(n30121), .B(n30120), .Z(n30122) );
  NANDN U48058 ( .A(n30123), .B(n30122), .Z(n30124) );
  AND U48059 ( .A(n30125), .B(n30124), .Z(n30127) );
  NAND U48060 ( .A(n30127), .B(n30126), .Z(n30129) );
  ANDN U48061 ( .B(n30129), .A(n30128), .Z(n30130) );
  NANDN U48062 ( .A(n30131), .B(n30130), .Z(n30135) );
  AND U48063 ( .A(n30133), .B(n30132), .Z(n30134) );
  NAND U48064 ( .A(n30135), .B(n30134), .Z(n30136) );
  NANDN U48065 ( .A(n30137), .B(n30136), .Z(n30139) );
  OR U48066 ( .A(n30139), .B(n30138), .Z(n30140) );
  AND U48067 ( .A(n30141), .B(n30140), .Z(n30143) );
  NOR U48068 ( .A(n30143), .B(n30142), .Z(n30144) );
  NANDN U48069 ( .A(n30145), .B(n30144), .Z(n30146) );
  AND U48070 ( .A(n30147), .B(n30146), .Z(n30149) );
  NAND U48071 ( .A(n30149), .B(n30148), .Z(n30151) );
  ANDN U48072 ( .B(n30151), .A(n30150), .Z(n30152) );
  NANDN U48073 ( .A(n30153), .B(n30152), .Z(n30157) );
  AND U48074 ( .A(n30155), .B(n30154), .Z(n30156) );
  NAND U48075 ( .A(n30157), .B(n30156), .Z(n30158) );
  NANDN U48076 ( .A(n30159), .B(n30158), .Z(n30161) );
  OR U48077 ( .A(n30161), .B(n30160), .Z(n30162) );
  AND U48078 ( .A(n30163), .B(n30162), .Z(n30165) );
  NOR U48079 ( .A(n30165), .B(n30164), .Z(n30166) );
  NANDN U48080 ( .A(n30167), .B(n30166), .Z(n30168) );
  AND U48081 ( .A(n30169), .B(n30168), .Z(n30171) );
  NAND U48082 ( .A(n30171), .B(n30170), .Z(n30173) );
  ANDN U48083 ( .B(n30173), .A(n30172), .Z(n30174) );
  NANDN U48084 ( .A(n30175), .B(n30174), .Z(n30179) );
  AND U48085 ( .A(n30177), .B(n30176), .Z(n30178) );
  NAND U48086 ( .A(n30179), .B(n30178), .Z(n30180) );
  NANDN U48087 ( .A(n30181), .B(n30180), .Z(n30183) );
  OR U48088 ( .A(n30183), .B(n30182), .Z(n30184) );
  AND U48089 ( .A(n30185), .B(n30184), .Z(n30187) );
  NOR U48090 ( .A(n30187), .B(n30186), .Z(n30188) );
  NANDN U48091 ( .A(n30189), .B(n30188), .Z(n30190) );
  AND U48092 ( .A(n30191), .B(n30190), .Z(n30193) );
  NAND U48093 ( .A(n30193), .B(n30192), .Z(n30195) );
  ANDN U48094 ( .B(n30195), .A(n30194), .Z(n30196) );
  NANDN U48095 ( .A(n30197), .B(n30196), .Z(n30201) );
  AND U48096 ( .A(n30199), .B(n30198), .Z(n30200) );
  NAND U48097 ( .A(n30201), .B(n30200), .Z(n30202) );
  NANDN U48098 ( .A(n30203), .B(n30202), .Z(n30205) );
  OR U48099 ( .A(n30205), .B(n30204), .Z(n30206) );
  AND U48100 ( .A(n30207), .B(n30206), .Z(n30209) );
  NOR U48101 ( .A(n30209), .B(n30208), .Z(n30210) );
  NANDN U48102 ( .A(n30211), .B(n30210), .Z(n30212) );
  AND U48103 ( .A(n30213), .B(n30212), .Z(n30215) );
  NAND U48104 ( .A(n30215), .B(n30214), .Z(n30217) );
  ANDN U48105 ( .B(n30217), .A(n30216), .Z(n30218) );
  NANDN U48106 ( .A(n30219), .B(n30218), .Z(n30223) );
  AND U48107 ( .A(n30221), .B(n30220), .Z(n30222) );
  NAND U48108 ( .A(n30223), .B(n30222), .Z(n30224) );
  NANDN U48109 ( .A(n30225), .B(n30224), .Z(n30227) );
  OR U48110 ( .A(n30227), .B(n30226), .Z(n30228) );
  AND U48111 ( .A(n30229), .B(n30228), .Z(n30231) );
  NOR U48112 ( .A(n30231), .B(n30230), .Z(n30232) );
  NANDN U48113 ( .A(n30233), .B(n30232), .Z(n30234) );
  AND U48114 ( .A(n30235), .B(n30234), .Z(n30237) );
  NAND U48115 ( .A(n30237), .B(n30236), .Z(n30239) );
  ANDN U48116 ( .B(n30239), .A(n30238), .Z(n30240) );
  NANDN U48117 ( .A(n30241), .B(n30240), .Z(n30245) );
  AND U48118 ( .A(n30243), .B(n30242), .Z(n30244) );
  NAND U48119 ( .A(n30245), .B(n30244), .Z(n30246) );
  NANDN U48120 ( .A(n30247), .B(n30246), .Z(n30249) );
  OR U48121 ( .A(n30249), .B(n30248), .Z(n30250) );
  AND U48122 ( .A(n30251), .B(n30250), .Z(n30253) );
  NOR U48123 ( .A(n30253), .B(n30252), .Z(n30254) );
  NANDN U48124 ( .A(n30255), .B(n30254), .Z(n30256) );
  AND U48125 ( .A(n30257), .B(n30256), .Z(n30259) );
  NAND U48126 ( .A(n30259), .B(n30258), .Z(n30261) );
  ANDN U48127 ( .B(n30261), .A(n30260), .Z(n30262) );
  NANDN U48128 ( .A(n30263), .B(n30262), .Z(n30267) );
  AND U48129 ( .A(n30265), .B(n30264), .Z(n30266) );
  NAND U48130 ( .A(n30267), .B(n30266), .Z(n30268) );
  NANDN U48131 ( .A(n30269), .B(n30268), .Z(n30271) );
  OR U48132 ( .A(n30271), .B(n30270), .Z(n30272) );
  AND U48133 ( .A(n30273), .B(n30272), .Z(n30275) );
  NOR U48134 ( .A(n30275), .B(n30274), .Z(n30276) );
  NANDN U48135 ( .A(n30277), .B(n30276), .Z(n30278) );
  AND U48136 ( .A(n30279), .B(n30278), .Z(n30281) );
  NAND U48137 ( .A(n30281), .B(n30280), .Z(n30283) );
  ANDN U48138 ( .B(n30283), .A(n30282), .Z(n30284) );
  NANDN U48139 ( .A(n30285), .B(n30284), .Z(n30289) );
  AND U48140 ( .A(n30287), .B(n30286), .Z(n30288) );
  NAND U48141 ( .A(n30289), .B(n30288), .Z(n30290) );
  NANDN U48142 ( .A(n30291), .B(n30290), .Z(n30293) );
  OR U48143 ( .A(n30293), .B(n30292), .Z(n30294) );
  AND U48144 ( .A(n30295), .B(n30294), .Z(n30297) );
  NOR U48145 ( .A(n30297), .B(n30296), .Z(n30298) );
  NANDN U48146 ( .A(n30299), .B(n30298), .Z(n30300) );
  AND U48147 ( .A(n30301), .B(n30300), .Z(n30303) );
  NAND U48148 ( .A(n30303), .B(n30302), .Z(n30305) );
  ANDN U48149 ( .B(n30305), .A(n30304), .Z(n30306) );
  NANDN U48150 ( .A(n30307), .B(n30306), .Z(n30311) );
  AND U48151 ( .A(n30309), .B(n30308), .Z(n30310) );
  NAND U48152 ( .A(n30311), .B(n30310), .Z(n30312) );
  NANDN U48153 ( .A(n30313), .B(n30312), .Z(n30315) );
  OR U48154 ( .A(n30315), .B(n30314), .Z(n30316) );
  AND U48155 ( .A(n30317), .B(n30316), .Z(n30319) );
  NOR U48156 ( .A(n30319), .B(n30318), .Z(n30320) );
  NANDN U48157 ( .A(n30321), .B(n30320), .Z(n30322) );
  AND U48158 ( .A(n30323), .B(n30322), .Z(n30325) );
  NAND U48159 ( .A(n30325), .B(n30324), .Z(n30327) );
  ANDN U48160 ( .B(n30327), .A(n30326), .Z(n30328) );
  NANDN U48161 ( .A(n30329), .B(n30328), .Z(n30333) );
  AND U48162 ( .A(n30331), .B(n30330), .Z(n30332) );
  NAND U48163 ( .A(n30333), .B(n30332), .Z(n30334) );
  NANDN U48164 ( .A(n30335), .B(n30334), .Z(n30337) );
  OR U48165 ( .A(n30337), .B(n30336), .Z(n30338) );
  AND U48166 ( .A(n30339), .B(n30338), .Z(n30341) );
  NOR U48167 ( .A(n30341), .B(n30340), .Z(n30342) );
  NANDN U48168 ( .A(n30343), .B(n30342), .Z(n30344) );
  AND U48169 ( .A(n30345), .B(n30344), .Z(n30347) );
  NAND U48170 ( .A(n30347), .B(n30346), .Z(n30349) );
  ANDN U48171 ( .B(n30349), .A(n30348), .Z(n30350) );
  NANDN U48172 ( .A(n30351), .B(n30350), .Z(n30355) );
  AND U48173 ( .A(n30353), .B(n30352), .Z(n30354) );
  NAND U48174 ( .A(n30355), .B(n30354), .Z(n30356) );
  NANDN U48175 ( .A(n30357), .B(n30356), .Z(n30359) );
  OR U48176 ( .A(n30359), .B(n30358), .Z(n30360) );
  AND U48177 ( .A(n30361), .B(n30360), .Z(n30363) );
  NOR U48178 ( .A(n30363), .B(n30362), .Z(n30364) );
  NANDN U48179 ( .A(n30365), .B(n30364), .Z(n30366) );
  AND U48180 ( .A(n30367), .B(n30366), .Z(n30369) );
  NAND U48181 ( .A(n30369), .B(n30368), .Z(n30371) );
  ANDN U48182 ( .B(n30371), .A(n30370), .Z(n30372) );
  NANDN U48183 ( .A(n30373), .B(n30372), .Z(n30377) );
  AND U48184 ( .A(n30375), .B(n30374), .Z(n30376) );
  NAND U48185 ( .A(n30377), .B(n30376), .Z(n30378) );
  NANDN U48186 ( .A(n30379), .B(n30378), .Z(n30381) );
  OR U48187 ( .A(n30381), .B(n30380), .Z(n30382) );
  AND U48188 ( .A(n30383), .B(n30382), .Z(n30385) );
  NOR U48189 ( .A(n30385), .B(n30384), .Z(n30386) );
  NANDN U48190 ( .A(n30387), .B(n30386), .Z(n30388) );
  AND U48191 ( .A(n30389), .B(n30388), .Z(n30391) );
  NAND U48192 ( .A(n30391), .B(n30390), .Z(n30393) );
  ANDN U48193 ( .B(n30393), .A(n30392), .Z(n30394) );
  NANDN U48194 ( .A(n30395), .B(n30394), .Z(n30399) );
  AND U48195 ( .A(n30397), .B(n30396), .Z(n30398) );
  NAND U48196 ( .A(n30399), .B(n30398), .Z(n30400) );
  NANDN U48197 ( .A(n30401), .B(n30400), .Z(n30403) );
  OR U48198 ( .A(n30403), .B(n30402), .Z(n30404) );
  AND U48199 ( .A(n30405), .B(n30404), .Z(n30407) );
  NOR U48200 ( .A(n30407), .B(n30406), .Z(n30408) );
  NANDN U48201 ( .A(n30409), .B(n30408), .Z(n30410) );
  AND U48202 ( .A(n30411), .B(n30410), .Z(n30413) );
  NAND U48203 ( .A(n30413), .B(n30412), .Z(n30415) );
  ANDN U48204 ( .B(n30415), .A(n30414), .Z(n30416) );
  NANDN U48205 ( .A(n30417), .B(n30416), .Z(n30421) );
  AND U48206 ( .A(n30419), .B(n30418), .Z(n30420) );
  NAND U48207 ( .A(n30421), .B(n30420), .Z(n30422) );
  NANDN U48208 ( .A(n30423), .B(n30422), .Z(n30425) );
  OR U48209 ( .A(n30425), .B(n30424), .Z(n30426) );
  AND U48210 ( .A(n30427), .B(n30426), .Z(n30429) );
  NOR U48211 ( .A(n30429), .B(n30428), .Z(n30430) );
  NANDN U48212 ( .A(n30431), .B(n30430), .Z(n30432) );
  AND U48213 ( .A(n30433), .B(n30432), .Z(n30435) );
  NAND U48214 ( .A(n30435), .B(n30434), .Z(n30437) );
  ANDN U48215 ( .B(n30437), .A(n30436), .Z(n30438) );
  NANDN U48216 ( .A(n30439), .B(n30438), .Z(n30443) );
  AND U48217 ( .A(n30441), .B(n30440), .Z(n30442) );
  NAND U48218 ( .A(n30443), .B(n30442), .Z(n30444) );
  NANDN U48219 ( .A(n30445), .B(n30444), .Z(n30448) );
  NANDN U48220 ( .A(y[526]), .B(n30448), .Z(n30447) );
  ANDN U48221 ( .B(n30447), .A(n30446), .Z(n30451) );
  XNOR U48222 ( .A(n30448), .B(y[526]), .Z(n30449) );
  NAND U48223 ( .A(n30449), .B(x[526]), .Z(n30450) );
  NAND U48224 ( .A(n30451), .B(n30450), .Z(n30452) );
  NAND U48225 ( .A(n30453), .B(n30452), .Z(n30454) );
  NANDN U48226 ( .A(n30455), .B(n30454), .Z(n30456) );
  AND U48227 ( .A(n30457), .B(n30456), .Z(n30458) );
  OR U48228 ( .A(n30459), .B(n30458), .Z(n30460) );
  NAND U48229 ( .A(n30461), .B(n30460), .Z(n30462) );
  NANDN U48230 ( .A(n30463), .B(n30462), .Z(n30464) );
  NAND U48231 ( .A(n30465), .B(n30464), .Z(n30466) );
  NANDN U48232 ( .A(n30467), .B(n30466), .Z(n30468) );
  AND U48233 ( .A(n30469), .B(n30468), .Z(n30470) );
  OR U48234 ( .A(n30471), .B(n30470), .Z(n30472) );
  NAND U48235 ( .A(n30473), .B(n30472), .Z(n30474) );
  NANDN U48236 ( .A(n30475), .B(n30474), .Z(n30479) );
  AND U48237 ( .A(n30477), .B(n30476), .Z(n30478) );
  NAND U48238 ( .A(n30479), .B(n30478), .Z(n30480) );
  NANDN U48239 ( .A(n30481), .B(n30480), .Z(n30483) );
  OR U48240 ( .A(n30483), .B(n30482), .Z(n30484) );
  AND U48241 ( .A(n30485), .B(n30484), .Z(n30486) );
  NOR U48242 ( .A(n30487), .B(n30486), .Z(n30488) );
  NANDN U48243 ( .A(n30489), .B(n30488), .Z(n30490) );
  AND U48244 ( .A(n30491), .B(n30490), .Z(n30493) );
  NANDN U48245 ( .A(x[542]), .B(y[542]), .Z(n30492) );
  NAND U48246 ( .A(n30493), .B(n30492), .Z(n30495) );
  ANDN U48247 ( .B(n30495), .A(n30494), .Z(n30496) );
  NANDN U48248 ( .A(n30497), .B(n30496), .Z(n30501) );
  AND U48249 ( .A(n30499), .B(n30498), .Z(n30500) );
  NAND U48250 ( .A(n30501), .B(n30500), .Z(n30502) );
  NANDN U48251 ( .A(n30503), .B(n30502), .Z(n30505) );
  OR U48252 ( .A(n30505), .B(n30504), .Z(n30506) );
  AND U48253 ( .A(n30507), .B(n30506), .Z(n30508) );
  NOR U48254 ( .A(n30509), .B(n30508), .Z(n30510) );
  NANDN U48255 ( .A(n30511), .B(n30510), .Z(n30512) );
  AND U48256 ( .A(n30513), .B(n30512), .Z(n30515) );
  NANDN U48257 ( .A(n30515), .B(n30514), .Z(n30516) );
  NANDN U48258 ( .A(n52438), .B(n30516), .Z(n30517) );
  AND U48259 ( .A(n52440), .B(n30517), .Z(n30518) );
  NOR U48260 ( .A(n52441), .B(n30518), .Z(n30519) );
  NANDN U48261 ( .A(n30520), .B(n30519), .Z(n30521) );
  AND U48262 ( .A(n30522), .B(n30521), .Z(n30523) );
  NOR U48263 ( .A(n52446), .B(n30523), .Z(n30524) );
  NANDN U48264 ( .A(n30525), .B(n30524), .Z(n30526) );
  AND U48265 ( .A(n52447), .B(n30526), .Z(n30529) );
  NANDN U48266 ( .A(x[556]), .B(y[556]), .Z(n30528) );
  NAND U48267 ( .A(n30528), .B(n30527), .Z(n52448) );
  OR U48268 ( .A(n30529), .B(n52448), .Z(n30530) );
  NAND U48269 ( .A(n52449), .B(n30530), .Z(n30531) );
  NANDN U48270 ( .A(n30532), .B(n30531), .Z(n30533) );
  OR U48271 ( .A(n30533), .B(n52450), .Z(n30534) );
  AND U48272 ( .A(n30535), .B(n30534), .Z(n30536) );
  NOR U48273 ( .A(n52454), .B(n30536), .Z(n30537) );
  NANDN U48274 ( .A(n30538), .B(n30537), .Z(n30539) );
  AND U48275 ( .A(n52455), .B(n30539), .Z(n30542) );
  NAND U48276 ( .A(n30541), .B(n30540), .Z(n52437) );
  OR U48277 ( .A(n30542), .B(n52437), .Z(n30543) );
  NAND U48278 ( .A(n52456), .B(n30543), .Z(n30544) );
  NANDN U48279 ( .A(n30545), .B(n30544), .Z(n30546) );
  OR U48280 ( .A(n30546), .B(n52457), .Z(n30547) );
  AND U48281 ( .A(n30548), .B(n30547), .Z(n30549) );
  NOR U48282 ( .A(n52462), .B(n30549), .Z(n30550) );
  NANDN U48283 ( .A(n30551), .B(n30550), .Z(n30552) );
  AND U48284 ( .A(n52463), .B(n30552), .Z(n30555) );
  NAND U48285 ( .A(n30554), .B(n30553), .Z(n52436) );
  OR U48286 ( .A(n30555), .B(n52436), .Z(n30556) );
  NAND U48287 ( .A(n52464), .B(n30556), .Z(n30557) );
  NANDN U48288 ( .A(n30558), .B(n30557), .Z(n30559) );
  OR U48289 ( .A(n30559), .B(n52465), .Z(n30560) );
  NAND U48290 ( .A(n52466), .B(n30560), .Z(n30561) );
  NANDN U48291 ( .A(n52434), .B(n30561), .Z(n30562) );
  NAND U48292 ( .A(n52467), .B(n30562), .Z(n30563) );
  NANDN U48293 ( .A(n52433), .B(n30563), .Z(n30564) );
  AND U48294 ( .A(n52468), .B(n30564), .Z(n30565) );
  NOR U48295 ( .A(n30565), .B(n52469), .Z(n30566) );
  NANDN U48296 ( .A(n30567), .B(n30566), .Z(n30568) );
  AND U48297 ( .A(n30569), .B(n30568), .Z(n30570) );
  NAND U48298 ( .A(n30570), .B(n52470), .Z(n30572) );
  ANDN U48299 ( .B(y[578]), .A(x[578]), .Z(n30571) );
  ANDN U48300 ( .B(n30572), .A(n30571), .Z(n30573) );
  NANDN U48301 ( .A(n52473), .B(n30573), .Z(n30574) );
  NAND U48302 ( .A(n52475), .B(n30574), .Z(n30575) );
  NANDN U48303 ( .A(n52432), .B(n30575), .Z(n30576) );
  AND U48304 ( .A(n52476), .B(n30576), .Z(n30577) );
  NOR U48305 ( .A(n52477), .B(n30577), .Z(n30578) );
  NANDN U48306 ( .A(n30579), .B(n30578), .Z(n30580) );
  AND U48307 ( .A(n30581), .B(n30580), .Z(n30582) );
  ANDN U48308 ( .B(n30583), .A(n30582), .Z(n30584) );
  NAND U48309 ( .A(n52481), .B(n30584), .Z(n30585) );
  NANDN U48310 ( .A(n52482), .B(n30585), .Z(n30586) );
  NAND U48311 ( .A(n52483), .B(n30586), .Z(n30587) );
  NANDN U48312 ( .A(n52484), .B(n30587), .Z(n30588) );
  AND U48313 ( .A(n30589), .B(n30588), .Z(n30590) );
  NAND U48314 ( .A(n30590), .B(n52485), .Z(n30591) );
  AND U48315 ( .A(n30592), .B(n30591), .Z(n30593) );
  NOR U48316 ( .A(n52489), .B(n30593), .Z(n30594) );
  NANDN U48317 ( .A(n30595), .B(n30594), .Z(n30596) );
  AND U48318 ( .A(n52490), .B(n30596), .Z(n30599) );
  NAND U48319 ( .A(n30598), .B(n30597), .Z(n52431) );
  OR U48320 ( .A(n30599), .B(n52431), .Z(n30600) );
  NAND U48321 ( .A(n52492), .B(n30600), .Z(n30601) );
  NANDN U48322 ( .A(n30602), .B(n30601), .Z(n30603) );
  OR U48323 ( .A(n30603), .B(n52493), .Z(n30604) );
  NAND U48324 ( .A(n30605), .B(n30604), .Z(n30606) );
  NANDN U48325 ( .A(n30607), .B(n30606), .Z(n30608) );
  OR U48326 ( .A(n30608), .B(n52497), .Z(n30609) );
  NAND U48327 ( .A(n52498), .B(n30609), .Z(n30610) );
  NANDN U48328 ( .A(n52499), .B(n30610), .Z(n30611) );
  NAND U48329 ( .A(n52500), .B(n30611), .Z(n30612) );
  ANDN U48330 ( .B(n30612), .A(n52501), .Z(n30613) );
  NANDN U48331 ( .A(n30614), .B(n30613), .Z(n30616) );
  AND U48332 ( .A(n52502), .B(n52504), .Z(n30615) );
  NAND U48333 ( .A(n30616), .B(n30615), .Z(n30617) );
  NANDN U48334 ( .A(n30618), .B(n30617), .Z(n30619) );
  OR U48335 ( .A(n30619), .B(n52505), .Z(n30620) );
  NAND U48336 ( .A(n52506), .B(n30620), .Z(n30621) );
  NANDN U48337 ( .A(n52430), .B(n30621), .Z(n30622) );
  NAND U48338 ( .A(n52507), .B(n30622), .Z(n30623) );
  ANDN U48339 ( .B(n30623), .A(n52508), .Z(n30624) );
  NANDN U48340 ( .A(n30625), .B(n30624), .Z(n30628) );
  AND U48341 ( .A(n30626), .B(n52510), .Z(n30627) );
  NAND U48342 ( .A(n30628), .B(n30627), .Z(n30629) );
  NANDN U48343 ( .A(n52513), .B(n30629), .Z(n30631) );
  ANDN U48344 ( .B(y[608]), .A(x[608]), .Z(n30630) );
  OR U48345 ( .A(n30631), .B(n30630), .Z(n30632) );
  NAND U48346 ( .A(n52514), .B(n30632), .Z(n30633) );
  NANDN U48347 ( .A(n52429), .B(n30633), .Z(n30634) );
  NAND U48348 ( .A(n52515), .B(n30634), .Z(n30635) );
  ANDN U48349 ( .B(n30635), .A(n52516), .Z(n30636) );
  NANDN U48350 ( .A(n30637), .B(n30636), .Z(n30638) );
  AND U48351 ( .A(n30638), .B(n52519), .Z(n30639) );
  NAND U48352 ( .A(n52517), .B(n30639), .Z(n30640) );
  AND U48353 ( .A(n30641), .B(n30640), .Z(n30642) );
  NANDN U48354 ( .A(n52520), .B(n30642), .Z(n30643) );
  NAND U48355 ( .A(n52521), .B(n30643), .Z(n30644) );
  NANDN U48356 ( .A(n52522), .B(n30644), .Z(n30645) );
  NAND U48357 ( .A(n52523), .B(n30645), .Z(n30646) );
  ANDN U48358 ( .B(n30646), .A(n52524), .Z(n30647) );
  NANDN U48359 ( .A(n30648), .B(n30647), .Z(n30649) );
  AND U48360 ( .A(n30649), .B(n52525), .Z(n30650) );
  NAND U48361 ( .A(n30651), .B(n30650), .Z(n30652) );
  AND U48362 ( .A(n30653), .B(n30652), .Z(n30654) );
  NANDN U48363 ( .A(n30655), .B(n30654), .Z(n30656) );
  AND U48364 ( .A(n30657), .B(n30656), .Z(n30659) );
  ANDN U48365 ( .B(y[622]), .A(x[622]), .Z(n30658) );
  NOR U48366 ( .A(n30659), .B(n30658), .Z(n30660) );
  NANDN U48367 ( .A(n30661), .B(n30660), .Z(n30662) );
  AND U48368 ( .A(n30663), .B(n30662), .Z(n30665) );
  NAND U48369 ( .A(n30665), .B(n30664), .Z(n30667) );
  ANDN U48370 ( .B(n30667), .A(n30666), .Z(n30668) );
  NANDN U48371 ( .A(n30669), .B(n30668), .Z(n30673) );
  AND U48372 ( .A(n30671), .B(n30670), .Z(n30672) );
  NAND U48373 ( .A(n30673), .B(n30672), .Z(n30674) );
  NANDN U48374 ( .A(n30675), .B(n30674), .Z(n30677) );
  OR U48375 ( .A(n30677), .B(n30676), .Z(n30678) );
  AND U48376 ( .A(n30679), .B(n30678), .Z(n30681) );
  ANDN U48377 ( .B(y[628]), .A(x[628]), .Z(n30680) );
  NOR U48378 ( .A(n30681), .B(n30680), .Z(n30682) );
  NANDN U48379 ( .A(n30683), .B(n30682), .Z(n30684) );
  AND U48380 ( .A(n30685), .B(n30684), .Z(n30687) );
  NAND U48381 ( .A(n30687), .B(n30686), .Z(n30689) );
  ANDN U48382 ( .B(n30689), .A(n30688), .Z(n30690) );
  NANDN U48383 ( .A(n30691), .B(n30690), .Z(n30695) );
  AND U48384 ( .A(n30693), .B(n30692), .Z(n30694) );
  NAND U48385 ( .A(n30695), .B(n30694), .Z(n30696) );
  NANDN U48386 ( .A(n30697), .B(n30696), .Z(n30699) );
  OR U48387 ( .A(n30699), .B(n30698), .Z(n30700) );
  AND U48388 ( .A(n30701), .B(n30700), .Z(n30703) );
  NOR U48389 ( .A(n30703), .B(n30702), .Z(n30704) );
  NANDN U48390 ( .A(n30705), .B(n30704), .Z(n30706) );
  AND U48391 ( .A(n30707), .B(n30706), .Z(n30709) );
  NAND U48392 ( .A(n30709), .B(n30708), .Z(n30711) );
  ANDN U48393 ( .B(n30711), .A(n30710), .Z(n30712) );
  NANDN U48394 ( .A(n30713), .B(n30712), .Z(n30717) );
  AND U48395 ( .A(n30715), .B(n30714), .Z(n30716) );
  NAND U48396 ( .A(n30717), .B(n30716), .Z(n30718) );
  NANDN U48397 ( .A(n30719), .B(n30718), .Z(n30721) );
  OR U48398 ( .A(n30721), .B(n30720), .Z(n30722) );
  AND U48399 ( .A(n30723), .B(n30722), .Z(n30725) );
  NOR U48400 ( .A(n30725), .B(n30724), .Z(n30726) );
  NANDN U48401 ( .A(n30727), .B(n30726), .Z(n30728) );
  AND U48402 ( .A(n30729), .B(n30728), .Z(n30731) );
  NAND U48403 ( .A(n30731), .B(n30730), .Z(n30733) );
  ANDN U48404 ( .B(y[642]), .A(x[642]), .Z(n30732) );
  ANDN U48405 ( .B(n30733), .A(n30732), .Z(n30734) );
  NANDN U48406 ( .A(n52571), .B(n30734), .Z(n30737) );
  AND U48407 ( .A(n30735), .B(n52572), .Z(n30736) );
  NAND U48408 ( .A(n30737), .B(n30736), .Z(n30738) );
  NANDN U48409 ( .A(n52428), .B(n30738), .Z(n30741) );
  AND U48410 ( .A(n30739), .B(n52427), .Z(n30740) );
  NAND U48411 ( .A(n30741), .B(n30740), .Z(n30742) );
  NANDN U48412 ( .A(n30743), .B(n30742), .Z(n30744) );
  OR U48413 ( .A(n30744), .B(n52573), .Z(n30745) );
  AND U48414 ( .A(n30746), .B(n30745), .Z(n30748) );
  NOR U48415 ( .A(n30748), .B(n30747), .Z(n30749) );
  NANDN U48416 ( .A(n30750), .B(n30749), .Z(n30751) );
  AND U48417 ( .A(n30752), .B(n30751), .Z(n30754) );
  NAND U48418 ( .A(n30754), .B(n30753), .Z(n30756) );
  ANDN U48419 ( .B(n30756), .A(n30755), .Z(n30757) );
  NANDN U48420 ( .A(n30758), .B(n30757), .Z(n30762) );
  AND U48421 ( .A(n30760), .B(n30759), .Z(n30761) );
  NAND U48422 ( .A(n30762), .B(n30761), .Z(n30763) );
  NANDN U48423 ( .A(n30764), .B(n30763), .Z(n30765) );
  OR U48424 ( .A(n30766), .B(n30765), .Z(n30767) );
  AND U48425 ( .A(n30768), .B(n30767), .Z(n30770) );
  NAND U48426 ( .A(n30770), .B(n30769), .Z(n30772) );
  ANDN U48427 ( .B(n30772), .A(n30771), .Z(n30773) );
  NANDN U48428 ( .A(n30774), .B(n30773), .Z(n30778) );
  AND U48429 ( .A(n30776), .B(n30775), .Z(n30777) );
  NAND U48430 ( .A(n30778), .B(n30777), .Z(n30779) );
  NANDN U48431 ( .A(n30780), .B(n30779), .Z(n30783) );
  NANDN U48432 ( .A(x[657]), .B(n30783), .Z(n30782) );
  ANDN U48433 ( .B(n30782), .A(n30781), .Z(n30786) );
  XNOR U48434 ( .A(n30783), .B(x[657]), .Z(n30784) );
  NAND U48435 ( .A(n30784), .B(y[657]), .Z(n30785) );
  NAND U48436 ( .A(n30786), .B(n30785), .Z(n30787) );
  NAND U48437 ( .A(n52587), .B(n30787), .Z(n30788) );
  NANDN U48438 ( .A(n52588), .B(n30788), .Z(n30789) );
  AND U48439 ( .A(n52589), .B(n30789), .Z(n30790) );
  OR U48440 ( .A(n52590), .B(n30790), .Z(n30791) );
  NAND U48441 ( .A(n52426), .B(n30791), .Z(n30792) );
  NANDN U48442 ( .A(n52425), .B(n30792), .Z(n30793) );
  NAND U48443 ( .A(n52424), .B(n30793), .Z(n30794) );
  NAND U48444 ( .A(n52591), .B(n30794), .Z(n30795) );
  AND U48445 ( .A(n30796), .B(n30795), .Z(n30797) );
  NAND U48446 ( .A(n52592), .B(n30797), .Z(n30799) );
  ANDN U48447 ( .B(n30799), .A(n30798), .Z(n30800) );
  NANDN U48448 ( .A(n52423), .B(n30800), .Z(n30804) );
  AND U48449 ( .A(n30802), .B(n30801), .Z(n30803) );
  NAND U48450 ( .A(n30804), .B(n30803), .Z(n30805) );
  NANDN U48451 ( .A(n30806), .B(n30805), .Z(n30808) );
  OR U48452 ( .A(n30808), .B(n30807), .Z(n30809) );
  AND U48453 ( .A(n30810), .B(n30809), .Z(n30812) );
  NOR U48454 ( .A(n30812), .B(n30811), .Z(n30813) );
  NANDN U48455 ( .A(n30814), .B(n30813), .Z(n30815) );
  AND U48456 ( .A(n30816), .B(n30815), .Z(n30818) );
  NAND U48457 ( .A(n30818), .B(n30817), .Z(n30820) );
  ANDN U48458 ( .B(n30820), .A(n30819), .Z(n30821) );
  NANDN U48459 ( .A(n30822), .B(n30821), .Z(n30825) );
  AND U48460 ( .A(n30823), .B(n52417), .Z(n30824) );
  NAND U48461 ( .A(n30825), .B(n30824), .Z(n30826) );
  NAND U48462 ( .A(n52597), .B(n30826), .Z(n30829) );
  AND U48463 ( .A(n30827), .B(n52598), .Z(n30828) );
  NAND U48464 ( .A(n30829), .B(n30828), .Z(n30830) );
  NANDN U48465 ( .A(n30831), .B(n30830), .Z(n30832) );
  OR U48466 ( .A(n30832), .B(n52416), .Z(n30833) );
  AND U48467 ( .A(n30834), .B(n30833), .Z(n30836) );
  NAND U48468 ( .A(n30836), .B(n30835), .Z(n30838) );
  ANDN U48469 ( .B(n30838), .A(n30837), .Z(n30839) );
  NANDN U48470 ( .A(n30840), .B(n30839), .Z(n30844) );
  AND U48471 ( .A(n30842), .B(n30841), .Z(n30843) );
  NAND U48472 ( .A(n30844), .B(n30843), .Z(n30845) );
  NANDN U48473 ( .A(n30846), .B(n30845), .Z(n30848) );
  OR U48474 ( .A(n30848), .B(n30847), .Z(n30849) );
  NAND U48475 ( .A(n30850), .B(n30849), .Z(n30854) );
  IV U48476 ( .A(n30851), .Z(n52603) );
  AND U48477 ( .A(n30852), .B(n52603), .Z(n30853) );
  NAND U48478 ( .A(n30854), .B(n30853), .Z(n30855) );
  NANDN U48479 ( .A(n30856), .B(n30855), .Z(n30857) );
  NANDN U48480 ( .A(n30857), .B(n52604), .Z(n30858) );
  AND U48481 ( .A(n52605), .B(n30858), .Z(n30860) );
  NAND U48482 ( .A(n52606), .B(n52607), .Z(n30859) );
  OR U48483 ( .A(n30860), .B(n30859), .Z(n30861) );
  AND U48484 ( .A(n30862), .B(n30861), .Z(n30864) );
  NANDN U48485 ( .A(x[686]), .B(y[686]), .Z(n30863) );
  NAND U48486 ( .A(n30864), .B(n30863), .Z(n30866) );
  ANDN U48487 ( .B(n30866), .A(n30865), .Z(n30867) );
  NANDN U48488 ( .A(n30868), .B(n30867), .Z(n30872) );
  AND U48489 ( .A(n30870), .B(n30869), .Z(n30871) );
  NAND U48490 ( .A(n30872), .B(n30871), .Z(n30873) );
  NANDN U48491 ( .A(n30874), .B(n30873), .Z(n30876) );
  OR U48492 ( .A(n30876), .B(n30875), .Z(n30877) );
  AND U48493 ( .A(n30878), .B(n30877), .Z(n30882) );
  NAND U48494 ( .A(n30880), .B(n30879), .Z(n30881) );
  OR U48495 ( .A(n30882), .B(n30881), .Z(n30883) );
  AND U48496 ( .A(n30884), .B(n30883), .Z(n30886) );
  NAND U48497 ( .A(n30886), .B(n30885), .Z(n30888) );
  ANDN U48498 ( .B(n30888), .A(n30887), .Z(n30889) );
  NANDN U48499 ( .A(n30890), .B(n30889), .Z(n30894) );
  AND U48500 ( .A(n30892), .B(n30891), .Z(n30893) );
  NAND U48501 ( .A(n30894), .B(n30893), .Z(n30895) );
  NANDN U48502 ( .A(n30896), .B(n30895), .Z(n30898) );
  NANDN U48503 ( .A(n30898), .B(n30897), .Z(n30899) );
  NAND U48504 ( .A(n30900), .B(n30899), .Z(n30904) );
  AND U48505 ( .A(n30902), .B(n30901), .Z(n30903) );
  NAND U48506 ( .A(n30904), .B(n30903), .Z(n30905) );
  NANDN U48507 ( .A(n30906), .B(n30905), .Z(n30907) );
  OR U48508 ( .A(n30908), .B(n30907), .Z(n30909) );
  AND U48509 ( .A(n30910), .B(n30909), .Z(n30911) );
  NANDN U48510 ( .A(n30912), .B(n30911), .Z(n30913) );
  AND U48511 ( .A(n30914), .B(n30913), .Z(n30916) );
  NAND U48512 ( .A(n30916), .B(n30915), .Z(n30918) );
  ANDN U48513 ( .B(n30918), .A(n30917), .Z(n30919) );
  NANDN U48514 ( .A(n30920), .B(n30919), .Z(n30924) );
  AND U48515 ( .A(n30922), .B(n30921), .Z(n30923) );
  NAND U48516 ( .A(n30924), .B(n30923), .Z(n30925) );
  NANDN U48517 ( .A(n30926), .B(n30925), .Z(n30927) );
  OR U48518 ( .A(n30928), .B(n30927), .Z(n30929) );
  AND U48519 ( .A(n30930), .B(n30929), .Z(n30931) );
  NAND U48520 ( .A(n30932), .B(n30931), .Z(n30933) );
  NAND U48521 ( .A(n30934), .B(n30933), .Z(n30935) );
  AND U48522 ( .A(n30936), .B(n30935), .Z(n30937) );
  OR U48523 ( .A(n52647), .B(n30937), .Z(n30938) );
  AND U48524 ( .A(n52649), .B(n30938), .Z(n30939) );
  OR U48525 ( .A(n30939), .B(n52651), .Z(n30940) );
  AND U48526 ( .A(n52652), .B(n30940), .Z(n30941) );
  OR U48527 ( .A(n52653), .B(n30941), .Z(n30942) );
  NAND U48528 ( .A(n30943), .B(n30942), .Z(n30944) );
  NANDN U48529 ( .A(n30945), .B(n30944), .Z(n30948) );
  AND U48530 ( .A(n30946), .B(n52656), .Z(n30947) );
  NAND U48531 ( .A(n30948), .B(n30947), .Z(n30949) );
  NANDN U48532 ( .A(n52657), .B(n30949), .Z(n30951) );
  OR U48533 ( .A(n30951), .B(n30950), .Z(n30952) );
  NAND U48534 ( .A(n52658), .B(n30952), .Z(n30953) );
  NANDN U48535 ( .A(n30954), .B(n30953), .Z(n30955) );
  NANDN U48536 ( .A(n30955), .B(n52659), .Z(n30956) );
  AND U48537 ( .A(n30957), .B(n30956), .Z(n30958) );
  NAND U48538 ( .A(n30958), .B(n52660), .Z(n30960) );
  ANDN U48539 ( .B(n30960), .A(n30959), .Z(n30961) );
  NANDN U48540 ( .A(n30962), .B(n30961), .Z(n30966) );
  AND U48541 ( .A(n30964), .B(n30963), .Z(n30965) );
  NAND U48542 ( .A(n30966), .B(n30965), .Z(n30967) );
  NANDN U48543 ( .A(n30968), .B(n30967), .Z(n30970) );
  OR U48544 ( .A(n30970), .B(n30969), .Z(n30971) );
  NAND U48545 ( .A(n30972), .B(n30971), .Z(n30976) );
  AND U48546 ( .A(n30974), .B(n30973), .Z(n30975) );
  NAND U48547 ( .A(n30976), .B(n30975), .Z(n30977) );
  NANDN U48548 ( .A(n30978), .B(n30977), .Z(n30979) );
  OR U48549 ( .A(n30979), .B(n52668), .Z(n30980) );
  NAND U48550 ( .A(n30981), .B(n30980), .Z(n30982) );
  NANDN U48551 ( .A(n52411), .B(n30982), .Z(n30984) );
  AND U48552 ( .A(n52671), .B(n52410), .Z(n30983) );
  NAND U48553 ( .A(n30984), .B(n30983), .Z(n30985) );
  NANDN U48554 ( .A(n30986), .B(n30985), .Z(n30988) );
  ANDN U48555 ( .B(y[726]), .A(x[726]), .Z(n30987) );
  OR U48556 ( .A(n30988), .B(n30987), .Z(n30989) );
  NAND U48557 ( .A(n30990), .B(n30989), .Z(n30991) );
  NANDN U48558 ( .A(n30992), .B(n30991), .Z(n30994) );
  ANDN U48559 ( .B(y[728]), .A(x[728]), .Z(n30993) );
  OR U48560 ( .A(n30994), .B(n30993), .Z(n30995) );
  NAND U48561 ( .A(n30996), .B(n30995), .Z(n31000) );
  AND U48562 ( .A(n30998), .B(n30997), .Z(n30999) );
  NAND U48563 ( .A(n31000), .B(n30999), .Z(n31001) );
  NANDN U48564 ( .A(n31002), .B(n31001), .Z(n31003) );
  OR U48565 ( .A(n31004), .B(n31003), .Z(n31005) );
  AND U48566 ( .A(n31006), .B(n31005), .Z(n31007) );
  NAND U48567 ( .A(n31007), .B(n52679), .Z(n31009) );
  IV U48568 ( .A(n31008), .Z(n52680) );
  ANDN U48569 ( .B(n31009), .A(n52680), .Z(n31010) );
  NANDN U48570 ( .A(n31011), .B(n31010), .Z(n31014) );
  AND U48571 ( .A(n52681), .B(n31012), .Z(n31013) );
  NAND U48572 ( .A(n31014), .B(n31013), .Z(n31015) );
  NANDN U48573 ( .A(n31016), .B(n31015), .Z(n31017) );
  NANDN U48574 ( .A(n31017), .B(n52682), .Z(n31018) );
  AND U48575 ( .A(n31019), .B(n31018), .Z(n31020) );
  NANDN U48576 ( .A(n31021), .B(n31020), .Z(n31022) );
  AND U48577 ( .A(n31023), .B(n31022), .Z(n31025) );
  NAND U48578 ( .A(n31025), .B(n31024), .Z(n31027) );
  ANDN U48579 ( .B(n31027), .A(n31026), .Z(n31028) );
  NANDN U48580 ( .A(n31029), .B(n31028), .Z(n31033) );
  AND U48581 ( .A(n31031), .B(n31030), .Z(n31032) );
  NAND U48582 ( .A(n31033), .B(n31032), .Z(n31034) );
  NANDN U48583 ( .A(n31035), .B(n31034), .Z(n31037) );
  OR U48584 ( .A(n31037), .B(n31036), .Z(n31038) );
  NAND U48585 ( .A(n31039), .B(n31038), .Z(n31042) );
  AND U48586 ( .A(n31040), .B(n52696), .Z(n31041) );
  NAND U48587 ( .A(n31042), .B(n31041), .Z(n31043) );
  NAND U48588 ( .A(n52697), .B(n31043), .Z(n31044) );
  OR U48589 ( .A(n31045), .B(n31044), .Z(n31046) );
  AND U48590 ( .A(n52700), .B(n31046), .Z(n31048) );
  NAND U48591 ( .A(n31048), .B(n31047), .Z(n31050) );
  ANDN U48592 ( .B(n31050), .A(n31049), .Z(n31051) );
  NANDN U48593 ( .A(n52702), .B(n31051), .Z(n31055) );
  AND U48594 ( .A(n31053), .B(n31052), .Z(n31054) );
  NAND U48595 ( .A(n31055), .B(n31054), .Z(n31056) );
  NANDN U48596 ( .A(n31057), .B(n31056), .Z(n31059) );
  OR U48597 ( .A(n31059), .B(n31058), .Z(n31060) );
  NAND U48598 ( .A(n31061), .B(n31060), .Z(n31065) );
  AND U48599 ( .A(n31063), .B(n31062), .Z(n31064) );
  NAND U48600 ( .A(n31065), .B(n31064), .Z(n31066) );
  NANDN U48601 ( .A(n31067), .B(n31066), .Z(n31069) );
  OR U48602 ( .A(n31069), .B(n31068), .Z(n31070) );
  NAND U48603 ( .A(n31071), .B(n31070), .Z(n31072) );
  NANDN U48604 ( .A(n31073), .B(n31072), .Z(n31077) );
  AND U48605 ( .A(n31075), .B(n31074), .Z(n31076) );
  NAND U48606 ( .A(n31077), .B(n31076), .Z(n31078) );
  NANDN U48607 ( .A(n31079), .B(n31078), .Z(n31081) );
  OR U48608 ( .A(n31081), .B(n31080), .Z(n31082) );
  NAND U48609 ( .A(n31083), .B(n31082), .Z(n31084) );
  NANDN U48610 ( .A(n31085), .B(n31084), .Z(n31089) );
  AND U48611 ( .A(n31087), .B(n31086), .Z(n31088) );
  NAND U48612 ( .A(n31089), .B(n31088), .Z(n31090) );
  NANDN U48613 ( .A(n31091), .B(n31090), .Z(n31093) );
  OR U48614 ( .A(n31093), .B(n31092), .Z(n31094) );
  NAND U48615 ( .A(n31095), .B(n31094), .Z(n31096) );
  NANDN U48616 ( .A(n31097), .B(n31096), .Z(n31101) );
  AND U48617 ( .A(n31099), .B(n31098), .Z(n31100) );
  NAND U48618 ( .A(n31101), .B(n31100), .Z(n31102) );
  NANDN U48619 ( .A(n31103), .B(n31102), .Z(n31104) );
  OR U48620 ( .A(n31104), .B(n52734), .Z(n31105) );
  NAND U48621 ( .A(n31106), .B(n31105), .Z(n31107) );
  NANDN U48622 ( .A(n52736), .B(n31107), .Z(n31110) );
  AND U48623 ( .A(n31108), .B(n52737), .Z(n31109) );
  NAND U48624 ( .A(n31110), .B(n31109), .Z(n31111) );
  NANDN U48625 ( .A(n31112), .B(n31111), .Z(n31114) );
  IV U48626 ( .A(n31113), .Z(n52738) );
  OR U48627 ( .A(n31114), .B(n52738), .Z(n31115) );
  AND U48628 ( .A(n31116), .B(n31115), .Z(n31118) );
  NAND U48629 ( .A(n31118), .B(n31117), .Z(n31120) );
  ANDN U48630 ( .B(n31120), .A(n31119), .Z(n31121) );
  NANDN U48631 ( .A(n31122), .B(n31121), .Z(n31126) );
  AND U48632 ( .A(n31124), .B(n31123), .Z(n31125) );
  NAND U48633 ( .A(n31126), .B(n31125), .Z(n31127) );
  NANDN U48634 ( .A(n31128), .B(n31127), .Z(n31130) );
  OR U48635 ( .A(n31130), .B(n31129), .Z(n31131) );
  NAND U48636 ( .A(n31132), .B(n31131), .Z(n31135) );
  AND U48637 ( .A(n31133), .B(n52406), .Z(n31134) );
  NAND U48638 ( .A(n31135), .B(n31134), .Z(n31136) );
  NANDN U48639 ( .A(n52745), .B(n31136), .Z(n31137) );
  OR U48640 ( .A(n31138), .B(n31137), .Z(n31139) );
  AND U48641 ( .A(n31139), .B(n52405), .Z(n31140) );
  NAND U48642 ( .A(n31141), .B(n31140), .Z(n31142) );
  AND U48643 ( .A(n31143), .B(n31142), .Z(n31144) );
  NAND U48644 ( .A(n31144), .B(n52746), .Z(n31148) );
  NANDN U48645 ( .A(x[776]), .B(y[776]), .Z(n31145) );
  AND U48646 ( .A(n31146), .B(n31145), .Z(n31147) );
  NAND U48647 ( .A(n31148), .B(n31147), .Z(n31149) );
  NANDN U48648 ( .A(n31150), .B(n31149), .Z(n31152) );
  OR U48649 ( .A(n31152), .B(n31151), .Z(n31153) );
  NAND U48650 ( .A(n31154), .B(n31153), .Z(n31155) );
  NANDN U48651 ( .A(n31156), .B(n31155), .Z(n31159) );
  NANDN U48652 ( .A(y[780]), .B(n31159), .Z(n31158) );
  ANDN U48653 ( .B(n31158), .A(n31157), .Z(n31162) );
  XNOR U48654 ( .A(n31159), .B(y[780]), .Z(n31160) );
  NAND U48655 ( .A(n31160), .B(x[780]), .Z(n31161) );
  NAND U48656 ( .A(n31162), .B(n31161), .Z(n31163) );
  NAND U48657 ( .A(n52749), .B(n31163), .Z(n31164) );
  NANDN U48658 ( .A(n52750), .B(n31164), .Z(n31165) );
  AND U48659 ( .A(n52752), .B(n31165), .Z(n31167) );
  IV U48660 ( .A(n31166), .Z(n52753) );
  OR U48661 ( .A(n31167), .B(n52753), .Z(n31168) );
  AND U48662 ( .A(n52754), .B(n31168), .Z(n31170) );
  NAND U48663 ( .A(n52400), .B(n52755), .Z(n31169) );
  OR U48664 ( .A(n31170), .B(n31169), .Z(n31171) );
  AND U48665 ( .A(n31172), .B(n31171), .Z(n31174) );
  NANDN U48666 ( .A(x[786]), .B(y[786]), .Z(n31173) );
  NAND U48667 ( .A(n31174), .B(n31173), .Z(n31176) );
  ANDN U48668 ( .B(n31176), .A(n31175), .Z(n31177) );
  NANDN U48669 ( .A(n31178), .B(n31177), .Z(n31182) );
  AND U48670 ( .A(n31180), .B(n31179), .Z(n31181) );
  NAND U48671 ( .A(n31182), .B(n31181), .Z(n31183) );
  NANDN U48672 ( .A(n31184), .B(n31183), .Z(n31186) );
  OR U48673 ( .A(n31186), .B(n31185), .Z(n31187) );
  NAND U48674 ( .A(n31188), .B(n31187), .Z(n31192) );
  AND U48675 ( .A(n31190), .B(n31189), .Z(n31191) );
  NAND U48676 ( .A(n31192), .B(n31191), .Z(n31193) );
  NANDN U48677 ( .A(n52763), .B(n31193), .Z(n31195) );
  OR U48678 ( .A(n31195), .B(n31194), .Z(n31196) );
  NAND U48679 ( .A(n31197), .B(n31196), .Z(n31198) );
  NANDN U48680 ( .A(n52399), .B(n31198), .Z(n31201) );
  AND U48681 ( .A(n31199), .B(n52398), .Z(n31200) );
  NAND U48682 ( .A(n31201), .B(n31200), .Z(n31202) );
  NANDN U48683 ( .A(n52766), .B(n31202), .Z(n31203) );
  OR U48684 ( .A(n31204), .B(n31203), .Z(n31205) );
  AND U48685 ( .A(n31206), .B(n31205), .Z(n31207) );
  NANDN U48686 ( .A(n31208), .B(n31207), .Z(n31209) );
  AND U48687 ( .A(n31210), .B(n31209), .Z(n31211) );
  ANDN U48688 ( .B(n31212), .A(n31211), .Z(n31213) );
  NAND U48689 ( .A(n31214), .B(n31213), .Z(n31215) );
  NANDN U48690 ( .A(n31216), .B(n31215), .Z(n31217) );
  OR U48691 ( .A(n31218), .B(n31217), .Z(n31219) );
  AND U48692 ( .A(n31220), .B(n31219), .Z(n31221) );
  NANDN U48693 ( .A(n31222), .B(n31221), .Z(n31223) );
  AND U48694 ( .A(n31224), .B(n31223), .Z(n31226) );
  NOR U48695 ( .A(n31226), .B(n31225), .Z(n31227) );
  NANDN U48696 ( .A(n31228), .B(n31227), .Z(n31229) );
  AND U48697 ( .A(n31230), .B(n31229), .Z(n31232) );
  AND U48698 ( .A(n31232), .B(n31231), .Z(n31236) );
  AND U48699 ( .A(n31234), .B(n31233), .Z(n31235) );
  NANDN U48700 ( .A(n31236), .B(n31235), .Z(n31237) );
  NAND U48701 ( .A(n31238), .B(n31237), .Z(n31242) );
  AND U48702 ( .A(n31240), .B(n31239), .Z(n31241) );
  NAND U48703 ( .A(n31242), .B(n31241), .Z(n31243) );
  NANDN U48704 ( .A(n31244), .B(n31243), .Z(n31246) );
  OR U48705 ( .A(n31246), .B(n31245), .Z(n31247) );
  NAND U48706 ( .A(n31248), .B(n31247), .Z(n31249) );
  NANDN U48707 ( .A(n31250), .B(n31249), .Z(n31254) );
  AND U48708 ( .A(n31252), .B(n31251), .Z(n31253) );
  NAND U48709 ( .A(n31254), .B(n31253), .Z(n31255) );
  NANDN U48710 ( .A(n31256), .B(n31255), .Z(n31257) );
  OR U48711 ( .A(n31257), .B(n52802), .Z(n31258) );
  NAND U48712 ( .A(n31259), .B(n31258), .Z(n31260) );
  NANDN U48713 ( .A(n52805), .B(n31260), .Z(n31262) );
  AND U48714 ( .A(n52811), .B(n52808), .Z(n31261) );
  NAND U48715 ( .A(n31262), .B(n31261), .Z(n31263) );
  NANDN U48716 ( .A(n31264), .B(n31263), .Z(n31266) );
  ANDN U48717 ( .B(y[816]), .A(x[816]), .Z(n31265) );
  OR U48718 ( .A(n31266), .B(n31265), .Z(n31267) );
  NAND U48719 ( .A(n31268), .B(n31267), .Z(n31272) );
  AND U48720 ( .A(n31270), .B(n31269), .Z(n31271) );
  NAND U48721 ( .A(n31272), .B(n31271), .Z(n31273) );
  NANDN U48722 ( .A(n31274), .B(n31273), .Z(n31276) );
  OR U48723 ( .A(n31276), .B(n31275), .Z(n31277) );
  NAND U48724 ( .A(n31278), .B(n31277), .Z(n31279) );
  NANDN U48725 ( .A(n31280), .B(n31279), .Z(n31284) );
  AND U48726 ( .A(n31282), .B(n31281), .Z(n31283) );
  NAND U48727 ( .A(n31284), .B(n31283), .Z(n31285) );
  NANDN U48728 ( .A(n31286), .B(n31285), .Z(n31287) );
  OR U48729 ( .A(n31288), .B(n31287), .Z(n31289) );
  AND U48730 ( .A(n31290), .B(n31289), .Z(n31292) );
  NAND U48731 ( .A(n31292), .B(n31291), .Z(n31293) );
  NANDN U48732 ( .A(n31294), .B(n31293), .Z(n31295) );
  AND U48733 ( .A(n31296), .B(n31295), .Z(n31297) );
  OR U48734 ( .A(n31298), .B(n31297), .Z(n31299) );
  NAND U48735 ( .A(n31300), .B(n31299), .Z(n31301) );
  NANDN U48736 ( .A(n31302), .B(n31301), .Z(n31304) );
  OR U48737 ( .A(n31304), .B(n31303), .Z(n31305) );
  NAND U48738 ( .A(n31306), .B(n31305), .Z(n31310) );
  AND U48739 ( .A(n31308), .B(n31307), .Z(n31309) );
  NAND U48740 ( .A(n31310), .B(n31309), .Z(n31311) );
  NANDN U48741 ( .A(n31312), .B(n31311), .Z(n31313) );
  OR U48742 ( .A(n31314), .B(n31313), .Z(n31315) );
  AND U48743 ( .A(n31316), .B(n31315), .Z(n31318) );
  NAND U48744 ( .A(n31318), .B(n31317), .Z(n31320) );
  ANDN U48745 ( .B(y[832]), .A(x[832]), .Z(n31319) );
  ANDN U48746 ( .B(n31320), .A(n31319), .Z(n31321) );
  NANDN U48747 ( .A(n52847), .B(n31321), .Z(n31324) );
  AND U48748 ( .A(n31322), .B(n52848), .Z(n31323) );
  NAND U48749 ( .A(n31324), .B(n31323), .Z(n31325) );
  NANDN U48750 ( .A(n52397), .B(n31325), .Z(n31328) );
  AND U48751 ( .A(n31326), .B(n52849), .Z(n31327) );
  NAND U48752 ( .A(n31328), .B(n31327), .Z(n31329) );
  NANDN U48753 ( .A(n52850), .B(n31329), .Z(n31331) );
  NAND U48754 ( .A(n31331), .B(n31330), .Z(n31332) );
  NANDN U48755 ( .A(n52852), .B(n31332), .Z(n31333) );
  AND U48756 ( .A(n31334), .B(n31333), .Z(n31335) );
  OR U48757 ( .A(n31336), .B(n31335), .Z(n31337) );
  NAND U48758 ( .A(n31338), .B(n31337), .Z(n31339) );
  NANDN U48759 ( .A(n31340), .B(n31339), .Z(n31344) );
  AND U48760 ( .A(n31342), .B(n31341), .Z(n31343) );
  NAND U48761 ( .A(n31344), .B(n31343), .Z(n31345) );
  NANDN U48762 ( .A(n31346), .B(n31345), .Z(n31347) );
  OR U48763 ( .A(n31347), .B(n52858), .Z(n31348) );
  NAND U48764 ( .A(n31349), .B(n31348), .Z(n31350) );
  NANDN U48765 ( .A(n52860), .B(n31350), .Z(n31351) );
  OR U48766 ( .A(n31352), .B(n31351), .Z(n31353) );
  AND U48767 ( .A(n31354), .B(n31353), .Z(n31355) );
  NANDN U48768 ( .A(n52861), .B(n31355), .Z(n31356) );
  AND U48769 ( .A(n31357), .B(n31356), .Z(n31359) );
  NOR U48770 ( .A(n31359), .B(n31358), .Z(n31360) );
  NANDN U48771 ( .A(n31361), .B(n31360), .Z(n31362) );
  AND U48772 ( .A(n31363), .B(n31362), .Z(n31364) );
  NANDN U48773 ( .A(n31365), .B(n31364), .Z(n31366) );
  NAND U48774 ( .A(n31367), .B(n31366), .Z(n31368) );
  NANDN U48775 ( .A(n31369), .B(n31368), .Z(n31373) );
  AND U48776 ( .A(n31371), .B(n31370), .Z(n31372) );
  NAND U48777 ( .A(n31373), .B(n31372), .Z(n31374) );
  NANDN U48778 ( .A(n31375), .B(n31374), .Z(n31376) );
  OR U48779 ( .A(n31377), .B(n31376), .Z(n31378) );
  AND U48780 ( .A(n31379), .B(n31378), .Z(n31381) );
  NAND U48781 ( .A(n31381), .B(n31380), .Z(n31383) );
  ANDN U48782 ( .B(n31383), .A(n31382), .Z(n31384) );
  NANDN U48783 ( .A(n31385), .B(n31384), .Z(n31389) );
  AND U48784 ( .A(n31387), .B(n31386), .Z(n31388) );
  NAND U48785 ( .A(n31389), .B(n31388), .Z(n31390) );
  NANDN U48786 ( .A(n31391), .B(n31390), .Z(n31393) );
  OR U48787 ( .A(n31393), .B(n31392), .Z(n31394) );
  AND U48788 ( .A(n31395), .B(n31394), .Z(n31399) );
  NAND U48789 ( .A(n31397), .B(n31396), .Z(n31398) );
  OR U48790 ( .A(n31399), .B(n31398), .Z(n31400) );
  AND U48791 ( .A(n31401), .B(n31400), .Z(n31403) );
  NAND U48792 ( .A(n31403), .B(n31402), .Z(n31405) );
  ANDN U48793 ( .B(n31405), .A(n31404), .Z(n31406) );
  NANDN U48794 ( .A(n31407), .B(n31406), .Z(n31411) );
  AND U48795 ( .A(n31409), .B(n31408), .Z(n31410) );
  NAND U48796 ( .A(n31411), .B(n31410), .Z(n31412) );
  NANDN U48797 ( .A(n31413), .B(n31412), .Z(n31414) );
  OR U48798 ( .A(n31414), .B(n52385), .Z(n31415) );
  AND U48799 ( .A(n31416), .B(n31415), .Z(n31417) );
  NAND U48800 ( .A(n52384), .B(n31417), .Z(n31418) );
  NAND U48801 ( .A(n52872), .B(n31418), .Z(n31419) );
  AND U48802 ( .A(n31420), .B(n31419), .Z(n31421) );
  NAND U48803 ( .A(n52873), .B(n31421), .Z(n31423) );
  ANDN U48804 ( .B(n31423), .A(n31422), .Z(n31424) );
  NANDN U48805 ( .A(n52383), .B(n31424), .Z(n31428) );
  AND U48806 ( .A(n31426), .B(n31425), .Z(n31427) );
  NAND U48807 ( .A(n31428), .B(n31427), .Z(n31429) );
  NANDN U48808 ( .A(n31430), .B(n31429), .Z(n31431) );
  OR U48809 ( .A(n31432), .B(n31431), .Z(n31433) );
  AND U48810 ( .A(n31434), .B(n31433), .Z(n31435) );
  NANDN U48811 ( .A(n31436), .B(n31435), .Z(n31437) );
  AND U48812 ( .A(n31438), .B(n31437), .Z(n31440) );
  NAND U48813 ( .A(n31440), .B(n31439), .Z(n31442) );
  ANDN U48814 ( .B(n31442), .A(n31441), .Z(n31443) );
  NANDN U48815 ( .A(n31444), .B(n31443), .Z(n31448) );
  IV U48816 ( .A(n31445), .Z(n52880) );
  AND U48817 ( .A(n31446), .B(n52880), .Z(n31447) );
  NAND U48818 ( .A(n31448), .B(n31447), .Z(n31449) );
  NANDN U48819 ( .A(n31450), .B(n31449), .Z(n31451) );
  NANDN U48820 ( .A(n31451), .B(n52881), .Z(n31452) );
  NAND U48821 ( .A(n52882), .B(n31452), .Z(n31453) );
  AND U48822 ( .A(n31454), .B(n31453), .Z(n31455) );
  NAND U48823 ( .A(n52883), .B(n31455), .Z(n31457) );
  ANDN U48824 ( .B(n31457), .A(n31456), .Z(n31458) );
  NANDN U48825 ( .A(n52884), .B(n31458), .Z(n31462) );
  AND U48826 ( .A(n31460), .B(n31459), .Z(n31461) );
  NAND U48827 ( .A(n31462), .B(n31461), .Z(n31463) );
  NANDN U48828 ( .A(n31464), .B(n31463), .Z(n31466) );
  OR U48829 ( .A(n31466), .B(n31465), .Z(n31467) );
  AND U48830 ( .A(n31468), .B(n31467), .Z(n31472) );
  NAND U48831 ( .A(n31470), .B(n31469), .Z(n31471) );
  OR U48832 ( .A(n31472), .B(n31471), .Z(n31473) );
  AND U48833 ( .A(n52888), .B(n31473), .Z(n31475) );
  NAND U48834 ( .A(n31475), .B(n31474), .Z(n31476) );
  NANDN U48835 ( .A(n31477), .B(n31476), .Z(n31478) );
  AND U48836 ( .A(n31478), .B(n52374), .Z(n31481) );
  NANDN U48837 ( .A(n31481), .B(n52889), .Z(n31482) );
  AND U48838 ( .A(n31483), .B(n31482), .Z(n31484) );
  NAND U48839 ( .A(n52890), .B(n31484), .Z(n31485) );
  AND U48840 ( .A(n52891), .B(n31485), .Z(n31491) );
  OR U48841 ( .A(n31487), .B(n31486), .Z(n31488) );
  AND U48842 ( .A(n31489), .B(n31488), .Z(n31490) );
  NANDN U48843 ( .A(n31491), .B(n31490), .Z(n31492) );
  NANDN U48844 ( .A(n52372), .B(n31492), .Z(n31493) );
  AND U48845 ( .A(n31493), .B(n52371), .Z(n31494) );
  OR U48846 ( .A(n31495), .B(n31494), .Z(n31496) );
  AND U48847 ( .A(n31497), .B(n31496), .Z(n31498) );
  ANDN U48848 ( .B(n31499), .A(n31498), .Z(n31500) );
  NAND U48849 ( .A(n31501), .B(n31500), .Z(n31502) );
  NANDN U48850 ( .A(n31503), .B(n31502), .Z(n31505) );
  OR U48851 ( .A(n31505), .B(n31504), .Z(n31506) );
  NAND U48852 ( .A(n31507), .B(n31506), .Z(n31508) );
  NANDN U48853 ( .A(n31509), .B(n31508), .Z(n31510) );
  AND U48854 ( .A(n31511), .B(n31510), .Z(n31512) );
  NAND U48855 ( .A(n31513), .B(n31512), .Z(n31514) );
  NANDN U48856 ( .A(n31515), .B(n31514), .Z(n31516) );
  OR U48857 ( .A(n31517), .B(n31516), .Z(n31518) );
  AND U48858 ( .A(n31519), .B(n31518), .Z(n31520) );
  NANDN U48859 ( .A(n31521), .B(n31520), .Z(n31522) );
  AND U48860 ( .A(n31523), .B(n31522), .Z(n31525) );
  NOR U48861 ( .A(n31525), .B(n31524), .Z(n31526) );
  NANDN U48862 ( .A(n31527), .B(n31526), .Z(n31528) );
  AND U48863 ( .A(n31529), .B(n31528), .Z(n31530) );
  NANDN U48864 ( .A(n31531), .B(n31530), .Z(n31532) );
  NAND U48865 ( .A(n31533), .B(n31532), .Z(n31534) );
  NANDN U48866 ( .A(n31535), .B(n31534), .Z(n31539) );
  AND U48867 ( .A(n31537), .B(n31536), .Z(n31538) );
  NAND U48868 ( .A(n31539), .B(n31538), .Z(n31540) );
  NANDN U48869 ( .A(n31541), .B(n31540), .Z(n31542) );
  OR U48870 ( .A(n31543), .B(n31542), .Z(n31544) );
  AND U48871 ( .A(n31545), .B(n31544), .Z(n31546) );
  NANDN U48872 ( .A(n31547), .B(n31546), .Z(n31548) );
  AND U48873 ( .A(n31549), .B(n31548), .Z(n31551) );
  NOR U48874 ( .A(n31551), .B(n31550), .Z(n31552) );
  NANDN U48875 ( .A(n31553), .B(n31552), .Z(n31554) );
  AND U48876 ( .A(n31555), .B(n31554), .Z(n31556) );
  NANDN U48877 ( .A(n31557), .B(n31556), .Z(n31558) );
  NAND U48878 ( .A(n31559), .B(n31558), .Z(n31560) );
  NANDN U48879 ( .A(n31561), .B(n31560), .Z(n31563) );
  OR U48880 ( .A(n31563), .B(n31562), .Z(n31564) );
  NAND U48881 ( .A(n31565), .B(n31564), .Z(n31569) );
  AND U48882 ( .A(n31567), .B(n31566), .Z(n31568) );
  NAND U48883 ( .A(n31569), .B(n31568), .Z(n31570) );
  NAND U48884 ( .A(n52912), .B(n31570), .Z(n31574) );
  IV U48885 ( .A(n31571), .Z(n52913) );
  NOR U48886 ( .A(n52913), .B(n31572), .Z(n31573) );
  NAND U48887 ( .A(n31574), .B(n31573), .Z(n31575) );
  AND U48888 ( .A(n31576), .B(n31575), .Z(n31577) );
  NAND U48889 ( .A(n52914), .B(n31577), .Z(n31579) );
  ANDN U48890 ( .B(n31579), .A(n31578), .Z(n31580) );
  NANDN U48891 ( .A(n31581), .B(n31580), .Z(n31585) );
  AND U48892 ( .A(n31583), .B(n31582), .Z(n31584) );
  NAND U48893 ( .A(n31585), .B(n31584), .Z(n31586) );
  NANDN U48894 ( .A(n31587), .B(n31586), .Z(n31589) );
  OR U48895 ( .A(n31589), .B(n31588), .Z(n31590) );
  NAND U48896 ( .A(n31591), .B(n31590), .Z(n31595) );
  AND U48897 ( .A(n31593), .B(n31592), .Z(n31594) );
  NAND U48898 ( .A(n31595), .B(n31594), .Z(n31596) );
  NANDN U48899 ( .A(n31597), .B(n31596), .Z(n31598) );
  OR U48900 ( .A(n31598), .B(n52921), .Z(n31599) );
  AND U48901 ( .A(n31599), .B(n52922), .Z(n31600) );
  NANDN U48902 ( .A(n31601), .B(n31600), .Z(n31602) );
  AND U48903 ( .A(n52923), .B(n31602), .Z(n31603) );
  NOR U48904 ( .A(n52924), .B(n31603), .Z(n31604) );
  NANDN U48905 ( .A(n31605), .B(n31604), .Z(n31606) );
  AND U48906 ( .A(n31606), .B(n52925), .Z(n31607) );
  OR U48907 ( .A(n31608), .B(n31607), .Z(n31610) );
  IV U48908 ( .A(n31609), .Z(n52927) );
  AND U48909 ( .A(n31610), .B(n52927), .Z(n31612) );
  IV U48910 ( .A(n31611), .Z(n52928) );
  OR U48911 ( .A(n31612), .B(n52928), .Z(n31613) );
  NAND U48912 ( .A(n52930), .B(n31613), .Z(n31614) );
  NANDN U48913 ( .A(n52931), .B(n31614), .Z(n31615) );
  NANDN U48914 ( .A(n31616), .B(n31615), .Z(n31617) );
  AND U48915 ( .A(n52932), .B(n31617), .Z(n31623) );
  NANDN U48916 ( .A(n31619), .B(n31618), .Z(n31621) );
  ANDN U48917 ( .B(n31621), .A(n31620), .Z(n31622) );
  OR U48918 ( .A(n31623), .B(n31622), .Z(n31624) );
  NAND U48919 ( .A(n52934), .B(n31624), .Z(n31625) );
  NAND U48920 ( .A(n52935), .B(n31625), .Z(n31628) );
  AND U48921 ( .A(n31626), .B(n52359), .Z(n31627) );
  NAND U48922 ( .A(n31628), .B(n31627), .Z(n31629) );
  NANDN U48923 ( .A(n31630), .B(n31629), .Z(n31631) );
  OR U48924 ( .A(n31631), .B(n52358), .Z(n31632) );
  AND U48925 ( .A(n31633), .B(n31632), .Z(n31637) );
  NAND U48926 ( .A(n31635), .B(n31634), .Z(n31636) );
  OR U48927 ( .A(n31637), .B(n31636), .Z(n31638) );
  AND U48928 ( .A(n31639), .B(n31638), .Z(n31641) );
  NAND U48929 ( .A(n31641), .B(n31640), .Z(n31643) );
  ANDN U48930 ( .B(n31643), .A(n31642), .Z(n31644) );
  NANDN U48931 ( .A(n31645), .B(n31644), .Z(n31649) );
  AND U48932 ( .A(n31647), .B(n31646), .Z(n31648) );
  NAND U48933 ( .A(n31649), .B(n31648), .Z(n31650) );
  NANDN U48934 ( .A(n31651), .B(n31650), .Z(n31652) );
  OR U48935 ( .A(n31652), .B(n52943), .Z(n31653) );
  AND U48936 ( .A(n31654), .B(n31653), .Z(n31657) );
  NAND U48937 ( .A(n31656), .B(n31655), .Z(n52357) );
  OR U48938 ( .A(n31657), .B(n52357), .Z(n31658) );
  AND U48939 ( .A(n31659), .B(n31658), .Z(n31660) );
  NAND U48940 ( .A(n52356), .B(n31660), .Z(n31662) );
  ANDN U48941 ( .B(n31662), .A(n31661), .Z(n31663) );
  NANDN U48942 ( .A(n52947), .B(n31663), .Z(n31667) );
  AND U48943 ( .A(n31665), .B(n31664), .Z(n31666) );
  NAND U48944 ( .A(n31667), .B(n31666), .Z(n31668) );
  NANDN U48945 ( .A(n31669), .B(n31668), .Z(n31671) );
  OR U48946 ( .A(n31671), .B(n31670), .Z(n31672) );
  NAND U48947 ( .A(n31673), .B(n31672), .Z(n31677) );
  AND U48948 ( .A(n31675), .B(n31674), .Z(n31676) );
  NAND U48949 ( .A(n31677), .B(n31676), .Z(n31678) );
  NANDN U48950 ( .A(n31679), .B(n31678), .Z(n31681) );
  OR U48951 ( .A(n31681), .B(n31680), .Z(n31682) );
  NAND U48952 ( .A(n31683), .B(n31682), .Z(n31684) );
  NANDN U48953 ( .A(n31685), .B(n31684), .Z(n31689) );
  AND U48954 ( .A(n31687), .B(n31686), .Z(n31688) );
  NAND U48955 ( .A(n31689), .B(n31688), .Z(n31690) );
  NANDN U48956 ( .A(n31691), .B(n31690), .Z(n31693) );
  OR U48957 ( .A(n31693), .B(n31692), .Z(n31694) );
  NAND U48958 ( .A(n31695), .B(n31694), .Z(n31696) );
  NANDN U48959 ( .A(n31697), .B(n31696), .Z(n31701) );
  AND U48960 ( .A(n31699), .B(n31698), .Z(n31700) );
  NAND U48961 ( .A(n31701), .B(n31700), .Z(n31702) );
  NANDN U48962 ( .A(n31703), .B(n31702), .Z(n31705) );
  OR U48963 ( .A(n31705), .B(n31704), .Z(n31706) );
  NAND U48964 ( .A(n31707), .B(n31706), .Z(n31708) );
  NANDN U48965 ( .A(n31709), .B(n31708), .Z(n31712) );
  AND U48966 ( .A(n31710), .B(n52966), .Z(n31711) );
  NAND U48967 ( .A(n31712), .B(n31711), .Z(n31713) );
  NANDN U48968 ( .A(n52967), .B(n31713), .Z(n31714) );
  OR U48969 ( .A(n31715), .B(n31714), .Z(n31718) );
  AND U48970 ( .A(n31717), .B(n31716), .Z(n52355) );
  AND U48971 ( .A(n31718), .B(n52355), .Z(n31720) );
  NAND U48972 ( .A(n52969), .B(n52968), .Z(n31719) );
  OR U48973 ( .A(n31720), .B(n31719), .Z(n31721) );
  AND U48974 ( .A(n31722), .B(n31721), .Z(n31724) );
  NANDN U48975 ( .A(x[966]), .B(y[966]), .Z(n31723) );
  NAND U48976 ( .A(n31724), .B(n31723), .Z(n31726) );
  ANDN U48977 ( .B(n31726), .A(n31725), .Z(n31727) );
  NANDN U48978 ( .A(n31728), .B(n31727), .Z(n31732) );
  AND U48979 ( .A(n31730), .B(n31729), .Z(n31731) );
  NAND U48980 ( .A(n31732), .B(n31731), .Z(n31733) );
  NANDN U48981 ( .A(n31734), .B(n31733), .Z(n31736) );
  OR U48982 ( .A(n31736), .B(n31735), .Z(n31737) );
  AND U48983 ( .A(n31738), .B(n31737), .Z(n31740) );
  NOR U48984 ( .A(n31740), .B(n31739), .Z(n31741) );
  NANDN U48985 ( .A(n31742), .B(n31741), .Z(n31743) );
  AND U48986 ( .A(n31744), .B(n31743), .Z(n31745) );
  NAND U48987 ( .A(n31745), .B(n52977), .Z(n31746) );
  NANDN U48988 ( .A(n31747), .B(n31746), .Z(n31748) );
  AND U48989 ( .A(n52980), .B(n31748), .Z(n31749) );
  ANDN U48990 ( .B(n52981), .A(n31749), .Z(n31750) );
  NANDN U48991 ( .A(n31751), .B(n31750), .Z(n31752) );
  AND U48992 ( .A(n31753), .B(n31752), .Z(n31754) );
  NAND U48993 ( .A(n31754), .B(n52982), .Z(n31756) );
  ANDN U48994 ( .B(n31756), .A(n31755), .Z(n31757) );
  NANDN U48995 ( .A(n31758), .B(n31757), .Z(n31762) );
  AND U48996 ( .A(n31760), .B(n31759), .Z(n31761) );
  NAND U48997 ( .A(n31762), .B(n31761), .Z(n31763) );
  NANDN U48998 ( .A(n31764), .B(n31763), .Z(n31766) );
  OR U48999 ( .A(n31766), .B(n31765), .Z(n31767) );
  NAND U49000 ( .A(n31768), .B(n31767), .Z(n31772) );
  AND U49001 ( .A(n31770), .B(n31769), .Z(n31771) );
  NAND U49002 ( .A(n31772), .B(n31771), .Z(n31773) );
  NANDN U49003 ( .A(n31774), .B(n31773), .Z(n31775) );
  OR U49004 ( .A(n52990), .B(n31775), .Z(n31776) );
  AND U49005 ( .A(n31776), .B(n52991), .Z(n31777) );
  NANDN U49006 ( .A(n31778), .B(n31777), .Z(n31779) );
  AND U49007 ( .A(n31780), .B(n31779), .Z(n31781) );
  NAND U49008 ( .A(n31781), .B(n52992), .Z(n31783) );
  ANDN U49009 ( .B(n31783), .A(n31782), .Z(n31784) );
  NAND U49010 ( .A(n52993), .B(n31784), .Z(n31788) );
  AND U49011 ( .A(n31786), .B(n31785), .Z(n31787) );
  NAND U49012 ( .A(n31788), .B(n31787), .Z(n31789) );
  NANDN U49013 ( .A(n31790), .B(n31789), .Z(n31791) );
  OR U49014 ( .A(n31792), .B(n31791), .Z(n31793) );
  AND U49015 ( .A(n31794), .B(n31793), .Z(n31795) );
  NANDN U49016 ( .A(n31796), .B(n31795), .Z(n31797) );
  AND U49017 ( .A(n31798), .B(n31797), .Z(n31800) );
  NAND U49018 ( .A(n31800), .B(n31799), .Z(n31802) );
  ANDN U49019 ( .B(n31802), .A(n31801), .Z(n31803) );
  NANDN U49020 ( .A(n31804), .B(n31803), .Z(n31808) );
  AND U49021 ( .A(n31806), .B(n31805), .Z(n31807) );
  NAND U49022 ( .A(n31808), .B(n31807), .Z(n31809) );
  NANDN U49023 ( .A(n31810), .B(n31809), .Z(n31811) );
  OR U49024 ( .A(n31811), .B(n53003), .Z(n31812) );
  AND U49025 ( .A(n31813), .B(n31812), .Z(n31816) );
  NAND U49026 ( .A(n31815), .B(n31814), .Z(n52354) );
  OR U49027 ( .A(n31816), .B(n52354), .Z(n31817) );
  AND U49028 ( .A(n53005), .B(n31817), .Z(n31818) );
  NAND U49029 ( .A(n52353), .B(n31818), .Z(n31820) );
  ANDN U49030 ( .B(y[996]), .A(x[996]), .Z(n31819) );
  ANDN U49031 ( .B(n31820), .A(n31819), .Z(n31821) );
  NANDN U49032 ( .A(n31822), .B(n31821), .Z(n31826) );
  AND U49033 ( .A(n31824), .B(n31823), .Z(n31825) );
  NAND U49034 ( .A(n31826), .B(n31825), .Z(n31827) );
  NANDN U49035 ( .A(n31828), .B(n31827), .Z(n31830) );
  OR U49036 ( .A(n31830), .B(n31829), .Z(n31831) );
  NAND U49037 ( .A(n31832), .B(n31831), .Z(n31836) );
  AND U49038 ( .A(n31834), .B(n31833), .Z(n31835) );
  NAND U49039 ( .A(n31836), .B(n31835), .Z(n31837) );
  NANDN U49040 ( .A(n31838), .B(n31837), .Z(n31840) );
  OR U49041 ( .A(n31840), .B(n31839), .Z(n31841) );
  NAND U49042 ( .A(n31842), .B(n31841), .Z(n31843) );
  NANDN U49043 ( .A(n31844), .B(n31843), .Z(n31848) );
  AND U49044 ( .A(n31846), .B(n31845), .Z(n31847) );
  NAND U49045 ( .A(n31848), .B(n31847), .Z(n31849) );
  NANDN U49046 ( .A(n31850), .B(n31849), .Z(n31851) );
  OR U49047 ( .A(n31852), .B(n31851), .Z(n31853) );
  AND U49048 ( .A(n31854), .B(n31853), .Z(n31855) );
  NAND U49049 ( .A(n31856), .B(n31855), .Z(n31857) );
  NAND U49050 ( .A(n31858), .B(n31857), .Z(n31859) );
  AND U49051 ( .A(n31860), .B(n31859), .Z(n31861) );
  OR U49052 ( .A(n31861), .B(n53019), .Z(n31862) );
  NAND U49053 ( .A(n53020), .B(n31862), .Z(n31863) );
  NANDN U49054 ( .A(n53021), .B(n31863), .Z(n31864) );
  AND U49055 ( .A(n53022), .B(n31864), .Z(n31865) );
  OR U49056 ( .A(n31866), .B(n31865), .Z(n31867) );
  NAND U49057 ( .A(n53024), .B(n31867), .Z(n31868) );
  NANDN U49058 ( .A(n31869), .B(n31868), .Z(n31871) );
  IV U49059 ( .A(n31870), .Z(n53025) );
  OR U49060 ( .A(n31871), .B(n53025), .Z(n31872) );
  AND U49061 ( .A(n53026), .B(n31872), .Z(n31873) );
  NOR U49062 ( .A(n53027), .B(n31873), .Z(n31874) );
  NANDN U49063 ( .A(n31875), .B(n31874), .Z(n31876) );
  AND U49064 ( .A(n31877), .B(n31876), .Z(n31878) );
  NAND U49065 ( .A(n53028), .B(n31878), .Z(n31880) );
  ANDN U49066 ( .B(n31880), .A(n31879), .Z(n31881) );
  NANDN U49067 ( .A(n31882), .B(n31881), .Z(n31886) );
  AND U49068 ( .A(n31884), .B(n31883), .Z(n31885) );
  NAND U49069 ( .A(n31886), .B(n31885), .Z(n31887) );
  NANDN U49070 ( .A(n31888), .B(n31887), .Z(n31890) );
  OR U49071 ( .A(n31890), .B(n31889), .Z(n31891) );
  NAND U49072 ( .A(n31892), .B(n31891), .Z(n31896) );
  AND U49073 ( .A(n31894), .B(n31893), .Z(n31895) );
  NAND U49074 ( .A(n31896), .B(n31895), .Z(n31897) );
  NANDN U49075 ( .A(n31898), .B(n31897), .Z(n31899) );
  OR U49076 ( .A(n31899), .B(n53036), .Z(n31900) );
  NAND U49077 ( .A(n31901), .B(n31900), .Z(n31902) );
  NANDN U49078 ( .A(n53038), .B(n31902), .Z(n31905) );
  AND U49079 ( .A(n31903), .B(n53039), .Z(n31904) );
  NAND U49080 ( .A(n31905), .B(n31904), .Z(n31906) );
  NANDN U49081 ( .A(n53040), .B(n31906), .Z(n31907) );
  OR U49082 ( .A(n31908), .B(n31907), .Z(n31909) );
  AND U49083 ( .A(n31910), .B(n31909), .Z(n31911) );
  NANDN U49084 ( .A(n31912), .B(n31911), .Z(n31913) );
  AND U49085 ( .A(n31914), .B(n31913), .Z(n31916) );
  NOR U49086 ( .A(n31916), .B(n31915), .Z(n31917) );
  NANDN U49087 ( .A(n31918), .B(n31917), .Z(n31919) );
  AND U49088 ( .A(n31920), .B(n31919), .Z(n31921) );
  NANDN U49089 ( .A(n31922), .B(n31921), .Z(n31923) );
  NAND U49090 ( .A(n31924), .B(n31923), .Z(n31925) );
  NANDN U49091 ( .A(n31926), .B(n31925), .Z(n31927) );
  OR U49092 ( .A(n31927), .B(n53048), .Z(n31928) );
  AND U49093 ( .A(n31929), .B(n31928), .Z(n31932) );
  NAND U49094 ( .A(n31931), .B(n31930), .Z(n53050) );
  OR U49095 ( .A(n31932), .B(n53050), .Z(n31933) );
  AND U49096 ( .A(n53052), .B(n31933), .Z(n31934) );
  NAND U49097 ( .A(n31934), .B(n53051), .Z(n31936) );
  ANDN U49098 ( .B(y[1036]), .A(x[1036]), .Z(n31935) );
  ANDN U49099 ( .B(n31936), .A(n31935), .Z(n31937) );
  NANDN U49100 ( .A(n31938), .B(n31937), .Z(n31942) );
  AND U49101 ( .A(n31940), .B(n31939), .Z(n31941) );
  NAND U49102 ( .A(n31942), .B(n31941), .Z(n31943) );
  NANDN U49103 ( .A(n31944), .B(n31943), .Z(n31946) );
  OR U49104 ( .A(n31946), .B(n31945), .Z(n31947) );
  NAND U49105 ( .A(n31948), .B(n31947), .Z(n31952) );
  AND U49106 ( .A(n31950), .B(n31949), .Z(n31951) );
  NAND U49107 ( .A(n31952), .B(n31951), .Z(n31953) );
  NANDN U49108 ( .A(n31954), .B(n31953), .Z(n31955) );
  OR U49109 ( .A(n31956), .B(n31955), .Z(n31957) );
  AND U49110 ( .A(n31958), .B(n31957), .Z(n31959) );
  NAND U49111 ( .A(n31959), .B(n53061), .Z(n31961) );
  IV U49112 ( .A(n31960), .Z(n53062) );
  ANDN U49113 ( .B(n31961), .A(n53062), .Z(n31962) );
  NANDN U49114 ( .A(n31963), .B(n31962), .Z(n31966) );
  AND U49115 ( .A(n53063), .B(n31964), .Z(n31965) );
  NAND U49116 ( .A(n31966), .B(n31965), .Z(n31967) );
  NAND U49117 ( .A(n53064), .B(n31967), .Z(n31969) );
  OR U49118 ( .A(n31969), .B(n31968), .Z(n31970) );
  AND U49119 ( .A(n31971), .B(n31970), .Z(n31972) );
  NANDN U49120 ( .A(n31973), .B(n31972), .Z(n31974) );
  AND U49121 ( .A(n31975), .B(n31974), .Z(n31977) );
  NAND U49122 ( .A(n31977), .B(n31976), .Z(n31979) );
  ANDN U49123 ( .B(n31979), .A(n31978), .Z(n31980) );
  NANDN U49124 ( .A(n31981), .B(n31980), .Z(n31985) );
  AND U49125 ( .A(n31983), .B(n31982), .Z(n31984) );
  NAND U49126 ( .A(n31985), .B(n31984), .Z(n31986) );
  NANDN U49127 ( .A(n31987), .B(n31986), .Z(n31988) );
  OR U49128 ( .A(n31989), .B(n31988), .Z(n31990) );
  AND U49129 ( .A(n31991), .B(n31990), .Z(n31992) );
  NANDN U49130 ( .A(n31993), .B(n31992), .Z(n31994) );
  AND U49131 ( .A(n31995), .B(n31994), .Z(n31997) );
  NAND U49132 ( .A(n31997), .B(n31996), .Z(n31999) );
  ANDN U49133 ( .B(n31999), .A(n31998), .Z(n32000) );
  NANDN U49134 ( .A(n32001), .B(n32000), .Z(n32005) );
  AND U49135 ( .A(n32003), .B(n32002), .Z(n32004) );
  NAND U49136 ( .A(n32005), .B(n32004), .Z(n32006) );
  NANDN U49137 ( .A(n32007), .B(n32006), .Z(n32009) );
  OR U49138 ( .A(n32009), .B(n32008), .Z(n32010) );
  AND U49139 ( .A(n32011), .B(n32010), .Z(n32015) );
  NAND U49140 ( .A(n32013), .B(n32012), .Z(n32014) );
  OR U49141 ( .A(n32015), .B(n32014), .Z(n32016) );
  AND U49142 ( .A(n32017), .B(n32016), .Z(n32019) );
  NAND U49143 ( .A(n32019), .B(n32018), .Z(n32021) );
  ANDN U49144 ( .B(n32021), .A(n32020), .Z(n32022) );
  NANDN U49145 ( .A(n32023), .B(n32022), .Z(n32027) );
  AND U49146 ( .A(n32025), .B(n32024), .Z(n32026) );
  NAND U49147 ( .A(n32027), .B(n32026), .Z(n32028) );
  NANDN U49148 ( .A(n32029), .B(n32028), .Z(n32030) );
  OR U49149 ( .A(n32031), .B(n32030), .Z(n32032) );
  AND U49150 ( .A(n32033), .B(n32032), .Z(n32034) );
  NANDN U49151 ( .A(n53080), .B(n32034), .Z(n32035) );
  NAND U49152 ( .A(n32036), .B(n32035), .Z(n32037) );
  NANDN U49153 ( .A(n53082), .B(n32037), .Z(n32040) );
  AND U49154 ( .A(n32038), .B(n53083), .Z(n32039) );
  NAND U49155 ( .A(n32040), .B(n32039), .Z(n32041) );
  NANDN U49156 ( .A(n53084), .B(n32041), .Z(n32043) );
  IV U49157 ( .A(n32042), .Z(n53087) );
  OR U49158 ( .A(n32043), .B(n53087), .Z(n32044) );
  AND U49159 ( .A(n32045), .B(n32044), .Z(n32046) );
  NAND U49160 ( .A(n53088), .B(n32046), .Z(n32047) );
  NANDN U49161 ( .A(n53089), .B(n32047), .Z(n32048) );
  AND U49162 ( .A(n53090), .B(n32048), .Z(n32051) );
  NAND U49163 ( .A(n32050), .B(n32049), .Z(n53091) );
  OR U49164 ( .A(n32051), .B(n53091), .Z(n32052) );
  AND U49165 ( .A(n32053), .B(n32052), .Z(n32054) );
  NAND U49166 ( .A(n32054), .B(n53092), .Z(n32056) );
  ANDN U49167 ( .B(n32056), .A(n32055), .Z(n32057) );
  NANDN U49168 ( .A(n53093), .B(n32057), .Z(n32061) );
  AND U49169 ( .A(n32059), .B(n32058), .Z(n32060) );
  NAND U49170 ( .A(n32061), .B(n32060), .Z(n32062) );
  NANDN U49171 ( .A(n32063), .B(n32062), .Z(n32065) );
  OR U49172 ( .A(n32065), .B(n32064), .Z(n32066) );
  NAND U49173 ( .A(n32067), .B(n32066), .Z(n32071) );
  AND U49174 ( .A(n32069), .B(n32068), .Z(n32070) );
  NAND U49175 ( .A(n32071), .B(n32070), .Z(n32072) );
  NANDN U49176 ( .A(n32073), .B(n32072), .Z(n32075) );
  OR U49177 ( .A(n32075), .B(n32074), .Z(n32076) );
  NAND U49178 ( .A(n32077), .B(n32076), .Z(n32078) );
  NANDN U49179 ( .A(n32079), .B(n32078), .Z(n32083) );
  AND U49180 ( .A(n32081), .B(n32080), .Z(n32082) );
  NAND U49181 ( .A(n32083), .B(n32082), .Z(n32084) );
  NANDN U49182 ( .A(n32085), .B(n32084), .Z(n32087) );
  OR U49183 ( .A(n32087), .B(n32086), .Z(n32088) );
  NAND U49184 ( .A(n32089), .B(n32088), .Z(n32090) );
  NANDN U49185 ( .A(n32091), .B(n32090), .Z(n32095) );
  AND U49186 ( .A(n32093), .B(n32092), .Z(n32094) );
  NAND U49187 ( .A(n32095), .B(n32094), .Z(n32096) );
  NANDN U49188 ( .A(n32097), .B(n32096), .Z(n32099) );
  OR U49189 ( .A(n32099), .B(n32098), .Z(n32100) );
  NAND U49190 ( .A(n32101), .B(n32100), .Z(n32102) );
  NANDN U49191 ( .A(n32103), .B(n32102), .Z(n32107) );
  AND U49192 ( .A(n32105), .B(n32104), .Z(n32106) );
  NAND U49193 ( .A(n32107), .B(n32106), .Z(n32108) );
  NANDN U49194 ( .A(n32109), .B(n32108), .Z(n32111) );
  OR U49195 ( .A(n32111), .B(n32110), .Z(n32112) );
  NAND U49196 ( .A(n32113), .B(n32112), .Z(n32114) );
  NANDN U49197 ( .A(n32115), .B(n32114), .Z(n32118) );
  AND U49198 ( .A(n32116), .B(n53116), .Z(n32117) );
  NAND U49199 ( .A(n32118), .B(n32117), .Z(n32119) );
  NANDN U49200 ( .A(n53117), .B(n32119), .Z(n32120) );
  OR U49201 ( .A(n32121), .B(n32120), .Z(n32122) );
  AND U49202 ( .A(n32123), .B(n32122), .Z(n32124) );
  NAND U49203 ( .A(n52346), .B(n32124), .Z(n32126) );
  ANDN U49204 ( .B(n32126), .A(n32125), .Z(n32127) );
  NANDN U49205 ( .A(n53118), .B(n32127), .Z(n32131) );
  AND U49206 ( .A(n32129), .B(n32128), .Z(n32130) );
  NAND U49207 ( .A(n32131), .B(n32130), .Z(n32132) );
  NANDN U49208 ( .A(n32133), .B(n32132), .Z(n32134) );
  OR U49209 ( .A(n32135), .B(n32134), .Z(n32136) );
  AND U49210 ( .A(n32137), .B(n32136), .Z(n32138) );
  NANDN U49211 ( .A(n32139), .B(n32138), .Z(n32140) );
  AND U49212 ( .A(n32141), .B(n32140), .Z(n32143) );
  NAND U49213 ( .A(n32143), .B(n32142), .Z(n32145) );
  ANDN U49214 ( .B(n32145), .A(n32144), .Z(n32146) );
  NANDN U49215 ( .A(n32147), .B(n32146), .Z(n32151) );
  AND U49216 ( .A(n32149), .B(n32148), .Z(n32150) );
  NAND U49217 ( .A(n32151), .B(n32150), .Z(n32152) );
  NANDN U49218 ( .A(n32153), .B(n32152), .Z(n32155) );
  OR U49219 ( .A(n32155), .B(n32154), .Z(n32156) );
  AND U49220 ( .A(n32157), .B(n32156), .Z(n32161) );
  NAND U49221 ( .A(n32159), .B(n32158), .Z(n32160) );
  OR U49222 ( .A(n32161), .B(n32160), .Z(n32162) );
  AND U49223 ( .A(n32163), .B(n32162), .Z(n32165) );
  NAND U49224 ( .A(n32165), .B(n32164), .Z(n32167) );
  ANDN U49225 ( .B(n32167), .A(n32166), .Z(n32168) );
  NANDN U49226 ( .A(n32169), .B(n32168), .Z(n32173) );
  AND U49227 ( .A(n32171), .B(n32170), .Z(n32172) );
  NAND U49228 ( .A(n32173), .B(n32172), .Z(n32174) );
  NANDN U49229 ( .A(n32175), .B(n32174), .Z(n32176) );
  OR U49230 ( .A(n32176), .B(n53146), .Z(n32177) );
  NAND U49231 ( .A(n32178), .B(n32177), .Z(n32179) );
  NANDN U49232 ( .A(n53150), .B(n32179), .Z(n32180) );
  NAND U49233 ( .A(n53152), .B(n32180), .Z(n32181) );
  ANDN U49234 ( .B(y[1112]), .A(x[1112]), .Z(n53154) );
  ANDN U49235 ( .B(n32181), .A(n53154), .Z(n32182) );
  NANDN U49236 ( .A(n32183), .B(n32182), .Z(n32186) );
  AND U49237 ( .A(n32184), .B(n53156), .Z(n32185) );
  NAND U49238 ( .A(n32186), .B(n32185), .Z(n32187) );
  NANDN U49239 ( .A(n32188), .B(n32187), .Z(n32189) );
  OR U49240 ( .A(n32190), .B(n32189), .Z(n32191) );
  AND U49241 ( .A(n32192), .B(n32191), .Z(n32194) );
  NAND U49242 ( .A(n32194), .B(n32193), .Z(n32196) );
  ANDN U49243 ( .B(n32196), .A(n32195), .Z(n32197) );
  NANDN U49244 ( .A(n32198), .B(n32197), .Z(n32202) );
  AND U49245 ( .A(n32200), .B(n32199), .Z(n32201) );
  NAND U49246 ( .A(n32202), .B(n32201), .Z(n32203) );
  NANDN U49247 ( .A(n32204), .B(n32203), .Z(n32205) );
  OR U49248 ( .A(n32205), .B(n53163), .Z(n32206) );
  NAND U49249 ( .A(n32207), .B(n32206), .Z(n32208) );
  NAND U49250 ( .A(n53165), .B(n32208), .Z(n32211) );
  AND U49251 ( .A(n32209), .B(n53166), .Z(n32210) );
  NAND U49252 ( .A(n32211), .B(n32210), .Z(n32212) );
  NANDN U49253 ( .A(n32213), .B(n32212), .Z(n32214) );
  OR U49254 ( .A(n32215), .B(n32214), .Z(n32216) );
  AND U49255 ( .A(n32217), .B(n32216), .Z(n32218) );
  NANDN U49256 ( .A(n32219), .B(n32218), .Z(n32220) );
  AND U49257 ( .A(n32221), .B(n32220), .Z(n32222) );
  ANDN U49258 ( .B(n32223), .A(n32222), .Z(n32224) );
  NAND U49259 ( .A(n32225), .B(n32224), .Z(n32226) );
  NANDN U49260 ( .A(n32227), .B(n32226), .Z(n32229) );
  OR U49261 ( .A(n32229), .B(n32228), .Z(n32230) );
  NAND U49262 ( .A(n32231), .B(n32230), .Z(n32232) );
  NANDN U49263 ( .A(n32233), .B(n32232), .Z(n32237) );
  AND U49264 ( .A(n32235), .B(n32234), .Z(n32236) );
  NAND U49265 ( .A(n32237), .B(n32236), .Z(n32238) );
  NANDN U49266 ( .A(n32239), .B(n32238), .Z(n32241) );
  OR U49267 ( .A(n32241), .B(n32240), .Z(n32242) );
  NAND U49268 ( .A(n32243), .B(n32242), .Z(n32244) );
  NANDN U49269 ( .A(n32245), .B(n32244), .Z(n32249) );
  AND U49270 ( .A(n32247), .B(n32246), .Z(n32248) );
  NAND U49271 ( .A(n32249), .B(n32248), .Z(n32250) );
  NANDN U49272 ( .A(n32251), .B(n32250), .Z(n32252) );
  OR U49273 ( .A(n32253), .B(n32252), .Z(n32254) );
  AND U49274 ( .A(n32255), .B(n32254), .Z(n32256) );
  NANDN U49275 ( .A(n32257), .B(n32256), .Z(n32258) );
  AND U49276 ( .A(n32259), .B(n32258), .Z(n32261) );
  NOR U49277 ( .A(n32261), .B(n32260), .Z(n32262) );
  NANDN U49278 ( .A(n32263), .B(n32262), .Z(n32264) );
  AND U49279 ( .A(n32265), .B(n32264), .Z(n32267) );
  AND U49280 ( .A(n32267), .B(n32266), .Z(n32271) );
  AND U49281 ( .A(n32269), .B(n32268), .Z(n32270) );
  NANDN U49282 ( .A(n32271), .B(n32270), .Z(n32272) );
  NAND U49283 ( .A(n32273), .B(n32272), .Z(n32277) );
  AND U49284 ( .A(n32275), .B(n32274), .Z(n32276) );
  NAND U49285 ( .A(n32277), .B(n32276), .Z(n32278) );
  NANDN U49286 ( .A(n32279), .B(n32278), .Z(n32280) );
  OR U49287 ( .A(n32281), .B(n32280), .Z(n32282) );
  AND U49288 ( .A(n32283), .B(n32282), .Z(n32285) );
  NAND U49289 ( .A(n32285), .B(n32284), .Z(n32287) );
  ANDN U49290 ( .B(n32287), .A(n32286), .Z(n32288) );
  NANDN U49291 ( .A(n53184), .B(n32288), .Z(n32291) );
  AND U49292 ( .A(n32289), .B(n53185), .Z(n32290) );
  NAND U49293 ( .A(n32291), .B(n32290), .Z(n32292) );
  NANDN U49294 ( .A(n53186), .B(n32292), .Z(n32295) );
  AND U49295 ( .A(n32293), .B(n53187), .Z(n32294) );
  NAND U49296 ( .A(n32295), .B(n32294), .Z(n32296) );
  NANDN U49297 ( .A(n32297), .B(n32296), .Z(n32298) );
  OR U49298 ( .A(n32298), .B(n53188), .Z(n32299) );
  NAND U49299 ( .A(n32300), .B(n32299), .Z(n32304) );
  AND U49300 ( .A(n32302), .B(n32301), .Z(n32303) );
  NAND U49301 ( .A(n32304), .B(n32303), .Z(n32305) );
  NANDN U49302 ( .A(n32306), .B(n32305), .Z(n32308) );
  OR U49303 ( .A(n32308), .B(n32307), .Z(n32309) );
  NAND U49304 ( .A(n32310), .B(n32309), .Z(n32311) );
  NANDN U49305 ( .A(n32312), .B(n32311), .Z(n32316) );
  AND U49306 ( .A(n32314), .B(n32313), .Z(n32315) );
  NAND U49307 ( .A(n32316), .B(n32315), .Z(n32317) );
  NANDN U49308 ( .A(n32318), .B(n32317), .Z(n32320) );
  OR U49309 ( .A(n32320), .B(n32319), .Z(n32321) );
  NAND U49310 ( .A(n32322), .B(n32321), .Z(n32323) );
  NANDN U49311 ( .A(n32324), .B(n32323), .Z(n32328) );
  AND U49312 ( .A(n32326), .B(n32325), .Z(n32327) );
  NAND U49313 ( .A(n32328), .B(n32327), .Z(n32329) );
  NANDN U49314 ( .A(n32330), .B(n32329), .Z(n32331) );
  OR U49315 ( .A(n32332), .B(n32331), .Z(n32333) );
  AND U49316 ( .A(n32334), .B(n32333), .Z(n32335) );
  NAND U49317 ( .A(n53202), .B(n32335), .Z(n32337) );
  ANDN U49318 ( .B(n32337), .A(n32336), .Z(n32338) );
  NANDN U49319 ( .A(n53203), .B(n32338), .Z(n32339) );
  NAND U49320 ( .A(n53204), .B(n32339), .Z(n32340) );
  NANDN U49321 ( .A(n53205), .B(n32340), .Z(n32341) );
  AND U49322 ( .A(n32342), .B(n32341), .Z(n32343) );
  NAND U49323 ( .A(n32343), .B(n53206), .Z(n32345) );
  ANDN U49324 ( .B(n32345), .A(n32344), .Z(n32346) );
  NANDN U49325 ( .A(n53207), .B(n32346), .Z(n32350) );
  NANDN U49326 ( .A(x[1166]), .B(y[1166]), .Z(n32347) );
  AND U49327 ( .A(n32348), .B(n32347), .Z(n32349) );
  NAND U49328 ( .A(n32350), .B(n32349), .Z(n32351) );
  NANDN U49329 ( .A(n32352), .B(n32351), .Z(n32354) );
  OR U49330 ( .A(n32354), .B(n32353), .Z(n32355) );
  NAND U49331 ( .A(n32356), .B(n32355), .Z(n32360) );
  AND U49332 ( .A(n32358), .B(n32357), .Z(n32359) );
  NAND U49333 ( .A(n32360), .B(n32359), .Z(n32361) );
  NANDN U49334 ( .A(n32362), .B(n32361), .Z(n32363) );
  OR U49335 ( .A(n32363), .B(n53214), .Z(n32364) );
  NAND U49336 ( .A(n32365), .B(n32364), .Z(n32366) );
  NANDN U49337 ( .A(n53216), .B(n32366), .Z(n32369) );
  AND U49338 ( .A(n32367), .B(n53217), .Z(n32368) );
  NAND U49339 ( .A(n32369), .B(n32368), .Z(n32370) );
  NANDN U49340 ( .A(n32371), .B(n32370), .Z(n32372) );
  OR U49341 ( .A(n32372), .B(n53218), .Z(n32373) );
  NAND U49342 ( .A(n32374), .B(n32373), .Z(n32378) );
  AND U49343 ( .A(n32376), .B(n32375), .Z(n32377) );
  NAND U49344 ( .A(n32378), .B(n32377), .Z(n32379) );
  NANDN U49345 ( .A(n32380), .B(n32379), .Z(n32382) );
  OR U49346 ( .A(n32382), .B(n32381), .Z(n32383) );
  NAND U49347 ( .A(n32384), .B(n32383), .Z(n32385) );
  NANDN U49348 ( .A(n32386), .B(n32385), .Z(n32387) );
  AND U49349 ( .A(n32388), .B(n32387), .Z(n32389) );
  NAND U49350 ( .A(n32390), .B(n32389), .Z(n32391) );
  NANDN U49351 ( .A(n32392), .B(n32391), .Z(n32393) );
  OR U49352 ( .A(n32394), .B(n32393), .Z(n32395) );
  AND U49353 ( .A(n32396), .B(n32395), .Z(n32397) );
  NANDN U49354 ( .A(n32398), .B(n32397), .Z(n32399) );
  AND U49355 ( .A(n32400), .B(n32399), .Z(n32402) );
  NOR U49356 ( .A(n32402), .B(n32401), .Z(n32403) );
  NANDN U49357 ( .A(n32404), .B(n32403), .Z(n32405) );
  AND U49358 ( .A(n32406), .B(n32405), .Z(n32407) );
  NANDN U49359 ( .A(n53231), .B(n32407), .Z(n32408) );
  AND U49360 ( .A(n32409), .B(n32408), .Z(n32410) );
  NAND U49361 ( .A(n32410), .B(n53232), .Z(n32411) );
  NANDN U49362 ( .A(n53233), .B(n32411), .Z(n32412) );
  AND U49363 ( .A(n53234), .B(n32412), .Z(n32415) );
  NANDN U49364 ( .A(n32415), .B(n53235), .Z(n32416) );
  AND U49365 ( .A(n32417), .B(n32416), .Z(n32418) );
  NAND U49366 ( .A(n52325), .B(n32418), .Z(n32420) );
  ANDN U49367 ( .B(n32420), .A(n32419), .Z(n32421) );
  NANDN U49368 ( .A(n32422), .B(n32421), .Z(n32426) );
  AND U49369 ( .A(n32424), .B(n32423), .Z(n32425) );
  NAND U49370 ( .A(n32426), .B(n32425), .Z(n32427) );
  NANDN U49371 ( .A(n32428), .B(n32427), .Z(n32430) );
  OR U49372 ( .A(n32430), .B(n32429), .Z(n32431) );
  NAND U49373 ( .A(n32432), .B(n32431), .Z(n32436) );
  AND U49374 ( .A(n32434), .B(n32433), .Z(n32435) );
  NAND U49375 ( .A(n32436), .B(n32435), .Z(n32437) );
  NANDN U49376 ( .A(n52322), .B(n32437), .Z(n32439) );
  ANDN U49377 ( .B(y[1196]), .A(x[1196]), .Z(n32438) );
  OR U49378 ( .A(n32439), .B(n32438), .Z(n32440) );
  NAND U49379 ( .A(n32441), .B(n32440), .Z(n32442) );
  NANDN U49380 ( .A(n52320), .B(n32442), .Z(n32444) );
  OR U49381 ( .A(n32444), .B(n32443), .Z(n32445) );
  NAND U49382 ( .A(n32446), .B(n32445), .Z(n32447) );
  NANDN U49383 ( .A(n53246), .B(n32447), .Z(n32448) );
  OR U49384 ( .A(n32449), .B(n32448), .Z(n32450) );
  AND U49385 ( .A(n32451), .B(n32450), .Z(n32453) );
  NAND U49386 ( .A(n32453), .B(n32452), .Z(n32454) );
  ANDN U49387 ( .B(y[1202]), .A(x[1202]), .Z(n53245) );
  ANDN U49388 ( .B(n32454), .A(n53245), .Z(n32455) );
  NANDN U49389 ( .A(n32456), .B(n32455), .Z(n32460) );
  AND U49390 ( .A(n32458), .B(n32457), .Z(n32459) );
  NAND U49391 ( .A(n32460), .B(n32459), .Z(n32461) );
  NANDN U49392 ( .A(n32462), .B(n32461), .Z(n32464) );
  OR U49393 ( .A(n32464), .B(n32463), .Z(n32465) );
  NAND U49394 ( .A(n32466), .B(n32465), .Z(n32470) );
  AND U49395 ( .A(n32468), .B(n32467), .Z(n32469) );
  NAND U49396 ( .A(n32470), .B(n32469), .Z(n32471) );
  NANDN U49397 ( .A(n32472), .B(n32471), .Z(n32473) );
  OR U49398 ( .A(n32474), .B(n32473), .Z(n32475) );
  AND U49399 ( .A(n32476), .B(n32475), .Z(n32478) );
  NANDN U49400 ( .A(x[1208]), .B(y[1208]), .Z(n32477) );
  NAND U49401 ( .A(n32478), .B(n32477), .Z(n32480) );
  ANDN U49402 ( .B(n32480), .A(n32479), .Z(n32481) );
  NANDN U49403 ( .A(n32482), .B(n32481), .Z(n32486) );
  NANDN U49404 ( .A(x[1210]), .B(y[1210]), .Z(n32483) );
  AND U49405 ( .A(n32484), .B(n32483), .Z(n32485) );
  NAND U49406 ( .A(n32486), .B(n32485), .Z(n32487) );
  NANDN U49407 ( .A(n32488), .B(n32487), .Z(n32490) );
  IV U49408 ( .A(n32489), .Z(n53257) );
  OR U49409 ( .A(n32490), .B(n53257), .Z(n32491) );
  AND U49410 ( .A(n32492), .B(n32491), .Z(n32493) );
  NAND U49411 ( .A(n53258), .B(n32493), .Z(n32494) );
  NANDN U49412 ( .A(n53259), .B(n32494), .Z(n32495) );
  AND U49413 ( .A(n53260), .B(n32495), .Z(n32496) );
  OR U49414 ( .A(n53261), .B(n32496), .Z(n32497) );
  NAND U49415 ( .A(n53262), .B(n32497), .Z(n32498) );
  NANDN U49416 ( .A(n32499), .B(n32498), .Z(n32500) );
  OR U49417 ( .A(n53263), .B(n32500), .Z(n32501) );
  AND U49418 ( .A(n32502), .B(n32501), .Z(n32503) );
  NAND U49419 ( .A(n32503), .B(n53264), .Z(n32505) );
  ANDN U49420 ( .B(n32505), .A(n32504), .Z(n32506) );
  NANDN U49421 ( .A(n32507), .B(n32506), .Z(n32511) );
  AND U49422 ( .A(n32509), .B(n32508), .Z(n32510) );
  NAND U49423 ( .A(n32511), .B(n32510), .Z(n32512) );
  NANDN U49424 ( .A(n32513), .B(n32512), .Z(n32514) );
  OR U49425 ( .A(n32515), .B(n32514), .Z(n32516) );
  AND U49426 ( .A(n32517), .B(n32516), .Z(n32518) );
  NANDN U49427 ( .A(n53270), .B(n32518), .Z(n32519) );
  NAND U49428 ( .A(n32520), .B(n32519), .Z(n32521) );
  NANDN U49429 ( .A(n52317), .B(n32521), .Z(n32524) );
  AND U49430 ( .A(n32522), .B(n52316), .Z(n32523) );
  NAND U49431 ( .A(n32524), .B(n32523), .Z(n32525) );
  NANDN U49432 ( .A(n53274), .B(n32525), .Z(n32526) );
  OR U49433 ( .A(n32527), .B(n32526), .Z(n32528) );
  AND U49434 ( .A(n32529), .B(n32528), .Z(n32530) );
  NANDN U49435 ( .A(n32531), .B(n32530), .Z(n32532) );
  AND U49436 ( .A(n32533), .B(n32532), .Z(n32534) );
  ANDN U49437 ( .B(n32535), .A(n32534), .Z(n32536) );
  NAND U49438 ( .A(n32537), .B(n32536), .Z(n32538) );
  NANDN U49439 ( .A(n32539), .B(n32538), .Z(n32541) );
  OR U49440 ( .A(n32541), .B(n32540), .Z(n32542) );
  NAND U49441 ( .A(n32543), .B(n32542), .Z(n32544) );
  NANDN U49442 ( .A(n32545), .B(n32544), .Z(n32549) );
  AND U49443 ( .A(n32547), .B(n32546), .Z(n32548) );
  NAND U49444 ( .A(n32549), .B(n32548), .Z(n32550) );
  NANDN U49445 ( .A(n32551), .B(n32550), .Z(n32552) );
  OR U49446 ( .A(n32553), .B(n32552), .Z(n32554) );
  AND U49447 ( .A(n32555), .B(n32554), .Z(n32557) );
  NAND U49448 ( .A(n32557), .B(n32556), .Z(n32559) );
  ANDN U49449 ( .B(n32559), .A(n32558), .Z(n32560) );
  NANDN U49450 ( .A(n32561), .B(n32560), .Z(n32565) );
  IV U49451 ( .A(n32562), .Z(n53286) );
  AND U49452 ( .A(n32563), .B(n53286), .Z(n32564) );
  NAND U49453 ( .A(n32565), .B(n32564), .Z(n32566) );
  NANDN U49454 ( .A(n32567), .B(n32566), .Z(n32569) );
  IV U49455 ( .A(n32568), .Z(n53287) );
  OR U49456 ( .A(n32569), .B(n53287), .Z(n32570) );
  AND U49457 ( .A(n53288), .B(n32570), .Z(n32573) );
  NAND U49458 ( .A(n32572), .B(n32571), .Z(n53289) );
  OR U49459 ( .A(n32573), .B(n53289), .Z(n32574) );
  AND U49460 ( .A(n53290), .B(n32574), .Z(n32575) );
  OR U49461 ( .A(n32576), .B(n32575), .Z(n32577) );
  NAND U49462 ( .A(n53292), .B(n32577), .Z(n32578) );
  NANDN U49463 ( .A(n32579), .B(n32578), .Z(n32583) );
  NAND U49464 ( .A(n32581), .B(n32580), .Z(n32582) );
  NANDN U49465 ( .A(n32583), .B(n32582), .Z(n32584) );
  AND U49466 ( .A(n53294), .B(n32584), .Z(n32585) );
  OR U49467 ( .A(n32586), .B(n32585), .Z(n32587) );
  AND U49468 ( .A(n32588), .B(n32587), .Z(n32589) );
  NOR U49469 ( .A(n32589), .B(n53297), .Z(n32590) );
  NANDN U49470 ( .A(n32591), .B(n32590), .Z(n32592) );
  AND U49471 ( .A(n53298), .B(n32592), .Z(n32594) );
  NAND U49472 ( .A(n32594), .B(n32593), .Z(n32595) );
  NANDN U49473 ( .A(n53299), .B(n32595), .Z(n32596) );
  AND U49474 ( .A(n32597), .B(n32596), .Z(n32598) );
  NAND U49475 ( .A(n32598), .B(n53300), .Z(n32600) );
  ANDN U49476 ( .B(n32600), .A(n32599), .Z(n32601) );
  NANDN U49477 ( .A(n53301), .B(n32601), .Z(n32605) );
  AND U49478 ( .A(n32603), .B(n32602), .Z(n32604) );
  NAND U49479 ( .A(n32605), .B(n32604), .Z(n32606) );
  NANDN U49480 ( .A(n32607), .B(n32606), .Z(n32609) );
  OR U49481 ( .A(n32609), .B(n32608), .Z(n32610) );
  NAND U49482 ( .A(n32611), .B(n32610), .Z(n32615) );
  AND U49483 ( .A(n32613), .B(n32612), .Z(n32614) );
  NAND U49484 ( .A(n32615), .B(n32614), .Z(n32616) );
  NANDN U49485 ( .A(n32617), .B(n32616), .Z(n32619) );
  OR U49486 ( .A(n32619), .B(n32618), .Z(n32620) );
  NAND U49487 ( .A(n32621), .B(n32620), .Z(n32622) );
  NANDN U49488 ( .A(n32623), .B(n32622), .Z(n32627) );
  AND U49489 ( .A(n32625), .B(n32624), .Z(n32626) );
  NAND U49490 ( .A(n32627), .B(n32626), .Z(n32628) );
  NANDN U49491 ( .A(n32629), .B(n32628), .Z(n32630) );
  OR U49492 ( .A(n32631), .B(n32630), .Z(n32632) );
  AND U49493 ( .A(n32633), .B(n32632), .Z(n32634) );
  NANDN U49494 ( .A(n32635), .B(n32634), .Z(n32636) );
  AND U49495 ( .A(n32637), .B(n32636), .Z(n32638) );
  NOR U49496 ( .A(n53314), .B(n32638), .Z(n32639) );
  NANDN U49497 ( .A(n32640), .B(n32639), .Z(n32641) );
  AND U49498 ( .A(n53315), .B(n32641), .Z(n32642) );
  OR U49499 ( .A(n53316), .B(n32642), .Z(n32643) );
  NAND U49500 ( .A(n53317), .B(n32643), .Z(n32644) );
  NANDN U49501 ( .A(n53318), .B(n32644), .Z(n32647) );
  AND U49502 ( .A(n32645), .B(n53320), .Z(n32646) );
  NAND U49503 ( .A(n32647), .B(n32646), .Z(n32648) );
  NANDN U49504 ( .A(n53321), .B(n32648), .Z(n32649) );
  OR U49505 ( .A(n32650), .B(n32649), .Z(n32651) );
  AND U49506 ( .A(n32652), .B(n32651), .Z(n32654) );
  NAND U49507 ( .A(n32654), .B(n32653), .Z(n32656) );
  AND U49508 ( .A(n32656), .B(n32655), .Z(n32657) );
  NAND U49509 ( .A(n32658), .B(n32657), .Z(n32659) );
  NAND U49510 ( .A(n32660), .B(n32659), .Z(n32661) );
  AND U49511 ( .A(n32662), .B(n32661), .Z(n32663) );
  OR U49512 ( .A(n32663), .B(n53325), .Z(n32664) );
  NAND U49513 ( .A(n53326), .B(n32664), .Z(n32665) );
  NANDN U49514 ( .A(n53327), .B(n32665), .Z(n32666) );
  NAND U49515 ( .A(n53328), .B(n32666), .Z(n32667) );
  ANDN U49516 ( .B(n32667), .A(n53329), .Z(n32668) );
  NANDN U49517 ( .A(n32669), .B(n32668), .Z(n32672) );
  AND U49518 ( .A(n32670), .B(n53330), .Z(n32671) );
  NAND U49519 ( .A(n32672), .B(n32671), .Z(n32673) );
  NANDN U49520 ( .A(n32674), .B(n32673), .Z(n32676) );
  OR U49521 ( .A(n32676), .B(n32675), .Z(n32677) );
  NAND U49522 ( .A(n32678), .B(n32677), .Z(n32682) );
  AND U49523 ( .A(n32680), .B(n32679), .Z(n32681) );
  NAND U49524 ( .A(n32682), .B(n32681), .Z(n32683) );
  NANDN U49525 ( .A(n32684), .B(n32683), .Z(n32686) );
  OR U49526 ( .A(n32686), .B(n32685), .Z(n32687) );
  NAND U49527 ( .A(n32688), .B(n32687), .Z(n32689) );
  NANDN U49528 ( .A(n32690), .B(n32689), .Z(n32694) );
  AND U49529 ( .A(n32692), .B(n32691), .Z(n32693) );
  NAND U49530 ( .A(n32694), .B(n32693), .Z(n32695) );
  NANDN U49531 ( .A(n32696), .B(n32695), .Z(n32698) );
  OR U49532 ( .A(n32698), .B(n32697), .Z(n32699) );
  NAND U49533 ( .A(n32700), .B(n32699), .Z(n32701) );
  NANDN U49534 ( .A(n32702), .B(n32701), .Z(n32706) );
  AND U49535 ( .A(n32704), .B(n32703), .Z(n32705) );
  NAND U49536 ( .A(n32706), .B(n32705), .Z(n32707) );
  NANDN U49537 ( .A(n32708), .B(n32707), .Z(n32709) );
  OR U49538 ( .A(n32710), .B(n32709), .Z(n32711) );
  AND U49539 ( .A(n32712), .B(n32711), .Z(n32713) );
  NANDN U49540 ( .A(n32714), .B(n32713), .Z(n32715) );
  AND U49541 ( .A(n32716), .B(n32715), .Z(n32717) );
  NOR U49542 ( .A(n32717), .B(n53347), .Z(n32718) );
  NANDN U49543 ( .A(n32719), .B(n32718), .Z(n32720) );
  AND U49544 ( .A(n32720), .B(n53348), .Z(n32722) );
  NAND U49545 ( .A(n32722), .B(n32721), .Z(n32723) );
  NANDN U49546 ( .A(n52309), .B(n32723), .Z(n32724) );
  AND U49547 ( .A(n32725), .B(n32724), .Z(n32726) );
  NAND U49548 ( .A(n52308), .B(n32726), .Z(n32728) );
  ANDN U49549 ( .B(n32728), .A(n32727), .Z(n32729) );
  NANDN U49550 ( .A(n53350), .B(n32729), .Z(n32733) );
  AND U49551 ( .A(n32731), .B(n32730), .Z(n32732) );
  NAND U49552 ( .A(n32733), .B(n32732), .Z(n32734) );
  NANDN U49553 ( .A(n32735), .B(n32734), .Z(n32736) );
  OR U49554 ( .A(n32737), .B(n32736), .Z(n32738) );
  AND U49555 ( .A(n32739), .B(n32738), .Z(n32740) );
  NANDN U49556 ( .A(n32741), .B(n32740), .Z(n32742) );
  AND U49557 ( .A(n32743), .B(n32742), .Z(n32745) );
  NAND U49558 ( .A(n32745), .B(n32744), .Z(n32747) );
  ANDN U49559 ( .B(n32747), .A(n32746), .Z(n32748) );
  NANDN U49560 ( .A(n32749), .B(n32748), .Z(n32752) );
  AND U49561 ( .A(n32750), .B(n53356), .Z(n32751) );
  NAND U49562 ( .A(n32752), .B(n32751), .Z(n32753) );
  NAND U49563 ( .A(n53357), .B(n32753), .Z(n32754) );
  NAND U49564 ( .A(n32755), .B(n32754), .Z(n32756) );
  NAND U49565 ( .A(n32757), .B(n32756), .Z(n32758) );
  NANDN U49566 ( .A(n32759), .B(n32758), .Z(n32760) );
  NANDN U49567 ( .A(n32760), .B(n52304), .Z(n32761) );
  NAND U49568 ( .A(n53360), .B(n32761), .Z(n32762) );
  AND U49569 ( .A(n32763), .B(n32762), .Z(n32764) );
  OR U49570 ( .A(n32764), .B(n53364), .Z(n32765) );
  AND U49571 ( .A(n32766), .B(n32765), .Z(n32767) );
  OR U49572 ( .A(n32768), .B(n32767), .Z(n32769) );
  AND U49573 ( .A(n32770), .B(n32769), .Z(n32772) );
  NAND U49574 ( .A(n32772), .B(n32771), .Z(n32774) );
  ANDN U49575 ( .B(n32774), .A(n32773), .Z(n32775) );
  NANDN U49576 ( .A(n32776), .B(n32775), .Z(n32780) );
  AND U49577 ( .A(n32778), .B(n32777), .Z(n32779) );
  NAND U49578 ( .A(n32780), .B(n32779), .Z(n32781) );
  NANDN U49579 ( .A(n32782), .B(n32781), .Z(n32784) );
  OR U49580 ( .A(n32784), .B(n32783), .Z(n32785) );
  AND U49581 ( .A(n32786), .B(n32785), .Z(n32790) );
  NAND U49582 ( .A(n32788), .B(n32787), .Z(n32789) );
  OR U49583 ( .A(n32790), .B(n32789), .Z(n32791) );
  AND U49584 ( .A(n32792), .B(n32791), .Z(n32794) );
  NAND U49585 ( .A(n32794), .B(n32793), .Z(n32796) );
  ANDN U49586 ( .B(n32796), .A(n32795), .Z(n32797) );
  NANDN U49587 ( .A(n32798), .B(n32797), .Z(n32802) );
  AND U49588 ( .A(n32800), .B(n32799), .Z(n32801) );
  NAND U49589 ( .A(n32802), .B(n32801), .Z(n32803) );
  NANDN U49590 ( .A(n32804), .B(n32803), .Z(n32806) );
  OR U49591 ( .A(n32806), .B(n32805), .Z(n32807) );
  NAND U49592 ( .A(n32808), .B(n32807), .Z(n32812) );
  AND U49593 ( .A(n32810), .B(n32809), .Z(n32811) );
  NAND U49594 ( .A(n32812), .B(n32811), .Z(n32813) );
  NANDN U49595 ( .A(n32814), .B(n32813), .Z(n32816) );
  OR U49596 ( .A(n32816), .B(n32815), .Z(n32817) );
  NAND U49597 ( .A(n32818), .B(n32817), .Z(n32819) );
  NANDN U49598 ( .A(n32820), .B(n32819), .Z(n32822) );
  OR U49599 ( .A(n32822), .B(n32821), .Z(n32823) );
  AND U49600 ( .A(n32824), .B(n32823), .Z(n32825) );
  OR U49601 ( .A(n32826), .B(n32825), .Z(n32827) );
  NAND U49602 ( .A(n32828), .B(n32827), .Z(n32829) );
  NANDN U49603 ( .A(n32830), .B(n32829), .Z(n32834) );
  AND U49604 ( .A(n32832), .B(n32831), .Z(n32833) );
  NAND U49605 ( .A(n32834), .B(n32833), .Z(n32835) );
  NANDN U49606 ( .A(n32836), .B(n32835), .Z(n32838) );
  OR U49607 ( .A(n32838), .B(n32837), .Z(n32839) );
  NAND U49608 ( .A(n32840), .B(n32839), .Z(n32841) );
  NANDN U49609 ( .A(n32842), .B(n32841), .Z(n32843) );
  OR U49610 ( .A(n32843), .B(n53408), .Z(n32844) );
  AND U49611 ( .A(n32845), .B(n32844), .Z(n32848) );
  NAND U49612 ( .A(n32847), .B(n32846), .Z(n53411) );
  OR U49613 ( .A(n32848), .B(n53411), .Z(n32849) );
  NAND U49614 ( .A(n32850), .B(n32849), .Z(n32851) );
  NANDN U49615 ( .A(n32852), .B(n32851), .Z(n32853) );
  OR U49616 ( .A(n32853), .B(n53410), .Z(n32854) );
  NAND U49617 ( .A(n32855), .B(n32854), .Z(n32859) );
  AND U49618 ( .A(n32857), .B(n32856), .Z(n32858) );
  NAND U49619 ( .A(n32859), .B(n32858), .Z(n32860) );
  NANDN U49620 ( .A(n32861), .B(n32860), .Z(n32863) );
  ANDN U49621 ( .B(y[1342]), .A(x[1342]), .Z(n32862) );
  OR U49622 ( .A(n32863), .B(n32862), .Z(n32864) );
  NAND U49623 ( .A(n32865), .B(n32864), .Z(n32866) );
  NANDN U49624 ( .A(n32867), .B(n32866), .Z(n32868) );
  OR U49625 ( .A(n32869), .B(n32868), .Z(n32870) );
  AND U49626 ( .A(n32871), .B(n32870), .Z(n32873) );
  NAND U49627 ( .A(n32873), .B(n32872), .Z(n32875) );
  ANDN U49628 ( .B(n32875), .A(n32874), .Z(n32876) );
  NANDN U49629 ( .A(n32877), .B(n32876), .Z(n32881) );
  AND U49630 ( .A(n32879), .B(n32878), .Z(n32880) );
  NAND U49631 ( .A(n32881), .B(n32880), .Z(n32882) );
  NANDN U49632 ( .A(n53423), .B(n32882), .Z(n32884) );
  OR U49633 ( .A(n32884), .B(n32883), .Z(n32885) );
  NAND U49634 ( .A(n32886), .B(n32885), .Z(n32887) );
  NANDN U49635 ( .A(n32888), .B(n32887), .Z(n32891) );
  AND U49636 ( .A(n32889), .B(n52300), .Z(n32890) );
  NAND U49637 ( .A(n32891), .B(n32890), .Z(n32892) );
  NANDN U49638 ( .A(n32893), .B(n32892), .Z(n32894) );
  OR U49639 ( .A(n32894), .B(n53425), .Z(n32895) );
  NAND U49640 ( .A(n32896), .B(n32895), .Z(n32897) );
  NANDN U49641 ( .A(n32898), .B(n32897), .Z(n32900) );
  OR U49642 ( .A(n32900), .B(n32899), .Z(n32901) );
  AND U49643 ( .A(n32902), .B(n32901), .Z(n32906) );
  NAND U49644 ( .A(n32904), .B(n32903), .Z(n32905) );
  OR U49645 ( .A(n32906), .B(n32905), .Z(n32907) );
  AND U49646 ( .A(n32908), .B(n32907), .Z(n32912) );
  NAND U49647 ( .A(n32910), .B(n32909), .Z(n32911) );
  OR U49648 ( .A(n32912), .B(n32911), .Z(n32913) );
  AND U49649 ( .A(n32914), .B(n32913), .Z(n32918) );
  NAND U49650 ( .A(n32916), .B(n32915), .Z(n32917) );
  OR U49651 ( .A(n32918), .B(n32917), .Z(n32919) );
  AND U49652 ( .A(n32920), .B(n32919), .Z(n32921) );
  ANDN U49653 ( .B(n32922), .A(n32921), .Z(n32923) );
  NAND U49654 ( .A(n32924), .B(n32923), .Z(n32925) );
  NANDN U49655 ( .A(n32926), .B(n32925), .Z(n32928) );
  OR U49656 ( .A(n32928), .B(n32927), .Z(n32929) );
  NAND U49657 ( .A(n32930), .B(n32929), .Z(n32931) );
  NANDN U49658 ( .A(n32932), .B(n32931), .Z(n32933) );
  OR U49659 ( .A(n32934), .B(n32933), .Z(n32935) );
  AND U49660 ( .A(n32936), .B(n32935), .Z(n32937) );
  NANDN U49661 ( .A(n32938), .B(n32937), .Z(n32939) );
  AND U49662 ( .A(n32940), .B(n32939), .Z(n32941) );
  OR U49663 ( .A(n32942), .B(n32941), .Z(n32943) );
  NAND U49664 ( .A(n32944), .B(n32943), .Z(n32948) );
  AND U49665 ( .A(n32946), .B(n32945), .Z(n32947) );
  NAND U49666 ( .A(n32948), .B(n32947), .Z(n32949) );
  NANDN U49667 ( .A(n32950), .B(n32949), .Z(n32952) );
  OR U49668 ( .A(n32952), .B(n32951), .Z(n32953) );
  NAND U49669 ( .A(n32954), .B(n32953), .Z(n32955) );
  NANDN U49670 ( .A(n32956), .B(n32955), .Z(n32957) );
  OR U49671 ( .A(n32958), .B(n32957), .Z(n32959) );
  AND U49672 ( .A(n32960), .B(n32959), .Z(n32962) );
  NAND U49673 ( .A(n32962), .B(n32961), .Z(n32964) );
  ANDN U49674 ( .B(n32964), .A(n32963), .Z(n32965) );
  NANDN U49675 ( .A(n32966), .B(n32965), .Z(n32970) );
  AND U49676 ( .A(n32968), .B(n32967), .Z(n32969) );
  NAND U49677 ( .A(n32970), .B(n32969), .Z(n32971) );
  NANDN U49678 ( .A(n32972), .B(n32971), .Z(n32974) );
  IV U49679 ( .A(n32973), .Z(n53444) );
  OR U49680 ( .A(n32974), .B(n53444), .Z(n32975) );
  AND U49681 ( .A(n32975), .B(n53445), .Z(n32977) );
  NAND U49682 ( .A(n32977), .B(n32976), .Z(n32978) );
  AND U49683 ( .A(n53446), .B(n32978), .Z(n32979) );
  OR U49684 ( .A(n32979), .B(n53447), .Z(n32980) );
  NAND U49685 ( .A(n53448), .B(n32980), .Z(n32981) );
  NANDN U49686 ( .A(n53449), .B(n32981), .Z(n32982) );
  AND U49687 ( .A(n32982), .B(n53452), .Z(n32983) );
  OR U49688 ( .A(n32983), .B(n52285), .Z(n32984) );
  NAND U49689 ( .A(n52284), .B(n32984), .Z(n32985) );
  NAND U49690 ( .A(n53453), .B(n32985), .Z(n32986) );
  NAND U49691 ( .A(n53454), .B(n32986), .Z(n32987) );
  NAND U49692 ( .A(n53455), .B(n32987), .Z(n32988) );
  AND U49693 ( .A(n32989), .B(n32988), .Z(n32992) );
  NAND U49694 ( .A(n53457), .B(n32990), .Z(n32991) );
  OR U49695 ( .A(n32992), .B(n32991), .Z(n32993) );
  AND U49696 ( .A(n32994), .B(n32993), .Z(n32998) );
  NAND U49697 ( .A(n32996), .B(n32995), .Z(n32997) );
  OR U49698 ( .A(n32998), .B(n32997), .Z(n32999) );
  AND U49699 ( .A(n33000), .B(n32999), .Z(n33002) );
  AND U49700 ( .A(n33002), .B(n33001), .Z(n33003) );
  OR U49701 ( .A(n33004), .B(n33003), .Z(n33005) );
  NAND U49702 ( .A(n33006), .B(n33005), .Z(n33010) );
  IV U49703 ( .A(n33007), .Z(n53465) );
  AND U49704 ( .A(n33008), .B(n53465), .Z(n33009) );
  NAND U49705 ( .A(n33010), .B(n33009), .Z(n33011) );
  NANDN U49706 ( .A(n33012), .B(n33011), .Z(n33014) );
  IV U49707 ( .A(n33013), .Z(n53466) );
  OR U49708 ( .A(n33014), .B(n53466), .Z(n33015) );
  AND U49709 ( .A(n53467), .B(n33015), .Z(n33016) );
  OR U49710 ( .A(n53468), .B(n33016), .Z(n33017) );
  NAND U49711 ( .A(n53469), .B(n33017), .Z(n33018) );
  NANDN U49712 ( .A(n33019), .B(n33018), .Z(n33021) );
  IV U49713 ( .A(n33020), .Z(n53470) );
  OR U49714 ( .A(n33021), .B(n53470), .Z(n33022) );
  AND U49715 ( .A(n33023), .B(n33022), .Z(n33024) );
  NANDN U49716 ( .A(n53471), .B(n33024), .Z(n33025) );
  NAND U49717 ( .A(n33026), .B(n33025), .Z(n33030) );
  NAND U49718 ( .A(n33028), .B(n33027), .Z(n33029) );
  ANDN U49719 ( .B(n33030), .A(n33029), .Z(n33034) );
  NAND U49720 ( .A(n33032), .B(n33031), .Z(n33033) );
  OR U49721 ( .A(n33034), .B(n33033), .Z(n33035) );
  AND U49722 ( .A(n33036), .B(n33035), .Z(n33042) );
  OR U49723 ( .A(n33038), .B(n33037), .Z(n33039) );
  AND U49724 ( .A(n33040), .B(n33039), .Z(n33041) );
  OR U49725 ( .A(n33042), .B(n33041), .Z(n33043) );
  AND U49726 ( .A(n53478), .B(n33043), .Z(n33044) );
  ANDN U49727 ( .B(n33045), .A(n33044), .Z(n33046) );
  OR U49728 ( .A(n33047), .B(n33046), .Z(n33048) );
  NAND U49729 ( .A(n33049), .B(n33048), .Z(n33050) );
  NANDN U49730 ( .A(n33051), .B(n33050), .Z(n33052) );
  OR U49731 ( .A(n33053), .B(n33052), .Z(n33054) );
  AND U49732 ( .A(n33055), .B(n33054), .Z(n33056) );
  NANDN U49733 ( .A(n53485), .B(n33056), .Z(n33057) );
  AND U49734 ( .A(n33058), .B(n33057), .Z(n33059) );
  OR U49735 ( .A(n53487), .B(n33059), .Z(n33060) );
  NAND U49736 ( .A(n33061), .B(n33060), .Z(n33062) );
  NANDN U49737 ( .A(n33063), .B(n33062), .Z(n33065) );
  IV U49738 ( .A(n33064), .Z(n53489) );
  OR U49739 ( .A(n33065), .B(n53489), .Z(n33066) );
  NAND U49740 ( .A(n33067), .B(n33066), .Z(n33070) );
  AND U49741 ( .A(n33068), .B(n53493), .Z(n33069) );
  NAND U49742 ( .A(n33070), .B(n33069), .Z(n33071) );
  NANDN U49743 ( .A(n33072), .B(n33071), .Z(n33073) );
  OR U49744 ( .A(n33073), .B(n52280), .Z(n33074) );
  AND U49745 ( .A(n53494), .B(n33074), .Z(n33076) );
  NANDN U49746 ( .A(n33076), .B(n53495), .Z(n33077) );
  NAND U49747 ( .A(n52279), .B(n33077), .Z(n33078) );
  NAND U49748 ( .A(n53497), .B(n33078), .Z(n33081) );
  AND U49749 ( .A(n33079), .B(n53498), .Z(n33080) );
  NAND U49750 ( .A(n33081), .B(n33080), .Z(n33082) );
  NANDN U49751 ( .A(n33083), .B(n33082), .Z(n33084) );
  OR U49752 ( .A(n33084), .B(n52278), .Z(n33085) );
  AND U49753 ( .A(n53501), .B(n33085), .Z(n33086) );
  NANDN U49754 ( .A(n33087), .B(n33086), .Z(n33091) );
  NANDN U49755 ( .A(n33089), .B(n33088), .Z(n33090) );
  AND U49756 ( .A(n33091), .B(n33090), .Z(n33092) );
  AND U49757 ( .A(n33092), .B(n53502), .Z(n33093) );
  OR U49758 ( .A(n53503), .B(n33093), .Z(n33094) );
  NAND U49759 ( .A(n53504), .B(n33094), .Z(n33095) );
  NAND U49760 ( .A(n53505), .B(n33095), .Z(n33096) );
  AND U49761 ( .A(n53506), .B(n33096), .Z(n33099) );
  NANDN U49762 ( .A(n33099), .B(n53507), .Z(n33100) );
  AND U49763 ( .A(n33101), .B(n33100), .Z(n33102) );
  NAND U49764 ( .A(n53508), .B(n33102), .Z(n33104) );
  ANDN U49765 ( .B(n33104), .A(n33103), .Z(n33105) );
  NANDN U49766 ( .A(n52277), .B(n33105), .Z(n33109) );
  AND U49767 ( .A(n33107), .B(n33106), .Z(n33108) );
  NAND U49768 ( .A(n33109), .B(n33108), .Z(n33110) );
  NANDN U49769 ( .A(n33111), .B(n33110), .Z(n33112) );
  OR U49770 ( .A(n53512), .B(n33112), .Z(n33113) );
  AND U49771 ( .A(n33114), .B(n33113), .Z(n33115) );
  NANDN U49772 ( .A(n53513), .B(n33115), .Z(n33116) );
  AND U49773 ( .A(n53514), .B(n33116), .Z(n33119) );
  NAND U49774 ( .A(n33118), .B(n33117), .Z(n52275) );
  OR U49775 ( .A(n33119), .B(n52275), .Z(n33120) );
  NAND U49776 ( .A(n33121), .B(n33120), .Z(n33122) );
  NANDN U49777 ( .A(n53516), .B(n33122), .Z(n33123) );
  AND U49778 ( .A(n33124), .B(n33123), .Z(n33126) );
  IV U49779 ( .A(n33125), .Z(n53517) );
  OR U49780 ( .A(n33126), .B(n53517), .Z(n33127) );
  NAND U49781 ( .A(n33128), .B(n33127), .Z(n33129) );
  NANDN U49782 ( .A(n33130), .B(n33129), .Z(n33134) );
  AND U49783 ( .A(n33132), .B(n33131), .Z(n33133) );
  NAND U49784 ( .A(n33134), .B(n33133), .Z(n33135) );
  NANDN U49785 ( .A(n33136), .B(n33135), .Z(n33137) );
  OR U49786 ( .A(n33138), .B(n33137), .Z(n33139) );
  AND U49787 ( .A(n33140), .B(n33139), .Z(n33142) );
  NAND U49788 ( .A(n33142), .B(n33141), .Z(n33144) );
  ANDN U49789 ( .B(n33144), .A(n33143), .Z(n33145) );
  NANDN U49790 ( .A(n33146), .B(n33145), .Z(n33147) );
  AND U49791 ( .A(n33148), .B(n33147), .Z(n33149) );
  OR U49792 ( .A(n33150), .B(n33149), .Z(n33151) );
  NAND U49793 ( .A(n33152), .B(n33151), .Z(n33153) );
  NANDN U49794 ( .A(n33154), .B(n33153), .Z(n33158) );
  AND U49795 ( .A(n33156), .B(n33155), .Z(n33157) );
  NAND U49796 ( .A(n33158), .B(n33157), .Z(n33159) );
  NANDN U49797 ( .A(n33160), .B(n33159), .Z(n33162) );
  ANDN U49798 ( .B(y[1456]), .A(x[1456]), .Z(n33161) );
  OR U49799 ( .A(n33162), .B(n33161), .Z(n33163) );
  NAND U49800 ( .A(n33164), .B(n33163), .Z(n33165) );
  NANDN U49801 ( .A(n33166), .B(n33165), .Z(n33167) );
  OR U49802 ( .A(n33168), .B(n33167), .Z(n33169) );
  AND U49803 ( .A(n33170), .B(n33169), .Z(n33172) );
  NAND U49804 ( .A(n33172), .B(n33171), .Z(n33174) );
  ANDN U49805 ( .B(n33174), .A(n33173), .Z(n33175) );
  NANDN U49806 ( .A(n33176), .B(n33175), .Z(n33180) );
  IV U49807 ( .A(n33177), .Z(n53529) );
  AND U49808 ( .A(n33178), .B(n53529), .Z(n33179) );
  NAND U49809 ( .A(n33180), .B(n33179), .Z(n33181) );
  NANDN U49810 ( .A(n53531), .B(n33181), .Z(n33183) );
  OR U49811 ( .A(n33183), .B(n33182), .Z(n33184) );
  NAND U49812 ( .A(n53532), .B(n33184), .Z(n33185) );
  NANDN U49813 ( .A(n33186), .B(n33185), .Z(n33189) );
  AND U49814 ( .A(n33187), .B(n53534), .Z(n33188) );
  NAND U49815 ( .A(n33189), .B(n33188), .Z(n33190) );
  NANDN U49816 ( .A(n33191), .B(n33190), .Z(n33192) );
  OR U49817 ( .A(n33193), .B(n33192), .Z(n33194) );
  AND U49818 ( .A(n33195), .B(n33194), .Z(n33196) );
  NANDN U49819 ( .A(n53537), .B(n33196), .Z(n33197) );
  AND U49820 ( .A(n33198), .B(n33197), .Z(n33199) );
  OR U49821 ( .A(n53539), .B(n33199), .Z(n33200) );
  NAND U49822 ( .A(n53540), .B(n33200), .Z(n33201) );
  NANDN U49823 ( .A(n33202), .B(n33201), .Z(n33203) );
  OR U49824 ( .A(n53541), .B(n33203), .Z(n33204) );
  AND U49825 ( .A(n33205), .B(n33204), .Z(n33206) );
  NAND U49826 ( .A(n33206), .B(n53542), .Z(n33208) );
  ANDN U49827 ( .B(n33208), .A(n33207), .Z(n33209) );
  NANDN U49828 ( .A(n33210), .B(n33209), .Z(n33214) );
  AND U49829 ( .A(n33212), .B(n33211), .Z(n33213) );
  NAND U49830 ( .A(n33214), .B(n33213), .Z(n33215) );
  NANDN U49831 ( .A(n33216), .B(n33215), .Z(n33217) );
  OR U49832 ( .A(n33218), .B(n33217), .Z(n33219) );
  AND U49833 ( .A(n33220), .B(n33219), .Z(n33221) );
  NANDN U49834 ( .A(n33222), .B(n33221), .Z(n33223) );
  AND U49835 ( .A(n53550), .B(n33223), .Z(n33225) );
  NAND U49836 ( .A(n33225), .B(n33224), .Z(n33226) );
  NAND U49837 ( .A(n33227), .B(n33226), .Z(n33228) );
  OR U49838 ( .A(n53551), .B(n33228), .Z(n33229) );
  AND U49839 ( .A(n33229), .B(n53552), .Z(n33232) );
  AND U49840 ( .A(n33231), .B(n33230), .Z(n53553) );
  NANDN U49841 ( .A(n33232), .B(n53553), .Z(n33233) );
  NAND U49842 ( .A(n33234), .B(n33233), .Z(n33235) );
  NANDN U49843 ( .A(n33236), .B(n33235), .Z(n33237) );
  OR U49844 ( .A(n33237), .B(n52265), .Z(n33238) );
  NAND U49845 ( .A(n33239), .B(n33238), .Z(n33243) );
  AND U49846 ( .A(n33241), .B(n33240), .Z(n33242) );
  NAND U49847 ( .A(n33243), .B(n33242), .Z(n33244) );
  NANDN U49848 ( .A(n33245), .B(n33244), .Z(n33247) );
  OR U49849 ( .A(n33247), .B(n33246), .Z(n33248) );
  NAND U49850 ( .A(n33249), .B(n33248), .Z(n33250) );
  NANDN U49851 ( .A(n33251), .B(n33250), .Z(n33253) );
  OR U49852 ( .A(n33253), .B(n33252), .Z(n33254) );
  AND U49853 ( .A(n33255), .B(n33254), .Z(n33259) );
  NAND U49854 ( .A(n33257), .B(n33256), .Z(n33258) );
  OR U49855 ( .A(n33259), .B(n33258), .Z(n33260) );
  AND U49856 ( .A(n33261), .B(n33260), .Z(n33265) );
  NAND U49857 ( .A(n33263), .B(n33262), .Z(n33264) );
  OR U49858 ( .A(n33265), .B(n33264), .Z(n33266) );
  AND U49859 ( .A(n33267), .B(n33266), .Z(n33271) );
  NAND U49860 ( .A(n33269), .B(n33268), .Z(n33270) );
  OR U49861 ( .A(n33271), .B(n33270), .Z(n33272) );
  AND U49862 ( .A(n33273), .B(n33272), .Z(n33274) );
  NOR U49863 ( .A(n52262), .B(n33274), .Z(n33275) );
  NANDN U49864 ( .A(n33276), .B(n33275), .Z(n33277) );
  AND U49865 ( .A(n53567), .B(n33277), .Z(n33278) );
  NANDN U49866 ( .A(n33279), .B(n33278), .Z(n33280) );
  NAND U49867 ( .A(n53568), .B(n33280), .Z(n33281) );
  NANDN U49868 ( .A(n33282), .B(n33281), .Z(n33285) );
  AND U49869 ( .A(n33283), .B(n53570), .Z(n33284) );
  NAND U49870 ( .A(n33285), .B(n33284), .Z(n33286) );
  NANDN U49871 ( .A(n33287), .B(n33286), .Z(n33288) );
  OR U49872 ( .A(n33289), .B(n33288), .Z(n33290) );
  AND U49873 ( .A(n33291), .B(n33290), .Z(n33292) );
  NANDN U49874 ( .A(n53574), .B(n33292), .Z(n33293) );
  AND U49875 ( .A(n33294), .B(n33293), .Z(n33295) );
  OR U49876 ( .A(n53576), .B(n33295), .Z(n33296) );
  NAND U49877 ( .A(n33297), .B(n33296), .Z(n33298) );
  NANDN U49878 ( .A(n33299), .B(n33298), .Z(n33301) );
  IV U49879 ( .A(n33300), .Z(n53579) );
  OR U49880 ( .A(n33301), .B(n53579), .Z(n33302) );
  AND U49881 ( .A(n33303), .B(n33302), .Z(n33304) );
  OR U49882 ( .A(n33305), .B(n33304), .Z(n33306) );
  NAND U49883 ( .A(n33307), .B(n33306), .Z(n33311) );
  AND U49884 ( .A(n33309), .B(n33308), .Z(n33310) );
  NAND U49885 ( .A(n33311), .B(n33310), .Z(n33312) );
  NANDN U49886 ( .A(n53584), .B(n33312), .Z(n33313) );
  OR U49887 ( .A(n33314), .B(n33313), .Z(n33315) );
  AND U49888 ( .A(n33316), .B(n33315), .Z(n33317) );
  NANDN U49889 ( .A(n53585), .B(n33317), .Z(n33318) );
  AND U49890 ( .A(n53586), .B(n33318), .Z(n33321) );
  NAND U49891 ( .A(n33320), .B(n33319), .Z(n52259) );
  OR U49892 ( .A(n33321), .B(n52259), .Z(n33322) );
  NAND U49893 ( .A(n53587), .B(n33322), .Z(n33323) );
  NANDN U49894 ( .A(n53588), .B(n33323), .Z(n33326) );
  AND U49895 ( .A(n33324), .B(n53589), .Z(n33325) );
  NAND U49896 ( .A(n33326), .B(n33325), .Z(n33327) );
  NANDN U49897 ( .A(n33328), .B(n33327), .Z(n33329) );
  OR U49898 ( .A(n33329), .B(n53590), .Z(n33330) );
  NAND U49899 ( .A(n33331), .B(n33330), .Z(n33334) );
  AND U49900 ( .A(n33332), .B(n53595), .Z(n33333) );
  NAND U49901 ( .A(n33334), .B(n33333), .Z(n33335) );
  NANDN U49902 ( .A(n33336), .B(n33335), .Z(n33337) );
  OR U49903 ( .A(n33337), .B(n52258), .Z(n33340) );
  AND U49904 ( .A(n33339), .B(n33338), .Z(n52257) );
  AND U49905 ( .A(n33340), .B(n52257), .Z(n33341) );
  OR U49906 ( .A(n53596), .B(n33341), .Z(n33342) );
  NAND U49907 ( .A(n53597), .B(n33342), .Z(n33343) );
  NANDN U49908 ( .A(n33344), .B(n33343), .Z(n33345) );
  OR U49909 ( .A(n53598), .B(n33345), .Z(n33346) );
  AND U49910 ( .A(n33347), .B(n33346), .Z(n33348) );
  NANDN U49911 ( .A(n53599), .B(n33348), .Z(n33349) );
  NAND U49912 ( .A(n33350), .B(n33349), .Z(n33351) );
  NANDN U49913 ( .A(n33352), .B(n33351), .Z(n33354) );
  OR U49914 ( .A(n33354), .B(n33353), .Z(n33355) );
  NAND U49915 ( .A(n33356), .B(n33355), .Z(n33357) );
  NANDN U49916 ( .A(n33358), .B(n33357), .Z(n33361) );
  NANDN U49917 ( .A(y[1532]), .B(n33361), .Z(n33360) );
  ANDN U49918 ( .B(n33360), .A(n33359), .Z(n33364) );
  XNOR U49919 ( .A(n33361), .B(y[1532]), .Z(n33362) );
  NAND U49920 ( .A(n33362), .B(x[1532]), .Z(n33363) );
  NAND U49921 ( .A(n33364), .B(n33363), .Z(n33365) );
  NAND U49922 ( .A(n53607), .B(n33365), .Z(n33366) );
  NANDN U49923 ( .A(n53608), .B(n33366), .Z(n33367) );
  AND U49924 ( .A(n33368), .B(n33367), .Z(n33369) );
  OR U49925 ( .A(n33370), .B(n33369), .Z(n33371) );
  AND U49926 ( .A(n33372), .B(n33371), .Z(n33373) );
  OR U49927 ( .A(n33374), .B(n33373), .Z(n33375) );
  NAND U49928 ( .A(n33376), .B(n33375), .Z(n33377) );
  NANDN U49929 ( .A(n33378), .B(n33377), .Z(n33379) );
  AND U49930 ( .A(n33380), .B(n33379), .Z(n33381) );
  NAND U49931 ( .A(n33382), .B(n33381), .Z(n33386) );
  NAND U49932 ( .A(n33384), .B(n33383), .Z(n33385) );
  ANDN U49933 ( .B(n33386), .A(n33385), .Z(n33387) );
  OR U49934 ( .A(n33388), .B(n33387), .Z(n33389) );
  NAND U49935 ( .A(n33390), .B(n33389), .Z(n33394) );
  AND U49936 ( .A(n33392), .B(n33391), .Z(n33393) );
  NAND U49937 ( .A(n33394), .B(n33393), .Z(n33395) );
  NANDN U49938 ( .A(n52255), .B(n33395), .Z(n33396) );
  OR U49939 ( .A(n33397), .B(n33396), .Z(n33398) );
  AND U49940 ( .A(n33399), .B(n33398), .Z(n33400) );
  NANDN U49941 ( .A(n33401), .B(n33400), .Z(n33402) );
  AND U49942 ( .A(n33403), .B(n33402), .Z(n33404) );
  OR U49943 ( .A(n33405), .B(n33404), .Z(n33406) );
  NAND U49944 ( .A(n33407), .B(n33406), .Z(n33408) );
  NANDN U49945 ( .A(n33409), .B(n33408), .Z(n33412) );
  AND U49946 ( .A(n33410), .B(n53626), .Z(n33411) );
  NAND U49947 ( .A(n33412), .B(n33411), .Z(n33413) );
  NANDN U49948 ( .A(n33414), .B(n33413), .Z(n33415) );
  OR U49949 ( .A(n33415), .B(n52253), .Z(n33418) );
  AND U49950 ( .A(n33417), .B(n33416), .Z(n52252) );
  AND U49951 ( .A(n33418), .B(n52252), .Z(n33421) );
  NANDN U49952 ( .A(n33421), .B(n53627), .Z(n33422) );
  NAND U49953 ( .A(n53628), .B(n33422), .Z(n33423) );
  NAND U49954 ( .A(n53629), .B(n33423), .Z(n33424) );
  NAND U49955 ( .A(n33425), .B(n33424), .Z(n33426) );
  AND U49956 ( .A(n33427), .B(n33426), .Z(n33428) );
  ANDN U49957 ( .B(n33429), .A(n33428), .Z(n33430) );
  NAND U49958 ( .A(n52250), .B(n33430), .Z(n33431) );
  NANDN U49959 ( .A(n53633), .B(n33431), .Z(n33433) );
  OR U49960 ( .A(n33433), .B(n33432), .Z(n33434) );
  NAND U49961 ( .A(n33435), .B(n33434), .Z(n33436) );
  NANDN U49962 ( .A(n33437), .B(n33436), .Z(n33439) );
  OR U49963 ( .A(n33439), .B(n33438), .Z(n33440) );
  NAND U49964 ( .A(n33441), .B(n33440), .Z(n33442) );
  AND U49965 ( .A(n53645), .B(n33442), .Z(n33443) );
  NAND U49966 ( .A(n33444), .B(n33443), .Z(n33445) );
  NANDN U49967 ( .A(n53647), .B(n33445), .Z(n33447) );
  OR U49968 ( .A(n33447), .B(n33446), .Z(n33448) );
  NAND U49969 ( .A(n53649), .B(n33448), .Z(n33449) );
  NANDN U49970 ( .A(n33450), .B(n33449), .Z(n33453) );
  AND U49971 ( .A(n33451), .B(n53653), .Z(n33452) );
  NAND U49972 ( .A(n33453), .B(n33452), .Z(n33454) );
  NANDN U49973 ( .A(n33455), .B(n33454), .Z(n33457) );
  OR U49974 ( .A(n33457), .B(n33456), .Z(n33458) );
  NAND U49975 ( .A(n33459), .B(n33458), .Z(n33460) );
  NANDN U49976 ( .A(n33461), .B(n33460), .Z(n33463) );
  OR U49977 ( .A(n33463), .B(n33462), .Z(n33464) );
  AND U49978 ( .A(n33465), .B(n33464), .Z(n33466) );
  OR U49979 ( .A(n33467), .B(n33466), .Z(n33468) );
  NAND U49980 ( .A(n33469), .B(n33468), .Z(n33470) );
  NANDN U49981 ( .A(n33471), .B(n33470), .Z(n33472) );
  AND U49982 ( .A(n33473), .B(n33472), .Z(n33474) );
  NAND U49983 ( .A(n33475), .B(n33474), .Z(n33476) );
  NANDN U49984 ( .A(n33477), .B(n33476), .Z(n33479) );
  OR U49985 ( .A(n33479), .B(n33478), .Z(n33480) );
  NAND U49986 ( .A(n33481), .B(n33480), .Z(n33482) );
  NANDN U49987 ( .A(n33483), .B(n33482), .Z(n33485) );
  OR U49988 ( .A(n33485), .B(n33484), .Z(n33486) );
  NAND U49989 ( .A(n33487), .B(n33486), .Z(n33491) );
  AND U49990 ( .A(n33489), .B(n33488), .Z(n33490) );
  NAND U49991 ( .A(n33491), .B(n33490), .Z(n33492) );
  NANDN U49992 ( .A(n33493), .B(n33492), .Z(n33496) );
  AND U49993 ( .A(n33494), .B(n53681), .Z(n33495) );
  NAND U49994 ( .A(n33496), .B(n33495), .Z(n33497) );
  NANDN U49995 ( .A(n33498), .B(n33497), .Z(n33499) );
  OR U49996 ( .A(n33500), .B(n33499), .Z(n33501) );
  AND U49997 ( .A(n33502), .B(n33501), .Z(n33503) );
  NANDN U49998 ( .A(n33504), .B(n33503), .Z(n33505) );
  NAND U49999 ( .A(n33506), .B(n33505), .Z(n33507) );
  NANDN U50000 ( .A(n52247), .B(n33507), .Z(n33508) );
  AND U50001 ( .A(n33509), .B(n33508), .Z(n33511) );
  OR U50002 ( .A(n33511), .B(n33510), .Z(n33512) );
  AND U50003 ( .A(n33512), .B(n53691), .Z(n33514) );
  IV U50004 ( .A(n33513), .Z(n53693) );
  NANDN U50005 ( .A(n33514), .B(n53693), .Z(n33515) );
  NANDN U50006 ( .A(n53694), .B(n33515), .Z(n33516) );
  AND U50007 ( .A(n33517), .B(n33516), .Z(n33518) );
  OR U50008 ( .A(n33519), .B(n33518), .Z(n33520) );
  NAND U50009 ( .A(n33521), .B(n33520), .Z(n33522) );
  NANDN U50010 ( .A(n33523), .B(n33522), .Z(n33524) );
  OR U50011 ( .A(n33524), .B(n53698), .Z(n33525) );
  AND U50012 ( .A(n33526), .B(n33525), .Z(n33529) );
  NAND U50013 ( .A(n33528), .B(n33527), .Z(n52246) );
  OR U50014 ( .A(n33529), .B(n52246), .Z(n33530) );
  NAND U50015 ( .A(n53700), .B(n33530), .Z(n33531) );
  NAND U50016 ( .A(n53701), .B(n33531), .Z(n33532) );
  NAND U50017 ( .A(n53702), .B(n33532), .Z(n33533) );
  ANDN U50018 ( .B(n33533), .A(n53703), .Z(n33534) );
  NANDN U50019 ( .A(n33535), .B(n33534), .Z(n33538) );
  AND U50020 ( .A(n33536), .B(n53704), .Z(n33537) );
  NAND U50021 ( .A(n33538), .B(n33537), .Z(n33539) );
  NANDN U50022 ( .A(n33540), .B(n33539), .Z(n33541) );
  OR U50023 ( .A(n33542), .B(n33541), .Z(n33543) );
  AND U50024 ( .A(n33544), .B(n33543), .Z(n33545) );
  NAND U50025 ( .A(n33545), .B(n53708), .Z(n33547) );
  ANDN U50026 ( .B(n33547), .A(n33546), .Z(n33548) );
  NANDN U50027 ( .A(n53710), .B(n33548), .Z(n33549) );
  AND U50028 ( .A(n53711), .B(n33549), .Z(n33552) );
  NANDN U50029 ( .A(x[1608]), .B(y[1608]), .Z(n33551) );
  NAND U50030 ( .A(n33551), .B(n33550), .Z(n53712) );
  OR U50031 ( .A(n33552), .B(n53712), .Z(n33553) );
  AND U50032 ( .A(n33554), .B(n33553), .Z(n33555) );
  NAND U50033 ( .A(n33555), .B(n53713), .Z(n33557) );
  ANDN U50034 ( .B(n33557), .A(n33556), .Z(n33558) );
  NANDN U50035 ( .A(n53714), .B(n33558), .Z(n33562) );
  AND U50036 ( .A(n33560), .B(n33559), .Z(n33561) );
  NAND U50037 ( .A(n33562), .B(n33561), .Z(n33563) );
  NANDN U50038 ( .A(n33564), .B(n33563), .Z(n33566) );
  OR U50039 ( .A(n33566), .B(n33565), .Z(n33567) );
  NAND U50040 ( .A(n33568), .B(n33567), .Z(n33569) );
  NANDN U50041 ( .A(n33570), .B(n33569), .Z(n33571) );
  OR U50042 ( .A(n33572), .B(n33571), .Z(n33573) );
  AND U50043 ( .A(n33574), .B(n33573), .Z(n33576) );
  NAND U50044 ( .A(n33576), .B(n33575), .Z(n33578) );
  ANDN U50045 ( .B(n33578), .A(n33577), .Z(n33579) );
  NANDN U50046 ( .A(n33580), .B(n33579), .Z(n33584) );
  AND U50047 ( .A(n33582), .B(n33581), .Z(n33583) );
  NAND U50048 ( .A(n33584), .B(n33583), .Z(n33585) );
  NANDN U50049 ( .A(n33586), .B(n33585), .Z(n33588) );
  OR U50050 ( .A(n33588), .B(n33587), .Z(n33589) );
  NAND U50051 ( .A(n33590), .B(n33589), .Z(n33591) );
  NANDN U50052 ( .A(n33592), .B(n33591), .Z(n33593) );
  OR U50053 ( .A(n33594), .B(n33593), .Z(n33595) );
  AND U50054 ( .A(n33596), .B(n33595), .Z(n33598) );
  NAND U50055 ( .A(n33598), .B(n33597), .Z(n33600) );
  ANDN U50056 ( .B(n33600), .A(n33599), .Z(n33601) );
  NANDN U50057 ( .A(n33602), .B(n33601), .Z(n33606) );
  AND U50058 ( .A(n33604), .B(n33603), .Z(n33605) );
  NAND U50059 ( .A(n33606), .B(n33605), .Z(n33607) );
  NANDN U50060 ( .A(n33608), .B(n33607), .Z(n33610) );
  OR U50061 ( .A(n33610), .B(n33609), .Z(n33611) );
  NAND U50062 ( .A(n33612), .B(n33611), .Z(n33613) );
  NANDN U50063 ( .A(n33614), .B(n33613), .Z(n33615) );
  OR U50064 ( .A(n33616), .B(n33615), .Z(n33617) );
  AND U50065 ( .A(n33618), .B(n33617), .Z(n33620) );
  NAND U50066 ( .A(n33620), .B(n33619), .Z(n33622) );
  ANDN U50067 ( .B(y[1628]), .A(x[1628]), .Z(n33621) );
  ANDN U50068 ( .B(n33622), .A(n33621), .Z(n33623) );
  NANDN U50069 ( .A(n33624), .B(n33623), .Z(n33627) );
  AND U50070 ( .A(n33625), .B(n53736), .Z(n33626) );
  NAND U50071 ( .A(n33627), .B(n33626), .Z(n33628) );
  NANDN U50072 ( .A(n33629), .B(n33628), .Z(n33631) );
  OR U50073 ( .A(n33631), .B(n33630), .Z(n33632) );
  NAND U50074 ( .A(n53740), .B(n33632), .Z(n33633) );
  NANDN U50075 ( .A(n33634), .B(n33633), .Z(n33637) );
  AND U50076 ( .A(n33635), .B(n53738), .Z(n33636) );
  NAND U50077 ( .A(n33637), .B(n33636), .Z(n33638) );
  NANDN U50078 ( .A(n33639), .B(n33638), .Z(n33640) );
  OR U50079 ( .A(n33641), .B(n33640), .Z(n33642) );
  AND U50080 ( .A(n33643), .B(n33642), .Z(n33644) );
  NANDN U50081 ( .A(n52244), .B(n33644), .Z(n33645) );
  AND U50082 ( .A(n33646), .B(n33645), .Z(n33649) );
  NANDN U50083 ( .A(n33649), .B(n53743), .Z(n33650) );
  NAND U50084 ( .A(n53745), .B(n33650), .Z(n33651) );
  NAND U50085 ( .A(n53746), .B(n33651), .Z(n33652) );
  NAND U50086 ( .A(n52242), .B(n33652), .Z(n33653) );
  AND U50087 ( .A(n33654), .B(n33653), .Z(n33655) );
  OR U50088 ( .A(n33656), .B(n33655), .Z(n33657) );
  NAND U50089 ( .A(n33658), .B(n33657), .Z(n33659) );
  NAND U50090 ( .A(n33660), .B(n33659), .Z(n33662) );
  AND U50091 ( .A(n33662), .B(n33661), .Z(n33663) );
  NAND U50092 ( .A(n33664), .B(n33663), .Z(n33665) );
  NAND U50093 ( .A(n33666), .B(n33665), .Z(n33667) );
  AND U50094 ( .A(n33668), .B(n33667), .Z(n33669) );
  OR U50095 ( .A(n33669), .B(n53750), .Z(n33670) );
  AND U50096 ( .A(n33671), .B(n33670), .Z(n33672) );
  NANDN U50097 ( .A(n53752), .B(n33672), .Z(n33673) );
  AND U50098 ( .A(n33674), .B(n33673), .Z(n33678) );
  NAND U50099 ( .A(n33676), .B(n33675), .Z(n33677) );
  OR U50100 ( .A(n33678), .B(n33677), .Z(n33679) );
  AND U50101 ( .A(n33680), .B(n33679), .Z(n33681) );
  OR U50102 ( .A(n33682), .B(n33681), .Z(n33683) );
  NAND U50103 ( .A(n33684), .B(n33683), .Z(n33685) );
  NANDN U50104 ( .A(n33686), .B(n33685), .Z(n33687) );
  AND U50105 ( .A(n33688), .B(n33687), .Z(n33689) );
  OR U50106 ( .A(n33690), .B(n33689), .Z(n33691) );
  NAND U50107 ( .A(n33692), .B(n33691), .Z(n33696) );
  AND U50108 ( .A(n33694), .B(n33693), .Z(n33695) );
  NAND U50109 ( .A(n33696), .B(n33695), .Z(n33697) );
  NANDN U50110 ( .A(n52236), .B(n33697), .Z(n33699) );
  OR U50111 ( .A(n33699), .B(n33698), .Z(n33700) );
  NAND U50112 ( .A(n33701), .B(n33700), .Z(n33702) );
  NANDN U50113 ( .A(n33703), .B(n33702), .Z(n33706) );
  AND U50114 ( .A(n33704), .B(n53779), .Z(n33705) );
  NAND U50115 ( .A(n33706), .B(n33705), .Z(n33707) );
  NANDN U50116 ( .A(n33708), .B(n33707), .Z(n33709) );
  OR U50117 ( .A(n33709), .B(n53783), .Z(n33710) );
  NAND U50118 ( .A(n33711), .B(n33710), .Z(n33712) );
  NANDN U50119 ( .A(n33713), .B(n33712), .Z(n33715) );
  OR U50120 ( .A(n33715), .B(n33714), .Z(n33716) );
  AND U50121 ( .A(n33717), .B(n33716), .Z(n33721) );
  NAND U50122 ( .A(n33719), .B(n33718), .Z(n33720) );
  OR U50123 ( .A(n33721), .B(n33720), .Z(n33722) );
  AND U50124 ( .A(n33723), .B(n33722), .Z(n33724) );
  NOR U50125 ( .A(n33725), .B(n33724), .Z(n33726) );
  NANDN U50126 ( .A(n33727), .B(n33726), .Z(n33728) );
  AND U50127 ( .A(n33729), .B(n33728), .Z(n33730) );
  OR U50128 ( .A(n53798), .B(n33730), .Z(n33731) );
  AND U50129 ( .A(n53799), .B(n33731), .Z(n33734) );
  NAND U50130 ( .A(n33733), .B(n33732), .Z(n52235) );
  OR U50131 ( .A(n33734), .B(n52235), .Z(n33735) );
  NAND U50132 ( .A(n33736), .B(n33735), .Z(n33737) );
  NANDN U50133 ( .A(n33738), .B(n33737), .Z(n33739) );
  OR U50134 ( .A(n53801), .B(n33739), .Z(n33740) );
  AND U50135 ( .A(n33741), .B(n33740), .Z(n33743) );
  NAND U50136 ( .A(n33743), .B(n33742), .Z(n33745) );
  ANDN U50137 ( .B(n33745), .A(n33744), .Z(n33746) );
  NANDN U50138 ( .A(n33747), .B(n33746), .Z(n33748) );
  NAND U50139 ( .A(n33749), .B(n33748), .Z(n33751) );
  ANDN U50140 ( .B(y[1680]), .A(x[1680]), .Z(n33750) );
  ANDN U50141 ( .B(n33751), .A(n33750), .Z(n33753) );
  ANDN U50142 ( .B(n33753), .A(n33752), .Z(n33757) );
  NAND U50143 ( .A(n33755), .B(n33754), .Z(n33756) );
  OR U50144 ( .A(n33757), .B(n33756), .Z(n33758) );
  AND U50145 ( .A(n33759), .B(n33758), .Z(n33760) );
  NOR U50146 ( .A(n33760), .B(n53811), .Z(n33761) );
  NANDN U50147 ( .A(n33762), .B(n33761), .Z(n33763) );
  AND U50148 ( .A(n33764), .B(n33763), .Z(n33765) );
  NAND U50149 ( .A(n53812), .B(n33765), .Z(n33766) );
  NANDN U50150 ( .A(n53813), .B(n33766), .Z(n33767) );
  AND U50151 ( .A(n33768), .B(n33767), .Z(n33770) );
  AND U50152 ( .A(n33769), .B(n52232), .Z(n53815) );
  NANDN U50153 ( .A(n33770), .B(n53815), .Z(n33771) );
  NAND U50154 ( .A(n33772), .B(n33771), .Z(n33773) );
  NAND U50155 ( .A(n53816), .B(n33773), .Z(n33774) );
  NAND U50156 ( .A(n53817), .B(n33774), .Z(n33775) );
  NANDN U50157 ( .A(n53818), .B(n33775), .Z(n33776) );
  AND U50158 ( .A(n33777), .B(n33776), .Z(n33780) );
  NAND U50159 ( .A(n53820), .B(n33778), .Z(n33779) );
  OR U50160 ( .A(n33780), .B(n33779), .Z(n33781) );
  AND U50161 ( .A(n33782), .B(n33781), .Z(n33786) );
  NAND U50162 ( .A(n33784), .B(n33783), .Z(n33785) );
  OR U50163 ( .A(n33786), .B(n33785), .Z(n33787) );
  AND U50164 ( .A(n33788), .B(n33787), .Z(n33792) );
  NAND U50165 ( .A(n33790), .B(n33789), .Z(n33791) );
  OR U50166 ( .A(n33792), .B(n33791), .Z(n33793) );
  AND U50167 ( .A(n33794), .B(n33793), .Z(n33798) );
  NAND U50168 ( .A(n33796), .B(n33795), .Z(n33797) );
  OR U50169 ( .A(n33798), .B(n33797), .Z(n33799) );
  AND U50170 ( .A(n33800), .B(n33799), .Z(n33804) );
  NAND U50171 ( .A(n33802), .B(n33801), .Z(n33803) );
  OR U50172 ( .A(n33804), .B(n33803), .Z(n33805) );
  AND U50173 ( .A(n33806), .B(n33805), .Z(n33810) );
  NAND U50174 ( .A(n33808), .B(n33807), .Z(n33809) );
  OR U50175 ( .A(n33810), .B(n33809), .Z(n33811) );
  AND U50176 ( .A(n33812), .B(n33811), .Z(n33813) );
  NOR U50177 ( .A(n33814), .B(n33813), .Z(n33815) );
  NAND U50178 ( .A(n33816), .B(n33815), .Z(n33817) );
  NANDN U50179 ( .A(n33818), .B(n33817), .Z(n33822) );
  AND U50180 ( .A(n33820), .B(n33819), .Z(n33821) );
  NAND U50181 ( .A(n33822), .B(n33821), .Z(n33823) );
  NANDN U50182 ( .A(n33824), .B(n33823), .Z(n33825) );
  OR U50183 ( .A(n33826), .B(n33825), .Z(n33827) );
  AND U50184 ( .A(n33828), .B(n33827), .Z(n33829) );
  NANDN U50185 ( .A(n33830), .B(n33829), .Z(n33831) );
  AND U50186 ( .A(n33832), .B(n33831), .Z(n33836) );
  NAND U50187 ( .A(n33834), .B(n33833), .Z(n33835) );
  OR U50188 ( .A(n33836), .B(n33835), .Z(n33837) );
  AND U50189 ( .A(n33838), .B(n33837), .Z(n33839) );
  ANDN U50190 ( .B(n33840), .A(n33839), .Z(n33841) );
  NAND U50191 ( .A(n53836), .B(n33841), .Z(n33842) );
  NANDN U50192 ( .A(n53837), .B(n33842), .Z(n33844) );
  OR U50193 ( .A(n33844), .B(n33843), .Z(n33845) );
  NAND U50194 ( .A(n53838), .B(n33845), .Z(n33846) );
  NANDN U50195 ( .A(n33847), .B(n33846), .Z(n33850) );
  AND U50196 ( .A(n33848), .B(n52220), .Z(n33849) );
  NAND U50197 ( .A(n33850), .B(n33849), .Z(n33851) );
  NANDN U50198 ( .A(n33852), .B(n33851), .Z(n33854) );
  ANDN U50199 ( .B(y[1718]), .A(x[1718]), .Z(n33853) );
  OR U50200 ( .A(n33854), .B(n33853), .Z(n33855) );
  NAND U50201 ( .A(n33856), .B(n33855), .Z(n33857) );
  NANDN U50202 ( .A(n53844), .B(n33857), .Z(n33859) );
  OR U50203 ( .A(n33859), .B(n33858), .Z(n33860) );
  NAND U50204 ( .A(n53845), .B(n33860), .Z(n33861) );
  NANDN U50205 ( .A(n53846), .B(n33861), .Z(n33864) );
  AND U50206 ( .A(n33862), .B(n53847), .Z(n33863) );
  NAND U50207 ( .A(n33864), .B(n33863), .Z(n33865) );
  NANDN U50208 ( .A(n53850), .B(n33865), .Z(n33866) );
  OR U50209 ( .A(n33866), .B(n53848), .Z(n33867) );
  NAND U50210 ( .A(n33868), .B(n33867), .Z(n33869) );
  AND U50211 ( .A(n33870), .B(n33869), .Z(n33871) );
  NAND U50212 ( .A(n53851), .B(n33871), .Z(n33872) );
  NANDN U50213 ( .A(n33873), .B(n33872), .Z(n33875) );
  OR U50214 ( .A(n33875), .B(n33874), .Z(n33876) );
  NAND U50215 ( .A(n33877), .B(n33876), .Z(n33878) );
  NANDN U50216 ( .A(n33879), .B(n33878), .Z(n33881) );
  OR U50217 ( .A(n33881), .B(n33880), .Z(n33882) );
  NAND U50218 ( .A(n33883), .B(n33882), .Z(n33884) );
  NAND U50219 ( .A(n33885), .B(n33884), .Z(n33886) );
  NANDN U50220 ( .A(n53860), .B(n33886), .Z(n33887) );
  AND U50221 ( .A(n53861), .B(n33887), .Z(n33890) );
  NAND U50222 ( .A(n33889), .B(n33888), .Z(n53862) );
  OR U50223 ( .A(n33890), .B(n53862), .Z(n33891) );
  NAND U50224 ( .A(n33892), .B(n33891), .Z(n33893) );
  NANDN U50225 ( .A(n52219), .B(n33893), .Z(n33895) );
  NAND U50226 ( .A(n33895), .B(n33894), .Z(n33896) );
  NANDN U50227 ( .A(n52217), .B(n33896), .Z(n33897) );
  AND U50228 ( .A(n33897), .B(n52216), .Z(n33898) );
  OR U50229 ( .A(n33898), .B(n53864), .Z(n33899) );
  AND U50230 ( .A(n33899), .B(n53865), .Z(n33900) );
  OR U50231 ( .A(n33900), .B(n52215), .Z(n33901) );
  AND U50232 ( .A(n33901), .B(n52214), .Z(n33902) );
  OR U50233 ( .A(n33903), .B(n33902), .Z(n33904) );
  NAND U50234 ( .A(n33905), .B(n33904), .Z(n33906) );
  NANDN U50235 ( .A(n53871), .B(n33906), .Z(n33907) );
  OR U50236 ( .A(n33908), .B(n33907), .Z(n33909) );
  AND U50237 ( .A(n53872), .B(n33909), .Z(n33911) );
  NAND U50238 ( .A(n33911), .B(n33910), .Z(n33912) );
  NAND U50239 ( .A(n33913), .B(n33912), .Z(n33915) );
  IV U50240 ( .A(n33914), .Z(n53874) );
  AND U50241 ( .A(n33915), .B(n53874), .Z(n33916) );
  OR U50242 ( .A(n33917), .B(n33916), .Z(n33918) );
  NAND U50243 ( .A(n33919), .B(n33918), .Z(n33920) );
  NAND U50244 ( .A(n33921), .B(n33920), .Z(n33922) );
  NAND U50245 ( .A(n33923), .B(n33922), .Z(n33924) );
  AND U50246 ( .A(n33924), .B(n53880), .Z(n33926) );
  NANDN U50247 ( .A(x[1756]), .B(y[1756]), .Z(n33925) );
  AND U50248 ( .A(n33926), .B(n33925), .Z(n33927) );
  OR U50249 ( .A(n53881), .B(n33927), .Z(n33928) );
  NAND U50250 ( .A(n33929), .B(n33928), .Z(n33930) );
  NANDN U50251 ( .A(n33931), .B(n33930), .Z(n33933) );
  IV U50252 ( .A(n33932), .Z(n53884) );
  OR U50253 ( .A(n33933), .B(n53884), .Z(n33934) );
  AND U50254 ( .A(n33935), .B(n33934), .Z(n33936) );
  OR U50255 ( .A(n33937), .B(n33936), .Z(n33938) );
  NAND U50256 ( .A(n33939), .B(n33938), .Z(n33940) );
  NANDN U50257 ( .A(n33941), .B(n33940), .Z(n33944) );
  AND U50258 ( .A(n52212), .B(n33942), .Z(n33943) );
  NAND U50259 ( .A(n33944), .B(n33943), .Z(n33945) );
  NANDN U50260 ( .A(n33946), .B(n33945), .Z(n33947) );
  OR U50261 ( .A(n53891), .B(n33947), .Z(n33948) );
  AND U50262 ( .A(n33949), .B(n33948), .Z(n33950) );
  OR U50263 ( .A(n33950), .B(n53893), .Z(n33953) );
  AND U50264 ( .A(n33952), .B(n33951), .Z(n52210) );
  AND U50265 ( .A(n33953), .B(n52210), .Z(n33956) );
  NANDN U50266 ( .A(n33956), .B(n53894), .Z(n33957) );
  NAND U50267 ( .A(n33958), .B(n33957), .Z(n33959) );
  NANDN U50268 ( .A(n33960), .B(n33959), .Z(n33961) );
  OR U50269 ( .A(n33961), .B(n52209), .Z(n33962) );
  AND U50270 ( .A(n33963), .B(n33962), .Z(n33964) );
  NANDN U50271 ( .A(n33965), .B(n33964), .Z(n33966) );
  ANDN U50272 ( .B(y[1782]), .A(x[1782]), .Z(n33974) );
  OR U50273 ( .A(n33975), .B(n33974), .Z(n33976) );
  AND U50274 ( .A(n33977), .B(n33976), .Z(n33978) );
  OR U50275 ( .A(n33979), .B(n33978), .Z(n33980) );
  NAND U50276 ( .A(n33981), .B(n33980), .Z(n33982) );
  NANDN U50277 ( .A(n33983), .B(n33982), .Z(n33984) );
  NAND U50278 ( .A(n53913), .B(n33984), .Z(n33985) );
  NANDN U50279 ( .A(n53916), .B(n33985), .Z(n33986) );
  AND U50280 ( .A(n33986), .B(n53918), .Z(n33987) );
  OR U50281 ( .A(n33987), .B(n52207), .Z(n33988) );
  AND U50282 ( .A(n33989), .B(n33988), .Z(n33990) );
  NAND U50283 ( .A(n33991), .B(n33990), .Z(n33992) );
  NAND U50284 ( .A(n53919), .B(n33992), .Z(n33993) );
  NANDN U50285 ( .A(n52205), .B(n33993), .Z(n33994) );
  NAND U50286 ( .A(n33995), .B(n33994), .Z(n33996) );
  NANDN U50287 ( .A(n33997), .B(n33996), .Z(n33998) );
  AND U50288 ( .A(n33999), .B(n33998), .Z(n34000) );
  OR U50289 ( .A(n34001), .B(n34000), .Z(n34002) );
  NAND U50290 ( .A(n34003), .B(n34002), .Z(n34004) );
  NANDN U50291 ( .A(n34005), .B(n34004), .Z(n34006) );
  AND U50292 ( .A(n34007), .B(n34006), .Z(n34009) );
  NANDN U50293 ( .A(n34009), .B(n34008), .Z(n34011) );
  IV U50294 ( .A(n34010), .Z(n53930) );
  AND U50295 ( .A(n34011), .B(n53930), .Z(n34012) );
  OR U50296 ( .A(n34013), .B(n34012), .Z(n34014) );
  NAND U50297 ( .A(n34015), .B(n34014), .Z(n34016) );
  NANDN U50298 ( .A(n34017), .B(n34016), .Z(n34019) );
  IV U50299 ( .A(n34018), .Z(n53933) );
  OR U50300 ( .A(n34019), .B(n53933), .Z(n34020) );
  AND U50301 ( .A(n34021), .B(n34020), .Z(n34022) );
  OR U50302 ( .A(n53935), .B(n34022), .Z(n34023) );
  NAND U50303 ( .A(n53936), .B(n34023), .Z(n34024) );
  NANDN U50304 ( .A(n53937), .B(n34024), .Z(n34025) );
  NAND U50305 ( .A(n53938), .B(n34025), .Z(n34026) );
  AND U50306 ( .A(n34027), .B(n34026), .Z(n34028) );
  OR U50307 ( .A(n34029), .B(n34028), .Z(n34030) );
  NAND U50308 ( .A(n34031), .B(n34030), .Z(n34032) );
  NANDN U50309 ( .A(n34033), .B(n34032), .Z(n34037) );
  AND U50310 ( .A(n34035), .B(n34034), .Z(n34036) );
  NAND U50311 ( .A(n34037), .B(n34036), .Z(n34038) );
  NANDN U50312 ( .A(n34039), .B(n34038), .Z(n34040) );
  OR U50313 ( .A(n34041), .B(n34040), .Z(n34042) );
  AND U50314 ( .A(n34043), .B(n34042), .Z(n34045) );
  NAND U50315 ( .A(n34045), .B(n34044), .Z(n34047) );
  ANDN U50316 ( .B(n34047), .A(n34046), .Z(n34048) );
  NANDN U50317 ( .A(n52200), .B(n34048), .Z(n34049) );
  AND U50318 ( .A(n34050), .B(n34049), .Z(n34053) );
  AND U50319 ( .A(n34052), .B(n34051), .Z(n53948) );
  NANDN U50320 ( .A(n34053), .B(n53948), .Z(n34054) );
  NANDN U50321 ( .A(n53949), .B(n34054), .Z(n34055) );
  AND U50322 ( .A(n53950), .B(n34055), .Z(n34056) );
  OR U50323 ( .A(n53951), .B(n34056), .Z(n34057) );
  NAND U50324 ( .A(n53952), .B(n34057), .Z(n34058) );
  NANDN U50325 ( .A(n34059), .B(n34058), .Z(n34062) );
  AND U50326 ( .A(n34060), .B(n53953), .Z(n34061) );
  NAND U50327 ( .A(n34062), .B(n34061), .Z(n34063) );
  NANDN U50328 ( .A(n34064), .B(n34063), .Z(n34066) );
  OR U50329 ( .A(n34066), .B(n34065), .Z(n34067) );
  NAND U50330 ( .A(n34068), .B(n34067), .Z(n34069) );
  NANDN U50331 ( .A(n34070), .B(n34069), .Z(n34071) );
  OR U50332 ( .A(n34072), .B(n34071), .Z(n34073) );
  AND U50333 ( .A(n34074), .B(n34073), .Z(n34076) );
  NAND U50334 ( .A(n34076), .B(n34075), .Z(n34078) );
  ANDN U50335 ( .B(n34078), .A(n34077), .Z(n34079) );
  NANDN U50336 ( .A(n34080), .B(n34079), .Z(n34081) );
  AND U50337 ( .A(n34082), .B(n34081), .Z(n34083) );
  NAND U50338 ( .A(n34084), .B(n34083), .Z(n34085) );
  NANDN U50339 ( .A(n34086), .B(n34085), .Z(n34087) );
  OR U50340 ( .A(n34088), .B(n34087), .Z(n34089) );
  AND U50341 ( .A(n34090), .B(n34089), .Z(n34091) );
  NANDN U50342 ( .A(n34092), .B(n34091), .Z(n34093) );
  AND U50343 ( .A(n34094), .B(n34093), .Z(n34095) );
  OR U50344 ( .A(n34096), .B(n34095), .Z(n34097) );
  NAND U50345 ( .A(n53967), .B(n34097), .Z(n34098) );
  NANDN U50346 ( .A(n34099), .B(n34098), .Z(n34100) );
  OR U50347 ( .A(n53968), .B(n34100), .Z(n34101) );
  AND U50348 ( .A(n34102), .B(n34101), .Z(n34103) );
  NAND U50349 ( .A(n53969), .B(n34103), .Z(n34105) );
  ANDN U50350 ( .B(n34105), .A(n34104), .Z(n34106) );
  NANDN U50351 ( .A(n34107), .B(n34106), .Z(n34111) );
  IV U50352 ( .A(n34108), .Z(n53973) );
  AND U50353 ( .A(n34109), .B(n53973), .Z(n34110) );
  NAND U50354 ( .A(n34111), .B(n34110), .Z(n34112) );
  NANDN U50355 ( .A(n34113), .B(n34112), .Z(n34114) );
  OR U50356 ( .A(n53974), .B(n34114), .Z(n34115) );
  AND U50357 ( .A(n53976), .B(n34115), .Z(n34116) );
  NOR U50358 ( .A(n53977), .B(n34116), .Z(n34117) );
  NAND U50359 ( .A(n34118), .B(n34117), .Z(n34119) );
  NANDN U50360 ( .A(n53978), .B(n34119), .Z(n34121) );
  OR U50361 ( .A(n34121), .B(n34120), .Z(n34122) );
  NAND U50362 ( .A(n34123), .B(n34122), .Z(n34124) );
  NANDN U50363 ( .A(n34125), .B(n34124), .Z(n34127) );
  OR U50364 ( .A(n34127), .B(n34126), .Z(n34128) );
  NAND U50365 ( .A(n34129), .B(n34128), .Z(n34133) );
  AND U50366 ( .A(n34131), .B(n34130), .Z(n34132) );
  NAND U50367 ( .A(n34133), .B(n34132), .Z(n34134) );
  NANDN U50368 ( .A(n53985), .B(n34134), .Z(n34135) );
  OR U50369 ( .A(n34136), .B(n34135), .Z(n34137) );
  AND U50370 ( .A(n34138), .B(n34137), .Z(n34139) );
  NANDN U50371 ( .A(n53986), .B(n34139), .Z(n34140) );
  AND U50372 ( .A(n53987), .B(n34140), .Z(n34143) );
  NANDN U50373 ( .A(y[1851]), .B(x[1851]), .Z(n34141) );
  NAND U50374 ( .A(n34142), .B(n34141), .Z(n52198) );
  OR U50375 ( .A(n34143), .B(n52198), .Z(n34145) );
  IV U50376 ( .A(n34144), .Z(n53988) );
  AND U50377 ( .A(n34145), .B(n53988), .Z(n34147) );
  IV U50378 ( .A(n34146), .Z(n53989) );
  OR U50379 ( .A(n34147), .B(n53989), .Z(n34148) );
  AND U50380 ( .A(n53990), .B(n34148), .Z(n34149) );
  OR U50381 ( .A(n34149), .B(n53991), .Z(n34150) );
  AND U50382 ( .A(n53992), .B(n34150), .Z(n34151) );
  OR U50383 ( .A(n53994), .B(n34151), .Z(n34152) );
  NAND U50384 ( .A(n53995), .B(n34152), .Z(n34153) );
  NANDN U50385 ( .A(n53996), .B(n34153), .Z(n34154) );
  NANDN U50386 ( .A(n52197), .B(n34154), .Z(n34155) );
  AND U50387 ( .A(n34156), .B(n34155), .Z(n34157) );
  NANDN U50388 ( .A(n53997), .B(n34157), .Z(n34158) );
  AND U50389 ( .A(n34159), .B(n34158), .Z(n34160) );
  OR U50390 ( .A(n34161), .B(n34160), .Z(n34162) );
  NAND U50391 ( .A(n34163), .B(n34162), .Z(n34164) );
  AND U50392 ( .A(n34165), .B(n34164), .Z(n34166) );
  OR U50393 ( .A(n34167), .B(n34166), .Z(n34168) );
  NAND U50394 ( .A(n34169), .B(n34168), .Z(n34170) );
  NANDN U50395 ( .A(n34171), .B(n34170), .Z(n34172) );
  AND U50396 ( .A(n34173), .B(n34172), .Z(n34174) );
  NAND U50397 ( .A(n34175), .B(n34174), .Z(n34179) );
  NAND U50398 ( .A(n34177), .B(n34176), .Z(n34178) );
  ANDN U50399 ( .B(n34179), .A(n34178), .Z(n34183) );
  NAND U50400 ( .A(n34181), .B(n34180), .Z(n34182) );
  OR U50401 ( .A(n34183), .B(n34182), .Z(n34184) );
  AND U50402 ( .A(n34185), .B(n34184), .Z(n34189) );
  NAND U50403 ( .A(n34187), .B(n34186), .Z(n34188) );
  OR U50404 ( .A(n34189), .B(n34188), .Z(n34190) );
  AND U50405 ( .A(n34191), .B(n34190), .Z(n34195) );
  NAND U50406 ( .A(n34193), .B(n34192), .Z(n34194) );
  OR U50407 ( .A(n34195), .B(n34194), .Z(n34196) );
  AND U50408 ( .A(n34197), .B(n34196), .Z(n34198) );
  ANDN U50409 ( .B(n34199), .A(n34198), .Z(n34200) );
  NAND U50410 ( .A(n34201), .B(n34200), .Z(n34202) );
  NANDN U50411 ( .A(n34203), .B(n34202), .Z(n34205) );
  OR U50412 ( .A(n34205), .B(n34204), .Z(n34206) );
  NAND U50413 ( .A(n34207), .B(n34206), .Z(n34208) );
  NANDN U50414 ( .A(n34209), .B(n34208), .Z(n34211) );
  OR U50415 ( .A(n34211), .B(n34210), .Z(n34212) );
  AND U50416 ( .A(n34213), .B(n34212), .Z(n34214) );
  OR U50417 ( .A(n34215), .B(n34214), .Z(n34216) );
  NAND U50418 ( .A(n54017), .B(n34216), .Z(n34217) );
  NANDN U50419 ( .A(n34218), .B(n34217), .Z(n34219) );
  OR U50420 ( .A(n34219), .B(n54018), .Z(n34220) );
  AND U50421 ( .A(n34221), .B(n34220), .Z(n34222) );
  OR U50422 ( .A(n34223), .B(n34222), .Z(n34224) );
  NAND U50423 ( .A(n34225), .B(n34224), .Z(n34226) );
  AND U50424 ( .A(n34226), .B(n54024), .Z(n34228) );
  NANDN U50425 ( .A(x[1888]), .B(y[1888]), .Z(n34227) );
  NAND U50426 ( .A(n34228), .B(n34227), .Z(n34229) );
  NANDN U50427 ( .A(n54025), .B(n34229), .Z(n34230) );
  AND U50428 ( .A(n54026), .B(n34230), .Z(n34231) );
  OR U50429 ( .A(n54027), .B(n34231), .Z(n34232) );
  NAND U50430 ( .A(n54028), .B(n34232), .Z(n34233) );
  NANDN U50431 ( .A(n34234), .B(n34233), .Z(n34237) );
  NANDN U50432 ( .A(x[1894]), .B(y[1894]), .Z(n54030) );
  AND U50433 ( .A(n34235), .B(n54030), .Z(n34236) );
  NAND U50434 ( .A(n34237), .B(n34236), .Z(n34238) );
  NANDN U50435 ( .A(n34239), .B(n34238), .Z(n34243) );
  AND U50436 ( .A(n34241), .B(n34240), .Z(n34242) );
  NAND U50437 ( .A(n34243), .B(n34242), .Z(n34244) );
  NANDN U50438 ( .A(n34245), .B(n34244), .Z(n34246) );
  OR U50439 ( .A(n34247), .B(n34246), .Z(n34248) );
  AND U50440 ( .A(n34249), .B(n34248), .Z(n34250) );
  NANDN U50441 ( .A(n34251), .B(n34250), .Z(n34252) );
  AND U50442 ( .A(n34253), .B(n34252), .Z(n34254) );
  OR U50443 ( .A(n34255), .B(n34254), .Z(n34256) );
  AND U50444 ( .A(n34257), .B(n34256), .Z(n34258) );
  OR U50445 ( .A(n34258), .B(n52188), .Z(n34259) );
  AND U50446 ( .A(n34259), .B(n52187), .Z(n34260) );
  OR U50447 ( .A(n34260), .B(n54037), .Z(n34261) );
  NAND U50448 ( .A(n54038), .B(n34261), .Z(n34262) );
  NANDN U50449 ( .A(n54039), .B(n34262), .Z(n34263) );
  AND U50450 ( .A(n34263), .B(n54040), .Z(n34264) );
  OR U50451 ( .A(n34264), .B(n52186), .Z(n34265) );
  NAND U50452 ( .A(n54041), .B(n34265), .Z(n34266) );
  NAND U50453 ( .A(n54042), .B(n34266), .Z(n34269) );
  AND U50454 ( .A(n34267), .B(n52185), .Z(n34268) );
  NAND U50455 ( .A(n34269), .B(n34268), .Z(n34270) );
  NANDN U50456 ( .A(n54043), .B(n34270), .Z(n34272) );
  OR U50457 ( .A(n34272), .B(n34271), .Z(n34273) );
  NAND U50458 ( .A(n34274), .B(n34273), .Z(n34275) );
  NANDN U50459 ( .A(n34276), .B(n34275), .Z(n34277) );
  OR U50460 ( .A(n34278), .B(n34277), .Z(n34279) );
  AND U50461 ( .A(n34280), .B(n34279), .Z(n34282) );
  NAND U50462 ( .A(n34282), .B(n34281), .Z(n34284) );
  ANDN U50463 ( .B(n34284), .A(n34283), .Z(n34285) );
  NANDN U50464 ( .A(n34286), .B(n34285), .Z(n34290) );
  AND U50465 ( .A(n34288), .B(n34287), .Z(n34289) );
  NAND U50466 ( .A(n34290), .B(n34289), .Z(n34291) );
  NANDN U50467 ( .A(n34292), .B(n34291), .Z(n34293) );
  OR U50468 ( .A(n34294), .B(n34293), .Z(n34295) );
  AND U50469 ( .A(n34296), .B(n34295), .Z(n34297) );
  NANDN U50470 ( .A(n54052), .B(n34297), .Z(n34298) );
  NAND U50471 ( .A(n34299), .B(n34298), .Z(n34300) );
  NANDN U50472 ( .A(n34301), .B(n34300), .Z(n34306) );
  NANDN U50473 ( .A(n34303), .B(n34302), .Z(n34304) );
  AND U50474 ( .A(n34305), .B(n34304), .Z(n54055) );
  OR U50475 ( .A(n34306), .B(n54055), .Z(n34307) );
  NAND U50476 ( .A(n34308), .B(n34307), .Z(n34309) );
  NANDN U50477 ( .A(n34310), .B(n34309), .Z(n34311) );
  OR U50478 ( .A(n34311), .B(n52182), .Z(n34312) );
  NAND U50479 ( .A(n34313), .B(n34312), .Z(n34314) );
  NANDN U50480 ( .A(n34315), .B(n34314), .Z(n34317) );
  OR U50481 ( .A(n34317), .B(n34316), .Z(n34318) );
  AND U50482 ( .A(n34319), .B(n34318), .Z(n34321) );
  NOR U50483 ( .A(n34321), .B(n34320), .Z(n34322) );
  NAND U50484 ( .A(n54061), .B(n34322), .Z(n34323) );
  AND U50485 ( .A(n34324), .B(n34323), .Z(n34325) );
  OR U50486 ( .A(n34325), .B(n54063), .Z(n34326) );
  AND U50487 ( .A(n34327), .B(n34326), .Z(n34328) );
  OR U50488 ( .A(n34329), .B(n34328), .Z(n34330) );
  NAND U50489 ( .A(n34331), .B(n34330), .Z(n34332) );
  NAND U50490 ( .A(n34333), .B(n34332), .Z(n34334) );
  NAND U50491 ( .A(n54068), .B(n34334), .Z(n34335) );
  AND U50492 ( .A(n54069), .B(n34335), .Z(n34338) );
  NANDN U50493 ( .A(n34338), .B(n54070), .Z(n34339) );
  NAND U50494 ( .A(n54071), .B(n34339), .Z(n34340) );
  NANDN U50495 ( .A(n34341), .B(n34340), .Z(n34342) );
  OR U50496 ( .A(n54072), .B(n34342), .Z(n34343) );
  AND U50497 ( .A(n34344), .B(n34343), .Z(n34345) );
  NANDN U50498 ( .A(n54074), .B(n34345), .Z(n34346) );
  NAND U50499 ( .A(n34347), .B(n34346), .Z(n34351) );
  NAND U50500 ( .A(n34349), .B(n34348), .Z(n34350) );
  ANDN U50501 ( .B(n34351), .A(n34350), .Z(n34355) );
  NAND U50502 ( .A(n34353), .B(n34352), .Z(n34354) );
  OR U50503 ( .A(n34355), .B(n34354), .Z(n34356) );
  AND U50504 ( .A(n34357), .B(n34356), .Z(n34361) );
  NAND U50505 ( .A(n34359), .B(n34358), .Z(n34360) );
  OR U50506 ( .A(n34361), .B(n34360), .Z(n34362) );
  AND U50507 ( .A(n34363), .B(n34362), .Z(n34367) );
  NAND U50508 ( .A(n34365), .B(n34364), .Z(n34366) );
  OR U50509 ( .A(n34367), .B(n34366), .Z(n34368) );
  AND U50510 ( .A(n34369), .B(n34368), .Z(n34373) );
  NAND U50511 ( .A(n34371), .B(n34370), .Z(n34372) );
  OR U50512 ( .A(n34373), .B(n34372), .Z(n34374) );
  AND U50513 ( .A(n34375), .B(n34374), .Z(n34379) );
  NAND U50514 ( .A(n34377), .B(n34376), .Z(n34378) );
  OR U50515 ( .A(n34379), .B(n34378), .Z(n34380) );
  AND U50516 ( .A(n34381), .B(n34380), .Z(n34385) );
  NAND U50517 ( .A(n34383), .B(n34382), .Z(n34384) );
  OR U50518 ( .A(n34385), .B(n34384), .Z(n34386) );
  AND U50519 ( .A(n34387), .B(n34386), .Z(n34388) );
  OR U50520 ( .A(n34389), .B(n34388), .Z(n34390) );
  NAND U50521 ( .A(n34391), .B(n34390), .Z(n34395) );
  AND U50522 ( .A(n34393), .B(n34392), .Z(n34394) );
  NAND U50523 ( .A(n34395), .B(n34394), .Z(n34396) );
  NANDN U50524 ( .A(n34397), .B(n34396), .Z(n34399) );
  OR U50525 ( .A(n34399), .B(n34398), .Z(n34400) );
  NAND U50526 ( .A(n34401), .B(n34400), .Z(n34402) );
  NANDN U50527 ( .A(n34403), .B(n34402), .Z(n34404) );
  OR U50528 ( .A(n34405), .B(n34404), .Z(n34406) );
  AND U50529 ( .A(n34407), .B(n34406), .Z(n34409) );
  NAND U50530 ( .A(n34409), .B(n34408), .Z(n34411) );
  AND U50531 ( .A(n34422), .B(n34421), .Z(n34423) );
  OR U50532 ( .A(n34424), .B(n34423), .Z(n34425) );
  NAND U50533 ( .A(n34426), .B(n34425), .Z(n34427) );
  NAND U50534 ( .A(n34428), .B(n34427), .Z(n34429) );
  NAND U50535 ( .A(n34430), .B(n34429), .Z(n34431) );
  AND U50536 ( .A(n34432), .B(n34431), .Z(n34434) );
  OR U50537 ( .A(n34434), .B(n34433), .Z(n34435) );
  NAND U50538 ( .A(n34436), .B(n34435), .Z(n34437) );
  NANDN U50539 ( .A(n34438), .B(n34437), .Z(n34439) );
  OR U50540 ( .A(n34439), .B(n54109), .Z(n34440) );
  AND U50541 ( .A(n34441), .B(n34440), .Z(n34445) );
  NAND U50542 ( .A(n34443), .B(n34442), .Z(n34444) );
  OR U50543 ( .A(n34445), .B(n34444), .Z(n34446) );
  AND U50544 ( .A(n34447), .B(n34446), .Z(n34448) );
  OR U50545 ( .A(n34449), .B(n34448), .Z(n34450) );
  NAND U50546 ( .A(n34451), .B(n34450), .Z(n34454) );
  AND U50547 ( .A(n34452), .B(n54114), .Z(n34453) );
  NAND U50548 ( .A(n34454), .B(n34453), .Z(n34455) );
  NANDN U50549 ( .A(n34456), .B(n34455), .Z(n34457) );
  OR U50550 ( .A(n34457), .B(n54117), .Z(n34458) );
  NAND U50551 ( .A(n54118), .B(n34458), .Z(n34459) );
  NANDN U50552 ( .A(n34460), .B(n34459), .Z(n34463) );
  AND U50553 ( .A(n34461), .B(n54120), .Z(n34462) );
  NAND U50554 ( .A(n34463), .B(n34462), .Z(n34464) );
  NANDN U50555 ( .A(n34465), .B(n34464), .Z(n34467) );
  OR U50556 ( .A(n34467), .B(n34466), .Z(n34468) );
  NAND U50557 ( .A(n34469), .B(n34468), .Z(n34470) );
  NANDN U50558 ( .A(n34471), .B(n34470), .Z(n34473) );
  OR U50559 ( .A(n34473), .B(n34472), .Z(n34474) );
  NAND U50560 ( .A(n34475), .B(n34474), .Z(n34476) );
  AND U50561 ( .A(n34477), .B(n34476), .Z(n34478) );
  OR U50562 ( .A(n34479), .B(n34478), .Z(n34480) );
  NAND U50563 ( .A(n34481), .B(n34480), .Z(n34482) );
  NANDN U50564 ( .A(n34483), .B(n34482), .Z(n34484) );
  NAND U50565 ( .A(n34485), .B(n34484), .Z(n34487) );
  ANDN U50566 ( .B(y[1998]), .A(x[1998]), .Z(n34486) );
  ANDN U50567 ( .B(n34487), .A(n34486), .Z(n34489) );
  ANDN U50568 ( .B(n34489), .A(n34488), .Z(n34493) );
  NAND U50569 ( .A(n34491), .B(n34490), .Z(n34492) );
  OR U50570 ( .A(n34493), .B(n34492), .Z(n34494) );
  AND U50571 ( .A(n34495), .B(n34494), .Z(n34496) );
  NOR U50572 ( .A(n54133), .B(n34496), .Z(n34497) );
  NANDN U50573 ( .A(n34498), .B(n34497), .Z(n34499) );
  AND U50574 ( .A(n34500), .B(n34499), .Z(n34501) );
  NANDN U50575 ( .A(n34502), .B(n34501), .Z(n34503) );
  NAND U50576 ( .A(n54134), .B(n34503), .Z(n34504) );
  NANDN U50577 ( .A(n34505), .B(n34504), .Z(n34508) );
  AND U50578 ( .A(n34506), .B(n52156), .Z(n34507) );
  NAND U50579 ( .A(n34508), .B(n34507), .Z(n34509) );
  NANDN U50580 ( .A(n34510), .B(n34509), .Z(n34511) );
  OR U50581 ( .A(n34512), .B(n34511), .Z(n34513) );
  AND U50582 ( .A(n34514), .B(n34513), .Z(n34515) );
  NAND U50583 ( .A(n34515), .B(n54139), .Z(n34517) );
  ANDN U50584 ( .B(n34517), .A(n34516), .Z(n34518) );
  NANDN U50585 ( .A(n54140), .B(n34518), .Z(n34519) );
  AND U50586 ( .A(n54141), .B(n34519), .Z(n34522) );
  NANDN U50587 ( .A(x[2010]), .B(y[2010]), .Z(n34521) );
  NAND U50588 ( .A(n34521), .B(n34520), .Z(n54142) );
  OR U50589 ( .A(n34522), .B(n54142), .Z(n34523) );
  AND U50590 ( .A(n34524), .B(n34523), .Z(n34525) );
  NAND U50591 ( .A(n34525), .B(n54143), .Z(n34527) );
  ANDN U50592 ( .B(n34527), .A(n34526), .Z(n34528) );
  NANDN U50593 ( .A(n54144), .B(n34528), .Z(n34532) );
  AND U50594 ( .A(n34530), .B(n34529), .Z(n34531) );
  NAND U50595 ( .A(n34532), .B(n34531), .Z(n34533) );
  NANDN U50596 ( .A(n34534), .B(n34533), .Z(n34536) );
  OR U50597 ( .A(n34536), .B(n34535), .Z(n34537) );
  NAND U50598 ( .A(n34538), .B(n34537), .Z(n34539) );
  NANDN U50599 ( .A(n34540), .B(n34539), .Z(n34541) );
  OR U50600 ( .A(n34541), .B(n54150), .Z(n34542) );
  AND U50601 ( .A(n34543), .B(n34542), .Z(n34544) );
  OR U50602 ( .A(n54152), .B(n34544), .Z(n34545) );
  NAND U50603 ( .A(n54153), .B(n34545), .Z(n34546) );
  NANDN U50604 ( .A(n54154), .B(n34546), .Z(n34547) );
  NAND U50605 ( .A(n54155), .B(n34547), .Z(n34549) );
  IV U50606 ( .A(n34548), .Z(n54156) );
  ANDN U50607 ( .B(n34549), .A(n54156), .Z(n34550) );
  NANDN U50608 ( .A(n34551), .B(n34550), .Z(n34554) );
  AND U50609 ( .A(n34552), .B(n54157), .Z(n34553) );
  NAND U50610 ( .A(n34554), .B(n34553), .Z(n34555) );
  NANDN U50611 ( .A(n34556), .B(n34555), .Z(n34558) );
  ANDN U50612 ( .B(y[2024]), .A(x[2024]), .Z(n34557) );
  OR U50613 ( .A(n34558), .B(n34557), .Z(n34559) );
  NAND U50614 ( .A(n34560), .B(n34559), .Z(n34561) );
  NANDN U50615 ( .A(n34562), .B(n34561), .Z(n34564) );
  OR U50616 ( .A(n34564), .B(n34563), .Z(n34565) );
  NAND U50617 ( .A(n54166), .B(n34565), .Z(n34566) );
  NANDN U50618 ( .A(n54165), .B(n34566), .Z(n34567) );
  OR U50619 ( .A(n34568), .B(n34567), .Z(n34569) );
  AND U50620 ( .A(n34570), .B(n34569), .Z(n34571) );
  NAND U50621 ( .A(n34571), .B(n54164), .Z(n34573) );
  ANDN U50622 ( .B(y[2030]), .A(x[2030]), .Z(n34572) );
  ANDN U50623 ( .B(n34573), .A(n34572), .Z(n34574) );
  NANDN U50624 ( .A(n34575), .B(n34574), .Z(n34576) );
  NAND U50625 ( .A(n34577), .B(n34576), .Z(n34578) );
  NANDN U50626 ( .A(n34579), .B(n34578), .Z(n34580) );
  AND U50627 ( .A(n34581), .B(n34580), .Z(n34582) );
  OR U50628 ( .A(n34583), .B(n34582), .Z(n34584) );
  NAND U50629 ( .A(n34585), .B(n34584), .Z(n34589) );
  NANDN U50630 ( .A(x[2036]), .B(y[2036]), .Z(n34586) );
  AND U50631 ( .A(n34587), .B(n34586), .Z(n34588) );
  NAND U50632 ( .A(n34589), .B(n34588), .Z(n34593) );
  NAND U50633 ( .A(n34591), .B(n34590), .Z(n34592) );
  ANDN U50634 ( .B(n34593), .A(n34592), .Z(n34597) );
  NAND U50635 ( .A(n34595), .B(n34594), .Z(n34596) );
  OR U50636 ( .A(n34597), .B(n34596), .Z(n34598) );
  AND U50637 ( .A(n34599), .B(n34598), .Z(n34603) );
  NAND U50638 ( .A(n34601), .B(n34600), .Z(n34602) );
  OR U50639 ( .A(n34603), .B(n34602), .Z(n34604) );
  AND U50640 ( .A(n34605), .B(n34604), .Z(n34606) );
  ANDN U50641 ( .B(n34607), .A(n34606), .Z(n34608) );
  NAND U50642 ( .A(n34609), .B(n34608), .Z(n34610) );
  NANDN U50643 ( .A(n34611), .B(n34610), .Z(n34613) );
  OR U50644 ( .A(n34613), .B(n34612), .Z(n34614) );
  NAND U50645 ( .A(n34615), .B(n34614), .Z(n34616) );
  NANDN U50646 ( .A(n34617), .B(n34616), .Z(n34618) );
  OR U50647 ( .A(n34619), .B(n34618), .Z(n34620) );
  AND U50648 ( .A(n34621), .B(n34620), .Z(n34623) );
  NAND U50649 ( .A(n34623), .B(n34622), .Z(n34625) );
  ANDN U50650 ( .B(n34625), .A(n34624), .Z(n34626) );
  NANDN U50651 ( .A(n34627), .B(n34626), .Z(n34628) );
  AND U50652 ( .A(n34629), .B(n34628), .Z(n34630) );
  NAND U50653 ( .A(n34631), .B(n34630), .Z(n34632) );
  NANDN U50654 ( .A(n54187), .B(n34632), .Z(n34634) );
  OR U50655 ( .A(n34634), .B(n34633), .Z(n34635) );
  NAND U50656 ( .A(n34636), .B(n34635), .Z(n34637) );
  NANDN U50657 ( .A(n54189), .B(n34637), .Z(n34640) );
  AND U50658 ( .A(n34638), .B(n54190), .Z(n34639) );
  NAND U50659 ( .A(n34640), .B(n34639), .Z(n34641) );
  NANDN U50660 ( .A(n34642), .B(n34641), .Z(n34643) );
  OR U50661 ( .A(n34643), .B(n54191), .Z(n34644) );
  NAND U50662 ( .A(n34645), .B(n34644), .Z(n34646) );
  NANDN U50663 ( .A(n34647), .B(n34646), .Z(n34648) );
  OR U50664 ( .A(n34648), .B(n54195), .Z(n34649) );
  AND U50665 ( .A(n34650), .B(n34649), .Z(n34659) );
  OR U50666 ( .A(n34652), .B(n34651), .Z(n34653) );
  NAND U50667 ( .A(n34654), .B(n34653), .Z(n34655) );
  NANDN U50668 ( .A(n34656), .B(n34655), .Z(n34658) );
  XNOR U50669 ( .A(y[2060]), .B(x[2060]), .Z(n34657) );
  NANDN U50670 ( .A(n34658), .B(n34657), .Z(n54199) );
  OR U50671 ( .A(n34659), .B(n54199), .Z(n34660) );
  NAND U50672 ( .A(n54200), .B(n34660), .Z(n34661) );
  NANDN U50673 ( .A(n34662), .B(n34661), .Z(n34664) );
  IV U50674 ( .A(n34663), .Z(n54201) );
  OR U50675 ( .A(n34664), .B(n54201), .Z(n34665) );
  NAND U50676 ( .A(n34666), .B(n34665), .Z(n34667) );
  NANDN U50677 ( .A(n34668), .B(n34667), .Z(n34670) );
  OR U50678 ( .A(n34670), .B(n34669), .Z(n34671) );
  NAND U50679 ( .A(n34672), .B(n34671), .Z(n34676) );
  AND U50680 ( .A(n34674), .B(n34673), .Z(n34675) );
  NAND U50681 ( .A(n34676), .B(n34675), .Z(n34677) );
  NANDN U50682 ( .A(n34678), .B(n34677), .Z(n34680) );
  OR U50683 ( .A(n34680), .B(n34679), .Z(n34681) );
  NAND U50684 ( .A(n34682), .B(n34681), .Z(n34683) );
  NANDN U50685 ( .A(n34684), .B(n34683), .Z(n34686) );
  OR U50686 ( .A(n34686), .B(n34685), .Z(n34687) );
  AND U50687 ( .A(n34688), .B(n34687), .Z(n34689) );
  OR U50688 ( .A(n34690), .B(n34689), .Z(n34691) );
  NAND U50689 ( .A(n34692), .B(n34691), .Z(n34693) );
  NANDN U50690 ( .A(n34694), .B(n34693), .Z(n34698) );
  AND U50691 ( .A(n34696), .B(n34695), .Z(n34697) );
  NAND U50692 ( .A(n34698), .B(n34697), .Z(n34699) );
  NANDN U50693 ( .A(n34700), .B(n34699), .Z(n34702) );
  OR U50694 ( .A(n34702), .B(n34701), .Z(n34703) );
  NAND U50695 ( .A(n34704), .B(n34703), .Z(n34705) );
  NANDN U50696 ( .A(n52149), .B(n34705), .Z(n34707) );
  OR U50697 ( .A(n34707), .B(n34706), .Z(n34708) );
  AND U50698 ( .A(n34709), .B(n34708), .Z(n34710) );
  OR U50699 ( .A(n34711), .B(n34710), .Z(n34712) );
  NAND U50700 ( .A(n54227), .B(n34712), .Z(n34713) );
  NANDN U50701 ( .A(n34714), .B(n34713), .Z(n34716) );
  NAND U50702 ( .A(n34716), .B(n34715), .Z(n34718) );
  ANDN U50703 ( .B(n34718), .A(n34717), .Z(n34719) );
  NANDN U50704 ( .A(n54233), .B(n34719), .Z(n34723) );
  IV U50705 ( .A(n34720), .Z(n54235) );
  AND U50706 ( .A(n34721), .B(n54235), .Z(n34722) );
  NAND U50707 ( .A(n34723), .B(n34722), .Z(n34724) );
  NANDN U50708 ( .A(n54238), .B(n34724), .Z(n34725) );
  OR U50709 ( .A(n34726), .B(n34725), .Z(n34727) );
  AND U50710 ( .A(n34728), .B(n34727), .Z(n34729) );
  OR U50711 ( .A(n34730), .B(n34729), .Z(n34731) );
  NAND U50712 ( .A(n54248), .B(n34731), .Z(n34732) );
  NANDN U50713 ( .A(n54250), .B(n34732), .Z(n34733) );
  AND U50714 ( .A(n54251), .B(n34733), .Z(n34736) );
  OR U50715 ( .A(n34736), .B(n54252), .Z(n34737) );
  AND U50716 ( .A(n34738), .B(n34737), .Z(n34739) );
  NAND U50717 ( .A(n34739), .B(n54253), .Z(n34741) );
  ANDN U50718 ( .B(n34741), .A(n34740), .Z(n34742) );
  NANDN U50719 ( .A(n54254), .B(n34742), .Z(n34746) );
  AND U50720 ( .A(n34744), .B(n34743), .Z(n34745) );
  NAND U50721 ( .A(n34746), .B(n34745), .Z(n34747) );
  NANDN U50722 ( .A(n34748), .B(n34747), .Z(n34750) );
  OR U50723 ( .A(n34750), .B(n34749), .Z(n34751) );
  NAND U50724 ( .A(n34752), .B(n34751), .Z(n34753) );
  NANDN U50725 ( .A(n34754), .B(n34753), .Z(n34755) );
  OR U50726 ( .A(n34756), .B(n34755), .Z(n34757) );
  AND U50727 ( .A(n34758), .B(n34757), .Z(n34760) );
  NAND U50728 ( .A(n34760), .B(n34759), .Z(n34762) );
  ANDN U50729 ( .B(n34762), .A(n34761), .Z(n34763) );
  NANDN U50730 ( .A(n34764), .B(n34763), .Z(n34768) );
  AND U50731 ( .A(n34766), .B(n34765), .Z(n34767) );
  NAND U50732 ( .A(n34768), .B(n34767), .Z(n34769) );
  NANDN U50733 ( .A(n34770), .B(n34769), .Z(n34772) );
  OR U50734 ( .A(n34772), .B(n34771), .Z(n34773) );
  NAND U50735 ( .A(n34774), .B(n34773), .Z(n34775) );
  NANDN U50736 ( .A(n34776), .B(n34775), .Z(n34777) );
  OR U50737 ( .A(n34778), .B(n34777), .Z(n34779) );
  AND U50738 ( .A(n34780), .B(n34779), .Z(n34782) );
  NAND U50739 ( .A(n34782), .B(n34781), .Z(n34784) );
  ANDN U50740 ( .B(n34784), .A(n34783), .Z(n34785) );
  NANDN U50741 ( .A(n34786), .B(n34785), .Z(n34790) );
  AND U50742 ( .A(n34788), .B(n34787), .Z(n34789) );
  NAND U50743 ( .A(n34790), .B(n34789), .Z(n34791) );
  NANDN U50744 ( .A(n34792), .B(n34791), .Z(n34795) );
  NANDN U50745 ( .A(x[2109]), .B(n34795), .Z(n34794) );
  ANDN U50746 ( .B(n34794), .A(n34793), .Z(n34798) );
  XNOR U50747 ( .A(n34795), .B(x[2109]), .Z(n34796) );
  NAND U50748 ( .A(n34796), .B(y[2109]), .Z(n34797) );
  NAND U50749 ( .A(n34798), .B(n34797), .Z(n34800) );
  IV U50750 ( .A(n34799), .Z(n54269) );
  AND U50751 ( .A(n34800), .B(n54269), .Z(n34802) );
  IV U50752 ( .A(n34801), .Z(n54270) );
  OR U50753 ( .A(n34802), .B(n54270), .Z(n34803) );
  NAND U50754 ( .A(n54271), .B(n34803), .Z(n34804) );
  NANDN U50755 ( .A(n54272), .B(n34804), .Z(n34805) );
  NAND U50756 ( .A(n54273), .B(n34805), .Z(n34806) );
  NANDN U50757 ( .A(n54274), .B(n34806), .Z(n34807) );
  AND U50758 ( .A(n34808), .B(n34807), .Z(n34809) );
  OR U50759 ( .A(n34810), .B(n34809), .Z(n34811) );
  NAND U50760 ( .A(n34812), .B(n34811), .Z(n34813) );
  NANDN U50761 ( .A(n34814), .B(n34813), .Z(n34815) );
  OR U50762 ( .A(n34816), .B(n34815), .Z(n34817) );
  AND U50763 ( .A(n34818), .B(n34817), .Z(n34820) );
  NAND U50764 ( .A(n34820), .B(n34819), .Z(n34822) );
  ANDN U50765 ( .B(n34822), .A(n34821), .Z(n34823) );
  NANDN U50766 ( .A(n34824), .B(n34823), .Z(n34828) );
  AND U50767 ( .A(n34826), .B(n34825), .Z(n34827) );
  NAND U50768 ( .A(n34828), .B(n34827), .Z(n34829) );
  NANDN U50769 ( .A(n34830), .B(n34829), .Z(n34832) );
  ANDN U50770 ( .B(y[2122]), .A(x[2122]), .Z(n34831) );
  OR U50771 ( .A(n34832), .B(n34831), .Z(n34833) );
  NAND U50772 ( .A(n34834), .B(n34833), .Z(n34835) );
  NANDN U50773 ( .A(n34836), .B(n34835), .Z(n34837) );
  OR U50774 ( .A(n34838), .B(n34837), .Z(n34839) );
  AND U50775 ( .A(n34840), .B(n34839), .Z(n34841) );
  NANDN U50776 ( .A(n34842), .B(n34841), .Z(n34843) );
  NAND U50777 ( .A(n34844), .B(n34843), .Z(n34845) );
  NANDN U50778 ( .A(n34846), .B(n34845), .Z(n34847) );
  AND U50779 ( .A(n54287), .B(n34847), .Z(n34848) );
  OR U50780 ( .A(n34849), .B(n34848), .Z(n34850) );
  NAND U50781 ( .A(n34851), .B(n34850), .Z(n34852) );
  NANDN U50782 ( .A(n34853), .B(n34852), .Z(n34854) );
  NAND U50783 ( .A(n34855), .B(n34854), .Z(n34857) );
  AND U50784 ( .A(n34857), .B(n34856), .Z(n34859) );
  OR U50785 ( .A(n34859), .B(n34858), .Z(n34860) );
  NAND U50786 ( .A(n34861), .B(n34860), .Z(n34862) );
  NANDN U50787 ( .A(n34863), .B(n34862), .Z(n34865) );
  OR U50788 ( .A(n34865), .B(n34864), .Z(n34866) );
  NAND U50789 ( .A(n34867), .B(n34866), .Z(n34868) );
  NANDN U50790 ( .A(n34869), .B(n34868), .Z(n34870) );
  OR U50791 ( .A(n34871), .B(n34870), .Z(n34872) );
  AND U50792 ( .A(n34873), .B(n34872), .Z(n34875) );
  NAND U50793 ( .A(n34875), .B(n34874), .Z(n34877) );
  ANDN U50794 ( .B(n34877), .A(n34876), .Z(n34878) );
  NANDN U50795 ( .A(n34879), .B(n34878), .Z(n34883) );
  AND U50796 ( .A(n34881), .B(n34880), .Z(n34882) );
  NAND U50797 ( .A(n34883), .B(n34882), .Z(n34884) );
  NANDN U50798 ( .A(n34885), .B(n34884), .Z(n34887) );
  OR U50799 ( .A(n34887), .B(n34886), .Z(n34888) );
  NAND U50800 ( .A(n34889), .B(n34888), .Z(n34890) );
  NANDN U50801 ( .A(n34891), .B(n34890), .Z(n34893) );
  OR U50802 ( .A(n34893), .B(n34892), .Z(n34894) );
  AND U50803 ( .A(n34895), .B(n34894), .Z(n34899) );
  NAND U50804 ( .A(n34897), .B(n34896), .Z(n34898) );
  OR U50805 ( .A(n34899), .B(n34898), .Z(n34900) );
  AND U50806 ( .A(n34901), .B(n34900), .Z(n34902) );
  ANDN U50807 ( .B(n34903), .A(n34902), .Z(n34904) );
  NAND U50808 ( .A(n34905), .B(n34904), .Z(n34906) );
  NANDN U50809 ( .A(n54306), .B(n34906), .Z(n34908) );
  OR U50810 ( .A(n34908), .B(n34907), .Z(n34909) );
  NAND U50811 ( .A(n34910), .B(n34909), .Z(n34911) );
  NAND U50812 ( .A(n54308), .B(n34911), .Z(n34912) );
  AND U50813 ( .A(n54309), .B(n34912), .Z(n34915) );
  NANDN U50814 ( .A(n34915), .B(n54310), .Z(n34916) );
  AND U50815 ( .A(n54311), .B(n34916), .Z(n34917) );
  ANDN U50816 ( .B(n34918), .A(n34917), .Z(n34919) );
  NAND U50817 ( .A(n54312), .B(n34919), .Z(n34920) );
  NANDN U50818 ( .A(n34921), .B(n34920), .Z(n34922) );
  OR U50819 ( .A(n54313), .B(n34922), .Z(n34923) );
  AND U50820 ( .A(n34924), .B(n34923), .Z(n34926) );
  NAND U50821 ( .A(n34926), .B(n34925), .Z(n34928) );
  ANDN U50822 ( .B(n34928), .A(n34927), .Z(n34929) );
  NANDN U50823 ( .A(n34930), .B(n34929), .Z(n34934) );
  AND U50824 ( .A(n34932), .B(n34931), .Z(n34933) );
  NAND U50825 ( .A(n34934), .B(n34933), .Z(n34935) );
  NANDN U50826 ( .A(n34936), .B(n34935), .Z(n34937) );
  OR U50827 ( .A(n54320), .B(n34937), .Z(n34938) );
  AND U50828 ( .A(n54321), .B(n34938), .Z(n34939) );
  NANDN U50829 ( .A(n34940), .B(n34939), .Z(n34941) );
  NAND U50830 ( .A(n54322), .B(n34941), .Z(n34942) );
  NANDN U50831 ( .A(n54323), .B(n34942), .Z(n34943) );
  AND U50832 ( .A(n54324), .B(n34943), .Z(n34944) );
  OR U50833 ( .A(n54325), .B(n34944), .Z(n34945) );
  NAND U50834 ( .A(n54326), .B(n34945), .Z(n34946) );
  NANDN U50835 ( .A(n34947), .B(n34946), .Z(n34949) );
  IV U50836 ( .A(n34948), .Z(n54327) );
  OR U50837 ( .A(n34949), .B(n54327), .Z(n34950) );
  AND U50838 ( .A(n34951), .B(n34950), .Z(n34955) );
  NAND U50839 ( .A(n34953), .B(n34952), .Z(n34954) );
  OR U50840 ( .A(n34955), .B(n34954), .Z(n34956) );
  AND U50841 ( .A(n34957), .B(n34956), .Z(n34959) );
  NOR U50842 ( .A(n34959), .B(n34958), .Z(n34960) );
  NANDN U50843 ( .A(n34961), .B(n34960), .Z(n34962) );
  AND U50844 ( .A(n34962), .B(n54334), .Z(n34963) );
  NANDN U50845 ( .A(n34964), .B(n34963), .Z(n34965) );
  AND U50846 ( .A(n34966), .B(n34965), .Z(n34967) );
  NANDN U50847 ( .A(n34968), .B(n34967), .Z(n34969) );
  AND U50848 ( .A(n54339), .B(n34969), .Z(n34970) );
  ANDN U50849 ( .B(n34971), .A(n34970), .Z(n34972) );
  NAND U50850 ( .A(n54338), .B(n34972), .Z(n34973) );
  NANDN U50851 ( .A(n54337), .B(n34973), .Z(n34975) );
  OR U50852 ( .A(n34975), .B(n34974), .Z(n34976) );
  NAND U50853 ( .A(n34977), .B(n34976), .Z(n34978) );
  NANDN U50854 ( .A(n34979), .B(n34978), .Z(n34981) );
  OR U50855 ( .A(n34981), .B(n34980), .Z(n34982) );
  NAND U50856 ( .A(n34983), .B(n34982), .Z(n34986) );
  AND U50857 ( .A(n34984), .B(n52143), .Z(n34985) );
  NAND U50858 ( .A(n34986), .B(n34985), .Z(n34987) );
  NANDN U50859 ( .A(n54345), .B(n34987), .Z(n34989) );
  OR U50860 ( .A(n34989), .B(n34988), .Z(n34990) );
  NAND U50861 ( .A(n34991), .B(n34990), .Z(n34992) );
  NANDN U50862 ( .A(n34993), .B(n34992), .Z(n34997) );
  IV U50863 ( .A(n34994), .Z(n54347) );
  AND U50864 ( .A(n34995), .B(n54347), .Z(n34996) );
  NAND U50865 ( .A(n34997), .B(n34996), .Z(n34998) );
  NANDN U50866 ( .A(n34999), .B(n34998), .Z(n35001) );
  OR U50867 ( .A(n35001), .B(n35000), .Z(n35002) );
  NAND U50868 ( .A(n35003), .B(n35002), .Z(n35004) );
  NANDN U50869 ( .A(n35005), .B(n35004), .Z(n35006) );
  OR U50870 ( .A(n35007), .B(n35006), .Z(n35008) );
  AND U50871 ( .A(n35009), .B(n35008), .Z(n35011) );
  NAND U50872 ( .A(n35011), .B(n35010), .Z(n35013) );
  ANDN U50873 ( .B(n35013), .A(n35012), .Z(n35014) );
  NANDN U50874 ( .A(n35015), .B(n35014), .Z(n35019) );
  NANDN U50875 ( .A(x[2186]), .B(y[2186]), .Z(n35016) );
  AND U50876 ( .A(n35017), .B(n35016), .Z(n35018) );
  NAND U50877 ( .A(n35019), .B(n35018), .Z(n35020) );
  NANDN U50878 ( .A(n35021), .B(n35020), .Z(n35022) );
  OR U50879 ( .A(n35023), .B(n35022), .Z(n35024) );
  AND U50880 ( .A(n35025), .B(n35024), .Z(n35027) );
  NANDN U50881 ( .A(x[2188]), .B(y[2188]), .Z(n35026) );
  AND U50882 ( .A(n35027), .B(n35026), .Z(n35031) );
  NAND U50883 ( .A(n35029), .B(n35028), .Z(n35030) );
  OR U50884 ( .A(n35031), .B(n35030), .Z(n35033) );
  IV U50885 ( .A(n35032), .Z(n54355) );
  AND U50886 ( .A(n35033), .B(n54355), .Z(n35035) );
  NANDN U50887 ( .A(x[2190]), .B(y[2190]), .Z(n35034) );
  AND U50888 ( .A(n35035), .B(n35034), .Z(n35036) );
  OR U50889 ( .A(n54356), .B(n35036), .Z(n35037) );
  NAND U50890 ( .A(n54357), .B(n35037), .Z(n35038) );
  NANDN U50891 ( .A(n54358), .B(n35038), .Z(n35039) );
  AND U50892 ( .A(n54360), .B(n35039), .Z(n35040) );
  OR U50893 ( .A(n54361), .B(n35040), .Z(n35041) );
  NAND U50894 ( .A(n54362), .B(n35041), .Z(n35042) );
  NANDN U50895 ( .A(n54363), .B(n35042), .Z(n35043) );
  NAND U50896 ( .A(n52134), .B(n35043), .Z(n35044) );
  ANDN U50897 ( .B(n35044), .A(n54364), .Z(n35045) );
  NANDN U50898 ( .A(n35046), .B(n35045), .Z(n35049) );
  AND U50899 ( .A(n35047), .B(n54365), .Z(n35048) );
  NAND U50900 ( .A(n35049), .B(n35048), .Z(n35050) );
  NANDN U50901 ( .A(n35051), .B(n35050), .Z(n35052) );
  OR U50902 ( .A(n35053), .B(n35052), .Z(n35054) );
  AND U50903 ( .A(n35055), .B(n35054), .Z(n35056) );
  NANDN U50904 ( .A(n35057), .B(n35056), .Z(n35058) );
  AND U50905 ( .A(n35059), .B(n35058), .Z(n35060) );
  NANDN U50906 ( .A(n35061), .B(n35060), .Z(n35062) );
  AND U50907 ( .A(n35063), .B(n35062), .Z(n35067) );
  NAND U50908 ( .A(n35065), .B(n35064), .Z(n35066) );
  OR U50909 ( .A(n35067), .B(n35066), .Z(n35068) );
  AND U50910 ( .A(n35069), .B(n35068), .Z(n35070) );
  ANDN U50911 ( .B(n35071), .A(n35070), .Z(n35072) );
  NAND U50912 ( .A(n35073), .B(n35072), .Z(n35074) );
  NANDN U50913 ( .A(n52130), .B(n35074), .Z(n35075) );
  OR U50914 ( .A(n35076), .B(n35075), .Z(n35077) );
  AND U50915 ( .A(n54375), .B(n35077), .Z(n35078) );
  NANDN U50916 ( .A(n35079), .B(n35078), .Z(n35080) );
  NAND U50917 ( .A(n52129), .B(n35080), .Z(n35081) );
  NANDN U50918 ( .A(n54376), .B(n35081), .Z(n35083) );
  IV U50919 ( .A(n35082), .Z(n54377) );
  AND U50920 ( .A(n35083), .B(n54377), .Z(n35085) );
  IV U50921 ( .A(n35084), .Z(n54378) );
  OR U50922 ( .A(n35085), .B(n54378), .Z(n35086) );
  NAND U50923 ( .A(n54379), .B(n35086), .Z(n35087) );
  NANDN U50924 ( .A(n35088), .B(n35087), .Z(n35090) );
  IV U50925 ( .A(n35089), .Z(n54380) );
  OR U50926 ( .A(n35090), .B(n54380), .Z(n35091) );
  NANDN U50927 ( .A(n54381), .B(n35091), .Z(n35092) );
  AND U50928 ( .A(n35093), .B(n35092), .Z(n35095) );
  IV U50929 ( .A(n35094), .Z(n54383) );
  NANDN U50930 ( .A(n35095), .B(n54383), .Z(n35096) );
  NANDN U50931 ( .A(n54384), .B(n35096), .Z(n35097) );
  AND U50932 ( .A(n35098), .B(n35097), .Z(n35099) );
  OR U50933 ( .A(n35100), .B(n35099), .Z(n35101) );
  NAND U50934 ( .A(n35102), .B(n35101), .Z(n35103) );
  NANDN U50935 ( .A(n35104), .B(n35103), .Z(n35106) );
  OR U50936 ( .A(n35106), .B(n35105), .Z(n35107) );
  AND U50937 ( .A(n35108), .B(n35107), .Z(n35109) );
  OR U50938 ( .A(n35110), .B(n35109), .Z(n35111) );
  NAND U50939 ( .A(n35112), .B(n35111), .Z(n35113) );
  AND U50940 ( .A(n35114), .B(n35113), .Z(n35115) );
  OR U50941 ( .A(n35116), .B(n35115), .Z(n35117) );
  NAND U50942 ( .A(n54391), .B(n35117), .Z(n35118) );
  NANDN U50943 ( .A(n54392), .B(n35118), .Z(n35119) );
  NAND U50944 ( .A(n54393), .B(n35119), .Z(n35120) );
  NAND U50945 ( .A(n35121), .B(n35120), .Z(n35122) );
  NANDN U50946 ( .A(n35123), .B(n35122), .Z(n35124) );
  AND U50947 ( .A(n35125), .B(n35124), .Z(n35126) );
  NAND U50948 ( .A(n35127), .B(n35126), .Z(n35128) );
  NANDN U50949 ( .A(n35129), .B(n35128), .Z(n35133) );
  AND U50950 ( .A(n35131), .B(n35130), .Z(n35132) );
  NAND U50951 ( .A(n35133), .B(n35132), .Z(n35134) );
  NANDN U50952 ( .A(n35135), .B(n35134), .Z(n35136) );
  OR U50953 ( .A(n35137), .B(n35136), .Z(n35138) );
  AND U50954 ( .A(n35139), .B(n35138), .Z(n35141) );
  NAND U50955 ( .A(n35141), .B(n35140), .Z(n35143) );
  ANDN U50956 ( .B(n35143), .A(n35142), .Z(n35144) );
  NANDN U50957 ( .A(n35145), .B(n35144), .Z(n35149) );
  IV U50958 ( .A(n35146), .Z(n54402) );
  AND U50959 ( .A(n35147), .B(n54402), .Z(n35148) );
  NAND U50960 ( .A(n35149), .B(n35148), .Z(n35150) );
  NANDN U50961 ( .A(n54404), .B(n35150), .Z(n35151) );
  OR U50962 ( .A(n35152), .B(n35151), .Z(n35153) );
  AND U50963 ( .A(n35154), .B(n35153), .Z(n35156) );
  NANDN U50964 ( .A(n35156), .B(n35155), .Z(n35157) );
  NANDN U50965 ( .A(n35158), .B(n35157), .Z(n35159) );
  AND U50966 ( .A(n35160), .B(n35159), .Z(n35162) );
  NANDN U50967 ( .A(n35162), .B(n35161), .Z(n35163) );
  AND U50968 ( .A(n35164), .B(n35163), .Z(n35165) );
  NANDN U50969 ( .A(n54406), .B(n35165), .Z(n35166) );
  AND U50970 ( .A(n35167), .B(n35166), .Z(n35168) );
  OR U50971 ( .A(n35169), .B(n35168), .Z(n35170) );
  NAND U50972 ( .A(n35171), .B(n35170), .Z(n35175) );
  IV U50973 ( .A(n35172), .Z(n54413) );
  AND U50974 ( .A(n35173), .B(n54413), .Z(n35174) );
  NAND U50975 ( .A(n35175), .B(n35174), .Z(n35176) );
  NANDN U50976 ( .A(n35177), .B(n35176), .Z(n35179) );
  IV U50977 ( .A(n35178), .Z(n54414) );
  OR U50978 ( .A(n35179), .B(n54414), .Z(n35180) );
  AND U50979 ( .A(n54415), .B(n35180), .Z(n35183) );
  NAND U50980 ( .A(n35182), .B(n35181), .Z(n54416) );
  OR U50981 ( .A(n35183), .B(n54416), .Z(n35184) );
  AND U50982 ( .A(n54417), .B(n35184), .Z(n35185) );
  OR U50983 ( .A(n54418), .B(n35185), .Z(n35186) );
  NAND U50984 ( .A(n35187), .B(n35186), .Z(n35188) );
  NANDN U50985 ( .A(n35189), .B(n35188), .Z(n35191) );
  IV U50986 ( .A(n35190), .Z(n54420) );
  OR U50987 ( .A(n35191), .B(n54420), .Z(n35192) );
  NAND U50988 ( .A(n35193), .B(n35192), .Z(n35194) );
  OR U50989 ( .A(n35195), .B(n35194), .Z(n35196) );
  AND U50990 ( .A(n35197), .B(n35196), .Z(n35199) );
  NANDN U50991 ( .A(x[2258]), .B(y[2258]), .Z(n35198) );
  NAND U50992 ( .A(n35199), .B(n35198), .Z(n35201) );
  ANDN U50993 ( .B(n35201), .A(n35200), .Z(n35202) );
  NANDN U50994 ( .A(n35203), .B(n35202), .Z(n35204) );
  AND U50995 ( .A(n35205), .B(n35204), .Z(n35206) );
  NOR U50996 ( .A(n35207), .B(n35206), .Z(n35209) );
  NAND U50997 ( .A(n35209), .B(n35208), .Z(n35213) );
  NANDN U50998 ( .A(x[2262]), .B(y[2262]), .Z(n35210) );
  AND U50999 ( .A(n35211), .B(n35210), .Z(n35212) );
  NAND U51000 ( .A(n35213), .B(n35212), .Z(n35217) );
  NAND U51001 ( .A(n35215), .B(n35214), .Z(n35216) );
  ANDN U51002 ( .B(n35217), .A(n35216), .Z(n35221) );
  NAND U51003 ( .A(n35219), .B(n35218), .Z(n35220) );
  OR U51004 ( .A(n35221), .B(n35220), .Z(n35222) );
  AND U51005 ( .A(n35223), .B(n35222), .Z(n35225) );
  NOR U51006 ( .A(n35225), .B(n35224), .Z(n35226) );
  NANDN U51007 ( .A(n35227), .B(n35226), .Z(n35229) );
  IV U51008 ( .A(n35228), .Z(n54433) );
  AND U51009 ( .A(n35229), .B(n54433), .Z(n35230) );
  NANDN U51010 ( .A(n35231), .B(n35230), .Z(n35232) );
  AND U51011 ( .A(n35233), .B(n35232), .Z(n35234) );
  NANDN U51012 ( .A(n54434), .B(n35234), .Z(n35235) );
  AND U51013 ( .A(n54435), .B(n35235), .Z(n35236) );
  OR U51014 ( .A(n54437), .B(n35236), .Z(n35237) );
  NAND U51015 ( .A(n54438), .B(n35237), .Z(n35238) );
  NANDN U51016 ( .A(n54439), .B(n35238), .Z(n35241) );
  AND U51017 ( .A(n35239), .B(n54440), .Z(n35240) );
  NAND U51018 ( .A(n35241), .B(n35240), .Z(n35242) );
  NANDN U51019 ( .A(n35243), .B(n35242), .Z(n35245) );
  IV U51020 ( .A(n35244), .Z(n54441) );
  OR U51021 ( .A(n35245), .B(n54441), .Z(n35246) );
  AND U51022 ( .A(n35247), .B(n35246), .Z(n35248) );
  OR U51023 ( .A(n35249), .B(n35248), .Z(n35250) );
  NAND U51024 ( .A(n35251), .B(n35250), .Z(n35255) );
  AND U51025 ( .A(n35253), .B(n35252), .Z(n35254) );
  NAND U51026 ( .A(n35255), .B(n35254), .Z(n35256) );
  NANDN U51027 ( .A(n54446), .B(n35256), .Z(n35257) );
  OR U51028 ( .A(n35258), .B(n35257), .Z(n35259) );
  AND U51029 ( .A(n35260), .B(n35259), .Z(n35261) );
  NANDN U51030 ( .A(n54447), .B(n35261), .Z(n35262) );
  AND U51031 ( .A(n54448), .B(n35262), .Z(n35265) );
  NANDN U51032 ( .A(x[2282]), .B(y[2282]), .Z(n35264) );
  NAND U51033 ( .A(n35264), .B(n35263), .Z(n54449) );
  OR U51034 ( .A(n35265), .B(n54449), .Z(n35266) );
  NAND U51035 ( .A(n54450), .B(n35266), .Z(n35267) );
  NANDN U51036 ( .A(n52112), .B(n35267), .Z(n35268) );
  AND U51037 ( .A(n35269), .B(n35268), .Z(n35272) );
  NAND U51038 ( .A(n54452), .B(n35270), .Z(n35271) );
  OR U51039 ( .A(n35272), .B(n35271), .Z(n35273) );
  AND U51040 ( .A(n35274), .B(n35273), .Z(n35276) );
  NAND U51041 ( .A(n35276), .B(n35275), .Z(n35277) );
  NANDN U51042 ( .A(n35278), .B(n35277), .Z(n35279) );
  AND U51043 ( .A(n35280), .B(n35279), .Z(n35281) );
  NOR U51044 ( .A(n54458), .B(n35281), .Z(n35282) );
  NANDN U51045 ( .A(n35283), .B(n35282), .Z(n35284) );
  AND U51046 ( .A(n35285), .B(n35284), .Z(n35286) );
  OR U51047 ( .A(n54460), .B(n35286), .Z(n35287) );
  NAND U51048 ( .A(n35288), .B(n35287), .Z(n35289) );
  NANDN U51049 ( .A(n35290), .B(n35289), .Z(n35292) );
  IV U51050 ( .A(n35291), .Z(n54462) );
  OR U51051 ( .A(n35292), .B(n54462), .Z(n35293) );
  AND U51052 ( .A(n35294), .B(n35293), .Z(n35295) );
  NANDN U51053 ( .A(n35296), .B(n35295), .Z(n35297) );
  AND U51054 ( .A(n35298), .B(n35297), .Z(n35300) );
  NOR U51055 ( .A(n35300), .B(n35299), .Z(n35301) );
  NANDN U51056 ( .A(n35302), .B(n35301), .Z(n35303) );
  AND U51057 ( .A(n54468), .B(n35303), .Z(n35305) );
  NAND U51058 ( .A(n35305), .B(n35304), .Z(n35306) );
  NAND U51059 ( .A(n54469), .B(n35306), .Z(n35308) );
  OR U51060 ( .A(n35308), .B(n35307), .Z(n35309) );
  AND U51061 ( .A(n35310), .B(n35309), .Z(n35314) );
  NAND U51062 ( .A(n35312), .B(n35311), .Z(n35313) );
  OR U51063 ( .A(n35314), .B(n35313), .Z(n35315) );
  AND U51064 ( .A(n35316), .B(n35315), .Z(n35318) );
  NOR U51065 ( .A(n35318), .B(n35317), .Z(n35319) );
  NANDN U51066 ( .A(n35320), .B(n35319), .Z(n35321) );
  AND U51067 ( .A(n52106), .B(n35321), .Z(n35323) );
  AND U51068 ( .A(n35323), .B(n35322), .Z(n35327) );
  NAND U51069 ( .A(n35325), .B(n35324), .Z(n35326) );
  OR U51070 ( .A(n35327), .B(n35326), .Z(n35328) );
  AND U51071 ( .A(n35329), .B(n35328), .Z(n35330) );
  NANDN U51072 ( .A(n52105), .B(n35330), .Z(n35331) );
  NAND U51073 ( .A(n35332), .B(n35331), .Z(n35333) );
  NANDN U51074 ( .A(n35334), .B(n35333), .Z(n35336) );
  OR U51075 ( .A(n35336), .B(n35335), .Z(n35337) );
  NAND U51076 ( .A(n35338), .B(n35337), .Z(n35342) );
  AND U51077 ( .A(n35340), .B(n35339), .Z(n35341) );
  NAND U51078 ( .A(n35342), .B(n35341), .Z(n35343) );
  NANDN U51079 ( .A(n54480), .B(n35343), .Z(n35344) );
  OR U51080 ( .A(n35345), .B(n35344), .Z(n35346) );
  AND U51081 ( .A(n35347), .B(n35346), .Z(n35348) );
  NANDN U51082 ( .A(n35349), .B(n35348), .Z(n35350) );
  AND U51083 ( .A(n54483), .B(n35350), .Z(n35351) );
  OR U51084 ( .A(n35352), .B(n35351), .Z(n35353) );
  NAND U51085 ( .A(n54484), .B(n35353), .Z(n35354) );
  NANDN U51086 ( .A(n35355), .B(n35354), .Z(n35356) );
  NANDN U51087 ( .A(n35356), .B(n54485), .Z(n35357) );
  NANDN U51088 ( .A(n54488), .B(n35357), .Z(n35359) );
  IV U51089 ( .A(n35358), .Z(n54489) );
  AND U51090 ( .A(n35359), .B(n54489), .Z(n35360) );
  ANDN U51091 ( .B(n35361), .A(n35360), .Z(n35362) );
  NAND U51092 ( .A(n52104), .B(n35362), .Z(n35363) );
  NANDN U51093 ( .A(n35364), .B(n35363), .Z(n35365) );
  OR U51094 ( .A(n35365), .B(n54490), .Z(n35366) );
  AND U51095 ( .A(n35367), .B(n35366), .Z(n35368) );
  NANDN U51096 ( .A(n35369), .B(n35368), .Z(n35370) );
  AND U51097 ( .A(n35371), .B(n35370), .Z(n35375) );
  NAND U51098 ( .A(n35373), .B(n35372), .Z(n35374) );
  OR U51099 ( .A(n35375), .B(n35374), .Z(n35376) );
  AND U51100 ( .A(n35377), .B(n35376), .Z(n35381) );
  NAND U51101 ( .A(n35379), .B(n35378), .Z(n35380) );
  OR U51102 ( .A(n35381), .B(n35380), .Z(n35382) );
  AND U51103 ( .A(n35383), .B(n35382), .Z(n35384) );
  ANDN U51104 ( .B(n35385), .A(n35384), .Z(n35386) );
  NAND U51105 ( .A(n35387), .B(n35386), .Z(n35388) );
  NANDN U51106 ( .A(n54498), .B(n35388), .Z(n35389) );
  OR U51107 ( .A(n35390), .B(n35389), .Z(n35391) );
  AND U51108 ( .A(n35392), .B(n35391), .Z(n35393) );
  NANDN U51109 ( .A(n54499), .B(n35393), .Z(n35396) );
  NANDN U51110 ( .A(x[2333]), .B(y[2333]), .Z(n35395) );
  AND U51111 ( .A(n35395), .B(n35394), .Z(n54500) );
  AND U51112 ( .A(n35396), .B(n54500), .Z(n35399) );
  NANDN U51113 ( .A(n35399), .B(n54501), .Z(n35400) );
  NAND U51114 ( .A(n52099), .B(n35400), .Z(n35401) );
  NANDN U51115 ( .A(n54502), .B(n35401), .Z(n35402) );
  NAND U51116 ( .A(n54504), .B(n35402), .Z(n35403) );
  ANDN U51117 ( .B(n35403), .A(n54505), .Z(n35404) );
  NANDN U51118 ( .A(n35405), .B(n35404), .Z(n35406) );
  AND U51119 ( .A(n35407), .B(n35406), .Z(n35408) );
  NAND U51120 ( .A(n54506), .B(n35408), .Z(n35412) );
  NAND U51121 ( .A(n35410), .B(n35409), .Z(n35411) );
  ANDN U51122 ( .B(n35412), .A(n35411), .Z(n35416) );
  NAND U51123 ( .A(n35414), .B(n35413), .Z(n35415) );
  OR U51124 ( .A(n35416), .B(n35415), .Z(n35417) );
  AND U51125 ( .A(n35418), .B(n35417), .Z(n35422) );
  NAND U51126 ( .A(n35420), .B(n35419), .Z(n35421) );
  OR U51127 ( .A(n35422), .B(n35421), .Z(n35423) );
  AND U51128 ( .A(n35424), .B(n35423), .Z(n35426) );
  AND U51129 ( .A(n35426), .B(n35425), .Z(n35427) );
  OR U51130 ( .A(n35428), .B(n35427), .Z(n35429) );
  NAND U51131 ( .A(n35430), .B(n35429), .Z(n35431) );
  AND U51132 ( .A(n35432), .B(n35431), .Z(n35433) );
  OR U51133 ( .A(n35434), .B(n35433), .Z(n35435) );
  NAND U51134 ( .A(n35436), .B(n35435), .Z(n35437) );
  NANDN U51135 ( .A(n35438), .B(n35437), .Z(n35442) );
  NANDN U51136 ( .A(x[2350]), .B(y[2350]), .Z(n35439) );
  AND U51137 ( .A(n35440), .B(n35439), .Z(n35441) );
  NAND U51138 ( .A(n35442), .B(n35441), .Z(n35446) );
  NAND U51139 ( .A(n35444), .B(n35443), .Z(n35445) );
  ANDN U51140 ( .B(n35446), .A(n35445), .Z(n35450) );
  NAND U51141 ( .A(n35448), .B(n35447), .Z(n35449) );
  OR U51142 ( .A(n35450), .B(n35449), .Z(n35451) );
  AND U51143 ( .A(n35452), .B(n35451), .Z(n35456) );
  NAND U51144 ( .A(n35454), .B(n35453), .Z(n35455) );
  OR U51145 ( .A(n35456), .B(n35455), .Z(n35457) );
  AND U51146 ( .A(n35458), .B(n35457), .Z(n35459) );
  OR U51147 ( .A(n35460), .B(n35459), .Z(n35461) );
  NAND U51148 ( .A(n35462), .B(n35461), .Z(n35463) );
  AND U51149 ( .A(n35464), .B(n35463), .Z(n35465) );
  OR U51150 ( .A(n54524), .B(n35465), .Z(n35466) );
  NAND U51151 ( .A(n54525), .B(n35466), .Z(n35467) );
  NANDN U51152 ( .A(n54526), .B(n35467), .Z(n35468) );
  NAND U51153 ( .A(n54527), .B(n35468), .Z(n35469) );
  NANDN U51154 ( .A(n54528), .B(n35469), .Z(n35470) );
  AND U51155 ( .A(n54529), .B(n35470), .Z(n35471) );
  OR U51156 ( .A(n35472), .B(n35471), .Z(n35473) );
  NAND U51157 ( .A(n35474), .B(n35473), .Z(n35478) );
  NAND U51158 ( .A(n35476), .B(n35475), .Z(n35477) );
  ANDN U51159 ( .B(n35478), .A(n35477), .Z(n35482) );
  NAND U51160 ( .A(n35480), .B(n35479), .Z(n35481) );
  OR U51161 ( .A(n35482), .B(n35481), .Z(n35483) );
  AND U51162 ( .A(n35484), .B(n35483), .Z(n35488) );
  NAND U51163 ( .A(n35486), .B(n35485), .Z(n35487) );
  OR U51164 ( .A(n35488), .B(n35487), .Z(n35489) );
  AND U51165 ( .A(n35490), .B(n35489), .Z(n35494) );
  NAND U51166 ( .A(n35492), .B(n35491), .Z(n35493) );
  OR U51167 ( .A(n35494), .B(n35493), .Z(n35495) );
  AND U51168 ( .A(n35496), .B(n35495), .Z(n35500) );
  NAND U51169 ( .A(n35498), .B(n35497), .Z(n35499) );
  OR U51170 ( .A(n35500), .B(n35499), .Z(n35501) );
  AND U51171 ( .A(n35502), .B(n35501), .Z(n35506) );
  NAND U51172 ( .A(n35504), .B(n35503), .Z(n35505) );
  OR U51173 ( .A(n35506), .B(n35505), .Z(n35507) );
  AND U51174 ( .A(n35508), .B(n35507), .Z(n35512) );
  NAND U51175 ( .A(n35510), .B(n35509), .Z(n35511) );
  OR U51176 ( .A(n35512), .B(n35511), .Z(n35513) );
  AND U51177 ( .A(n35514), .B(n35513), .Z(n35516) );
  NOR U51178 ( .A(n35516), .B(n35515), .Z(n35517) );
  NANDN U51179 ( .A(n35518), .B(n35517), .Z(n35519) );
  AND U51180 ( .A(n35520), .B(n35519), .Z(n35521) );
  NANDN U51181 ( .A(n35522), .B(n35521), .Z(n35523) );
  AND U51182 ( .A(n35524), .B(n35523), .Z(n35526) );
  NANDN U51183 ( .A(x[2382]), .B(y[2382]), .Z(n35525) );
  NAND U51184 ( .A(n35526), .B(n35525), .Z(n35528) );
  ANDN U51185 ( .B(n35528), .A(n35527), .Z(n35529) );
  NANDN U51186 ( .A(n54547), .B(n35529), .Z(n35530) );
  AND U51187 ( .A(n35531), .B(n35530), .Z(n35534) );
  NANDN U51188 ( .A(n35534), .B(n54551), .Z(n35535) );
  NANDN U51189 ( .A(n54552), .B(n35535), .Z(n35536) );
  AND U51190 ( .A(n54553), .B(n35536), .Z(n35539) );
  NANDN U51191 ( .A(x[2389]), .B(y[2389]), .Z(n35538) );
  NAND U51192 ( .A(n35538), .B(n35537), .Z(n52090) );
  OR U51193 ( .A(n35539), .B(n52090), .Z(n35540) );
  AND U51194 ( .A(n54554), .B(n35540), .Z(n35541) );
  OR U51195 ( .A(n35541), .B(n54555), .Z(n35543) );
  IV U51196 ( .A(n35542), .Z(n54556) );
  AND U51197 ( .A(n35543), .B(n54556), .Z(n35545) );
  IV U51198 ( .A(n35544), .Z(n54557) );
  OR U51199 ( .A(n35545), .B(n54557), .Z(n35546) );
  AND U51200 ( .A(n54558), .B(n35546), .Z(n35549) );
  NAND U51201 ( .A(n35548), .B(n35547), .Z(n54559) );
  OR U51202 ( .A(n35549), .B(n54559), .Z(n35550) );
  NAND U51203 ( .A(n35551), .B(n35550), .Z(n35552) );
  NANDN U51204 ( .A(n35553), .B(n35552), .Z(n35554) );
  OR U51205 ( .A(n54561), .B(n35554), .Z(n35555) );
  AND U51206 ( .A(n35556), .B(n35555), .Z(n35558) );
  NAND U51207 ( .A(n35558), .B(n35557), .Z(n35560) );
  ANDN U51208 ( .B(n35560), .A(n35559), .Z(n35561) );
  NANDN U51209 ( .A(n35562), .B(n35561), .Z(n35566) );
  AND U51210 ( .A(n35564), .B(n35563), .Z(n35565) );
  NAND U51211 ( .A(n35566), .B(n35565), .Z(n35567) );
  NANDN U51212 ( .A(n35568), .B(n35567), .Z(n35570) );
  IV U51213 ( .A(n35569), .Z(n54569) );
  OR U51214 ( .A(n35570), .B(n54569), .Z(n35571) );
  AND U51215 ( .A(n35572), .B(n35571), .Z(n35573) );
  NANDN U51216 ( .A(n54570), .B(n35573), .Z(n35576) );
  AND U51217 ( .A(n35575), .B(n35574), .Z(n54571) );
  AND U51218 ( .A(n35576), .B(n54571), .Z(n35579) );
  NANDN U51219 ( .A(n35579), .B(n54572), .Z(n35580) );
  NAND U51220 ( .A(n54573), .B(n35580), .Z(n35581) );
  NAND U51221 ( .A(n54574), .B(n35581), .Z(n35582) );
  NAND U51222 ( .A(n54575), .B(n35582), .Z(n35583) );
  ANDN U51223 ( .B(n35583), .A(n54576), .Z(n35584) );
  NANDN U51224 ( .A(n35585), .B(n35584), .Z(n35588) );
  AND U51225 ( .A(n35586), .B(n52089), .Z(n35587) );
  NAND U51226 ( .A(n35588), .B(n35587), .Z(n35589) );
  NANDN U51227 ( .A(n35590), .B(n35589), .Z(n35592) );
  OR U51228 ( .A(n35592), .B(n35591), .Z(n35593) );
  NAND U51229 ( .A(n35594), .B(n35593), .Z(n35595) );
  NANDN U51230 ( .A(n35596), .B(n35595), .Z(n35598) );
  OR U51231 ( .A(n35598), .B(n35597), .Z(n35599) );
  NAND U51232 ( .A(n35600), .B(n35599), .Z(n35601) );
  AND U51233 ( .A(n35602), .B(n35601), .Z(n35606) );
  NANDN U51234 ( .A(n35606), .B(n54584), .Z(n35607) );
  NAND U51235 ( .A(n54585), .B(n35607), .Z(n35608) );
  NANDN U51236 ( .A(n54586), .B(n35608), .Z(n35609) );
  NAND U51237 ( .A(n54587), .B(n35609), .Z(n35610) );
  NAND U51238 ( .A(n54588), .B(n35610), .Z(n35611) );
  NANDN U51239 ( .A(n54589), .B(n35611), .Z(n35613) );
  IV U51240 ( .A(n35612), .Z(n54590) );
  AND U51241 ( .A(n35613), .B(n54590), .Z(n35615) );
  IV U51242 ( .A(n35614), .Z(n54591) );
  OR U51243 ( .A(n35615), .B(n54591), .Z(n35616) );
  NAND U51244 ( .A(n35617), .B(n35616), .Z(n35618) );
  NANDN U51245 ( .A(n35619), .B(n35618), .Z(n35620) );
  AND U51246 ( .A(n35621), .B(n35620), .Z(n35622) );
  NAND U51247 ( .A(n35623), .B(n35622), .Z(n35624) );
  NANDN U51248 ( .A(n35625), .B(n35624), .Z(n35626) );
  OR U51249 ( .A(n35627), .B(n35626), .Z(n35628) );
  AND U51250 ( .A(n54595), .B(n35628), .Z(n35630) );
  NANDN U51251 ( .A(x[2426]), .B(y[2426]), .Z(n35629) );
  NAND U51252 ( .A(n35630), .B(n35629), .Z(n35632) );
  ANDN U51253 ( .B(n35632), .A(n35631), .Z(n35633) );
  NANDN U51254 ( .A(n35634), .B(n35633), .Z(n35636) );
  AND U51255 ( .A(n35636), .B(n35635), .Z(n35637) );
  NANDN U51256 ( .A(x[2428]), .B(y[2428]), .Z(n54596) );
  AND U51257 ( .A(n35637), .B(n54596), .Z(n35638) );
  NOR U51258 ( .A(n35639), .B(n35638), .Z(n35641) );
  NAND U51259 ( .A(n35641), .B(n35640), .Z(n35643) );
  AND U51260 ( .A(n35643), .B(n35642), .Z(n35644) );
  NANDN U51261 ( .A(n35645), .B(n35644), .Z(n35646) );
  NAND U51262 ( .A(n35647), .B(n35646), .Z(n35651) );
  AND U51263 ( .A(n35649), .B(n35648), .Z(n35650) );
  NAND U51264 ( .A(n35651), .B(n35650), .Z(n35652) );
  NANDN U51265 ( .A(n54605), .B(n35652), .Z(n35653) );
  OR U51266 ( .A(n35654), .B(n35653), .Z(n35655) );
  AND U51267 ( .A(n35656), .B(n35655), .Z(n35657) );
  NANDN U51268 ( .A(n54606), .B(n35657), .Z(n35658) );
  AND U51269 ( .A(n54607), .B(n35658), .Z(n35659) );
  OR U51270 ( .A(n54608), .B(n35659), .Z(n35660) );
  NAND U51271 ( .A(n35661), .B(n35660), .Z(n35662) );
  NANDN U51272 ( .A(n35663), .B(n35662), .Z(n35664) );
  OR U51273 ( .A(n35664), .B(n54610), .Z(n35665) );
  AND U51274 ( .A(n35666), .B(n35665), .Z(n35668) );
  NOR U51275 ( .A(n35668), .B(n35667), .Z(n35669) );
  NANDN U51276 ( .A(n35670), .B(n35669), .Z(n35671) );
  AND U51277 ( .A(n35672), .B(n35671), .Z(n35674) );
  NAND U51278 ( .A(n35674), .B(n35673), .Z(n35675) );
  NAND U51279 ( .A(n35676), .B(n35675), .Z(n35677) );
  AND U51280 ( .A(n35678), .B(n35677), .Z(n35679) );
  OR U51281 ( .A(n35680), .B(n35679), .Z(n35681) );
  NAND U51282 ( .A(n35682), .B(n35681), .Z(n35686) );
  NANDN U51283 ( .A(x[2446]), .B(y[2446]), .Z(n35684) );
  IV U51284 ( .A(n35683), .Z(n54620) );
  AND U51285 ( .A(n35684), .B(n54620), .Z(n35685) );
  NAND U51286 ( .A(n35686), .B(n35685), .Z(n35687) );
  NANDN U51287 ( .A(n35688), .B(n35687), .Z(n35689) );
  OR U51288 ( .A(n35690), .B(n35689), .Z(n35691) );
  AND U51289 ( .A(n35692), .B(n35691), .Z(n35693) );
  NANDN U51290 ( .A(x[2448]), .B(y[2448]), .Z(n54621) );
  NAND U51291 ( .A(n35693), .B(n54621), .Z(n35695) );
  ANDN U51292 ( .B(n35695), .A(n35694), .Z(n35696) );
  NANDN U51293 ( .A(n35697), .B(n35696), .Z(n35701) );
  NANDN U51294 ( .A(x[2450]), .B(y[2450]), .Z(n35698) );
  AND U51295 ( .A(n35699), .B(n35698), .Z(n35700) );
  NAND U51296 ( .A(n35701), .B(n35700), .Z(n35702) );
  NANDN U51297 ( .A(n35703), .B(n35702), .Z(n35706) );
  AND U51298 ( .A(n35704), .B(n54625), .Z(n35705) );
  NAND U51299 ( .A(n35706), .B(n35705), .Z(n35707) );
  NANDN U51300 ( .A(n35708), .B(n35707), .Z(n35709) );
  OR U51301 ( .A(n54626), .B(n35709), .Z(n35710) );
  AND U51302 ( .A(n54627), .B(n35710), .Z(n35713) );
  NAND U51303 ( .A(n35712), .B(n35711), .Z(n52081) );
  OR U51304 ( .A(n35713), .B(n52081), .Z(n35714) );
  NAND U51305 ( .A(n54629), .B(n35714), .Z(n35715) );
  NANDN U51306 ( .A(n54630), .B(n35715), .Z(n35716) );
  NAND U51307 ( .A(n54631), .B(n35716), .Z(n35717) );
  AND U51308 ( .A(n35718), .B(n35717), .Z(n35719) );
  OR U51309 ( .A(n35720), .B(n35719), .Z(n35721) );
  NAND U51310 ( .A(n35722), .B(n35721), .Z(n35723) );
  NANDN U51311 ( .A(n35724), .B(n35723), .Z(n35728) );
  NOR U51312 ( .A(n35726), .B(n35725), .Z(n35727) );
  NAND U51313 ( .A(n35728), .B(n35727), .Z(n35729) );
  AND U51314 ( .A(n35730), .B(n35729), .Z(n35733) );
  NANDN U51315 ( .A(y[2465]), .B(n35733), .Z(n35732) );
  ANDN U51316 ( .B(n35732), .A(n35731), .Z(n35736) );
  XNOR U51317 ( .A(n35733), .B(y[2465]), .Z(n35734) );
  NAND U51318 ( .A(n35734), .B(x[2465]), .Z(n35735) );
  NAND U51319 ( .A(n35736), .B(n35735), .Z(n35740) );
  NANDN U51320 ( .A(x[2466]), .B(y[2466]), .Z(n35737) );
  AND U51321 ( .A(n35738), .B(n35737), .Z(n35739) );
  NAND U51322 ( .A(n35740), .B(n35739), .Z(n35744) );
  NAND U51323 ( .A(n35742), .B(n35741), .Z(n35743) );
  ANDN U51324 ( .B(n35744), .A(n35743), .Z(n35745) );
  OR U51325 ( .A(n35746), .B(n35745), .Z(n35747) );
  NAND U51326 ( .A(n35748), .B(n35747), .Z(n35752) );
  NANDN U51327 ( .A(x[2470]), .B(y[2470]), .Z(n35749) );
  AND U51328 ( .A(n35750), .B(n35749), .Z(n35751) );
  NAND U51329 ( .A(n35752), .B(n35751), .Z(n35756) );
  NAND U51330 ( .A(n35754), .B(n35753), .Z(n35755) );
  ANDN U51331 ( .B(n35756), .A(n35755), .Z(n35757) );
  OR U51332 ( .A(n35758), .B(n35757), .Z(n35759) );
  NAND U51333 ( .A(n35760), .B(n35759), .Z(n35761) );
  AND U51334 ( .A(n54650), .B(n35761), .Z(n35762) );
  NAND U51335 ( .A(n35763), .B(n35762), .Z(n35764) );
  NANDN U51336 ( .A(n54651), .B(n35764), .Z(n35766) );
  OR U51337 ( .A(n35766), .B(n35765), .Z(n35767) );
  NAND U51338 ( .A(n35768), .B(n35767), .Z(n35769) );
  NANDN U51339 ( .A(n35770), .B(n35769), .Z(n35774) );
  IV U51340 ( .A(n35771), .Z(n52076) );
  AND U51341 ( .A(n35772), .B(n52076), .Z(n35773) );
  NAND U51342 ( .A(n35774), .B(n35773), .Z(n35775) );
  NANDN U51343 ( .A(n35776), .B(n35775), .Z(n35778) );
  OR U51344 ( .A(n35778), .B(n35777), .Z(n35779) );
  NAND U51345 ( .A(n35780), .B(n35779), .Z(n35781) );
  NANDN U51346 ( .A(n35782), .B(n35781), .Z(n35784) );
  OR U51347 ( .A(n35784), .B(n35783), .Z(n35785) );
  NAND U51348 ( .A(n35786), .B(n35785), .Z(n35787) );
  NAND U51349 ( .A(n35788), .B(n35787), .Z(n35790) );
  ANDN U51350 ( .B(y[2484]), .A(x[2484]), .Z(n35789) );
  ANDN U51351 ( .B(n35790), .A(n35789), .Z(n35792) );
  ANDN U51352 ( .B(n35792), .A(n35791), .Z(n35793) );
  OR U51353 ( .A(n35794), .B(n35793), .Z(n35795) );
  NAND U51354 ( .A(n35796), .B(n35795), .Z(n35800) );
  AND U51355 ( .A(n35798), .B(n35797), .Z(n35799) );
  NAND U51356 ( .A(n35800), .B(n35799), .Z(n35801) );
  NANDN U51357 ( .A(n35802), .B(n35801), .Z(n35804) );
  ANDN U51358 ( .B(y[2488]), .A(x[2488]), .Z(n35803) );
  OR U51359 ( .A(n35804), .B(n35803), .Z(n35805) );
  NAND U51360 ( .A(n35806), .B(n35805), .Z(n35807) );
  NANDN U51361 ( .A(n35808), .B(n35807), .Z(n35809) );
  OR U51362 ( .A(n35810), .B(n35809), .Z(n35811) );
  AND U51363 ( .A(n35812), .B(n35811), .Z(n35813) );
  NANDN U51364 ( .A(n35814), .B(n35813), .Z(n35815) );
  AND U51365 ( .A(n35816), .B(n35815), .Z(n35817) );
  NOR U51366 ( .A(n35818), .B(n35817), .Z(n35819) );
  NANDN U51367 ( .A(n35820), .B(n35819), .Z(n35821) );
  AND U51368 ( .A(n35822), .B(n35821), .Z(n35824) );
  NANDN U51369 ( .A(x[2494]), .B(y[2494]), .Z(n35823) );
  NAND U51370 ( .A(n35824), .B(n35823), .Z(n35825) );
  NAND U51371 ( .A(n35826), .B(n35825), .Z(n35828) );
  OR U51372 ( .A(n35828), .B(n35827), .Z(n35829) );
  AND U51373 ( .A(n35830), .B(n35829), .Z(n35834) );
  NAND U51374 ( .A(n35832), .B(n35831), .Z(n35833) );
  OR U51375 ( .A(n35834), .B(n35833), .Z(n35835) );
  AND U51376 ( .A(n35836), .B(n35835), .Z(n35840) );
  NAND U51377 ( .A(n35838), .B(n35837), .Z(n35839) );
  OR U51378 ( .A(n35840), .B(n35839), .Z(n35841) );
  AND U51379 ( .A(n35842), .B(n35841), .Z(n35843) );
  NANDN U51380 ( .A(n35844), .B(n35843), .Z(n35845) );
  NAND U51381 ( .A(n35846), .B(n35845), .Z(n35847) );
  NANDN U51382 ( .A(n35848), .B(n35847), .Z(n35850) );
  ANDN U51383 ( .B(y[2502]), .A(x[2502]), .Z(n35849) );
  OR U51384 ( .A(n35850), .B(n35849), .Z(n35851) );
  NAND U51385 ( .A(n35852), .B(n35851), .Z(n35853) );
  NANDN U51386 ( .A(n35854), .B(n35853), .Z(n35856) );
  ANDN U51387 ( .B(y[2504]), .A(x[2504]), .Z(n35855) );
  OR U51388 ( .A(n35856), .B(n35855), .Z(n35857) );
  NAND U51389 ( .A(n35858), .B(n35857), .Z(n35862) );
  AND U51390 ( .A(n35860), .B(n35859), .Z(n35861) );
  NAND U51391 ( .A(n35862), .B(n35861), .Z(n35863) );
  NANDN U51392 ( .A(n35864), .B(n35863), .Z(n35866) );
  OR U51393 ( .A(n35866), .B(n35865), .Z(n35867) );
  NAND U51394 ( .A(n35868), .B(n35867), .Z(n35869) );
  NANDN U51395 ( .A(n35870), .B(n35869), .Z(n35872) );
  OR U51396 ( .A(n35872), .B(n35871), .Z(n35873) );
  NAND U51397 ( .A(n35874), .B(n35873), .Z(n35875) );
  NAND U51398 ( .A(n35876), .B(n35875), .Z(n35877) );
  NAND U51399 ( .A(n54685), .B(n35877), .Z(n35878) );
  AND U51400 ( .A(n54686), .B(n35878), .Z(n35881) );
  NANDN U51401 ( .A(n35881), .B(n54688), .Z(n35882) );
  NAND U51402 ( .A(n54689), .B(n35882), .Z(n35883) );
  NAND U51403 ( .A(n54690), .B(n35883), .Z(n35886) );
  AND U51404 ( .A(n35884), .B(n54691), .Z(n35885) );
  NAND U51405 ( .A(n35886), .B(n35885), .Z(n35887) );
  NANDN U51406 ( .A(n35888), .B(n35887), .Z(n35889) );
  OR U51407 ( .A(n35889), .B(n54692), .Z(n35890) );
  NAND U51408 ( .A(n35891), .B(n35890), .Z(n35895) );
  NANDN U51409 ( .A(x[2520]), .B(y[2520]), .Z(n35892) );
  AND U51410 ( .A(n35893), .B(n35892), .Z(n35894) );
  NAND U51411 ( .A(n35895), .B(n35894), .Z(n35896) );
  NANDN U51412 ( .A(n35897), .B(n35896), .Z(n35901) );
  AND U51413 ( .A(n35899), .B(n35898), .Z(n35900) );
  NAND U51414 ( .A(n35901), .B(n35900), .Z(n35902) );
  NANDN U51415 ( .A(n35903), .B(n35902), .Z(n35904) );
  OR U51416 ( .A(n35905), .B(n35904), .Z(n35906) );
  AND U51417 ( .A(n35907), .B(n35906), .Z(n35909) );
  NAND U51418 ( .A(n35909), .B(n35908), .Z(n35911) );
  ANDN U51419 ( .B(n35911), .A(n35910), .Z(n35912) );
  NANDN U51420 ( .A(n35913), .B(n35912), .Z(n35916) );
  AND U51421 ( .A(n35914), .B(n52067), .Z(n35915) );
  NAND U51422 ( .A(n35916), .B(n35915), .Z(n35917) );
  NANDN U51423 ( .A(n35918), .B(n35917), .Z(n35919) );
  OR U51424 ( .A(n35919), .B(n52066), .Z(n35920) );
  NAND U51425 ( .A(n52065), .B(n35920), .Z(n35921) );
  NANDN U51426 ( .A(n35922), .B(n35921), .Z(n35925) );
  AND U51427 ( .A(n35923), .B(n54702), .Z(n35924) );
  NAND U51428 ( .A(n35925), .B(n35924), .Z(n35926) );
  NANDN U51429 ( .A(n35927), .B(n35926), .Z(n35929) );
  OR U51430 ( .A(n35929), .B(n35928), .Z(n35930) );
  NAND U51431 ( .A(n35931), .B(n35930), .Z(n35932) );
  NANDN U51432 ( .A(n35933), .B(n35932), .Z(n35935) );
  OR U51433 ( .A(n35935), .B(n35934), .Z(n35936) );
  AND U51434 ( .A(n35937), .B(n35936), .Z(n35938) );
  OR U51435 ( .A(n35939), .B(n35938), .Z(n35940) );
  NAND U51436 ( .A(n52062), .B(n35940), .Z(n35941) );
  NANDN U51437 ( .A(n52061), .B(n35941), .Z(n35942) );
  NANDN U51438 ( .A(n35942), .B(n52063), .Z(n35943) );
  NAND U51439 ( .A(n35944), .B(n35943), .Z(n35948) );
  AND U51440 ( .A(n35946), .B(n35945), .Z(n35947) );
  NAND U51441 ( .A(n35948), .B(n35947), .Z(n35949) );
  NANDN U51442 ( .A(n35950), .B(n35949), .Z(n35952) );
  ANDN U51443 ( .B(y[2540]), .A(x[2540]), .Z(n35951) );
  OR U51444 ( .A(n35952), .B(n35951), .Z(n35953) );
  NAND U51445 ( .A(n35954), .B(n35953), .Z(n35955) );
  NANDN U51446 ( .A(n35956), .B(n35955), .Z(n35958) );
  ANDN U51447 ( .B(y[2542]), .A(x[2542]), .Z(n35957) );
  OR U51448 ( .A(n35958), .B(n35957), .Z(n35959) );
  NAND U51449 ( .A(n35960), .B(n35959), .Z(n35961) );
  AND U51450 ( .A(n35962), .B(n35961), .Z(n35963) );
  NAND U51451 ( .A(n35964), .B(n35963), .Z(n35965) );
  NANDN U51452 ( .A(n35966), .B(n35965), .Z(n35967) );
  OR U51453 ( .A(n35968), .B(n35967), .Z(n35969) );
  AND U51454 ( .A(n35970), .B(n35969), .Z(n35972) );
  NANDN U51455 ( .A(x[2546]), .B(y[2546]), .Z(n35971) );
  AND U51456 ( .A(n35972), .B(n35971), .Z(n35976) );
  NAND U51457 ( .A(n35974), .B(n35973), .Z(n35975) );
  OR U51458 ( .A(n35976), .B(n35975), .Z(n35977) );
  AND U51459 ( .A(n52058), .B(n35977), .Z(n35979) );
  NANDN U51460 ( .A(x[2548]), .B(y[2548]), .Z(n35978) );
  NAND U51461 ( .A(n35979), .B(n35978), .Z(n35981) );
  ANDN U51462 ( .B(n35981), .A(n35980), .Z(n35982) );
  NANDN U51463 ( .A(n35983), .B(n35982), .Z(n35985) );
  AND U51464 ( .A(n35985), .B(n35984), .Z(n35986) );
  NANDN U51465 ( .A(x[2550]), .B(y[2550]), .Z(n52059) );
  AND U51466 ( .A(n35986), .B(n52059), .Z(n35987) );
  OR U51467 ( .A(n35988), .B(n35987), .Z(n35989) );
  AND U51468 ( .A(n35990), .B(n35989), .Z(n35991) );
  NOR U51469 ( .A(n35992), .B(n35991), .Z(n35993) );
  NANDN U51470 ( .A(n35994), .B(n35993), .Z(n35995) );
  AND U51471 ( .A(n35996), .B(n35995), .Z(n35998) );
  NANDN U51472 ( .A(x[2554]), .B(y[2554]), .Z(n35997) );
  NAND U51473 ( .A(n35998), .B(n35997), .Z(n35999) );
  NAND U51474 ( .A(n36000), .B(n35999), .Z(n36002) );
  OR U51475 ( .A(n36002), .B(n36001), .Z(n36003) );
  AND U51476 ( .A(n36004), .B(n36003), .Z(n36007) );
  NANDN U51477 ( .A(n36007), .B(n54729), .Z(n36008) );
  NAND U51478 ( .A(n36009), .B(n36008), .Z(n36010) );
  NANDN U51479 ( .A(n36011), .B(n36010), .Z(n36012) );
  OR U51480 ( .A(n54731), .B(n36012), .Z(n36013) );
  AND U51481 ( .A(n36014), .B(n36013), .Z(n36016) );
  NAND U51482 ( .A(n36016), .B(n36015), .Z(n36018) );
  ANDN U51483 ( .B(n36018), .A(n36017), .Z(n36019) );
  NANDN U51484 ( .A(n36020), .B(n36019), .Z(n36023) );
  AND U51485 ( .A(n36021), .B(n52057), .Z(n36022) );
  NAND U51486 ( .A(n36023), .B(n36022), .Z(n36024) );
  NANDN U51487 ( .A(n54737), .B(n36024), .Z(n36026) );
  OR U51488 ( .A(n36026), .B(n36025), .Z(n36027) );
  NAND U51489 ( .A(n54738), .B(n36027), .Z(n36028) );
  NANDN U51490 ( .A(n36029), .B(n36028), .Z(n36032) );
  AND U51491 ( .A(n36030), .B(n54740), .Z(n36031) );
  NAND U51492 ( .A(n36032), .B(n36031), .Z(n36033) );
  NANDN U51493 ( .A(n36034), .B(n36033), .Z(n36036) );
  OR U51494 ( .A(n36036), .B(n36035), .Z(n36037) );
  NAND U51495 ( .A(n36038), .B(n36037), .Z(n36039) );
  NANDN U51496 ( .A(n36040), .B(n36039), .Z(n36042) );
  OR U51497 ( .A(n36042), .B(n36041), .Z(n36043) );
  AND U51498 ( .A(n36044), .B(n36043), .Z(n36045) );
  OR U51499 ( .A(n36046), .B(n36045), .Z(n36047) );
  NAND U51500 ( .A(n36048), .B(n36047), .Z(n36052) );
  AND U51501 ( .A(n36050), .B(n36049), .Z(n36051) );
  NAND U51502 ( .A(n36052), .B(n36051), .Z(n36053) );
  NANDN U51503 ( .A(n36054), .B(n36053), .Z(n36055) );
  OR U51504 ( .A(n54748), .B(n36055), .Z(n36056) );
  AND U51505 ( .A(n36057), .B(n36056), .Z(n36058) );
  NANDN U51506 ( .A(n54750), .B(n36058), .Z(n36059) );
  AND U51507 ( .A(n54751), .B(n36059), .Z(n36060) );
  OR U51508 ( .A(n54752), .B(n36060), .Z(n36061) );
  NAND U51509 ( .A(n54753), .B(n36061), .Z(n36062) );
  NANDN U51510 ( .A(n54754), .B(n36062), .Z(n36063) );
  NAND U51511 ( .A(n54755), .B(n36063), .Z(n36065) );
  IV U51512 ( .A(n36064), .Z(n54756) );
  ANDN U51513 ( .B(n36065), .A(n54756), .Z(n36066) );
  NANDN U51514 ( .A(n36067), .B(n36066), .Z(n36070) );
  AND U51515 ( .A(n36068), .B(n54757), .Z(n36069) );
  NAND U51516 ( .A(n36070), .B(n36069), .Z(n36071) );
  NANDN U51517 ( .A(n36072), .B(n36071), .Z(n36073) );
  OR U51518 ( .A(n36074), .B(n36073), .Z(n36075) );
  AND U51519 ( .A(n36076), .B(n36075), .Z(n36079) );
  NANDN U51520 ( .A(y[2585]), .B(n36079), .Z(n36078) );
  ANDN U51521 ( .B(n36078), .A(n36077), .Z(n36082) );
  XNOR U51522 ( .A(n36079), .B(y[2585]), .Z(n36080) );
  NAND U51523 ( .A(n36080), .B(x[2585]), .Z(n36081) );
  NAND U51524 ( .A(n36082), .B(n36081), .Z(n36083) );
  AND U51525 ( .A(n36084), .B(n36083), .Z(n36085) );
  NAND U51526 ( .A(n36086), .B(n36085), .Z(n36087) );
  NANDN U51527 ( .A(n36088), .B(n36087), .Z(n36090) );
  OR U51528 ( .A(n36090), .B(n36089), .Z(n36091) );
  NAND U51529 ( .A(n36092), .B(n36091), .Z(n36093) );
  NANDN U51530 ( .A(n36094), .B(n36093), .Z(n36096) );
  NANDN U51531 ( .A(n36096), .B(n36095), .Z(n36097) );
  NAND U51532 ( .A(n36098), .B(n36097), .Z(n36099) );
  NAND U51533 ( .A(n36100), .B(n36099), .Z(n36101) );
  AND U51534 ( .A(n36102), .B(n36101), .Z(n36103) );
  NAND U51535 ( .A(n36104), .B(n36103), .Z(n36105) );
  NANDN U51536 ( .A(n36106), .B(n36105), .Z(n36107) );
  OR U51537 ( .A(n36108), .B(n36107), .Z(n36109) );
  NAND U51538 ( .A(n36110), .B(n36109), .Z(n36111) );
  NANDN U51539 ( .A(n36112), .B(n36111), .Z(n36113) );
  NANDN U51540 ( .A(y[2596]), .B(n36113), .Z(n36116) );
  XNOR U51541 ( .A(y[2596]), .B(n36113), .Z(n36114) );
  NAND U51542 ( .A(n36114), .B(x[2596]), .Z(n36115) );
  NAND U51543 ( .A(n36116), .B(n36115), .Z(n36117) );
  AND U51544 ( .A(n36118), .B(n36117), .Z(n36122) );
  NAND U51545 ( .A(n36120), .B(n36119), .Z(n36121) );
  OR U51546 ( .A(n36122), .B(n36121), .Z(n36123) );
  AND U51547 ( .A(n36124), .B(n36123), .Z(n36128) );
  NAND U51548 ( .A(n36126), .B(n36125), .Z(n36127) );
  OR U51549 ( .A(n36128), .B(n36127), .Z(n36129) );
  AND U51550 ( .A(n36130), .B(n36129), .Z(n36134) );
  NAND U51551 ( .A(n36132), .B(n36131), .Z(n36133) );
  OR U51552 ( .A(n36134), .B(n36133), .Z(n36135) );
  AND U51553 ( .A(n36136), .B(n36135), .Z(n36140) );
  NAND U51554 ( .A(n36138), .B(n36137), .Z(n36139) );
  OR U51555 ( .A(n36140), .B(n36139), .Z(n36141) );
  AND U51556 ( .A(n36142), .B(n36141), .Z(n36144) );
  NOR U51557 ( .A(n36144), .B(n36143), .Z(n36145) );
  NANDN U51558 ( .A(n36146), .B(n36145), .Z(n36147) );
  AND U51559 ( .A(n36148), .B(n36147), .Z(n36150) );
  NANDN U51560 ( .A(x[2606]), .B(y[2606]), .Z(n36149) );
  NAND U51561 ( .A(n36150), .B(n36149), .Z(n36151) );
  NAND U51562 ( .A(n36152), .B(n36151), .Z(n36154) );
  OR U51563 ( .A(n36154), .B(n36153), .Z(n36155) );
  AND U51564 ( .A(n36156), .B(n36155), .Z(n36160) );
  NAND U51565 ( .A(n36158), .B(n36157), .Z(n36159) );
  OR U51566 ( .A(n36160), .B(n36159), .Z(n36161) );
  AND U51567 ( .A(n36162), .B(n36161), .Z(n36166) );
  NAND U51568 ( .A(n36164), .B(n36163), .Z(n36165) );
  OR U51569 ( .A(n36166), .B(n36165), .Z(n36167) );
  AND U51570 ( .A(n36168), .B(n36167), .Z(n36169) );
  NOR U51571 ( .A(n36170), .B(n36169), .Z(n36171) );
  NANDN U51572 ( .A(n36172), .B(n36171), .Z(n36173) );
  AND U51573 ( .A(n36173), .B(n54790), .Z(n36175) );
  NANDN U51574 ( .A(x[2614]), .B(y[2614]), .Z(n36174) );
  NAND U51575 ( .A(n36175), .B(n36174), .Z(n36176) );
  NAND U51576 ( .A(n36177), .B(n36176), .Z(n36179) );
  OR U51577 ( .A(n36179), .B(n36178), .Z(n36180) );
  AND U51578 ( .A(n36181), .B(n36180), .Z(n36182) );
  ANDN U51579 ( .B(n36183), .A(n36182), .Z(n36184) );
  NAND U51580 ( .A(n36185), .B(n36184), .Z(n36186) );
  NANDN U51581 ( .A(n52050), .B(n36186), .Z(n36188) );
  OR U51582 ( .A(n36188), .B(n36187), .Z(n36189) );
  NAND U51583 ( .A(n36190), .B(n36189), .Z(n36191) );
  NANDN U51584 ( .A(n36192), .B(n36191), .Z(n36194) );
  OR U51585 ( .A(n36194), .B(n36193), .Z(n36195) );
  AND U51586 ( .A(n36196), .B(n36195), .Z(n36197) );
  OR U51587 ( .A(n36198), .B(n36197), .Z(n36199) );
  NAND U51588 ( .A(n36200), .B(n36199), .Z(n36201) );
  NANDN U51589 ( .A(n36202), .B(n36201), .Z(n36206) );
  AND U51590 ( .A(n36204), .B(n36203), .Z(n36205) );
  NAND U51591 ( .A(n36206), .B(n36205), .Z(n36207) );
  NANDN U51592 ( .A(n36208), .B(n36207), .Z(n36210) );
  OR U51593 ( .A(n36210), .B(n36209), .Z(n36211) );
  NAND U51594 ( .A(n36212), .B(n36211), .Z(n36213) );
  NANDN U51595 ( .A(n52048), .B(n36213), .Z(n36215) );
  OR U51596 ( .A(n36215), .B(n36214), .Z(n36216) );
  NAND U51597 ( .A(n36217), .B(n36216), .Z(n36219) );
  NANDN U51598 ( .A(x[2630]), .B(y[2630]), .Z(n52049) );
  AND U51599 ( .A(n54806), .B(n52049), .Z(n36218) );
  NAND U51600 ( .A(n36219), .B(n36218), .Z(n36220) );
  NANDN U51601 ( .A(n36221), .B(n36220), .Z(n36222) );
  OR U51602 ( .A(n36223), .B(n36222), .Z(n36224) );
  AND U51603 ( .A(n36225), .B(n36224), .Z(n36226) );
  NAND U51604 ( .A(n52047), .B(n36226), .Z(n36228) );
  ANDN U51605 ( .B(n36228), .A(n36227), .Z(n36229) );
  NANDN U51606 ( .A(n36230), .B(n36229), .Z(n36231) );
  NAND U51607 ( .A(n36232), .B(n36231), .Z(n36233) );
  NANDN U51608 ( .A(n36234), .B(n36233), .Z(n36235) );
  AND U51609 ( .A(n36236), .B(n36235), .Z(n36237) );
  ANDN U51610 ( .B(n36238), .A(n36237), .Z(n36239) );
  NAND U51611 ( .A(n36240), .B(n36239), .Z(n36241) );
  NANDN U51612 ( .A(n36242), .B(n36241), .Z(n36243) );
  OR U51613 ( .A(n36244), .B(n36243), .Z(n36245) );
  AND U51614 ( .A(n36246), .B(n36245), .Z(n36248) );
  NAND U51615 ( .A(n36248), .B(n36247), .Z(n36249) );
  NAND U51616 ( .A(n36250), .B(n36249), .Z(n36251) );
  NANDN U51617 ( .A(n36252), .B(n36251), .Z(n36253) );
  AND U51618 ( .A(n36254), .B(n36253), .Z(n36256) );
  NAND U51619 ( .A(n36256), .B(n36255), .Z(n36257) );
  NANDN U51620 ( .A(n36258), .B(n36257), .Z(n36259) );
  AND U51621 ( .A(n36260), .B(n36259), .Z(n36261) );
  NANDN U51622 ( .A(n36262), .B(n36261), .Z(n36263) );
  NAND U51623 ( .A(n36264), .B(n36263), .Z(n36265) );
  NANDN U51624 ( .A(n36266), .B(n36265), .Z(n36268) );
  ANDN U51625 ( .B(y[2646]), .A(x[2646]), .Z(n36267) );
  OR U51626 ( .A(n36268), .B(n36267), .Z(n36269) );
  NANDN U51627 ( .A(n36270), .B(n36269), .Z(n36271) );
  AND U51628 ( .A(n36272), .B(n36271), .Z(n36276) );
  NAND U51629 ( .A(n36274), .B(n36273), .Z(n36275) );
  OR U51630 ( .A(n36276), .B(n36275), .Z(n36277) );
  AND U51631 ( .A(n36278), .B(n36277), .Z(n36279) );
  OR U51632 ( .A(n36280), .B(n36279), .Z(n36281) );
  NAND U51633 ( .A(n36282), .B(n36281), .Z(n36283) );
  AND U51634 ( .A(n36284), .B(n36283), .Z(n36285) );
  OR U51635 ( .A(n36286), .B(n36285), .Z(n36287) );
  NAND U51636 ( .A(n36288), .B(n36287), .Z(n36292) );
  NAND U51637 ( .A(n36290), .B(n36289), .Z(n36291) );
  ANDN U51638 ( .B(n36292), .A(n36291), .Z(n36296) );
  NAND U51639 ( .A(n36294), .B(n36293), .Z(n36295) );
  OR U51640 ( .A(n36296), .B(n36295), .Z(n36297) );
  AND U51641 ( .A(n36298), .B(n36297), .Z(n36302) );
  NAND U51642 ( .A(n36300), .B(n36299), .Z(n36301) );
  OR U51643 ( .A(n36302), .B(n36301), .Z(n36303) );
  AND U51644 ( .A(n36304), .B(n36303), .Z(n36308) );
  NAND U51645 ( .A(n36306), .B(n36305), .Z(n36307) );
  OR U51646 ( .A(n36308), .B(n36307), .Z(n36309) );
  AND U51647 ( .A(n36310), .B(n36309), .Z(n36314) );
  NAND U51648 ( .A(n36312), .B(n36311), .Z(n36313) );
  OR U51649 ( .A(n36314), .B(n36313), .Z(n36315) );
  AND U51650 ( .A(n36316), .B(n36315), .Z(n36320) );
  NAND U51651 ( .A(n36318), .B(n36317), .Z(n36319) );
  OR U51652 ( .A(n36320), .B(n36319), .Z(n36321) );
  AND U51653 ( .A(n36322), .B(n36321), .Z(n36326) );
  NAND U51654 ( .A(n36324), .B(n36323), .Z(n36325) );
  OR U51655 ( .A(n36326), .B(n36325), .Z(n36327) );
  AND U51656 ( .A(n36328), .B(n36327), .Z(n36329) );
  ANDN U51657 ( .B(n36330), .A(n36329), .Z(n36331) );
  NAND U51658 ( .A(n36332), .B(n36331), .Z(n36333) );
  NANDN U51659 ( .A(n54836), .B(n36333), .Z(n36334) );
  OR U51660 ( .A(n36335), .B(n36334), .Z(n36336) );
  AND U51661 ( .A(n36337), .B(n36336), .Z(n36339) );
  NAND U51662 ( .A(n36339), .B(n36338), .Z(n36340) );
  NANDN U51663 ( .A(n36341), .B(n36340), .Z(n36342) );
  AND U51664 ( .A(n36343), .B(n36342), .Z(n36345) );
  NAND U51665 ( .A(n36345), .B(n36344), .Z(n36346) );
  NANDN U51666 ( .A(n36347), .B(n36346), .Z(n36348) );
  AND U51667 ( .A(n36349), .B(n36348), .Z(n36351) );
  AND U51668 ( .A(n36351), .B(n36350), .Z(n36355) );
  NAND U51669 ( .A(n36353), .B(n36352), .Z(n36354) );
  OR U51670 ( .A(n36355), .B(n36354), .Z(n36356) );
  AND U51671 ( .A(n36357), .B(n36356), .Z(n36361) );
  NAND U51672 ( .A(n36359), .B(n36358), .Z(n36360) );
  OR U51673 ( .A(n36361), .B(n36360), .Z(n36362) );
  AND U51674 ( .A(n36363), .B(n36362), .Z(n36367) );
  NAND U51675 ( .A(n36365), .B(n36364), .Z(n36366) );
  OR U51676 ( .A(n36367), .B(n36366), .Z(n36368) );
  AND U51677 ( .A(n36369), .B(n36368), .Z(n36373) );
  NAND U51678 ( .A(n36371), .B(n36370), .Z(n36372) );
  OR U51679 ( .A(n36373), .B(n36372), .Z(n36374) );
  AND U51680 ( .A(n36375), .B(n36374), .Z(n36379) );
  NAND U51681 ( .A(n36377), .B(n36376), .Z(n36378) );
  OR U51682 ( .A(n36379), .B(n36378), .Z(n36380) );
  AND U51683 ( .A(n36381), .B(n36380), .Z(n36385) );
  NAND U51684 ( .A(n36383), .B(n36382), .Z(n36384) );
  OR U51685 ( .A(n36385), .B(n36384), .Z(n36386) );
  AND U51686 ( .A(n36387), .B(n36386), .Z(n36391) );
  NANDN U51687 ( .A(x[2688]), .B(y[2688]), .Z(n36389) );
  NAND U51688 ( .A(n36389), .B(n36388), .Z(n36390) );
  OR U51689 ( .A(n36391), .B(n36390), .Z(n36392) );
  AND U51690 ( .A(n36393), .B(n36392), .Z(n36394) );
  OR U51691 ( .A(n36395), .B(n36394), .Z(n36396) );
  NAND U51692 ( .A(n36397), .B(n36396), .Z(n36398) );
  AND U51693 ( .A(n36399), .B(n36398), .Z(n36400) );
  OR U51694 ( .A(n36401), .B(n36400), .Z(n36402) );
  NAND U51695 ( .A(n36403), .B(n36402), .Z(n36407) );
  NAND U51696 ( .A(n36405), .B(n36404), .Z(n36406) );
  ANDN U51697 ( .B(n36407), .A(n36406), .Z(n36411) );
  NAND U51698 ( .A(n36409), .B(n36408), .Z(n36410) );
  OR U51699 ( .A(n36411), .B(n36410), .Z(n36412) );
  AND U51700 ( .A(n36413), .B(n36412), .Z(n36417) );
  NAND U51701 ( .A(n36415), .B(n36414), .Z(n36416) );
  OR U51702 ( .A(n36417), .B(n36416), .Z(n36418) );
  AND U51703 ( .A(n36419), .B(n36418), .Z(n36422) );
  NAND U51704 ( .A(n36420), .B(n54867), .Z(n36421) );
  OR U51705 ( .A(n36422), .B(n36421), .Z(n36423) );
  AND U51706 ( .A(n36424), .B(n36423), .Z(n36427) );
  NANDN U51707 ( .A(x[2702]), .B(y[2702]), .Z(n54868) );
  AND U51708 ( .A(n36425), .B(n54868), .Z(n36426) );
  NANDN U51709 ( .A(n36427), .B(n36426), .Z(n36428) );
  NANDN U51710 ( .A(n36429), .B(n36428), .Z(n36430) );
  AND U51711 ( .A(n36431), .B(n36430), .Z(n36433) );
  NOR U51712 ( .A(n36433), .B(n36432), .Z(n36434) );
  NANDN U51713 ( .A(n36435), .B(n36434), .Z(n36436) );
  AND U51714 ( .A(n36437), .B(n36436), .Z(n36439) );
  NAND U51715 ( .A(n36439), .B(n36438), .Z(n36440) );
  NANDN U51716 ( .A(n36441), .B(n36440), .Z(n36442) );
  AND U51717 ( .A(n52024), .B(n36442), .Z(n36443) );
  NANDN U51718 ( .A(n36444), .B(n36443), .Z(n36445) );
  AND U51719 ( .A(n36446), .B(n36445), .Z(n36448) );
  NAND U51720 ( .A(n36448), .B(n36447), .Z(n36449) );
  ANDN U51721 ( .B(y[2710]), .A(x[2710]), .Z(n52023) );
  ANDN U51722 ( .B(n36449), .A(n52023), .Z(n36451) );
  ANDN U51723 ( .B(n36451), .A(n36450), .Z(n36452) );
  OR U51724 ( .A(n36453), .B(n36452), .Z(n36454) );
  NAND U51725 ( .A(n36455), .B(n36454), .Z(n36456) );
  AND U51726 ( .A(n36457), .B(n36456), .Z(n36458) );
  NOR U51727 ( .A(n54881), .B(n36458), .Z(n36459) );
  NANDN U51728 ( .A(n54883), .B(n36459), .Z(n36460) );
  AND U51729 ( .A(n36461), .B(n36460), .Z(n36463) );
  NAND U51730 ( .A(n36463), .B(n36462), .Z(n36464) );
  NANDN U51731 ( .A(n36465), .B(n36464), .Z(n36466) );
  AND U51732 ( .A(n36467), .B(n36466), .Z(n36469) );
  NAND U51733 ( .A(n36469), .B(n36468), .Z(n36470) );
  NANDN U51734 ( .A(n36471), .B(n36470), .Z(n36472) );
  AND U51735 ( .A(n36473), .B(n36472), .Z(n36475) );
  AND U51736 ( .A(n36475), .B(n36474), .Z(n36479) );
  NAND U51737 ( .A(n36477), .B(n36476), .Z(n36478) );
  OR U51738 ( .A(n36479), .B(n36478), .Z(n36480) );
  AND U51739 ( .A(n36481), .B(n36480), .Z(n36485) );
  NAND U51740 ( .A(n36483), .B(n36482), .Z(n36484) );
  OR U51741 ( .A(n36485), .B(n36484), .Z(n36486) );
  AND U51742 ( .A(n36487), .B(n36486), .Z(n36491) );
  NAND U51743 ( .A(n36489), .B(n36488), .Z(n36490) );
  OR U51744 ( .A(n36491), .B(n36490), .Z(n36492) );
  AND U51745 ( .A(n36493), .B(n36492), .Z(n36497) );
  NAND U51746 ( .A(n36495), .B(n36494), .Z(n36496) );
  OR U51747 ( .A(n36497), .B(n36496), .Z(n36498) );
  AND U51748 ( .A(n36499), .B(n36498), .Z(n36503) );
  NAND U51749 ( .A(n36501), .B(n36500), .Z(n36502) );
  OR U51750 ( .A(n36503), .B(n36502), .Z(n36504) );
  AND U51751 ( .A(n36505), .B(n36504), .Z(n36509) );
  NAND U51752 ( .A(n36507), .B(n36506), .Z(n36508) );
  OR U51753 ( .A(n36509), .B(n36508), .Z(n36510) );
  AND U51754 ( .A(n36511), .B(n36510), .Z(n36515) );
  NAND U51755 ( .A(n36513), .B(n36512), .Z(n36514) );
  OR U51756 ( .A(n36515), .B(n36514), .Z(n36516) );
  AND U51757 ( .A(n36517), .B(n36516), .Z(n36520) );
  NAND U51758 ( .A(n52022), .B(n36518), .Z(n36519) );
  OR U51759 ( .A(n36520), .B(n36519), .Z(n36521) );
  AND U51760 ( .A(n36522), .B(n36521), .Z(n36523) );
  OR U51761 ( .A(n54928), .B(n36523), .Z(n36524) );
  NAND U51762 ( .A(n36525), .B(n36524), .Z(n36526) );
  NANDN U51763 ( .A(n36527), .B(n36526), .Z(n36529) );
  IV U51764 ( .A(n36528), .Z(n54930) );
  OR U51765 ( .A(n36529), .B(n54930), .Z(n36530) );
  NANDN U51766 ( .A(n36531), .B(n36530), .Z(n36532) );
  AND U51767 ( .A(n36533), .B(n36532), .Z(n36538) );
  OR U51768 ( .A(n36535), .B(n36534), .Z(n36536) );
  AND U51769 ( .A(n54934), .B(n36536), .Z(n36537) );
  NANDN U51770 ( .A(n36538), .B(n36537), .Z(n36539) );
  AND U51771 ( .A(n36540), .B(n36539), .Z(n36541) );
  OR U51772 ( .A(n36542), .B(n36541), .Z(n36543) );
  NAND U51773 ( .A(n36544), .B(n36543), .Z(n36545) );
  NANDN U51774 ( .A(n36546), .B(n36545), .Z(n36548) );
  OR U51775 ( .A(n36548), .B(n36547), .Z(n36549) );
  NAND U51776 ( .A(n36550), .B(n36549), .Z(n36551) );
  NANDN U51777 ( .A(n36552), .B(n36551), .Z(n36553) );
  AND U51778 ( .A(n36554), .B(n36553), .Z(n36555) );
  NOR U51779 ( .A(n36556), .B(n36555), .Z(n36558) );
  NAND U51780 ( .A(n36558), .B(n36557), .Z(n36560) );
  AND U51781 ( .A(n36560), .B(n36559), .Z(n36561) );
  NANDN U51782 ( .A(x[2750]), .B(y[2750]), .Z(n52020) );
  NAND U51783 ( .A(n36561), .B(n52020), .Z(n36562) );
  NANDN U51784 ( .A(n36563), .B(n36562), .Z(n36564) );
  AND U51785 ( .A(n36565), .B(n36564), .Z(n36567) );
  NAND U51786 ( .A(n36567), .B(n36566), .Z(n36568) );
  NANDN U51787 ( .A(n36569), .B(n36568), .Z(n36570) );
  AND U51788 ( .A(n36571), .B(n36570), .Z(n36573) );
  NAND U51789 ( .A(n36573), .B(n36572), .Z(n36574) );
  NANDN U51790 ( .A(n36575), .B(n36574), .Z(n36576) );
  AND U51791 ( .A(n36577), .B(n36576), .Z(n36579) );
  NAND U51792 ( .A(n36579), .B(n36578), .Z(n36580) );
  NANDN U51793 ( .A(n36581), .B(n36580), .Z(n36582) );
  AND U51794 ( .A(n36583), .B(n36582), .Z(n36585) );
  AND U51795 ( .A(n36585), .B(n36584), .Z(n36589) );
  NAND U51796 ( .A(n36587), .B(n36586), .Z(n36588) );
  OR U51797 ( .A(n36589), .B(n36588), .Z(n36590) );
  AND U51798 ( .A(n36591), .B(n36590), .Z(n36595) );
  NAND U51799 ( .A(n36593), .B(n36592), .Z(n36594) );
  OR U51800 ( .A(n36595), .B(n36594), .Z(n36596) );
  AND U51801 ( .A(n36597), .B(n36596), .Z(n36598) );
  ANDN U51802 ( .B(n36599), .A(n36598), .Z(n36600) );
  NAND U51803 ( .A(n36601), .B(n36600), .Z(n36602) );
  NANDN U51804 ( .A(n36603), .B(n36602), .Z(n36604) );
  OR U51805 ( .A(n36605), .B(n36604), .Z(n36606) );
  AND U51806 ( .A(n36607), .B(n36606), .Z(n36609) );
  NAND U51807 ( .A(n36609), .B(n36608), .Z(n36610) );
  NANDN U51808 ( .A(n36611), .B(n36610), .Z(n36612) );
  AND U51809 ( .A(n36613), .B(n36612), .Z(n36615) );
  NAND U51810 ( .A(n36615), .B(n36614), .Z(n36616) );
  NANDN U51811 ( .A(n36617), .B(n36616), .Z(n36618) );
  AND U51812 ( .A(n36619), .B(n36618), .Z(n36621) );
  AND U51813 ( .A(n36621), .B(n36620), .Z(n36625) );
  NAND U51814 ( .A(n36623), .B(n36622), .Z(n36624) );
  OR U51815 ( .A(n36625), .B(n36624), .Z(n36626) );
  AND U51816 ( .A(n36627), .B(n36626), .Z(n36631) );
  NAND U51817 ( .A(n36629), .B(n36628), .Z(n36630) );
  OR U51818 ( .A(n36631), .B(n36630), .Z(n36632) );
  AND U51819 ( .A(n36633), .B(n36632), .Z(n36634) );
  OR U51820 ( .A(n36635), .B(n36634), .Z(n36636) );
  NAND U51821 ( .A(n36637), .B(n36636), .Z(n36638) );
  NANDN U51822 ( .A(n54984), .B(n36638), .Z(n36639) );
  ANDN U51823 ( .B(y[2776]), .A(x[2776]), .Z(n54980) );
  OR U51824 ( .A(n36639), .B(n54980), .Z(n36640) );
  NAND U51825 ( .A(n36641), .B(n36640), .Z(n36642) );
  NANDN U51826 ( .A(n36643), .B(n36642), .Z(n36644) );
  ANDN U51827 ( .B(y[2778]), .A(x[2778]), .Z(n54986) );
  OR U51828 ( .A(n36644), .B(n54986), .Z(n36645) );
  NAND U51829 ( .A(n36646), .B(n36645), .Z(n36647) );
  NANDN U51830 ( .A(n36648), .B(n36647), .Z(n36650) );
  OR U51831 ( .A(n36650), .B(n36649), .Z(n36651) );
  NAND U51832 ( .A(n36652), .B(n36651), .Z(n36656) );
  NAND U51833 ( .A(n36654), .B(n36653), .Z(n36655) );
  ANDN U51834 ( .B(n36656), .A(n36655), .Z(n36660) );
  NAND U51835 ( .A(n36658), .B(n36657), .Z(n36659) );
  OR U51836 ( .A(n36660), .B(n36659), .Z(n36661) );
  AND U51837 ( .A(n36662), .B(n36661), .Z(n36666) );
  NAND U51838 ( .A(n36664), .B(n36663), .Z(n36665) );
  OR U51839 ( .A(n36666), .B(n36665), .Z(n36667) );
  AND U51840 ( .A(n36668), .B(n36667), .Z(n36670) );
  AND U51841 ( .A(n36670), .B(n36669), .Z(n36674) );
  NAND U51842 ( .A(n36672), .B(n36671), .Z(n36673) );
  OR U51843 ( .A(n36674), .B(n36673), .Z(n36675) );
  AND U51844 ( .A(n36676), .B(n36675), .Z(n36680) );
  AND U51845 ( .A(n36678), .B(n36677), .Z(n36679) );
  NANDN U51846 ( .A(n36680), .B(n36679), .Z(n36681) );
  NAND U51847 ( .A(n36682), .B(n36681), .Z(n36683) );
  AND U51848 ( .A(n36684), .B(n36683), .Z(n36685) );
  NOR U51849 ( .A(n36686), .B(n36685), .Z(n36687) );
  NANDN U51850 ( .A(n36688), .B(n36687), .Z(n36689) );
  AND U51851 ( .A(n36690), .B(n36689), .Z(n36692) );
  NAND U51852 ( .A(n36692), .B(n36691), .Z(n36693) );
  NANDN U51853 ( .A(n36694), .B(n36693), .Z(n36695) );
  NAND U51854 ( .A(n36696), .B(n36695), .Z(n36697) );
  AND U51855 ( .A(n36698), .B(n36697), .Z(n36699) );
  OR U51856 ( .A(n55010), .B(n36699), .Z(n36700) );
  NAND U51857 ( .A(n36701), .B(n36700), .Z(n36702) );
  NANDN U51858 ( .A(n36703), .B(n36702), .Z(n36704) );
  NAND U51859 ( .A(n36705), .B(n36704), .Z(n36706) );
  NANDN U51860 ( .A(n36707), .B(n36706), .Z(n36708) );
  AND U51861 ( .A(n36709), .B(n36708), .Z(n36711) );
  NAND U51862 ( .A(n36711), .B(n36710), .Z(n36712) );
  NANDN U51863 ( .A(n36713), .B(n36712), .Z(n36714) );
  AND U51864 ( .A(n36715), .B(n36714), .Z(n36717) );
  NAND U51865 ( .A(n36717), .B(n36716), .Z(n36718) );
  NANDN U51866 ( .A(n36719), .B(n36718), .Z(n36720) );
  AND U51867 ( .A(n36721), .B(n36720), .Z(n36723) );
  AND U51868 ( .A(n36723), .B(n36722), .Z(n36727) );
  NAND U51869 ( .A(n36725), .B(n36724), .Z(n36726) );
  OR U51870 ( .A(n36727), .B(n36726), .Z(n36728) );
  AND U51871 ( .A(n36729), .B(n36728), .Z(n36733) );
  NAND U51872 ( .A(n36731), .B(n36730), .Z(n36732) );
  OR U51873 ( .A(n36733), .B(n36732), .Z(n36734) );
  AND U51874 ( .A(n36735), .B(n36734), .Z(n36739) );
  NAND U51875 ( .A(n36737), .B(n36736), .Z(n36738) );
  OR U51876 ( .A(n36739), .B(n36738), .Z(n36740) );
  AND U51877 ( .A(n36741), .B(n36740), .Z(n36745) );
  NAND U51878 ( .A(n36743), .B(n36742), .Z(n36744) );
  OR U51879 ( .A(n36745), .B(n36744), .Z(n36746) );
  AND U51880 ( .A(n36747), .B(n36746), .Z(n36751) );
  NAND U51881 ( .A(n36749), .B(n36748), .Z(n36750) );
  OR U51882 ( .A(n36751), .B(n36750), .Z(n36752) );
  AND U51883 ( .A(n36753), .B(n36752), .Z(n36757) );
  NAND U51884 ( .A(n36755), .B(n36754), .Z(n36756) );
  OR U51885 ( .A(n36757), .B(n36756), .Z(n36758) );
  AND U51886 ( .A(n36759), .B(n36758), .Z(n36760) );
  OR U51887 ( .A(n36761), .B(n36760), .Z(n36762) );
  NAND U51888 ( .A(n36763), .B(n36762), .Z(n36764) );
  NAND U51889 ( .A(n36765), .B(n36764), .Z(n36766) );
  NANDN U51890 ( .A(n36767), .B(n36766), .Z(n36768) );
  AND U51891 ( .A(n36769), .B(n36768), .Z(n36771) );
  NAND U51892 ( .A(n36771), .B(n36770), .Z(n36772) );
  NANDN U51893 ( .A(n36773), .B(n36772), .Z(n36774) );
  AND U51894 ( .A(n36775), .B(n36774), .Z(n36776) );
  NANDN U51895 ( .A(n36777), .B(n36776), .Z(n36778) );
  NAND U51896 ( .A(n36779), .B(n36778), .Z(n36780) );
  NANDN U51897 ( .A(n36781), .B(n36780), .Z(n36782) );
  AND U51898 ( .A(n36783), .B(n36782), .Z(n36784) );
  NAND U51899 ( .A(n36785), .B(n36784), .Z(n36789) );
  NAND U51900 ( .A(n36787), .B(n36786), .Z(n36788) );
  ANDN U51901 ( .B(n36789), .A(n36788), .Z(n36793) );
  NAND U51902 ( .A(n36791), .B(n36790), .Z(n36792) );
  OR U51903 ( .A(n36793), .B(n36792), .Z(n36794) );
  AND U51904 ( .A(n36795), .B(n36794), .Z(n36799) );
  NAND U51905 ( .A(n36797), .B(n36796), .Z(n36798) );
  OR U51906 ( .A(n36799), .B(n36798), .Z(n36800) );
  AND U51907 ( .A(n36801), .B(n36800), .Z(n36805) );
  NAND U51908 ( .A(n36803), .B(n36802), .Z(n36804) );
  OR U51909 ( .A(n36805), .B(n36804), .Z(n36806) );
  AND U51910 ( .A(n36807), .B(n36806), .Z(n36810) );
  NAND U51911 ( .A(n36808), .B(n55052), .Z(n36809) );
  OR U51912 ( .A(n36810), .B(n36809), .Z(n36811) );
  AND U51913 ( .A(n36812), .B(n36811), .Z(n36813) );
  OR U51914 ( .A(n36814), .B(n36813), .Z(n36815) );
  NAND U51915 ( .A(n36816), .B(n36815), .Z(n36820) );
  NANDN U51916 ( .A(x[2838]), .B(y[2838]), .Z(n36817) );
  AND U51917 ( .A(n36818), .B(n36817), .Z(n36819) );
  NAND U51918 ( .A(n36820), .B(n36819), .Z(n36821) );
  NANDN U51919 ( .A(n36822), .B(n36821), .Z(n36823) );
  NAND U51920 ( .A(n36824), .B(n36823), .Z(n36825) );
  NAND U51921 ( .A(n36826), .B(n36825), .Z(n36827) );
  NANDN U51922 ( .A(n36828), .B(n36827), .Z(n36830) );
  ANDN U51923 ( .B(y[2842]), .A(x[2842]), .Z(n36829) );
  OR U51924 ( .A(n36830), .B(n36829), .Z(n36831) );
  NAND U51925 ( .A(n36832), .B(n36831), .Z(n36833) );
  NANDN U51926 ( .A(n36834), .B(n36833), .Z(n36836) );
  ANDN U51927 ( .B(y[2844]), .A(x[2844]), .Z(n36835) );
  OR U51928 ( .A(n36836), .B(n36835), .Z(n36837) );
  NAND U51929 ( .A(n36838), .B(n36837), .Z(n36839) );
  NANDN U51930 ( .A(n36840), .B(n36839), .Z(n36841) );
  AND U51931 ( .A(n36842), .B(n36841), .Z(n36843) );
  NAND U51932 ( .A(n36844), .B(n36843), .Z(n36848) );
  NAND U51933 ( .A(n36846), .B(n36845), .Z(n36847) );
  ANDN U51934 ( .B(n36848), .A(n36847), .Z(n36852) );
  NAND U51935 ( .A(n36850), .B(n36849), .Z(n36851) );
  OR U51936 ( .A(n36852), .B(n36851), .Z(n36853) );
  AND U51937 ( .A(n36854), .B(n36853), .Z(n36858) );
  NAND U51938 ( .A(n36856), .B(n36855), .Z(n36857) );
  OR U51939 ( .A(n36858), .B(n36857), .Z(n36859) );
  AND U51940 ( .A(n36860), .B(n36859), .Z(n36864) );
  NAND U51941 ( .A(n36862), .B(n36861), .Z(n36863) );
  OR U51942 ( .A(n36864), .B(n36863), .Z(n36865) );
  AND U51943 ( .A(n36866), .B(n36865), .Z(n36867) );
  ANDN U51944 ( .B(n36868), .A(n36867), .Z(n36869) );
  NAND U51945 ( .A(n36870), .B(n36869), .Z(n36871) );
  NANDN U51946 ( .A(n36872), .B(n36871), .Z(n36873) );
  OR U51947 ( .A(n36874), .B(n36873), .Z(n36875) );
  AND U51948 ( .A(n36876), .B(n36875), .Z(n36878) );
  NAND U51949 ( .A(n36878), .B(n36877), .Z(n36879) );
  NANDN U51950 ( .A(n36880), .B(n36879), .Z(n36881) );
  AND U51951 ( .A(n36882), .B(n36881), .Z(n36884) );
  NAND U51952 ( .A(n36884), .B(n36883), .Z(n36885) );
  NANDN U51953 ( .A(n36886), .B(n36885), .Z(n36887) );
  AND U51954 ( .A(n36888), .B(n36887), .Z(n36890) );
  AND U51955 ( .A(n36890), .B(n36889), .Z(n36894) );
  NAND U51956 ( .A(n36892), .B(n36891), .Z(n36893) );
  OR U51957 ( .A(n36894), .B(n36893), .Z(n36895) );
  AND U51958 ( .A(n36896), .B(n36895), .Z(n36900) );
  NAND U51959 ( .A(n36898), .B(n36897), .Z(n36899) );
  OR U51960 ( .A(n36900), .B(n36899), .Z(n36901) );
  AND U51961 ( .A(n36902), .B(n36901), .Z(n36906) );
  NAND U51962 ( .A(n36904), .B(n36903), .Z(n36905) );
  OR U51963 ( .A(n36906), .B(n36905), .Z(n36907) );
  AND U51964 ( .A(n36908), .B(n36907), .Z(n36912) );
  NAND U51965 ( .A(n36910), .B(n36909), .Z(n36911) );
  OR U51966 ( .A(n36912), .B(n36911), .Z(n36913) );
  AND U51967 ( .A(n36914), .B(n36913), .Z(n36918) );
  NAND U51968 ( .A(n36916), .B(n36915), .Z(n36917) );
  OR U51969 ( .A(n36918), .B(n36917), .Z(n36919) );
  AND U51970 ( .A(n36920), .B(n36919), .Z(n36921) );
  OR U51971 ( .A(n36922), .B(n36921), .Z(n36923) );
  NAND U51972 ( .A(n36924), .B(n36923), .Z(n36928) );
  NANDN U51973 ( .A(x[2874]), .B(y[2874]), .Z(n36925) );
  AND U51974 ( .A(n36926), .B(n36925), .Z(n36927) );
  NAND U51975 ( .A(n36928), .B(n36927), .Z(n36929) );
  NANDN U51976 ( .A(n36930), .B(n36929), .Z(n36931) );
  NAND U51977 ( .A(n36932), .B(n36931), .Z(n36933) );
  NANDN U51978 ( .A(n36934), .B(n36933), .Z(n36935) );
  AND U51979 ( .A(n36936), .B(n36935), .Z(n36938) );
  NANDN U51980 ( .A(x[2878]), .B(y[2878]), .Z(n36937) );
  NAND U51981 ( .A(n36938), .B(n36937), .Z(n36939) );
  NANDN U51982 ( .A(n36940), .B(n36939), .Z(n36941) );
  AND U51983 ( .A(n36942), .B(n36941), .Z(n36944) );
  NAND U51984 ( .A(n36944), .B(n36943), .Z(n36945) );
  NANDN U51985 ( .A(n36946), .B(n36945), .Z(n36947) );
  AND U51986 ( .A(n36948), .B(n36947), .Z(n36950) );
  NAND U51987 ( .A(n36950), .B(n36949), .Z(n36951) );
  NANDN U51988 ( .A(n36952), .B(n36951), .Z(n36953) );
  AND U51989 ( .A(n36954), .B(n36953), .Z(n36956) );
  NAND U51990 ( .A(n36956), .B(n36955), .Z(n36957) );
  AND U51991 ( .A(n36958), .B(n36957), .Z(n36959) );
  ANDN U51992 ( .B(n36960), .A(n36959), .Z(n36961) );
  OR U51993 ( .A(n36962), .B(n36961), .Z(n36963) );
  NAND U51994 ( .A(n51993), .B(n36963), .Z(n36964) );
  NANDN U51995 ( .A(n36965), .B(n36964), .Z(n36966) );
  OR U51996 ( .A(n36966), .B(n55095), .Z(n36967) );
  NANDN U51997 ( .A(n36968), .B(n36967), .Z(n36969) );
  AND U51998 ( .A(n36970), .B(n36969), .Z(n36974) );
  NAND U51999 ( .A(n36972), .B(n36971), .Z(n36973) );
  OR U52000 ( .A(n36974), .B(n36973), .Z(n36975) );
  AND U52001 ( .A(n36976), .B(n36975), .Z(n36980) );
  NAND U52002 ( .A(n36978), .B(n36977), .Z(n36979) );
  OR U52003 ( .A(n36980), .B(n36979), .Z(n36981) );
  AND U52004 ( .A(n36982), .B(n36981), .Z(n36986) );
  NAND U52005 ( .A(n36984), .B(n36983), .Z(n36985) );
  OR U52006 ( .A(n36986), .B(n36985), .Z(n36987) );
  AND U52007 ( .A(n36988), .B(n36987), .Z(n36992) );
  NAND U52008 ( .A(n36990), .B(n36989), .Z(n36991) );
  OR U52009 ( .A(n36992), .B(n36991), .Z(n36993) );
  AND U52010 ( .A(n36994), .B(n36993), .Z(n36998) );
  NAND U52011 ( .A(n36996), .B(n36995), .Z(n36997) );
  OR U52012 ( .A(n36998), .B(n36997), .Z(n36999) );
  AND U52013 ( .A(n37000), .B(n36999), .Z(n37001) );
  OR U52014 ( .A(n37002), .B(n37001), .Z(n37003) );
  NAND U52015 ( .A(n37004), .B(n37003), .Z(n37005) );
  AND U52016 ( .A(n37006), .B(n37005), .Z(n37007) );
  NOR U52017 ( .A(n37008), .B(n37007), .Z(n37010) );
  NAND U52018 ( .A(n37010), .B(n37009), .Z(n37014) );
  NANDN U52019 ( .A(x[2906]), .B(y[2906]), .Z(n37011) );
  AND U52020 ( .A(n37012), .B(n37011), .Z(n37013) );
  NAND U52021 ( .A(n37014), .B(n37013), .Z(n37015) );
  NANDN U52022 ( .A(n37016), .B(n37015), .Z(n37017) );
  NAND U52023 ( .A(n37018), .B(n37017), .Z(n37019) );
  NAND U52024 ( .A(n37020), .B(n37019), .Z(n37021) );
  NANDN U52025 ( .A(n37022), .B(n37021), .Z(n37024) );
  ANDN U52026 ( .B(y[2910]), .A(x[2910]), .Z(n37023) );
  OR U52027 ( .A(n37024), .B(n37023), .Z(n37025) );
  NAND U52028 ( .A(n37026), .B(n37025), .Z(n37027) );
  NANDN U52029 ( .A(n37028), .B(n37027), .Z(n37030) );
  OR U52030 ( .A(n37030), .B(n37029), .Z(n37031) );
  NANDN U52031 ( .A(n37032), .B(n37031), .Z(n37033) );
  AND U52032 ( .A(n37034), .B(n37033), .Z(n37038) );
  NAND U52033 ( .A(n37036), .B(n37035), .Z(n37037) );
  OR U52034 ( .A(n37038), .B(n37037), .Z(n37039) );
  AND U52035 ( .A(n37040), .B(n37039), .Z(n37044) );
  NAND U52036 ( .A(n37042), .B(n37041), .Z(n37043) );
  OR U52037 ( .A(n37044), .B(n37043), .Z(n37045) );
  AND U52038 ( .A(n37046), .B(n37045), .Z(n37050) );
  NAND U52039 ( .A(n37048), .B(n37047), .Z(n37049) );
  OR U52040 ( .A(n37050), .B(n37049), .Z(n37051) );
  AND U52041 ( .A(n37052), .B(n37051), .Z(n37056) );
  NAND U52042 ( .A(n37054), .B(n37053), .Z(n37055) );
  OR U52043 ( .A(n37056), .B(n37055), .Z(n37057) );
  AND U52044 ( .A(n37058), .B(n37057), .Z(n37062) );
  NAND U52045 ( .A(n37060), .B(n37059), .Z(n37061) );
  OR U52046 ( .A(n37062), .B(n37061), .Z(n37063) );
  AND U52047 ( .A(n37064), .B(n37063), .Z(n37068) );
  NAND U52048 ( .A(n37066), .B(n37065), .Z(n37067) );
  OR U52049 ( .A(n37068), .B(n37067), .Z(n37069) );
  AND U52050 ( .A(n37070), .B(n37069), .Z(n37074) );
  NAND U52051 ( .A(n37072), .B(n37071), .Z(n37073) );
  OR U52052 ( .A(n37074), .B(n37073), .Z(n37075) );
  AND U52053 ( .A(n37076), .B(n37075), .Z(n37080) );
  NAND U52054 ( .A(n37078), .B(n37077), .Z(n37079) );
  OR U52055 ( .A(n37080), .B(n37079), .Z(n37081) );
  AND U52056 ( .A(n37082), .B(n37081), .Z(n37086) );
  NAND U52057 ( .A(n37084), .B(n37083), .Z(n37085) );
  OR U52058 ( .A(n37086), .B(n37085), .Z(n37087) );
  AND U52059 ( .A(n37088), .B(n37087), .Z(n37092) );
  NAND U52060 ( .A(n37090), .B(n37089), .Z(n37091) );
  OR U52061 ( .A(n37092), .B(n37091), .Z(n37093) );
  AND U52062 ( .A(n37094), .B(n37093), .Z(n37098) );
  NAND U52063 ( .A(n37096), .B(n37095), .Z(n37097) );
  OR U52064 ( .A(n37098), .B(n37097), .Z(n37099) );
  AND U52065 ( .A(n37100), .B(n37099), .Z(n37104) );
  NAND U52066 ( .A(n37102), .B(n37101), .Z(n37103) );
  OR U52067 ( .A(n37104), .B(n37103), .Z(n37105) );
  AND U52068 ( .A(n37106), .B(n37105), .Z(n37110) );
  NAND U52069 ( .A(n37108), .B(n37107), .Z(n37109) );
  OR U52070 ( .A(n37110), .B(n37109), .Z(n37111) );
  AND U52071 ( .A(n37112), .B(n37111), .Z(n37113) );
  NOR U52072 ( .A(n37114), .B(n37113), .Z(n37115) );
  NAND U52073 ( .A(n37116), .B(n37115), .Z(n37117) );
  NANDN U52074 ( .A(n37118), .B(n37117), .Z(n37119) );
  NAND U52075 ( .A(n37120), .B(n37119), .Z(n37121) );
  NANDN U52076 ( .A(n37122), .B(n37121), .Z(n37123) );
  AND U52077 ( .A(n37124), .B(n37123), .Z(n37126) );
  NAND U52078 ( .A(n37126), .B(n37125), .Z(n37127) );
  NANDN U52079 ( .A(n37128), .B(n37127), .Z(n37129) );
  AND U52080 ( .A(n37130), .B(n37129), .Z(n37132) );
  NAND U52081 ( .A(n37132), .B(n37131), .Z(n37133) );
  NANDN U52082 ( .A(n37134), .B(n37133), .Z(n37135) );
  AND U52083 ( .A(n37136), .B(n37135), .Z(n37138) );
  AND U52084 ( .A(n37138), .B(n37137), .Z(n37139) );
  OR U52085 ( .A(n37140), .B(n37139), .Z(n37141) );
  NAND U52086 ( .A(n37142), .B(n37141), .Z(n37143) );
  AND U52087 ( .A(n37144), .B(n37143), .Z(n37145) );
  ANDN U52088 ( .B(n37146), .A(n37145), .Z(n37147) );
  OR U52089 ( .A(n37148), .B(n37147), .Z(n37149) );
  NAND U52090 ( .A(n37150), .B(n37149), .Z(n37151) );
  NAND U52091 ( .A(n37152), .B(n37151), .Z(n37153) );
  NANDN U52092 ( .A(n37154), .B(n37153), .Z(n37155) );
  AND U52093 ( .A(n37156), .B(n37155), .Z(n37158) );
  NAND U52094 ( .A(n37158), .B(n37157), .Z(n37159) );
  NANDN U52095 ( .A(n37160), .B(n37159), .Z(n37161) );
  AND U52096 ( .A(n37162), .B(n37161), .Z(n37164) );
  NAND U52097 ( .A(n37164), .B(n37163), .Z(n37165) );
  NANDN U52098 ( .A(n37166), .B(n37165), .Z(n37167) );
  AND U52099 ( .A(n55171), .B(n37167), .Z(n37169) );
  AND U52100 ( .A(n37169), .B(n37168), .Z(n37173) );
  NAND U52101 ( .A(n37171), .B(n37170), .Z(n37172) );
  OR U52102 ( .A(n37173), .B(n37172), .Z(n37174) );
  AND U52103 ( .A(n37175), .B(n37174), .Z(n37179) );
  NAND U52104 ( .A(n37177), .B(n37176), .Z(n37178) );
  OR U52105 ( .A(n37179), .B(n37178), .Z(n37180) );
  AND U52106 ( .A(n37181), .B(n37180), .Z(n37185) );
  NAND U52107 ( .A(n37183), .B(n37182), .Z(n37184) );
  OR U52108 ( .A(n37185), .B(n37184), .Z(n37186) );
  AND U52109 ( .A(n37187), .B(n37186), .Z(n37191) );
  NAND U52110 ( .A(n37189), .B(n37188), .Z(n37190) );
  OR U52111 ( .A(n37191), .B(n37190), .Z(n37192) );
  AND U52112 ( .A(n37193), .B(n37192), .Z(n37197) );
  NAND U52113 ( .A(n37195), .B(n37194), .Z(n37196) );
  OR U52114 ( .A(n37197), .B(n37196), .Z(n37198) );
  AND U52115 ( .A(n37199), .B(n37198), .Z(n37203) );
  NAND U52116 ( .A(n37201), .B(n37200), .Z(n37202) );
  OR U52117 ( .A(n37203), .B(n37202), .Z(n37204) );
  AND U52118 ( .A(n37205), .B(n37204), .Z(n37209) );
  NAND U52119 ( .A(n37207), .B(n37206), .Z(n37208) );
  OR U52120 ( .A(n37209), .B(n37208), .Z(n37210) );
  AND U52121 ( .A(n37211), .B(n37210), .Z(n37212) );
  OR U52122 ( .A(n37213), .B(n37212), .Z(n37214) );
  NAND U52123 ( .A(n37215), .B(n37214), .Z(n37216) );
  AND U52124 ( .A(n37217), .B(n37216), .Z(n37218) );
  ANDN U52125 ( .B(n37219), .A(n37218), .Z(n37220) );
  OR U52126 ( .A(n37221), .B(n37220), .Z(n37222) );
  NAND U52127 ( .A(n37223), .B(n37222), .Z(n37224) );
  AND U52128 ( .A(n37225), .B(n37224), .Z(n37226) );
  OR U52129 ( .A(n37227), .B(n37226), .Z(n37228) );
  NAND U52130 ( .A(n37229), .B(n37228), .Z(n37230) );
  NANDN U52131 ( .A(n37231), .B(n37230), .Z(n37233) );
  OR U52132 ( .A(n37233), .B(n37232), .Z(n37234) );
  NAND U52133 ( .A(n37235), .B(n37234), .Z(n37239) );
  NAND U52134 ( .A(n37237), .B(n37236), .Z(n37238) );
  ANDN U52135 ( .B(n37239), .A(n37238), .Z(n37243) );
  NAND U52136 ( .A(n37241), .B(n37240), .Z(n37242) );
  OR U52137 ( .A(n37243), .B(n37242), .Z(n37244) );
  AND U52138 ( .A(n37245), .B(n37244), .Z(n37249) );
  NAND U52139 ( .A(n37247), .B(n37246), .Z(n37248) );
  OR U52140 ( .A(n37249), .B(n37248), .Z(n37250) );
  AND U52141 ( .A(n37251), .B(n37250), .Z(n37255) );
  NAND U52142 ( .A(n37253), .B(n37252), .Z(n37254) );
  OR U52143 ( .A(n37255), .B(n37254), .Z(n37256) );
  AND U52144 ( .A(n37257), .B(n37256), .Z(n37261) );
  NAND U52145 ( .A(n37259), .B(n37258), .Z(n37260) );
  OR U52146 ( .A(n37261), .B(n37260), .Z(n37262) );
  AND U52147 ( .A(n37263), .B(n37262), .Z(n37267) );
  NAND U52148 ( .A(n37265), .B(n37264), .Z(n37266) );
  OR U52149 ( .A(n37267), .B(n37266), .Z(n37268) );
  AND U52150 ( .A(n37269), .B(n37268), .Z(n37273) );
  NAND U52151 ( .A(n37271), .B(n37270), .Z(n37272) );
  OR U52152 ( .A(n37273), .B(n37272), .Z(n37274) );
  AND U52153 ( .A(n37275), .B(n37274), .Z(n37279) );
  NAND U52154 ( .A(n37277), .B(n37276), .Z(n37278) );
  OR U52155 ( .A(n37279), .B(n37278), .Z(n37280) );
  AND U52156 ( .A(n37281), .B(n37280), .Z(n37285) );
  NAND U52157 ( .A(n37283), .B(n37282), .Z(n37284) );
  OR U52158 ( .A(n37285), .B(n37284), .Z(n37286) );
  AND U52159 ( .A(n37287), .B(n37286), .Z(n37291) );
  NAND U52160 ( .A(n37289), .B(n37288), .Z(n37290) );
  OR U52161 ( .A(n37291), .B(n37290), .Z(n37292) );
  AND U52162 ( .A(n37293), .B(n37292), .Z(n37297) );
  NAND U52163 ( .A(n37295), .B(n37294), .Z(n37296) );
  OR U52164 ( .A(n37297), .B(n37296), .Z(n37298) );
  AND U52165 ( .A(n37299), .B(n37298), .Z(n37303) );
  NAND U52166 ( .A(n37301), .B(n37300), .Z(n37302) );
  OR U52167 ( .A(n37303), .B(n37302), .Z(n37304) );
  AND U52168 ( .A(n37305), .B(n37304), .Z(n37306) );
  ANDN U52169 ( .B(n37307), .A(n37306), .Z(n37308) );
  NAND U52170 ( .A(n37309), .B(n37308), .Z(n37310) );
  NANDN U52171 ( .A(n37311), .B(n37310), .Z(n37312) );
  OR U52172 ( .A(n51977), .B(n37312), .Z(n37313) );
  AND U52173 ( .A(n37314), .B(n37313), .Z(n37316) );
  NAND U52174 ( .A(n37316), .B(n37315), .Z(n37317) );
  NANDN U52175 ( .A(n37318), .B(n37317), .Z(n37319) );
  AND U52176 ( .A(n37320), .B(n37319), .Z(n37322) );
  NAND U52177 ( .A(n37322), .B(n37321), .Z(n37324) );
  ANDN U52178 ( .B(n37324), .A(n37323), .Z(n37325) );
  NANDN U52179 ( .A(n37326), .B(n37325), .Z(n37330) );
  NOR U52180 ( .A(n37328), .B(n37327), .Z(n37329) );
  NAND U52181 ( .A(n37330), .B(n37329), .Z(n37331) );
  AND U52182 ( .A(n37332), .B(n37331), .Z(n37334) );
  NAND U52183 ( .A(n37334), .B(n37333), .Z(n37335) );
  NANDN U52184 ( .A(n37336), .B(n37335), .Z(n37337) );
  AND U52185 ( .A(n37338), .B(n37337), .Z(n37340) );
  NAND U52186 ( .A(n37340), .B(n37339), .Z(n37341) );
  NANDN U52187 ( .A(n37342), .B(n37341), .Z(n37343) );
  AND U52188 ( .A(n37344), .B(n37343), .Z(n37346) );
  AND U52189 ( .A(n37346), .B(n37345), .Z(n37350) );
  NAND U52190 ( .A(n37348), .B(n37347), .Z(n37349) );
  OR U52191 ( .A(n37350), .B(n37349), .Z(n37351) );
  AND U52192 ( .A(n37352), .B(n37351), .Z(n37356) );
  NAND U52193 ( .A(n37354), .B(n37353), .Z(n37355) );
  OR U52194 ( .A(n37356), .B(n37355), .Z(n37357) );
  AND U52195 ( .A(n37358), .B(n37357), .Z(n37362) );
  NAND U52196 ( .A(n37360), .B(n37359), .Z(n37361) );
  OR U52197 ( .A(n37362), .B(n37361), .Z(n37363) );
  AND U52198 ( .A(n37364), .B(n37363), .Z(n37365) );
  NOR U52199 ( .A(n37366), .B(n37365), .Z(n37367) );
  NAND U52200 ( .A(n37368), .B(n37367), .Z(n37372) );
  NANDN U52201 ( .A(x[3030]), .B(y[3030]), .Z(n37370) );
  NAND U52202 ( .A(n37370), .B(n37369), .Z(n37371) );
  ANDN U52203 ( .B(n37372), .A(n37371), .Z(n37376) );
  NAND U52204 ( .A(n37374), .B(n37373), .Z(n37375) );
  OR U52205 ( .A(n37376), .B(n37375), .Z(n37377) );
  AND U52206 ( .A(n37378), .B(n37377), .Z(n37382) );
  NAND U52207 ( .A(n37380), .B(n37379), .Z(n37381) );
  OR U52208 ( .A(n37382), .B(n37381), .Z(n37383) );
  AND U52209 ( .A(n37384), .B(n37383), .Z(n37388) );
  NAND U52210 ( .A(n37386), .B(n37385), .Z(n37387) );
  OR U52211 ( .A(n37388), .B(n37387), .Z(n37389) );
  AND U52212 ( .A(n37390), .B(n37389), .Z(n37394) );
  NAND U52213 ( .A(n37392), .B(n37391), .Z(n37393) );
  OR U52214 ( .A(n37394), .B(n37393), .Z(n37395) );
  AND U52215 ( .A(n37395), .B(n55268), .Z(n37397) );
  AND U52216 ( .A(n37397), .B(n37396), .Z(n37398) );
  OR U52217 ( .A(n37399), .B(n37398), .Z(n37400) );
  NAND U52218 ( .A(n37401), .B(n37400), .Z(n37402) );
  AND U52219 ( .A(n37403), .B(n37402), .Z(n37404) );
  OR U52220 ( .A(n37405), .B(n37404), .Z(n37406) );
  NANDN U52221 ( .A(n37407), .B(n37406), .Z(n37408) );
  AND U52222 ( .A(n37408), .B(n55277), .Z(n37409) );
  OR U52223 ( .A(n37410), .B(n37409), .Z(n37411) );
  NAND U52224 ( .A(n55279), .B(n37411), .Z(n37412) );
  NANDN U52225 ( .A(n37413), .B(n37412), .Z(n37414) );
  OR U52226 ( .A(n37415), .B(n37414), .Z(n37416) );
  AND U52227 ( .A(n37417), .B(n37416), .Z(n37418) );
  NANDN U52228 ( .A(x[3046]), .B(y[3046]), .Z(n55280) );
  AND U52229 ( .A(n37418), .B(n55280), .Z(n37419) );
  OR U52230 ( .A(n37420), .B(n37419), .Z(n37421) );
  NAND U52231 ( .A(n37422), .B(n37421), .Z(n37423) );
  NANDN U52232 ( .A(n37424), .B(n37423), .Z(n37426) );
  NAND U52233 ( .A(n37426), .B(n37425), .Z(n37427) );
  ANDN U52234 ( .B(y[3050]), .A(x[3050]), .Z(n55285) );
  OR U52235 ( .A(n37427), .B(n55285), .Z(n37428) );
  NAND U52236 ( .A(n37429), .B(n37428), .Z(n37430) );
  NANDN U52237 ( .A(n37431), .B(n37430), .Z(n37433) );
  OR U52238 ( .A(n37433), .B(n37432), .Z(n37434) );
  NANDN U52239 ( .A(n37435), .B(n37434), .Z(n37436) );
  AND U52240 ( .A(n37437), .B(n37436), .Z(n37441) );
  NAND U52241 ( .A(n37439), .B(n37438), .Z(n37440) );
  OR U52242 ( .A(n37441), .B(n37440), .Z(n37442) );
  AND U52243 ( .A(n37443), .B(n37442), .Z(n37447) );
  NAND U52244 ( .A(n37445), .B(n37444), .Z(n37446) );
  OR U52245 ( .A(n37447), .B(n37446), .Z(n37448) );
  AND U52246 ( .A(n37449), .B(n37448), .Z(n37453) );
  NAND U52247 ( .A(n37451), .B(n37450), .Z(n37452) );
  OR U52248 ( .A(n37453), .B(n37452), .Z(n37454) );
  AND U52249 ( .A(n37455), .B(n37454), .Z(n37459) );
  NAND U52250 ( .A(n37457), .B(n37456), .Z(n37458) );
  OR U52251 ( .A(n37459), .B(n37458), .Z(n37460) );
  AND U52252 ( .A(n37461), .B(n37460), .Z(n37465) );
  NAND U52253 ( .A(n37463), .B(n37462), .Z(n37464) );
  OR U52254 ( .A(n37465), .B(n37464), .Z(n37466) );
  AND U52255 ( .A(n37467), .B(n37466), .Z(n37468) );
  OR U52256 ( .A(n37469), .B(n37468), .Z(n37470) );
  NAND U52257 ( .A(n37471), .B(n37470), .Z(n37472) );
  NAND U52258 ( .A(n37473), .B(n37472), .Z(n37474) );
  NANDN U52259 ( .A(n37475), .B(n37474), .Z(n37476) );
  AND U52260 ( .A(n37477), .B(n37476), .Z(n37479) );
  NAND U52261 ( .A(n37479), .B(n37478), .Z(n37480) );
  NANDN U52262 ( .A(n37481), .B(n37480), .Z(n37482) );
  AND U52263 ( .A(n37483), .B(n37482), .Z(n37485) );
  NAND U52264 ( .A(n37485), .B(n37484), .Z(n37486) );
  NANDN U52265 ( .A(n37487), .B(n37486), .Z(n37488) );
  AND U52266 ( .A(n37489), .B(n37488), .Z(n37491) );
  NAND U52267 ( .A(n37491), .B(n37490), .Z(n37492) );
  NANDN U52268 ( .A(n37493), .B(n37492), .Z(n37494) );
  AND U52269 ( .A(n37495), .B(n37494), .Z(n37497) );
  NAND U52270 ( .A(n37497), .B(n37496), .Z(n37498) );
  NANDN U52271 ( .A(n37499), .B(n37498), .Z(n37500) );
  ANDN U52272 ( .B(y[3076]), .A(x[3076]), .Z(n55307) );
  OR U52273 ( .A(n37500), .B(n55307), .Z(n37501) );
  NAND U52274 ( .A(n37502), .B(n37501), .Z(n37503) );
  NANDN U52275 ( .A(n55311), .B(n37503), .Z(n37505) );
  OR U52276 ( .A(n37505), .B(n37504), .Z(n37506) );
  NANDN U52277 ( .A(n37507), .B(n37506), .Z(n37508) );
  AND U52278 ( .A(n37509), .B(n37508), .Z(n37513) );
  NAND U52279 ( .A(n37511), .B(n37510), .Z(n37512) );
  OR U52280 ( .A(n37513), .B(n37512), .Z(n37514) );
  AND U52281 ( .A(n37515), .B(n37514), .Z(n37519) );
  NAND U52282 ( .A(n37517), .B(n37516), .Z(n37518) );
  OR U52283 ( .A(n37519), .B(n37518), .Z(n37520) );
  AND U52284 ( .A(n37521), .B(n37520), .Z(n37525) );
  NAND U52285 ( .A(n37523), .B(n37522), .Z(n37524) );
  OR U52286 ( .A(n37525), .B(n37524), .Z(n37526) );
  AND U52287 ( .A(n37527), .B(n37526), .Z(n37531) );
  AND U52288 ( .A(n37529), .B(n37528), .Z(n37530) );
  NANDN U52289 ( .A(n37531), .B(n37530), .Z(n37532) );
  NANDN U52290 ( .A(n37533), .B(n37532), .Z(n37534) );
  AND U52291 ( .A(n37535), .B(n37534), .Z(n37537) );
  NAND U52292 ( .A(n37537), .B(n37536), .Z(n37538) );
  NANDN U52293 ( .A(n37539), .B(n37538), .Z(n37540) );
  AND U52294 ( .A(n37541), .B(n37540), .Z(n37543) );
  NAND U52295 ( .A(n37543), .B(n37542), .Z(n37544) );
  NANDN U52296 ( .A(n37545), .B(n37544), .Z(n37546) );
  AND U52297 ( .A(n37547), .B(n37546), .Z(n37549) );
  NAND U52298 ( .A(n37549), .B(n37548), .Z(n37550) );
  NANDN U52299 ( .A(n37551), .B(n37550), .Z(n37552) );
  AND U52300 ( .A(n37553), .B(n37552), .Z(n37555) );
  AND U52301 ( .A(n37555), .B(n37554), .Z(n37559) );
  NAND U52302 ( .A(n37557), .B(n37556), .Z(n37558) );
  OR U52303 ( .A(n37559), .B(n37558), .Z(n37560) );
  AND U52304 ( .A(n37561), .B(n37560), .Z(n37562) );
  OR U52305 ( .A(n37563), .B(n37562), .Z(n37564) );
  NAND U52306 ( .A(n37565), .B(n37564), .Z(n37566) );
  AND U52307 ( .A(n37567), .B(n37566), .Z(n37568) );
  NOR U52308 ( .A(n37569), .B(n37568), .Z(n37571) );
  NAND U52309 ( .A(n37571), .B(n37570), .Z(n37575) );
  NANDN U52310 ( .A(x[3102]), .B(y[3102]), .Z(n37572) );
  AND U52311 ( .A(n37573), .B(n37572), .Z(n37574) );
  NAND U52312 ( .A(n37575), .B(n37574), .Z(n37576) );
  NANDN U52313 ( .A(n37577), .B(n37576), .Z(n37578) );
  NAND U52314 ( .A(n37579), .B(n37578), .Z(n37580) );
  NANDN U52315 ( .A(n37581), .B(n37580), .Z(n37582) );
  AND U52316 ( .A(n37583), .B(n37582), .Z(n37585) );
  NAND U52317 ( .A(n37585), .B(n37584), .Z(n37586) );
  NANDN U52318 ( .A(n37587), .B(n37586), .Z(n37588) );
  AND U52319 ( .A(n37589), .B(n37588), .Z(n37591) );
  NAND U52320 ( .A(n37591), .B(n37590), .Z(n37592) );
  NANDN U52321 ( .A(n37593), .B(n37592), .Z(n37594) );
  AND U52322 ( .A(n37595), .B(n37594), .Z(n37596) );
  NANDN U52323 ( .A(n37597), .B(n37596), .Z(n37598) );
  NAND U52324 ( .A(n37599), .B(n37598), .Z(n37600) );
  NANDN U52325 ( .A(n37601), .B(n37600), .Z(n37602) );
  NAND U52326 ( .A(n37603), .B(n37602), .Z(n37604) );
  NANDN U52327 ( .A(n37605), .B(n37604), .Z(n37606) );
  AND U52328 ( .A(n37607), .B(n37606), .Z(n37608) );
  NAND U52329 ( .A(n37608), .B(n55370), .Z(n37612) );
  AND U52330 ( .A(n37610), .B(n37609), .Z(n37611) );
  ANDN U52331 ( .B(n37612), .A(n37611), .Z(n37613) );
  NANDN U52332 ( .A(n55371), .B(n37613), .Z(n37614) );
  AND U52333 ( .A(n37615), .B(n37614), .Z(n37617) );
  XNOR U52334 ( .A(x[3119]), .B(y[3119]), .Z(n37616) );
  NANDN U52335 ( .A(n37617), .B(n37616), .Z(n37618) );
  AND U52336 ( .A(n37619), .B(n37618), .Z(n37620) );
  OR U52337 ( .A(n37621), .B(n37620), .Z(n37622) );
  NAND U52338 ( .A(n37623), .B(n37622), .Z(n37624) );
  NAND U52339 ( .A(n37625), .B(n37624), .Z(n37626) );
  NANDN U52340 ( .A(n37627), .B(n37626), .Z(n37628) );
  AND U52341 ( .A(n37629), .B(n37628), .Z(n37631) );
  NAND U52342 ( .A(n37631), .B(n37630), .Z(n37632) );
  NANDN U52343 ( .A(n37633), .B(n37632), .Z(n37634) );
  AND U52344 ( .A(n37635), .B(n37634), .Z(n37637) );
  NAND U52345 ( .A(n37637), .B(n37636), .Z(n37638) );
  NANDN U52346 ( .A(n37639), .B(n37638), .Z(n37640) );
  AND U52347 ( .A(n37641), .B(n37640), .Z(n37643) );
  AND U52348 ( .A(n37643), .B(n37642), .Z(n37647) );
  NAND U52349 ( .A(n37645), .B(n37644), .Z(n37646) );
  OR U52350 ( .A(n37647), .B(n37646), .Z(n37648) );
  AND U52351 ( .A(n37649), .B(n37648), .Z(n37653) );
  NAND U52352 ( .A(n37651), .B(n37650), .Z(n37652) );
  OR U52353 ( .A(n37653), .B(n37652), .Z(n37654) );
  AND U52354 ( .A(n37655), .B(n37654), .Z(n37659) );
  NAND U52355 ( .A(n37657), .B(n37656), .Z(n37658) );
  OR U52356 ( .A(n37659), .B(n37658), .Z(n37660) );
  AND U52357 ( .A(n37661), .B(n37660), .Z(n37665) );
  NAND U52358 ( .A(n37663), .B(n37662), .Z(n37664) );
  OR U52359 ( .A(n37665), .B(n37664), .Z(n37666) );
  AND U52360 ( .A(n37667), .B(n37666), .Z(n37671) );
  NAND U52361 ( .A(n37669), .B(n37668), .Z(n37670) );
  OR U52362 ( .A(n37671), .B(n37670), .Z(n37672) );
  AND U52363 ( .A(n37673), .B(n37672), .Z(n37674) );
  OR U52364 ( .A(n37675), .B(n37674), .Z(n37676) );
  NAND U52365 ( .A(n37677), .B(n37676), .Z(n37678) );
  AND U52366 ( .A(n37679), .B(n37678), .Z(n37680) );
  ANDN U52367 ( .B(n37681), .A(n37680), .Z(n37685) );
  NAND U52368 ( .A(n37683), .B(n37682), .Z(n37684) );
  OR U52369 ( .A(n37685), .B(n37684), .Z(n37686) );
  AND U52370 ( .A(n37687), .B(n37686), .Z(n37691) );
  NAND U52371 ( .A(n37689), .B(n37688), .Z(n37690) );
  OR U52372 ( .A(n37691), .B(n37690), .Z(n37692) );
  AND U52373 ( .A(n37693), .B(n37692), .Z(n37697) );
  NAND U52374 ( .A(n37695), .B(n37694), .Z(n37696) );
  OR U52375 ( .A(n37697), .B(n37696), .Z(n37698) );
  AND U52376 ( .A(n37699), .B(n37698), .Z(n37703) );
  NAND U52377 ( .A(n37701), .B(n37700), .Z(n37702) );
  OR U52378 ( .A(n37703), .B(n37702), .Z(n37704) );
  AND U52379 ( .A(n37705), .B(n37704), .Z(n37706) );
  NOR U52380 ( .A(n37707), .B(n37706), .Z(n37708) );
  NAND U52381 ( .A(n37709), .B(n37708), .Z(n37713) );
  NAND U52382 ( .A(n37711), .B(n37710), .Z(n37712) );
  ANDN U52383 ( .B(n37713), .A(n37712), .Z(n37717) );
  NAND U52384 ( .A(n37715), .B(n37714), .Z(n37716) );
  OR U52385 ( .A(n37717), .B(n37716), .Z(n37718) );
  AND U52386 ( .A(n37719), .B(n37718), .Z(n37723) );
  NAND U52387 ( .A(n37721), .B(n37720), .Z(n37722) );
  OR U52388 ( .A(n37723), .B(n37722), .Z(n37724) );
  AND U52389 ( .A(n37725), .B(n37724), .Z(n37729) );
  NAND U52390 ( .A(n37727), .B(n37726), .Z(n37728) );
  OR U52391 ( .A(n37729), .B(n37728), .Z(n37730) );
  AND U52392 ( .A(n37731), .B(n37730), .Z(n37735) );
  NAND U52393 ( .A(n37733), .B(n37732), .Z(n37734) );
  OR U52394 ( .A(n37735), .B(n37734), .Z(n37736) );
  AND U52395 ( .A(n37737), .B(n37736), .Z(n37738) );
  OR U52396 ( .A(n37739), .B(n37738), .Z(n37740) );
  NAND U52397 ( .A(n37741), .B(n37740), .Z(n37742) );
  AND U52398 ( .A(n37743), .B(n37742), .Z(n37744) );
  NOR U52399 ( .A(n55420), .B(n37744), .Z(n37745) );
  NANDN U52400 ( .A(n37746), .B(n37745), .Z(n37747) );
  AND U52401 ( .A(n37748), .B(n37747), .Z(n37750) );
  NAND U52402 ( .A(n37750), .B(n37749), .Z(n37751) );
  NANDN U52403 ( .A(n37752), .B(n37751), .Z(n37753) );
  AND U52404 ( .A(n37754), .B(n37753), .Z(n37756) );
  NAND U52405 ( .A(n37756), .B(n37755), .Z(n37757) );
  NANDN U52406 ( .A(n37758), .B(n37757), .Z(n37759) );
  AND U52407 ( .A(n37760), .B(n37759), .Z(n37762) );
  AND U52408 ( .A(n37762), .B(n37761), .Z(n37766) );
  NAND U52409 ( .A(n37764), .B(n37763), .Z(n37765) );
  OR U52410 ( .A(n37766), .B(n37765), .Z(n37767) );
  AND U52411 ( .A(n37768), .B(n37767), .Z(n37772) );
  NAND U52412 ( .A(n37770), .B(n37769), .Z(n37771) );
  OR U52413 ( .A(n37772), .B(n37771), .Z(n37773) );
  AND U52414 ( .A(n37774), .B(n37773), .Z(n37778) );
  NAND U52415 ( .A(n37776), .B(n37775), .Z(n37777) );
  OR U52416 ( .A(n37778), .B(n37777), .Z(n37779) );
  AND U52417 ( .A(n37780), .B(n37779), .Z(n37781) );
  OR U52418 ( .A(n37782), .B(n37781), .Z(n37783) );
  NAND U52419 ( .A(n37784), .B(n37783), .Z(n37785) );
  NANDN U52420 ( .A(n37786), .B(n37785), .Z(n37788) );
  ANDN U52421 ( .B(y[3178]), .A(x[3178]), .Z(n37787) );
  OR U52422 ( .A(n37788), .B(n37787), .Z(n37789) );
  NAND U52423 ( .A(n37790), .B(n37789), .Z(n37791) );
  AND U52424 ( .A(n37792), .B(n37791), .Z(n37793) );
  OR U52425 ( .A(n37794), .B(n37793), .Z(n37795) );
  NAND U52426 ( .A(n37796), .B(n37795), .Z(n37800) );
  NAND U52427 ( .A(n37798), .B(n37797), .Z(n37799) );
  ANDN U52428 ( .B(n37800), .A(n37799), .Z(n37804) );
  NAND U52429 ( .A(n37802), .B(n37801), .Z(n37803) );
  OR U52430 ( .A(n37804), .B(n37803), .Z(n37805) );
  AND U52431 ( .A(n37806), .B(n37805), .Z(n37810) );
  NAND U52432 ( .A(n37808), .B(n37807), .Z(n37809) );
  OR U52433 ( .A(n37810), .B(n37809), .Z(n37811) );
  AND U52434 ( .A(n37812), .B(n37811), .Z(n37813) );
  OR U52435 ( .A(n37814), .B(n37813), .Z(n37815) );
  NAND U52436 ( .A(n37816), .B(n37815), .Z(n37819) );
  NANDN U52437 ( .A(x[3190]), .B(y[3190]), .Z(n51957) );
  IV U52438 ( .A(n37817), .Z(n55445) );
  AND U52439 ( .A(n51957), .B(n55445), .Z(n37818) );
  NAND U52440 ( .A(n37819), .B(n37818), .Z(n37820) );
  NANDN U52441 ( .A(n37821), .B(n37820), .Z(n37822) );
  AND U52442 ( .A(n37823), .B(n37822), .Z(n37826) );
  NAND U52443 ( .A(n51954), .B(n37824), .Z(n37825) );
  OR U52444 ( .A(n37826), .B(n37825), .Z(n37827) );
  AND U52445 ( .A(n37828), .B(n37827), .Z(n37830) );
  NAND U52446 ( .A(n37830), .B(n37829), .Z(n37831) );
  NANDN U52447 ( .A(n37832), .B(n37831), .Z(n37833) );
  AND U52448 ( .A(n37834), .B(n37833), .Z(n37836) );
  NAND U52449 ( .A(n37836), .B(n37835), .Z(n37837) );
  NANDN U52450 ( .A(n37838), .B(n37837), .Z(n37839) );
  AND U52451 ( .A(n37840), .B(n37839), .Z(n37844) );
  NAND U52452 ( .A(n37842), .B(n37841), .Z(n37843) );
  OR U52453 ( .A(n37844), .B(n37843), .Z(n37845) );
  AND U52454 ( .A(n37846), .B(n37845), .Z(n37850) );
  NAND U52455 ( .A(n37848), .B(n37847), .Z(n37849) );
  OR U52456 ( .A(n37850), .B(n37849), .Z(n37851) );
  AND U52457 ( .A(n37852), .B(n37851), .Z(n37856) );
  NAND U52458 ( .A(n37854), .B(n37853), .Z(n37855) );
  OR U52459 ( .A(n37856), .B(n37855), .Z(n37857) );
  AND U52460 ( .A(n37858), .B(n37857), .Z(n37862) );
  NAND U52461 ( .A(n37860), .B(n37859), .Z(n37861) );
  OR U52462 ( .A(n37862), .B(n37861), .Z(n37863) );
  AND U52463 ( .A(n37864), .B(n37863), .Z(n37868) );
  NAND U52464 ( .A(n37866), .B(n37865), .Z(n37867) );
  OR U52465 ( .A(n37868), .B(n37867), .Z(n37869) );
  AND U52466 ( .A(n37870), .B(n37869), .Z(n37874) );
  NAND U52467 ( .A(n37872), .B(n37871), .Z(n37873) );
  OR U52468 ( .A(n37874), .B(n37873), .Z(n37875) );
  AND U52469 ( .A(n37876), .B(n37875), .Z(n37880) );
  NAND U52470 ( .A(n37878), .B(n37877), .Z(n37879) );
  OR U52471 ( .A(n37880), .B(n37879), .Z(n37881) );
  AND U52472 ( .A(n37882), .B(n37881), .Z(n37886) );
  NAND U52473 ( .A(n37884), .B(n37883), .Z(n37885) );
  OR U52474 ( .A(n37886), .B(n37885), .Z(n37887) );
  AND U52475 ( .A(n37888), .B(n37887), .Z(n37892) );
  NAND U52476 ( .A(n37890), .B(n37889), .Z(n37891) );
  OR U52477 ( .A(n37892), .B(n37891), .Z(n37893) );
  AND U52478 ( .A(n37894), .B(n37893), .Z(n37898) );
  NAND U52479 ( .A(n37896), .B(n37895), .Z(n37897) );
  OR U52480 ( .A(n37898), .B(n37897), .Z(n37899) );
  AND U52481 ( .A(n37900), .B(n37899), .Z(n37904) );
  AND U52482 ( .A(n37902), .B(n37901), .Z(n37903) );
  NANDN U52483 ( .A(n37904), .B(n37903), .Z(n37905) );
  AND U52484 ( .A(n37906), .B(n37905), .Z(n37910) );
  NAND U52485 ( .A(n37908), .B(n37907), .Z(n37909) );
  OR U52486 ( .A(n37910), .B(n37909), .Z(n37911) );
  AND U52487 ( .A(n37912), .B(n37911), .Z(n37916) );
  NAND U52488 ( .A(n37914), .B(n37913), .Z(n37915) );
  OR U52489 ( .A(n37916), .B(n37915), .Z(n37917) );
  AND U52490 ( .A(n37918), .B(n37917), .Z(n37922) );
  NAND U52491 ( .A(n37920), .B(n37919), .Z(n37921) );
  OR U52492 ( .A(n37922), .B(n37921), .Z(n37923) );
  AND U52493 ( .A(n37924), .B(n37923), .Z(n37928) );
  NAND U52494 ( .A(n37926), .B(n37925), .Z(n37927) );
  OR U52495 ( .A(n37928), .B(n37927), .Z(n37929) );
  AND U52496 ( .A(n37930), .B(n37929), .Z(n37931) );
  OR U52497 ( .A(n37932), .B(n37931), .Z(n37933) );
  NAND U52498 ( .A(n37934), .B(n37933), .Z(n37935) );
  AND U52499 ( .A(n37936), .B(n37935), .Z(n37937) );
  NOR U52500 ( .A(n55480), .B(n37937), .Z(n37938) );
  NANDN U52501 ( .A(n37939), .B(n37938), .Z(n37940) );
  AND U52502 ( .A(n37941), .B(n37940), .Z(n37943) );
  NAND U52503 ( .A(n37943), .B(n37942), .Z(n37944) );
  NANDN U52504 ( .A(n37945), .B(n37944), .Z(n37946) );
  AND U52505 ( .A(n37947), .B(n37946), .Z(n37949) );
  NAND U52506 ( .A(n37949), .B(n37948), .Z(n37950) );
  NANDN U52507 ( .A(n37951), .B(n37950), .Z(n37952) );
  AND U52508 ( .A(n37953), .B(n37952), .Z(n37955) );
  NAND U52509 ( .A(n37955), .B(n37954), .Z(n37956) );
  NANDN U52510 ( .A(n37957), .B(n37956), .Z(n37958) );
  AND U52511 ( .A(n37959), .B(n37958), .Z(n37961) );
  AND U52512 ( .A(n37961), .B(n37960), .Z(n37965) );
  NAND U52513 ( .A(n37963), .B(n37962), .Z(n37964) );
  OR U52514 ( .A(n37965), .B(n37964), .Z(n37966) );
  AND U52515 ( .A(n37967), .B(n37966), .Z(n37971) );
  NAND U52516 ( .A(n37969), .B(n37968), .Z(n37970) );
  OR U52517 ( .A(n37971), .B(n37970), .Z(n37972) );
  AND U52518 ( .A(n37973), .B(n37972), .Z(n37974) );
  NOR U52519 ( .A(n37975), .B(n37974), .Z(n37976) );
  NAND U52520 ( .A(n37977), .B(n37976), .Z(n37978) );
  NANDN U52521 ( .A(n37979), .B(n37978), .Z(n37980) );
  NAND U52522 ( .A(n37981), .B(n37980), .Z(n37982) );
  NANDN U52523 ( .A(n37983), .B(n37982), .Z(n37984) );
  AND U52524 ( .A(n37985), .B(n37984), .Z(n37987) );
  NAND U52525 ( .A(n37987), .B(n37986), .Z(n37988) );
  NANDN U52526 ( .A(n37989), .B(n37988), .Z(n37990) );
  AND U52527 ( .A(n37991), .B(n37990), .Z(n37993) );
  NAND U52528 ( .A(n37993), .B(n37992), .Z(n37994) );
  NANDN U52529 ( .A(n37995), .B(n37994), .Z(n37996) );
  AND U52530 ( .A(n37997), .B(n37996), .Z(n37999) );
  NANDN U52531 ( .A(x[3252]), .B(y[3252]), .Z(n37998) );
  AND U52532 ( .A(n37999), .B(n37998), .Z(n38003) );
  NAND U52533 ( .A(n38001), .B(n38000), .Z(n38002) );
  OR U52534 ( .A(n38003), .B(n38002), .Z(n38004) );
  AND U52535 ( .A(n38005), .B(n38004), .Z(n38009) );
  NAND U52536 ( .A(n38007), .B(n38006), .Z(n38008) );
  OR U52537 ( .A(n38009), .B(n38008), .Z(n38010) );
  AND U52538 ( .A(n38011), .B(n38010), .Z(n38015) );
  NAND U52539 ( .A(n38013), .B(n38012), .Z(n38014) );
  OR U52540 ( .A(n38015), .B(n38014), .Z(n38016) );
  AND U52541 ( .A(n38017), .B(n38016), .Z(n38021) );
  NAND U52542 ( .A(n38019), .B(n38018), .Z(n38020) );
  OR U52543 ( .A(n38021), .B(n38020), .Z(n38022) );
  AND U52544 ( .A(n38023), .B(n38022), .Z(n38027) );
  NAND U52545 ( .A(n38025), .B(n38024), .Z(n38026) );
  OR U52546 ( .A(n38027), .B(n38026), .Z(n38028) );
  AND U52547 ( .A(n38029), .B(n38028), .Z(n38033) );
  NAND U52548 ( .A(n38031), .B(n38030), .Z(n38032) );
  OR U52549 ( .A(n38033), .B(n38032), .Z(n38034) );
  AND U52550 ( .A(n38035), .B(n38034), .Z(n38039) );
  NAND U52551 ( .A(n38037), .B(n38036), .Z(n38038) );
  OR U52552 ( .A(n38039), .B(n38038), .Z(n38040) );
  AND U52553 ( .A(n38041), .B(n38040), .Z(n38042) );
  OR U52554 ( .A(n38043), .B(n38042), .Z(n38044) );
  NAND U52555 ( .A(n38045), .B(n38044), .Z(n38046) );
  AND U52556 ( .A(n38047), .B(n38046), .Z(n38048) );
  OR U52557 ( .A(n38049), .B(n38048), .Z(n38050) );
  NAND U52558 ( .A(n38051), .B(n38050), .Z(n38055) );
  NAND U52559 ( .A(n38053), .B(n38052), .Z(n38054) );
  ANDN U52560 ( .B(n38055), .A(n38054), .Z(n38059) );
  NAND U52561 ( .A(n38057), .B(n38056), .Z(n38058) );
  OR U52562 ( .A(n38059), .B(n38058), .Z(n38060) );
  AND U52563 ( .A(n38061), .B(n38060), .Z(n38065) );
  NAND U52564 ( .A(n38063), .B(n38062), .Z(n38064) );
  OR U52565 ( .A(n38065), .B(n38064), .Z(n38066) );
  AND U52566 ( .A(n38067), .B(n38066), .Z(n38071) );
  NAND U52567 ( .A(n38069), .B(n38068), .Z(n38070) );
  OR U52568 ( .A(n38071), .B(n38070), .Z(n38072) );
  AND U52569 ( .A(n38073), .B(n38072), .Z(n38077) );
  NAND U52570 ( .A(n38075), .B(n38074), .Z(n38076) );
  OR U52571 ( .A(n38077), .B(n38076), .Z(n38078) );
  AND U52572 ( .A(n38079), .B(n38078), .Z(n38083) );
  NAND U52573 ( .A(n38081), .B(n38080), .Z(n38082) );
  OR U52574 ( .A(n38083), .B(n38082), .Z(n38084) );
  AND U52575 ( .A(n38085), .B(n38084), .Z(n38089) );
  NAND U52576 ( .A(n38087), .B(n38086), .Z(n38088) );
  OR U52577 ( .A(n38089), .B(n38088), .Z(n38090) );
  AND U52578 ( .A(n38091), .B(n38090), .Z(n38095) );
  NAND U52579 ( .A(n38093), .B(n38092), .Z(n38094) );
  OR U52580 ( .A(n38095), .B(n38094), .Z(n38096) );
  AND U52581 ( .A(n38097), .B(n38096), .Z(n38101) );
  NAND U52582 ( .A(n38099), .B(n38098), .Z(n38100) );
  OR U52583 ( .A(n38101), .B(n38100), .Z(n38102) );
  AND U52584 ( .A(n38103), .B(n38102), .Z(n38107) );
  NAND U52585 ( .A(n38105), .B(n38104), .Z(n38106) );
  OR U52586 ( .A(n38107), .B(n38106), .Z(n38108) );
  AND U52587 ( .A(n38109), .B(n38108), .Z(n38113) );
  NAND U52588 ( .A(n38111), .B(n38110), .Z(n38112) );
  OR U52589 ( .A(n38113), .B(n38112), .Z(n38114) );
  AND U52590 ( .A(n38115), .B(n38114), .Z(n38119) );
  NAND U52591 ( .A(n38117), .B(n38116), .Z(n38118) );
  OR U52592 ( .A(n38119), .B(n38118), .Z(n38120) );
  AND U52593 ( .A(n38121), .B(n38120), .Z(n38125) );
  NAND U52594 ( .A(n38123), .B(n38122), .Z(n38124) );
  OR U52595 ( .A(n38125), .B(n38124), .Z(n38126) );
  AND U52596 ( .A(n38127), .B(n38126), .Z(n38131) );
  NAND U52597 ( .A(n38129), .B(n38128), .Z(n38130) );
  OR U52598 ( .A(n38131), .B(n38130), .Z(n38132) );
  AND U52599 ( .A(n38133), .B(n38132), .Z(n38137) );
  NAND U52600 ( .A(n38135), .B(n38134), .Z(n38136) );
  OR U52601 ( .A(n38137), .B(n38136), .Z(n38138) );
  AND U52602 ( .A(n38139), .B(n38138), .Z(n38143) );
  NAND U52603 ( .A(n38141), .B(n38140), .Z(n38142) );
  OR U52604 ( .A(n38143), .B(n38142), .Z(n38144) );
  AND U52605 ( .A(n38145), .B(n38144), .Z(n38149) );
  NAND U52606 ( .A(n38147), .B(n38146), .Z(n38148) );
  OR U52607 ( .A(n38149), .B(n38148), .Z(n38150) );
  AND U52608 ( .A(n38151), .B(n38150), .Z(n38155) );
  NAND U52609 ( .A(n38153), .B(n38152), .Z(n38154) );
  OR U52610 ( .A(n38155), .B(n38154), .Z(n38156) );
  AND U52611 ( .A(n38157), .B(n38156), .Z(n38161) );
  NAND U52612 ( .A(n38159), .B(n38158), .Z(n38160) );
  OR U52613 ( .A(n38161), .B(n38160), .Z(n38162) );
  AND U52614 ( .A(n38163), .B(n38162), .Z(n38167) );
  NAND U52615 ( .A(n38165), .B(n38164), .Z(n38166) );
  OR U52616 ( .A(n38167), .B(n38166), .Z(n38168) );
  AND U52617 ( .A(n38169), .B(n38168), .Z(n38173) );
  NAND U52618 ( .A(n38171), .B(n38170), .Z(n38172) );
  OR U52619 ( .A(n38173), .B(n38172), .Z(n38174) );
  AND U52620 ( .A(n38175), .B(n38174), .Z(n38179) );
  NAND U52621 ( .A(n38177), .B(n38176), .Z(n38178) );
  OR U52622 ( .A(n38179), .B(n38178), .Z(n38180) );
  AND U52623 ( .A(n38181), .B(n38180), .Z(n38185) );
  NAND U52624 ( .A(n38183), .B(n38182), .Z(n38184) );
  OR U52625 ( .A(n38185), .B(n38184), .Z(n38186) );
  AND U52626 ( .A(n38187), .B(n38186), .Z(n38191) );
  NAND U52627 ( .A(n38189), .B(n38188), .Z(n38190) );
  OR U52628 ( .A(n38191), .B(n38190), .Z(n38192) );
  AND U52629 ( .A(n38193), .B(n38192), .Z(n38197) );
  NAND U52630 ( .A(n38195), .B(n38194), .Z(n38196) );
  OR U52631 ( .A(n38197), .B(n38196), .Z(n38198) );
  AND U52632 ( .A(n38199), .B(n38198), .Z(n38203) );
  NAND U52633 ( .A(n38201), .B(n38200), .Z(n38202) );
  OR U52634 ( .A(n38203), .B(n38202), .Z(n38204) );
  AND U52635 ( .A(n38205), .B(n38204), .Z(n38209) );
  NAND U52636 ( .A(n38207), .B(n38206), .Z(n38208) );
  OR U52637 ( .A(n38209), .B(n38208), .Z(n38210) );
  AND U52638 ( .A(n38211), .B(n38210), .Z(n38212) );
  NOR U52639 ( .A(n38213), .B(n38212), .Z(n38214) );
  NAND U52640 ( .A(n38215), .B(n38214), .Z(n38219) );
  NAND U52641 ( .A(n38217), .B(n38216), .Z(n38218) );
  ANDN U52642 ( .B(n38219), .A(n38218), .Z(n38223) );
  NAND U52643 ( .A(n38221), .B(n38220), .Z(n38222) );
  OR U52644 ( .A(n38223), .B(n38222), .Z(n38224) );
  AND U52645 ( .A(n38225), .B(n38224), .Z(n38229) );
  NAND U52646 ( .A(n38227), .B(n38226), .Z(n38228) );
  OR U52647 ( .A(n38229), .B(n38228), .Z(n38230) );
  AND U52648 ( .A(n38231), .B(n38230), .Z(n38235) );
  NAND U52649 ( .A(n38233), .B(n38232), .Z(n38234) );
  OR U52650 ( .A(n38235), .B(n38234), .Z(n38236) );
  AND U52651 ( .A(n38237), .B(n38236), .Z(n38241) );
  NAND U52652 ( .A(n38239), .B(n38238), .Z(n38240) );
  OR U52653 ( .A(n38241), .B(n38240), .Z(n38242) );
  AND U52654 ( .A(n38243), .B(n38242), .Z(n38247) );
  NAND U52655 ( .A(n38245), .B(n38244), .Z(n38246) );
  OR U52656 ( .A(n38247), .B(n38246), .Z(n38248) );
  AND U52657 ( .A(n38249), .B(n38248), .Z(n38253) );
  NAND U52658 ( .A(n38251), .B(n38250), .Z(n38252) );
  OR U52659 ( .A(n38253), .B(n38252), .Z(n38254) );
  AND U52660 ( .A(n38255), .B(n38254), .Z(n38256) );
  OR U52661 ( .A(n38257), .B(n38256), .Z(n38258) );
  NAND U52662 ( .A(n38259), .B(n38258), .Z(n38260) );
  NAND U52663 ( .A(n38261), .B(n38260), .Z(n38262) );
  NANDN U52664 ( .A(n38263), .B(n38262), .Z(n38264) );
  AND U52665 ( .A(n55573), .B(n38264), .Z(n38266) );
  NAND U52666 ( .A(n38266), .B(n38265), .Z(n38267) );
  NANDN U52667 ( .A(n38268), .B(n38267), .Z(n38269) );
  AND U52668 ( .A(n38270), .B(n38269), .Z(n38271) );
  NANDN U52669 ( .A(n55574), .B(n38271), .Z(n38272) );
  NAND U52670 ( .A(n38273), .B(n38272), .Z(n38274) );
  NANDN U52671 ( .A(n38275), .B(n38274), .Z(n38276) );
  AND U52672 ( .A(n38277), .B(n38276), .Z(n38278) );
  NAND U52673 ( .A(n38279), .B(n38278), .Z(n38280) );
  NANDN U52674 ( .A(n38281), .B(n38280), .Z(n38282) );
  NAND U52675 ( .A(n38283), .B(n38282), .Z(n38284) );
  NANDN U52676 ( .A(n38285), .B(n38284), .Z(n38286) );
  AND U52677 ( .A(n51900), .B(n38286), .Z(n38288) );
  NAND U52678 ( .A(n38288), .B(n38287), .Z(n38289) );
  NANDN U52679 ( .A(n38290), .B(n38289), .Z(n38291) );
  AND U52680 ( .A(n38292), .B(n38291), .Z(n38293) );
  NANDN U52681 ( .A(x[3354]), .B(y[3354]), .Z(n51901) );
  NAND U52682 ( .A(n38293), .B(n51901), .Z(n38294) );
  NANDN U52683 ( .A(n38295), .B(n38294), .Z(n38296) );
  AND U52684 ( .A(n38297), .B(n38296), .Z(n38301) );
  NAND U52685 ( .A(n38299), .B(n38298), .Z(n38300) );
  OR U52686 ( .A(n38301), .B(n38300), .Z(n38302) );
  AND U52687 ( .A(n38303), .B(n38302), .Z(n38307) );
  NAND U52688 ( .A(n38305), .B(n38304), .Z(n38306) );
  OR U52689 ( .A(n38307), .B(n38306), .Z(n38308) );
  AND U52690 ( .A(n38309), .B(n38308), .Z(n38313) );
  NAND U52691 ( .A(n38311), .B(n38310), .Z(n38312) );
  OR U52692 ( .A(n38313), .B(n38312), .Z(n38314) );
  AND U52693 ( .A(n38315), .B(n38314), .Z(n38319) );
  NAND U52694 ( .A(n38317), .B(n38316), .Z(n38318) );
  OR U52695 ( .A(n38319), .B(n38318), .Z(n38320) );
  AND U52696 ( .A(n38321), .B(n38320), .Z(n38325) );
  NAND U52697 ( .A(n38323), .B(n38322), .Z(n38324) );
  OR U52698 ( .A(n38325), .B(n38324), .Z(n38326) );
  AND U52699 ( .A(n38327), .B(n38326), .Z(n38331) );
  NAND U52700 ( .A(n38329), .B(n38328), .Z(n38330) );
  OR U52701 ( .A(n38331), .B(n38330), .Z(n38332) );
  AND U52702 ( .A(n38333), .B(n38332), .Z(n38337) );
  NAND U52703 ( .A(n38335), .B(n38334), .Z(n38336) );
  OR U52704 ( .A(n38337), .B(n38336), .Z(n38338) );
  AND U52705 ( .A(n38339), .B(n38338), .Z(n38343) );
  NAND U52706 ( .A(n38341), .B(n38340), .Z(n38342) );
  OR U52707 ( .A(n38343), .B(n38342), .Z(n38344) );
  AND U52708 ( .A(n38345), .B(n38344), .Z(n38349) );
  NAND U52709 ( .A(n38347), .B(n38346), .Z(n38348) );
  OR U52710 ( .A(n38349), .B(n38348), .Z(n38350) );
  AND U52711 ( .A(n38351), .B(n38350), .Z(n38352) );
  NOR U52712 ( .A(n38353), .B(n38352), .Z(n38354) );
  NAND U52713 ( .A(n38355), .B(n38354), .Z(n38359) );
  NAND U52714 ( .A(n38357), .B(n38356), .Z(n38358) );
  ANDN U52715 ( .B(n38359), .A(n38358), .Z(n38363) );
  NAND U52716 ( .A(n38361), .B(n38360), .Z(n38362) );
  OR U52717 ( .A(n38363), .B(n38362), .Z(n38364) );
  AND U52718 ( .A(n38365), .B(n38364), .Z(n38369) );
  NAND U52719 ( .A(n38367), .B(n38366), .Z(n38368) );
  OR U52720 ( .A(n38369), .B(n38368), .Z(n38370) );
  AND U52721 ( .A(n38371), .B(n38370), .Z(n38372) );
  ANDN U52722 ( .B(n38373), .A(n38372), .Z(n38374) );
  NAND U52723 ( .A(n38375), .B(n38374), .Z(n38376) );
  NANDN U52724 ( .A(n38377), .B(n38376), .Z(n38378) );
  OR U52725 ( .A(n55605), .B(n38378), .Z(n38379) );
  AND U52726 ( .A(n38380), .B(n38379), .Z(n38382) );
  NAND U52727 ( .A(n38382), .B(n38381), .Z(n38383) );
  NANDN U52728 ( .A(n38384), .B(n38383), .Z(n38385) );
  AND U52729 ( .A(n38386), .B(n38385), .Z(n38388) );
  NAND U52730 ( .A(n38388), .B(n38387), .Z(n38389) );
  NANDN U52731 ( .A(n38390), .B(n38389), .Z(n38391) );
  AND U52732 ( .A(n38392), .B(n38391), .Z(n38393) );
  OR U52733 ( .A(n38394), .B(n38393), .Z(n38395) );
  NAND U52734 ( .A(n38396), .B(n38395), .Z(n38399) );
  NANDN U52735 ( .A(x[3390]), .B(y[3390]), .Z(n55611) );
  AND U52736 ( .A(n38397), .B(n55611), .Z(n38398) );
  NAND U52737 ( .A(n38399), .B(n38398), .Z(n38400) );
  NANDN U52738 ( .A(n38401), .B(n38400), .Z(n38402) );
  NAND U52739 ( .A(n38403), .B(n38402), .Z(n38404) );
  NANDN U52740 ( .A(n38405), .B(n38404), .Z(n38406) );
  AND U52741 ( .A(n55618), .B(n38406), .Z(n38408) );
  NAND U52742 ( .A(n38408), .B(n38407), .Z(n38409) );
  NANDN U52743 ( .A(n38410), .B(n38409), .Z(n38411) );
  AND U52744 ( .A(n38412), .B(n38411), .Z(n38416) );
  NAND U52745 ( .A(n38414), .B(n38413), .Z(n38415) );
  OR U52746 ( .A(n38416), .B(n38415), .Z(n38417) );
  AND U52747 ( .A(n38418), .B(n38417), .Z(n38422) );
  NAND U52748 ( .A(n38420), .B(n38419), .Z(n38421) );
  OR U52749 ( .A(n38422), .B(n38421), .Z(n38423) );
  AND U52750 ( .A(n38424), .B(n38423), .Z(n38428) );
  NAND U52751 ( .A(n38426), .B(n38425), .Z(n38427) );
  OR U52752 ( .A(n38428), .B(n38427), .Z(n38429) );
  AND U52753 ( .A(n38430), .B(n38429), .Z(n38434) );
  NAND U52754 ( .A(n38432), .B(n38431), .Z(n38433) );
  OR U52755 ( .A(n38434), .B(n38433), .Z(n38435) );
  AND U52756 ( .A(n38436), .B(n38435), .Z(n38440) );
  NAND U52757 ( .A(n38438), .B(n38437), .Z(n38439) );
  OR U52758 ( .A(n38440), .B(n38439), .Z(n38441) );
  AND U52759 ( .A(n38442), .B(n38441), .Z(n38446) );
  NAND U52760 ( .A(n38444), .B(n38443), .Z(n38445) );
  OR U52761 ( .A(n38446), .B(n38445), .Z(n38447) );
  AND U52762 ( .A(n38448), .B(n38447), .Z(n38452) );
  NAND U52763 ( .A(n38450), .B(n38449), .Z(n38451) );
  OR U52764 ( .A(n38452), .B(n38451), .Z(n38453) );
  AND U52765 ( .A(n38454), .B(n38453), .Z(n38458) );
  NAND U52766 ( .A(n38456), .B(n38455), .Z(n38457) );
  OR U52767 ( .A(n38458), .B(n38457), .Z(n38459) );
  AND U52768 ( .A(n38460), .B(n38459), .Z(n38464) );
  NAND U52769 ( .A(n38462), .B(n38461), .Z(n38463) );
  OR U52770 ( .A(n38464), .B(n38463), .Z(n38465) );
  AND U52771 ( .A(n38466), .B(n38465), .Z(n38467) );
  OR U52772 ( .A(n38468), .B(n38467), .Z(n38469) );
  NAND U52773 ( .A(n38470), .B(n38469), .Z(n38471) );
  AND U52774 ( .A(n38472), .B(n38471), .Z(n38473) );
  NOR U52775 ( .A(n55642), .B(n38473), .Z(n38474) );
  NANDN U52776 ( .A(n38475), .B(n38474), .Z(n38476) );
  AND U52777 ( .A(n38477), .B(n38476), .Z(n38479) );
  NAND U52778 ( .A(n38479), .B(n38478), .Z(n38480) );
  NANDN U52779 ( .A(n38481), .B(n38480), .Z(n38482) );
  AND U52780 ( .A(n38483), .B(n38482), .Z(n38485) );
  NAND U52781 ( .A(n38485), .B(n38484), .Z(n38486) );
  NANDN U52782 ( .A(n38487), .B(n38486), .Z(n38488) );
  AND U52783 ( .A(n38489), .B(n38488), .Z(n38491) );
  NAND U52784 ( .A(n38491), .B(n38490), .Z(n38494) );
  NANDN U52785 ( .A(x[3424]), .B(y[3424]), .Z(n55650) );
  AND U52786 ( .A(n38492), .B(n55650), .Z(n38493) );
  NAND U52787 ( .A(n38494), .B(n38493), .Z(n38498) );
  NAND U52788 ( .A(n38496), .B(n38495), .Z(n38497) );
  ANDN U52789 ( .B(n38498), .A(n38497), .Z(n38502) );
  NAND U52790 ( .A(n38500), .B(n38499), .Z(n38501) );
  OR U52791 ( .A(n38502), .B(n38501), .Z(n38503) );
  AND U52792 ( .A(n38504), .B(n38503), .Z(n38505) );
  OR U52793 ( .A(n38506), .B(n38505), .Z(n38507) );
  NAND U52794 ( .A(n38508), .B(n38507), .Z(n38509) );
  AND U52795 ( .A(n38510), .B(n38509), .Z(n38511) );
  NOR U52796 ( .A(n38512), .B(n38511), .Z(n38514) );
  NAND U52797 ( .A(n38514), .B(n38513), .Z(n38516) );
  AND U52798 ( .A(n38516), .B(n38515), .Z(n38517) );
  NANDN U52799 ( .A(x[3432]), .B(y[3432]), .Z(n55659) );
  AND U52800 ( .A(n38517), .B(n55659), .Z(n38518) );
  ANDN U52801 ( .B(n38519), .A(n38518), .Z(n38523) );
  NAND U52802 ( .A(n38521), .B(n38520), .Z(n38522) );
  OR U52803 ( .A(n38523), .B(n38522), .Z(n38524) );
  AND U52804 ( .A(n38525), .B(n38524), .Z(n38529) );
  NANDN U52805 ( .A(x[3436]), .B(y[3436]), .Z(n38527) );
  NAND U52806 ( .A(n38527), .B(n38526), .Z(n38528) );
  OR U52807 ( .A(n38529), .B(n38528), .Z(n38530) );
  AND U52808 ( .A(n38531), .B(n38530), .Z(n38533) );
  NAND U52809 ( .A(n38533), .B(n38532), .Z(n38534) );
  NANDN U52810 ( .A(n38535), .B(n38534), .Z(n38536) );
  AND U52811 ( .A(n38537), .B(n38536), .Z(n38541) );
  NAND U52812 ( .A(n38539), .B(n38538), .Z(n38540) );
  OR U52813 ( .A(n38541), .B(n38540), .Z(n38542) );
  AND U52814 ( .A(n38543), .B(n38542), .Z(n38544) );
  NOR U52815 ( .A(n38545), .B(n38544), .Z(n38546) );
  NAND U52816 ( .A(n38547), .B(n38546), .Z(n38548) );
  NANDN U52817 ( .A(n38549), .B(n38548), .Z(n38550) );
  NAND U52818 ( .A(n38551), .B(n38550), .Z(n38552) );
  NANDN U52819 ( .A(n38553), .B(n38552), .Z(n38554) );
  AND U52820 ( .A(n38555), .B(n38554), .Z(n38557) );
  NAND U52821 ( .A(n38557), .B(n38556), .Z(n38558) );
  NANDN U52822 ( .A(n38559), .B(n38558), .Z(n38560) );
  AND U52823 ( .A(n38561), .B(n38560), .Z(n38563) );
  NAND U52824 ( .A(n38563), .B(n38562), .Z(n38564) );
  NANDN U52825 ( .A(n38565), .B(n38564), .Z(n38566) );
  AND U52826 ( .A(n38567), .B(n38566), .Z(n38569) );
  NANDN U52827 ( .A(x[3450]), .B(y[3450]), .Z(n38568) );
  NAND U52828 ( .A(n38569), .B(n38568), .Z(n38570) );
  NANDN U52829 ( .A(n38571), .B(n38570), .Z(n38572) );
  AND U52830 ( .A(n38573), .B(n38572), .Z(n38574) );
  OR U52831 ( .A(n38575), .B(n38574), .Z(n38576) );
  NAND U52832 ( .A(n38577), .B(n38576), .Z(n38578) );
  AND U52833 ( .A(n38579), .B(n38578), .Z(n38580) );
  OR U52834 ( .A(n38581), .B(n38580), .Z(n38582) );
  NAND U52835 ( .A(n38583), .B(n38582), .Z(n38584) );
  NANDN U52836 ( .A(n38585), .B(n38584), .Z(n38586) );
  AND U52837 ( .A(n38587), .B(n38586), .Z(n38588) );
  ANDN U52838 ( .B(n38589), .A(n38588), .Z(n38593) );
  AND U52839 ( .A(n38591), .B(n38590), .Z(n38592) );
  NANDN U52840 ( .A(n38593), .B(n38592), .Z(n38594) );
  NANDN U52841 ( .A(n38595), .B(n38594), .Z(n38596) );
  AND U52842 ( .A(n38597), .B(n38596), .Z(n38599) );
  NAND U52843 ( .A(n38599), .B(n38598), .Z(n38600) );
  NANDN U52844 ( .A(n38601), .B(n38600), .Z(n38602) );
  AND U52845 ( .A(n38603), .B(n38602), .Z(n38605) );
  NAND U52846 ( .A(n38605), .B(n38604), .Z(n38606) );
  NANDN U52847 ( .A(n38607), .B(n38606), .Z(n38608) );
  AND U52848 ( .A(n38609), .B(n38608), .Z(n38611) );
  NAND U52849 ( .A(n38611), .B(n38610), .Z(n38612) );
  NANDN U52850 ( .A(n38613), .B(n38612), .Z(n38614) );
  AND U52851 ( .A(n38615), .B(n38614), .Z(n38617) );
  NAND U52852 ( .A(n38617), .B(n38616), .Z(n38618) );
  NANDN U52853 ( .A(n38619), .B(n38618), .Z(n38620) );
  AND U52854 ( .A(n38621), .B(n38620), .Z(n38623) );
  AND U52855 ( .A(n38623), .B(n38622), .Z(n38627) );
  NAND U52856 ( .A(n38625), .B(n38624), .Z(n38626) );
  OR U52857 ( .A(n38627), .B(n38626), .Z(n38628) );
  AND U52858 ( .A(n38629), .B(n38628), .Z(n38630) );
  OR U52859 ( .A(n38631), .B(n38630), .Z(n38632) );
  NAND U52860 ( .A(n38633), .B(n38632), .Z(n38634) );
  AND U52861 ( .A(n38635), .B(n38634), .Z(n38639) );
  AND U52862 ( .A(n38637), .B(n38636), .Z(n38638) );
  NANDN U52863 ( .A(n38639), .B(n38638), .Z(n38642) );
  NANDN U52864 ( .A(x[3478]), .B(y[3478]), .Z(n51882) );
  AND U52865 ( .A(n38640), .B(n51882), .Z(n38641) );
  NAND U52866 ( .A(n38642), .B(n38641), .Z(n38643) );
  NANDN U52867 ( .A(n38644), .B(n38643), .Z(n38645) );
  NAND U52868 ( .A(n38646), .B(n38645), .Z(n38647) );
  NANDN U52869 ( .A(n38648), .B(n38647), .Z(n38649) );
  AND U52870 ( .A(n38650), .B(n38649), .Z(n38652) );
  NAND U52871 ( .A(n38652), .B(n38651), .Z(n38653) );
  NANDN U52872 ( .A(n38654), .B(n38653), .Z(n38655) );
  AND U52873 ( .A(n38656), .B(n38655), .Z(n38658) );
  NANDN U52874 ( .A(x[3484]), .B(y[3484]), .Z(n38657) );
  AND U52875 ( .A(n38658), .B(n38657), .Z(n38662) );
  NAND U52876 ( .A(n38660), .B(n38659), .Z(n38661) );
  OR U52877 ( .A(n38662), .B(n38661), .Z(n38663) );
  AND U52878 ( .A(n38664), .B(n38663), .Z(n38666) );
  NANDN U52879 ( .A(x[3486]), .B(y[3486]), .Z(n38665) );
  NAND U52880 ( .A(n38666), .B(n38665), .Z(n38667) );
  NANDN U52881 ( .A(n38668), .B(n38667), .Z(n38669) );
  AND U52882 ( .A(n38670), .B(n38669), .Z(n38674) );
  NAND U52883 ( .A(n38672), .B(n38671), .Z(n38673) );
  OR U52884 ( .A(n38674), .B(n38673), .Z(n38675) );
  AND U52885 ( .A(n38676), .B(n38675), .Z(n38680) );
  NAND U52886 ( .A(n38678), .B(n38677), .Z(n38679) );
  OR U52887 ( .A(n38680), .B(n38679), .Z(n38681) );
  AND U52888 ( .A(n38682), .B(n38681), .Z(n38683) );
  OR U52889 ( .A(n38684), .B(n38683), .Z(n38685) );
  NAND U52890 ( .A(n38686), .B(n38685), .Z(n38687) );
  AND U52891 ( .A(n38688), .B(n38687), .Z(n38689) );
  ANDN U52892 ( .B(n51877), .A(n38689), .Z(n38690) );
  OR U52893 ( .A(n38691), .B(n38690), .Z(n38692) );
  NAND U52894 ( .A(n38693), .B(n38692), .Z(n38694) );
  NAND U52895 ( .A(n38695), .B(n38694), .Z(n38696) );
  NANDN U52896 ( .A(n38697), .B(n38696), .Z(n38698) );
  AND U52897 ( .A(n38699), .B(n38698), .Z(n38701) );
  NAND U52898 ( .A(n38701), .B(n38700), .Z(n38702) );
  NANDN U52899 ( .A(n38703), .B(n38702), .Z(n38704) );
  AND U52900 ( .A(n38705), .B(n38704), .Z(n38707) );
  NAND U52901 ( .A(n38707), .B(n38706), .Z(n38708) );
  NANDN U52902 ( .A(n38709), .B(n38708), .Z(n38710) );
  AND U52903 ( .A(n38711), .B(n38710), .Z(n38713) );
  NAND U52904 ( .A(n38713), .B(n38712), .Z(n38716) );
  NANDN U52905 ( .A(x[3506]), .B(y[3506]), .Z(n55775) );
  AND U52906 ( .A(n38714), .B(n55775), .Z(n38715) );
  NAND U52907 ( .A(n38716), .B(n38715), .Z(n38717) );
  NANDN U52908 ( .A(n38718), .B(n38717), .Z(n38719) );
  NAND U52909 ( .A(n38720), .B(n38719), .Z(n38721) );
  NANDN U52910 ( .A(n38722), .B(n38721), .Z(n38723) );
  AND U52911 ( .A(n38724), .B(n38723), .Z(n38726) );
  NAND U52912 ( .A(n38726), .B(n38725), .Z(n38727) );
  NANDN U52913 ( .A(n38728), .B(n38727), .Z(n38729) );
  AND U52914 ( .A(n38730), .B(n38729), .Z(n38732) );
  NAND U52915 ( .A(n38732), .B(n38731), .Z(n38733) );
  NANDN U52916 ( .A(n38734), .B(n38733), .Z(n38735) );
  AND U52917 ( .A(n38736), .B(n38735), .Z(n38738) );
  NAND U52918 ( .A(n38738), .B(n38737), .Z(n38739) );
  NANDN U52919 ( .A(n38740), .B(n38739), .Z(n38741) );
  AND U52920 ( .A(n38742), .B(n38741), .Z(n38744) );
  NANDN U52921 ( .A(x[3516]), .B(y[3516]), .Z(n38743) );
  AND U52922 ( .A(n38744), .B(n38743), .Z(n38748) );
  NAND U52923 ( .A(n38746), .B(n38745), .Z(n38747) );
  OR U52924 ( .A(n38748), .B(n38747), .Z(n38749) );
  AND U52925 ( .A(n38750), .B(n38749), .Z(n38754) );
  NAND U52926 ( .A(n38752), .B(n38751), .Z(n38753) );
  OR U52927 ( .A(n38754), .B(n38753), .Z(n38755) );
  AND U52928 ( .A(n38756), .B(n38755), .Z(n38758) );
  AND U52929 ( .A(n38758), .B(n38757), .Z(n38762) );
  NAND U52930 ( .A(n38760), .B(n38759), .Z(n38761) );
  OR U52931 ( .A(n38762), .B(n38761), .Z(n38763) );
  AND U52932 ( .A(n38764), .B(n38763), .Z(n38765) );
  OR U52933 ( .A(n38766), .B(n38765), .Z(n38767) );
  NAND U52934 ( .A(n38768), .B(n38767), .Z(n38769) );
  AND U52935 ( .A(n38770), .B(n38769), .Z(n38771) );
  NOR U52936 ( .A(n55794), .B(n38771), .Z(n38772) );
  NANDN U52937 ( .A(n38773), .B(n38772), .Z(n38774) );
  AND U52938 ( .A(n38775), .B(n38774), .Z(n38777) );
  NAND U52939 ( .A(n38777), .B(n38776), .Z(n38778) );
  NANDN U52940 ( .A(n38779), .B(n38778), .Z(n38780) );
  AND U52941 ( .A(n38781), .B(n38780), .Z(n38783) );
  NAND U52942 ( .A(n38783), .B(n38782), .Z(n38784) );
  NANDN U52943 ( .A(n38785), .B(n38784), .Z(n38786) );
  AND U52944 ( .A(n38787), .B(n38786), .Z(n38789) );
  NAND U52945 ( .A(n38789), .B(n38788), .Z(n38792) );
  NANDN U52946 ( .A(x[3532]), .B(y[3532]), .Z(n51870) );
  AND U52947 ( .A(n38790), .B(n51870), .Z(n38791) );
  NAND U52948 ( .A(n38792), .B(n38791), .Z(n38793) );
  NANDN U52949 ( .A(n38794), .B(n38793), .Z(n38795) );
  NAND U52950 ( .A(n38796), .B(n38795), .Z(n38797) );
  NAND U52951 ( .A(n38798), .B(n38797), .Z(n38799) );
  NANDN U52952 ( .A(n38800), .B(n38799), .Z(n38801) );
  NANDN U52953 ( .A(x[3536]), .B(y[3536]), .Z(n55801) );
  NANDN U52954 ( .A(n38801), .B(n55801), .Z(n38802) );
  NAND U52955 ( .A(n38803), .B(n38802), .Z(n38804) );
  NANDN U52956 ( .A(n38805), .B(n38804), .Z(n38807) );
  OR U52957 ( .A(n38807), .B(n38806), .Z(n38808) );
  NANDN U52958 ( .A(n38809), .B(n38808), .Z(n38810) );
  AND U52959 ( .A(n38811), .B(n38810), .Z(n38815) );
  NAND U52960 ( .A(n38813), .B(n38812), .Z(n38814) );
  OR U52961 ( .A(n38815), .B(n38814), .Z(n38816) );
  AND U52962 ( .A(n38817), .B(n38816), .Z(n38821) );
  NAND U52963 ( .A(n38819), .B(n38818), .Z(n38820) );
  OR U52964 ( .A(n38821), .B(n38820), .Z(n38822) );
  AND U52965 ( .A(n38823), .B(n38822), .Z(n38824) );
  NOR U52966 ( .A(n38825), .B(n38824), .Z(n38826) );
  NAND U52967 ( .A(n38827), .B(n38826), .Z(n38828) );
  NANDN U52968 ( .A(n38829), .B(n38828), .Z(n38830) );
  AND U52969 ( .A(n38831), .B(n38830), .Z(n38834) );
  AND U52970 ( .A(n38832), .B(n55814), .Z(n38833) );
  NANDN U52971 ( .A(n38834), .B(n38833), .Z(n38835) );
  NAND U52972 ( .A(n38836), .B(n38835), .Z(n38838) );
  OR U52973 ( .A(n38838), .B(n38837), .Z(n38839) );
  NAND U52974 ( .A(n38840), .B(n38839), .Z(n38841) );
  NANDN U52975 ( .A(n38842), .B(n38841), .Z(n38844) );
  OR U52976 ( .A(n38844), .B(n38843), .Z(n38845) );
  NAND U52977 ( .A(n38846), .B(n38845), .Z(n38847) );
  NANDN U52978 ( .A(n38848), .B(n38847), .Z(n38849) );
  AND U52979 ( .A(n38850), .B(n38849), .Z(n38851) );
  NAND U52980 ( .A(n38852), .B(n38851), .Z(n38856) );
  NAND U52981 ( .A(n38854), .B(n38853), .Z(n38855) );
  ANDN U52982 ( .B(n38856), .A(n38855), .Z(n38860) );
  NAND U52983 ( .A(n38858), .B(n38857), .Z(n38859) );
  OR U52984 ( .A(n38860), .B(n38859), .Z(n38861) );
  AND U52985 ( .A(n38862), .B(n38861), .Z(n38866) );
  NAND U52986 ( .A(n38864), .B(n38863), .Z(n38865) );
  OR U52987 ( .A(n38866), .B(n38865), .Z(n38867) );
  AND U52988 ( .A(n38868), .B(n38867), .Z(n38872) );
  NAND U52989 ( .A(n38870), .B(n38869), .Z(n38871) );
  OR U52990 ( .A(n38872), .B(n38871), .Z(n38873) );
  AND U52991 ( .A(n38874), .B(n38873), .Z(n38878) );
  NAND U52992 ( .A(n38876), .B(n38875), .Z(n38877) );
  OR U52993 ( .A(n38878), .B(n38877), .Z(n38879) );
  AND U52994 ( .A(n38880), .B(n38879), .Z(n38881) );
  OR U52995 ( .A(n38882), .B(n38881), .Z(n38883) );
  NAND U52996 ( .A(n38884), .B(n38883), .Z(n38885) );
  AND U52997 ( .A(n38886), .B(n38885), .Z(n38887) );
  NOR U52998 ( .A(n38888), .B(n38887), .Z(n38890) );
  NAND U52999 ( .A(n38890), .B(n38889), .Z(n38893) );
  NANDN U53000 ( .A(x[3568]), .B(y[3568]), .Z(n55832) );
  AND U53001 ( .A(n38891), .B(n55832), .Z(n38892) );
  NAND U53002 ( .A(n38893), .B(n38892), .Z(n38894) );
  NANDN U53003 ( .A(n38895), .B(n38894), .Z(n38896) );
  NAND U53004 ( .A(n38897), .B(n38896), .Z(n38898) );
  NANDN U53005 ( .A(n38899), .B(n38898), .Z(n38900) );
  AND U53006 ( .A(n38901), .B(n38900), .Z(n38902) );
  NANDN U53007 ( .A(x[3572]), .B(y[3572]), .Z(n55837) );
  NAND U53008 ( .A(n38902), .B(n55837), .Z(n38903) );
  AND U53009 ( .A(n38904), .B(n38903), .Z(n38908) );
  NAND U53010 ( .A(n38906), .B(n38905), .Z(n38907) );
  OR U53011 ( .A(n38908), .B(n38907), .Z(n38909) );
  AND U53012 ( .A(n38910), .B(n38909), .Z(n38914) );
  NAND U53013 ( .A(n38912), .B(n38911), .Z(n38913) );
  OR U53014 ( .A(n38914), .B(n38913), .Z(n38915) );
  AND U53015 ( .A(n38916), .B(n38915), .Z(n38917) );
  ANDN U53016 ( .B(n38918), .A(n38917), .Z(n38919) );
  NAND U53017 ( .A(n38920), .B(n38919), .Z(n38921) );
  NANDN U53018 ( .A(n38922), .B(n38921), .Z(n38923) );
  OR U53019 ( .A(n38924), .B(n38923), .Z(n38925) );
  AND U53020 ( .A(n38926), .B(n38925), .Z(n38928) );
  NAND U53021 ( .A(n38928), .B(n38927), .Z(n38929) );
  NANDN U53022 ( .A(n38930), .B(n38929), .Z(n38931) );
  AND U53023 ( .A(n38932), .B(n38931), .Z(n38936) );
  NAND U53024 ( .A(n38934), .B(n38933), .Z(n38935) );
  OR U53025 ( .A(n38936), .B(n38935), .Z(n38937) );
  AND U53026 ( .A(n38938), .B(n38937), .Z(n38942) );
  NAND U53027 ( .A(n38940), .B(n38939), .Z(n38941) );
  OR U53028 ( .A(n38942), .B(n38941), .Z(n38943) );
  AND U53029 ( .A(n38944), .B(n38943), .Z(n38945) );
  ANDN U53030 ( .B(n38946), .A(n38945), .Z(n38947) );
  NAND U53031 ( .A(n38948), .B(n38947), .Z(n38949) );
  NANDN U53032 ( .A(n38950), .B(n38949), .Z(n38952) );
  ANDN U53033 ( .B(y[3588]), .A(x[3588]), .Z(n38951) );
  OR U53034 ( .A(n38952), .B(n38951), .Z(n38953) );
  NAND U53035 ( .A(n38954), .B(n38953), .Z(n38958) );
  NAND U53036 ( .A(n38956), .B(n38955), .Z(n38957) );
  ANDN U53037 ( .B(n38958), .A(n38957), .Z(n38962) );
  NAND U53038 ( .A(n38960), .B(n38959), .Z(n38961) );
  OR U53039 ( .A(n38962), .B(n38961), .Z(n38963) );
  AND U53040 ( .A(n38964), .B(n38963), .Z(n38968) );
  AND U53041 ( .A(n38966), .B(n38965), .Z(n38967) );
  NANDN U53042 ( .A(n38968), .B(n38967), .Z(n38969) );
  NAND U53043 ( .A(n38970), .B(n38969), .Z(n38971) );
  AND U53044 ( .A(n38972), .B(n38971), .Z(n38976) );
  NAND U53045 ( .A(n38974), .B(n38973), .Z(n38975) );
  OR U53046 ( .A(n38976), .B(n38975), .Z(n38977) );
  AND U53047 ( .A(n38978), .B(n38977), .Z(n38980) );
  NAND U53048 ( .A(n38980), .B(n38979), .Z(n38981) );
  NANDN U53049 ( .A(n38982), .B(n38981), .Z(n38983) );
  AND U53050 ( .A(n38984), .B(n38983), .Z(n38986) );
  NAND U53051 ( .A(n38986), .B(n38985), .Z(n38987) );
  NANDN U53052 ( .A(n38988), .B(n38987), .Z(n38989) );
  AND U53053 ( .A(n38990), .B(n38989), .Z(n38992) );
  NAND U53054 ( .A(n38992), .B(n38991), .Z(n38993) );
  NANDN U53055 ( .A(n38994), .B(n38993), .Z(n38995) );
  AND U53056 ( .A(n38996), .B(n38995), .Z(n38998) );
  AND U53057 ( .A(n38998), .B(n38997), .Z(n39002) );
  NAND U53058 ( .A(n39000), .B(n38999), .Z(n39001) );
  OR U53059 ( .A(n39002), .B(n39001), .Z(n39003) );
  AND U53060 ( .A(n39004), .B(n39003), .Z(n39008) );
  NAND U53061 ( .A(n39006), .B(n39005), .Z(n39007) );
  OR U53062 ( .A(n39008), .B(n39007), .Z(n39009) );
  AND U53063 ( .A(n39010), .B(n39009), .Z(n39014) );
  NAND U53064 ( .A(n39012), .B(n39011), .Z(n39013) );
  OR U53065 ( .A(n39014), .B(n39013), .Z(n39015) );
  AND U53066 ( .A(n39016), .B(n39015), .Z(n39020) );
  NAND U53067 ( .A(n39018), .B(n39017), .Z(n39019) );
  OR U53068 ( .A(n39020), .B(n39019), .Z(n39021) );
  AND U53069 ( .A(n39022), .B(n39021), .Z(n39025) );
  AND U53070 ( .A(n39023), .B(n51852), .Z(n39024) );
  NANDN U53071 ( .A(n39025), .B(n39024), .Z(n39026) );
  NANDN U53072 ( .A(n39027), .B(n39026), .Z(n39028) );
  AND U53073 ( .A(n39029), .B(n39028), .Z(n39030) );
  NANDN U53074 ( .A(x[3614]), .B(y[3614]), .Z(n51853) );
  AND U53075 ( .A(n39030), .B(n51853), .Z(n39031) );
  OR U53076 ( .A(n39032), .B(n39031), .Z(n39033) );
  NAND U53077 ( .A(n39034), .B(n39033), .Z(n39038) );
  NAND U53078 ( .A(n39036), .B(n39035), .Z(n39037) );
  ANDN U53079 ( .B(n39038), .A(n39037), .Z(n39042) );
  NAND U53080 ( .A(n39040), .B(n39039), .Z(n39041) );
  OR U53081 ( .A(n39042), .B(n39041), .Z(n39043) );
  AND U53082 ( .A(n39044), .B(n39043), .Z(n39048) );
  NAND U53083 ( .A(n39046), .B(n39045), .Z(n39047) );
  OR U53084 ( .A(n39048), .B(n39047), .Z(n39049) );
  AND U53085 ( .A(n39050), .B(n39049), .Z(n39054) );
  AND U53086 ( .A(n39052), .B(n39051), .Z(n39053) );
  NANDN U53087 ( .A(n39054), .B(n39053), .Z(n39055) );
  NANDN U53088 ( .A(n39056), .B(n39055), .Z(n39057) );
  AND U53089 ( .A(n39058), .B(n39057), .Z(n39060) );
  NAND U53090 ( .A(n39060), .B(n39059), .Z(n39061) );
  NANDN U53091 ( .A(n39062), .B(n39061), .Z(n39063) );
  AND U53092 ( .A(n39064), .B(n39063), .Z(n39066) );
  NAND U53093 ( .A(n39066), .B(n39065), .Z(n39067) );
  NANDN U53094 ( .A(n39068), .B(n39067), .Z(n39070) );
  IV U53095 ( .A(n39069), .Z(n51844) );
  AND U53096 ( .A(n39070), .B(n51844), .Z(n39072) );
  AND U53097 ( .A(n39072), .B(n39071), .Z(n39076) );
  NAND U53098 ( .A(n39074), .B(n39073), .Z(n39075) );
  OR U53099 ( .A(n39076), .B(n39075), .Z(n39077) );
  AND U53100 ( .A(n39078), .B(n39077), .Z(n39082) );
  NAND U53101 ( .A(n39080), .B(n39079), .Z(n39081) );
  OR U53102 ( .A(n39082), .B(n39081), .Z(n39083) );
  AND U53103 ( .A(n39084), .B(n39083), .Z(n39088) );
  NAND U53104 ( .A(n39086), .B(n39085), .Z(n39087) );
  OR U53105 ( .A(n39088), .B(n39087), .Z(n39089) );
  AND U53106 ( .A(n39090), .B(n39089), .Z(n39094) );
  NAND U53107 ( .A(n39092), .B(n39091), .Z(n39093) );
  OR U53108 ( .A(n39094), .B(n39093), .Z(n39095) );
  AND U53109 ( .A(n39096), .B(n39095), .Z(n39100) );
  NAND U53110 ( .A(n39098), .B(n39097), .Z(n39099) );
  OR U53111 ( .A(n39100), .B(n39099), .Z(n39101) );
  AND U53112 ( .A(n39102), .B(n39101), .Z(n39103) );
  ANDN U53113 ( .B(n39104), .A(n39103), .Z(n39105) );
  NAND U53114 ( .A(n39106), .B(n39105), .Z(n39107) );
  NANDN U53115 ( .A(n39108), .B(n39107), .Z(n39109) );
  OR U53116 ( .A(n39110), .B(n39109), .Z(n39111) );
  AND U53117 ( .A(n39112), .B(n39111), .Z(n39114) );
  NAND U53118 ( .A(n39114), .B(n39113), .Z(n39115) );
  NANDN U53119 ( .A(n39116), .B(n39115), .Z(n39117) );
  AND U53120 ( .A(n39118), .B(n39117), .Z(n39120) );
  NAND U53121 ( .A(n39120), .B(n39119), .Z(n39121) );
  NANDN U53122 ( .A(n39122), .B(n39121), .Z(n39123) );
  AND U53123 ( .A(n39124), .B(n39123), .Z(n39126) );
  NAND U53124 ( .A(n39126), .B(n39125), .Z(n39128) );
  NANDN U53125 ( .A(x[3646]), .B(y[3646]), .Z(n51836) );
  AND U53126 ( .A(n55904), .B(n51836), .Z(n39127) );
  NAND U53127 ( .A(n39128), .B(n39127), .Z(n39129) );
  NANDN U53128 ( .A(n39130), .B(n39129), .Z(n39131) );
  NAND U53129 ( .A(n39132), .B(n39131), .Z(n39133) );
  NAND U53130 ( .A(n39134), .B(n39133), .Z(n39135) );
  NANDN U53131 ( .A(n39136), .B(n39135), .Z(n39138) );
  ANDN U53132 ( .B(y[3650]), .A(x[3650]), .Z(n39137) );
  OR U53133 ( .A(n39138), .B(n39137), .Z(n39139) );
  NAND U53134 ( .A(n39140), .B(n39139), .Z(n39141) );
  NANDN U53135 ( .A(n39142), .B(n39141), .Z(n39144) );
  OR U53136 ( .A(n39144), .B(n39143), .Z(n39145) );
  NANDN U53137 ( .A(n39146), .B(n39145), .Z(n39147) );
  AND U53138 ( .A(n39148), .B(n39147), .Z(n39149) );
  OR U53139 ( .A(n39150), .B(n39149), .Z(n39151) );
  NAND U53140 ( .A(n39152), .B(n39151), .Z(n39153) );
  AND U53141 ( .A(n39154), .B(n39153), .Z(n39155) );
  ANDN U53142 ( .B(n39156), .A(n39155), .Z(n39157) );
  OR U53143 ( .A(n39158), .B(n39157), .Z(n39159) );
  NAND U53144 ( .A(n39160), .B(n39159), .Z(n39161) );
  NAND U53145 ( .A(n39162), .B(n39161), .Z(n39163) );
  ANDN U53146 ( .B(y[3662]), .A(x[3662]), .Z(n55919) );
  ANDN U53147 ( .B(n39163), .A(n55919), .Z(n39164) );
  NANDN U53148 ( .A(n39165), .B(n39164), .Z(n39166) );
  NAND U53149 ( .A(n39167), .B(n39166), .Z(n39168) );
  NANDN U53150 ( .A(n39169), .B(n39168), .Z(n39170) );
  AND U53151 ( .A(n39171), .B(n39170), .Z(n39173) );
  NAND U53152 ( .A(n39173), .B(n39172), .Z(n39174) );
  NANDN U53153 ( .A(n39175), .B(n39174), .Z(n39176) );
  AND U53154 ( .A(n39177), .B(n39176), .Z(n39179) );
  NAND U53155 ( .A(n39179), .B(n39178), .Z(n39180) );
  NANDN U53156 ( .A(n39181), .B(n39180), .Z(n39182) );
  AND U53157 ( .A(n39183), .B(n39182), .Z(n39185) );
  NAND U53158 ( .A(n39185), .B(n39184), .Z(n39189) );
  NANDN U53159 ( .A(x[3670]), .B(y[3670]), .Z(n39186) );
  AND U53160 ( .A(n39187), .B(n39186), .Z(n39188) );
  NAND U53161 ( .A(n39189), .B(n39188), .Z(n39190) );
  NANDN U53162 ( .A(n39191), .B(n39190), .Z(n39192) );
  AND U53163 ( .A(n39193), .B(n39192), .Z(n39194) );
  ANDN U53164 ( .B(n39195), .A(n39194), .Z(n39196) );
  OR U53165 ( .A(n39197), .B(n39196), .Z(n39198) );
  NAND U53166 ( .A(n39199), .B(n39198), .Z(n39200) );
  AND U53167 ( .A(n39201), .B(n39200), .Z(n39202) );
  NAND U53168 ( .A(n39203), .B(n39202), .Z(n39204) );
  NANDN U53169 ( .A(n39205), .B(n39204), .Z(n39206) );
  AND U53170 ( .A(n39207), .B(n39206), .Z(n39208) );
  OR U53171 ( .A(n39209), .B(n39208), .Z(n39210) );
  NAND U53172 ( .A(n39211), .B(n39210), .Z(n39215) );
  NAND U53173 ( .A(n39213), .B(n39212), .Z(n39214) );
  ANDN U53174 ( .B(n39215), .A(n39214), .Z(n39219) );
  NAND U53175 ( .A(n39217), .B(n39216), .Z(n39218) );
  OR U53176 ( .A(n39219), .B(n39218), .Z(n39220) );
  AND U53177 ( .A(n39221), .B(n39220), .Z(n39225) );
  NAND U53178 ( .A(n39223), .B(n39222), .Z(n39224) );
  OR U53179 ( .A(n39225), .B(n39224), .Z(n39226) );
  AND U53180 ( .A(n39227), .B(n39226), .Z(n39231) );
  NAND U53181 ( .A(n39229), .B(n39228), .Z(n39230) );
  OR U53182 ( .A(n39231), .B(n39230), .Z(n39232) );
  AND U53183 ( .A(n39233), .B(n39232), .Z(n39237) );
  NAND U53184 ( .A(n39235), .B(n39234), .Z(n39236) );
  OR U53185 ( .A(n39237), .B(n39236), .Z(n39238) );
  AND U53186 ( .A(n39239), .B(n39238), .Z(n39240) );
  OR U53187 ( .A(n39241), .B(n39240), .Z(n39242) );
  NAND U53188 ( .A(n39243), .B(n39242), .Z(n39244) );
  AND U53189 ( .A(n39245), .B(n39244), .Z(n39246) );
  NOR U53190 ( .A(n39247), .B(n39246), .Z(n39249) );
  NAND U53191 ( .A(n39249), .B(n39248), .Z(n39252) );
  NANDN U53192 ( .A(x[3694]), .B(y[3694]), .Z(n55947) );
  AND U53193 ( .A(n39250), .B(n55947), .Z(n39251) );
  NAND U53194 ( .A(n39252), .B(n39251), .Z(n39253) );
  NANDN U53195 ( .A(n39254), .B(n39253), .Z(n39255) );
  NAND U53196 ( .A(n39256), .B(n39255), .Z(n39257) );
  NANDN U53197 ( .A(n39258), .B(n39257), .Z(n39259) );
  AND U53198 ( .A(n39260), .B(n39259), .Z(n39262) );
  NAND U53199 ( .A(n39262), .B(n39261), .Z(n39263) );
  NANDN U53200 ( .A(n39264), .B(n39263), .Z(n39265) );
  AND U53201 ( .A(n39266), .B(n39265), .Z(n39267) );
  NANDN U53202 ( .A(n39268), .B(n39267), .Z(n39269) );
  NAND U53203 ( .A(n39270), .B(n39269), .Z(n39271) );
  NANDN U53204 ( .A(n39272), .B(n39271), .Z(n39273) );
  NAND U53205 ( .A(n39274), .B(n39273), .Z(n39275) );
  NAND U53206 ( .A(n39276), .B(n39275), .Z(n39277) );
  NANDN U53207 ( .A(n39278), .B(n39277), .Z(n39281) );
  NANDN U53208 ( .A(x[3706]), .B(y[3706]), .Z(n55956) );
  ANDN U53209 ( .B(n55956), .A(n39279), .Z(n39280) );
  NAND U53210 ( .A(n39281), .B(n39280), .Z(n39282) );
  AND U53211 ( .A(n39283), .B(n39282), .Z(n39285) );
  NAND U53212 ( .A(n39285), .B(n39284), .Z(n39286) );
  NANDN U53213 ( .A(n39287), .B(n39286), .Z(n39288) );
  AND U53214 ( .A(n39289), .B(n39288), .Z(n39291) );
  NAND U53215 ( .A(n39291), .B(n39290), .Z(n39292) );
  NANDN U53216 ( .A(n39293), .B(n39292), .Z(n39294) );
  AND U53217 ( .A(n39295), .B(n39294), .Z(n39297) );
  AND U53218 ( .A(n39297), .B(n39296), .Z(n39301) );
  NAND U53219 ( .A(n39299), .B(n39298), .Z(n39300) );
  OR U53220 ( .A(n39301), .B(n39300), .Z(n39302) );
  AND U53221 ( .A(n39303), .B(n39302), .Z(n39307) );
  NAND U53222 ( .A(n39305), .B(n39304), .Z(n39306) );
  OR U53223 ( .A(n39307), .B(n39306), .Z(n39308) );
  AND U53224 ( .A(n39309), .B(n39308), .Z(n39313) );
  NAND U53225 ( .A(n39311), .B(n39310), .Z(n39312) );
  OR U53226 ( .A(n39313), .B(n39312), .Z(n39314) );
  AND U53227 ( .A(n39315), .B(n39314), .Z(n39319) );
  NAND U53228 ( .A(n39317), .B(n39316), .Z(n39318) );
  OR U53229 ( .A(n39319), .B(n39318), .Z(n39320) );
  AND U53230 ( .A(n39321), .B(n39320), .Z(n39322) );
  ANDN U53231 ( .B(n39323), .A(n39322), .Z(n39324) );
  OR U53232 ( .A(n39325), .B(n39324), .Z(n39326) );
  NAND U53233 ( .A(n39327), .B(n39326), .Z(n39328) );
  NANDN U53234 ( .A(n39329), .B(n39328), .Z(n39330) );
  OR U53235 ( .A(n39331), .B(n39330), .Z(n39332) );
  AND U53236 ( .A(n55975), .B(n39332), .Z(n39334) );
  NAND U53237 ( .A(n39334), .B(n39333), .Z(n39335) );
  NANDN U53238 ( .A(n39336), .B(n39335), .Z(n39337) );
  AND U53239 ( .A(n39338), .B(n39337), .Z(n39340) );
  NAND U53240 ( .A(n39340), .B(n39339), .Z(n39341) );
  NANDN U53241 ( .A(n39342), .B(n39341), .Z(n39343) );
  AND U53242 ( .A(n39344), .B(n39343), .Z(n39348) );
  NAND U53243 ( .A(n39346), .B(n39345), .Z(n39347) );
  OR U53244 ( .A(n39348), .B(n39347), .Z(n39349) );
  AND U53245 ( .A(n39350), .B(n39349), .Z(n39354) );
  NAND U53246 ( .A(n39352), .B(n39351), .Z(n39353) );
  OR U53247 ( .A(n39354), .B(n39353), .Z(n39355) );
  AND U53248 ( .A(n39356), .B(n39355), .Z(n39360) );
  NAND U53249 ( .A(n39358), .B(n39357), .Z(n39359) );
  OR U53250 ( .A(n39360), .B(n39359), .Z(n39361) );
  AND U53251 ( .A(n39362), .B(n39361), .Z(n39366) );
  NAND U53252 ( .A(n39364), .B(n39363), .Z(n39365) );
  OR U53253 ( .A(n39366), .B(n39365), .Z(n39367) );
  AND U53254 ( .A(n39368), .B(n39367), .Z(n39369) );
  NOR U53255 ( .A(n39370), .B(n39369), .Z(n39371) );
  NAND U53256 ( .A(n39372), .B(n39371), .Z(n39373) );
  NANDN U53257 ( .A(n39374), .B(n39373), .Z(n39375) );
  NAND U53258 ( .A(n39376), .B(n39375), .Z(n39377) );
  NANDN U53259 ( .A(n39378), .B(n39377), .Z(n39379) );
  AND U53260 ( .A(n39380), .B(n39379), .Z(n39382) );
  NAND U53261 ( .A(n39382), .B(n39381), .Z(n39383) );
  NANDN U53262 ( .A(n39384), .B(n39383), .Z(n39385) );
  AND U53263 ( .A(n39386), .B(n39385), .Z(n39388) );
  NAND U53264 ( .A(n39388), .B(n39387), .Z(n39389) );
  NANDN U53265 ( .A(n39390), .B(n39389), .Z(n39391) );
  AND U53266 ( .A(n39392), .B(n39391), .Z(n39394) );
  AND U53267 ( .A(n39394), .B(n39393), .Z(n39395) );
  OR U53268 ( .A(n39396), .B(n39395), .Z(n39397) );
  NAND U53269 ( .A(n39398), .B(n39397), .Z(n39399) );
  AND U53270 ( .A(n39400), .B(n39399), .Z(n39401) );
  NOR U53271 ( .A(n39402), .B(n39401), .Z(n39404) );
  NAND U53272 ( .A(n39404), .B(n39403), .Z(n39408) );
  NANDN U53273 ( .A(x[3750]), .B(y[3750]), .Z(n39405) );
  AND U53274 ( .A(n39406), .B(n39405), .Z(n39407) );
  NAND U53275 ( .A(n39408), .B(n39407), .Z(n39409) );
  NANDN U53276 ( .A(n39410), .B(n39409), .Z(n39411) );
  NAND U53277 ( .A(n39412), .B(n39411), .Z(n39413) );
  NAND U53278 ( .A(n39414), .B(n39413), .Z(n39415) );
  NANDN U53279 ( .A(n39416), .B(n39415), .Z(n39418) );
  ANDN U53280 ( .B(y[3754]), .A(x[3754]), .Z(n39417) );
  OR U53281 ( .A(n39418), .B(n39417), .Z(n39419) );
  NAND U53282 ( .A(n39420), .B(n39419), .Z(n39421) );
  NANDN U53283 ( .A(n39422), .B(n39421), .Z(n39424) );
  ANDN U53284 ( .B(y[3756]), .A(x[3756]), .Z(n39423) );
  OR U53285 ( .A(n39424), .B(n39423), .Z(n39425) );
  NAND U53286 ( .A(n39426), .B(n39425), .Z(n39427) );
  NANDN U53287 ( .A(n39428), .B(n39427), .Z(n39430) );
  OR U53288 ( .A(n39430), .B(n39429), .Z(n39431) );
  NAND U53289 ( .A(n39432), .B(n39431), .Z(n39436) );
  NAND U53290 ( .A(n39434), .B(n39433), .Z(n39435) );
  ANDN U53291 ( .B(n39436), .A(n39435), .Z(n39440) );
  NAND U53292 ( .A(n39438), .B(n39437), .Z(n39439) );
  OR U53293 ( .A(n39440), .B(n39439), .Z(n39441) );
  AND U53294 ( .A(n39442), .B(n39441), .Z(n39446) );
  NAND U53295 ( .A(n39444), .B(n39443), .Z(n39445) );
  OR U53296 ( .A(n39446), .B(n39445), .Z(n39447) );
  AND U53297 ( .A(n39448), .B(n39447), .Z(n39449) );
  NOR U53298 ( .A(n39450), .B(n39449), .Z(n39451) );
  NAND U53299 ( .A(n39452), .B(n39451), .Z(n39453) );
  NANDN U53300 ( .A(n39454), .B(n39453), .Z(n39455) );
  AND U53301 ( .A(n39456), .B(n39455), .Z(n39457) );
  OR U53302 ( .A(n39458), .B(n39457), .Z(n39459) );
  NAND U53303 ( .A(n39460), .B(n39459), .Z(n39463) );
  NAND U53304 ( .A(n39461), .B(n56016), .Z(n39462) );
  ANDN U53305 ( .B(n39463), .A(n39462), .Z(n39467) );
  NAND U53306 ( .A(n39465), .B(n39464), .Z(n39466) );
  OR U53307 ( .A(n39467), .B(n39466), .Z(n39468) );
  AND U53308 ( .A(n39469), .B(n39468), .Z(n39473) );
  NAND U53309 ( .A(n39471), .B(n39470), .Z(n39472) );
  OR U53310 ( .A(n39473), .B(n39472), .Z(n39474) );
  AND U53311 ( .A(n39475), .B(n39474), .Z(n39476) );
  OR U53312 ( .A(n39477), .B(n39476), .Z(n39478) );
  NAND U53313 ( .A(n39479), .B(n39478), .Z(n39480) );
  AND U53314 ( .A(n39481), .B(n39480), .Z(n39482) );
  NOR U53315 ( .A(n56024), .B(n39482), .Z(n39483) );
  NANDN U53316 ( .A(n56026), .B(n39483), .Z(n39484) );
  AND U53317 ( .A(n39485), .B(n39484), .Z(n39487) );
  NAND U53318 ( .A(n39487), .B(n39486), .Z(n39488) );
  NANDN U53319 ( .A(n39489), .B(n39488), .Z(n39490) );
  AND U53320 ( .A(n39491), .B(n39490), .Z(n39493) );
  NAND U53321 ( .A(n39493), .B(n39492), .Z(n39494) );
  NANDN U53322 ( .A(n39495), .B(n39494), .Z(n39496) );
  AND U53323 ( .A(n39497), .B(n39496), .Z(n39499) );
  AND U53324 ( .A(n39499), .B(n39498), .Z(n39503) );
  NAND U53325 ( .A(n39501), .B(n39500), .Z(n39502) );
  OR U53326 ( .A(n39503), .B(n39502), .Z(n39504) );
  AND U53327 ( .A(n39505), .B(n39504), .Z(n39506) );
  OR U53328 ( .A(n39507), .B(n39506), .Z(n39508) );
  NAND U53329 ( .A(n39509), .B(n39508), .Z(n39510) );
  AND U53330 ( .A(n39511), .B(n39510), .Z(n39512) );
  NOR U53331 ( .A(n39513), .B(n39512), .Z(n39515) );
  NAND U53332 ( .A(n39515), .B(n39514), .Z(n39519) );
  NANDN U53333 ( .A(x[3790]), .B(y[3790]), .Z(n39516) );
  AND U53334 ( .A(n39517), .B(n39516), .Z(n39518) );
  NAND U53335 ( .A(n39519), .B(n39518), .Z(n39520) );
  NANDN U53336 ( .A(n39521), .B(n39520), .Z(n39522) );
  NAND U53337 ( .A(n39523), .B(n39522), .Z(n39524) );
  NANDN U53338 ( .A(n39525), .B(n39524), .Z(n39526) );
  AND U53339 ( .A(n39527), .B(n39526), .Z(n39529) );
  NAND U53340 ( .A(n39529), .B(n39528), .Z(n39530) );
  NANDN U53341 ( .A(n39531), .B(n39530), .Z(n39532) );
  AND U53342 ( .A(n39533), .B(n39532), .Z(n39534) );
  NAND U53343 ( .A(n39534), .B(n51798), .Z(n39535) );
  NANDN U53344 ( .A(n39536), .B(n39535), .Z(n39537) );
  AND U53345 ( .A(n39538), .B(n39537), .Z(n39539) );
  OR U53346 ( .A(n39540), .B(n39539), .Z(n39541) );
  NAND U53347 ( .A(n56051), .B(n39541), .Z(n39542) );
  NANDN U53348 ( .A(n39543), .B(n39542), .Z(n39544) );
  OR U53349 ( .A(n39544), .B(n56050), .Z(n39545) );
  NAND U53350 ( .A(n39546), .B(n39545), .Z(n39547) );
  NANDN U53351 ( .A(n39548), .B(n39547), .Z(n39549) );
  AND U53352 ( .A(n39550), .B(n39549), .Z(n39551) );
  NAND U53353 ( .A(n39552), .B(n39551), .Z(n39556) );
  NAND U53354 ( .A(n39554), .B(n39553), .Z(n39555) );
  ANDN U53355 ( .B(n39556), .A(n39555), .Z(n39560) );
  NAND U53356 ( .A(n39558), .B(n39557), .Z(n39559) );
  OR U53357 ( .A(n39560), .B(n39559), .Z(n39561) );
  AND U53358 ( .A(n39562), .B(n39561), .Z(n39566) );
  NAND U53359 ( .A(n39564), .B(n39563), .Z(n39565) );
  OR U53360 ( .A(n39566), .B(n39565), .Z(n39567) );
  AND U53361 ( .A(n39568), .B(n39567), .Z(n39572) );
  NAND U53362 ( .A(n39570), .B(n39569), .Z(n39571) );
  OR U53363 ( .A(n39572), .B(n39571), .Z(n39573) );
  AND U53364 ( .A(n39574), .B(n39573), .Z(n39578) );
  NAND U53365 ( .A(n39576), .B(n39575), .Z(n39577) );
  OR U53366 ( .A(n39578), .B(n39577), .Z(n39579) );
  AND U53367 ( .A(n39580), .B(n39579), .Z(n39581) );
  ANDN U53368 ( .B(n39582), .A(n39581), .Z(n39583) );
  NAND U53369 ( .A(n39584), .B(n39583), .Z(n39585) );
  NANDN U53370 ( .A(n39586), .B(n39585), .Z(n39587) );
  OR U53371 ( .A(n39588), .B(n39587), .Z(n39589) );
  AND U53372 ( .A(n39590), .B(n39589), .Z(n39592) );
  NAND U53373 ( .A(n39592), .B(n39591), .Z(n39593) );
  NANDN U53374 ( .A(n39594), .B(n39593), .Z(n39595) );
  AND U53375 ( .A(n39596), .B(n39595), .Z(n39598) );
  NANDN U53376 ( .A(x[3818]), .B(y[3818]), .Z(n39597) );
  AND U53377 ( .A(n39598), .B(n39597), .Z(n39599) );
  OR U53378 ( .A(n39600), .B(n39599), .Z(n39601) );
  AND U53379 ( .A(n39602), .B(n39601), .Z(n39606) );
  NAND U53380 ( .A(n39604), .B(n39603), .Z(n39605) );
  OR U53381 ( .A(n39606), .B(n39605), .Z(n39607) );
  AND U53382 ( .A(n39608), .B(n39607), .Z(n39612) );
  NAND U53383 ( .A(n39610), .B(n39609), .Z(n39611) );
  OR U53384 ( .A(n39612), .B(n39611), .Z(n39613) );
  AND U53385 ( .A(n39614), .B(n39613), .Z(n39618) );
  NAND U53386 ( .A(n39616), .B(n39615), .Z(n39617) );
  OR U53387 ( .A(n39618), .B(n39617), .Z(n39619) );
  AND U53388 ( .A(n39620), .B(n39619), .Z(n39624) );
  NAND U53389 ( .A(n39622), .B(n39621), .Z(n39623) );
  OR U53390 ( .A(n39624), .B(n39623), .Z(n39625) );
  AND U53391 ( .A(n39626), .B(n39625), .Z(n39630) );
  NAND U53392 ( .A(n39628), .B(n39627), .Z(n39629) );
  OR U53393 ( .A(n39630), .B(n39629), .Z(n39631) );
  AND U53394 ( .A(n39632), .B(n39631), .Z(n39633) );
  OR U53395 ( .A(n39634), .B(n39633), .Z(n39635) );
  NAND U53396 ( .A(n39636), .B(n39635), .Z(n39637) );
  AND U53397 ( .A(n39638), .B(n39637), .Z(n39639) );
  NOR U53398 ( .A(n51785), .B(n39639), .Z(n39640) );
  NAND U53399 ( .A(n56080), .B(n39640), .Z(n39641) );
  AND U53400 ( .A(n39642), .B(n39641), .Z(n39644) );
  NAND U53401 ( .A(n39644), .B(n39643), .Z(n39645) );
  NANDN U53402 ( .A(n39646), .B(n39645), .Z(n39647) );
  AND U53403 ( .A(n39648), .B(n39647), .Z(n39650) );
  NAND U53404 ( .A(n39650), .B(n39649), .Z(n39651) );
  NANDN U53405 ( .A(n39652), .B(n39651), .Z(n39653) );
  AND U53406 ( .A(n39654), .B(n39653), .Z(n39656) );
  NAND U53407 ( .A(n39656), .B(n39655), .Z(n39657) );
  AND U53408 ( .A(n39657), .B(n56090), .Z(n39658) );
  NANDN U53409 ( .A(x[3840]), .B(y[3840]), .Z(n56087) );
  AND U53410 ( .A(n39658), .B(n56087), .Z(n39662) );
  AND U53411 ( .A(n39660), .B(n39659), .Z(n39661) );
  NANDN U53412 ( .A(n39662), .B(n39661), .Z(n39665) );
  NANDN U53413 ( .A(x[3842]), .B(y[3842]), .Z(n56091) );
  AND U53414 ( .A(n39663), .B(n56091), .Z(n39664) );
  NAND U53415 ( .A(n39665), .B(n39664), .Z(n39666) );
  NANDN U53416 ( .A(n39667), .B(n39666), .Z(n39668) );
  NAND U53417 ( .A(n39669), .B(n39668), .Z(n39670) );
  NANDN U53418 ( .A(n39671), .B(n39670), .Z(n39672) );
  AND U53419 ( .A(n39673), .B(n39672), .Z(n39675) );
  NAND U53420 ( .A(n39675), .B(n39674), .Z(n39676) );
  NANDN U53421 ( .A(n39677), .B(n39676), .Z(n39678) );
  AND U53422 ( .A(n39679), .B(n39678), .Z(n39680) );
  NANDN U53423 ( .A(n39681), .B(n39680), .Z(n39682) );
  AND U53424 ( .A(n39683), .B(n39682), .Z(n39684) );
  NANDN U53425 ( .A(n39685), .B(n39684), .Z(n39686) );
  AND U53426 ( .A(n39687), .B(n39686), .Z(n39688) );
  OR U53427 ( .A(n39689), .B(n39688), .Z(n39690) );
  NAND U53428 ( .A(n39691), .B(n39690), .Z(n39692) );
  AND U53429 ( .A(n39693), .B(n39692), .Z(n39694) );
  NOR U53430 ( .A(n56102), .B(n39694), .Z(n39695) );
  NANDN U53431 ( .A(n39696), .B(n39695), .Z(n39697) );
  AND U53432 ( .A(n39698), .B(n39697), .Z(n39700) );
  NAND U53433 ( .A(n39700), .B(n39699), .Z(n39701) );
  NANDN U53434 ( .A(n39702), .B(n39701), .Z(n39703) );
  AND U53435 ( .A(n39704), .B(n39703), .Z(n39706) );
  NAND U53436 ( .A(n39706), .B(n39705), .Z(n39707) );
  NANDN U53437 ( .A(n39708), .B(n39707), .Z(n39709) );
  AND U53438 ( .A(n39710), .B(n39709), .Z(n39712) );
  NAND U53439 ( .A(n39712), .B(n39711), .Z(n39713) );
  NANDN U53440 ( .A(n39714), .B(n39713), .Z(n39715) );
  AND U53441 ( .A(n39716), .B(n39715), .Z(n39718) );
  NAND U53442 ( .A(n39718), .B(n39717), .Z(n39722) );
  NANDN U53443 ( .A(x[3862]), .B(y[3862]), .Z(n39719) );
  AND U53444 ( .A(n39720), .B(n39719), .Z(n39721) );
  NAND U53445 ( .A(n39722), .B(n39721), .Z(n39723) );
  NANDN U53446 ( .A(n39724), .B(n39723), .Z(n39725) );
  NAND U53447 ( .A(n39726), .B(n39725), .Z(n39727) );
  NANDN U53448 ( .A(n39728), .B(n39727), .Z(n39729) );
  AND U53449 ( .A(n39730), .B(n39729), .Z(n39732) );
  NAND U53450 ( .A(n39732), .B(n39731), .Z(n39733) );
  NANDN U53451 ( .A(n39734), .B(n39733), .Z(n39735) );
  AND U53452 ( .A(n39736), .B(n39735), .Z(n39737) );
  NANDN U53453 ( .A(n39738), .B(n39737), .Z(n39739) );
  NAND U53454 ( .A(n39740), .B(n39739), .Z(n39741) );
  NANDN U53455 ( .A(n39742), .B(n39741), .Z(n39743) );
  AND U53456 ( .A(n39744), .B(n39743), .Z(n39745) );
  NAND U53457 ( .A(n39746), .B(n39745), .Z(n39749) );
  NAND U53458 ( .A(n39747), .B(n56121), .Z(n39748) );
  ANDN U53459 ( .B(n39749), .A(n39748), .Z(n39753) );
  NAND U53460 ( .A(n39751), .B(n39750), .Z(n39752) );
  OR U53461 ( .A(n39753), .B(n39752), .Z(n39754) );
  AND U53462 ( .A(n39755), .B(n39754), .Z(n39756) );
  OR U53463 ( .A(n39757), .B(n39756), .Z(n39758) );
  NAND U53464 ( .A(n39759), .B(n39758), .Z(n39760) );
  AND U53465 ( .A(n39761), .B(n39760), .Z(n39762) );
  ANDN U53466 ( .B(n51775), .A(n39762), .Z(n39763) );
  NANDN U53467 ( .A(n56127), .B(n39763), .Z(n39764) );
  AND U53468 ( .A(n39765), .B(n39764), .Z(n39767) );
  NAND U53469 ( .A(n39767), .B(n39766), .Z(n39768) );
  NANDN U53470 ( .A(n39769), .B(n39768), .Z(n39770) );
  AND U53471 ( .A(n39771), .B(n39770), .Z(n39773) );
  NAND U53472 ( .A(n39773), .B(n39772), .Z(n39774) );
  NANDN U53473 ( .A(n39775), .B(n39774), .Z(n39776) );
  AND U53474 ( .A(n39777), .B(n39776), .Z(n39778) );
  OR U53475 ( .A(n39779), .B(n39778), .Z(n39780) );
  NAND U53476 ( .A(n39781), .B(n39780), .Z(n39782) );
  AND U53477 ( .A(n39783), .B(n39782), .Z(n39787) );
  AND U53478 ( .A(n39785), .B(n39784), .Z(n39786) );
  NANDN U53479 ( .A(n39787), .B(n39786), .Z(n39790) );
  NANDN U53480 ( .A(x[3888]), .B(y[3888]), .Z(n56137) );
  AND U53481 ( .A(n39788), .B(n56137), .Z(n39789) );
  NAND U53482 ( .A(n39790), .B(n39789), .Z(n39791) );
  NANDN U53483 ( .A(n39792), .B(n39791), .Z(n39793) );
  NAND U53484 ( .A(n39794), .B(n39793), .Z(n39795) );
  NAND U53485 ( .A(n39796), .B(n39795), .Z(n39797) );
  NANDN U53486 ( .A(n39798), .B(n39797), .Z(n39800) );
  OR U53487 ( .A(n39800), .B(n39799), .Z(n39801) );
  NAND U53488 ( .A(n39802), .B(n39801), .Z(n39804) );
  ANDN U53489 ( .B(n39804), .A(n39803), .Z(n39806) );
  NAND U53490 ( .A(n39806), .B(n39805), .Z(n39807) );
  NANDN U53491 ( .A(n39808), .B(n39807), .Z(n39809) );
  AND U53492 ( .A(n39810), .B(n39809), .Z(n39811) );
  NANDN U53493 ( .A(n39812), .B(n39811), .Z(n39813) );
  NAND U53494 ( .A(n39814), .B(n39813), .Z(n39815) );
  NANDN U53495 ( .A(n39816), .B(n39815), .Z(n39817) );
  AND U53496 ( .A(n39818), .B(n39817), .Z(n39819) );
  NAND U53497 ( .A(n39820), .B(n39819), .Z(n39824) );
  NAND U53498 ( .A(n39822), .B(n39821), .Z(n39823) );
  ANDN U53499 ( .B(n39824), .A(n39823), .Z(n39828) );
  NAND U53500 ( .A(n39826), .B(n39825), .Z(n39827) );
  OR U53501 ( .A(n39828), .B(n39827), .Z(n39829) );
  AND U53502 ( .A(n39830), .B(n39829), .Z(n39834) );
  NAND U53503 ( .A(n39832), .B(n39831), .Z(n39833) );
  OR U53504 ( .A(n39834), .B(n39833), .Z(n39835) );
  AND U53505 ( .A(n39836), .B(n39835), .Z(n39840) );
  NAND U53506 ( .A(n39838), .B(n39837), .Z(n39839) );
  OR U53507 ( .A(n39840), .B(n39839), .Z(n39841) );
  AND U53508 ( .A(n39842), .B(n39841), .Z(n39846) );
  NAND U53509 ( .A(n39844), .B(n39843), .Z(n39845) );
  OR U53510 ( .A(n39846), .B(n39845), .Z(n39847) );
  AND U53511 ( .A(n39848), .B(n39847), .Z(n39852) );
  NAND U53512 ( .A(n39850), .B(n39849), .Z(n39851) );
  OR U53513 ( .A(n39852), .B(n39851), .Z(n39853) );
  AND U53514 ( .A(n39854), .B(n39853), .Z(n39855) );
  NOR U53515 ( .A(n39856), .B(n39855), .Z(n39857) );
  NAND U53516 ( .A(n39858), .B(n39857), .Z(n39859) );
  NANDN U53517 ( .A(n39860), .B(n39859), .Z(n39861) );
  NAND U53518 ( .A(n39862), .B(n39861), .Z(n39863) );
  NANDN U53519 ( .A(n39864), .B(n39863), .Z(n39865) );
  AND U53520 ( .A(n39866), .B(n39865), .Z(n39868) );
  NAND U53521 ( .A(n39868), .B(n39867), .Z(n39869) );
  NANDN U53522 ( .A(n39870), .B(n39869), .Z(n39871) );
  AND U53523 ( .A(n39872), .B(n39871), .Z(n39874) );
  NAND U53524 ( .A(n39874), .B(n39873), .Z(n39875) );
  NANDN U53525 ( .A(n39876), .B(n39875), .Z(n39877) );
  AND U53526 ( .A(n39878), .B(n39877), .Z(n39880) );
  AND U53527 ( .A(n39880), .B(n39879), .Z(n39884) );
  NAND U53528 ( .A(n39882), .B(n39881), .Z(n39883) );
  OR U53529 ( .A(n39884), .B(n39883), .Z(n39885) );
  AND U53530 ( .A(n39886), .B(n39885), .Z(n39890) );
  NAND U53531 ( .A(n39888), .B(n39887), .Z(n39889) );
  OR U53532 ( .A(n39890), .B(n39889), .Z(n39891) );
  AND U53533 ( .A(n39892), .B(n39891), .Z(n39896) );
  NAND U53534 ( .A(n39894), .B(n39893), .Z(n39895) );
  OR U53535 ( .A(n39896), .B(n39895), .Z(n39897) );
  AND U53536 ( .A(n39898), .B(n39897), .Z(n39902) );
  NAND U53537 ( .A(n39900), .B(n39899), .Z(n39901) );
  OR U53538 ( .A(n39902), .B(n39901), .Z(n39903) );
  AND U53539 ( .A(n39904), .B(n39903), .Z(n39905) );
  OR U53540 ( .A(n39906), .B(n39905), .Z(n39907) );
  NAND U53541 ( .A(n39908), .B(n39907), .Z(n39909) );
  AND U53542 ( .A(n39910), .B(n39909), .Z(n39911) );
  NOR U53543 ( .A(n39912), .B(n39911), .Z(n39914) );
  NAND U53544 ( .A(n39914), .B(n39913), .Z(n39915) );
  AND U53545 ( .A(n39915), .B(n56178), .Z(n39916) );
  NANDN U53546 ( .A(x[3932]), .B(y[3932]), .Z(n51762) );
  AND U53547 ( .A(n39916), .B(n51762), .Z(n39920) );
  AND U53548 ( .A(n39918), .B(n39917), .Z(n39919) );
  NANDN U53549 ( .A(n39920), .B(n39919), .Z(n39923) );
  NANDN U53550 ( .A(x[3934]), .B(y[3934]), .Z(n56179) );
  AND U53551 ( .A(n39921), .B(n56179), .Z(n39922) );
  NAND U53552 ( .A(n39923), .B(n39922), .Z(n39924) );
  NANDN U53553 ( .A(n39925), .B(n39924), .Z(n39926) );
  NAND U53554 ( .A(n39927), .B(n39926), .Z(n39928) );
  NANDN U53555 ( .A(n39929), .B(n39928), .Z(n39930) );
  AND U53556 ( .A(n39931), .B(n39930), .Z(n39933) );
  NAND U53557 ( .A(n39933), .B(n39932), .Z(n39934) );
  NANDN U53558 ( .A(n39935), .B(n39934), .Z(n39936) );
  AND U53559 ( .A(n39937), .B(n39936), .Z(n39939) );
  NAND U53560 ( .A(n39939), .B(n39938), .Z(n39940) );
  AND U53561 ( .A(n39941), .B(n39940), .Z(n39942) );
  OR U53562 ( .A(n39943), .B(n39942), .Z(n39944) );
  NAND U53563 ( .A(n39945), .B(n39944), .Z(n39946) );
  NANDN U53564 ( .A(n39947), .B(n39946), .Z(n39949) );
  ANDN U53565 ( .B(y[3944]), .A(x[3944]), .Z(n39948) );
  OR U53566 ( .A(n39949), .B(n39948), .Z(n39950) );
  NAND U53567 ( .A(n39951), .B(n39950), .Z(n39952) );
  NANDN U53568 ( .A(n39953), .B(n39952), .Z(n39955) );
  ANDN U53569 ( .B(y[3946]), .A(x[3946]), .Z(n39954) );
  OR U53570 ( .A(n39955), .B(n39954), .Z(n39956) );
  NANDN U53571 ( .A(n39957), .B(n39956), .Z(n39958) );
  AND U53572 ( .A(n39959), .B(n39958), .Z(n39960) );
  OR U53573 ( .A(n39961), .B(n39960), .Z(n39962) );
  NAND U53574 ( .A(n39963), .B(n39962), .Z(n39964) );
  NAND U53575 ( .A(n39965), .B(n39964), .Z(n39966) );
  NAND U53576 ( .A(n51753), .B(n39966), .Z(n39967) );
  AND U53577 ( .A(n39968), .B(n39967), .Z(n39969) );
  NAND U53578 ( .A(n51752), .B(n39969), .Z(n39970) );
  NANDN U53579 ( .A(n39971), .B(n39970), .Z(n39972) );
  AND U53580 ( .A(n39973), .B(n39972), .Z(n39975) );
  NAND U53581 ( .A(n39975), .B(n39974), .Z(n39976) );
  AND U53582 ( .A(n39977), .B(n39976), .Z(n39978) );
  NOR U53583 ( .A(n39979), .B(n39978), .Z(n39981) );
  NAND U53584 ( .A(n39981), .B(n39980), .Z(n39984) );
  NANDN U53585 ( .A(x[3958]), .B(y[3958]), .Z(n56200) );
  AND U53586 ( .A(n39982), .B(n56200), .Z(n39983) );
  NAND U53587 ( .A(n39984), .B(n39983), .Z(n39985) );
  NANDN U53588 ( .A(n39986), .B(n39985), .Z(n39987) );
  NAND U53589 ( .A(n39988), .B(n39987), .Z(n39989) );
  NANDN U53590 ( .A(n39990), .B(n39989), .Z(n39991) );
  AND U53591 ( .A(n56206), .B(n39991), .Z(n39993) );
  NAND U53592 ( .A(n39993), .B(n39992), .Z(n39994) );
  NANDN U53593 ( .A(n39995), .B(n39994), .Z(n39996) );
  AND U53594 ( .A(n39997), .B(n39996), .Z(n39998) );
  NANDN U53595 ( .A(n56207), .B(n39998), .Z(n39999) );
  NAND U53596 ( .A(n40000), .B(n39999), .Z(n40001) );
  NANDN U53597 ( .A(n40002), .B(n40001), .Z(n40003) );
  AND U53598 ( .A(n40004), .B(n40003), .Z(n40005) );
  NAND U53599 ( .A(n40006), .B(n40005), .Z(n40010) );
  NAND U53600 ( .A(n40008), .B(n40007), .Z(n40009) );
  ANDN U53601 ( .B(n40010), .A(n40009), .Z(n40014) );
  NAND U53602 ( .A(n40012), .B(n40011), .Z(n40013) );
  OR U53603 ( .A(n40014), .B(n40013), .Z(n40015) );
  AND U53604 ( .A(n40016), .B(n40015), .Z(n40017) );
  OR U53605 ( .A(n40018), .B(n40017), .Z(n40019) );
  NAND U53606 ( .A(n40020), .B(n40019), .Z(n40021) );
  AND U53607 ( .A(n40022), .B(n40021), .Z(n40023) );
  NOR U53608 ( .A(n40024), .B(n40023), .Z(n40025) );
  NANDN U53609 ( .A(n40026), .B(n40025), .Z(n40027) );
  AND U53610 ( .A(n40028), .B(n40027), .Z(n40030) );
  NAND U53611 ( .A(n40030), .B(n40029), .Z(n40031) );
  NANDN U53612 ( .A(n40032), .B(n40031), .Z(n40033) );
  AND U53613 ( .A(n40034), .B(n40033), .Z(n40036) );
  NAND U53614 ( .A(n40036), .B(n40035), .Z(n40037) );
  NANDN U53615 ( .A(n40038), .B(n40037), .Z(n40039) );
  AND U53616 ( .A(n40040), .B(n40039), .Z(n40042) );
  NAND U53617 ( .A(n40042), .B(n40041), .Z(n40043) );
  NANDN U53618 ( .A(n40044), .B(n40043), .Z(n40045) );
  AND U53619 ( .A(n40046), .B(n40045), .Z(n40048) );
  NAND U53620 ( .A(n40048), .B(n40047), .Z(n40049) );
  NAND U53621 ( .A(n40050), .B(n40049), .Z(n40051) );
  NANDN U53622 ( .A(n40052), .B(n40051), .Z(n40053) );
  NANDN U53623 ( .A(x[3984]), .B(y[3984]), .Z(n56226) );
  AND U53624 ( .A(n40053), .B(n56226), .Z(n40055) );
  NAND U53625 ( .A(n40055), .B(n40054), .Z(n40056) );
  NANDN U53626 ( .A(n40057), .B(n40056), .Z(n40058) );
  AND U53627 ( .A(n51745), .B(n40058), .Z(n40059) );
  NANDN U53628 ( .A(n40060), .B(n40059), .Z(n40061) );
  NAND U53629 ( .A(n40062), .B(n40061), .Z(n40063) );
  NANDN U53630 ( .A(n40064), .B(n40063), .Z(n40065) );
  AND U53631 ( .A(n40066), .B(n40065), .Z(n40069) );
  AND U53632 ( .A(n40067), .B(n56235), .Z(n40068) );
  NANDN U53633 ( .A(n40069), .B(n40068), .Z(n40070) );
  NANDN U53634 ( .A(n40071), .B(n40070), .Z(n40072) );
  AND U53635 ( .A(n51743), .B(n40072), .Z(n40073) );
  NANDN U53636 ( .A(x[3992]), .B(y[3992]), .Z(n56236) );
  AND U53637 ( .A(n40073), .B(n56236), .Z(n40077) );
  NAND U53638 ( .A(n40075), .B(n40074), .Z(n40076) );
  OR U53639 ( .A(n40077), .B(n40076), .Z(n40078) );
  AND U53640 ( .A(n40079), .B(n40078), .Z(n40080) );
  OR U53641 ( .A(n40081), .B(n40080), .Z(n40082) );
  NAND U53642 ( .A(n40083), .B(n40082), .Z(n40084) );
  AND U53643 ( .A(n40085), .B(n40084), .Z(n40086) );
  ANDN U53644 ( .B(n51741), .A(n40086), .Z(n40087) );
  NAND U53645 ( .A(n56242), .B(n40087), .Z(n40088) );
  NANDN U53646 ( .A(n40089), .B(n40088), .Z(n40091) );
  OR U53647 ( .A(n40091), .B(n40090), .Z(n40092) );
  NAND U53648 ( .A(n40093), .B(n40092), .Z(n40094) );
  NANDN U53649 ( .A(n40095), .B(n40094), .Z(n40098) );
  NANDN U53650 ( .A(x[4002]), .B(y[4002]), .Z(n56246) );
  AND U53651 ( .A(n40096), .B(n56246), .Z(n40097) );
  NAND U53652 ( .A(n40098), .B(n40097), .Z(n40099) );
  NANDN U53653 ( .A(n40100), .B(n40099), .Z(n40101) );
  NAND U53654 ( .A(n40102), .B(n40101), .Z(n40103) );
  NANDN U53655 ( .A(n40104), .B(n40103), .Z(n40105) );
  AND U53656 ( .A(n40106), .B(n40105), .Z(n40108) );
  NAND U53657 ( .A(n40108), .B(n40107), .Z(n40109) );
  NANDN U53658 ( .A(n40110), .B(n40109), .Z(n40111) );
  AND U53659 ( .A(n40112), .B(n40111), .Z(n40113) );
  NANDN U53660 ( .A(n40114), .B(n40113), .Z(n40115) );
  NAND U53661 ( .A(n40116), .B(n40115), .Z(n40117) );
  NANDN U53662 ( .A(n40118), .B(n40117), .Z(n40120) );
  OR U53663 ( .A(n40120), .B(n40119), .Z(n40121) );
  NAND U53664 ( .A(n40122), .B(n40121), .Z(n40126) );
  NANDN U53665 ( .A(x[4012]), .B(y[4012]), .Z(n40124) );
  NAND U53666 ( .A(n40124), .B(n40123), .Z(n40125) );
  ANDN U53667 ( .B(n40126), .A(n40125), .Z(n40130) );
  NAND U53668 ( .A(n40128), .B(n40127), .Z(n40129) );
  OR U53669 ( .A(n40130), .B(n40129), .Z(n40131) );
  AND U53670 ( .A(n40132), .B(n40131), .Z(n40136) );
  NAND U53671 ( .A(n40134), .B(n40133), .Z(n40135) );
  OR U53672 ( .A(n40136), .B(n40135), .Z(n40137) );
  AND U53673 ( .A(n40138), .B(n40137), .Z(n40142) );
  NAND U53674 ( .A(n40140), .B(n40139), .Z(n40141) );
  OR U53675 ( .A(n40142), .B(n40141), .Z(n40143) );
  AND U53676 ( .A(n40144), .B(n40143), .Z(n40148) );
  NAND U53677 ( .A(n40146), .B(n40145), .Z(n40147) );
  OR U53678 ( .A(n40148), .B(n40147), .Z(n40149) );
  AND U53679 ( .A(n40150), .B(n40149), .Z(n40154) );
  NAND U53680 ( .A(n40152), .B(n40151), .Z(n40153) );
  OR U53681 ( .A(n40154), .B(n40153), .Z(n40155) );
  AND U53682 ( .A(n40156), .B(n40155), .Z(n40160) );
  NAND U53683 ( .A(n40158), .B(n40157), .Z(n40159) );
  OR U53684 ( .A(n40160), .B(n40159), .Z(n40161) );
  AND U53685 ( .A(n40162), .B(n40161), .Z(n40166) );
  NAND U53686 ( .A(n40164), .B(n40163), .Z(n40165) );
  OR U53687 ( .A(n40166), .B(n40165), .Z(n40167) );
  AND U53688 ( .A(n40168), .B(n40167), .Z(n40169) );
  OR U53689 ( .A(n40170), .B(n40169), .Z(n40171) );
  NAND U53690 ( .A(n40172), .B(n40171), .Z(n40173) );
  NAND U53691 ( .A(n40174), .B(n40173), .Z(n40175) );
  AND U53692 ( .A(n40176), .B(n40175), .Z(n40180) );
  NAND U53693 ( .A(n40178), .B(n40177), .Z(n40179) );
  OR U53694 ( .A(n40180), .B(n40179), .Z(n40181) );
  AND U53695 ( .A(n40182), .B(n40181), .Z(n40186) );
  NAND U53696 ( .A(n40184), .B(n40183), .Z(n40185) );
  OR U53697 ( .A(n40186), .B(n40185), .Z(n40187) );
  AND U53698 ( .A(n40188), .B(n40187), .Z(n40192) );
  NAND U53699 ( .A(n40190), .B(n40189), .Z(n40191) );
  OR U53700 ( .A(n40192), .B(n40191), .Z(n40193) );
  AND U53701 ( .A(n40194), .B(n40193), .Z(n40195) );
  NOR U53702 ( .A(n40196), .B(n40195), .Z(n40197) );
  NAND U53703 ( .A(n40198), .B(n40197), .Z(n40199) );
  NANDN U53704 ( .A(n40200), .B(n40199), .Z(n40201) );
  NAND U53705 ( .A(n40202), .B(n40201), .Z(n40203) );
  NANDN U53706 ( .A(n40204), .B(n40203), .Z(n40205) );
  AND U53707 ( .A(n40206), .B(n40205), .Z(n40208) );
  NAND U53708 ( .A(n40208), .B(n40207), .Z(n40209) );
  NANDN U53709 ( .A(n40210), .B(n40209), .Z(n40211) );
  AND U53710 ( .A(n40212), .B(n40211), .Z(n40214) );
  NAND U53711 ( .A(n40214), .B(n40213), .Z(n40215) );
  NANDN U53712 ( .A(n40216), .B(n40215), .Z(n40217) );
  AND U53713 ( .A(n40218), .B(n40217), .Z(n40220) );
  NAND U53714 ( .A(n40220), .B(n40219), .Z(n40224) );
  NANDN U53715 ( .A(x[4046]), .B(y[4046]), .Z(n40221) );
  AND U53716 ( .A(n40222), .B(n40221), .Z(n40223) );
  NAND U53717 ( .A(n40224), .B(n40223), .Z(n40225) );
  NANDN U53718 ( .A(n40226), .B(n40225), .Z(n40227) );
  NAND U53719 ( .A(n40228), .B(n40227), .Z(n40229) );
  NANDN U53720 ( .A(n40230), .B(n40229), .Z(n40231) );
  AND U53721 ( .A(n40232), .B(n40231), .Z(n40234) );
  NAND U53722 ( .A(n40234), .B(n40233), .Z(n40235) );
  NANDN U53723 ( .A(n40236), .B(n40235), .Z(n40237) );
  AND U53724 ( .A(n40238), .B(n40237), .Z(n40240) );
  NANDN U53725 ( .A(x[4052]), .B(y[4052]), .Z(n40239) );
  NAND U53726 ( .A(n40240), .B(n40239), .Z(n40241) );
  NANDN U53727 ( .A(n40242), .B(n40241), .Z(n40243) );
  AND U53728 ( .A(n40244), .B(n40243), .Z(n40246) );
  AND U53729 ( .A(n40246), .B(n40245), .Z(n40250) );
  NAND U53730 ( .A(n40248), .B(n40247), .Z(n40249) );
  OR U53731 ( .A(n40250), .B(n40249), .Z(n40251) );
  AND U53732 ( .A(n40252), .B(n40251), .Z(n40256) );
  NAND U53733 ( .A(n40254), .B(n40253), .Z(n40255) );
  OR U53734 ( .A(n40256), .B(n40255), .Z(n40257) );
  AND U53735 ( .A(n40258), .B(n40257), .Z(n40260) );
  AND U53736 ( .A(n40260), .B(n40259), .Z(n40264) );
  NAND U53737 ( .A(n40262), .B(n40261), .Z(n40263) );
  OR U53738 ( .A(n40264), .B(n40263), .Z(n40265) );
  AND U53739 ( .A(n40266), .B(n40265), .Z(n40270) );
  NAND U53740 ( .A(n40268), .B(n40267), .Z(n40269) );
  OR U53741 ( .A(n40270), .B(n40269), .Z(n40271) );
  AND U53742 ( .A(n40272), .B(n40271), .Z(n40273) );
  NOR U53743 ( .A(n40274), .B(n40273), .Z(n40275) );
  NAND U53744 ( .A(n40276), .B(n40275), .Z(n40277) );
  NANDN U53745 ( .A(n40278), .B(n40277), .Z(n40279) );
  NAND U53746 ( .A(n40280), .B(n40279), .Z(n40281) );
  NANDN U53747 ( .A(n40282), .B(n40281), .Z(n40283) );
  AND U53748 ( .A(n40284), .B(n40283), .Z(n40286) );
  NAND U53749 ( .A(n40286), .B(n40285), .Z(n40287) );
  NANDN U53750 ( .A(n40288), .B(n40287), .Z(n40289) );
  AND U53751 ( .A(n40290), .B(n40289), .Z(n40292) );
  NAND U53752 ( .A(n40292), .B(n40291), .Z(n40293) );
  NANDN U53753 ( .A(n40294), .B(n40293), .Z(n40295) );
  AND U53754 ( .A(n40296), .B(n40295), .Z(n40298) );
  NAND U53755 ( .A(n40298), .B(n40297), .Z(n40299) );
  NANDN U53756 ( .A(n40300), .B(n40299), .Z(n40301) );
  AND U53757 ( .A(n40302), .B(n40301), .Z(n40304) );
  AND U53758 ( .A(n40304), .B(n40303), .Z(n40308) );
  NAND U53759 ( .A(n40306), .B(n40305), .Z(n40307) );
  OR U53760 ( .A(n40308), .B(n40307), .Z(n40309) );
  AND U53761 ( .A(n40310), .B(n40309), .Z(n40311) );
  OR U53762 ( .A(n40312), .B(n40311), .Z(n40313) );
  NAND U53763 ( .A(n40314), .B(n40313), .Z(n40315) );
  AND U53764 ( .A(n40316), .B(n40315), .Z(n40317) );
  NOR U53765 ( .A(n40318), .B(n40317), .Z(n40320) );
  NAND U53766 ( .A(n40320), .B(n40319), .Z(n40321) );
  AND U53767 ( .A(n40321), .B(n56320), .Z(n40322) );
  NANDN U53768 ( .A(n40323), .B(n40322), .Z(n40324) );
  NAND U53769 ( .A(n40325), .B(n40324), .Z(n40326) );
  NANDN U53770 ( .A(n56321), .B(n40326), .Z(n40327) );
  ANDN U53771 ( .B(y[4082]), .A(x[4082]), .Z(n56319) );
  OR U53772 ( .A(n40327), .B(n56319), .Z(n40328) );
  NAND U53773 ( .A(n40329), .B(n40328), .Z(n40330) );
  NANDN U53774 ( .A(n40331), .B(n40330), .Z(n40332) );
  ANDN U53775 ( .B(y[4084]), .A(x[4084]), .Z(n51716) );
  OR U53776 ( .A(n40332), .B(n51716), .Z(n40333) );
  NAND U53777 ( .A(n40334), .B(n40333), .Z(n40335) );
  NANDN U53778 ( .A(n40336), .B(n40335), .Z(n40337) );
  ANDN U53779 ( .B(n40338), .A(n40337), .Z(n40342) );
  NAND U53780 ( .A(n40340), .B(n40339), .Z(n40341) );
  OR U53781 ( .A(n40342), .B(n40341), .Z(n40343) );
  AND U53782 ( .A(n40344), .B(n40343), .Z(n40348) );
  NAND U53783 ( .A(n40346), .B(n40345), .Z(n40347) );
  OR U53784 ( .A(n40348), .B(n40347), .Z(n40349) );
  AND U53785 ( .A(n40350), .B(n40349), .Z(n40351) );
  OR U53786 ( .A(n40352), .B(n40351), .Z(n40353) );
  NAND U53787 ( .A(n40354), .B(n40353), .Z(n40355) );
  NAND U53788 ( .A(n40356), .B(n40355), .Z(n40357) );
  NANDN U53789 ( .A(n40358), .B(n40357), .Z(n40359) );
  AND U53790 ( .A(n40360), .B(n40359), .Z(n40362) );
  NAND U53791 ( .A(n40362), .B(n40361), .Z(n40363) );
  NANDN U53792 ( .A(n40364), .B(n40363), .Z(n40365) );
  AND U53793 ( .A(n40366), .B(n40365), .Z(n40368) );
  NAND U53794 ( .A(n40368), .B(n40367), .Z(n40369) );
  NANDN U53795 ( .A(n40370), .B(n40369), .Z(n40371) );
  AND U53796 ( .A(n40372), .B(n40371), .Z(n40374) );
  AND U53797 ( .A(n40374), .B(n40373), .Z(n40378) );
  NAND U53798 ( .A(n40376), .B(n40375), .Z(n40377) );
  OR U53799 ( .A(n40378), .B(n40377), .Z(n40379) );
  AND U53800 ( .A(n40380), .B(n40379), .Z(n40384) );
  NAND U53801 ( .A(n40382), .B(n40381), .Z(n40383) );
  OR U53802 ( .A(n40384), .B(n40383), .Z(n40385) );
  AND U53803 ( .A(n40386), .B(n40385), .Z(n40390) );
  NAND U53804 ( .A(n40388), .B(n40387), .Z(n40389) );
  OR U53805 ( .A(n40390), .B(n40389), .Z(n40391) );
  AND U53806 ( .A(n40392), .B(n40391), .Z(n40396) );
  NAND U53807 ( .A(n40394), .B(n40393), .Z(n40395) );
  OR U53808 ( .A(n40396), .B(n40395), .Z(n40397) );
  AND U53809 ( .A(n40398), .B(n40397), .Z(n40402) );
  NANDN U53810 ( .A(x[4108]), .B(y[4108]), .Z(n40400) );
  NAND U53811 ( .A(n40400), .B(n40399), .Z(n40401) );
  OR U53812 ( .A(n40402), .B(n40401), .Z(n40403) );
  AND U53813 ( .A(n40404), .B(n40403), .Z(n40408) );
  NAND U53814 ( .A(n40406), .B(n40405), .Z(n40407) );
  OR U53815 ( .A(n40408), .B(n40407), .Z(n40409) );
  AND U53816 ( .A(n40410), .B(n40409), .Z(n40414) );
  NAND U53817 ( .A(n40412), .B(n40411), .Z(n40413) );
  OR U53818 ( .A(n40414), .B(n40413), .Z(n40415) );
  AND U53819 ( .A(n40416), .B(n40415), .Z(n40420) );
  NAND U53820 ( .A(n40418), .B(n40417), .Z(n40419) );
  OR U53821 ( .A(n40420), .B(n40419), .Z(n40421) );
  AND U53822 ( .A(n40422), .B(n40421), .Z(n40423) );
  ANDN U53823 ( .B(n40424), .A(n40423), .Z(n40425) );
  NAND U53824 ( .A(n40426), .B(n40425), .Z(n40427) );
  NANDN U53825 ( .A(n40428), .B(n40427), .Z(n40429) );
  OR U53826 ( .A(n40430), .B(n40429), .Z(n40431) );
  AND U53827 ( .A(n40432), .B(n40431), .Z(n40434) );
  NAND U53828 ( .A(n40434), .B(n40433), .Z(n40435) );
  NANDN U53829 ( .A(n40436), .B(n40435), .Z(n40437) );
  AND U53830 ( .A(n40438), .B(n40437), .Z(n40440) );
  NAND U53831 ( .A(n40440), .B(n40439), .Z(n40441) );
  NANDN U53832 ( .A(n40442), .B(n40441), .Z(n40443) );
  AND U53833 ( .A(n40444), .B(n40443), .Z(n40446) );
  NAND U53834 ( .A(n40446), .B(n40445), .Z(n40447) );
  NANDN U53835 ( .A(n40448), .B(n40447), .Z(n40449) );
  AND U53836 ( .A(n40450), .B(n40449), .Z(n40452) );
  NAND U53837 ( .A(n40452), .B(n40451), .Z(n40453) );
  NAND U53838 ( .A(n40454), .B(n40453), .Z(n40455) );
  AND U53839 ( .A(n40456), .B(n40455), .Z(n40460) );
  NAND U53840 ( .A(n40458), .B(n40457), .Z(n40459) );
  OR U53841 ( .A(n40460), .B(n40459), .Z(n40461) );
  AND U53842 ( .A(n40462), .B(n40461), .Z(n40466) );
  NAND U53843 ( .A(n40464), .B(n40463), .Z(n40465) );
  OR U53844 ( .A(n40466), .B(n40465), .Z(n40467) );
  AND U53845 ( .A(n40468), .B(n40467), .Z(n40470) );
  AND U53846 ( .A(n40470), .B(n40469), .Z(n40474) );
  NAND U53847 ( .A(n40472), .B(n40471), .Z(n40473) );
  OR U53848 ( .A(n40474), .B(n40473), .Z(n40475) );
  AND U53849 ( .A(n40476), .B(n40475), .Z(n40480) );
  AND U53850 ( .A(n40478), .B(n40477), .Z(n40479) );
  NANDN U53851 ( .A(n40480), .B(n40479), .Z(n40481) );
  NAND U53852 ( .A(n40482), .B(n40481), .Z(n40483) );
  NAND U53853 ( .A(n40484), .B(n40483), .Z(n40485) );
  NANDN U53854 ( .A(n40486), .B(n40485), .Z(n40487) );
  AND U53855 ( .A(n40488), .B(n40487), .Z(n40490) );
  NAND U53856 ( .A(n40490), .B(n40489), .Z(n40491) );
  NANDN U53857 ( .A(n40492), .B(n40491), .Z(n40493) );
  AND U53858 ( .A(n40494), .B(n40493), .Z(n40496) );
  NAND U53859 ( .A(n40496), .B(n40495), .Z(n40497) );
  NANDN U53860 ( .A(n40498), .B(n40497), .Z(n40499) );
  AND U53861 ( .A(n40500), .B(n40499), .Z(n40502) );
  AND U53862 ( .A(n40502), .B(n40501), .Z(n40506) );
  NAND U53863 ( .A(n40504), .B(n40503), .Z(n40505) );
  OR U53864 ( .A(n40506), .B(n40505), .Z(n40507) );
  AND U53865 ( .A(n40508), .B(n40507), .Z(n40512) );
  NAND U53866 ( .A(n40510), .B(n40509), .Z(n40511) );
  OR U53867 ( .A(n40512), .B(n40511), .Z(n40513) );
  AND U53868 ( .A(n40514), .B(n40513), .Z(n40515) );
  NOR U53869 ( .A(n40516), .B(n40515), .Z(n40517) );
  NAND U53870 ( .A(n51695), .B(n40517), .Z(n40518) );
  NANDN U53871 ( .A(n40519), .B(n40518), .Z(n40521) );
  AND U53872 ( .A(n40521), .B(n40520), .Z(n40522) );
  NANDN U53873 ( .A(x[4148]), .B(y[4148]), .Z(n51696) );
  NAND U53874 ( .A(n40522), .B(n51696), .Z(n40523) );
  NANDN U53875 ( .A(n40524), .B(n40523), .Z(n40526) );
  IV U53876 ( .A(n40525), .Z(n56380) );
  AND U53877 ( .A(n40526), .B(n56380), .Z(n40528) );
  NAND U53878 ( .A(n40528), .B(n40527), .Z(n40529) );
  NANDN U53879 ( .A(n40530), .B(n40529), .Z(n40531) );
  AND U53880 ( .A(n40532), .B(n40531), .Z(n40536) );
  NAND U53881 ( .A(n40534), .B(n40533), .Z(n40535) );
  OR U53882 ( .A(n40536), .B(n40535), .Z(n40537) );
  AND U53883 ( .A(n40538), .B(n40537), .Z(n40542) );
  NAND U53884 ( .A(n40540), .B(n40539), .Z(n40541) );
  OR U53885 ( .A(n40542), .B(n40541), .Z(n40543) );
  AND U53886 ( .A(n40544), .B(n40543), .Z(n40548) );
  NAND U53887 ( .A(n40546), .B(n40545), .Z(n40547) );
  OR U53888 ( .A(n40548), .B(n40547), .Z(n40549) );
  AND U53889 ( .A(n40550), .B(n40549), .Z(n40554) );
  NAND U53890 ( .A(n40552), .B(n40551), .Z(n40553) );
  OR U53891 ( .A(n40554), .B(n40553), .Z(n40555) );
  AND U53892 ( .A(n40556), .B(n40555), .Z(n40560) );
  NAND U53893 ( .A(n40558), .B(n40557), .Z(n40559) );
  OR U53894 ( .A(n40560), .B(n40559), .Z(n40561) );
  AND U53895 ( .A(n40562), .B(n40561), .Z(n40563) );
  OR U53896 ( .A(n40564), .B(n40563), .Z(n40565) );
  NAND U53897 ( .A(n40566), .B(n40565), .Z(n40567) );
  NAND U53898 ( .A(n40568), .B(n40567), .Z(n40570) );
  ANDN U53899 ( .B(y[4166]), .A(x[4166]), .Z(n40569) );
  ANDN U53900 ( .B(n40570), .A(n40569), .Z(n40572) );
  ANDN U53901 ( .B(n40572), .A(n40571), .Z(n40576) );
  NAND U53902 ( .A(n40574), .B(n40573), .Z(n40575) );
  OR U53903 ( .A(n40576), .B(n40575), .Z(n40577) );
  AND U53904 ( .A(n40578), .B(n40577), .Z(n40582) );
  NAND U53905 ( .A(n40580), .B(n40579), .Z(n40581) );
  OR U53906 ( .A(n40582), .B(n40581), .Z(n40583) );
  AND U53907 ( .A(n40584), .B(n40583), .Z(n40588) );
  NAND U53908 ( .A(n40586), .B(n40585), .Z(n40587) );
  OR U53909 ( .A(n40588), .B(n40587), .Z(n40589) );
  AND U53910 ( .A(n40590), .B(n40589), .Z(n40591) );
  ANDN U53911 ( .B(n40592), .A(n40591), .Z(n40593) );
  NAND U53912 ( .A(n40594), .B(n40593), .Z(n40595) );
  NANDN U53913 ( .A(n40596), .B(n40595), .Z(n40597) );
  OR U53914 ( .A(n40598), .B(n40597), .Z(n40599) );
  AND U53915 ( .A(n40600), .B(n40599), .Z(n40602) );
  NAND U53916 ( .A(n40602), .B(n40601), .Z(n40603) );
  NANDN U53917 ( .A(n40604), .B(n40603), .Z(n40605) );
  AND U53918 ( .A(n40606), .B(n40605), .Z(n40608) );
  NAND U53919 ( .A(n40608), .B(n40607), .Z(n40609) );
  NANDN U53920 ( .A(n40610), .B(n40609), .Z(n40611) );
  AND U53921 ( .A(n40612), .B(n40611), .Z(n40614) );
  AND U53922 ( .A(n40614), .B(n40613), .Z(n40618) );
  NANDN U53923 ( .A(x[4180]), .B(y[4180]), .Z(n40616) );
  NAND U53924 ( .A(n40616), .B(n40615), .Z(n40617) );
  OR U53925 ( .A(n40618), .B(n40617), .Z(n40619) );
  AND U53926 ( .A(n40620), .B(n40619), .Z(n40624) );
  NAND U53927 ( .A(n40622), .B(n40621), .Z(n40623) );
  OR U53928 ( .A(n40624), .B(n40623), .Z(n40625) );
  AND U53929 ( .A(n40626), .B(n40625), .Z(n40630) );
  NAND U53930 ( .A(n40628), .B(n40627), .Z(n40629) );
  OR U53931 ( .A(n40630), .B(n40629), .Z(n40631) );
  AND U53932 ( .A(n40632), .B(n40631), .Z(n40636) );
  NAND U53933 ( .A(n40634), .B(n40633), .Z(n40635) );
  OR U53934 ( .A(n40636), .B(n40635), .Z(n40637) );
  AND U53935 ( .A(n40638), .B(n40637), .Z(n40639) );
  ANDN U53936 ( .B(n40640), .A(n40639), .Z(n40641) );
  NAND U53937 ( .A(n40642), .B(n40641), .Z(n40643) );
  NANDN U53938 ( .A(n40644), .B(n40643), .Z(n40645) );
  OR U53939 ( .A(n40646), .B(n40645), .Z(n40647) );
  AND U53940 ( .A(n40648), .B(n40647), .Z(n40650) );
  NAND U53941 ( .A(n40650), .B(n40649), .Z(n40651) );
  NANDN U53942 ( .A(n40652), .B(n40651), .Z(n40653) );
  AND U53943 ( .A(n40654), .B(n40653), .Z(n40656) );
  NANDN U53944 ( .A(x[4192]), .B(y[4192]), .Z(n40655) );
  AND U53945 ( .A(n40656), .B(n40655), .Z(n40660) );
  AND U53946 ( .A(n40658), .B(n40657), .Z(n40659) );
  NANDN U53947 ( .A(n40660), .B(n40659), .Z(n40662) );
  NAND U53948 ( .A(n40662), .B(n40661), .Z(n40664) );
  ANDN U53949 ( .B(y[4194]), .A(x[4194]), .Z(n40663) );
  OR U53950 ( .A(n40664), .B(n40663), .Z(n40665) );
  NAND U53951 ( .A(n40666), .B(n40665), .Z(n40668) );
  ANDN U53952 ( .B(n40668), .A(n40667), .Z(n40670) );
  NAND U53953 ( .A(n40670), .B(n40669), .Z(n40671) );
  NANDN U53954 ( .A(n40672), .B(n40671), .Z(n40673) );
  AND U53955 ( .A(n40674), .B(n40673), .Z(n40675) );
  NANDN U53956 ( .A(n40676), .B(n40675), .Z(n40677) );
  NAND U53957 ( .A(n40678), .B(n40677), .Z(n40679) );
  NANDN U53958 ( .A(n51680), .B(n40679), .Z(n40680) );
  ANDN U53959 ( .B(n40681), .A(n40680), .Z(n40685) );
  NAND U53960 ( .A(n40683), .B(n40682), .Z(n40684) );
  OR U53961 ( .A(n40685), .B(n40684), .Z(n40686) );
  AND U53962 ( .A(n40687), .B(n40686), .Z(n40691) );
  NAND U53963 ( .A(n40689), .B(n40688), .Z(n40690) );
  OR U53964 ( .A(n40691), .B(n40690), .Z(n40692) );
  AND U53965 ( .A(n40693), .B(n40692), .Z(n40697) );
  NAND U53966 ( .A(n40695), .B(n40694), .Z(n40696) );
  OR U53967 ( .A(n40697), .B(n40696), .Z(n40698) );
  AND U53968 ( .A(n40699), .B(n40698), .Z(n40703) );
  NAND U53969 ( .A(n40701), .B(n40700), .Z(n40702) );
  OR U53970 ( .A(n40703), .B(n40702), .Z(n40704) );
  AND U53971 ( .A(n40705), .B(n40704), .Z(n40709) );
  NAND U53972 ( .A(n40707), .B(n40706), .Z(n40708) );
  OR U53973 ( .A(n40709), .B(n40708), .Z(n40710) );
  AND U53974 ( .A(n40711), .B(n40710), .Z(n40712) );
  OR U53975 ( .A(n40713), .B(n40712), .Z(n40714) );
  NAND U53976 ( .A(n40715), .B(n40714), .Z(n40716) );
  AND U53977 ( .A(n40717), .B(n40716), .Z(n40718) );
  NOR U53978 ( .A(n51678), .B(n40718), .Z(n40719) );
  NANDN U53979 ( .A(n40720), .B(n40719), .Z(n40721) );
  AND U53980 ( .A(n40722), .B(n40721), .Z(n40724) );
  NAND U53981 ( .A(n40724), .B(n40723), .Z(n40725) );
  NANDN U53982 ( .A(n40726), .B(n40725), .Z(n40727) );
  AND U53983 ( .A(n40728), .B(n40727), .Z(n40730) );
  NAND U53984 ( .A(n40730), .B(n40729), .Z(n40731) );
  NANDN U53985 ( .A(n40732), .B(n40731), .Z(n40733) );
  AND U53986 ( .A(n40734), .B(n40733), .Z(n40735) );
  NANDN U53987 ( .A(n40736), .B(n40735), .Z(n40737) );
  AND U53988 ( .A(n40738), .B(n40737), .Z(n40740) );
  NANDN U53989 ( .A(x[4220]), .B(y[4220]), .Z(n40739) );
  NAND U53990 ( .A(n40740), .B(n40739), .Z(n40742) );
  ANDN U53991 ( .B(n40742), .A(n40741), .Z(n40743) );
  NANDN U53992 ( .A(n40744), .B(n40743), .Z(n40745) );
  NAND U53993 ( .A(n40746), .B(n40745), .Z(n40747) );
  NANDN U53994 ( .A(n40748), .B(n40747), .Z(n40749) );
  AND U53995 ( .A(n40750), .B(n40749), .Z(n40752) );
  NAND U53996 ( .A(n40752), .B(n40751), .Z(n40753) );
  NANDN U53997 ( .A(n40754), .B(n40753), .Z(n40755) );
  AND U53998 ( .A(n40756), .B(n40755), .Z(n40758) );
  NAND U53999 ( .A(n40758), .B(n40757), .Z(n40759) );
  NANDN U54000 ( .A(n40760), .B(n40759), .Z(n40761) );
  AND U54001 ( .A(n40762), .B(n40761), .Z(n40764) );
  AND U54002 ( .A(n40764), .B(n40763), .Z(n40768) );
  NAND U54003 ( .A(n40766), .B(n40765), .Z(n40767) );
  OR U54004 ( .A(n40768), .B(n40767), .Z(n40769) );
  AND U54005 ( .A(n40770), .B(n40769), .Z(n40771) );
  OR U54006 ( .A(n40772), .B(n40771), .Z(n40773) );
  NAND U54007 ( .A(n40774), .B(n40773), .Z(n40775) );
  NAND U54008 ( .A(n40776), .B(n40775), .Z(n40777) );
  NANDN U54009 ( .A(n40778), .B(n40777), .Z(n40779) );
  AND U54010 ( .A(n40780), .B(n40779), .Z(n40782) );
  NAND U54011 ( .A(n40782), .B(n40781), .Z(n40783) );
  NANDN U54012 ( .A(n40784), .B(n40783), .Z(n40785) );
  AND U54013 ( .A(n40786), .B(n40785), .Z(n40787) );
  NANDN U54014 ( .A(n40788), .B(n40787), .Z(n40789) );
  NAND U54015 ( .A(n40790), .B(n40789), .Z(n40791) );
  NANDN U54016 ( .A(n40792), .B(n40791), .Z(n40793) );
  AND U54017 ( .A(n40794), .B(n40793), .Z(n40795) );
  NAND U54018 ( .A(n40796), .B(n40795), .Z(n40800) );
  NAND U54019 ( .A(n40798), .B(n40797), .Z(n40799) );
  ANDN U54020 ( .B(n40800), .A(n40799), .Z(n40801) );
  OR U54021 ( .A(n40802), .B(n40801), .Z(n40803) );
  NAND U54022 ( .A(n40804), .B(n40803), .Z(n40805) );
  AND U54023 ( .A(n40806), .B(n40805), .Z(n40807) );
  NOR U54024 ( .A(n40808), .B(n40807), .Z(n40810) );
  NAND U54025 ( .A(n40810), .B(n40809), .Z(n40811) );
  AND U54026 ( .A(n40811), .B(n51674), .Z(n40813) );
  NANDN U54027 ( .A(x[4246]), .B(y[4246]), .Z(n40812) );
  AND U54028 ( .A(n40813), .B(n40812), .Z(n40814) );
  NOR U54029 ( .A(n40815), .B(n40814), .Z(n40817) );
  NAND U54030 ( .A(n40817), .B(n40816), .Z(n40819) );
  AND U54031 ( .A(n40819), .B(n40818), .Z(n40820) );
  NANDN U54032 ( .A(x[4248]), .B(y[4248]), .Z(n51675) );
  AND U54033 ( .A(n40820), .B(n51675), .Z(n40821) );
  OR U54034 ( .A(n40822), .B(n40821), .Z(n40823) );
  NAND U54035 ( .A(n40824), .B(n40823), .Z(n40828) );
  NAND U54036 ( .A(n40826), .B(n40825), .Z(n40827) );
  ANDN U54037 ( .B(n40828), .A(n40827), .Z(n40832) );
  NAND U54038 ( .A(n40830), .B(n40829), .Z(n40831) );
  OR U54039 ( .A(n40832), .B(n40831), .Z(n40833) );
  AND U54040 ( .A(n40834), .B(n40833), .Z(n40838) );
  NAND U54041 ( .A(n40836), .B(n40835), .Z(n40837) );
  OR U54042 ( .A(n40838), .B(n40837), .Z(n40839) );
  AND U54043 ( .A(n40840), .B(n40839), .Z(n40841) );
  ANDN U54044 ( .B(n56502), .A(n40841), .Z(n40842) );
  NAND U54045 ( .A(n40843), .B(n40842), .Z(n40844) );
  NANDN U54046 ( .A(n40845), .B(n40844), .Z(n40847) );
  OR U54047 ( .A(n40847), .B(n40846), .Z(n40848) );
  AND U54048 ( .A(n40849), .B(n40848), .Z(n40850) );
  NANDN U54049 ( .A(x[4258]), .B(y[4258]), .Z(n56503) );
  AND U54050 ( .A(n40850), .B(n56503), .Z(n40854) );
  NAND U54051 ( .A(n40852), .B(n40851), .Z(n40853) );
  OR U54052 ( .A(n40854), .B(n40853), .Z(n40855) );
  AND U54053 ( .A(n40856), .B(n40855), .Z(n40857) );
  NANDN U54054 ( .A(n40858), .B(n40857), .Z(n40859) );
  AND U54055 ( .A(n40860), .B(n40859), .Z(n40861) );
  OR U54056 ( .A(n40862), .B(n40861), .Z(n40863) );
  NAND U54057 ( .A(n40864), .B(n40863), .Z(n40865) );
  NANDN U54058 ( .A(n40866), .B(n40865), .Z(n40868) );
  ANDN U54059 ( .B(y[4264]), .A(x[4264]), .Z(n40867) );
  OR U54060 ( .A(n40868), .B(n40867), .Z(n40869) );
  NANDN U54061 ( .A(n40870), .B(n40869), .Z(n40871) );
  AND U54062 ( .A(n40872), .B(n40871), .Z(n40874) );
  NANDN U54063 ( .A(x[4266]), .B(y[4266]), .Z(n40873) );
  NAND U54064 ( .A(n40874), .B(n40873), .Z(n40875) );
  AND U54065 ( .A(n40876), .B(n40875), .Z(n40877) );
  OR U54066 ( .A(n40878), .B(n40877), .Z(n40879) );
  NAND U54067 ( .A(n40880), .B(n40879), .Z(n40881) );
  NANDN U54068 ( .A(n40882), .B(n40881), .Z(n40883) );
  NAND U54069 ( .A(n40884), .B(n40883), .Z(n40885) );
  NANDN U54070 ( .A(n40886), .B(n40885), .Z(n40887) );
  AND U54071 ( .A(n40888), .B(n40887), .Z(n40890) );
  NAND U54072 ( .A(n40890), .B(n40889), .Z(n40891) );
  NANDN U54073 ( .A(n40892), .B(n40891), .Z(n40893) );
  AND U54074 ( .A(n40894), .B(n40893), .Z(n40896) );
  NAND U54075 ( .A(n40896), .B(n40895), .Z(n40897) );
  NANDN U54076 ( .A(n40898), .B(n40897), .Z(n40899) );
  AND U54077 ( .A(n40900), .B(n40899), .Z(n40902) );
  NAND U54078 ( .A(n40902), .B(n40901), .Z(n40903) );
  AND U54079 ( .A(n40904), .B(n40903), .Z(n40905) );
  NOR U54080 ( .A(n40906), .B(n40905), .Z(n40908) );
  NAND U54081 ( .A(n40908), .B(n40907), .Z(n40912) );
  NANDN U54082 ( .A(x[4280]), .B(y[4280]), .Z(n40909) );
  AND U54083 ( .A(n40910), .B(n40909), .Z(n40911) );
  NAND U54084 ( .A(n40912), .B(n40911), .Z(n40913) );
  NANDN U54085 ( .A(n40914), .B(n40913), .Z(n40915) );
  NAND U54086 ( .A(n40916), .B(n40915), .Z(n40917) );
  NANDN U54087 ( .A(n40918), .B(n40917), .Z(n40919) );
  AND U54088 ( .A(n40920), .B(n40919), .Z(n40922) );
  NAND U54089 ( .A(n40922), .B(n40921), .Z(n40923) );
  NANDN U54090 ( .A(n40924), .B(n40923), .Z(n40925) );
  AND U54091 ( .A(n40926), .B(n40925), .Z(n40927) );
  NANDN U54092 ( .A(n40928), .B(n40927), .Z(n40929) );
  NAND U54093 ( .A(n40930), .B(n40929), .Z(n40931) );
  NANDN U54094 ( .A(n40932), .B(n40931), .Z(n40934) );
  OR U54095 ( .A(n40934), .B(n40933), .Z(n40935) );
  NAND U54096 ( .A(n40936), .B(n40935), .Z(n40940) );
  NAND U54097 ( .A(n40938), .B(n40937), .Z(n40939) );
  ANDN U54098 ( .B(n40940), .A(n40939), .Z(n40944) );
  NAND U54099 ( .A(n40942), .B(n40941), .Z(n40943) );
  OR U54100 ( .A(n40944), .B(n40943), .Z(n40945) );
  AND U54101 ( .A(n40946), .B(n40945), .Z(n40950) );
  AND U54102 ( .A(n40948), .B(n40947), .Z(n40949) );
  NANDN U54103 ( .A(n40950), .B(n40949), .Z(n40951) );
  NAND U54104 ( .A(n40952), .B(n40951), .Z(n40953) );
  NAND U54105 ( .A(n40954), .B(n40953), .Z(n40955) );
  NAND U54106 ( .A(n40956), .B(n40955), .Z(n40957) );
  NANDN U54107 ( .A(n40958), .B(n40957), .Z(n40960) );
  OR U54108 ( .A(n40960), .B(n40959), .Z(n40961) );
  NAND U54109 ( .A(n40962), .B(n40961), .Z(n40963) );
  NANDN U54110 ( .A(n40964), .B(n40963), .Z(n40966) );
  OR U54111 ( .A(n40966), .B(n40965), .Z(n40967) );
  NAND U54112 ( .A(n40968), .B(n40967), .Z(n40969) );
  NANDN U54113 ( .A(n40970), .B(n40969), .Z(n40971) );
  AND U54114 ( .A(n40971), .B(n51661), .Z(n40972) );
  NANDN U54115 ( .A(x[4302]), .B(y[4302]), .Z(n56546) );
  AND U54116 ( .A(n40972), .B(n56546), .Z(n40973) );
  NOR U54117 ( .A(n40974), .B(n40973), .Z(n40976) );
  NAND U54118 ( .A(n40976), .B(n40975), .Z(n40978) );
  AND U54119 ( .A(n40978), .B(n40977), .Z(n40979) );
  NANDN U54120 ( .A(x[4304]), .B(y[4304]), .Z(n51662) );
  AND U54121 ( .A(n40979), .B(n51662), .Z(n40980) );
  OR U54122 ( .A(n40981), .B(n40980), .Z(n40982) );
  NAND U54123 ( .A(n40983), .B(n40982), .Z(n40987) );
  NAND U54124 ( .A(n40985), .B(n40984), .Z(n40986) );
  ANDN U54125 ( .B(n40987), .A(n40986), .Z(n40991) );
  NAND U54126 ( .A(n40989), .B(n40988), .Z(n40990) );
  OR U54127 ( .A(n40991), .B(n40990), .Z(n40992) );
  AND U54128 ( .A(n40993), .B(n40992), .Z(n40997) );
  NAND U54129 ( .A(n40995), .B(n40994), .Z(n40996) );
  OR U54130 ( .A(n40997), .B(n40996), .Z(n40998) );
  AND U54131 ( .A(n40999), .B(n40998), .Z(n41003) );
  NAND U54132 ( .A(n41001), .B(n41000), .Z(n41002) );
  OR U54133 ( .A(n41003), .B(n41002), .Z(n41004) );
  AND U54134 ( .A(n41005), .B(n41004), .Z(n41009) );
  NAND U54135 ( .A(n41007), .B(n41006), .Z(n41008) );
  OR U54136 ( .A(n41009), .B(n41008), .Z(n41010) );
  AND U54137 ( .A(n41011), .B(n41010), .Z(n41012) );
  NOR U54138 ( .A(n41013), .B(n41012), .Z(n41014) );
  NAND U54139 ( .A(n41015), .B(n41014), .Z(n41019) );
  NAND U54140 ( .A(n41017), .B(n41016), .Z(n41018) );
  ANDN U54141 ( .B(n41019), .A(n41018), .Z(n41023) );
  NANDN U54142 ( .A(x[4318]), .B(y[4318]), .Z(n41021) );
  NAND U54143 ( .A(n41021), .B(n41020), .Z(n41022) );
  OR U54144 ( .A(n41023), .B(n41022), .Z(n41024) );
  AND U54145 ( .A(n41025), .B(n41024), .Z(n41028) );
  NAND U54146 ( .A(n41026), .B(n56564), .Z(n41027) );
  OR U54147 ( .A(n41028), .B(n41027), .Z(n41029) );
  AND U54148 ( .A(n41030), .B(n41029), .Z(n41032) );
  NAND U54149 ( .A(n41032), .B(n41031), .Z(n41034) );
  AND U54150 ( .A(n41034), .B(n41033), .Z(n41035) );
  NANDN U54151 ( .A(x[4322]), .B(y[4322]), .Z(n56565) );
  AND U54152 ( .A(n41035), .B(n56565), .Z(n41039) );
  AND U54153 ( .A(n41037), .B(n41036), .Z(n41038) );
  NANDN U54154 ( .A(n41039), .B(n41038), .Z(n41041) );
  AND U54155 ( .A(n41041), .B(n41040), .Z(n41043) );
  NANDN U54156 ( .A(x[4324]), .B(y[4324]), .Z(n41042) );
  AND U54157 ( .A(n41043), .B(n41042), .Z(n41044) );
  NOR U54158 ( .A(n41045), .B(n41044), .Z(n41047) );
  NAND U54159 ( .A(n41047), .B(n41046), .Z(n41051) );
  NANDN U54160 ( .A(x[4326]), .B(y[4326]), .Z(n41048) );
  AND U54161 ( .A(n41049), .B(n41048), .Z(n41050) );
  NAND U54162 ( .A(n41051), .B(n41050), .Z(n41052) );
  NANDN U54163 ( .A(n41053), .B(n41052), .Z(n41054) );
  NAND U54164 ( .A(n41055), .B(n41054), .Z(n41056) );
  NANDN U54165 ( .A(n41057), .B(n41056), .Z(n41058) );
  AND U54166 ( .A(n41059), .B(n41058), .Z(n41061) );
  NAND U54167 ( .A(n41061), .B(n41060), .Z(n41062) );
  NANDN U54168 ( .A(n41063), .B(n41062), .Z(n41064) );
  AND U54169 ( .A(n41065), .B(n41064), .Z(n41067) );
  NAND U54170 ( .A(n41067), .B(n41066), .Z(n41068) );
  NANDN U54171 ( .A(n41069), .B(n41068), .Z(n41070) );
  AND U54172 ( .A(n41070), .B(n51657), .Z(n41072) );
  AND U54173 ( .A(n41072), .B(n41071), .Z(n41076) );
  NAND U54174 ( .A(n41074), .B(n41073), .Z(n41075) );
  OR U54175 ( .A(n41076), .B(n41075), .Z(n41077) );
  AND U54176 ( .A(n41078), .B(n41077), .Z(n41082) );
  NAND U54177 ( .A(n41080), .B(n41079), .Z(n41081) );
  OR U54178 ( .A(n41082), .B(n41081), .Z(n41083) );
  AND U54179 ( .A(n41084), .B(n41083), .Z(n41088) );
  NAND U54180 ( .A(n41086), .B(n41085), .Z(n41087) );
  OR U54181 ( .A(n41088), .B(n41087), .Z(n41089) );
  AND U54182 ( .A(n41090), .B(n41089), .Z(n41094) );
  NAND U54183 ( .A(n41092), .B(n41091), .Z(n41093) );
  OR U54184 ( .A(n41094), .B(n41093), .Z(n41095) );
  AND U54185 ( .A(n41096), .B(n41095), .Z(n41100) );
  NAND U54186 ( .A(n41098), .B(n41097), .Z(n41099) );
  OR U54187 ( .A(n41100), .B(n41099), .Z(n41101) );
  AND U54188 ( .A(n41102), .B(n41101), .Z(n41106) );
  NAND U54189 ( .A(n41104), .B(n41103), .Z(n41105) );
  OR U54190 ( .A(n41106), .B(n41105), .Z(n41107) );
  AND U54191 ( .A(n41108), .B(n41107), .Z(n41112) );
  NAND U54192 ( .A(n41110), .B(n41109), .Z(n41111) );
  OR U54193 ( .A(n41112), .B(n41111), .Z(n41113) );
  AND U54194 ( .A(n41114), .B(n41113), .Z(n41115) );
  OR U54195 ( .A(n41116), .B(n41115), .Z(n41117) );
  NAND U54196 ( .A(n41118), .B(n41117), .Z(n41119) );
  NANDN U54197 ( .A(n41120), .B(n41119), .Z(n41121) );
  AND U54198 ( .A(n41121), .B(n56594), .Z(n41122) );
  OR U54199 ( .A(n41122), .B(n56596), .Z(n41123) );
  NAND U54200 ( .A(n41124), .B(n41123), .Z(n41125) );
  NANDN U54201 ( .A(n41126), .B(n41125), .Z(n41127) );
  AND U54202 ( .A(n41128), .B(n41127), .Z(n41132) );
  NAND U54203 ( .A(n41130), .B(n41129), .Z(n41131) );
  OR U54204 ( .A(n41132), .B(n41131), .Z(n41133) );
  AND U54205 ( .A(n41134), .B(n41133), .Z(n41136) );
  NAND U54206 ( .A(n41136), .B(n41135), .Z(n41137) );
  NANDN U54207 ( .A(n41138), .B(n41137), .Z(n41139) );
  AND U54208 ( .A(n41139), .B(n56600), .Z(n41141) );
  NANDN U54209 ( .A(x[4358]), .B(y[4358]), .Z(n41140) );
  AND U54210 ( .A(n41141), .B(n41140), .Z(n41142) );
  OR U54211 ( .A(n41143), .B(n41142), .Z(n41144) );
  AND U54212 ( .A(n41145), .B(n41144), .Z(n41149) );
  NAND U54213 ( .A(n41147), .B(n41146), .Z(n41148) );
  OR U54214 ( .A(n41149), .B(n41148), .Z(n41150) );
  AND U54215 ( .A(n41151), .B(n41150), .Z(n41152) );
  OR U54216 ( .A(n41153), .B(n41152), .Z(n41154) );
  NAND U54217 ( .A(n41155), .B(n41154), .Z(n41156) );
  AND U54218 ( .A(n41157), .B(n41156), .Z(n41158) );
  NOR U54219 ( .A(n51646), .B(n41158), .Z(n41159) );
  NAND U54220 ( .A(n41160), .B(n41159), .Z(n41161) );
  NANDN U54221 ( .A(n41162), .B(n41161), .Z(n41164) );
  OR U54222 ( .A(n41164), .B(n41163), .Z(n41165) );
  NAND U54223 ( .A(n41166), .B(n41165), .Z(n41167) );
  NANDN U54224 ( .A(n41168), .B(n41167), .Z(n41170) );
  OR U54225 ( .A(n41170), .B(n41169), .Z(n41171) );
  NAND U54226 ( .A(n41172), .B(n41171), .Z(n41173) );
  NANDN U54227 ( .A(n41174), .B(n41173), .Z(n41175) );
  AND U54228 ( .A(n41176), .B(n41175), .Z(n41177) );
  NOR U54229 ( .A(n41178), .B(n41177), .Z(n41180) );
  NAND U54230 ( .A(n41180), .B(n41179), .Z(n41183) );
  NANDN U54231 ( .A(x[4374]), .B(y[4374]), .Z(n51644) );
  AND U54232 ( .A(n41181), .B(n51644), .Z(n41182) );
  NAND U54233 ( .A(n41183), .B(n41182), .Z(n41184) );
  NANDN U54234 ( .A(n41185), .B(n41184), .Z(n41186) );
  NAND U54235 ( .A(n41187), .B(n41186), .Z(n41188) );
  NANDN U54236 ( .A(n41189), .B(n41188), .Z(n41190) );
  AND U54237 ( .A(n41191), .B(n41190), .Z(n41193) );
  NAND U54238 ( .A(n41193), .B(n41192), .Z(n41194) );
  NANDN U54239 ( .A(n41195), .B(n41194), .Z(n41196) );
  AND U54240 ( .A(n41197), .B(n41196), .Z(n41198) );
  NANDN U54241 ( .A(n41199), .B(n41198), .Z(n41200) );
  AND U54242 ( .A(n41201), .B(n41200), .Z(n41202) );
  NAND U54243 ( .A(n41203), .B(n41202), .Z(n41205) );
  ANDN U54244 ( .B(n41205), .A(n41204), .Z(n41206) );
  NANDN U54245 ( .A(n41207), .B(n41206), .Z(n41208) );
  AND U54246 ( .A(n41209), .B(n41208), .Z(n41210) );
  NOR U54247 ( .A(n41211), .B(n41210), .Z(n41212) );
  NANDN U54248 ( .A(n41213), .B(n41212), .Z(n41214) );
  AND U54249 ( .A(n41215), .B(n41214), .Z(n41217) );
  NAND U54250 ( .A(n41217), .B(n41216), .Z(n41218) );
  NANDN U54251 ( .A(n41219), .B(n41218), .Z(n41220) );
  AND U54252 ( .A(n41221), .B(n41220), .Z(n41223) );
  NAND U54253 ( .A(n41223), .B(n41222), .Z(n41224) );
  NANDN U54254 ( .A(n41225), .B(n41224), .Z(n41226) );
  AND U54255 ( .A(n41227), .B(n41226), .Z(n41228) );
  NAND U54256 ( .A(n41228), .B(y[4390]), .Z(n41231) );
  XOR U54257 ( .A(n41228), .B(y[4390]), .Z(n41229) );
  NANDN U54258 ( .A(x[4390]), .B(n41229), .Z(n41230) );
  NAND U54259 ( .A(n41231), .B(n41230), .Z(n41232) );
  OR U54260 ( .A(n41233), .B(n41232), .Z(n41234) );
  AND U54261 ( .A(n41235), .B(n41234), .Z(n41238) );
  AND U54262 ( .A(n41236), .B(n56633), .Z(n41237) );
  NANDN U54263 ( .A(n41238), .B(n41237), .Z(n41239) );
  NANDN U54264 ( .A(n41240), .B(n41239), .Z(n41241) );
  AND U54265 ( .A(n41242), .B(n41241), .Z(n41243) );
  NANDN U54266 ( .A(x[4394]), .B(y[4394]), .Z(n56634) );
  NAND U54267 ( .A(n41243), .B(n56634), .Z(n41244) );
  AND U54268 ( .A(n41245), .B(n41244), .Z(n41247) );
  NANDN U54269 ( .A(n41247), .B(n41246), .Z(n41249) );
  ANDN U54270 ( .B(y[4396]), .A(x[4396]), .Z(n41248) );
  OR U54271 ( .A(n41249), .B(n41248), .Z(n41250) );
  NAND U54272 ( .A(n41251), .B(n41250), .Z(n41252) );
  NANDN U54273 ( .A(n41253), .B(n41252), .Z(n41254) );
  OR U54274 ( .A(n41255), .B(n41254), .Z(n41256) );
  AND U54275 ( .A(n41257), .B(n41256), .Z(n41258) );
  NANDN U54276 ( .A(n41259), .B(n41258), .Z(n41260) );
  AND U54277 ( .A(n41261), .B(n41260), .Z(n41265) );
  NAND U54278 ( .A(n41263), .B(n41262), .Z(n41264) );
  OR U54279 ( .A(n41265), .B(n41264), .Z(n41266) );
  AND U54280 ( .A(n41267), .B(n41266), .Z(n41268) );
  OR U54281 ( .A(n41269), .B(n41268), .Z(n41270) );
  NAND U54282 ( .A(n41271), .B(n41270), .Z(n41272) );
  AND U54283 ( .A(n41273), .B(n41272), .Z(n41274) );
  NOR U54284 ( .A(n56647), .B(n41274), .Z(n41275) );
  NANDN U54285 ( .A(n51634), .B(n41275), .Z(n41276) );
  AND U54286 ( .A(n41277), .B(n41276), .Z(n41279) );
  NAND U54287 ( .A(n41279), .B(n41278), .Z(n41280) );
  NANDN U54288 ( .A(n41281), .B(n41280), .Z(n41282) );
  AND U54289 ( .A(n41283), .B(n41282), .Z(n41285) );
  NAND U54290 ( .A(n41285), .B(n41284), .Z(n41286) );
  NANDN U54291 ( .A(n41287), .B(n41286), .Z(n41288) );
  AND U54292 ( .A(n41289), .B(n41288), .Z(n41291) );
  NAND U54293 ( .A(n41291), .B(n41290), .Z(n41292) );
  AND U54294 ( .A(n41292), .B(n56655), .Z(n41293) );
  ANDN U54295 ( .B(y[4412]), .A(x[4412]), .Z(n56653) );
  ANDN U54296 ( .B(n41293), .A(n56653), .Z(n41297) );
  AND U54297 ( .A(n41295), .B(n41294), .Z(n41296) );
  NANDN U54298 ( .A(n41297), .B(n41296), .Z(n41300) );
  NANDN U54299 ( .A(x[4414]), .B(y[4414]), .Z(n56656) );
  AND U54300 ( .A(n41298), .B(n56656), .Z(n41299) );
  NAND U54301 ( .A(n41300), .B(n41299), .Z(n41301) );
  NANDN U54302 ( .A(n41302), .B(n41301), .Z(n41303) );
  NAND U54303 ( .A(n41304), .B(n41303), .Z(n41305) );
  NANDN U54304 ( .A(n41306), .B(n41305), .Z(n41307) );
  AND U54305 ( .A(n41308), .B(n41307), .Z(n41310) );
  NAND U54306 ( .A(n41310), .B(n41309), .Z(n41311) );
  NANDN U54307 ( .A(n41312), .B(n41311), .Z(n41313) );
  AND U54308 ( .A(n41314), .B(n41313), .Z(n41316) );
  NAND U54309 ( .A(n41316), .B(n41315), .Z(n41317) );
  NANDN U54310 ( .A(n41318), .B(n41317), .Z(n41319) );
  AND U54311 ( .A(n41320), .B(n41319), .Z(n41322) );
  NANDN U54312 ( .A(x[4422]), .B(y[4422]), .Z(n41321) );
  AND U54313 ( .A(n41322), .B(n41321), .Z(n41323) );
  OR U54314 ( .A(n41324), .B(n41323), .Z(n41325) );
  AND U54315 ( .A(n41326), .B(n41325), .Z(n41327) );
  OR U54316 ( .A(n41328), .B(n41327), .Z(n41329) );
  NAND U54317 ( .A(n41330), .B(n41329), .Z(n41331) );
  AND U54318 ( .A(n41332), .B(n41331), .Z(n41333) );
  NOR U54319 ( .A(n56666), .B(n41333), .Z(n41334) );
  NANDN U54320 ( .A(n56668), .B(n41334), .Z(n41335) );
  AND U54321 ( .A(n41336), .B(n41335), .Z(n41338) );
  NAND U54322 ( .A(n41338), .B(n41337), .Z(n41339) );
  NANDN U54323 ( .A(n41340), .B(n41339), .Z(n41341) );
  AND U54324 ( .A(n41342), .B(n41341), .Z(n41344) );
  NAND U54325 ( .A(n41344), .B(n41343), .Z(n41345) );
  NANDN U54326 ( .A(n41346), .B(n41345), .Z(n41347) );
  AND U54327 ( .A(n41348), .B(n41347), .Z(n41350) );
  NAND U54328 ( .A(n41350), .B(n41349), .Z(n41352) );
  AND U54329 ( .A(n41352), .B(n41351), .Z(n41354) );
  NANDN U54330 ( .A(x[4434]), .B(y[4434]), .Z(n41353) );
  AND U54331 ( .A(n41354), .B(n41353), .Z(n41355) );
  NOR U54332 ( .A(n41356), .B(n41355), .Z(n41358) );
  NAND U54333 ( .A(n41358), .B(n41357), .Z(n41360) );
  AND U54334 ( .A(n41360), .B(n41359), .Z(n41362) );
  NANDN U54335 ( .A(x[4436]), .B(y[4436]), .Z(n41361) );
  AND U54336 ( .A(n41362), .B(n41361), .Z(n41363) );
  NOR U54337 ( .A(n41364), .B(n41363), .Z(n41366) );
  NAND U54338 ( .A(n41366), .B(n41365), .Z(n41368) );
  AND U54339 ( .A(n41368), .B(n41367), .Z(n41370) );
  NANDN U54340 ( .A(x[4438]), .B(y[4438]), .Z(n41369) );
  AND U54341 ( .A(n41370), .B(n41369), .Z(n41371) );
  NOR U54342 ( .A(n41372), .B(n41371), .Z(n41374) );
  NAND U54343 ( .A(n41374), .B(n41373), .Z(n41376) );
  AND U54344 ( .A(n41376), .B(n41375), .Z(n41378) );
  NANDN U54345 ( .A(x[4440]), .B(y[4440]), .Z(n41377) );
  AND U54346 ( .A(n41378), .B(n41377), .Z(n41382) );
  AND U54347 ( .A(n41380), .B(n41379), .Z(n41381) );
  NANDN U54348 ( .A(n41382), .B(n41381), .Z(n41384) );
  AND U54349 ( .A(n41384), .B(n41383), .Z(n41386) );
  NANDN U54350 ( .A(x[4442]), .B(y[4442]), .Z(n41385) );
  AND U54351 ( .A(n41386), .B(n41385), .Z(n41387) );
  NOR U54352 ( .A(n41388), .B(n41387), .Z(n41390) );
  NAND U54353 ( .A(n41390), .B(n41389), .Z(n41392) );
  AND U54354 ( .A(n41392), .B(n41391), .Z(n41393) );
  NANDN U54355 ( .A(n41394), .B(n41393), .Z(n41395) );
  NAND U54356 ( .A(n41396), .B(n41395), .Z(n41398) );
  AND U54357 ( .A(n41398), .B(n41397), .Z(n41400) );
  NANDN U54358 ( .A(x[4446]), .B(y[4446]), .Z(n41399) );
  AND U54359 ( .A(n41400), .B(n41399), .Z(n41401) );
  NOR U54360 ( .A(n41402), .B(n41401), .Z(n41404) );
  NAND U54361 ( .A(n41404), .B(n41403), .Z(n41405) );
  AND U54362 ( .A(n41405), .B(n56688), .Z(n41406) );
  NANDN U54363 ( .A(n41407), .B(n41406), .Z(n41408) );
  NAND U54364 ( .A(n41409), .B(n41408), .Z(n41411) );
  AND U54365 ( .A(n41411), .B(n41410), .Z(n41412) );
  NANDN U54366 ( .A(x[4450]), .B(y[4450]), .Z(n56689) );
  AND U54367 ( .A(n41412), .B(n56689), .Z(n41416) );
  AND U54368 ( .A(n41414), .B(n41413), .Z(n41415) );
  NANDN U54369 ( .A(n41416), .B(n41415), .Z(n41420) );
  NANDN U54370 ( .A(x[4452]), .B(y[4452]), .Z(n41417) );
  AND U54371 ( .A(n41418), .B(n41417), .Z(n41419) );
  NAND U54372 ( .A(n41420), .B(n41419), .Z(n41421) );
  NANDN U54373 ( .A(n41422), .B(n41421), .Z(n41423) );
  AND U54374 ( .A(n41424), .B(n41423), .Z(n41428) );
  AND U54375 ( .A(n41426), .B(n41425), .Z(n41427) );
  NANDN U54376 ( .A(n41428), .B(n41427), .Z(n41430) );
  AND U54377 ( .A(n41430), .B(n41429), .Z(n41431) );
  NANDN U54378 ( .A(n41432), .B(n41431), .Z(n41433) );
  AND U54379 ( .A(n41434), .B(n41433), .Z(n41435) );
  OR U54380 ( .A(n41436), .B(n41435), .Z(n41437) );
  NAND U54381 ( .A(n41438), .B(n41437), .Z(n41439) );
  NANDN U54382 ( .A(n41440), .B(n41439), .Z(n41444) );
  AND U54383 ( .A(n41442), .B(n41441), .Z(n41443) );
  NAND U54384 ( .A(n41444), .B(n41443), .Z(n41445) );
  NANDN U54385 ( .A(n41446), .B(n41445), .Z(n41447) );
  ANDN U54386 ( .B(y[4462]), .A(x[4462]), .Z(n56700) );
  OR U54387 ( .A(n41447), .B(n56700), .Z(n41448) );
  NAND U54388 ( .A(n41449), .B(n41448), .Z(n41450) );
  NANDN U54389 ( .A(n41451), .B(n41450), .Z(n41453) );
  OR U54390 ( .A(n41453), .B(n41452), .Z(n41454) );
  NANDN U54391 ( .A(n41455), .B(n41454), .Z(n41456) );
  AND U54392 ( .A(n41457), .B(n41456), .Z(n41461) );
  NAND U54393 ( .A(n41459), .B(n41458), .Z(n41460) );
  OR U54394 ( .A(n41461), .B(n41460), .Z(n41462) );
  AND U54395 ( .A(n41463), .B(n41462), .Z(n41467) );
  NAND U54396 ( .A(n41465), .B(n41464), .Z(n41466) );
  OR U54397 ( .A(n41467), .B(n41466), .Z(n41468) );
  AND U54398 ( .A(n41469), .B(n41468), .Z(n41470) );
  ANDN U54399 ( .B(n41471), .A(n41470), .Z(n41472) );
  NAND U54400 ( .A(n41473), .B(n41472), .Z(n41474) );
  NANDN U54401 ( .A(n41475), .B(n41474), .Z(n41476) );
  OR U54402 ( .A(n41477), .B(n41476), .Z(n41478) );
  AND U54403 ( .A(n41479), .B(n41478), .Z(n41481) );
  NAND U54404 ( .A(n41481), .B(n41480), .Z(n41482) );
  NANDN U54405 ( .A(n41483), .B(n41482), .Z(n41484) );
  AND U54406 ( .A(n41485), .B(n41484), .Z(n41487) );
  NAND U54407 ( .A(n41487), .B(n41486), .Z(n41488) );
  NANDN U54408 ( .A(n41489), .B(n41488), .Z(n41490) );
  AND U54409 ( .A(n41491), .B(n41490), .Z(n41493) );
  NAND U54410 ( .A(n41493), .B(n41492), .Z(n41496) );
  NANDN U54411 ( .A(x[4478]), .B(y[4478]), .Z(n51613) );
  AND U54412 ( .A(n41494), .B(n51613), .Z(n41495) );
  NAND U54413 ( .A(n41496), .B(n41495), .Z(n41497) );
  NANDN U54414 ( .A(n41498), .B(n41497), .Z(n41499) );
  NAND U54415 ( .A(n41500), .B(n41499), .Z(n41501) );
  NAND U54416 ( .A(n41502), .B(n41501), .Z(n41503) );
  NANDN U54417 ( .A(n41504), .B(n41503), .Z(n41506) );
  ANDN U54418 ( .B(y[4482]), .A(x[4482]), .Z(n41505) );
  OR U54419 ( .A(n41506), .B(n41505), .Z(n41507) );
  NAND U54420 ( .A(n41508), .B(n41507), .Z(n41509) );
  NAND U54421 ( .A(n56723), .B(n41509), .Z(n41511) );
  ANDN U54422 ( .B(y[4484]), .A(x[4484]), .Z(n41510) );
  OR U54423 ( .A(n41511), .B(n41510), .Z(n41512) );
  NAND U54424 ( .A(n41513), .B(n41512), .Z(n41514) );
  NANDN U54425 ( .A(n41515), .B(n41514), .Z(n41516) );
  ANDN U54426 ( .B(n56722), .A(n41516), .Z(n41517) );
  OR U54427 ( .A(n41518), .B(n41517), .Z(n41519) );
  NAND U54428 ( .A(n41520), .B(n41519), .Z(n41521) );
  NAND U54429 ( .A(n56729), .B(n41521), .Z(n41522) );
  NANDN U54430 ( .A(n56730), .B(n41522), .Z(n41523) );
  AND U54431 ( .A(n41524), .B(n41523), .Z(n41525) );
  OR U54432 ( .A(n41526), .B(n41525), .Z(n41527) );
  NAND U54433 ( .A(n41528), .B(n41527), .Z(n41529) );
  AND U54434 ( .A(n41530), .B(n41529), .Z(n41531) );
  NOR U54435 ( .A(n41532), .B(n41531), .Z(n41534) );
  NAND U54436 ( .A(n41534), .B(n41533), .Z(n41536) );
  AND U54437 ( .A(n41536), .B(n41535), .Z(n41538) );
  NANDN U54438 ( .A(x[4496]), .B(y[4496]), .Z(n41537) );
  AND U54439 ( .A(n41538), .B(n41537), .Z(n41542) );
  AND U54440 ( .A(n41540), .B(n41539), .Z(n41541) );
  NANDN U54441 ( .A(n41542), .B(n41541), .Z(n41544) );
  AND U54442 ( .A(n41544), .B(n41543), .Z(n41546) );
  NANDN U54443 ( .A(x[4498]), .B(y[4498]), .Z(n41545) );
  AND U54444 ( .A(n41546), .B(n41545), .Z(n41547) );
  NOR U54445 ( .A(n41548), .B(n41547), .Z(n41550) );
  NAND U54446 ( .A(n41550), .B(n41549), .Z(n41552) );
  AND U54447 ( .A(n41552), .B(n41551), .Z(n41554) );
  NANDN U54448 ( .A(x[4500]), .B(y[4500]), .Z(n41553) );
  AND U54449 ( .A(n41554), .B(n41553), .Z(n41555) );
  NOR U54450 ( .A(n41556), .B(n41555), .Z(n41558) );
  NAND U54451 ( .A(n41558), .B(n41557), .Z(n41562) );
  NANDN U54452 ( .A(x[4502]), .B(y[4502]), .Z(n41559) );
  AND U54453 ( .A(n41560), .B(n41559), .Z(n41561) );
  NAND U54454 ( .A(n41562), .B(n41561), .Z(n41563) );
  NANDN U54455 ( .A(n41564), .B(n41563), .Z(n41565) );
  NAND U54456 ( .A(n41566), .B(n41565), .Z(n41567) );
  NANDN U54457 ( .A(n41568), .B(n41567), .Z(n41569) );
  AND U54458 ( .A(n41570), .B(n41569), .Z(n41572) );
  NAND U54459 ( .A(n41572), .B(n41571), .Z(n41573) );
  NANDN U54460 ( .A(n41574), .B(n41573), .Z(n41575) );
  AND U54461 ( .A(n41576), .B(n41575), .Z(n41578) );
  NAND U54462 ( .A(n41578), .B(n41577), .Z(n41579) );
  NANDN U54463 ( .A(n41580), .B(n41579), .Z(n41581) );
  AND U54464 ( .A(n41582), .B(n41581), .Z(n41584) );
  NANDN U54465 ( .A(x[4510]), .B(y[4510]), .Z(n41583) );
  AND U54466 ( .A(n41584), .B(n41583), .Z(n41588) );
  NAND U54467 ( .A(n41586), .B(n41585), .Z(n41587) );
  OR U54468 ( .A(n41588), .B(n41587), .Z(n41589) );
  AND U54469 ( .A(n41590), .B(n41589), .Z(n41594) );
  NAND U54470 ( .A(n41592), .B(n41591), .Z(n41593) );
  OR U54471 ( .A(n41594), .B(n41593), .Z(n41595) );
  AND U54472 ( .A(n41596), .B(n41595), .Z(n41597) );
  OR U54473 ( .A(n41598), .B(n41597), .Z(n41599) );
  NAND U54474 ( .A(n41600), .B(n41599), .Z(n41601) );
  NAND U54475 ( .A(n41602), .B(n41601), .Z(n41603) );
  ANDN U54476 ( .B(y[4518]), .A(x[4518]), .Z(n56756) );
  ANDN U54477 ( .B(n41603), .A(n56756), .Z(n41605) );
  ANDN U54478 ( .B(n41605), .A(n41604), .Z(n41609) );
  NAND U54479 ( .A(n41607), .B(n41606), .Z(n41608) );
  OR U54480 ( .A(n41609), .B(n41608), .Z(n41610) );
  AND U54481 ( .A(n41611), .B(n41610), .Z(n41615) );
  NAND U54482 ( .A(n41613), .B(n41612), .Z(n41614) );
  OR U54483 ( .A(n41615), .B(n41614), .Z(n41616) );
  AND U54484 ( .A(n41617), .B(n41616), .Z(n41618) );
  ANDN U54485 ( .B(n41619), .A(n41618), .Z(n41620) );
  NAND U54486 ( .A(n41621), .B(n41620), .Z(n41622) );
  NANDN U54487 ( .A(n41623), .B(n41622), .Z(n41624) );
  OR U54488 ( .A(n41625), .B(n41624), .Z(n41626) );
  AND U54489 ( .A(n41627), .B(n41626), .Z(n41629) );
  NAND U54490 ( .A(n41629), .B(n41628), .Z(n41630) );
  NANDN U54491 ( .A(n41631), .B(n41630), .Z(n41632) );
  AND U54492 ( .A(n41633), .B(n41632), .Z(n41635) );
  NAND U54493 ( .A(n41635), .B(n41634), .Z(n41636) );
  NANDN U54494 ( .A(n41637), .B(n41636), .Z(n41638) );
  AND U54495 ( .A(n41639), .B(n41638), .Z(n41641) );
  NAND U54496 ( .A(n41641), .B(n41640), .Z(n41642) );
  AND U54497 ( .A(n41642), .B(n56774), .Z(n41643) );
  NANDN U54498 ( .A(x[4530]), .B(y[4530]), .Z(n56768) );
  AND U54499 ( .A(n41643), .B(n56768), .Z(n41644) );
  NOR U54500 ( .A(n41645), .B(n41644), .Z(n41647) );
  NAND U54501 ( .A(n41647), .B(n41646), .Z(n41649) );
  AND U54502 ( .A(n41649), .B(n41648), .Z(n41650) );
  NANDN U54503 ( .A(x[4532]), .B(y[4532]), .Z(n56775) );
  NAND U54504 ( .A(n41650), .B(n56775), .Z(n41651) );
  NANDN U54505 ( .A(n41652), .B(n41651), .Z(n41653) );
  AND U54506 ( .A(n41654), .B(n41653), .Z(n41656) );
  NAND U54507 ( .A(n41656), .B(n41655), .Z(n41657) );
  NANDN U54508 ( .A(n41658), .B(n41657), .Z(n41659) );
  AND U54509 ( .A(n56788), .B(n41659), .Z(n41661) );
  NANDN U54510 ( .A(x[4536]), .B(y[4536]), .Z(n41660) );
  AND U54511 ( .A(n41661), .B(n41660), .Z(n41662) );
  OR U54512 ( .A(n41663), .B(n41662), .Z(n41664) );
  AND U54513 ( .A(n41665), .B(n41664), .Z(n41669) );
  NAND U54514 ( .A(n41667), .B(n41666), .Z(n41668) );
  OR U54515 ( .A(n41669), .B(n41668), .Z(n41670) );
  AND U54516 ( .A(n41671), .B(n41670), .Z(n41675) );
  NAND U54517 ( .A(n41673), .B(n41672), .Z(n41674) );
  OR U54518 ( .A(n41675), .B(n41674), .Z(n41676) );
  AND U54519 ( .A(n41677), .B(n41676), .Z(n41681) );
  NAND U54520 ( .A(n41679), .B(n41678), .Z(n41680) );
  OR U54521 ( .A(n41681), .B(n41680), .Z(n41682) );
  AND U54522 ( .A(n41683), .B(n41682), .Z(n41687) );
  NAND U54523 ( .A(n41685), .B(n41684), .Z(n41686) );
  OR U54524 ( .A(n41687), .B(n41686), .Z(n41688) );
  AND U54525 ( .A(n41689), .B(n41688), .Z(n41690) );
  OR U54526 ( .A(n41691), .B(n41690), .Z(n41692) );
  NAND U54527 ( .A(n41693), .B(n41692), .Z(n41694) );
  AND U54528 ( .A(n41695), .B(n41694), .Z(n41696) );
  NOR U54529 ( .A(n56812), .B(n41696), .Z(n41697) );
  NANDN U54530 ( .A(n51603), .B(n41697), .Z(n41698) );
  AND U54531 ( .A(n41699), .B(n41698), .Z(n41701) );
  NAND U54532 ( .A(n41701), .B(n41700), .Z(n41702) );
  NANDN U54533 ( .A(n41703), .B(n41702), .Z(n41704) );
  AND U54534 ( .A(n41705), .B(n41704), .Z(n41706) );
  NANDN U54535 ( .A(n41707), .B(n41706), .Z(n41708) );
  AND U54536 ( .A(n41709), .B(n41708), .Z(n41711) );
  NANDN U54537 ( .A(x[4554]), .B(y[4554]), .Z(n41710) );
  NAND U54538 ( .A(n41711), .B(n41710), .Z(n41713) );
  ANDN U54539 ( .B(n41713), .A(n41712), .Z(n41715) );
  ANDN U54540 ( .B(n41715), .A(n41714), .Z(n41716) );
  OR U54541 ( .A(n41717), .B(n41716), .Z(n41718) );
  NAND U54542 ( .A(n41719), .B(n41718), .Z(n41720) );
  NANDN U54543 ( .A(n41721), .B(n41720), .Z(n41725) );
  AND U54544 ( .A(n41723), .B(n41722), .Z(n41724) );
  NAND U54545 ( .A(n41725), .B(n41724), .Z(n41726) );
  NANDN U54546 ( .A(n41727), .B(n41726), .Z(n41729) );
  ANDN U54547 ( .B(y[4560]), .A(x[4560]), .Z(n41728) );
  OR U54548 ( .A(n41729), .B(n41728), .Z(n41730) );
  NAND U54549 ( .A(n41731), .B(n41730), .Z(n41732) );
  NANDN U54550 ( .A(n51601), .B(n41732), .Z(n41734) );
  ANDN U54551 ( .B(y[4562]), .A(x[4562]), .Z(n41733) );
  OR U54552 ( .A(n41734), .B(n41733), .Z(n41735) );
  NAND U54553 ( .A(n41736), .B(n41735), .Z(n41737) );
  NAND U54554 ( .A(n51602), .B(n41737), .Z(n41738) );
  NANDN U54555 ( .A(n41738), .B(n56828), .Z(n41739) );
  AND U54556 ( .A(n41740), .B(n41739), .Z(n41741) );
  OR U54557 ( .A(n41742), .B(n41741), .Z(n41743) );
  NAND U54558 ( .A(n41744), .B(n41743), .Z(n41745) );
  NANDN U54559 ( .A(n56833), .B(n41745), .Z(n41746) );
  ANDN U54560 ( .B(y[4568]), .A(x[4568]), .Z(n56831) );
  OR U54561 ( .A(n41746), .B(n56831), .Z(n41747) );
  AND U54562 ( .A(n41748), .B(n41747), .Z(n41750) );
  NAND U54563 ( .A(n41750), .B(n41749), .Z(n41751) );
  NANDN U54564 ( .A(n41752), .B(n41751), .Z(n41753) );
  AND U54565 ( .A(n41754), .B(n41753), .Z(n41756) );
  NAND U54566 ( .A(n41756), .B(n41755), .Z(n41757) );
  NANDN U54567 ( .A(n41758), .B(n41757), .Z(n41759) );
  AND U54568 ( .A(n41760), .B(n41759), .Z(n41762) );
  NAND U54569 ( .A(n41762), .B(n41761), .Z(n41764) );
  AND U54570 ( .A(n41764), .B(n41763), .Z(n41765) );
  NANDN U54571 ( .A(x[4574]), .B(y[4574]), .Z(n56839) );
  AND U54572 ( .A(n41765), .B(n56839), .Z(n41766) );
  NOR U54573 ( .A(n41767), .B(n41766), .Z(n41769) );
  NAND U54574 ( .A(n41769), .B(n41768), .Z(n41771) );
  AND U54575 ( .A(n41771), .B(n41770), .Z(n41773) );
  NANDN U54576 ( .A(x[4576]), .B(y[4576]), .Z(n41772) );
  AND U54577 ( .A(n41773), .B(n41772), .Z(n41777) );
  AND U54578 ( .A(n41775), .B(n41774), .Z(n41776) );
  NANDN U54579 ( .A(n41777), .B(n41776), .Z(n41779) );
  AND U54580 ( .A(n41779), .B(n41778), .Z(n41781) );
  NANDN U54581 ( .A(x[4578]), .B(y[4578]), .Z(n41780) );
  AND U54582 ( .A(n41781), .B(n41780), .Z(n41782) );
  NOR U54583 ( .A(n41783), .B(n41782), .Z(n41785) );
  NAND U54584 ( .A(n41785), .B(n41784), .Z(n41787) );
  AND U54585 ( .A(n41787), .B(n41786), .Z(n41789) );
  NANDN U54586 ( .A(x[4580]), .B(y[4580]), .Z(n41788) );
  AND U54587 ( .A(n41789), .B(n41788), .Z(n41790) );
  NOR U54588 ( .A(n41791), .B(n41790), .Z(n41793) );
  NAND U54589 ( .A(n41793), .B(n41792), .Z(n41795) );
  AND U54590 ( .A(n41795), .B(n41794), .Z(n41797) );
  NANDN U54591 ( .A(x[4582]), .B(y[4582]), .Z(n41796) );
  AND U54592 ( .A(n41797), .B(n41796), .Z(n41798) );
  NOR U54593 ( .A(n41799), .B(n41798), .Z(n41801) );
  NAND U54594 ( .A(n41801), .B(n41800), .Z(n41802) );
  AND U54595 ( .A(n41802), .B(n56854), .Z(n41803) );
  NANDN U54596 ( .A(n41804), .B(n41803), .Z(n41805) );
  NAND U54597 ( .A(n41806), .B(n41805), .Z(n41807) );
  NANDN U54598 ( .A(n56856), .B(n41807), .Z(n41808) );
  ANDN U54599 ( .B(y[4586]), .A(x[4586]), .Z(n56853) );
  OR U54600 ( .A(n41808), .B(n56853), .Z(n41809) );
  NAND U54601 ( .A(n41810), .B(n41809), .Z(n41811) );
  NANDN U54602 ( .A(n41812), .B(n41811), .Z(n41813) );
  ANDN U54603 ( .B(y[4588]), .A(x[4588]), .Z(n56857) );
  OR U54604 ( .A(n41813), .B(n56857), .Z(n41814) );
  NAND U54605 ( .A(n41815), .B(n41814), .Z(n41816) );
  NANDN U54606 ( .A(n41817), .B(n41816), .Z(n41818) );
  ANDN U54607 ( .B(n41819), .A(n41818), .Z(n41823) );
  NAND U54608 ( .A(n41821), .B(n41820), .Z(n41822) );
  OR U54609 ( .A(n41823), .B(n41822), .Z(n41824) );
  AND U54610 ( .A(n41825), .B(n41824), .Z(n41829) );
  NAND U54611 ( .A(n41827), .B(n41826), .Z(n41828) );
  OR U54612 ( .A(n41829), .B(n41828), .Z(n41830) );
  AND U54613 ( .A(n41831), .B(n41830), .Z(n41832) );
  OR U54614 ( .A(n41833), .B(n41832), .Z(n41834) );
  NAND U54615 ( .A(n41835), .B(n41834), .Z(n41836) );
  AND U54616 ( .A(n41837), .B(n41836), .Z(n41841) );
  NANDN U54617 ( .A(x[4598]), .B(y[4598]), .Z(n41839) );
  AND U54618 ( .A(n41839), .B(n41838), .Z(n41840) );
  NANDN U54619 ( .A(n41841), .B(n41840), .Z(n41842) );
  NANDN U54620 ( .A(n41843), .B(n41842), .Z(n41844) );
  AND U54621 ( .A(n41845), .B(n41844), .Z(n41847) );
  NANDN U54622 ( .A(x[4600]), .B(y[4600]), .Z(n41846) );
  AND U54623 ( .A(n41847), .B(n41846), .Z(n41851) );
  NAND U54624 ( .A(n41849), .B(n41848), .Z(n41850) );
  OR U54625 ( .A(n41851), .B(n41850), .Z(n41852) );
  AND U54626 ( .A(n41853), .B(n41852), .Z(n41857) );
  NAND U54627 ( .A(n41855), .B(n41854), .Z(n41856) );
  OR U54628 ( .A(n41857), .B(n41856), .Z(n41858) );
  AND U54629 ( .A(n41859), .B(n41858), .Z(n41863) );
  NAND U54630 ( .A(n41861), .B(n41860), .Z(n41862) );
  OR U54631 ( .A(n41863), .B(n41862), .Z(n41864) );
  AND U54632 ( .A(n41865), .B(n41864), .Z(n41869) );
  NAND U54633 ( .A(n41867), .B(n41866), .Z(n41868) );
  OR U54634 ( .A(n41869), .B(n41868), .Z(n41870) );
  AND U54635 ( .A(n41871), .B(n41870), .Z(n41872) );
  OR U54636 ( .A(n41873), .B(n41872), .Z(n41874) );
  NAND U54637 ( .A(n41875), .B(n41874), .Z(n41876) );
  AND U54638 ( .A(n41877), .B(n41876), .Z(n41878) );
  NOR U54639 ( .A(n51595), .B(n41878), .Z(n41879) );
  NANDN U54640 ( .A(n41880), .B(n41879), .Z(n41881) );
  AND U54641 ( .A(n41882), .B(n41881), .Z(n41884) );
  NAND U54642 ( .A(n41884), .B(n41883), .Z(n41885) );
  NANDN U54643 ( .A(n41886), .B(n41885), .Z(n41887) );
  AND U54644 ( .A(n41888), .B(n41887), .Z(n41889) );
  NANDN U54645 ( .A(n41890), .B(n41889), .Z(n41891) );
  NAND U54646 ( .A(n41892), .B(n41891), .Z(n41893) );
  NANDN U54647 ( .A(n41894), .B(n41893), .Z(n41895) );
  AND U54648 ( .A(n41895), .B(n56889), .Z(n41896) );
  NANDN U54649 ( .A(x[4618]), .B(y[4618]), .Z(n51593) );
  AND U54650 ( .A(n41896), .B(n51593), .Z(n41897) );
  NOR U54651 ( .A(n41898), .B(n41897), .Z(n41900) );
  NAND U54652 ( .A(n41900), .B(n41899), .Z(n41902) );
  AND U54653 ( .A(n41902), .B(n41901), .Z(n41903) );
  NANDN U54654 ( .A(x[4620]), .B(y[4620]), .Z(n56890) );
  AND U54655 ( .A(n41903), .B(n56890), .Z(n41907) );
  AND U54656 ( .A(n41905), .B(n41904), .Z(n41906) );
  NANDN U54657 ( .A(n41907), .B(n41906), .Z(n41909) );
  AND U54658 ( .A(n41909), .B(n41908), .Z(n41910) );
  NANDN U54659 ( .A(n41911), .B(n41910), .Z(n41912) );
  NAND U54660 ( .A(n41913), .B(n41912), .Z(n41915) );
  AND U54661 ( .A(n41915), .B(n41914), .Z(n41917) );
  NANDN U54662 ( .A(x[4624]), .B(y[4624]), .Z(n41916) );
  AND U54663 ( .A(n41917), .B(n41916), .Z(n41918) );
  NOR U54664 ( .A(n41919), .B(n41918), .Z(n41921) );
  NAND U54665 ( .A(n41921), .B(n41920), .Z(n41923) );
  AND U54666 ( .A(n41923), .B(n41922), .Z(n41925) );
  NANDN U54667 ( .A(x[4626]), .B(y[4626]), .Z(n41924) );
  AND U54668 ( .A(n41925), .B(n41924), .Z(n41926) );
  NOR U54669 ( .A(n41927), .B(n41926), .Z(n41929) );
  NAND U54670 ( .A(n41929), .B(n41928), .Z(n41931) );
  AND U54671 ( .A(n41931), .B(n41930), .Z(n41933) );
  NANDN U54672 ( .A(x[4628]), .B(y[4628]), .Z(n41932) );
  AND U54673 ( .A(n41933), .B(n41932), .Z(n41934) );
  NOR U54674 ( .A(n41935), .B(n41934), .Z(n41937) );
  NAND U54675 ( .A(n41937), .B(n41936), .Z(n41939) );
  AND U54676 ( .A(n41939), .B(n41938), .Z(n41941) );
  NANDN U54677 ( .A(x[4630]), .B(y[4630]), .Z(n41940) );
  AND U54678 ( .A(n41941), .B(n41940), .Z(n41942) );
  NOR U54679 ( .A(n41943), .B(n41942), .Z(n41945) );
  NAND U54680 ( .A(n41945), .B(n41944), .Z(n41947) );
  AND U54681 ( .A(n41947), .B(n41946), .Z(n41949) );
  NANDN U54682 ( .A(x[4632]), .B(y[4632]), .Z(n41948) );
  AND U54683 ( .A(n41949), .B(n41948), .Z(n41953) );
  AND U54684 ( .A(n41951), .B(n41950), .Z(n41952) );
  NANDN U54685 ( .A(n41953), .B(n41952), .Z(n41957) );
  NANDN U54686 ( .A(x[4634]), .B(y[4634]), .Z(n41954) );
  AND U54687 ( .A(n41955), .B(n41954), .Z(n41956) );
  NAND U54688 ( .A(n41957), .B(n41956), .Z(n41958) );
  NANDN U54689 ( .A(n41959), .B(n41958), .Z(n41960) );
  AND U54690 ( .A(n41961), .B(n41960), .Z(n41964) );
  NAND U54691 ( .A(n41963), .B(n41962), .Z(n56907) );
  OR U54692 ( .A(n41964), .B(n56907), .Z(n41965) );
  AND U54693 ( .A(n41966), .B(n41965), .Z(n41967) );
  NAND U54694 ( .A(n41967), .B(n56908), .Z(n41968) );
  NANDN U54695 ( .A(n41969), .B(n41968), .Z(n41970) );
  AND U54696 ( .A(n41971), .B(n41970), .Z(n41975) );
  AND U54697 ( .A(n41973), .B(n41972), .Z(n41974) );
  NANDN U54698 ( .A(n41975), .B(n41974), .Z(n41976) );
  AND U54699 ( .A(n41977), .B(n41976), .Z(n41981) );
  NAND U54700 ( .A(n41979), .B(n41978), .Z(n41980) );
  OR U54701 ( .A(n41981), .B(n41980), .Z(n41982) );
  AND U54702 ( .A(n41983), .B(n41982), .Z(n41984) );
  OR U54703 ( .A(n41985), .B(n41984), .Z(n41986) );
  NAND U54704 ( .A(n41987), .B(n41986), .Z(n41988) );
  AND U54705 ( .A(n56919), .B(n41988), .Z(n41991) );
  NANDN U54706 ( .A(x[4648]), .B(y[4648]), .Z(n51583) );
  NAND U54707 ( .A(n51583), .B(n41989), .Z(n41990) );
  OR U54708 ( .A(n41991), .B(n41990), .Z(n41992) );
  AND U54709 ( .A(n41993), .B(n41992), .Z(n41994) );
  NANDN U54710 ( .A(n56920), .B(n41994), .Z(n41995) );
  NAND U54711 ( .A(n41996), .B(n41995), .Z(n41997) );
  NANDN U54712 ( .A(n41998), .B(n41997), .Z(n42000) );
  AND U54713 ( .A(n42000), .B(n41999), .Z(n42001) );
  NANDN U54714 ( .A(x[4652]), .B(y[4652]), .Z(n56925) );
  AND U54715 ( .A(n42001), .B(n56925), .Z(n42002) );
  NOR U54716 ( .A(n42003), .B(n42002), .Z(n42005) );
  NAND U54717 ( .A(n42005), .B(n42004), .Z(n42007) );
  AND U54718 ( .A(n42007), .B(n42006), .Z(n42009) );
  NANDN U54719 ( .A(x[4654]), .B(y[4654]), .Z(n42008) );
  AND U54720 ( .A(n42009), .B(n42008), .Z(n42010) );
  NOR U54721 ( .A(n42011), .B(n42010), .Z(n42013) );
  NAND U54722 ( .A(n42013), .B(n42012), .Z(n42015) );
  AND U54723 ( .A(n42015), .B(n42014), .Z(n42017) );
  NANDN U54724 ( .A(x[4656]), .B(y[4656]), .Z(n42016) );
  AND U54725 ( .A(n42017), .B(n42016), .Z(n42018) );
  NOR U54726 ( .A(n42019), .B(n42018), .Z(n42021) );
  NAND U54727 ( .A(n42021), .B(n42020), .Z(n42023) );
  AND U54728 ( .A(n42023), .B(n42022), .Z(n42024) );
  NANDN U54729 ( .A(n42025), .B(n42024), .Z(n42026) );
  NAND U54730 ( .A(n42027), .B(n42026), .Z(n42028) );
  NANDN U54731 ( .A(n56935), .B(n42028), .Z(n42030) );
  ANDN U54732 ( .B(y[4660]), .A(x[4660]), .Z(n42029) );
  OR U54733 ( .A(n42030), .B(n42029), .Z(n42031) );
  NAND U54734 ( .A(n42032), .B(n42031), .Z(n42033) );
  NANDN U54735 ( .A(n42034), .B(n42033), .Z(n42035) );
  ANDN U54736 ( .B(y[4662]), .A(x[4662]), .Z(n51581) );
  OR U54737 ( .A(n42035), .B(n51581), .Z(n42036) );
  NAND U54738 ( .A(n42037), .B(n42036), .Z(n42038) );
  NANDN U54739 ( .A(n42039), .B(n42038), .Z(n42041) );
  OR U54740 ( .A(n42041), .B(n42040), .Z(n42042) );
  NAND U54741 ( .A(n42043), .B(n42042), .Z(n42047) );
  NAND U54742 ( .A(n42045), .B(n42044), .Z(n42046) );
  ANDN U54743 ( .B(n42047), .A(n42046), .Z(n42051) );
  NAND U54744 ( .A(n42049), .B(n42048), .Z(n42050) );
  OR U54745 ( .A(n42051), .B(n42050), .Z(n42052) );
  AND U54746 ( .A(n42053), .B(n42052), .Z(n42057) );
  NAND U54747 ( .A(n42055), .B(n42054), .Z(n42056) );
  OR U54748 ( .A(n42057), .B(n42056), .Z(n42058) );
  AND U54749 ( .A(n42059), .B(n42058), .Z(n42063) );
  NAND U54750 ( .A(n42061), .B(n42060), .Z(n42062) );
  OR U54751 ( .A(n42063), .B(n42062), .Z(n42064) );
  AND U54752 ( .A(n42065), .B(n42064), .Z(n42069) );
  NAND U54753 ( .A(n42067), .B(n42066), .Z(n42068) );
  OR U54754 ( .A(n42069), .B(n42068), .Z(n42070) );
  AND U54755 ( .A(n42071), .B(n42070), .Z(n42075) );
  NAND U54756 ( .A(n42073), .B(n42072), .Z(n42074) );
  OR U54757 ( .A(n42075), .B(n42074), .Z(n42076) );
  AND U54758 ( .A(n42077), .B(n42076), .Z(n42081) );
  AND U54759 ( .A(n42079), .B(n42078), .Z(n42080) );
  NANDN U54760 ( .A(n42081), .B(n42080), .Z(n42082) );
  NAND U54761 ( .A(n42083), .B(n42082), .Z(n42084) );
  AND U54762 ( .A(n42085), .B(n42084), .Z(n42087) );
  NANDN U54763 ( .A(x[4680]), .B(y[4680]), .Z(n56954) );
  NAND U54764 ( .A(n56954), .B(n51577), .Z(n42086) );
  OR U54765 ( .A(n42087), .B(n42086), .Z(n42088) );
  AND U54766 ( .A(n42089), .B(n42088), .Z(n42091) );
  NAND U54767 ( .A(n42091), .B(n42090), .Z(n42092) );
  NANDN U54768 ( .A(n42093), .B(n42092), .Z(n42094) );
  AND U54769 ( .A(n42095), .B(n42094), .Z(n42096) );
  NANDN U54770 ( .A(n42097), .B(n42096), .Z(n42098) );
  NAND U54771 ( .A(n42099), .B(n42098), .Z(n42100) );
  NANDN U54772 ( .A(n42101), .B(n42100), .Z(n42103) );
  IV U54773 ( .A(n42102), .Z(n51575) );
  AND U54774 ( .A(n42103), .B(n51575), .Z(n42104) );
  NANDN U54775 ( .A(n42105), .B(n42104), .Z(n42106) );
  AND U54776 ( .A(n42107), .B(n42106), .Z(n42108) );
  ANDN U54777 ( .B(n56965), .A(n42108), .Z(n42109) );
  NANDN U54778 ( .A(x[4688]), .B(y[4688]), .Z(n51576) );
  AND U54779 ( .A(n42109), .B(n51576), .Z(n42110) );
  NOR U54780 ( .A(n42111), .B(n42110), .Z(n42113) );
  NAND U54781 ( .A(n42113), .B(n42112), .Z(n42115) );
  IV U54782 ( .A(n42114), .Z(n56967) );
  AND U54783 ( .A(n42115), .B(n56967), .Z(n42116) );
  NANDN U54784 ( .A(n56964), .B(n42116), .Z(n42117) );
  NAND U54785 ( .A(n42118), .B(n42117), .Z(n42119) );
  NANDN U54786 ( .A(n42120), .B(n42119), .Z(n42121) );
  ANDN U54787 ( .B(y[4692]), .A(x[4692]), .Z(n56968) );
  OR U54788 ( .A(n42121), .B(n56968), .Z(n42122) );
  NAND U54789 ( .A(n42123), .B(n42122), .Z(n42124) );
  NANDN U54790 ( .A(n56974), .B(n42124), .Z(n42126) );
  ANDN U54791 ( .B(y[4694]), .A(x[4694]), .Z(n42125) );
  OR U54792 ( .A(n42126), .B(n42125), .Z(n42127) );
  NAND U54793 ( .A(n42128), .B(n42127), .Z(n42129) );
  NANDN U54794 ( .A(n42130), .B(n42129), .Z(n42131) );
  NAND U54795 ( .A(n42132), .B(n42131), .Z(n42134) );
  ANDN U54796 ( .B(y[4698]), .A(x[4698]), .Z(n42133) );
  ANDN U54797 ( .B(n42134), .A(n42133), .Z(n42136) );
  ANDN U54798 ( .B(n42136), .A(n42135), .Z(n42140) );
  NAND U54799 ( .A(n42138), .B(n42137), .Z(n42139) );
  OR U54800 ( .A(n42140), .B(n42139), .Z(n42141) );
  AND U54801 ( .A(n42142), .B(n42141), .Z(n42146) );
  NAND U54802 ( .A(n42144), .B(n42143), .Z(n42145) );
  OR U54803 ( .A(n42146), .B(n42145), .Z(n42147) );
  AND U54804 ( .A(n42148), .B(n42147), .Z(n42152) );
  NAND U54805 ( .A(n42150), .B(n42149), .Z(n42151) );
  OR U54806 ( .A(n42152), .B(n42151), .Z(n42153) );
  AND U54807 ( .A(n42154), .B(n42153), .Z(n42155) );
  OR U54808 ( .A(n42156), .B(n42155), .Z(n42157) );
  NAND U54809 ( .A(n42158), .B(n42157), .Z(n42159) );
  AND U54810 ( .A(n42160), .B(n42159), .Z(n42161) );
  NOR U54811 ( .A(n56987), .B(n42161), .Z(n42162) );
  NANDN U54812 ( .A(n56989), .B(n42162), .Z(n42163) );
  AND U54813 ( .A(n42164), .B(n42163), .Z(n42166) );
  NAND U54814 ( .A(n42166), .B(n42165), .Z(n42167) );
  NANDN U54815 ( .A(n42168), .B(n42167), .Z(n42169) );
  AND U54816 ( .A(n42170), .B(n42169), .Z(n42171) );
  NANDN U54817 ( .A(n42172), .B(n42171), .Z(n42173) );
  NAND U54818 ( .A(n42174), .B(n42173), .Z(n42175) );
  NANDN U54819 ( .A(n42176), .B(n42175), .Z(n42178) );
  AND U54820 ( .A(n42178), .B(n42177), .Z(n42180) );
  NANDN U54821 ( .A(x[4714]), .B(y[4714]), .Z(n42179) );
  AND U54822 ( .A(n42180), .B(n42179), .Z(n42181) );
  NOR U54823 ( .A(n42182), .B(n42181), .Z(n42184) );
  NAND U54824 ( .A(n42184), .B(n42183), .Z(n42188) );
  NANDN U54825 ( .A(x[4716]), .B(y[4716]), .Z(n42185) );
  AND U54826 ( .A(n42186), .B(n42185), .Z(n42187) );
  NAND U54827 ( .A(n42188), .B(n42187), .Z(n42189) );
  NANDN U54828 ( .A(n42190), .B(n42189), .Z(n42191) );
  NAND U54829 ( .A(n42192), .B(n42191), .Z(n42193) );
  NANDN U54830 ( .A(n42194), .B(n42193), .Z(n42195) );
  AND U54831 ( .A(n42196), .B(n42195), .Z(n42198) );
  NANDN U54832 ( .A(x[4720]), .B(y[4720]), .Z(n42197) );
  NAND U54833 ( .A(n42198), .B(n42197), .Z(n42199) );
  NANDN U54834 ( .A(n42200), .B(n42199), .Z(n42201) );
  AND U54835 ( .A(n57005), .B(n42201), .Z(n42203) );
  NAND U54836 ( .A(n42203), .B(n42202), .Z(n42204) );
  NANDN U54837 ( .A(n42205), .B(n42204), .Z(n42206) );
  AND U54838 ( .A(n42207), .B(n42206), .Z(n42208) );
  OR U54839 ( .A(n42209), .B(n42208), .Z(n42210) );
  NAND U54840 ( .A(n42211), .B(n42210), .Z(n42212) );
  AND U54841 ( .A(n42213), .B(n42212), .Z(n42214) );
  ANDN U54842 ( .B(n51572), .A(n42214), .Z(n42215) );
  NAND U54843 ( .A(n57014), .B(n42215), .Z(n42216) );
  NANDN U54844 ( .A(n42217), .B(n42216), .Z(n42218) );
  OR U54845 ( .A(n42219), .B(n42218), .Z(n42220) );
  NAND U54846 ( .A(n42221), .B(n42220), .Z(n42222) );
  NANDN U54847 ( .A(n42223), .B(n42222), .Z(n42225) );
  AND U54848 ( .A(n42225), .B(n42224), .Z(n42226) );
  NANDN U54849 ( .A(x[4732]), .B(y[4732]), .Z(n57016) );
  AND U54850 ( .A(n42226), .B(n57016), .Z(n42227) );
  NOR U54851 ( .A(n42228), .B(n42227), .Z(n42230) );
  NAND U54852 ( .A(n42230), .B(n42229), .Z(n42232) );
  AND U54853 ( .A(n42232), .B(n42231), .Z(n42234) );
  NANDN U54854 ( .A(x[4734]), .B(y[4734]), .Z(n42233) );
  AND U54855 ( .A(n42234), .B(n42233), .Z(n42235) );
  NOR U54856 ( .A(n42236), .B(n42235), .Z(n42238) );
  NAND U54857 ( .A(n42238), .B(n42237), .Z(n42240) );
  AND U54858 ( .A(n42240), .B(n42239), .Z(n42242) );
  NANDN U54859 ( .A(x[4736]), .B(y[4736]), .Z(n42241) );
  AND U54860 ( .A(n42242), .B(n42241), .Z(n42243) );
  NOR U54861 ( .A(n42244), .B(n42243), .Z(n42246) );
  NAND U54862 ( .A(n42246), .B(n42245), .Z(n42248) );
  AND U54863 ( .A(n42248), .B(n42247), .Z(n42250) );
  NANDN U54864 ( .A(x[4738]), .B(y[4738]), .Z(n42249) );
  NAND U54865 ( .A(n42250), .B(n42249), .Z(n42251) );
  NAND U54866 ( .A(n42252), .B(n42251), .Z(n42254) );
  AND U54867 ( .A(n42254), .B(n42253), .Z(n42256) );
  NANDN U54868 ( .A(x[4740]), .B(y[4740]), .Z(n42255) );
  AND U54869 ( .A(n42256), .B(n42255), .Z(n42257) );
  NOR U54870 ( .A(n42258), .B(n42257), .Z(n42260) );
  NAND U54871 ( .A(n42260), .B(n42259), .Z(n42261) );
  AND U54872 ( .A(n42261), .B(n57028), .Z(n42263) );
  NANDN U54873 ( .A(x[4742]), .B(y[4742]), .Z(n42262) );
  AND U54874 ( .A(n42263), .B(n42262), .Z(n42264) );
  NOR U54875 ( .A(n42265), .B(n42264), .Z(n42267) );
  NAND U54876 ( .A(n42267), .B(n42266), .Z(n42269) );
  AND U54877 ( .A(n42269), .B(n42268), .Z(n42270) );
  NANDN U54878 ( .A(x[4744]), .B(y[4744]), .Z(n57029) );
  NAND U54879 ( .A(n42270), .B(n57029), .Z(n42271) );
  NANDN U54880 ( .A(n42272), .B(n42271), .Z(n42273) );
  AND U54881 ( .A(n57034), .B(n42273), .Z(n42275) );
  NAND U54882 ( .A(n42275), .B(n42274), .Z(n42276) );
  NANDN U54883 ( .A(n42277), .B(n42276), .Z(n42278) );
  AND U54884 ( .A(n42279), .B(n42278), .Z(n42280) );
  NANDN U54885 ( .A(x[4748]), .B(y[4748]), .Z(n57035) );
  AND U54886 ( .A(n42280), .B(n57035), .Z(n42281) );
  OR U54887 ( .A(n42282), .B(n42281), .Z(n42283) );
  AND U54888 ( .A(n42284), .B(n42283), .Z(n42288) );
  NAND U54889 ( .A(n42286), .B(n42285), .Z(n42287) );
  OR U54890 ( .A(n42288), .B(n42287), .Z(n42289) );
  AND U54891 ( .A(n42290), .B(n42289), .Z(n42294) );
  NAND U54892 ( .A(n42292), .B(n42291), .Z(n42293) );
  OR U54893 ( .A(n42294), .B(n42293), .Z(n42295) );
  AND U54894 ( .A(n42296), .B(n42295), .Z(n42300) );
  NAND U54895 ( .A(n42298), .B(n42297), .Z(n42299) );
  OR U54896 ( .A(n42300), .B(n42299), .Z(n42301) );
  AND U54897 ( .A(n42302), .B(n42301), .Z(n42306) );
  NAND U54898 ( .A(n42304), .B(n42303), .Z(n42305) );
  OR U54899 ( .A(n42306), .B(n42305), .Z(n42307) );
  AND U54900 ( .A(n42308), .B(n42307), .Z(n42312) );
  NAND U54901 ( .A(n42310), .B(n42309), .Z(n42311) );
  OR U54902 ( .A(n42312), .B(n42311), .Z(n42313) );
  AND U54903 ( .A(n42314), .B(n42313), .Z(n42318) );
  AND U54904 ( .A(n42316), .B(n42315), .Z(n42317) );
  NANDN U54905 ( .A(n42318), .B(n42317), .Z(n42319) );
  AND U54906 ( .A(n42320), .B(n42319), .Z(n42324) );
  NAND U54907 ( .A(n42322), .B(n42321), .Z(n42323) );
  OR U54908 ( .A(n42324), .B(n42323), .Z(n42325) );
  AND U54909 ( .A(n42326), .B(n42325), .Z(n42330) );
  NAND U54910 ( .A(n42328), .B(n42327), .Z(n42329) );
  OR U54911 ( .A(n42330), .B(n42329), .Z(n42331) );
  AND U54912 ( .A(n42332), .B(n42331), .Z(n42333) );
  NANDN U54913 ( .A(x[4766]), .B(y[4766]), .Z(n51563) );
  AND U54914 ( .A(n42333), .B(n51563), .Z(n42337) );
  NAND U54915 ( .A(n42335), .B(n42334), .Z(n42336) );
  OR U54916 ( .A(n42337), .B(n42336), .Z(n42338) );
  AND U54917 ( .A(n42339), .B(n42338), .Z(n42340) );
  OR U54918 ( .A(n42341), .B(n42340), .Z(n42342) );
  NAND U54919 ( .A(n42343), .B(n42342), .Z(n42344) );
  AND U54920 ( .A(n42345), .B(n42344), .Z(n42346) );
  ANDN U54921 ( .B(n42347), .A(n42346), .Z(n42351) );
  NAND U54922 ( .A(n42349), .B(n42348), .Z(n42350) );
  OR U54923 ( .A(n42351), .B(n42350), .Z(n42352) );
  AND U54924 ( .A(n42353), .B(n42352), .Z(n42357) );
  NAND U54925 ( .A(n42355), .B(n42354), .Z(n42356) );
  OR U54926 ( .A(n42357), .B(n42356), .Z(n42358) );
  AND U54927 ( .A(n42359), .B(n42358), .Z(n42360) );
  OR U54928 ( .A(n42361), .B(n42360), .Z(n42362) );
  NAND U54929 ( .A(n42363), .B(n42362), .Z(n42364) );
  AND U54930 ( .A(n42365), .B(n42364), .Z(n42366) );
  ANDN U54931 ( .B(n42367), .A(n42366), .Z(n42369) );
  NANDN U54932 ( .A(x[4780]), .B(y[4780]), .Z(n42368) );
  AND U54933 ( .A(n42369), .B(n42368), .Z(n42373) );
  NAND U54934 ( .A(n42371), .B(n42370), .Z(n42372) );
  OR U54935 ( .A(n42373), .B(n42372), .Z(n42374) );
  AND U54936 ( .A(n42375), .B(n42374), .Z(n42379) );
  NAND U54937 ( .A(n42377), .B(n42376), .Z(n42378) );
  OR U54938 ( .A(n42379), .B(n42378), .Z(n42380) );
  AND U54939 ( .A(n42381), .B(n42380), .Z(n42385) );
  NAND U54940 ( .A(n42383), .B(n42382), .Z(n42384) );
  OR U54941 ( .A(n42385), .B(n42384), .Z(n42386) );
  AND U54942 ( .A(n42387), .B(n42386), .Z(n42391) );
  NAND U54943 ( .A(n42389), .B(n42388), .Z(n42390) );
  OR U54944 ( .A(n42391), .B(n42390), .Z(n42392) );
  AND U54945 ( .A(n42393), .B(n42392), .Z(n42397) );
  NAND U54946 ( .A(n42395), .B(n42394), .Z(n42396) );
  OR U54947 ( .A(n42397), .B(n42396), .Z(n42398) );
  AND U54948 ( .A(n42399), .B(n42398), .Z(n42403) );
  NAND U54949 ( .A(n42401), .B(n42400), .Z(n42402) );
  OR U54950 ( .A(n42403), .B(n42402), .Z(n42404) );
  AND U54951 ( .A(n42405), .B(n42404), .Z(n42408) );
  NAND U54952 ( .A(n57080), .B(n42406), .Z(n42407) );
  OR U54953 ( .A(n42408), .B(n42407), .Z(n42409) );
  AND U54954 ( .A(n42410), .B(n42409), .Z(n42413) );
  NAND U54955 ( .A(n51556), .B(n42411), .Z(n42412) );
  OR U54956 ( .A(n42413), .B(n42412), .Z(n42414) );
  AND U54957 ( .A(n42415), .B(n42414), .Z(n42419) );
  NAND U54958 ( .A(n42417), .B(n42416), .Z(n42418) );
  OR U54959 ( .A(n42419), .B(n42418), .Z(n42420) );
  AND U54960 ( .A(n42421), .B(n42420), .Z(n42425) );
  NAND U54961 ( .A(n42423), .B(n42422), .Z(n42424) );
  OR U54962 ( .A(n42425), .B(n42424), .Z(n42426) );
  AND U54963 ( .A(n42427), .B(n42426), .Z(n42428) );
  OR U54964 ( .A(n42429), .B(n42428), .Z(n42430) );
  NAND U54965 ( .A(n42431), .B(n42430), .Z(n42432) );
  AND U54966 ( .A(n42433), .B(n42432), .Z(n42434) );
  ANDN U54967 ( .B(n42435), .A(n42434), .Z(n42436) );
  OR U54968 ( .A(n57094), .B(n42436), .Z(n42437) );
  NAND U54969 ( .A(n57095), .B(n42437), .Z(n42438) );
  NANDN U54970 ( .A(n42439), .B(n42438), .Z(n42440) );
  AND U54971 ( .A(n42440), .B(n51554), .Z(n42441) );
  NANDN U54972 ( .A(x[4808]), .B(y[4808]), .Z(n57096) );
  AND U54973 ( .A(n42441), .B(n57096), .Z(n42442) );
  NOR U54974 ( .A(n42443), .B(n42442), .Z(n42445) );
  NAND U54975 ( .A(n42445), .B(n42444), .Z(n42447) );
  NAND U54976 ( .A(n42447), .B(n42446), .Z(n42448) );
  ANDN U54977 ( .B(y[4810]), .A(x[4810]), .Z(n51552) );
  OR U54978 ( .A(n42448), .B(n51552), .Z(n42449) );
  NAND U54979 ( .A(n42450), .B(n42449), .Z(n42451) );
  AND U54980 ( .A(n42452), .B(n42451), .Z(n42453) );
  OR U54981 ( .A(n42454), .B(n42453), .Z(n42455) );
  NAND U54982 ( .A(n42456), .B(n42455), .Z(n42457) );
  NANDN U54983 ( .A(n42458), .B(n42457), .Z(n42460) );
  NANDN U54984 ( .A(n42460), .B(n42459), .Z(n42461) );
  AND U54985 ( .A(n42462), .B(n42461), .Z(n42463) );
  OR U54986 ( .A(n42464), .B(n42463), .Z(n42465) );
  NAND U54987 ( .A(n42466), .B(n42465), .Z(n42467) );
  NANDN U54988 ( .A(n42468), .B(n42467), .Z(n42470) );
  NANDN U54989 ( .A(n42470), .B(n42469), .Z(n42471) );
  NAND U54990 ( .A(n42472), .B(n42471), .Z(n42473) );
  AND U54991 ( .A(n42474), .B(n42473), .Z(n42475) );
  ANDN U54992 ( .B(n42476), .A(n42475), .Z(n42477) );
  NAND U54993 ( .A(n51549), .B(n42477), .Z(n42478) );
  NANDN U54994 ( .A(n42479), .B(n42478), .Z(n42480) );
  AND U54995 ( .A(n42481), .B(n42480), .Z(n42482) );
  OR U54996 ( .A(n42483), .B(n42482), .Z(n42484) );
  NAND U54997 ( .A(n42485), .B(n42484), .Z(n42486) );
  NANDN U54998 ( .A(n42487), .B(n42486), .Z(n42489) );
  AND U54999 ( .A(n42489), .B(n42488), .Z(n42490) );
  NANDN U55000 ( .A(x[4828]), .B(y[4828]), .Z(n51547) );
  AND U55001 ( .A(n42490), .B(n51547), .Z(n42491) );
  OR U55002 ( .A(n42492), .B(n42491), .Z(n42493) );
  NAND U55003 ( .A(n42494), .B(n42493), .Z(n42495) );
  NANDN U55004 ( .A(n42496), .B(n42495), .Z(n42498) );
  AND U55005 ( .A(n42498), .B(n42497), .Z(n42500) );
  NANDN U55006 ( .A(x[4832]), .B(y[4832]), .Z(n42499) );
  AND U55007 ( .A(n42500), .B(n42499), .Z(n42501) );
  OR U55008 ( .A(n42502), .B(n42501), .Z(n42503) );
  NAND U55009 ( .A(n42504), .B(n42503), .Z(n42505) );
  NANDN U55010 ( .A(n42506), .B(n42505), .Z(n42508) );
  AND U55011 ( .A(n42508), .B(n42507), .Z(n42509) );
  NANDN U55012 ( .A(x[4836]), .B(y[4836]), .Z(n57122) );
  AND U55013 ( .A(n42509), .B(n57122), .Z(n42510) );
  OR U55014 ( .A(n42511), .B(n42510), .Z(n42512) );
  NAND U55015 ( .A(n42513), .B(n42512), .Z(n42514) );
  NANDN U55016 ( .A(n42515), .B(n42514), .Z(n42517) );
  OR U55017 ( .A(n42517), .B(n42516), .Z(n42518) );
  AND U55018 ( .A(n42518), .B(n57130), .Z(n42519) );
  NANDN U55019 ( .A(x[4840]), .B(y[4840]), .Z(n57127) );
  NAND U55020 ( .A(n42519), .B(n57127), .Z(n42520) );
  AND U55021 ( .A(n42521), .B(n42520), .Z(n42523) );
  NANDN U55022 ( .A(x[4842]), .B(y[4842]), .Z(n57129) );
  AND U55023 ( .A(n57132), .B(n57129), .Z(n42522) );
  NANDN U55024 ( .A(n42523), .B(n42522), .Z(n42524) );
  NANDN U55025 ( .A(n42525), .B(n42524), .Z(n42527) );
  IV U55026 ( .A(n42526), .Z(n57135) );
  AND U55027 ( .A(n42527), .B(n57135), .Z(n42528) );
  NANDN U55028 ( .A(x[4844]), .B(y[4844]), .Z(n57133) );
  NAND U55029 ( .A(n42528), .B(n57133), .Z(n42529) );
  NAND U55030 ( .A(n42530), .B(n42529), .Z(n42533) );
  NANDN U55031 ( .A(x[4846]), .B(y[4846]), .Z(n57136) );
  AND U55032 ( .A(n42531), .B(n57136), .Z(n42532) );
  NAND U55033 ( .A(n42533), .B(n42532), .Z(n42534) );
  NANDN U55034 ( .A(n42535), .B(n42534), .Z(n42536) );
  NAND U55035 ( .A(n42537), .B(n42536), .Z(n42538) );
  AND U55036 ( .A(n42539), .B(n42538), .Z(n42540) );
  ANDN U55037 ( .B(n42541), .A(n42540), .Z(n42542) );
  NAND U55038 ( .A(n57142), .B(n42542), .Z(n42543) );
  NANDN U55039 ( .A(n42544), .B(n42543), .Z(n42545) );
  NAND U55040 ( .A(n42546), .B(n42545), .Z(n42547) );
  AND U55041 ( .A(n42548), .B(n42547), .Z(n42549) );
  ANDN U55042 ( .B(n57149), .A(n42549), .Z(n42550) );
  NAND U55043 ( .A(n51543), .B(n42550), .Z(n42551) );
  NANDN U55044 ( .A(n42552), .B(n42551), .Z(n42553) );
  AND U55045 ( .A(n42553), .B(n57152), .Z(n42554) );
  NANDN U55046 ( .A(x[4856]), .B(y[4856]), .Z(n57150) );
  NAND U55047 ( .A(n42554), .B(n57150), .Z(n42555) );
  NAND U55048 ( .A(n42556), .B(n42555), .Z(n42559) );
  NANDN U55049 ( .A(x[4858]), .B(y[4858]), .Z(n57153) );
  IV U55050 ( .A(n42557), .Z(n57155) );
  AND U55051 ( .A(n57153), .B(n57155), .Z(n42558) );
  NAND U55052 ( .A(n42559), .B(n42558), .Z(n42560) );
  NANDN U55053 ( .A(n42561), .B(n42560), .Z(n42562) );
  AND U55054 ( .A(n42562), .B(n51540), .Z(n42563) );
  NANDN U55055 ( .A(x[4860]), .B(y[4860]), .Z(n57156) );
  NAND U55056 ( .A(n42563), .B(n57156), .Z(n42564) );
  AND U55057 ( .A(n42565), .B(n42564), .Z(n42566) );
  ANDN U55058 ( .B(n57160), .A(n42566), .Z(n42567) );
  NAND U55059 ( .A(n51541), .B(n42567), .Z(n42568) );
  NANDN U55060 ( .A(n42569), .B(n42568), .Z(n42571) );
  IV U55061 ( .A(n42570), .Z(n57162) );
  AND U55062 ( .A(n42571), .B(n57162), .Z(n42572) );
  NANDN U55063 ( .A(x[4864]), .B(y[4864]), .Z(n57161) );
  NAND U55064 ( .A(n42572), .B(n57161), .Z(n42573) );
  AND U55065 ( .A(n42574), .B(n42573), .Z(n42575) );
  NOR U55066 ( .A(n57163), .B(n42575), .Z(n42576) );
  NAND U55067 ( .A(n57165), .B(n42576), .Z(n42577) );
  NANDN U55068 ( .A(n42578), .B(n42577), .Z(n42580) );
  NANDN U55069 ( .A(n42580), .B(n42579), .Z(n42581) );
  AND U55070 ( .A(n42581), .B(n51537), .Z(n42582) );
  NANDN U55071 ( .A(x[4868]), .B(y[4868]), .Z(n57166) );
  NAND U55072 ( .A(n42582), .B(n57166), .Z(n42583) );
  AND U55073 ( .A(n42584), .B(n42583), .Z(n42585) );
  ANDN U55074 ( .B(n57171), .A(n42585), .Z(n42586) );
  NAND U55075 ( .A(n51538), .B(n42586), .Z(n42587) );
  NANDN U55076 ( .A(n42588), .B(n42587), .Z(n42589) );
  AND U55077 ( .A(n42589), .B(n57175), .Z(n42590) );
  NANDN U55078 ( .A(x[4872]), .B(y[4872]), .Z(n57173) );
  NAND U55079 ( .A(n42590), .B(n57173), .Z(n42591) );
  AND U55080 ( .A(n42592), .B(n42591), .Z(n42593) );
  ANDN U55081 ( .B(n57178), .A(n42593), .Z(n42594) );
  NAND U55082 ( .A(n57176), .B(n42594), .Z(n42595) );
  NANDN U55083 ( .A(n42596), .B(n42595), .Z(n42598) );
  AND U55084 ( .A(n42598), .B(n42597), .Z(n42599) );
  NANDN U55085 ( .A(x[4876]), .B(y[4876]), .Z(n57179) );
  AND U55086 ( .A(n42599), .B(n57179), .Z(n42600) );
  OR U55087 ( .A(n42601), .B(n42600), .Z(n42602) );
  NAND U55088 ( .A(n42603), .B(n42602), .Z(n42604) );
  NANDN U55089 ( .A(n42605), .B(n42604), .Z(n42607) );
  AND U55090 ( .A(n42607), .B(n42606), .Z(n42609) );
  NANDN U55091 ( .A(x[4880]), .B(y[4880]), .Z(n42608) );
  AND U55092 ( .A(n42609), .B(n42608), .Z(n42610) );
  OR U55093 ( .A(n42611), .B(n42610), .Z(n42612) );
  NAND U55094 ( .A(n42613), .B(n42612), .Z(n42614) );
  NANDN U55095 ( .A(n42615), .B(n42614), .Z(n42616) );
  NAND U55096 ( .A(n42617), .B(n42616), .Z(n42618) );
  AND U55097 ( .A(n42619), .B(n42618), .Z(n42620) );
  ANDN U55098 ( .B(n42621), .A(n42620), .Z(n42622) );
  NAND U55099 ( .A(n57190), .B(n42622), .Z(n42623) );
  NANDN U55100 ( .A(n42624), .B(n42623), .Z(n42625) );
  AND U55101 ( .A(n42626), .B(n42625), .Z(n42627) );
  OR U55102 ( .A(n42628), .B(n42627), .Z(n42629) );
  NAND U55103 ( .A(n42630), .B(n42629), .Z(n42631) );
  NANDN U55104 ( .A(n42632), .B(n42631), .Z(n42634) );
  NANDN U55105 ( .A(n42634), .B(n42633), .Z(n42635) );
  AND U55106 ( .A(n42636), .B(n42635), .Z(n42637) );
  OR U55107 ( .A(n42638), .B(n42637), .Z(n42639) );
  NAND U55108 ( .A(n42640), .B(n42639), .Z(n42641) );
  NANDN U55109 ( .A(n42642), .B(n42641), .Z(n42644) );
  NANDN U55110 ( .A(n42644), .B(n42643), .Z(n42645) );
  AND U55111 ( .A(n42646), .B(n42645), .Z(n42647) );
  OR U55112 ( .A(n42648), .B(n42647), .Z(n42649) );
  NAND U55113 ( .A(n42650), .B(n42649), .Z(n42651) );
  NANDN U55114 ( .A(n42652), .B(n42651), .Z(n42654) );
  NANDN U55115 ( .A(n42654), .B(n42653), .Z(n42655) );
  AND U55116 ( .A(n42656), .B(n42655), .Z(n42657) );
  OR U55117 ( .A(n42658), .B(n42657), .Z(n42659) );
  NAND U55118 ( .A(n42660), .B(n42659), .Z(n42661) );
  NANDN U55119 ( .A(n42662), .B(n42661), .Z(n42664) );
  NANDN U55120 ( .A(n42664), .B(n42663), .Z(n42665) );
  AND U55121 ( .A(n42666), .B(n42665), .Z(n42667) );
  OR U55122 ( .A(n42668), .B(n42667), .Z(n42669) );
  NAND U55123 ( .A(n42670), .B(n42669), .Z(n42671) );
  NANDN U55124 ( .A(n42672), .B(n42671), .Z(n42673) );
  AND U55125 ( .A(n42674), .B(n42673), .Z(n42675) );
  OR U55126 ( .A(n42676), .B(n42675), .Z(n42677) );
  NAND U55127 ( .A(n42678), .B(n42677), .Z(n42679) );
  NANDN U55128 ( .A(n42680), .B(n42679), .Z(n42682) );
  NANDN U55129 ( .A(n42682), .B(n42681), .Z(n42683) );
  NAND U55130 ( .A(n42684), .B(n42683), .Z(n42685) );
  AND U55131 ( .A(n42686), .B(n42685), .Z(n42687) );
  ANDN U55132 ( .B(n57220), .A(n42687), .Z(n42688) );
  NAND U55133 ( .A(n57217), .B(n42688), .Z(n42689) );
  NANDN U55134 ( .A(n42690), .B(n42689), .Z(n42691) );
  AND U55135 ( .A(n42691), .B(n57223), .Z(n42692) );
  NANDN U55136 ( .A(x[4916]), .B(y[4916]), .Z(n57221) );
  NAND U55137 ( .A(n42692), .B(n57221), .Z(n42693) );
  AND U55138 ( .A(n42694), .B(n42693), .Z(n42695) );
  ANDN U55139 ( .B(n42696), .A(n42695), .Z(n42697) );
  NAND U55140 ( .A(n51530), .B(n42697), .Z(n42698) );
  NANDN U55141 ( .A(n42699), .B(n42698), .Z(n42700) );
  AND U55142 ( .A(n42701), .B(n42700), .Z(n42702) );
  OR U55143 ( .A(n42703), .B(n42702), .Z(n42704) );
  NAND U55144 ( .A(n42705), .B(n42704), .Z(n42706) );
  NANDN U55145 ( .A(n42707), .B(n42706), .Z(n42709) );
  NANDN U55146 ( .A(n42709), .B(n42708), .Z(n42711) );
  IV U55147 ( .A(n42710), .Z(n51525) );
  AND U55148 ( .A(n42711), .B(n51525), .Z(n42712) );
  NANDN U55149 ( .A(x[4924]), .B(y[4924]), .Z(n57229) );
  NAND U55150 ( .A(n42712), .B(n57229), .Z(n42713) );
  AND U55151 ( .A(n42714), .B(n42713), .Z(n42715) );
  ANDN U55152 ( .B(n57232), .A(n42715), .Z(n42716) );
  NAND U55153 ( .A(n51526), .B(n42716), .Z(n42717) );
  NANDN U55154 ( .A(n42718), .B(n42717), .Z(n42719) );
  AND U55155 ( .A(n42719), .B(n57235), .Z(n42720) );
  NANDN U55156 ( .A(n57233), .B(n42720), .Z(n42721) );
  NAND U55157 ( .A(n42722), .B(n42721), .Z(n42723) );
  NANDN U55158 ( .A(n42724), .B(n42723), .Z(n42725) );
  ANDN U55159 ( .B(y[4930]), .A(x[4930]), .Z(n57236) );
  OR U55160 ( .A(n42725), .B(n57236), .Z(n42726) );
  NAND U55161 ( .A(n42727), .B(n42726), .Z(n42728) );
  AND U55162 ( .A(n42729), .B(n42728), .Z(n42730) );
  OR U55163 ( .A(n42731), .B(n42730), .Z(n42732) );
  NAND U55164 ( .A(n42733), .B(n42732), .Z(n42734) );
  NANDN U55165 ( .A(n42735), .B(n42734), .Z(n42736) );
  AND U55166 ( .A(n42737), .B(n42736), .Z(n42738) );
  NANDN U55167 ( .A(x[4936]), .B(y[4936]), .Z(n51523) );
  AND U55168 ( .A(n42738), .B(n51523), .Z(n42739) );
  OR U55169 ( .A(n42740), .B(n42739), .Z(n42741) );
  NAND U55170 ( .A(n42742), .B(n42741), .Z(n42743) );
  NANDN U55171 ( .A(n42744), .B(n42743), .Z(n42746) );
  OR U55172 ( .A(n42746), .B(n42745), .Z(n42747) );
  NAND U55173 ( .A(n42748), .B(n42747), .Z(n42749) );
  NAND U55174 ( .A(n42750), .B(n42749), .Z(n42751) );
  AND U55175 ( .A(n42751), .B(n57254), .Z(n42752) );
  NANDN U55176 ( .A(x[4942]), .B(y[4942]), .Z(n57251) );
  AND U55177 ( .A(n42752), .B(n57251), .Z(n42756) );
  AND U55178 ( .A(n42754), .B(n42753), .Z(n42755) );
  NANDN U55179 ( .A(n42756), .B(n42755), .Z(n42757) );
  NAND U55180 ( .A(n42758), .B(n42757), .Z(n42759) );
  NAND U55181 ( .A(n42760), .B(n42759), .Z(n42761) );
  AND U55182 ( .A(n42761), .B(n57259), .Z(n42762) );
  NANDN U55183 ( .A(x[4946]), .B(y[4946]), .Z(n51522) );
  AND U55184 ( .A(n42762), .B(n51522), .Z(n42766) );
  AND U55185 ( .A(n42764), .B(n42763), .Z(n42765) );
  NANDN U55186 ( .A(n42766), .B(n42765), .Z(n42767) );
  NAND U55187 ( .A(n42768), .B(n42767), .Z(n42769) );
  AND U55188 ( .A(n42770), .B(n42769), .Z(n42771) );
  OR U55189 ( .A(n42772), .B(n42771), .Z(n42773) );
  NAND U55190 ( .A(n42774), .B(n42773), .Z(n42775) );
  NANDN U55191 ( .A(n42776), .B(n42775), .Z(n42777) );
  NAND U55192 ( .A(n42778), .B(n42777), .Z(n42780) );
  IV U55193 ( .A(n42779), .Z(n57269) );
  AND U55194 ( .A(n42780), .B(n57269), .Z(n42781) );
  ANDN U55195 ( .B(y[4954]), .A(x[4954]), .Z(n57265) );
  ANDN U55196 ( .B(n42781), .A(n57265), .Z(n42785) );
  AND U55197 ( .A(n42783), .B(n42782), .Z(n42784) );
  NANDN U55198 ( .A(n42785), .B(n42784), .Z(n42786) );
  NAND U55199 ( .A(n42787), .B(n42786), .Z(n42788) );
  AND U55200 ( .A(n42789), .B(n42788), .Z(n42790) );
  ANDN U55201 ( .B(n51517), .A(n42790), .Z(n42791) );
  NANDN U55202 ( .A(x[4958]), .B(y[4958]), .Z(n57273) );
  AND U55203 ( .A(n42791), .B(n57273), .Z(n42792) );
  OR U55204 ( .A(n42793), .B(n42792), .Z(n42794) );
  NAND U55205 ( .A(n42795), .B(n42794), .Z(n42796) );
  NAND U55206 ( .A(n42797), .B(n42796), .Z(n42799) );
  IV U55207 ( .A(n42798), .Z(n57277) );
  AND U55208 ( .A(n42799), .B(n57277), .Z(n42800) );
  NANDN U55209 ( .A(x[4962]), .B(y[4962]), .Z(n51515) );
  AND U55210 ( .A(n42800), .B(n51515), .Z(n42804) );
  AND U55211 ( .A(n42802), .B(n42801), .Z(n42803) );
  NANDN U55212 ( .A(n42804), .B(n42803), .Z(n42805) );
  NAND U55213 ( .A(n42806), .B(n42805), .Z(n42807) );
  NAND U55214 ( .A(n42808), .B(n42807), .Z(n42810) );
  AND U55215 ( .A(n42810), .B(n42809), .Z(n42811) );
  NANDN U55216 ( .A(n57281), .B(n42811), .Z(n42812) );
  NAND U55217 ( .A(n42813), .B(n42812), .Z(n42814) );
  NANDN U55218 ( .A(n42815), .B(n42814), .Z(n42816) );
  AND U55219 ( .A(n42817), .B(n42816), .Z(n42818) );
  OR U55220 ( .A(n42819), .B(n42818), .Z(n42820) );
  NAND U55221 ( .A(n42821), .B(n42820), .Z(n42822) );
  NANDN U55222 ( .A(n42823), .B(n42822), .Z(n42824) );
  AND U55223 ( .A(n42825), .B(n42824), .Z(n42826) );
  OR U55224 ( .A(n42827), .B(n42826), .Z(n42828) );
  NAND U55225 ( .A(n42829), .B(n42828), .Z(n42830) );
  NANDN U55226 ( .A(n42831), .B(n42830), .Z(n42832) );
  NAND U55227 ( .A(n42833), .B(n42832), .Z(n42834) );
  AND U55228 ( .A(n42834), .B(n51511), .Z(n42836) );
  NANDN U55229 ( .A(x[4978]), .B(y[4978]), .Z(n42835) );
  AND U55230 ( .A(n42836), .B(n42835), .Z(n42840) );
  AND U55231 ( .A(n42838), .B(n42837), .Z(n42839) );
  NANDN U55232 ( .A(n42840), .B(n42839), .Z(n42841) );
  NAND U55233 ( .A(n42842), .B(n42841), .Z(n42843) );
  NAND U55234 ( .A(n42844), .B(n42843), .Z(n42845) );
  AND U55235 ( .A(n42845), .B(n57303), .Z(n42846) );
  NANDN U55236 ( .A(x[4982]), .B(y[4982]), .Z(n57301) );
  AND U55237 ( .A(n42846), .B(n57301), .Z(n42850) );
  AND U55238 ( .A(n42848), .B(n42847), .Z(n42849) );
  NANDN U55239 ( .A(n42850), .B(n42849), .Z(n42851) );
  NAND U55240 ( .A(n42852), .B(n42851), .Z(n42853) );
  NAND U55241 ( .A(n42854), .B(n42853), .Z(n42855) );
  AND U55242 ( .A(n42855), .B(n57310), .Z(n42856) );
  NANDN U55243 ( .A(x[4986]), .B(y[4986]), .Z(n57307) );
  AND U55244 ( .A(n42856), .B(n57307), .Z(n42860) );
  AND U55245 ( .A(n42858), .B(n42857), .Z(n42859) );
  NANDN U55246 ( .A(n42860), .B(n42859), .Z(n42861) );
  NAND U55247 ( .A(n42862), .B(n42861), .Z(n42863) );
  NAND U55248 ( .A(n42864), .B(n42863), .Z(n42866) );
  IV U55249 ( .A(n42865), .Z(n57314) );
  AND U55250 ( .A(n42866), .B(n57314), .Z(n42867) );
  NANDN U55251 ( .A(x[4990]), .B(y[4990]), .Z(n57312) );
  AND U55252 ( .A(n42867), .B(n57312), .Z(n42871) );
  AND U55253 ( .A(n42869), .B(n42868), .Z(n42870) );
  NANDN U55254 ( .A(n42871), .B(n42870), .Z(n42872) );
  NAND U55255 ( .A(n42873), .B(n42872), .Z(n42874) );
  AND U55256 ( .A(n42875), .B(n42874), .Z(n42879) );
  IV U55257 ( .A(n42876), .Z(n57320) );
  AND U55258 ( .A(n42877), .B(n57320), .Z(n42878) );
  NANDN U55259 ( .A(n42879), .B(n42878), .Z(n42880) );
  NAND U55260 ( .A(n42881), .B(n42880), .Z(n42883) );
  OR U55261 ( .A(n42883), .B(n42882), .Z(n42884) );
  NAND U55262 ( .A(n42885), .B(n42884), .Z(n42886) );
  AND U55263 ( .A(n42887), .B(n42886), .Z(n42888) );
  ANDN U55264 ( .B(n42889), .A(n42888), .Z(n42890) );
  NAND U55265 ( .A(n57324), .B(n42890), .Z(n42891) );
  NANDN U55266 ( .A(n42892), .B(n42891), .Z(n42893) );
  NAND U55267 ( .A(n42894), .B(n42893), .Z(n42895) );
  NAND U55268 ( .A(n42896), .B(n42895), .Z(n42898) );
  IV U55269 ( .A(n42897), .Z(n57330) );
  AND U55270 ( .A(n42898), .B(n57330), .Z(n42899) );
  NANDN U55271 ( .A(x[5002]), .B(y[5002]), .Z(n57328) );
  AND U55272 ( .A(n42899), .B(n57328), .Z(n42903) );
  AND U55273 ( .A(n42901), .B(n42900), .Z(n42902) );
  NANDN U55274 ( .A(n42903), .B(n42902), .Z(n42904) );
  NAND U55275 ( .A(n42905), .B(n42904), .Z(n42906) );
  NAND U55276 ( .A(n42907), .B(n42906), .Z(n42908) );
  AND U55277 ( .A(n42909), .B(n42908), .Z(n42913) );
  AND U55278 ( .A(n42911), .B(n42910), .Z(n42912) );
  NANDN U55279 ( .A(n42913), .B(n42912), .Z(n42914) );
  NAND U55280 ( .A(n42915), .B(n42914), .Z(n42916) );
  AND U55281 ( .A(n42917), .B(n42916), .Z(n42918) );
  OR U55282 ( .A(n42919), .B(n42918), .Z(n42920) );
  NAND U55283 ( .A(n42921), .B(n42920), .Z(n42922) );
  NANDN U55284 ( .A(n42923), .B(n42922), .Z(n42924) );
  NAND U55285 ( .A(n42925), .B(n42924), .Z(n42926) );
  AND U55286 ( .A(n42927), .B(n42926), .Z(n42931) );
  AND U55287 ( .A(n42929), .B(n42928), .Z(n42930) );
  NANDN U55288 ( .A(n42931), .B(n42930), .Z(n42932) );
  NAND U55289 ( .A(n42933), .B(n42932), .Z(n42934) );
  NAND U55290 ( .A(n42935), .B(n42934), .Z(n42937) );
  AND U55291 ( .A(n42937), .B(n42936), .Z(n42938) );
  NANDN U55292 ( .A(n57351), .B(n42938), .Z(n42939) );
  NAND U55293 ( .A(n42940), .B(n42939), .Z(n42941) );
  NANDN U55294 ( .A(n42942), .B(n42941), .Z(n42943) );
  AND U55295 ( .A(n42944), .B(n42943), .Z(n42946) );
  NANDN U55296 ( .A(x[5022]), .B(y[5022]), .Z(n57353) );
  AND U55297 ( .A(n57356), .B(n57353), .Z(n42945) );
  NANDN U55298 ( .A(n42946), .B(n42945), .Z(n42947) );
  NAND U55299 ( .A(n42948), .B(n42947), .Z(n42949) );
  ANDN U55300 ( .B(y[5024]), .A(x[5024]), .Z(n57357) );
  ANDN U55301 ( .B(n42949), .A(n57357), .Z(n42950) );
  NANDN U55302 ( .A(n42951), .B(n42950), .Z(n42952) );
  NAND U55303 ( .A(n42953), .B(n42952), .Z(n42954) );
  AND U55304 ( .A(n42954), .B(n57360), .Z(n42956) );
  NANDN U55305 ( .A(x[5026]), .B(y[5026]), .Z(n42955) );
  AND U55306 ( .A(n42956), .B(n42955), .Z(n42960) );
  AND U55307 ( .A(n42958), .B(n42957), .Z(n42959) );
  NANDN U55308 ( .A(n42960), .B(n42959), .Z(n42961) );
  NAND U55309 ( .A(n42962), .B(n42961), .Z(n42963) );
  AND U55310 ( .A(n42964), .B(n42963), .Z(n42965) );
  OR U55311 ( .A(n42966), .B(n42965), .Z(n42967) );
  NAND U55312 ( .A(n42968), .B(n42967), .Z(n42969) );
  NANDN U55313 ( .A(n42970), .B(n42969), .Z(n42971) );
  AND U55314 ( .A(n42972), .B(n42971), .Z(n42973) );
  OR U55315 ( .A(n42974), .B(n42973), .Z(n42975) );
  NAND U55316 ( .A(n42976), .B(n42975), .Z(n42978) );
  ANDN U55317 ( .B(n42978), .A(n42977), .Z(n42979) );
  NAND U55318 ( .A(n42979), .B(n51501), .Z(n42980) );
  AND U55319 ( .A(n42981), .B(n42980), .Z(n42982) );
  OR U55320 ( .A(n42983), .B(n42982), .Z(n42984) );
  NAND U55321 ( .A(n42985), .B(n42984), .Z(n42986) );
  NANDN U55322 ( .A(n42987), .B(n42986), .Z(n42988) );
  NAND U55323 ( .A(n42989), .B(n42988), .Z(n42991) );
  AND U55324 ( .A(n42991), .B(n42990), .Z(n42992) );
  NANDN U55325 ( .A(n57378), .B(n42992), .Z(n42993) );
  NAND U55326 ( .A(n42994), .B(n42993), .Z(n42995) );
  NANDN U55327 ( .A(n42996), .B(n42995), .Z(n42997) );
  AND U55328 ( .A(n42998), .B(n42997), .Z(n42999) );
  OR U55329 ( .A(n43000), .B(n42999), .Z(n43001) );
  NAND U55330 ( .A(n43002), .B(n43001), .Z(n43003) );
  NANDN U55331 ( .A(n43004), .B(n43003), .Z(n43005) );
  NAND U55332 ( .A(n43006), .B(n43005), .Z(n43007) );
  AND U55333 ( .A(n43007), .B(n57387), .Z(n43008) );
  NANDN U55334 ( .A(x[5050]), .B(y[5050]), .Z(n51498) );
  AND U55335 ( .A(n43008), .B(n51498), .Z(n43012) );
  AND U55336 ( .A(n43010), .B(n43009), .Z(n43011) );
  NANDN U55337 ( .A(n43012), .B(n43011), .Z(n43013) );
  NAND U55338 ( .A(n43014), .B(n43013), .Z(n43015) );
  AND U55339 ( .A(n43016), .B(n43015), .Z(n43017) );
  OR U55340 ( .A(n43018), .B(n43017), .Z(n43019) );
  NAND U55341 ( .A(n43020), .B(n43019), .Z(n43021) );
  NANDN U55342 ( .A(n43022), .B(n43021), .Z(n43023) );
  NAND U55343 ( .A(n43024), .B(n43023), .Z(n43025) );
  AND U55344 ( .A(n43026), .B(n43025), .Z(n43030) );
  AND U55345 ( .A(n43028), .B(n43027), .Z(n43029) );
  NANDN U55346 ( .A(n43030), .B(n43029), .Z(n43031) );
  NAND U55347 ( .A(n43032), .B(n43031), .Z(n43033) );
  NAND U55348 ( .A(n43034), .B(n43033), .Z(n43035) );
  AND U55349 ( .A(n43035), .B(n57403), .Z(n43036) );
  NANDN U55350 ( .A(x[5062]), .B(y[5062]), .Z(n51495) );
  AND U55351 ( .A(n43036), .B(n51495), .Z(n43040) );
  AND U55352 ( .A(n43038), .B(n43037), .Z(n43039) );
  NANDN U55353 ( .A(n43040), .B(n43039), .Z(n43041) );
  NAND U55354 ( .A(n43042), .B(n43041), .Z(n43043) );
  NAND U55355 ( .A(n43044), .B(n43043), .Z(n43045) );
  AND U55356 ( .A(n43045), .B(n57409), .Z(n43046) );
  NANDN U55357 ( .A(x[5066]), .B(y[5066]), .Z(n57406) );
  AND U55358 ( .A(n43046), .B(n57406), .Z(n43050) );
  AND U55359 ( .A(n43048), .B(n43047), .Z(n43049) );
  NANDN U55360 ( .A(n43050), .B(n43049), .Z(n43051) );
  NAND U55361 ( .A(n43052), .B(n43051), .Z(n43053) );
  AND U55362 ( .A(n43054), .B(n43053), .Z(n43055) );
  OR U55363 ( .A(n43056), .B(n43055), .Z(n43057) );
  NAND U55364 ( .A(n43058), .B(n43057), .Z(n43059) );
  NANDN U55365 ( .A(n43060), .B(n43059), .Z(n43061) );
  NAND U55366 ( .A(n43062), .B(n43061), .Z(n43063) );
  AND U55367 ( .A(n43064), .B(n43063), .Z(n43068) );
  AND U55368 ( .A(n43066), .B(n43065), .Z(n43067) );
  NANDN U55369 ( .A(n43068), .B(n43067), .Z(n43069) );
  NAND U55370 ( .A(n43070), .B(n43069), .Z(n43071) );
  NAND U55371 ( .A(n43072), .B(n43071), .Z(n43073) );
  AND U55372 ( .A(n43074), .B(n43073), .Z(n43078) );
  AND U55373 ( .A(n43076), .B(n43075), .Z(n43077) );
  NANDN U55374 ( .A(n43078), .B(n43077), .Z(n43079) );
  NAND U55375 ( .A(n43080), .B(n43079), .Z(n43081) );
  NAND U55376 ( .A(n43082), .B(n43081), .Z(n43083) );
  AND U55377 ( .A(n43083), .B(n57427), .Z(n43084) );
  NANDN U55378 ( .A(x[5082]), .B(y[5082]), .Z(n51491) );
  AND U55379 ( .A(n43084), .B(n51491), .Z(n43088) );
  AND U55380 ( .A(n43086), .B(n43085), .Z(n43087) );
  NANDN U55381 ( .A(n43088), .B(n43087), .Z(n43089) );
  NAND U55382 ( .A(n43090), .B(n43089), .Z(n43091) );
  AND U55383 ( .A(n43092), .B(n43091), .Z(n43093) );
  OR U55384 ( .A(n43094), .B(n43093), .Z(n43095) );
  NAND U55385 ( .A(n43096), .B(n43095), .Z(n43097) );
  NANDN U55386 ( .A(n43098), .B(n43097), .Z(n43099) );
  AND U55387 ( .A(n43100), .B(n43099), .Z(n43101) );
  OR U55388 ( .A(n43102), .B(n43101), .Z(n43103) );
  NAND U55389 ( .A(n43104), .B(n43103), .Z(n43105) );
  NANDN U55390 ( .A(n43106), .B(n43105), .Z(n43107) );
  NAND U55391 ( .A(n43108), .B(n43107), .Z(n43110) );
  IV U55392 ( .A(n43109), .Z(n51488) );
  AND U55393 ( .A(n43110), .B(n51488), .Z(n43111) );
  NANDN U55394 ( .A(x[5094]), .B(y[5094]), .Z(n57442) );
  AND U55395 ( .A(n43111), .B(n57442), .Z(n43115) );
  AND U55396 ( .A(n43113), .B(n43112), .Z(n43114) );
  NANDN U55397 ( .A(n43115), .B(n43114), .Z(n43116) );
  NAND U55398 ( .A(n43117), .B(n43116), .Z(n43118) );
  AND U55399 ( .A(n43119), .B(n43118), .Z(n43123) );
  AND U55400 ( .A(n43121), .B(n43120), .Z(n43122) );
  NANDN U55401 ( .A(n43123), .B(n43122), .Z(n43124) );
  NANDN U55402 ( .A(n43125), .B(n43124), .Z(n43126) );
  AND U55403 ( .A(n43127), .B(n43126), .Z(n43129) );
  NAND U55404 ( .A(n43129), .B(n43128), .Z(n43130) );
  AND U55405 ( .A(n43131), .B(n43130), .Z(n43132) );
  OR U55406 ( .A(n43133), .B(n43132), .Z(n43134) );
  NAND U55407 ( .A(n43135), .B(n43134), .Z(n43136) );
  NANDN U55408 ( .A(n43137), .B(n43136), .Z(n43138) );
  NAND U55409 ( .A(n43139), .B(n43138), .Z(n43140) );
  AND U55410 ( .A(n43140), .B(n51486), .Z(n43141) );
  NANDN U55411 ( .A(x[5106]), .B(y[5106]), .Z(n57455) );
  AND U55412 ( .A(n43141), .B(n57455), .Z(n43142) );
  OR U55413 ( .A(n43143), .B(n43142), .Z(n43144) );
  NAND U55414 ( .A(n43145), .B(n43144), .Z(n43146) );
  NAND U55415 ( .A(n43147), .B(n43146), .Z(n43149) );
  IV U55416 ( .A(n43148), .Z(n57459) );
  AND U55417 ( .A(n43149), .B(n57459), .Z(n43150) );
  NANDN U55418 ( .A(x[5110]), .B(y[5110]), .Z(n51485) );
  AND U55419 ( .A(n43150), .B(n51485), .Z(n43154) );
  AND U55420 ( .A(n43152), .B(n43151), .Z(n43153) );
  NANDN U55421 ( .A(n43154), .B(n43153), .Z(n43155) );
  NAND U55422 ( .A(n43156), .B(n43155), .Z(n43157) );
  AND U55423 ( .A(n43158), .B(n43157), .Z(n43159) );
  ANDN U55424 ( .B(n51482), .A(n43159), .Z(n43160) );
  NANDN U55425 ( .A(x[5114]), .B(y[5114]), .Z(n57463) );
  AND U55426 ( .A(n43160), .B(n57463), .Z(n43161) );
  OR U55427 ( .A(n43162), .B(n43161), .Z(n43163) );
  NAND U55428 ( .A(n43164), .B(n43163), .Z(n43165) );
  AND U55429 ( .A(n43166), .B(n43165), .Z(n43167) );
  OR U55430 ( .A(n43168), .B(n43167), .Z(n43169) );
  NAND U55431 ( .A(n43170), .B(n43169), .Z(n43171) );
  NANDN U55432 ( .A(n43172), .B(n43171), .Z(n43173) );
  AND U55433 ( .A(n43174), .B(n43173), .Z(n43175) );
  OR U55434 ( .A(n43176), .B(n43175), .Z(n43177) );
  NAND U55435 ( .A(n43178), .B(n43177), .Z(n43179) );
  NANDN U55436 ( .A(n43180), .B(n43179), .Z(n43181) );
  NAND U55437 ( .A(n43182), .B(n43181), .Z(n43183) );
  AND U55438 ( .A(n43183), .B(n51480), .Z(n43185) );
  NANDN U55439 ( .A(x[5126]), .B(y[5126]), .Z(n43184) );
  AND U55440 ( .A(n43185), .B(n43184), .Z(n43189) );
  AND U55441 ( .A(n43187), .B(n43186), .Z(n43188) );
  NANDN U55442 ( .A(n43189), .B(n43188), .Z(n43190) );
  NAND U55443 ( .A(n43191), .B(n43190), .Z(n43192) );
  NAND U55444 ( .A(n43193), .B(n43192), .Z(n43195) );
  IV U55445 ( .A(n43194), .Z(n57484) );
  AND U55446 ( .A(n43195), .B(n57484), .Z(n43196) );
  NANDN U55447 ( .A(x[5130]), .B(y[5130]), .Z(n57480) );
  AND U55448 ( .A(n43196), .B(n57480), .Z(n43200) );
  AND U55449 ( .A(n43198), .B(n43197), .Z(n43199) );
  NANDN U55450 ( .A(n43200), .B(n43199), .Z(n43201) );
  NAND U55451 ( .A(n43202), .B(n43201), .Z(n43203) );
  NAND U55452 ( .A(n43204), .B(n43203), .Z(n43206) );
  IV U55453 ( .A(n43205), .Z(n51477) );
  AND U55454 ( .A(n43206), .B(n51477), .Z(n43207) );
  NANDN U55455 ( .A(x[5134]), .B(y[5134]), .Z(n57488) );
  AND U55456 ( .A(n43207), .B(n57488), .Z(n43211) );
  AND U55457 ( .A(n43209), .B(n43208), .Z(n43210) );
  NANDN U55458 ( .A(n43211), .B(n43210), .Z(n43212) );
  NAND U55459 ( .A(n43213), .B(n43212), .Z(n43214) );
  AND U55460 ( .A(n43215), .B(n43214), .Z(n43216) );
  OR U55461 ( .A(n43217), .B(n43216), .Z(n43218) );
  NAND U55462 ( .A(n43219), .B(n43218), .Z(n43220) );
  NANDN U55463 ( .A(n43221), .B(n43220), .Z(n43222) );
  AND U55464 ( .A(n43223), .B(n43222), .Z(n43224) );
  OR U55465 ( .A(n43225), .B(n43224), .Z(n43226) );
  NAND U55466 ( .A(n43227), .B(n43226), .Z(n43228) );
  NANDN U55467 ( .A(n43229), .B(n43228), .Z(n43230) );
  NAND U55468 ( .A(n43231), .B(n43230), .Z(n43233) );
  IV U55469 ( .A(n43232), .Z(n51473) );
  AND U55470 ( .A(n43233), .B(n51473), .Z(n43234) );
  NANDN U55471 ( .A(x[5146]), .B(y[5146]), .Z(n57501) );
  AND U55472 ( .A(n43234), .B(n57501), .Z(n43238) );
  AND U55473 ( .A(n43236), .B(n43235), .Z(n43237) );
  NANDN U55474 ( .A(n43238), .B(n43237), .Z(n43239) );
  NAND U55475 ( .A(n43240), .B(n43239), .Z(n43241) );
  AND U55476 ( .A(n43242), .B(n43241), .Z(n43245) );
  AND U55477 ( .A(n43243), .B(n57505), .Z(n43244) );
  NANDN U55478 ( .A(n43245), .B(n43244), .Z(n43246) );
  NAND U55479 ( .A(n43247), .B(n43246), .Z(n43248) );
  OR U55480 ( .A(n43249), .B(n43248), .Z(n43250) );
  AND U55481 ( .A(n43251), .B(n43250), .Z(n43252) );
  OR U55482 ( .A(n43253), .B(n43252), .Z(n43254) );
  NAND U55483 ( .A(n43255), .B(n43254), .Z(n43256) );
  NANDN U55484 ( .A(n43257), .B(n43256), .Z(n43258) );
  AND U55485 ( .A(n43258), .B(n57513), .Z(n43259) );
  NANDN U55486 ( .A(x[5156]), .B(y[5156]), .Z(n57511) );
  NAND U55487 ( .A(n43259), .B(n57511), .Z(n43260) );
  AND U55488 ( .A(n43261), .B(n43260), .Z(n43264) );
  NANDN U55489 ( .A(x[5158]), .B(y[5158]), .Z(n57514) );
  AND U55490 ( .A(n57514), .B(n43262), .Z(n43263) );
  NANDN U55491 ( .A(n43264), .B(n43263), .Z(n43265) );
  NANDN U55492 ( .A(n43266), .B(n43265), .Z(n43267) );
  AND U55493 ( .A(n43268), .B(n43267), .Z(n43270) );
  NAND U55494 ( .A(n43270), .B(n43269), .Z(n43271) );
  AND U55495 ( .A(n43272), .B(n43271), .Z(n43273) );
  OR U55496 ( .A(n43274), .B(n43273), .Z(n43275) );
  NAND U55497 ( .A(n43276), .B(n43275), .Z(n43277) );
  NANDN U55498 ( .A(n43278), .B(n43277), .Z(n43279) );
  NAND U55499 ( .A(n43280), .B(n43279), .Z(n43282) );
  AND U55500 ( .A(n43282), .B(n43281), .Z(n43283) );
  NAND U55501 ( .A(n51469), .B(n43283), .Z(n43284) );
  NAND U55502 ( .A(n43285), .B(n43284), .Z(n43286) );
  NANDN U55503 ( .A(n43287), .B(n43286), .Z(n43288) );
  NAND U55504 ( .A(n43289), .B(n43288), .Z(n43290) );
  AND U55505 ( .A(n43290), .B(n51466), .Z(n43291) );
  NANDN U55506 ( .A(x[5170]), .B(y[5170]), .Z(n57528) );
  AND U55507 ( .A(n43291), .B(n57528), .Z(n43295) );
  AND U55508 ( .A(n43293), .B(n43292), .Z(n43294) );
  NANDN U55509 ( .A(n43295), .B(n43294), .Z(n43296) );
  NAND U55510 ( .A(n43297), .B(n43296), .Z(n43298) );
  NAND U55511 ( .A(n43299), .B(n43298), .Z(n43301) );
  IV U55512 ( .A(n43300), .Z(n57534) );
  AND U55513 ( .A(n43301), .B(n57534), .Z(n43302) );
  NANDN U55514 ( .A(x[5174]), .B(y[5174]), .Z(n57531) );
  AND U55515 ( .A(n43302), .B(n57531), .Z(n43306) );
  AND U55516 ( .A(n43304), .B(n43303), .Z(n43305) );
  NANDN U55517 ( .A(n43306), .B(n43305), .Z(n43307) );
  NAND U55518 ( .A(n43308), .B(n43307), .Z(n43309) );
  NAND U55519 ( .A(n43310), .B(n43309), .Z(n43311) );
  AND U55520 ( .A(n43312), .B(n43311), .Z(n43316) );
  AND U55521 ( .A(n43314), .B(n43313), .Z(n43315) );
  NANDN U55522 ( .A(n43316), .B(n43315), .Z(n43317) );
  NAND U55523 ( .A(n43318), .B(n43317), .Z(n43319) );
  AND U55524 ( .A(n43320), .B(n43319), .Z(n43321) );
  NOR U55525 ( .A(n57544), .B(n43321), .Z(n43322) );
  NAND U55526 ( .A(n57546), .B(n43322), .Z(n43323) );
  NANDN U55527 ( .A(n43324), .B(n43323), .Z(n43325) );
  OR U55528 ( .A(n43326), .B(n43325), .Z(n43327) );
  NAND U55529 ( .A(n43328), .B(n43327), .Z(n43329) );
  NAND U55530 ( .A(n43330), .B(n43329), .Z(n43331) );
  AND U55531 ( .A(n43332), .B(n43331), .Z(n43336) );
  AND U55532 ( .A(n43334), .B(n43333), .Z(n43335) );
  NANDN U55533 ( .A(n43336), .B(n43335), .Z(n43337) );
  NAND U55534 ( .A(n43338), .B(n43337), .Z(n43339) );
  AND U55535 ( .A(n43340), .B(n43339), .Z(n43341) );
  OR U55536 ( .A(n43342), .B(n43341), .Z(n43343) );
  NAND U55537 ( .A(n43344), .B(n43343), .Z(n43345) );
  AND U55538 ( .A(n57557), .B(n43345), .Z(n43346) );
  NAND U55539 ( .A(n51461), .B(n43346), .Z(n43347) );
  NAND U55540 ( .A(n43348), .B(n43347), .Z(n43350) );
  IV U55541 ( .A(n43349), .Z(n57558) );
  AND U55542 ( .A(n43350), .B(n57558), .Z(n43351) );
  NANDN U55543 ( .A(x[5194]), .B(y[5194]), .Z(n57556) );
  AND U55544 ( .A(n43351), .B(n57556), .Z(n43355) );
  AND U55545 ( .A(n43353), .B(n43352), .Z(n43354) );
  NANDN U55546 ( .A(n43355), .B(n43354), .Z(n43356) );
  NAND U55547 ( .A(n43357), .B(n43356), .Z(n43358) );
  NAND U55548 ( .A(n43359), .B(n43358), .Z(n43361) );
  IV U55549 ( .A(n43360), .Z(n51457) );
  AND U55550 ( .A(n43361), .B(n51457), .Z(n43362) );
  NANDN U55551 ( .A(x[5198]), .B(y[5198]), .Z(n57562) );
  AND U55552 ( .A(n43362), .B(n57562), .Z(n43366) );
  AND U55553 ( .A(n43364), .B(n43363), .Z(n43365) );
  NANDN U55554 ( .A(n43366), .B(n43365), .Z(n43367) );
  NAND U55555 ( .A(n43368), .B(n43367), .Z(n43369) );
  AND U55556 ( .A(n43370), .B(n43369), .Z(n43371) );
  OR U55557 ( .A(n43372), .B(n43371), .Z(n43373) );
  NAND U55558 ( .A(n43374), .B(n43373), .Z(n43375) );
  NANDN U55559 ( .A(n43376), .B(n43375), .Z(n43377) );
  NAND U55560 ( .A(n43378), .B(n43377), .Z(n43379) );
  AND U55561 ( .A(n43380), .B(n43379), .Z(n43384) );
  AND U55562 ( .A(n43382), .B(n43381), .Z(n43383) );
  NANDN U55563 ( .A(n43384), .B(n43383), .Z(n43385) );
  NAND U55564 ( .A(n43386), .B(n43385), .Z(n43387) );
  NAND U55565 ( .A(n43388), .B(n43387), .Z(n43389) );
  AND U55566 ( .A(n43389), .B(n51450), .Z(n43390) );
  NANDN U55567 ( .A(x[5210]), .B(y[5210]), .Z(n57575) );
  AND U55568 ( .A(n43390), .B(n57575), .Z(n43394) );
  AND U55569 ( .A(n43392), .B(n43391), .Z(n43393) );
  NANDN U55570 ( .A(n43394), .B(n43393), .Z(n43395) );
  NAND U55571 ( .A(n43396), .B(n43395), .Z(n43397) );
  AND U55572 ( .A(n43398), .B(n43397), .Z(n43399) );
  OR U55573 ( .A(n43400), .B(n43399), .Z(n43401) );
  NAND U55574 ( .A(n43402), .B(n43401), .Z(n43403) );
  NANDN U55575 ( .A(n43404), .B(n43403), .Z(n43405) );
  NAND U55576 ( .A(n43406), .B(n43405), .Z(n43407) );
  AND U55577 ( .A(n43407), .B(n57586), .Z(n43409) );
  NANDN U55578 ( .A(x[5218]), .B(y[5218]), .Z(n43408) );
  AND U55579 ( .A(n43409), .B(n43408), .Z(n43413) );
  AND U55580 ( .A(n43411), .B(n43410), .Z(n43412) );
  NANDN U55581 ( .A(n43413), .B(n43412), .Z(n43414) );
  NAND U55582 ( .A(n43415), .B(n43414), .Z(n43416) );
  NAND U55583 ( .A(n43417), .B(n43416), .Z(n43418) );
  AND U55584 ( .A(n43418), .B(n51444), .Z(n43420) );
  NANDN U55585 ( .A(x[5222]), .B(y[5222]), .Z(n43419) );
  AND U55586 ( .A(n43420), .B(n43419), .Z(n43424) );
  AND U55587 ( .A(n43422), .B(n43421), .Z(n43423) );
  NANDN U55588 ( .A(n43424), .B(n43423), .Z(n43425) );
  NAND U55589 ( .A(n43426), .B(n43425), .Z(n43427) );
  AND U55590 ( .A(n43428), .B(n43427), .Z(n43429) );
  OR U55591 ( .A(n43430), .B(n43429), .Z(n43431) );
  NAND U55592 ( .A(n43432), .B(n43431), .Z(n43433) );
  NANDN U55593 ( .A(n43434), .B(n43433), .Z(n43435) );
  NAND U55594 ( .A(n43436), .B(n43435), .Z(n43437) );
  AND U55595 ( .A(n43437), .B(n57598), .Z(n43438) );
  NANDN U55596 ( .A(x[5230]), .B(y[5230]), .Z(n51442) );
  AND U55597 ( .A(n43438), .B(n51442), .Z(n43442) );
  AND U55598 ( .A(n43440), .B(n43439), .Z(n43441) );
  NANDN U55599 ( .A(n43442), .B(n43441), .Z(n43443) );
  NAND U55600 ( .A(n43444), .B(n43443), .Z(n43445) );
  NAND U55601 ( .A(n43446), .B(n43445), .Z(n43447) );
  AND U55602 ( .A(n43448), .B(n43447), .Z(n43452) );
  AND U55603 ( .A(n43450), .B(n43449), .Z(n43451) );
  NANDN U55604 ( .A(n43452), .B(n43451), .Z(n43453) );
  NAND U55605 ( .A(n43454), .B(n43453), .Z(n43455) );
  NAND U55606 ( .A(n43456), .B(n43455), .Z(n43457) );
  AND U55607 ( .A(n43457), .B(n57608), .Z(n43458) );
  NANDN U55608 ( .A(x[5238]), .B(y[5238]), .Z(n57605) );
  AND U55609 ( .A(n43458), .B(n57605), .Z(n43462) );
  AND U55610 ( .A(n43460), .B(n43459), .Z(n43461) );
  NANDN U55611 ( .A(n43462), .B(n43461), .Z(n43463) );
  NAND U55612 ( .A(n43464), .B(n43463), .Z(n43465) );
  AND U55613 ( .A(n43466), .B(n43465), .Z(n43467) );
  OR U55614 ( .A(n43468), .B(n43467), .Z(n43469) );
  NAND U55615 ( .A(n43470), .B(n43469), .Z(n43471) );
  NANDN U55616 ( .A(n43472), .B(n43471), .Z(n43473) );
  AND U55617 ( .A(n43474), .B(n43473), .Z(n43477) );
  NANDN U55618 ( .A(x[5246]), .B(y[5246]), .Z(n57617) );
  IV U55619 ( .A(n43475), .Z(n57620) );
  AND U55620 ( .A(n57617), .B(n57620), .Z(n43476) );
  NANDN U55621 ( .A(n43477), .B(n43476), .Z(n43478) );
  NANDN U55622 ( .A(n43479), .B(n43478), .Z(n43480) );
  NANDN U55623 ( .A(x[5248]), .B(y[5248]), .Z(n51440) );
  AND U55624 ( .A(n43480), .B(n51440), .Z(n43482) );
  NAND U55625 ( .A(n43482), .B(n43481), .Z(n43483) );
  AND U55626 ( .A(n43484), .B(n43483), .Z(n43485) );
  OR U55627 ( .A(n43486), .B(n43485), .Z(n43487) );
  NAND U55628 ( .A(n43488), .B(n43487), .Z(n43489) );
  NANDN U55629 ( .A(n43490), .B(n43489), .Z(n43491) );
  NAND U55630 ( .A(n43492), .B(n43491), .Z(n43494) );
  IV U55631 ( .A(n43493), .Z(n57629) );
  AND U55632 ( .A(n43494), .B(n57629), .Z(n43495) );
  NANDN U55633 ( .A(x[5254]), .B(y[5254]), .Z(n57627) );
  AND U55634 ( .A(n43495), .B(n57627), .Z(n43499) );
  AND U55635 ( .A(n43497), .B(n43496), .Z(n43498) );
  NANDN U55636 ( .A(n43499), .B(n43498), .Z(n43500) );
  NAND U55637 ( .A(n43501), .B(n43500), .Z(n43502) );
  NAND U55638 ( .A(n43503), .B(n43502), .Z(n43504) );
  AND U55639 ( .A(n43505), .B(n43504), .Z(n43509) );
  AND U55640 ( .A(n43507), .B(n43506), .Z(n43508) );
  NANDN U55641 ( .A(n43509), .B(n43508), .Z(n43510) );
  NAND U55642 ( .A(n43511), .B(n43510), .Z(n43512) );
  NAND U55643 ( .A(n43513), .B(n43512), .Z(n43515) );
  IV U55644 ( .A(n43514), .Z(n51437) );
  AND U55645 ( .A(n43515), .B(n51437), .Z(n43516) );
  NANDN U55646 ( .A(x[5262]), .B(y[5262]), .Z(n57639) );
  AND U55647 ( .A(n43516), .B(n57639), .Z(n43520) );
  AND U55648 ( .A(n43518), .B(n43517), .Z(n43519) );
  NANDN U55649 ( .A(n43520), .B(n43519), .Z(n43521) );
  NAND U55650 ( .A(n43522), .B(n43521), .Z(n43523) );
  AND U55651 ( .A(n43524), .B(n43523), .Z(n43525) );
  OR U55652 ( .A(n43526), .B(n43525), .Z(n43527) );
  NAND U55653 ( .A(n43528), .B(n43527), .Z(n43529) );
  NANDN U55654 ( .A(n43530), .B(n43529), .Z(n43531) );
  AND U55655 ( .A(n43532), .B(n43531), .Z(n43533) );
  NOR U55656 ( .A(n43534), .B(n43533), .Z(n43535) );
  NAND U55657 ( .A(n57650), .B(n43535), .Z(n43536) );
  NANDN U55658 ( .A(n43537), .B(n43536), .Z(n43538) );
  OR U55659 ( .A(n43539), .B(n43538), .Z(n43540) );
  NAND U55660 ( .A(n43541), .B(n43540), .Z(n43542) );
  AND U55661 ( .A(n43543), .B(n43542), .Z(n43544) );
  OR U55662 ( .A(n43545), .B(n43544), .Z(n43546) );
  NAND U55663 ( .A(n43547), .B(n43546), .Z(n43548) );
  NANDN U55664 ( .A(n43549), .B(n43548), .Z(n43550) );
  NAND U55665 ( .A(n43551), .B(n43550), .Z(n43553) );
  AND U55666 ( .A(n43553), .B(n43552), .Z(n43554) );
  NANDN U55667 ( .A(n57657), .B(n43554), .Z(n43555) );
  NAND U55668 ( .A(n43556), .B(n43555), .Z(n43557) );
  NANDN U55669 ( .A(n43558), .B(n43557), .Z(n43559) );
  NAND U55670 ( .A(n43560), .B(n43559), .Z(n43561) );
  AND U55671 ( .A(n43562), .B(n43561), .Z(n43566) );
  AND U55672 ( .A(n43564), .B(n43563), .Z(n43565) );
  NANDN U55673 ( .A(n43566), .B(n43565), .Z(n43567) );
  NAND U55674 ( .A(n43568), .B(n43567), .Z(n43569) );
  AND U55675 ( .A(n43570), .B(n43569), .Z(n43571) );
  OR U55676 ( .A(n43572), .B(n43571), .Z(n43573) );
  NAND U55677 ( .A(n43574), .B(n43573), .Z(n43575) );
  NANDN U55678 ( .A(n43576), .B(n43575), .Z(n43578) );
  NANDN U55679 ( .A(n43578), .B(n43577), .Z(n43579) );
  AND U55680 ( .A(n43580), .B(n43579), .Z(n43581) );
  OR U55681 ( .A(n43582), .B(n43581), .Z(n43583) );
  NAND U55682 ( .A(n43584), .B(n43583), .Z(n43585) );
  NANDN U55683 ( .A(n43586), .B(n43585), .Z(n43587) );
  AND U55684 ( .A(n43588), .B(n43587), .Z(n43589) );
  OR U55685 ( .A(n43590), .B(n43589), .Z(n43591) );
  NAND U55686 ( .A(n43592), .B(n43591), .Z(n43593) );
  NANDN U55687 ( .A(n43594), .B(n43593), .Z(n43595) );
  NAND U55688 ( .A(n43596), .B(n43595), .Z(n43597) );
  AND U55689 ( .A(n43598), .B(n43597), .Z(n43602) );
  AND U55690 ( .A(n43600), .B(n43599), .Z(n43601) );
  NANDN U55691 ( .A(n43602), .B(n43601), .Z(n43603) );
  NAND U55692 ( .A(n43604), .B(n43603), .Z(n43605) );
  NAND U55693 ( .A(n43606), .B(n43605), .Z(n43607) );
  AND U55694 ( .A(n43608), .B(n43607), .Z(n43612) );
  AND U55695 ( .A(n43610), .B(n43609), .Z(n43611) );
  NANDN U55696 ( .A(n43612), .B(n43611), .Z(n43613) );
  NAND U55697 ( .A(n43614), .B(n43613), .Z(n43615) );
  AND U55698 ( .A(n43616), .B(n43615), .Z(n43617) );
  ANDN U55699 ( .B(n43618), .A(n43617), .Z(n43619) );
  OR U55700 ( .A(n43620), .B(n43619), .Z(n43621) );
  AND U55701 ( .A(n43622), .B(n43621), .Z(n43623) );
  OR U55702 ( .A(n43624), .B(n43623), .Z(n43625) );
  NAND U55703 ( .A(n43626), .B(n43625), .Z(n43627) );
  NANDN U55704 ( .A(n43628), .B(n43627), .Z(n43629) );
  OR U55705 ( .A(n43630), .B(n43629), .Z(n43631) );
  NAND U55706 ( .A(n43632), .B(n43631), .Z(n43633) );
  NAND U55707 ( .A(n43634), .B(n43633), .Z(n43635) );
  AND U55708 ( .A(n43636), .B(n43635), .Z(n43637) );
  OR U55709 ( .A(n43638), .B(n43637), .Z(n43639) );
  NAND U55710 ( .A(n43640), .B(n43639), .Z(n43641) );
  AND U55711 ( .A(n43642), .B(n43641), .Z(n43645) );
  NANDN U55712 ( .A(x[5318]), .B(y[5318]), .Z(n51419) );
  AND U55713 ( .A(n51419), .B(n43643), .Z(n43644) );
  NANDN U55714 ( .A(n43645), .B(n43644), .Z(n43646) );
  NANDN U55715 ( .A(n43647), .B(n43646), .Z(n43648) );
  AND U55716 ( .A(n43649), .B(n43648), .Z(n43650) );
  NAND U55717 ( .A(n57701), .B(n43650), .Z(n43651) );
  NAND U55718 ( .A(n43652), .B(n43651), .Z(n43653) );
  AND U55719 ( .A(n43653), .B(n51416), .Z(n43654) );
  NANDN U55720 ( .A(x[5322]), .B(y[5322]), .Z(n57702) );
  AND U55721 ( .A(n43654), .B(n57702), .Z(n43658) );
  XNOR U55722 ( .A(x[5324]), .B(y[5324]), .Z(n43656) );
  AND U55723 ( .A(n43656), .B(n43655), .Z(n43657) );
  NANDN U55724 ( .A(n43658), .B(n43657), .Z(n43659) );
  NAND U55725 ( .A(n43660), .B(n43659), .Z(n43661) );
  NAND U55726 ( .A(n43662), .B(n43661), .Z(n43663) );
  AND U55727 ( .A(n43663), .B(n57708), .Z(n43664) );
  NANDN U55728 ( .A(x[5326]), .B(y[5326]), .Z(n57705) );
  AND U55729 ( .A(n43664), .B(n57705), .Z(n43668) );
  AND U55730 ( .A(n43666), .B(n43665), .Z(n43667) );
  NANDN U55731 ( .A(n43668), .B(n43667), .Z(n43669) );
  NAND U55732 ( .A(n43670), .B(n43669), .Z(n43671) );
  NAND U55733 ( .A(n43672), .B(n43671), .Z(n43674) );
  AND U55734 ( .A(n43674), .B(n43673), .Z(n43675) );
  NANDN U55735 ( .A(n57714), .B(n43675), .Z(n43676) );
  NAND U55736 ( .A(n43677), .B(n43676), .Z(n43678) );
  NANDN U55737 ( .A(n43679), .B(n43678), .Z(n43680) );
  AND U55738 ( .A(n43681), .B(n43680), .Z(n43682) );
  OR U55739 ( .A(n43683), .B(n43682), .Z(n43684) );
  NAND U55740 ( .A(n43685), .B(n43684), .Z(n43686) );
  NANDN U55741 ( .A(n43687), .B(n43686), .Z(n43688) );
  NAND U55742 ( .A(n43689), .B(n43688), .Z(n43690) );
  AND U55743 ( .A(n43691), .B(n43690), .Z(n43695) );
  AND U55744 ( .A(n43693), .B(n43692), .Z(n43694) );
  NANDN U55745 ( .A(n43695), .B(n43694), .Z(n43696) );
  NAND U55746 ( .A(n43697), .B(n43696), .Z(n43698) );
  AND U55747 ( .A(n43699), .B(n43698), .Z(n43700) );
  OR U55748 ( .A(n43701), .B(n43700), .Z(n43702) );
  NAND U55749 ( .A(n43703), .B(n43702), .Z(n43704) );
  NANDN U55750 ( .A(n43705), .B(n43704), .Z(n43706) );
  AND U55751 ( .A(n43707), .B(n43706), .Z(n43708) );
  OR U55752 ( .A(n43709), .B(n43708), .Z(n43710) );
  NAND U55753 ( .A(n43711), .B(n43710), .Z(n43712) );
  NANDN U55754 ( .A(n43713), .B(n43712), .Z(n43714) );
  NAND U55755 ( .A(n43715), .B(n43714), .Z(n43716) );
  AND U55756 ( .A(n43716), .B(n57738), .Z(n43717) );
  NANDN U55757 ( .A(x[5350]), .B(y[5350]), .Z(n57734) );
  AND U55758 ( .A(n43717), .B(n57734), .Z(n43721) );
  AND U55759 ( .A(n43719), .B(n43718), .Z(n43720) );
  NANDN U55760 ( .A(n43721), .B(n43720), .Z(n43722) );
  NAND U55761 ( .A(n43723), .B(n43722), .Z(n43724) );
  AND U55762 ( .A(n43725), .B(n43724), .Z(n43726) );
  OR U55763 ( .A(n43727), .B(n43726), .Z(n43728) );
  NAND U55764 ( .A(n43729), .B(n43728), .Z(n43730) );
  NANDN U55765 ( .A(n57743), .B(n43730), .Z(n43732) );
  NANDN U55766 ( .A(n43732), .B(n43731), .Z(n43733) );
  NAND U55767 ( .A(n43734), .B(n43733), .Z(n43736) );
  IV U55768 ( .A(n43735), .Z(n57744) );
  AND U55769 ( .A(n43736), .B(n57744), .Z(n43737) );
  NANDN U55770 ( .A(x[5358]), .B(y[5358]), .Z(n57742) );
  AND U55771 ( .A(n43737), .B(n57742), .Z(n43741) );
  AND U55772 ( .A(n43739), .B(n43738), .Z(n43740) );
  NANDN U55773 ( .A(n43741), .B(n43740), .Z(n43742) );
  NAND U55774 ( .A(n43743), .B(n43742), .Z(n43744) );
  NAND U55775 ( .A(n43745), .B(n43744), .Z(n43746) );
  AND U55776 ( .A(n43746), .B(n57750), .Z(n43747) );
  NANDN U55777 ( .A(x[5362]), .B(y[5362]), .Z(n51403) );
  AND U55778 ( .A(n43747), .B(n51403), .Z(n43751) );
  AND U55779 ( .A(n43749), .B(n43748), .Z(n43750) );
  NANDN U55780 ( .A(n43751), .B(n43750), .Z(n43752) );
  NAND U55781 ( .A(n43753), .B(n43752), .Z(n43754) );
  AND U55782 ( .A(n43755), .B(n43754), .Z(n43756) );
  OR U55783 ( .A(n43757), .B(n43756), .Z(n43758) );
  NAND U55784 ( .A(n43759), .B(n43758), .Z(n43760) );
  NANDN U55785 ( .A(n43761), .B(n43760), .Z(n43762) );
  NAND U55786 ( .A(n43763), .B(n43762), .Z(n43764) );
  AND U55787 ( .A(n43764), .B(n57758), .Z(n43766) );
  NANDN U55788 ( .A(x[5370]), .B(y[5370]), .Z(n43765) );
  AND U55789 ( .A(n43766), .B(n43765), .Z(n43770) );
  AND U55790 ( .A(n43768), .B(n43767), .Z(n43769) );
  NANDN U55791 ( .A(n43770), .B(n43769), .Z(n43771) );
  NAND U55792 ( .A(n43772), .B(n43771), .Z(n43773) );
  AND U55793 ( .A(n43774), .B(n43773), .Z(n43775) );
  OR U55794 ( .A(n43776), .B(n43775), .Z(n43777) );
  NAND U55795 ( .A(n43778), .B(n43777), .Z(n43779) );
  NANDN U55796 ( .A(n43780), .B(n43779), .Z(n43781) );
  NAND U55797 ( .A(n43782), .B(n43781), .Z(n43783) );
  AND U55798 ( .A(n43784), .B(n43783), .Z(n43788) );
  AND U55799 ( .A(n43786), .B(n43785), .Z(n43787) );
  NANDN U55800 ( .A(n43788), .B(n43787), .Z(n43789) );
  NAND U55801 ( .A(n43790), .B(n43789), .Z(n43791) );
  NAND U55802 ( .A(n43792), .B(n43791), .Z(n43793) );
  AND U55803 ( .A(n43793), .B(n57773), .Z(n43794) );
  NANDN U55804 ( .A(x[5382]), .B(y[5382]), .Z(n57769) );
  AND U55805 ( .A(n43794), .B(n57769), .Z(n43798) );
  AND U55806 ( .A(n43796), .B(n43795), .Z(n43797) );
  NANDN U55807 ( .A(n43798), .B(n43797), .Z(n43799) );
  NAND U55808 ( .A(n43800), .B(n43799), .Z(n43801) );
  NAND U55809 ( .A(n43802), .B(n43801), .Z(n43803) );
  AND U55810 ( .A(n43803), .B(n57778), .Z(n43805) );
  NANDN U55811 ( .A(x[5386]), .B(y[5386]), .Z(n43804) );
  AND U55812 ( .A(n43805), .B(n43804), .Z(n43809) );
  AND U55813 ( .A(n43807), .B(n43806), .Z(n43808) );
  NANDN U55814 ( .A(n43809), .B(n43808), .Z(n43810) );
  NAND U55815 ( .A(n43811), .B(n43810), .Z(n43812) );
  NAND U55816 ( .A(n43813), .B(n43812), .Z(n43815) );
  IV U55817 ( .A(n43814), .Z(n57783) );
  AND U55818 ( .A(n43815), .B(n57783), .Z(n43816) );
  NANDN U55819 ( .A(x[5390]), .B(y[5390]), .Z(n57781) );
  AND U55820 ( .A(n43816), .B(n57781), .Z(n43820) );
  AND U55821 ( .A(n43818), .B(n43817), .Z(n43819) );
  NANDN U55822 ( .A(n43820), .B(n43819), .Z(n43821) );
  NAND U55823 ( .A(n43822), .B(n43821), .Z(n43823) );
  AND U55824 ( .A(n43824), .B(n43823), .Z(n43825) );
  ANDN U55825 ( .B(n43826), .A(n43825), .Z(n43827) );
  OR U55826 ( .A(n43828), .B(n43827), .Z(n43829) );
  NAND U55827 ( .A(n43830), .B(n43829), .Z(n43831) );
  AND U55828 ( .A(n43832), .B(n43831), .Z(n43833) );
  OR U55829 ( .A(n43834), .B(n43833), .Z(n43835) );
  NAND U55830 ( .A(n43836), .B(n43835), .Z(n43837) );
  NANDN U55831 ( .A(n43838), .B(n43837), .Z(n43839) );
  NAND U55832 ( .A(n43840), .B(n43839), .Z(n43841) );
  AND U55833 ( .A(n43842), .B(n43841), .Z(n43846) );
  AND U55834 ( .A(n43844), .B(n43843), .Z(n43845) );
  NANDN U55835 ( .A(n43846), .B(n43845), .Z(n43847) );
  NAND U55836 ( .A(n43848), .B(n43847), .Z(n43849) );
  NAND U55837 ( .A(n43850), .B(n43849), .Z(n43852) );
  IV U55838 ( .A(n43851), .Z(n57806) );
  AND U55839 ( .A(n43852), .B(n57806), .Z(n43853) );
  NANDN U55840 ( .A(x[5406]), .B(y[5406]), .Z(n57804) );
  AND U55841 ( .A(n43853), .B(n57804), .Z(n43857) );
  AND U55842 ( .A(n43855), .B(n43854), .Z(n43856) );
  NANDN U55843 ( .A(n43857), .B(n43856), .Z(n43858) );
  NAND U55844 ( .A(n43859), .B(n43858), .Z(n43860) );
  NAND U55845 ( .A(n43861), .B(n43860), .Z(n43862) );
  AND U55846 ( .A(n43862), .B(n57810), .Z(n43863) );
  NANDN U55847 ( .A(x[5410]), .B(y[5410]), .Z(n51390) );
  AND U55848 ( .A(n43863), .B(n51390), .Z(n43867) );
  AND U55849 ( .A(n43865), .B(n43864), .Z(n43866) );
  NANDN U55850 ( .A(n43867), .B(n43866), .Z(n43868) );
  NAND U55851 ( .A(n43869), .B(n43868), .Z(n43870) );
  NAND U55852 ( .A(n43871), .B(n43870), .Z(n43872) );
  AND U55853 ( .A(n43872), .B(n57817), .Z(n43873) );
  NANDN U55854 ( .A(x[5414]), .B(y[5414]), .Z(n57814) );
  AND U55855 ( .A(n43873), .B(n57814), .Z(n43877) );
  AND U55856 ( .A(n43875), .B(n43874), .Z(n43876) );
  NANDN U55857 ( .A(n43877), .B(n43876), .Z(n43878) );
  NAND U55858 ( .A(n43879), .B(n43878), .Z(n43880) );
  NAND U55859 ( .A(n43881), .B(n43880), .Z(n43882) );
  AND U55860 ( .A(n43882), .B(n57823), .Z(n43883) );
  NANDN U55861 ( .A(x[5418]), .B(y[5418]), .Z(n51387) );
  AND U55862 ( .A(n43883), .B(n51387), .Z(n43887) );
  AND U55863 ( .A(n43885), .B(n43884), .Z(n43886) );
  NANDN U55864 ( .A(n43887), .B(n43886), .Z(n43888) );
  NAND U55865 ( .A(n43889), .B(n43888), .Z(n43890) );
  AND U55866 ( .A(n43891), .B(n43890), .Z(n43892) );
  ANDN U55867 ( .B(n57827), .A(n43892), .Z(n43893) );
  NAND U55868 ( .A(n57826), .B(n43893), .Z(n43894) );
  NANDN U55869 ( .A(n43895), .B(n43894), .Z(n43896) );
  OR U55870 ( .A(n43897), .B(n43896), .Z(n43898) );
  NAND U55871 ( .A(n43899), .B(n43898), .Z(n43900) );
  NAND U55872 ( .A(n43901), .B(n43900), .Z(n43903) );
  IV U55873 ( .A(n43902), .Z(n57834) );
  AND U55874 ( .A(n43903), .B(n57834), .Z(n43904) );
  NANDN U55875 ( .A(x[5426]), .B(y[5426]), .Z(n51384) );
  AND U55876 ( .A(n43904), .B(n51384), .Z(n43905) );
  OR U55877 ( .A(n43906), .B(n43905), .Z(n43907) );
  NAND U55878 ( .A(n43908), .B(n43907), .Z(n43909) );
  NAND U55879 ( .A(n43910), .B(n43909), .Z(n43911) );
  AND U55880 ( .A(n43911), .B(n57839), .Z(n43912) );
  NANDN U55881 ( .A(x[5430]), .B(y[5430]), .Z(n57837) );
  AND U55882 ( .A(n43912), .B(n57837), .Z(n43916) );
  AND U55883 ( .A(n43914), .B(n43913), .Z(n43915) );
  NANDN U55884 ( .A(n43916), .B(n43915), .Z(n43917) );
  NAND U55885 ( .A(n43918), .B(n43917), .Z(n43919) );
  NAND U55886 ( .A(n43920), .B(n43919), .Z(n43921) );
  AND U55887 ( .A(n43921), .B(n57844), .Z(n43922) );
  NANDN U55888 ( .A(x[5434]), .B(y[5434]), .Z(n51382) );
  AND U55889 ( .A(n43922), .B(n51382), .Z(n43926) );
  AND U55890 ( .A(n43924), .B(n43923), .Z(n43925) );
  NANDN U55891 ( .A(n43926), .B(n43925), .Z(n43927) );
  NAND U55892 ( .A(n43928), .B(n43927), .Z(n43929) );
  NAND U55893 ( .A(n43930), .B(n43929), .Z(n43931) );
  AND U55894 ( .A(n43931), .B(n57850), .Z(n43932) );
  NANDN U55895 ( .A(x[5438]), .B(y[5438]), .Z(n57847) );
  AND U55896 ( .A(n43932), .B(n57847), .Z(n43936) );
  AND U55897 ( .A(n43934), .B(n43933), .Z(n43935) );
  NANDN U55898 ( .A(n43936), .B(n43935), .Z(n43937) );
  NAND U55899 ( .A(n43938), .B(n43937), .Z(n43939) );
  NAND U55900 ( .A(n43940), .B(n43939), .Z(n43941) );
  AND U55901 ( .A(n43941), .B(n57855), .Z(n43942) );
  NANDN U55902 ( .A(x[5442]), .B(y[5442]), .Z(n51380) );
  AND U55903 ( .A(n43942), .B(n51380), .Z(n43946) );
  AND U55904 ( .A(n43944), .B(n43943), .Z(n43945) );
  NANDN U55905 ( .A(n43946), .B(n43945), .Z(n43947) );
  NAND U55906 ( .A(n43948), .B(n43947), .Z(n43949) );
  NAND U55907 ( .A(n43950), .B(n43949), .Z(n43951) );
  AND U55908 ( .A(n43951), .B(n57860), .Z(n43952) );
  NANDN U55909 ( .A(x[5446]), .B(y[5446]), .Z(n57858) );
  AND U55910 ( .A(n43952), .B(n57858), .Z(n43956) );
  AND U55911 ( .A(n43954), .B(n43953), .Z(n43955) );
  NANDN U55912 ( .A(n43956), .B(n43955), .Z(n43957) );
  NAND U55913 ( .A(n43958), .B(n43957), .Z(n43959) );
  AND U55914 ( .A(n43960), .B(n43959), .Z(n43961) );
  ANDN U55915 ( .B(n57865), .A(n43961), .Z(n43962) );
  NAND U55916 ( .A(n51378), .B(n43962), .Z(n43963) );
  NANDN U55917 ( .A(n43964), .B(n43963), .Z(n43965) );
  AND U55918 ( .A(n43965), .B(n57869), .Z(n43966) );
  NANDN U55919 ( .A(x[5452]), .B(y[5452]), .Z(n57866) );
  NAND U55920 ( .A(n43966), .B(n57866), .Z(n43967) );
  NAND U55921 ( .A(n43968), .B(n43967), .Z(n43969) );
  AND U55922 ( .A(n43969), .B(n57872), .Z(n43970) );
  NANDN U55923 ( .A(x[5454]), .B(y[5454]), .Z(n57870) );
  AND U55924 ( .A(n43970), .B(n57870), .Z(n43974) );
  AND U55925 ( .A(n43972), .B(n43971), .Z(n43973) );
  NANDN U55926 ( .A(n43974), .B(n43973), .Z(n43975) );
  NAND U55927 ( .A(n43976), .B(n43975), .Z(n43977) );
  NAND U55928 ( .A(n43978), .B(n43977), .Z(n43979) );
  AND U55929 ( .A(n43979), .B(n57877), .Z(n43980) );
  NANDN U55930 ( .A(x[5458]), .B(y[5458]), .Z(n51376) );
  AND U55931 ( .A(n43980), .B(n51376), .Z(n43984) );
  AND U55932 ( .A(n43982), .B(n43981), .Z(n43983) );
  NANDN U55933 ( .A(n43984), .B(n43983), .Z(n43985) );
  NAND U55934 ( .A(n43986), .B(n43985), .Z(n43987) );
  AND U55935 ( .A(n43988), .B(n43987), .Z(n43989) );
  OR U55936 ( .A(n43990), .B(n43989), .Z(n43991) );
  NAND U55937 ( .A(n43992), .B(n43991), .Z(n43993) );
  NANDN U55938 ( .A(n43994), .B(n43993), .Z(n43995) );
  NAND U55939 ( .A(n43996), .B(n43995), .Z(n43998) );
  IV U55940 ( .A(n43997), .Z(n57884) );
  AND U55941 ( .A(n43998), .B(n57884), .Z(n44000) );
  NANDN U55942 ( .A(x[5466]), .B(y[5466]), .Z(n43999) );
  AND U55943 ( .A(n44000), .B(n43999), .Z(n44004) );
  AND U55944 ( .A(n44002), .B(n44001), .Z(n44003) );
  NANDN U55945 ( .A(n44004), .B(n44003), .Z(n44005) );
  NAND U55946 ( .A(n44006), .B(n44005), .Z(n44007) );
  NAND U55947 ( .A(n44008), .B(n44007), .Z(n44009) );
  AND U55948 ( .A(n44009), .B(n57888), .Z(n44010) );
  NANDN U55949 ( .A(x[5470]), .B(y[5470]), .Z(n51371) );
  AND U55950 ( .A(n44010), .B(n51371), .Z(n44014) );
  AND U55951 ( .A(n44012), .B(n44011), .Z(n44013) );
  NANDN U55952 ( .A(n44014), .B(n44013), .Z(n44015) );
  NAND U55953 ( .A(n44016), .B(n44015), .Z(n44017) );
  AND U55954 ( .A(n44018), .B(n44017), .Z(n44019) );
  OR U55955 ( .A(n44020), .B(n44019), .Z(n44021) );
  NAND U55956 ( .A(n44022), .B(n44021), .Z(n44023) );
  NANDN U55957 ( .A(n57896), .B(n44023), .Z(n44025) );
  NANDN U55958 ( .A(n44025), .B(n44024), .Z(n44026) );
  AND U55959 ( .A(n44027), .B(n44026), .Z(n44028) );
  OR U55960 ( .A(n44029), .B(n44028), .Z(n44030) );
  NAND U55961 ( .A(n44031), .B(n44030), .Z(n44032) );
  NANDN U55962 ( .A(n44033), .B(n44032), .Z(n44034) );
  AND U55963 ( .A(n44035), .B(n44034), .Z(n44036) );
  OR U55964 ( .A(n44037), .B(n44036), .Z(n44038) );
  NAND U55965 ( .A(n44039), .B(n44038), .Z(n44040) );
  NAND U55966 ( .A(n44041), .B(n44040), .Z(n44042) );
  AND U55967 ( .A(n44043), .B(n44042), .Z(n44046) );
  NANDN U55968 ( .A(x[5486]), .B(y[5486]), .Z(n57903) );
  AND U55969 ( .A(n57903), .B(n44044), .Z(n44045) );
  NANDN U55970 ( .A(n44046), .B(n44045), .Z(n44047) );
  NANDN U55971 ( .A(n44048), .B(n44047), .Z(n44049) );
  AND U55972 ( .A(n44050), .B(n44049), .Z(n44051) );
  NAND U55973 ( .A(n57909), .B(n44051), .Z(n44052) );
  NAND U55974 ( .A(n44053), .B(n44052), .Z(n44055) );
  IV U55975 ( .A(n44054), .Z(n57910) );
  AND U55976 ( .A(n44055), .B(n57910), .Z(n44056) );
  NANDN U55977 ( .A(x[5490]), .B(y[5490]), .Z(n57908) );
  AND U55978 ( .A(n44056), .B(n57908), .Z(n44060) );
  AND U55979 ( .A(n44058), .B(n44057), .Z(n44059) );
  NANDN U55980 ( .A(n44060), .B(n44059), .Z(n44061) );
  NAND U55981 ( .A(n44062), .B(n44061), .Z(n44063) );
  NAND U55982 ( .A(n44064), .B(n44063), .Z(n44066) );
  AND U55983 ( .A(n44066), .B(n44065), .Z(n44067) );
  NANDN U55984 ( .A(n57914), .B(n44067), .Z(n44068) );
  NAND U55985 ( .A(n44069), .B(n44068), .Z(n44070) );
  NANDN U55986 ( .A(n44071), .B(n44070), .Z(n44072) );
  AND U55987 ( .A(n44073), .B(n44072), .Z(n44074) );
  OR U55988 ( .A(n44075), .B(n44074), .Z(n44076) );
  NAND U55989 ( .A(n44077), .B(n44076), .Z(n44078) );
  NANDN U55990 ( .A(n44079), .B(n44078), .Z(n44080) );
  NAND U55991 ( .A(n44081), .B(n44080), .Z(n44082) );
  AND U55992 ( .A(n44082), .B(n57926), .Z(n44084) );
  NANDN U55993 ( .A(x[5502]), .B(y[5502]), .Z(n44083) );
  AND U55994 ( .A(n44084), .B(n44083), .Z(n44088) );
  AND U55995 ( .A(n44086), .B(n44085), .Z(n44087) );
  NANDN U55996 ( .A(n44088), .B(n44087), .Z(n44089) );
  NAND U55997 ( .A(n44090), .B(n44089), .Z(n44091) );
  NAND U55998 ( .A(n44092), .B(n44091), .Z(n44093) );
  AND U55999 ( .A(n44093), .B(n57931), .Z(n44094) );
  NANDN U56000 ( .A(x[5506]), .B(y[5506]), .Z(n57928) );
  AND U56001 ( .A(n44094), .B(n57928), .Z(n44098) );
  AND U56002 ( .A(n44096), .B(n44095), .Z(n44097) );
  NANDN U56003 ( .A(n44098), .B(n44097), .Z(n44099) );
  NAND U56004 ( .A(n44100), .B(n44099), .Z(n44101) );
  AND U56005 ( .A(n44102), .B(n44101), .Z(n44103) );
  ANDN U56006 ( .B(n51359), .A(n44103), .Z(n44104) );
  NAND U56007 ( .A(n44105), .B(n44104), .Z(n44106) );
  NANDN U56008 ( .A(n44107), .B(n44106), .Z(n44108) );
  AND U56009 ( .A(n44108), .B(n57937), .Z(n44109) );
  NANDN U56010 ( .A(x[5512]), .B(y[5512]), .Z(n51360) );
  NAND U56011 ( .A(n44109), .B(n51360), .Z(n44110) );
  AND U56012 ( .A(n44111), .B(n44110), .Z(n44114) );
  NANDN U56013 ( .A(x[5514]), .B(y[5514]), .Z(n51358) );
  AND U56014 ( .A(n44112), .B(n51358), .Z(n44113) );
  NANDN U56015 ( .A(n44114), .B(n44113), .Z(n44115) );
  NANDN U56016 ( .A(n44116), .B(n44115), .Z(n44117) );
  AND U56017 ( .A(n44118), .B(n44117), .Z(n44119) );
  NAND U56018 ( .A(n57939), .B(n44119), .Z(n44120) );
  NAND U56019 ( .A(n44121), .B(n44120), .Z(n44122) );
  AND U56020 ( .A(n57946), .B(n44122), .Z(n44123) );
  OR U56021 ( .A(n44124), .B(n44123), .Z(n44125) );
  NAND U56022 ( .A(n44126), .B(n44125), .Z(n44127) );
  NAND U56023 ( .A(n44128), .B(n44127), .Z(n44130) );
  IV U56024 ( .A(n44129), .Z(n51354) );
  AND U56025 ( .A(n44130), .B(n51354), .Z(n44131) );
  NANDN U56026 ( .A(x[5522]), .B(y[5522]), .Z(n57949) );
  AND U56027 ( .A(n44131), .B(n57949), .Z(n44135) );
  AND U56028 ( .A(n44133), .B(n44132), .Z(n44134) );
  NANDN U56029 ( .A(n44135), .B(n44134), .Z(n44136) );
  NAND U56030 ( .A(n44137), .B(n44136), .Z(n44138) );
  NAND U56031 ( .A(n44139), .B(n44138), .Z(n44141) );
  AND U56032 ( .A(n44141), .B(n44140), .Z(n44142) );
  NANDN U56033 ( .A(x[5526]), .B(y[5526]), .Z(n57952) );
  AND U56034 ( .A(n44142), .B(n57952), .Z(n44143) );
  OR U56035 ( .A(n44144), .B(n44143), .Z(n44145) );
  NAND U56036 ( .A(n44146), .B(n44145), .Z(n44147) );
  AND U56037 ( .A(n44148), .B(n44147), .Z(n44149) );
  ANDN U56038 ( .B(n57959), .A(n44149), .Z(n44150) );
  NANDN U56039 ( .A(x[5530]), .B(y[5530]), .Z(n51352) );
  AND U56040 ( .A(n44150), .B(n51352), .Z(n44151) );
  OR U56041 ( .A(n44152), .B(n44151), .Z(n44153) );
  NAND U56042 ( .A(n44154), .B(n44153), .Z(n44155) );
  NAND U56043 ( .A(n44156), .B(n44155), .Z(n44157) );
  AND U56044 ( .A(n44157), .B(n57964), .Z(n44158) );
  NANDN U56045 ( .A(x[5534]), .B(y[5534]), .Z(n57962) );
  AND U56046 ( .A(n44158), .B(n57962), .Z(n44162) );
  AND U56047 ( .A(n44160), .B(n44159), .Z(n44161) );
  NANDN U56048 ( .A(n44162), .B(n44161), .Z(n44163) );
  NAND U56049 ( .A(n44164), .B(n44163), .Z(n44165) );
  AND U56050 ( .A(n44166), .B(n44165), .Z(n44167) );
  OR U56051 ( .A(n44168), .B(n44167), .Z(n44169) );
  NAND U56052 ( .A(n44170), .B(n44169), .Z(n44171) );
  NANDN U56053 ( .A(n57972), .B(n44171), .Z(n44173) );
  NANDN U56054 ( .A(x[5540]), .B(y[5540]), .Z(n44172) );
  NANDN U56055 ( .A(n44173), .B(n44172), .Z(n44174) );
  AND U56056 ( .A(n44175), .B(n44174), .Z(n44176) );
  OR U56057 ( .A(n44177), .B(n44176), .Z(n44178) );
  NAND U56058 ( .A(n44179), .B(n44178), .Z(n44180) );
  NANDN U56059 ( .A(n44181), .B(n44180), .Z(n44182) );
  NAND U56060 ( .A(n44183), .B(n44182), .Z(n44185) );
  IV U56061 ( .A(n44184), .Z(n57977) );
  AND U56062 ( .A(n44185), .B(n57977), .Z(n44186) );
  NANDN U56063 ( .A(x[5546]), .B(y[5546]), .Z(n51349) );
  AND U56064 ( .A(n44186), .B(n51349), .Z(n44190) );
  AND U56065 ( .A(n44188), .B(n44187), .Z(n44189) );
  NANDN U56066 ( .A(n44190), .B(n44189), .Z(n44191) );
  NAND U56067 ( .A(n44192), .B(n44191), .Z(n44193) );
  NAND U56068 ( .A(n44194), .B(n44193), .Z(n44196) );
  IV U56069 ( .A(n44195), .Z(n51346) );
  AND U56070 ( .A(n44196), .B(n51346), .Z(n44197) );
  NANDN U56071 ( .A(x[5550]), .B(y[5550]), .Z(n57981) );
  AND U56072 ( .A(n44197), .B(n57981), .Z(n44201) );
  AND U56073 ( .A(n44199), .B(n44198), .Z(n44200) );
  NANDN U56074 ( .A(n44201), .B(n44200), .Z(n44202) );
  NAND U56075 ( .A(n44203), .B(n44202), .Z(n44204) );
  NAND U56076 ( .A(n44205), .B(n44204), .Z(n44206) );
  AND U56077 ( .A(n44206), .B(n57988), .Z(n44207) );
  NANDN U56078 ( .A(x[5554]), .B(y[5554]), .Z(n57985) );
  AND U56079 ( .A(n44207), .B(n57985), .Z(n44211) );
  AND U56080 ( .A(n44209), .B(n44208), .Z(n44210) );
  NANDN U56081 ( .A(n44211), .B(n44210), .Z(n44212) );
  NAND U56082 ( .A(n44213), .B(n44212), .Z(n44214) );
  NAND U56083 ( .A(n44215), .B(n44214), .Z(n44217) );
  IV U56084 ( .A(n44216), .Z(n51344) );
  AND U56085 ( .A(n44217), .B(n51344), .Z(n44218) );
  NANDN U56086 ( .A(x[5558]), .B(y[5558]), .Z(n57992) );
  AND U56087 ( .A(n44218), .B(n57992), .Z(n44222) );
  AND U56088 ( .A(n44220), .B(n44219), .Z(n44221) );
  NANDN U56089 ( .A(n44222), .B(n44221), .Z(n44223) );
  NAND U56090 ( .A(n44224), .B(n44223), .Z(n44225) );
  NAND U56091 ( .A(n44226), .B(n44225), .Z(n44227) );
  AND U56092 ( .A(n44227), .B(n58000), .Z(n44228) );
  NANDN U56093 ( .A(x[5562]), .B(y[5562]), .Z(n57996) );
  AND U56094 ( .A(n44228), .B(n57996), .Z(n44232) );
  AND U56095 ( .A(n44230), .B(n44229), .Z(n44231) );
  NANDN U56096 ( .A(n44232), .B(n44231), .Z(n44233) );
  NAND U56097 ( .A(n44234), .B(n44233), .Z(n44235) );
  NAND U56098 ( .A(n44236), .B(n44235), .Z(n44238) );
  AND U56099 ( .A(n44238), .B(n44237), .Z(n44239) );
  NANDN U56100 ( .A(n58004), .B(n44239), .Z(n44240) );
  NAND U56101 ( .A(n44241), .B(n44240), .Z(n44242) );
  NANDN U56102 ( .A(n44243), .B(n44242), .Z(n44244) );
  AND U56103 ( .A(n44245), .B(n44244), .Z(n44246) );
  OR U56104 ( .A(n44247), .B(n44246), .Z(n44248) );
  NAND U56105 ( .A(n44249), .B(n44248), .Z(n44250) );
  NANDN U56106 ( .A(n44251), .B(n44250), .Z(n44253) );
  NANDN U56107 ( .A(x[5572]), .B(y[5572]), .Z(n44252) );
  NANDN U56108 ( .A(n44253), .B(n44252), .Z(n44254) );
  NAND U56109 ( .A(n44255), .B(n44254), .Z(n44257) );
  AND U56110 ( .A(n44257), .B(n44256), .Z(n44259) );
  NANDN U56111 ( .A(x[5574]), .B(y[5574]), .Z(n44258) );
  NAND U56112 ( .A(n44259), .B(n44258), .Z(n44260) );
  NAND U56113 ( .A(n44261), .B(n44260), .Z(n44267) );
  NAND U56114 ( .A(n44263), .B(n44262), .Z(n44264) );
  NAND U56115 ( .A(n44265), .B(n44264), .Z(n44266) );
  AND U56116 ( .A(n44267), .B(n44266), .Z(n44268) );
  OR U56117 ( .A(n44269), .B(n44268), .Z(n44270) );
  NAND U56118 ( .A(n44271), .B(n44270), .Z(n44272) );
  NANDN U56119 ( .A(n44273), .B(n44272), .Z(n44275) );
  NANDN U56120 ( .A(n44275), .B(n44274), .Z(n44277) );
  AND U56121 ( .A(n44277), .B(n44276), .Z(n44278) );
  NANDN U56122 ( .A(x[5580]), .B(y[5580]), .Z(n58019) );
  NAND U56123 ( .A(n44278), .B(n58019), .Z(n44279) );
  AND U56124 ( .A(n44280), .B(n44279), .Z(n44281) );
  ANDN U56125 ( .B(n51343), .A(n44281), .Z(n44282) );
  NAND U56126 ( .A(n44283), .B(n44282), .Z(n44284) );
  NANDN U56127 ( .A(n44285), .B(n44284), .Z(n44286) );
  AND U56128 ( .A(n44286), .B(n58026), .Z(n44287) );
  NANDN U56129 ( .A(x[5584]), .B(y[5584]), .Z(n51342) );
  AND U56130 ( .A(n44287), .B(n51342), .Z(n44288) );
  OR U56131 ( .A(n44289), .B(n44288), .Z(n44290) );
  NAND U56132 ( .A(n44291), .B(n44290), .Z(n44292) );
  NANDN U56133 ( .A(n44293), .B(n44292), .Z(n44294) );
  NAND U56134 ( .A(n44295), .B(n44294), .Z(n44296) );
  AND U56135 ( .A(n44297), .B(n44296), .Z(n44298) );
  ANDN U56136 ( .B(n44299), .A(n44298), .Z(n44300) );
  NAND U56137 ( .A(n51341), .B(n44300), .Z(n44301) );
  NANDN U56138 ( .A(n44302), .B(n44301), .Z(n44303) );
  AND U56139 ( .A(n44304), .B(n44303), .Z(n44305) );
  OR U56140 ( .A(n44306), .B(n44305), .Z(n44307) );
  NAND U56141 ( .A(n44308), .B(n44307), .Z(n44309) );
  NANDN U56142 ( .A(n44310), .B(n44309), .Z(n44311) );
  AND U56143 ( .A(n44311), .B(n58039), .Z(n44313) );
  NANDN U56144 ( .A(x[5596]), .B(y[5596]), .Z(n44312) );
  AND U56145 ( .A(n44313), .B(n44312), .Z(n44314) );
  OR U56146 ( .A(n44315), .B(n44314), .Z(n44316) );
  NAND U56147 ( .A(n44317), .B(n44316), .Z(n44318) );
  NANDN U56148 ( .A(n44319), .B(n44318), .Z(n44320) );
  AND U56149 ( .A(n44321), .B(n44320), .Z(n44322) );
  OR U56150 ( .A(n44323), .B(n44322), .Z(n44324) );
  NAND U56151 ( .A(n44325), .B(n44324), .Z(n44326) );
  NANDN U56152 ( .A(n44327), .B(n44326), .Z(n44329) );
  AND U56153 ( .A(n44329), .B(n44328), .Z(n44330) );
  NANDN U56154 ( .A(x[5604]), .B(y[5604]), .Z(n58046) );
  NAND U56155 ( .A(n44330), .B(n58046), .Z(n44331) );
  AND U56156 ( .A(n44332), .B(n44331), .Z(n44333) );
  OR U56157 ( .A(n44334), .B(n44333), .Z(n44335) );
  NAND U56158 ( .A(n44336), .B(n44335), .Z(n44338) );
  AND U56159 ( .A(n44338), .B(n44337), .Z(n44339) );
  NANDN U56160 ( .A(x[5608]), .B(y[5608]), .Z(n51337) );
  AND U56161 ( .A(n44339), .B(n51337), .Z(n44340) );
  OR U56162 ( .A(n44341), .B(n44340), .Z(n44342) );
  NAND U56163 ( .A(n44343), .B(n44342), .Z(n44344) );
  NANDN U56164 ( .A(n44345), .B(n44344), .Z(n44347) );
  NANDN U56165 ( .A(n44347), .B(n44346), .Z(n44349) );
  IV U56166 ( .A(n44348), .Z(n51334) );
  AND U56167 ( .A(n44349), .B(n51334), .Z(n44350) );
  NANDN U56168 ( .A(x[5612]), .B(y[5612]), .Z(n58055) );
  NAND U56169 ( .A(n44350), .B(n58055), .Z(n44351) );
  NAND U56170 ( .A(n44352), .B(n44351), .Z(n44355) );
  NANDN U56171 ( .A(x[5614]), .B(y[5614]), .Z(n51335) );
  AND U56172 ( .A(n44353), .B(n51335), .Z(n44354) );
  NAND U56173 ( .A(n44355), .B(n44354), .Z(n44356) );
  NANDN U56174 ( .A(n44357), .B(n44356), .Z(n44359) );
  AND U56175 ( .A(n44359), .B(n44358), .Z(n44361) );
  NANDN U56176 ( .A(x[5616]), .B(y[5616]), .Z(n44360) );
  AND U56177 ( .A(n44361), .B(n44360), .Z(n44362) );
  OR U56178 ( .A(n44363), .B(n44362), .Z(n44364) );
  NAND U56179 ( .A(n44365), .B(n44364), .Z(n44366) );
  NANDN U56180 ( .A(n44367), .B(n44366), .Z(n44369) );
  AND U56181 ( .A(n44369), .B(n44368), .Z(n44370) );
  NANDN U56182 ( .A(x[5620]), .B(y[5620]), .Z(n51331) );
  AND U56183 ( .A(n44370), .B(n51331), .Z(n44371) );
  OR U56184 ( .A(n44372), .B(n44371), .Z(n44373) );
  NAND U56185 ( .A(n44374), .B(n44373), .Z(n44375) );
  NANDN U56186 ( .A(n44376), .B(n44375), .Z(n44377) );
  AND U56187 ( .A(n44377), .B(n51328), .Z(n44378) );
  NANDN U56188 ( .A(x[5624]), .B(y[5624]), .Z(n58066) );
  NAND U56189 ( .A(n44378), .B(n58066), .Z(n44379) );
  NAND U56190 ( .A(n44380), .B(n44379), .Z(n44382) );
  NANDN U56191 ( .A(x[5626]), .B(y[5626]), .Z(n51329) );
  AND U56192 ( .A(n58070), .B(n51329), .Z(n44381) );
  NAND U56193 ( .A(n44382), .B(n44381), .Z(n44383) );
  NANDN U56194 ( .A(n44384), .B(n44383), .Z(n44385) );
  AND U56195 ( .A(n44385), .B(n58073), .Z(n44386) );
  NANDN U56196 ( .A(x[5628]), .B(y[5628]), .Z(n58069) );
  NAND U56197 ( .A(n44386), .B(n58069), .Z(n44387) );
  AND U56198 ( .A(n44388), .B(n44387), .Z(n44389) );
  NOR U56199 ( .A(n58074), .B(n44389), .Z(n44390) );
  NAND U56200 ( .A(n58077), .B(n44390), .Z(n44391) );
  NANDN U56201 ( .A(n44392), .B(n44391), .Z(n44394) );
  NANDN U56202 ( .A(n44394), .B(n44393), .Z(n44396) );
  IV U56203 ( .A(n44395), .Z(n51326) );
  AND U56204 ( .A(n44396), .B(n51326), .Z(n44397) );
  NANDN U56205 ( .A(x[5632]), .B(y[5632]), .Z(n58078) );
  NAND U56206 ( .A(n44397), .B(n58078), .Z(n44398) );
  AND U56207 ( .A(n44399), .B(n44398), .Z(n44400) );
  ANDN U56208 ( .B(n58082), .A(n44400), .Z(n44401) );
  NAND U56209 ( .A(n51327), .B(n44401), .Z(n44402) );
  NANDN U56210 ( .A(n44403), .B(n44402), .Z(n44404) );
  AND U56211 ( .A(n44404), .B(n58084), .Z(n44405) );
  NANDN U56212 ( .A(x[5636]), .B(y[5636]), .Z(n58081) );
  NAND U56213 ( .A(n44405), .B(n58081), .Z(n44406) );
  AND U56214 ( .A(n44407), .B(n44406), .Z(n44408) );
  ANDN U56215 ( .B(n58087), .A(n44408), .Z(n44409) );
  NAND U56216 ( .A(n58085), .B(n44409), .Z(n44410) );
  NANDN U56217 ( .A(n44411), .B(n44410), .Z(n44413) );
  IV U56218 ( .A(n44412), .Z(n51324) );
  AND U56219 ( .A(n44413), .B(n51324), .Z(n44414) );
  NANDN U56220 ( .A(x[5640]), .B(y[5640]), .Z(n58088) );
  NAND U56221 ( .A(n44414), .B(n58088), .Z(n44415) );
  AND U56222 ( .A(n44416), .B(n44415), .Z(n44417) );
  ANDN U56223 ( .B(n58094), .A(n44417), .Z(n44418) );
  NAND U56224 ( .A(n51325), .B(n44418), .Z(n44419) );
  NANDN U56225 ( .A(n44420), .B(n44419), .Z(n44421) );
  AND U56226 ( .A(n44421), .B(n58096), .Z(n44422) );
  NANDN U56227 ( .A(x[5644]), .B(y[5644]), .Z(n58093) );
  NAND U56228 ( .A(n44422), .B(n58093), .Z(n44423) );
  AND U56229 ( .A(n44424), .B(n44423), .Z(n44425) );
  ANDN U56230 ( .B(n58099), .A(n44425), .Z(n44426) );
  NAND U56231 ( .A(n58097), .B(n44426), .Z(n44427) );
  NANDN U56232 ( .A(n44428), .B(n44427), .Z(n44429) );
  AND U56233 ( .A(n44429), .B(n51322), .Z(n44430) );
  NANDN U56234 ( .A(x[5648]), .B(y[5648]), .Z(n58100) );
  AND U56235 ( .A(n44430), .B(n58100), .Z(n44431) );
  OR U56236 ( .A(n44432), .B(n44431), .Z(n44433) );
  NAND U56237 ( .A(n44434), .B(n44433), .Z(n44435) );
  NANDN U56238 ( .A(n44436), .B(n44435), .Z(n44437) );
  AND U56239 ( .A(n44437), .B(n58105), .Z(n44439) );
  NANDN U56240 ( .A(x[5652]), .B(y[5652]), .Z(n44438) );
  NAND U56241 ( .A(n44439), .B(n44438), .Z(n44440) );
  AND U56242 ( .A(n44441), .B(n44440), .Z(n44442) );
  ANDN U56243 ( .B(n51320), .A(n44442), .Z(n44443) );
  NAND U56244 ( .A(n58106), .B(n44443), .Z(n44444) );
  NANDN U56245 ( .A(n44445), .B(n44444), .Z(n44447) );
  NANDN U56246 ( .A(n44447), .B(n44446), .Z(n44448) );
  AND U56247 ( .A(n44448), .B(n58112), .Z(n44449) );
  NANDN U56248 ( .A(x[5656]), .B(y[5656]), .Z(n51321) );
  NAND U56249 ( .A(n44449), .B(n51321), .Z(n44450) );
  AND U56250 ( .A(n44451), .B(n44450), .Z(n44452) );
  ANDN U56251 ( .B(n58113), .A(n44452), .Z(n44453) );
  NAND U56252 ( .A(n58111), .B(n44453), .Z(n44454) );
  NANDN U56253 ( .A(n44455), .B(n44454), .Z(n44456) );
  AND U56254 ( .A(n44456), .B(n58116), .Z(n44457) );
  NANDN U56255 ( .A(x[5660]), .B(y[5660]), .Z(n58114) );
  NAND U56256 ( .A(n44457), .B(n58114), .Z(n44458) );
  AND U56257 ( .A(n44459), .B(n44458), .Z(n44460) );
  ANDN U56258 ( .B(n51317), .A(n44460), .Z(n44461) );
  NAND U56259 ( .A(n58117), .B(n44461), .Z(n44462) );
  NANDN U56260 ( .A(n44463), .B(n44462), .Z(n44465) );
  AND U56261 ( .A(n44465), .B(n44464), .Z(n44466) );
  NANDN U56262 ( .A(x[5664]), .B(y[5664]), .Z(n51318) );
  AND U56263 ( .A(n44466), .B(n51318), .Z(n44467) );
  OR U56264 ( .A(n44468), .B(n44467), .Z(n44469) );
  NAND U56265 ( .A(n44470), .B(n44469), .Z(n44471) );
  NANDN U56266 ( .A(n44472), .B(n44471), .Z(n44474) );
  IV U56267 ( .A(n44473), .Z(n51315) );
  AND U56268 ( .A(n44474), .B(n51315), .Z(n44475) );
  NANDN U56269 ( .A(x[5668]), .B(y[5668]), .Z(n58124) );
  NAND U56270 ( .A(n44475), .B(n58124), .Z(n44476) );
  AND U56271 ( .A(n44477), .B(n44476), .Z(n44478) );
  ANDN U56272 ( .B(n44479), .A(n44478), .Z(n44480) );
  NAND U56273 ( .A(n51316), .B(n44480), .Z(n44481) );
  NANDN U56274 ( .A(n44482), .B(n44481), .Z(n44483) );
  NAND U56275 ( .A(n44484), .B(n44483), .Z(n44485) );
  NAND U56276 ( .A(n44486), .B(n44485), .Z(n44488) );
  NANDN U56277 ( .A(x[5674]), .B(y[5674]), .Z(n51312) );
  AND U56278 ( .A(n58129), .B(n51312), .Z(n44487) );
  NAND U56279 ( .A(n44488), .B(n44487), .Z(n44489) );
  NANDN U56280 ( .A(n44490), .B(n44489), .Z(n44491) );
  AND U56281 ( .A(n44491), .B(n58135), .Z(n44492) );
  NANDN U56282 ( .A(x[5676]), .B(y[5676]), .Z(n58130) );
  NAND U56283 ( .A(n44492), .B(n58130), .Z(n44493) );
  AND U56284 ( .A(n44494), .B(n44493), .Z(n44495) );
  ANDN U56285 ( .B(n58138), .A(n44495), .Z(n44496) );
  NAND U56286 ( .A(n58134), .B(n44496), .Z(n44497) );
  NANDN U56287 ( .A(n44498), .B(n44497), .Z(n44500) );
  IV U56288 ( .A(n44499), .Z(n58141) );
  AND U56289 ( .A(n44500), .B(n58141), .Z(n44501) );
  NANDN U56290 ( .A(x[5680]), .B(y[5680]), .Z(n58139) );
  NAND U56291 ( .A(n44501), .B(n58139), .Z(n44502) );
  AND U56292 ( .A(n44503), .B(n44502), .Z(n44504) );
  NOR U56293 ( .A(n58142), .B(n44504), .Z(n44505) );
  NAND U56294 ( .A(n51310), .B(n44505), .Z(n44506) );
  NANDN U56295 ( .A(n44507), .B(n44506), .Z(n44509) );
  NANDN U56296 ( .A(n44509), .B(n44508), .Z(n44510) );
  AND U56297 ( .A(n44510), .B(n58146), .Z(n44511) );
  NANDN U56298 ( .A(x[5684]), .B(y[5684]), .Z(n51311) );
  NAND U56299 ( .A(n44511), .B(n51311), .Z(n44512) );
  AND U56300 ( .A(n44513), .B(n44512), .Z(n44514) );
  ANDN U56301 ( .B(n58147), .A(n44514), .Z(n44515) );
  NAND U56302 ( .A(n58145), .B(n44515), .Z(n44516) );
  NANDN U56303 ( .A(n44517), .B(n44516), .Z(n44518) );
  AND U56304 ( .A(n44518), .B(n58151), .Z(n44519) );
  NANDN U56305 ( .A(x[5688]), .B(y[5688]), .Z(n58149) );
  NAND U56306 ( .A(n44519), .B(n58149), .Z(n44520) );
  AND U56307 ( .A(n44521), .B(n44520), .Z(n44522) );
  ANDN U56308 ( .B(n44523), .A(n44522), .Z(n44524) );
  NAND U56309 ( .A(n58152), .B(n44524), .Z(n44525) );
  NANDN U56310 ( .A(n44526), .B(n44525), .Z(n44527) );
  NAND U56311 ( .A(n44528), .B(n44527), .Z(n44529) );
  AND U56312 ( .A(n44530), .B(n44529), .Z(n44531) );
  ANDN U56313 ( .B(n58156), .A(n44531), .Z(n44532) );
  NAND U56314 ( .A(n51308), .B(n44532), .Z(n44533) );
  NANDN U56315 ( .A(n44534), .B(n44533), .Z(n44535) );
  AND U56316 ( .A(n44535), .B(n51304), .Z(n44536) );
  NANDN U56317 ( .A(x[5696]), .B(y[5696]), .Z(n58157) );
  AND U56318 ( .A(n44536), .B(n58157), .Z(n44537) );
  OR U56319 ( .A(n44538), .B(n44537), .Z(n44539) );
  NAND U56320 ( .A(n44540), .B(n44539), .Z(n44541) );
  NANDN U56321 ( .A(n44542), .B(n44541), .Z(n44543) );
  AND U56322 ( .A(n44543), .B(n58163), .Z(n44545) );
  NANDN U56323 ( .A(x[5700]), .B(y[5700]), .Z(n44544) );
  NAND U56324 ( .A(n44545), .B(n44544), .Z(n44546) );
  AND U56325 ( .A(n44547), .B(n44546), .Z(n44548) );
  ANDN U56326 ( .B(n44549), .A(n44548), .Z(n44550) );
  NAND U56327 ( .A(n58164), .B(n44550), .Z(n44551) );
  NANDN U56328 ( .A(n44552), .B(n44551), .Z(n44553) );
  AND U56329 ( .A(n44554), .B(n44553), .Z(n44555) );
  OR U56330 ( .A(n44556), .B(n44555), .Z(n44557) );
  NAND U56331 ( .A(n44558), .B(n44557), .Z(n44559) );
  NANDN U56332 ( .A(n44560), .B(n44559), .Z(n44562) );
  NANDN U56333 ( .A(n44562), .B(n44561), .Z(n44563) );
  AND U56334 ( .A(n44563), .B(n51302), .Z(n44564) );
  NANDN U56335 ( .A(x[5708]), .B(y[5708]), .Z(n58171) );
  AND U56336 ( .A(n44564), .B(n58171), .Z(n44565) );
  OR U56337 ( .A(n44566), .B(n44565), .Z(n44567) );
  NAND U56338 ( .A(n44568), .B(n44567), .Z(n44569) );
  NANDN U56339 ( .A(n44570), .B(n44569), .Z(n44571) );
  OR U56340 ( .A(n44572), .B(n44571), .Z(n44574) );
  IV U56341 ( .A(n44573), .Z(n58178) );
  AND U56342 ( .A(n44574), .B(n58178), .Z(n44575) );
  NANDN U56343 ( .A(x[5712]), .B(y[5712]), .Z(n58175) );
  NAND U56344 ( .A(n44575), .B(n58175), .Z(n44576) );
  AND U56345 ( .A(n44577), .B(n44576), .Z(n44580) );
  NANDN U56346 ( .A(x[5714]), .B(y[5714]), .Z(n51300) );
  AND U56347 ( .A(n44578), .B(n51300), .Z(n44579) );
  NANDN U56348 ( .A(n44580), .B(n44579), .Z(n44581) );
  NANDN U56349 ( .A(n44582), .B(n44581), .Z(n44583) );
  AND U56350 ( .A(n58181), .B(n44583), .Z(n44585) );
  NANDN U56351 ( .A(x[5716]), .B(y[5716]), .Z(n44584) );
  NAND U56352 ( .A(n44585), .B(n44584), .Z(n44586) );
  AND U56353 ( .A(n44587), .B(n44586), .Z(n44589) );
  NANDN U56354 ( .A(x[5718]), .B(y[5718]), .Z(n58180) );
  AND U56355 ( .A(n58182), .B(n58180), .Z(n44588) );
  NANDN U56356 ( .A(n44589), .B(n44588), .Z(n44590) );
  NANDN U56357 ( .A(n44591), .B(n44590), .Z(n44592) );
  AND U56358 ( .A(n58185), .B(n44592), .Z(n44593) );
  NANDN U56359 ( .A(x[5720]), .B(y[5720]), .Z(n58183) );
  NAND U56360 ( .A(n44593), .B(n58183), .Z(n44594) );
  AND U56361 ( .A(n44595), .B(n44594), .Z(n44597) );
  NANDN U56362 ( .A(x[5722]), .B(y[5722]), .Z(n58186) );
  AND U56363 ( .A(n58186), .B(n51295), .Z(n44596) );
  NANDN U56364 ( .A(n44597), .B(n44596), .Z(n44598) );
  NANDN U56365 ( .A(n44599), .B(n44598), .Z(n44600) );
  AND U56366 ( .A(n44600), .B(n58190), .Z(n44601) );
  NANDN U56367 ( .A(x[5724]), .B(y[5724]), .Z(n51296) );
  NAND U56368 ( .A(n44601), .B(n51296), .Z(n44602) );
  AND U56369 ( .A(n44603), .B(n44602), .Z(n44606) );
  NANDN U56370 ( .A(x[5726]), .B(y[5726]), .Z(n58191) );
  IV U56371 ( .A(n44604), .Z(n58192) );
  AND U56372 ( .A(n58191), .B(n58192), .Z(n44605) );
  NANDN U56373 ( .A(n44606), .B(n44605), .Z(n44607) );
  NANDN U56374 ( .A(n44608), .B(n44607), .Z(n44609) );
  AND U56375 ( .A(n58195), .B(n44609), .Z(n44610) );
  NANDN U56376 ( .A(x[5728]), .B(y[5728]), .Z(n58193) );
  NAND U56377 ( .A(n44610), .B(n58193), .Z(n44611) );
  NAND U56378 ( .A(n44612), .B(n44611), .Z(n44614) );
  AND U56379 ( .A(n44614), .B(n44613), .Z(n44615) );
  NANDN U56380 ( .A(x[5730]), .B(y[5730]), .Z(n58196) );
  AND U56381 ( .A(n44615), .B(n58196), .Z(n44616) );
  NOR U56382 ( .A(n44617), .B(n44616), .Z(n44619) );
  NAND U56383 ( .A(n44619), .B(n44618), .Z(n44621) );
  IV U56384 ( .A(n44620), .Z(n58198) );
  AND U56385 ( .A(n44621), .B(n58198), .Z(n44623) );
  NANDN U56386 ( .A(x[5732]), .B(y[5732]), .Z(n44622) );
  AND U56387 ( .A(n44623), .B(n44622), .Z(n44627) );
  AND U56388 ( .A(n44625), .B(n44624), .Z(n44626) );
  NANDN U56389 ( .A(n44627), .B(n44626), .Z(n44628) );
  NAND U56390 ( .A(n44629), .B(n44628), .Z(n44633) );
  ANDN U56391 ( .B(n44631), .A(n44630), .Z(n44632) );
  NAND U56392 ( .A(n44633), .B(n44632), .Z(n44634) );
  AND U56393 ( .A(n51290), .B(n44634), .Z(n44635) );
  NANDN U56394 ( .A(x[5736]), .B(y[5736]), .Z(n58203) );
  NAND U56395 ( .A(n44635), .B(n58203), .Z(n44636) );
  AND U56396 ( .A(n44637), .B(n44636), .Z(n44639) );
  NANDN U56397 ( .A(x[5738]), .B(y[5738]), .Z(n51291) );
  AND U56398 ( .A(n51291), .B(n58206), .Z(n44638) );
  NANDN U56399 ( .A(n44639), .B(n44638), .Z(n44640) );
  NANDN U56400 ( .A(n44641), .B(n44640), .Z(n44642) );
  AND U56401 ( .A(n58209), .B(n44642), .Z(n44643) );
  NANDN U56402 ( .A(x[5740]), .B(y[5740]), .Z(n58207) );
  NAND U56403 ( .A(n44643), .B(n58207), .Z(n44644) );
  AND U56404 ( .A(n44645), .B(n44644), .Z(n44647) );
  NANDN U56405 ( .A(x[5742]), .B(y[5742]), .Z(n51289) );
  AND U56406 ( .A(n58211), .B(n51289), .Z(n44646) );
  NANDN U56407 ( .A(n44647), .B(n44646), .Z(n44648) );
  NANDN U56408 ( .A(n44649), .B(n44648), .Z(n44650) );
  AND U56409 ( .A(n51287), .B(n44650), .Z(n44651) );
  NANDN U56410 ( .A(x[5744]), .B(y[5744]), .Z(n58212) );
  NAND U56411 ( .A(n44651), .B(n58212), .Z(n44652) );
  AND U56412 ( .A(n44653), .B(n44652), .Z(n44656) );
  NANDN U56413 ( .A(x[5746]), .B(y[5746]), .Z(n51288) );
  AND U56414 ( .A(n51288), .B(n44654), .Z(n44655) );
  NANDN U56415 ( .A(n44656), .B(n44655), .Z(n44657) );
  NANDN U56416 ( .A(n44658), .B(n44657), .Z(n44660) );
  IV U56417 ( .A(n44659), .Z(n58217) );
  AND U56418 ( .A(n44660), .B(n58217), .Z(n44662) );
  NAND U56419 ( .A(n44662), .B(n44661), .Z(n44663) );
  AND U56420 ( .A(n44664), .B(n44663), .Z(n44666) );
  NANDN U56421 ( .A(x[5750]), .B(y[5750]), .Z(n58218) );
  AND U56422 ( .A(n58218), .B(n51284), .Z(n44665) );
  NANDN U56423 ( .A(n44666), .B(n44665), .Z(n44667) );
  NANDN U56424 ( .A(n44668), .B(n44667), .Z(n44669) );
  AND U56425 ( .A(n44669), .B(n58222), .Z(n44670) );
  NANDN U56426 ( .A(x[5752]), .B(y[5752]), .Z(n51285) );
  NAND U56427 ( .A(n44670), .B(n51285), .Z(n44671) );
  AND U56428 ( .A(n44672), .B(n44671), .Z(n44674) );
  NANDN U56429 ( .A(x[5754]), .B(y[5754]), .Z(n58221) );
  AND U56430 ( .A(n58225), .B(n58221), .Z(n44673) );
  NANDN U56431 ( .A(n44674), .B(n44673), .Z(n44675) );
  NANDN U56432 ( .A(n44676), .B(n44675), .Z(n44678) );
  IV U56433 ( .A(n44677), .Z(n58228) );
  AND U56434 ( .A(n44678), .B(n58228), .Z(n44679) );
  NANDN U56435 ( .A(x[5756]), .B(y[5756]), .Z(n58226) );
  NAND U56436 ( .A(n44679), .B(n58226), .Z(n44680) );
  AND U56437 ( .A(n44681), .B(n44680), .Z(n44684) );
  NANDN U56438 ( .A(x[5758]), .B(y[5758]), .Z(n58229) );
  IV U56439 ( .A(n44682), .Z(n51282) );
  AND U56440 ( .A(n58229), .B(n51282), .Z(n44683) );
  NANDN U56441 ( .A(n44684), .B(n44683), .Z(n44685) );
  NANDN U56442 ( .A(n44686), .B(n44685), .Z(n44687) );
  AND U56443 ( .A(n44688), .B(n44687), .Z(n44689) );
  NANDN U56444 ( .A(x[5760]), .B(y[5760]), .Z(n51283) );
  AND U56445 ( .A(n44689), .B(n51283), .Z(n44690) );
  OR U56446 ( .A(n44691), .B(n44690), .Z(n44692) );
  NAND U56447 ( .A(n44693), .B(n44692), .Z(n44694) );
  NAND U56448 ( .A(n44695), .B(n44694), .Z(n44696) );
  AND U56449 ( .A(n44697), .B(n44696), .Z(n44698) );
  OR U56450 ( .A(n44699), .B(n44698), .Z(n44700) );
  NAND U56451 ( .A(n44701), .B(n44700), .Z(n44702) );
  NANDN U56452 ( .A(n44703), .B(n44702), .Z(n44705) );
  NANDN U56453 ( .A(n44705), .B(n44704), .Z(n44706) );
  AND U56454 ( .A(n44707), .B(n44706), .Z(n44711) );
  AND U56455 ( .A(n44709), .B(n44708), .Z(n44710) );
  NANDN U56456 ( .A(n44711), .B(n44710), .Z(n44712) );
  NANDN U56457 ( .A(n44713), .B(n44712), .Z(n44714) );
  AND U56458 ( .A(n44715), .B(n44714), .Z(n44717) );
  NAND U56459 ( .A(n44717), .B(n44716), .Z(n44718) );
  AND U56460 ( .A(n44719), .B(n44718), .Z(n44720) );
  OR U56461 ( .A(n44721), .B(n44720), .Z(n44722) );
  NAND U56462 ( .A(n44723), .B(n44722), .Z(n44724) );
  NANDN U56463 ( .A(n44725), .B(n44724), .Z(n44726) );
  AND U56464 ( .A(n44727), .B(n44726), .Z(n44728) );
  OR U56465 ( .A(n44729), .B(n44728), .Z(n44730) );
  NAND U56466 ( .A(n44731), .B(n44730), .Z(n44732) );
  NANDN U56467 ( .A(n44733), .B(n44732), .Z(n44734) );
  AND U56468 ( .A(n44734), .B(n51276), .Z(n44735) );
  NANDN U56469 ( .A(x[5780]), .B(y[5780]), .Z(n58251) );
  NAND U56470 ( .A(n44735), .B(n58251), .Z(n44736) );
  NAND U56471 ( .A(n44737), .B(n44736), .Z(n44739) );
  NANDN U56472 ( .A(x[5782]), .B(y[5782]), .Z(n51275) );
  AND U56473 ( .A(n58255), .B(n51275), .Z(n44738) );
  NAND U56474 ( .A(n44739), .B(n44738), .Z(n44740) );
  NANDN U56475 ( .A(n44741), .B(n44740), .Z(n44742) );
  AND U56476 ( .A(n44742), .B(n58257), .Z(n44743) );
  NANDN U56477 ( .A(x[5784]), .B(y[5784]), .Z(n58254) );
  NAND U56478 ( .A(n44743), .B(n58254), .Z(n44744) );
  AND U56479 ( .A(n44745), .B(n44744), .Z(n44746) );
  ANDN U56480 ( .B(n58260), .A(n44746), .Z(n44747) );
  NAND U56481 ( .A(n58258), .B(n44747), .Z(n44748) );
  NANDN U56482 ( .A(n44749), .B(n44748), .Z(n44751) );
  IV U56483 ( .A(n44750), .Z(n51273) );
  AND U56484 ( .A(n44751), .B(n51273), .Z(n44752) );
  NANDN U56485 ( .A(x[5788]), .B(y[5788]), .Z(n58261) );
  AND U56486 ( .A(n44752), .B(n58261), .Z(n44756) );
  AND U56487 ( .A(n44754), .B(n44753), .Z(n44755) );
  NANDN U56488 ( .A(n44756), .B(n44755), .Z(n44757) );
  AND U56489 ( .A(n44757), .B(n51271), .Z(n44758) );
  NANDN U56490 ( .A(x[5790]), .B(y[5790]), .Z(n51274) );
  AND U56491 ( .A(n44758), .B(n51274), .Z(n44759) );
  NOR U56492 ( .A(n44760), .B(n44759), .Z(n44762) );
  NAND U56493 ( .A(n44762), .B(n44761), .Z(n44763) );
  AND U56494 ( .A(n44763), .B(n58266), .Z(n44764) );
  NANDN U56495 ( .A(x[5792]), .B(y[5792]), .Z(n51272) );
  NAND U56496 ( .A(n44764), .B(n51272), .Z(n44765) );
  AND U56497 ( .A(n44766), .B(n44765), .Z(n44767) );
  ANDN U56498 ( .B(n58269), .A(n44767), .Z(n44768) );
  NAND U56499 ( .A(n58267), .B(n44768), .Z(n44769) );
  NANDN U56500 ( .A(n44770), .B(n44769), .Z(n44772) );
  IV U56501 ( .A(n44771), .Z(n58272) );
  AND U56502 ( .A(n44772), .B(n58272), .Z(n44773) );
  NANDN U56503 ( .A(x[5796]), .B(y[5796]), .Z(n58270) );
  AND U56504 ( .A(n44773), .B(n58270), .Z(n44774) );
  OR U56505 ( .A(n44775), .B(n44774), .Z(n44776) );
  NAND U56506 ( .A(n44777), .B(n44776), .Z(n44778) );
  NANDN U56507 ( .A(n44779), .B(n44778), .Z(n44781) );
  OR U56508 ( .A(n44781), .B(n44780), .Z(n44782) );
  AND U56509 ( .A(n58278), .B(n44782), .Z(n44783) );
  NANDN U56510 ( .A(x[5800]), .B(y[5800]), .Z(n58275) );
  NAND U56511 ( .A(n44783), .B(n58275), .Z(n44784) );
  AND U56512 ( .A(n44785), .B(n44784), .Z(n44787) );
  NANDN U56513 ( .A(x[5802]), .B(y[5802]), .Z(n58279) );
  AND U56514 ( .A(n58279), .B(n58281), .Z(n44786) );
  NANDN U56515 ( .A(n44787), .B(n44786), .Z(n44788) );
  NANDN U56516 ( .A(n44789), .B(n44788), .Z(n44791) );
  IV U56517 ( .A(n44790), .Z(n51268) );
  AND U56518 ( .A(n44791), .B(n51268), .Z(n44792) );
  NANDN U56519 ( .A(x[5804]), .B(y[5804]), .Z(n58282) );
  NAND U56520 ( .A(n44792), .B(n58282), .Z(n44793) );
  AND U56521 ( .A(n44794), .B(n44793), .Z(n44796) );
  NANDN U56522 ( .A(x[5806]), .B(y[5806]), .Z(n51269) );
  AND U56523 ( .A(n51269), .B(n58292), .Z(n44795) );
  NANDN U56524 ( .A(n44796), .B(n44795), .Z(n44797) );
  NANDN U56525 ( .A(n44798), .B(n44797), .Z(n44799) );
  AND U56526 ( .A(n58298), .B(n44799), .Z(n44800) );
  NANDN U56527 ( .A(x[5808]), .B(y[5808]), .Z(n58291) );
  NAND U56528 ( .A(n44800), .B(n58291), .Z(n44801) );
  AND U56529 ( .A(n44802), .B(n44801), .Z(n44804) );
  NANDN U56530 ( .A(x[5810]), .B(y[5810]), .Z(n58299) );
  AND U56531 ( .A(n58299), .B(n58304), .Z(n44803) );
  NANDN U56532 ( .A(n44804), .B(n44803), .Z(n44805) );
  NANDN U56533 ( .A(n44806), .B(n44805), .Z(n44807) );
  AND U56534 ( .A(n44808), .B(n44807), .Z(n44809) );
  NANDN U56535 ( .A(x[5812]), .B(y[5812]), .Z(n58305) );
  NAND U56536 ( .A(n44809), .B(n58305), .Z(n44810) );
  AND U56537 ( .A(n44811), .B(n44810), .Z(n44814) );
  NAND U56538 ( .A(n44812), .B(n51266), .Z(n44813) );
  OR U56539 ( .A(n44814), .B(n44813), .Z(n44815) );
  NAND U56540 ( .A(n44816), .B(n44815), .Z(n44818) );
  AND U56541 ( .A(n44818), .B(n44817), .Z(n44819) );
  NANDN U56542 ( .A(x[5816]), .B(y[5816]), .Z(n51267) );
  AND U56543 ( .A(n44819), .B(n51267), .Z(n44820) );
  OR U56544 ( .A(n44821), .B(n44820), .Z(n44822) );
  NAND U56545 ( .A(n44823), .B(n44822), .Z(n44824) );
  NANDN U56546 ( .A(n44825), .B(n44824), .Z(n44827) );
  IV U56547 ( .A(n44826), .Z(n58323) );
  AND U56548 ( .A(n44827), .B(n58323), .Z(n44828) );
  NANDN U56549 ( .A(x[5820]), .B(y[5820]), .Z(n51263) );
  AND U56550 ( .A(n44828), .B(n51263), .Z(n44829) );
  OR U56551 ( .A(n44830), .B(n44829), .Z(n44831) );
  NAND U56552 ( .A(n44832), .B(n44831), .Z(n44833) );
  NAND U56553 ( .A(n44834), .B(n44833), .Z(n44835) );
  NAND U56554 ( .A(n44836), .B(n44835), .Z(n44837) );
  AND U56555 ( .A(n44838), .B(n44837), .Z(n44839) );
  NOR U56556 ( .A(n51261), .B(n44839), .Z(n44840) );
  NAND U56557 ( .A(n58329), .B(n44840), .Z(n44841) );
  NANDN U56558 ( .A(n44842), .B(n44841), .Z(n44844) );
  XNOR U56559 ( .A(x[5828]), .B(y[5828]), .Z(n44843) );
  NANDN U56560 ( .A(n44844), .B(n44843), .Z(n44846) );
  IV U56561 ( .A(n44845), .Z(n58330) );
  AND U56562 ( .A(n44846), .B(n58330), .Z(n44847) );
  NANDN U56563 ( .A(x[5828]), .B(y[5828]), .Z(n58328) );
  NAND U56564 ( .A(n44847), .B(n58328), .Z(n44848) );
  AND U56565 ( .A(n44849), .B(n44848), .Z(n44850) );
  ANDN U56566 ( .B(n58333), .A(n44850), .Z(n44851) );
  NAND U56567 ( .A(n58331), .B(n44851), .Z(n44852) );
  NANDN U56568 ( .A(n44853), .B(n44852), .Z(n44855) );
  AND U56569 ( .A(n44855), .B(n44854), .Z(n44856) );
  NANDN U56570 ( .A(x[5832]), .B(y[5832]), .Z(n58334) );
  AND U56571 ( .A(n44856), .B(n58334), .Z(n44857) );
  OR U56572 ( .A(n44858), .B(n44857), .Z(n44859) );
  NAND U56573 ( .A(n44860), .B(n44859), .Z(n44861) );
  NANDN U56574 ( .A(n44862), .B(n44861), .Z(n44864) );
  IV U56575 ( .A(n44863), .Z(n58341) );
  AND U56576 ( .A(n44864), .B(n58341), .Z(n44865) );
  NANDN U56577 ( .A(x[5836]), .B(y[5836]), .Z(n58339) );
  NAND U56578 ( .A(n44865), .B(n58339), .Z(n44866) );
  AND U56579 ( .A(n44867), .B(n44866), .Z(n44868) );
  ANDN U56580 ( .B(n58344), .A(n44868), .Z(n44869) );
  NAND U56581 ( .A(n58342), .B(n44869), .Z(n44870) );
  NANDN U56582 ( .A(n44871), .B(n44870), .Z(n44872) );
  AND U56583 ( .A(n44872), .B(n51257), .Z(n44873) );
  NANDN U56584 ( .A(x[5840]), .B(y[5840]), .Z(n58345) );
  NAND U56585 ( .A(n44873), .B(n58345), .Z(n44874) );
  AND U56586 ( .A(n44875), .B(n44874), .Z(n44876) );
  ANDN U56587 ( .B(n58349), .A(n44876), .Z(n44877) );
  NAND U56588 ( .A(n51258), .B(n44877), .Z(n44878) );
  NANDN U56589 ( .A(n44879), .B(n44878), .Z(n44881) );
  IV U56590 ( .A(n44880), .Z(n58351) );
  AND U56591 ( .A(n44881), .B(n58351), .Z(n44882) );
  NANDN U56592 ( .A(x[5844]), .B(y[5844]), .Z(n58348) );
  NAND U56593 ( .A(n44882), .B(n58348), .Z(n44883) );
  AND U56594 ( .A(n44884), .B(n44883), .Z(n44885) );
  ANDN U56595 ( .B(n58354), .A(n44885), .Z(n44886) );
  NAND U56596 ( .A(n58352), .B(n44886), .Z(n44887) );
  NANDN U56597 ( .A(n44888), .B(n44887), .Z(n44889) );
  AND U56598 ( .A(n44889), .B(n51254), .Z(n44890) );
  NANDN U56599 ( .A(x[5848]), .B(y[5848]), .Z(n58355) );
  AND U56600 ( .A(n44890), .B(n58355), .Z(n44891) );
  OR U56601 ( .A(n44892), .B(n44891), .Z(n44893) );
  NAND U56602 ( .A(n44894), .B(n44893), .Z(n44895) );
  NANDN U56603 ( .A(n44896), .B(n44895), .Z(n44897) );
  OR U56604 ( .A(n44898), .B(n44897), .Z(n44900) );
  IV U56605 ( .A(n44899), .Z(n58360) );
  AND U56606 ( .A(n44900), .B(n58360), .Z(n44901) );
  NANDN U56607 ( .A(x[5852]), .B(y[5852]), .Z(n58358) );
  NAND U56608 ( .A(n44901), .B(n58358), .Z(n44902) );
  AND U56609 ( .A(n44903), .B(n44902), .Z(n44905) );
  NANDN U56610 ( .A(x[5854]), .B(y[5854]), .Z(n58361) );
  AND U56611 ( .A(n58361), .B(n58363), .Z(n44904) );
  NANDN U56612 ( .A(n44905), .B(n44904), .Z(n44906) );
  NANDN U56613 ( .A(n44907), .B(n44906), .Z(n44908) );
  AND U56614 ( .A(n44909), .B(n44908), .Z(n44910) );
  NANDN U56615 ( .A(x[5856]), .B(y[5856]), .Z(n58364) );
  NAND U56616 ( .A(n44910), .B(n58364), .Z(n44911) );
  AND U56617 ( .A(n44912), .B(n44911), .Z(n44913) );
  OR U56618 ( .A(n44914), .B(n44913), .Z(n44915) );
  NAND U56619 ( .A(n44916), .B(n44915), .Z(n44917) );
  NAND U56620 ( .A(n44918), .B(n44917), .Z(n44919) );
  AND U56621 ( .A(n44920), .B(n44919), .Z(n44921) );
  ANDN U56622 ( .B(n58374), .A(n44921), .Z(n44922) );
  NAND U56623 ( .A(n58372), .B(n44922), .Z(n44923) );
  NANDN U56624 ( .A(n44924), .B(n44923), .Z(n44926) );
  AND U56625 ( .A(n44926), .B(n44925), .Z(n44927) );
  NANDN U56626 ( .A(x[5864]), .B(y[5864]), .Z(n58373) );
  AND U56627 ( .A(n44927), .B(n58373), .Z(n44928) );
  OR U56628 ( .A(n44929), .B(n44928), .Z(n44930) );
  NAND U56629 ( .A(n44931), .B(n44930), .Z(n44932) );
  NANDN U56630 ( .A(n44933), .B(n44932), .Z(n44935) );
  IV U56631 ( .A(n44934), .Z(n51249) );
  AND U56632 ( .A(n44935), .B(n51249), .Z(n44936) );
  NANDN U56633 ( .A(x[5868]), .B(y[5868]), .Z(n58378) );
  NAND U56634 ( .A(n44936), .B(n58378), .Z(n44937) );
  AND U56635 ( .A(n44938), .B(n44937), .Z(n44939) );
  ANDN U56636 ( .B(n44940), .A(n44939), .Z(n44941) );
  NAND U56637 ( .A(n51250), .B(n44941), .Z(n44942) );
  NANDN U56638 ( .A(n44943), .B(n44942), .Z(n44944) );
  NAND U56639 ( .A(n44945), .B(n44944), .Z(n44946) );
  AND U56640 ( .A(n44947), .B(n44946), .Z(n44948) );
  ANDN U56641 ( .B(n51245), .A(n44948), .Z(n44949) );
  NAND U56642 ( .A(n58383), .B(n44949), .Z(n44950) );
  NANDN U56643 ( .A(n44951), .B(n44950), .Z(n44952) );
  AND U56644 ( .A(n44952), .B(n58386), .Z(n44953) );
  NANDN U56645 ( .A(x[5876]), .B(y[5876]), .Z(n51246) );
  AND U56646 ( .A(n44953), .B(n51246), .Z(n44957) );
  AND U56647 ( .A(n44955), .B(n44954), .Z(n44956) );
  NANDN U56648 ( .A(n44957), .B(n44956), .Z(n44958) );
  NAND U56649 ( .A(n44959), .B(n44958), .Z(n44960) );
  NANDN U56650 ( .A(n44961), .B(n44960), .Z(n44963) );
  IV U56651 ( .A(n44962), .Z(n58393) );
  AND U56652 ( .A(n44963), .B(n58393), .Z(n44964) );
  NANDN U56653 ( .A(x[5880]), .B(y[5880]), .Z(n58391) );
  NAND U56654 ( .A(n44964), .B(n58391), .Z(n44965) );
  AND U56655 ( .A(n44966), .B(n44965), .Z(n44968) );
  NANDN U56656 ( .A(x[5882]), .B(y[5882]), .Z(n58394) );
  AND U56657 ( .A(n58394), .B(n51243), .Z(n44967) );
  NANDN U56658 ( .A(n44968), .B(n44967), .Z(n44969) );
  NANDN U56659 ( .A(n44970), .B(n44969), .Z(n44971) );
  AND U56660 ( .A(n44971), .B(n58398), .Z(n44972) );
  NANDN U56661 ( .A(x[5884]), .B(y[5884]), .Z(n51244) );
  NAND U56662 ( .A(n44972), .B(n51244), .Z(n44973) );
  AND U56663 ( .A(n44974), .B(n44973), .Z(n44976) );
  NANDN U56664 ( .A(x[5886]), .B(y[5886]), .Z(n58397) );
  AND U56665 ( .A(n58400), .B(n58397), .Z(n44975) );
  NANDN U56666 ( .A(n44976), .B(n44975), .Z(n44977) );
  NANDN U56667 ( .A(n44978), .B(n44977), .Z(n44980) );
  IV U56668 ( .A(n44979), .Z(n58403) );
  AND U56669 ( .A(n44980), .B(n58403), .Z(n44981) );
  NANDN U56670 ( .A(x[5888]), .B(y[5888]), .Z(n58401) );
  NAND U56671 ( .A(n44981), .B(n58401), .Z(n44982) );
  AND U56672 ( .A(n44983), .B(n44982), .Z(n44985) );
  NANDN U56673 ( .A(x[5890]), .B(y[5890]), .Z(n58405) );
  AND U56674 ( .A(n58405), .B(n51241), .Z(n44984) );
  NANDN U56675 ( .A(n44985), .B(n44984), .Z(n44986) );
  NANDN U56676 ( .A(n44987), .B(n44986), .Z(n44988) );
  AND U56677 ( .A(n44988), .B(n58409), .Z(n44989) );
  NANDN U56678 ( .A(x[5892]), .B(y[5892]), .Z(n51242) );
  NAND U56679 ( .A(n44989), .B(n51242), .Z(n44990) );
  AND U56680 ( .A(n44991), .B(n44990), .Z(n44993) );
  NANDN U56681 ( .A(x[5894]), .B(y[5894]), .Z(n58408) );
  AND U56682 ( .A(n58411), .B(n58408), .Z(n44992) );
  NANDN U56683 ( .A(n44993), .B(n44992), .Z(n44994) );
  NANDN U56684 ( .A(n44995), .B(n44994), .Z(n44997) );
  IV U56685 ( .A(n44996), .Z(n58414) );
  AND U56686 ( .A(n44997), .B(n58414), .Z(n44998) );
  NANDN U56687 ( .A(x[5896]), .B(y[5896]), .Z(n58412) );
  NAND U56688 ( .A(n44998), .B(n58412), .Z(n44999) );
  AND U56689 ( .A(n45000), .B(n44999), .Z(n45002) );
  NANDN U56690 ( .A(x[5898]), .B(y[5898]), .Z(n58415) );
  AND U56691 ( .A(n58415), .B(n51239), .Z(n45001) );
  NANDN U56692 ( .A(n45002), .B(n45001), .Z(n45003) );
  NANDN U56693 ( .A(n45004), .B(n45003), .Z(n45005) );
  AND U56694 ( .A(n45005), .B(n58422), .Z(n45006) );
  NANDN U56695 ( .A(x[5900]), .B(y[5900]), .Z(n51240) );
  NAND U56696 ( .A(n45006), .B(n51240), .Z(n45007) );
  AND U56697 ( .A(n45008), .B(n45007), .Z(n45010) );
  NANDN U56698 ( .A(x[5902]), .B(y[5902]), .Z(n58420) );
  AND U56699 ( .A(n58424), .B(n58420), .Z(n45009) );
  NANDN U56700 ( .A(n45010), .B(n45009), .Z(n45011) );
  NANDN U56701 ( .A(n45012), .B(n45011), .Z(n45014) );
  IV U56702 ( .A(n45013), .Z(n58427) );
  AND U56703 ( .A(n45014), .B(n58427), .Z(n45015) );
  NANDN U56704 ( .A(x[5904]), .B(y[5904]), .Z(n58425) );
  NAND U56705 ( .A(n45015), .B(n58425), .Z(n45016) );
  AND U56706 ( .A(n45017), .B(n45016), .Z(n45019) );
  NANDN U56707 ( .A(x[5906]), .B(y[5906]), .Z(n58428) );
  AND U56708 ( .A(n58428), .B(n51237), .Z(n45018) );
  NANDN U56709 ( .A(n45019), .B(n45018), .Z(n45020) );
  NANDN U56710 ( .A(n45021), .B(n45020), .Z(n45022) );
  AND U56711 ( .A(n58432), .B(n45022), .Z(n45023) );
  NANDN U56712 ( .A(x[5908]), .B(y[5908]), .Z(n51238) );
  NAND U56713 ( .A(n45023), .B(n51238), .Z(n45024) );
  AND U56714 ( .A(n45025), .B(n45024), .Z(n45027) );
  NANDN U56715 ( .A(x[5910]), .B(y[5910]), .Z(n58431) );
  AND U56716 ( .A(n58431), .B(n58434), .Z(n45026) );
  NANDN U56717 ( .A(n45027), .B(n45026), .Z(n45028) );
  NANDN U56718 ( .A(n45029), .B(n45028), .Z(n45031) );
  IV U56719 ( .A(n45030), .Z(n58439) );
  AND U56720 ( .A(n45031), .B(n58439), .Z(n45032) );
  NANDN U56721 ( .A(x[5912]), .B(y[5912]), .Z(n58435) );
  NAND U56722 ( .A(n45032), .B(n58435), .Z(n45033) );
  AND U56723 ( .A(n45034), .B(n45033), .Z(n45036) );
  NANDN U56724 ( .A(x[5914]), .B(y[5914]), .Z(n58440) );
  AND U56725 ( .A(n58440), .B(n51235), .Z(n45035) );
  NANDN U56726 ( .A(n45036), .B(n45035), .Z(n45037) );
  NANDN U56727 ( .A(n45038), .B(n45037), .Z(n45039) );
  AND U56728 ( .A(n45039), .B(n58443), .Z(n45040) );
  NANDN U56729 ( .A(x[5916]), .B(y[5916]), .Z(n51236) );
  NAND U56730 ( .A(n45040), .B(n51236), .Z(n45041) );
  AND U56731 ( .A(n45042), .B(n45041), .Z(n45045) );
  NANDN U56732 ( .A(x[5918]), .B(y[5918]), .Z(n58444) );
  AND U56733 ( .A(n45043), .B(n58444), .Z(n45044) );
  NANDN U56734 ( .A(n45045), .B(n45044), .Z(n45046) );
  NANDN U56735 ( .A(n45047), .B(n45046), .Z(n45048) );
  AND U56736 ( .A(n45049), .B(n45048), .Z(n45051) );
  NANDN U56737 ( .A(x[5920]), .B(y[5920]), .Z(n45050) );
  NAND U56738 ( .A(n45051), .B(n45050), .Z(n45052) );
  AND U56739 ( .A(n45053), .B(n45052), .Z(n45054) );
  OR U56740 ( .A(n45055), .B(n45054), .Z(n45056) );
  NAND U56741 ( .A(n45057), .B(n45056), .Z(n45058) );
  AND U56742 ( .A(n45058), .B(n58452), .Z(n45059) );
  NANDN U56743 ( .A(x[5924]), .B(y[5924]), .Z(n58448) );
  NAND U56744 ( .A(n45059), .B(n58448), .Z(n45060) );
  AND U56745 ( .A(n45061), .B(n45060), .Z(n45062) );
  ANDN U56746 ( .B(n58455), .A(n45062), .Z(n45063) );
  NAND U56747 ( .A(n58453), .B(n45063), .Z(n45064) );
  NANDN U56748 ( .A(n45065), .B(n45064), .Z(n45067) );
  IV U56749 ( .A(n45066), .Z(n51231) );
  AND U56750 ( .A(n45067), .B(n51231), .Z(n45068) );
  NANDN U56751 ( .A(x[5928]), .B(y[5928]), .Z(n58456) );
  AND U56752 ( .A(n45068), .B(n58456), .Z(n45069) );
  OR U56753 ( .A(n45070), .B(n45069), .Z(n45071) );
  NAND U56754 ( .A(n45072), .B(n45071), .Z(n45076) );
  ANDN U56755 ( .B(n45074), .A(n45073), .Z(n45075) );
  NAND U56756 ( .A(n45076), .B(n45075), .Z(n45077) );
  AND U56757 ( .A(n58462), .B(n45077), .Z(n45078) );
  NANDN U56758 ( .A(x[5932]), .B(y[5932]), .Z(n58460) );
  NAND U56759 ( .A(n45078), .B(n58460), .Z(n45079) );
  AND U56760 ( .A(n45080), .B(n45079), .Z(n45083) );
  NANDN U56761 ( .A(x[5934]), .B(y[5934]), .Z(n51230) );
  AND U56762 ( .A(n45081), .B(n51230), .Z(n45082) );
  NANDN U56763 ( .A(n45083), .B(n45082), .Z(n45084) );
  NANDN U56764 ( .A(n45085), .B(n45084), .Z(n45086) );
  AND U56765 ( .A(n45086), .B(n58466), .Z(n45088) );
  NANDN U56766 ( .A(x[5936]), .B(y[5936]), .Z(n45087) );
  NAND U56767 ( .A(n45088), .B(n45087), .Z(n45089) );
  AND U56768 ( .A(n45090), .B(n45089), .Z(n45092) );
  NANDN U56769 ( .A(x[5938]), .B(y[5938]), .Z(n58465) );
  AND U56770 ( .A(n58468), .B(n58465), .Z(n45091) );
  NANDN U56771 ( .A(n45092), .B(n45091), .Z(n45093) );
  NANDN U56772 ( .A(n45094), .B(n45093), .Z(n45096) );
  IV U56773 ( .A(n45095), .Z(n58471) );
  AND U56774 ( .A(n45096), .B(n58471), .Z(n45097) );
  NANDN U56775 ( .A(x[5940]), .B(y[5940]), .Z(n58469) );
  NAND U56776 ( .A(n45097), .B(n58469), .Z(n45098) );
  AND U56777 ( .A(n45099), .B(n45098), .Z(n45101) );
  NANDN U56778 ( .A(x[5942]), .B(y[5942]), .Z(n58472) );
  AND U56779 ( .A(n58472), .B(n51226), .Z(n45100) );
  NANDN U56780 ( .A(n45101), .B(n45100), .Z(n45102) );
  NANDN U56781 ( .A(n45103), .B(n45102), .Z(n45104) );
  AND U56782 ( .A(n45104), .B(n58477), .Z(n45105) );
  NANDN U56783 ( .A(x[5944]), .B(y[5944]), .Z(n51227) );
  NAND U56784 ( .A(n45105), .B(n51227), .Z(n45106) );
  AND U56785 ( .A(n45107), .B(n45106), .Z(n45110) );
  NANDN U56786 ( .A(x[5946]), .B(y[5946]), .Z(n58479) );
  IV U56787 ( .A(n45108), .Z(n58481) );
  AND U56788 ( .A(n58479), .B(n58481), .Z(n45109) );
  NANDN U56789 ( .A(n45110), .B(n45109), .Z(n45111) );
  NANDN U56790 ( .A(n45112), .B(n45111), .Z(n45114) );
  IV U56791 ( .A(n45113), .Z(n58484) );
  AND U56792 ( .A(n45114), .B(n58484), .Z(n45115) );
  NANDN U56793 ( .A(x[5948]), .B(y[5948]), .Z(n58482) );
  NAND U56794 ( .A(n45115), .B(n58482), .Z(n45116) );
  NAND U56795 ( .A(n45117), .B(n45116), .Z(n45118) );
  AND U56796 ( .A(n45118), .B(n51224), .Z(n45119) );
  NANDN U56797 ( .A(x[5950]), .B(y[5950]), .Z(n58485) );
  AND U56798 ( .A(n45119), .B(n58485), .Z(n45123) );
  AND U56799 ( .A(n45121), .B(n45120), .Z(n45122) );
  NANDN U56800 ( .A(n45123), .B(n45122), .Z(n45125) );
  AND U56801 ( .A(n45125), .B(n45124), .Z(n45126) );
  NANDN U56802 ( .A(x[5952]), .B(y[5952]), .Z(n51225) );
  AND U56803 ( .A(n45126), .B(n51225), .Z(n45127) );
  OR U56804 ( .A(n45128), .B(n45127), .Z(n45129) );
  NAND U56805 ( .A(n45130), .B(n45129), .Z(n45131) );
  NANDN U56806 ( .A(n45132), .B(n45131), .Z(n45134) );
  NANDN U56807 ( .A(n45134), .B(n45133), .Z(n45135) );
  AND U56808 ( .A(n45135), .B(n51222), .Z(n45136) );
  NANDN U56809 ( .A(x[5956]), .B(y[5956]), .Z(n58491) );
  NAND U56810 ( .A(n45136), .B(n58491), .Z(n45137) );
  AND U56811 ( .A(n45138), .B(n45137), .Z(n45139) );
  ANDN U56812 ( .B(n45140), .A(n45139), .Z(n45141) );
  NAND U56813 ( .A(n51223), .B(n45141), .Z(n45142) );
  NANDN U56814 ( .A(n45143), .B(n45142), .Z(n45144) );
  NAND U56815 ( .A(n45145), .B(n45144), .Z(n45146) );
  AND U56816 ( .A(n45147), .B(n45146), .Z(n45148) );
  ANDN U56817 ( .B(n51219), .A(n45148), .Z(n45149) );
  NAND U56818 ( .A(n58497), .B(n45149), .Z(n45150) );
  NANDN U56819 ( .A(n45151), .B(n45150), .Z(n45153) );
  AND U56820 ( .A(n45153), .B(n45152), .Z(n45154) );
  NANDN U56821 ( .A(x[5964]), .B(y[5964]), .Z(n51220) );
  AND U56822 ( .A(n45154), .B(n51220), .Z(n45155) );
  OR U56823 ( .A(n45156), .B(n45155), .Z(n45157) );
  NAND U56824 ( .A(n45158), .B(n45157), .Z(n45159) );
  NANDN U56825 ( .A(n45160), .B(n45159), .Z(n45162) );
  NANDN U56826 ( .A(n45162), .B(n45161), .Z(n45163) );
  NAND U56827 ( .A(n45164), .B(n45163), .Z(n45165) );
  AND U56828 ( .A(n45166), .B(n45165), .Z(n45167) );
  ANDN U56829 ( .B(n58507), .A(n45167), .Z(n45168) );
  NAND U56830 ( .A(n51218), .B(n45168), .Z(n45169) );
  NANDN U56831 ( .A(n45170), .B(n45169), .Z(n45171) );
  AND U56832 ( .A(n45171), .B(n58511), .Z(n45172) );
  NANDN U56833 ( .A(x[5972]), .B(y[5972]), .Z(n58508) );
  NAND U56834 ( .A(n45172), .B(n58508), .Z(n45173) );
  AND U56835 ( .A(n45174), .B(n45173), .Z(n45175) );
  ANDN U56836 ( .B(n58514), .A(n45175), .Z(n45176) );
  NAND U56837 ( .A(n58512), .B(n45176), .Z(n45177) );
  NANDN U56838 ( .A(n45178), .B(n45177), .Z(n45179) );
  AND U56839 ( .A(n45179), .B(n51215), .Z(n45180) );
  NANDN U56840 ( .A(x[5976]), .B(y[5976]), .Z(n58515) );
  NAND U56841 ( .A(n45180), .B(n58515), .Z(n45181) );
  AND U56842 ( .A(n45182), .B(n45181), .Z(n45183) );
  ANDN U56843 ( .B(n58519), .A(n45183), .Z(n45184) );
  NAND U56844 ( .A(n51216), .B(n45184), .Z(n45185) );
  NANDN U56845 ( .A(n45186), .B(n45185), .Z(n45188) );
  IV U56846 ( .A(n45187), .Z(n58520) );
  AND U56847 ( .A(n45188), .B(n58520), .Z(n45189) );
  NANDN U56848 ( .A(n58518), .B(n45189), .Z(n45190) );
  NAND U56849 ( .A(n45191), .B(n45190), .Z(n45192) );
  NANDN U56850 ( .A(n58525), .B(n45192), .Z(n45193) );
  ANDN U56851 ( .B(y[5982]), .A(x[5982]), .Z(n58521) );
  OR U56852 ( .A(n45193), .B(n58521), .Z(n45194) );
  NAND U56853 ( .A(n45195), .B(n45194), .Z(n45196) );
  ANDN U56854 ( .B(n45196), .A(n51212), .Z(n45197) );
  NANDN U56855 ( .A(x[5984]), .B(y[5984]), .Z(n58527) );
  NAND U56856 ( .A(n45197), .B(n58527), .Z(n45198) );
  AND U56857 ( .A(n45199), .B(n45198), .Z(n45201) );
  NANDN U56858 ( .A(x[5986]), .B(y[5986]), .Z(n51213) );
  AND U56859 ( .A(n51213), .B(n58530), .Z(n45200) );
  NANDN U56860 ( .A(n45201), .B(n45200), .Z(n45202) );
  NANDN U56861 ( .A(n45203), .B(n45202), .Z(n45205) );
  IV U56862 ( .A(n45204), .Z(n58532) );
  AND U56863 ( .A(n45205), .B(n58532), .Z(n45206) );
  NANDN U56864 ( .A(x[5988]), .B(y[5988]), .Z(n58531) );
  NAND U56865 ( .A(n45206), .B(n58531), .Z(n45207) );
  AND U56866 ( .A(n45208), .B(n45207), .Z(n45209) );
  ANDN U56867 ( .B(n58535), .A(n45209), .Z(n45210) );
  NAND U56868 ( .A(n58533), .B(n45210), .Z(n45211) );
  NANDN U56869 ( .A(n45212), .B(n45211), .Z(n45213) );
  AND U56870 ( .A(n45213), .B(n51209), .Z(n45214) );
  NANDN U56871 ( .A(x[5992]), .B(y[5992]), .Z(n58536) );
  NAND U56872 ( .A(n45214), .B(n58536), .Z(n45215) );
  AND U56873 ( .A(n45216), .B(n45215), .Z(n45218) );
  NANDN U56874 ( .A(x[5994]), .B(y[5994]), .Z(n51210) );
  AND U56875 ( .A(n51210), .B(n58540), .Z(n45217) );
  NANDN U56876 ( .A(n45218), .B(n45217), .Z(n45219) );
  NANDN U56877 ( .A(n45220), .B(n45219), .Z(n45222) );
  IV U56878 ( .A(n45221), .Z(n58542) );
  AND U56879 ( .A(n45222), .B(n58542), .Z(n45223) );
  NANDN U56880 ( .A(x[5996]), .B(y[5996]), .Z(n58541) );
  NAND U56881 ( .A(n45223), .B(n58541), .Z(n45224) );
  AND U56882 ( .A(n45225), .B(n45224), .Z(n45228) );
  NANDN U56883 ( .A(x[5998]), .B(y[5998]), .Z(n58543) );
  IV U56884 ( .A(n45226), .Z(n58545) );
  AND U56885 ( .A(n58543), .B(n58545), .Z(n45227) );
  NANDN U56886 ( .A(n45228), .B(n45227), .Z(n45229) );
  NANDN U56887 ( .A(n45230), .B(n45229), .Z(n45231) );
  AND U56888 ( .A(n51206), .B(n45231), .Z(n45232) );
  NANDN U56889 ( .A(x[6000]), .B(y[6000]), .Z(n58546) );
  NAND U56890 ( .A(n45232), .B(n58546), .Z(n45233) );
  AND U56891 ( .A(n45234), .B(n45233), .Z(n45236) );
  NANDN U56892 ( .A(x[6002]), .B(y[6002]), .Z(n51207) );
  AND U56893 ( .A(n51207), .B(n58549), .Z(n45235) );
  NANDN U56894 ( .A(n45236), .B(n45235), .Z(n45237) );
  NANDN U56895 ( .A(n45238), .B(n45237), .Z(n45240) );
  IV U56896 ( .A(n45239), .Z(n58553) );
  AND U56897 ( .A(n45240), .B(n58553), .Z(n45241) );
  NANDN U56898 ( .A(x[6004]), .B(y[6004]), .Z(n58550) );
  NAND U56899 ( .A(n45241), .B(n58550), .Z(n45242) );
  AND U56900 ( .A(n45243), .B(n45242), .Z(n45246) );
  NANDN U56901 ( .A(x[6006]), .B(y[6006]), .Z(n58554) );
  IV U56902 ( .A(n45244), .Z(n58556) );
  AND U56903 ( .A(n58554), .B(n58556), .Z(n45245) );
  NANDN U56904 ( .A(n45246), .B(n45245), .Z(n45247) );
  NANDN U56905 ( .A(n45248), .B(n45247), .Z(n45249) );
  AND U56906 ( .A(n51203), .B(n45249), .Z(n45250) );
  NANDN U56907 ( .A(x[6008]), .B(y[6008]), .Z(n58557) );
  NAND U56908 ( .A(n45250), .B(n58557), .Z(n45251) );
  AND U56909 ( .A(n45252), .B(n45251), .Z(n45254) );
  NANDN U56910 ( .A(x[6010]), .B(y[6010]), .Z(n51204) );
  AND U56911 ( .A(n51204), .B(n58560), .Z(n45253) );
  NANDN U56912 ( .A(n45254), .B(n45253), .Z(n45255) );
  NANDN U56913 ( .A(n45256), .B(n45255), .Z(n45258) );
  IV U56914 ( .A(n45257), .Z(n58562) );
  AND U56915 ( .A(n45258), .B(n58562), .Z(n45259) );
  NANDN U56916 ( .A(x[6012]), .B(y[6012]), .Z(n58561) );
  NAND U56917 ( .A(n45259), .B(n58561), .Z(n45260) );
  AND U56918 ( .A(n45261), .B(n45260), .Z(n45264) );
  NANDN U56919 ( .A(x[6014]), .B(y[6014]), .Z(n58563) );
  IV U56920 ( .A(n45262), .Z(n58566) );
  AND U56921 ( .A(n58563), .B(n58566), .Z(n45263) );
  NANDN U56922 ( .A(n45264), .B(n45263), .Z(n45265) );
  NANDN U56923 ( .A(n45266), .B(n45265), .Z(n45267) );
  AND U56924 ( .A(n51200), .B(n45267), .Z(n45268) );
  NANDN U56925 ( .A(x[6016]), .B(y[6016]), .Z(n58567) );
  NAND U56926 ( .A(n45268), .B(n58567), .Z(n45269) );
  NAND U56927 ( .A(n45270), .B(n45269), .Z(n45271) );
  AND U56928 ( .A(n45271), .B(n58571), .Z(n45272) );
  NANDN U56929 ( .A(x[6018]), .B(y[6018]), .Z(n51201) );
  AND U56930 ( .A(n45272), .B(n51201), .Z(n45273) );
  NOR U56931 ( .A(n45274), .B(n45273), .Z(n45276) );
  NAND U56932 ( .A(n45276), .B(n45275), .Z(n45278) );
  AND U56933 ( .A(n45278), .B(n45277), .Z(n45279) );
  NANDN U56934 ( .A(x[6020]), .B(y[6020]), .Z(n58570) );
  AND U56935 ( .A(n45279), .B(n58570), .Z(n45280) );
  OR U56936 ( .A(n45281), .B(n45280), .Z(n45282) );
  NAND U56937 ( .A(n45283), .B(n45282), .Z(n45284) );
  NANDN U56938 ( .A(n45285), .B(n45284), .Z(n45286) );
  AND U56939 ( .A(n45286), .B(n58580), .Z(n45287) );
  NANDN U56940 ( .A(x[6024]), .B(y[6024]), .Z(n51199) );
  NAND U56941 ( .A(n45287), .B(n51199), .Z(n45288) );
  AND U56942 ( .A(n45289), .B(n45288), .Z(n45290) );
  ANDN U56943 ( .B(n58582), .A(n45290), .Z(n45291) );
  NAND U56944 ( .A(n58578), .B(n45291), .Z(n45292) );
  NANDN U56945 ( .A(n45293), .B(n45292), .Z(n45294) );
  AND U56946 ( .A(n45294), .B(n58585), .Z(n45295) );
  NANDN U56947 ( .A(x[6028]), .B(y[6028]), .Z(n58583) );
  NAND U56948 ( .A(n45295), .B(n58583), .Z(n45296) );
  NAND U56949 ( .A(n45297), .B(n45296), .Z(n45298) );
  AND U56950 ( .A(n45298), .B(n51196), .Z(n45299) );
  NANDN U56951 ( .A(x[6030]), .B(y[6030]), .Z(n58586) );
  AND U56952 ( .A(n45299), .B(n58586), .Z(n45300) );
  NOR U56953 ( .A(n45301), .B(n45300), .Z(n45303) );
  NAND U56954 ( .A(n45303), .B(n45302), .Z(n45304) );
  AND U56955 ( .A(n45304), .B(n58590), .Z(n45305) );
  NANDN U56956 ( .A(x[6032]), .B(y[6032]), .Z(n51197) );
  NAND U56957 ( .A(n45305), .B(n51197), .Z(n45306) );
  AND U56958 ( .A(n45307), .B(n45306), .Z(n45308) );
  ANDN U56959 ( .B(n58592), .A(n45308), .Z(n45309) );
  NAND U56960 ( .A(n58589), .B(n45309), .Z(n45310) );
  NANDN U56961 ( .A(n45311), .B(n45310), .Z(n45313) );
  AND U56962 ( .A(n45313), .B(n45312), .Z(n45314) );
  NANDN U56963 ( .A(x[6036]), .B(y[6036]), .Z(n51195) );
  AND U56964 ( .A(n45314), .B(n51195), .Z(n45318) );
  AND U56965 ( .A(n45316), .B(n45315), .Z(n45317) );
  NANDN U56966 ( .A(n45318), .B(n45317), .Z(n45319) );
  NANDN U56967 ( .A(n45320), .B(n45319), .Z(n45321) );
  AND U56968 ( .A(n45322), .B(n45321), .Z(n45324) );
  NAND U56969 ( .A(n45324), .B(n45323), .Z(n45325) );
  AND U56970 ( .A(n45325), .B(n58600), .Z(n45326) );
  NANDN U56971 ( .A(x[6040]), .B(y[6040]), .Z(n58597) );
  NAND U56972 ( .A(n45326), .B(n58597), .Z(n45327) );
  AND U56973 ( .A(n45328), .B(n45327), .Z(n45329) );
  ANDN U56974 ( .B(n58603), .A(n45329), .Z(n45330) );
  NAND U56975 ( .A(n58601), .B(n45330), .Z(n45331) );
  NANDN U56976 ( .A(n45332), .B(n45331), .Z(n45333) );
  AND U56977 ( .A(n45333), .B(n51193), .Z(n45334) );
  NANDN U56978 ( .A(x[6044]), .B(y[6044]), .Z(n58604) );
  NAND U56979 ( .A(n45334), .B(n58604), .Z(n45335) );
  AND U56980 ( .A(n45336), .B(n45335), .Z(n45337) );
  ANDN U56981 ( .B(n58608), .A(n45337), .Z(n45338) );
  NAND U56982 ( .A(n51194), .B(n45338), .Z(n45339) );
  NANDN U56983 ( .A(n45340), .B(n45339), .Z(n45342) );
  AND U56984 ( .A(n45342), .B(n45341), .Z(n45343) );
  NANDN U56985 ( .A(x[6048]), .B(y[6048]), .Z(n58607) );
  AND U56986 ( .A(n45343), .B(n58607), .Z(n45344) );
  OR U56987 ( .A(n45345), .B(n45344), .Z(n45346) );
  NAND U56988 ( .A(n45347), .B(n45346), .Z(n45348) );
  NANDN U56989 ( .A(n45349), .B(n45348), .Z(n45350) );
  AND U56990 ( .A(n45351), .B(n45350), .Z(n45352) );
  OR U56991 ( .A(n45353), .B(n45352), .Z(n45354) );
  NAND U56992 ( .A(n45355), .B(n45354), .Z(n45356) );
  NANDN U56993 ( .A(n45357), .B(n45356), .Z(n45358) );
  AND U56994 ( .A(n45358), .B(n51191), .Z(n45359) );
  NANDN U56995 ( .A(x[6056]), .B(y[6056]), .Z(n58618) );
  NAND U56996 ( .A(n45359), .B(n58618), .Z(n45360) );
  AND U56997 ( .A(n45361), .B(n45360), .Z(n45362) );
  ANDN U56998 ( .B(n45363), .A(n45362), .Z(n45364) );
  NAND U56999 ( .A(n51192), .B(n45364), .Z(n45365) );
  NANDN U57000 ( .A(n45366), .B(n45365), .Z(n45367) );
  AND U57001 ( .A(n45368), .B(n45367), .Z(n45369) );
  OR U57002 ( .A(n45370), .B(n45369), .Z(n45371) );
  NAND U57003 ( .A(n45372), .B(n45371), .Z(n45373) );
  NANDN U57004 ( .A(n45374), .B(n45373), .Z(n45376) );
  AND U57005 ( .A(n45376), .B(n45375), .Z(n45377) );
  NANDN U57006 ( .A(x[6064]), .B(y[6064]), .Z(n51190) );
  AND U57007 ( .A(n45377), .B(n51190), .Z(n45378) );
  OR U57008 ( .A(n45379), .B(n45378), .Z(n45380) );
  NAND U57009 ( .A(n45381), .B(n45380), .Z(n45382) );
  NANDN U57010 ( .A(n45383), .B(n45382), .Z(n45384) );
  NAND U57011 ( .A(n45385), .B(n45384), .Z(n45386) );
  NAND U57012 ( .A(n45387), .B(n45386), .Z(n45389) );
  NANDN U57013 ( .A(x[6070]), .B(y[6070]), .Z(n51188) );
  AND U57014 ( .A(n58633), .B(n51188), .Z(n45388) );
  NAND U57015 ( .A(n45389), .B(n45388), .Z(n45390) );
  NANDN U57016 ( .A(n45391), .B(n45390), .Z(n45392) );
  AND U57017 ( .A(n45392), .B(n58635), .Z(n45393) );
  NANDN U57018 ( .A(x[6072]), .B(y[6072]), .Z(n58632) );
  AND U57019 ( .A(n45393), .B(n58632), .Z(n45394) );
  OR U57020 ( .A(n45395), .B(n45394), .Z(n45396) );
  NAND U57021 ( .A(n45397), .B(n45396), .Z(n45398) );
  NANDN U57022 ( .A(n45399), .B(n45398), .Z(n45400) );
  AND U57023 ( .A(n45400), .B(n51185), .Z(n45401) );
  NANDN U57024 ( .A(x[6076]), .B(y[6076]), .Z(n58639) );
  NAND U57025 ( .A(n45401), .B(n58639), .Z(n45402) );
  NAND U57026 ( .A(n45403), .B(n45402), .Z(n45405) );
  NANDN U57027 ( .A(x[6078]), .B(y[6078]), .Z(n51186) );
  AND U57028 ( .A(n51186), .B(n58644), .Z(n45404) );
  NAND U57029 ( .A(n45405), .B(n45404), .Z(n45406) );
  NANDN U57030 ( .A(n45407), .B(n45406), .Z(n45408) );
  AND U57031 ( .A(n45408), .B(n58648), .Z(n45409) );
  NANDN U57032 ( .A(x[6080]), .B(y[6080]), .Z(n58646) );
  NAND U57033 ( .A(n45409), .B(n58646), .Z(n45410) );
  AND U57034 ( .A(n45411), .B(n45410), .Z(n45412) );
  ANDN U57035 ( .B(n58651), .A(n45412), .Z(n45413) );
  NAND U57036 ( .A(n58649), .B(n45413), .Z(n45414) );
  NANDN U57037 ( .A(n45415), .B(n45414), .Z(n45416) );
  AND U57038 ( .A(n45416), .B(n51183), .Z(n45417) );
  NANDN U57039 ( .A(x[6084]), .B(y[6084]), .Z(n58652) );
  NAND U57040 ( .A(n45417), .B(n58652), .Z(n45418) );
  AND U57041 ( .A(n45419), .B(n45418), .Z(n45420) );
  ANDN U57042 ( .B(n58656), .A(n45420), .Z(n45421) );
  NAND U57043 ( .A(n51184), .B(n45421), .Z(n45422) );
  NANDN U57044 ( .A(n45423), .B(n45422), .Z(n45424) );
  AND U57045 ( .A(n45424), .B(n58658), .Z(n45425) );
  NANDN U57046 ( .A(x[6088]), .B(y[6088]), .Z(n58655) );
  NAND U57047 ( .A(n45425), .B(n58655), .Z(n45426) );
  AND U57048 ( .A(n45427), .B(n45426), .Z(n45428) );
  ANDN U57049 ( .B(n58662), .A(n45428), .Z(n45429) );
  NAND U57050 ( .A(n58659), .B(n45429), .Z(n45430) );
  NANDN U57051 ( .A(n45431), .B(n45430), .Z(n45432) );
  AND U57052 ( .A(n45432), .B(n51181), .Z(n45433) );
  NANDN U57053 ( .A(x[6092]), .B(y[6092]), .Z(n58663) );
  AND U57054 ( .A(n45433), .B(n58663), .Z(n45434) );
  OR U57055 ( .A(n45435), .B(n45434), .Z(n45436) );
  NAND U57056 ( .A(n45437), .B(n45436), .Z(n45441) );
  ANDN U57057 ( .B(n45439), .A(n45438), .Z(n45440) );
  NAND U57058 ( .A(n45441), .B(n45440), .Z(n45442) );
  AND U57059 ( .A(n58666), .B(n45442), .Z(n45443) );
  NANDN U57060 ( .A(x[6096]), .B(y[6096]), .Z(n51180) );
  NAND U57061 ( .A(n45443), .B(n51180), .Z(n45444) );
  AND U57062 ( .A(n45445), .B(n45444), .Z(n45447) );
  NANDN U57063 ( .A(x[6098]), .B(y[6098]), .Z(n58667) );
  AND U57064 ( .A(n58667), .B(n58669), .Z(n45446) );
  NANDN U57065 ( .A(n45447), .B(n45446), .Z(n45448) );
  NANDN U57066 ( .A(n45449), .B(n45448), .Z(n45450) );
  AND U57067 ( .A(n51176), .B(n45450), .Z(n45451) );
  NANDN U57068 ( .A(x[6100]), .B(y[6100]), .Z(n58670) );
  NAND U57069 ( .A(n45451), .B(n58670), .Z(n45452) );
  AND U57070 ( .A(n45453), .B(n45452), .Z(n45455) );
  NANDN U57071 ( .A(x[6102]), .B(y[6102]), .Z(n51177) );
  AND U57072 ( .A(n51177), .B(n58674), .Z(n45454) );
  NANDN U57073 ( .A(n45455), .B(n45454), .Z(n45456) );
  NANDN U57074 ( .A(n45457), .B(n45456), .Z(n45458) );
  AND U57075 ( .A(n58678), .B(n45458), .Z(n45459) );
  NANDN U57076 ( .A(x[6104]), .B(y[6104]), .Z(n58673) );
  NAND U57077 ( .A(n45459), .B(n58673), .Z(n45460) );
  AND U57078 ( .A(n45461), .B(n45460), .Z(n45463) );
  NANDN U57079 ( .A(x[6106]), .B(y[6106]), .Z(n58679) );
  AND U57080 ( .A(n58679), .B(n58680), .Z(n45462) );
  NANDN U57081 ( .A(n45463), .B(n45462), .Z(n45464) );
  NANDN U57082 ( .A(n45465), .B(n45464), .Z(n45467) );
  IV U57083 ( .A(n45466), .Z(n51173) );
  AND U57084 ( .A(n45467), .B(n51173), .Z(n45468) );
  NANDN U57085 ( .A(x[6108]), .B(y[6108]), .Z(n58681) );
  NAND U57086 ( .A(n45468), .B(n58681), .Z(n45469) );
  AND U57087 ( .A(n45470), .B(n45469), .Z(n45472) );
  NANDN U57088 ( .A(x[6110]), .B(y[6110]), .Z(n51174) );
  AND U57089 ( .A(n51174), .B(n58685), .Z(n45471) );
  NANDN U57090 ( .A(n45472), .B(n45471), .Z(n45473) );
  NANDN U57091 ( .A(n45474), .B(n45473), .Z(n45475) );
  AND U57092 ( .A(n58687), .B(n45475), .Z(n45476) );
  NANDN U57093 ( .A(x[6112]), .B(y[6112]), .Z(n58684) );
  NAND U57094 ( .A(n45476), .B(n58684), .Z(n45477) );
  AND U57095 ( .A(n45478), .B(n45477), .Z(n45480) );
  NANDN U57096 ( .A(x[6114]), .B(y[6114]), .Z(n58688) );
  AND U57097 ( .A(n58688), .B(n58691), .Z(n45479) );
  NANDN U57098 ( .A(n45480), .B(n45479), .Z(n45481) );
  NANDN U57099 ( .A(n45482), .B(n45481), .Z(n45483) );
  AND U57100 ( .A(n51171), .B(n45483), .Z(n45484) );
  NANDN U57101 ( .A(x[6116]), .B(y[6116]), .Z(n58692) );
  NAND U57102 ( .A(n45484), .B(n58692), .Z(n45485) );
  AND U57103 ( .A(n45486), .B(n45485), .Z(n45488) );
  NANDN U57104 ( .A(x[6118]), .B(y[6118]), .Z(n51172) );
  AND U57105 ( .A(n51172), .B(n58696), .Z(n45487) );
  NANDN U57106 ( .A(n45488), .B(n45487), .Z(n45489) );
  NANDN U57107 ( .A(n45490), .B(n45489), .Z(n45491) );
  AND U57108 ( .A(n58698), .B(n45491), .Z(n45492) );
  NANDN U57109 ( .A(x[6120]), .B(y[6120]), .Z(n58695) );
  NAND U57110 ( .A(n45492), .B(n58695), .Z(n45493) );
  AND U57111 ( .A(n45494), .B(n45493), .Z(n45495) );
  NOR U57112 ( .A(n58699), .B(n45495), .Z(n45496) );
  NAND U57113 ( .A(n45497), .B(n45496), .Z(n45498) );
  NANDN U57114 ( .A(n45499), .B(n45498), .Z(n45501) );
  OR U57115 ( .A(n45501), .B(n45500), .Z(n45502) );
  AND U57116 ( .A(n58704), .B(n45502), .Z(n45504) );
  NANDN U57117 ( .A(x[6124]), .B(y[6124]), .Z(n45503) );
  NAND U57118 ( .A(n45504), .B(n45503), .Z(n45505) );
  AND U57119 ( .A(n45506), .B(n45505), .Z(n45509) );
  NANDN U57120 ( .A(x[6126]), .B(y[6126]), .Z(n58703) );
  IV U57121 ( .A(n45507), .Z(n58705) );
  AND U57122 ( .A(n58703), .B(n58705), .Z(n45508) );
  NANDN U57123 ( .A(n45509), .B(n45508), .Z(n45510) );
  NANDN U57124 ( .A(n45511), .B(n45510), .Z(n45512) );
  AND U57125 ( .A(n58709), .B(n45512), .Z(n45513) );
  NANDN U57126 ( .A(x[6128]), .B(y[6128]), .Z(n58706) );
  NAND U57127 ( .A(n45513), .B(n58706), .Z(n45514) );
  AND U57128 ( .A(n45515), .B(n45514), .Z(n45517) );
  NANDN U57129 ( .A(x[6130]), .B(y[6130]), .Z(n58710) );
  AND U57130 ( .A(n58710), .B(n51168), .Z(n45516) );
  NANDN U57131 ( .A(n45517), .B(n45516), .Z(n45518) );
  NANDN U57132 ( .A(n45519), .B(n45518), .Z(n45520) );
  AND U57133 ( .A(n58714), .B(n45520), .Z(n45521) );
  NANDN U57134 ( .A(x[6132]), .B(y[6132]), .Z(n51169) );
  NAND U57135 ( .A(n45521), .B(n51169), .Z(n45522) );
  AND U57136 ( .A(n45523), .B(n45522), .Z(n45526) );
  NANDN U57137 ( .A(x[6134]), .B(y[6134]), .Z(n58713) );
  IV U57138 ( .A(n45524), .Z(n58715) );
  AND U57139 ( .A(n58713), .B(n58715), .Z(n45525) );
  NANDN U57140 ( .A(n45526), .B(n45525), .Z(n45527) );
  NANDN U57141 ( .A(n45528), .B(n45527), .Z(n45530) );
  IV U57142 ( .A(n45529), .Z(n58718) );
  AND U57143 ( .A(n45530), .B(n58718), .Z(n45531) );
  NANDN U57144 ( .A(x[6136]), .B(y[6136]), .Z(n58716) );
  NAND U57145 ( .A(n45531), .B(n58716), .Z(n45532) );
  AND U57146 ( .A(n45533), .B(n45532), .Z(n45534) );
  OR U57147 ( .A(n45535), .B(n45534), .Z(n45536) );
  NAND U57148 ( .A(n45537), .B(n45536), .Z(n45538) );
  NANDN U57149 ( .A(n58724), .B(n45538), .Z(n45540) );
  ANDN U57150 ( .B(y[6140]), .A(x[6140]), .Z(n45539) );
  OR U57151 ( .A(n45540), .B(n45539), .Z(n45541) );
  NAND U57152 ( .A(n45542), .B(n45541), .Z(n45543) );
  NANDN U57153 ( .A(n58728), .B(n45543), .Z(n45544) );
  ANDN U57154 ( .B(y[6142]), .A(x[6142]), .Z(n58723) );
  OR U57155 ( .A(n45544), .B(n58723), .Z(n45545) );
  NAND U57156 ( .A(n45546), .B(n45545), .Z(n45547) );
  NANDN U57157 ( .A(n45548), .B(n45547), .Z(n45549) );
  NAND U57158 ( .A(n45550), .B(n45549), .Z(n45551) );
  NAND U57159 ( .A(n45552), .B(n45551), .Z(n45553) );
  NAND U57160 ( .A(n45554), .B(n45553), .Z(n45555) );
  ANDN U57161 ( .B(y[6148]), .A(x[6148]), .Z(n58731) );
  ANDN U57162 ( .B(n45555), .A(n58731), .Z(n45556) );
  NANDN U57163 ( .A(n58733), .B(n45556), .Z(n45557) );
  NAND U57164 ( .A(n45558), .B(n45557), .Z(n45559) );
  AND U57165 ( .A(n45559), .B(n58736), .Z(n45560) );
  NANDN U57166 ( .A(x[6150]), .B(y[6150]), .Z(n58734) );
  AND U57167 ( .A(n45560), .B(n58734), .Z(n45564) );
  AND U57168 ( .A(n45562), .B(n45561), .Z(n45563) );
  NANDN U57169 ( .A(n45564), .B(n45563), .Z(n45565) );
  NAND U57170 ( .A(n45566), .B(n45565), .Z(n45567) );
  NAND U57171 ( .A(n45568), .B(n45567), .Z(n45569) );
  AND U57172 ( .A(n45569), .B(n58742), .Z(n45570) );
  NANDN U57173 ( .A(x[6154]), .B(y[6154]), .Z(n51163) );
  AND U57174 ( .A(n45570), .B(n51163), .Z(n45574) );
  AND U57175 ( .A(n45572), .B(n45571), .Z(n45573) );
  NANDN U57176 ( .A(n45574), .B(n45573), .Z(n45575) );
  NAND U57177 ( .A(n45576), .B(n45575), .Z(n45577) );
  NAND U57178 ( .A(n45578), .B(n45577), .Z(n45579) );
  AND U57179 ( .A(n45579), .B(n58746), .Z(n45580) );
  NANDN U57180 ( .A(x[6158]), .B(y[6158]), .Z(n58744) );
  AND U57181 ( .A(n45580), .B(n58744), .Z(n45584) );
  AND U57182 ( .A(n45582), .B(n45581), .Z(n45583) );
  NANDN U57183 ( .A(n45584), .B(n45583), .Z(n45585) );
  NAND U57184 ( .A(n45586), .B(n45585), .Z(n45587) );
  NAND U57185 ( .A(n45588), .B(n45587), .Z(n45590) );
  AND U57186 ( .A(n45590), .B(n45589), .Z(n45591) );
  NAND U57187 ( .A(n51160), .B(n45591), .Z(n45592) );
  NAND U57188 ( .A(n45593), .B(n45592), .Z(n45594) );
  NANDN U57189 ( .A(n45595), .B(n45594), .Z(n45596) );
  AND U57190 ( .A(n45597), .B(n45596), .Z(n45598) );
  OR U57191 ( .A(n45599), .B(n45598), .Z(n45600) );
  NAND U57192 ( .A(n45601), .B(n45600), .Z(n45602) );
  NANDN U57193 ( .A(n45603), .B(n45602), .Z(n45604) );
  AND U57194 ( .A(n45605), .B(n45604), .Z(n45606) );
  ANDN U57195 ( .B(n58758), .A(n45606), .Z(n45607) );
  NANDN U57196 ( .A(x[6170]), .B(y[6170]), .Z(n58756) );
  AND U57197 ( .A(n45607), .B(n58756), .Z(n45608) );
  OR U57198 ( .A(n45609), .B(n45608), .Z(n45610) );
  NAND U57199 ( .A(n45611), .B(n45610), .Z(n45612) );
  NAND U57200 ( .A(n45613), .B(n45612), .Z(n45614) );
  AND U57201 ( .A(n45614), .B(n51155), .Z(n45615) );
  NANDN U57202 ( .A(x[6174]), .B(y[6174]), .Z(n58762) );
  AND U57203 ( .A(n45615), .B(n58762), .Z(n45619) );
  AND U57204 ( .A(n45617), .B(n45616), .Z(n45618) );
  NANDN U57205 ( .A(n45619), .B(n45618), .Z(n45620) );
  NAND U57206 ( .A(n45621), .B(n45620), .Z(n45622) );
  NAND U57207 ( .A(n45623), .B(n45622), .Z(n45625) );
  IV U57208 ( .A(n45624), .Z(n58771) );
  AND U57209 ( .A(n45625), .B(n58771), .Z(n45626) );
  NANDN U57210 ( .A(x[6178]), .B(y[6178]), .Z(n58768) );
  AND U57211 ( .A(n45626), .B(n58768), .Z(n45630) );
  AND U57212 ( .A(n45628), .B(n45627), .Z(n45629) );
  NANDN U57213 ( .A(n45630), .B(n45629), .Z(n45631) );
  NAND U57214 ( .A(n45632), .B(n45631), .Z(n45633) );
  NAND U57215 ( .A(n45634), .B(n45633), .Z(n45635) );
  AND U57216 ( .A(n45635), .B(n51152), .Z(n45636) );
  NANDN U57217 ( .A(x[6182]), .B(y[6182]), .Z(n58775) );
  AND U57218 ( .A(n45636), .B(n58775), .Z(n45640) );
  AND U57219 ( .A(n45638), .B(n45637), .Z(n45639) );
  NANDN U57220 ( .A(n45640), .B(n45639), .Z(n45641) );
  NAND U57221 ( .A(n45642), .B(n45641), .Z(n45643) );
  NAND U57222 ( .A(n45644), .B(n45643), .Z(n45646) );
  IV U57223 ( .A(n45645), .Z(n58781) );
  AND U57224 ( .A(n45646), .B(n58781), .Z(n45647) );
  NANDN U57225 ( .A(x[6186]), .B(y[6186]), .Z(n58778) );
  AND U57226 ( .A(n45647), .B(n58778), .Z(n45651) );
  AND U57227 ( .A(n45649), .B(n45648), .Z(n45650) );
  NANDN U57228 ( .A(n45651), .B(n45650), .Z(n45652) );
  NAND U57229 ( .A(n45653), .B(n45652), .Z(n45654) );
  NAND U57230 ( .A(n45655), .B(n45654), .Z(n45656) );
  AND U57231 ( .A(n45656), .B(n51149), .Z(n45657) );
  NANDN U57232 ( .A(x[6190]), .B(y[6190]), .Z(n58785) );
  AND U57233 ( .A(n45657), .B(n58785), .Z(n45661) );
  AND U57234 ( .A(n45659), .B(n45658), .Z(n45660) );
  NANDN U57235 ( .A(n45661), .B(n45660), .Z(n45662) );
  NAND U57236 ( .A(n45663), .B(n45662), .Z(n45664) );
  NAND U57237 ( .A(n45665), .B(n45664), .Z(n45667) );
  IV U57238 ( .A(n45666), .Z(n58790) );
  AND U57239 ( .A(n45667), .B(n58790), .Z(n45668) );
  NANDN U57240 ( .A(x[6194]), .B(y[6194]), .Z(n58788) );
  AND U57241 ( .A(n45668), .B(n58788), .Z(n45672) );
  AND U57242 ( .A(n45670), .B(n45669), .Z(n45671) );
  NANDN U57243 ( .A(n45672), .B(n45671), .Z(n45673) );
  NAND U57244 ( .A(n45674), .B(n45673), .Z(n45675) );
  NAND U57245 ( .A(n45676), .B(n45675), .Z(n45677) );
  AND U57246 ( .A(n45677), .B(n51145), .Z(n45678) );
  NANDN U57247 ( .A(x[6198]), .B(y[6198]), .Z(n58794) );
  AND U57248 ( .A(n45678), .B(n58794), .Z(n45682) );
  AND U57249 ( .A(n45680), .B(n45679), .Z(n45681) );
  NANDN U57250 ( .A(n45682), .B(n45681), .Z(n45683) );
  NAND U57251 ( .A(n45684), .B(n45683), .Z(n45685) );
  NAND U57252 ( .A(n45686), .B(n45685), .Z(n45688) );
  IV U57253 ( .A(n45687), .Z(n58799) );
  AND U57254 ( .A(n45688), .B(n58799), .Z(n45689) );
  NANDN U57255 ( .A(x[6202]), .B(y[6202]), .Z(n58797) );
  AND U57256 ( .A(n45689), .B(n58797), .Z(n45693) );
  AND U57257 ( .A(n45691), .B(n45690), .Z(n45692) );
  NANDN U57258 ( .A(n45693), .B(n45692), .Z(n45694) );
  NAND U57259 ( .A(n45695), .B(n45694), .Z(n45696) );
  NAND U57260 ( .A(n45697), .B(n45696), .Z(n45698) );
  AND U57261 ( .A(n45698), .B(n51141), .Z(n45699) );
  NANDN U57262 ( .A(x[6206]), .B(y[6206]), .Z(n58802) );
  AND U57263 ( .A(n45699), .B(n58802), .Z(n45703) );
  AND U57264 ( .A(n45701), .B(n45700), .Z(n45702) );
  NANDN U57265 ( .A(n45703), .B(n45702), .Z(n45704) );
  NAND U57266 ( .A(n45705), .B(n45704), .Z(n45706) );
  NAND U57267 ( .A(n45707), .B(n45706), .Z(n45709) );
  IV U57268 ( .A(n45708), .Z(n58807) );
  AND U57269 ( .A(n45709), .B(n58807), .Z(n45710) );
  NANDN U57270 ( .A(x[6210]), .B(y[6210]), .Z(n58806) );
  AND U57271 ( .A(n45710), .B(n58806), .Z(n45714) );
  AND U57272 ( .A(n45712), .B(n45711), .Z(n45713) );
  NANDN U57273 ( .A(n45714), .B(n45713), .Z(n45715) );
  NAND U57274 ( .A(n45716), .B(n45715), .Z(n45717) );
  NAND U57275 ( .A(n45718), .B(n45717), .Z(n45719) );
  AND U57276 ( .A(n45719), .B(n51137), .Z(n45720) );
  NANDN U57277 ( .A(x[6214]), .B(y[6214]), .Z(n58811) );
  AND U57278 ( .A(n45720), .B(n58811), .Z(n45724) );
  AND U57279 ( .A(n45722), .B(n45721), .Z(n45723) );
  NANDN U57280 ( .A(n45724), .B(n45723), .Z(n45725) );
  NAND U57281 ( .A(n45726), .B(n45725), .Z(n45727) );
  NAND U57282 ( .A(n45728), .B(n45727), .Z(n45730) );
  IV U57283 ( .A(n45729), .Z(n58818) );
  AND U57284 ( .A(n45730), .B(n58818), .Z(n45731) );
  NANDN U57285 ( .A(x[6218]), .B(y[6218]), .Z(n58815) );
  AND U57286 ( .A(n45731), .B(n58815), .Z(n45735) );
  AND U57287 ( .A(n45733), .B(n45732), .Z(n45734) );
  NANDN U57288 ( .A(n45735), .B(n45734), .Z(n45736) );
  NAND U57289 ( .A(n45737), .B(n45736), .Z(n45738) );
  AND U57290 ( .A(n45739), .B(n45738), .Z(n45740) );
  ANDN U57291 ( .B(n45741), .A(n45740), .Z(n45742) );
  OR U57292 ( .A(n45743), .B(n45742), .Z(n45744) );
  NAND U57293 ( .A(n45745), .B(n45744), .Z(n45746) );
  NAND U57294 ( .A(n45747), .B(n45746), .Z(n45748) );
  AND U57295 ( .A(n45748), .B(n58827), .Z(n45750) );
  NANDN U57296 ( .A(x[6226]), .B(y[6226]), .Z(n45749) );
  AND U57297 ( .A(n45750), .B(n45749), .Z(n45754) );
  AND U57298 ( .A(n45752), .B(n45751), .Z(n45753) );
  NANDN U57299 ( .A(n45754), .B(n45753), .Z(n45755) );
  NAND U57300 ( .A(n45756), .B(n45755), .Z(n45757) );
  NAND U57301 ( .A(n45758), .B(n45757), .Z(n45759) );
  AND U57302 ( .A(n45759), .B(n58834), .Z(n45760) );
  NANDN U57303 ( .A(x[6230]), .B(y[6230]), .Z(n51132) );
  AND U57304 ( .A(n45760), .B(n51132), .Z(n45764) );
  AND U57305 ( .A(n45762), .B(n45761), .Z(n45763) );
  NANDN U57306 ( .A(n45764), .B(n45763), .Z(n45765) );
  NAND U57307 ( .A(n45766), .B(n45765), .Z(n45767) );
  NAND U57308 ( .A(n45768), .B(n45767), .Z(n45769) );
  AND U57309 ( .A(n45769), .B(n58838), .Z(n45770) );
  NANDN U57310 ( .A(x[6234]), .B(y[6234]), .Z(n58836) );
  AND U57311 ( .A(n45770), .B(n58836), .Z(n45774) );
  AND U57312 ( .A(n45772), .B(n45771), .Z(n45773) );
  NANDN U57313 ( .A(n45774), .B(n45773), .Z(n45775) );
  NAND U57314 ( .A(n45776), .B(n45775), .Z(n45777) );
  AND U57315 ( .A(n45778), .B(n45777), .Z(n45779) );
  OR U57316 ( .A(n45780), .B(n45779), .Z(n45781) );
  NAND U57317 ( .A(n45782), .B(n45781), .Z(n45783) );
  NANDN U57318 ( .A(n45784), .B(n45783), .Z(n45785) );
  AND U57319 ( .A(n45786), .B(n45785), .Z(n45787) );
  OR U57320 ( .A(n45788), .B(n45787), .Z(n45789) );
  NAND U57321 ( .A(n45790), .B(n45789), .Z(n45791) );
  NANDN U57322 ( .A(n45792), .B(n45791), .Z(n45793) );
  NAND U57323 ( .A(n45794), .B(n45793), .Z(n45796) );
  IV U57324 ( .A(n45795), .Z(n51125) );
  AND U57325 ( .A(n45796), .B(n51125), .Z(n45797) );
  NANDN U57326 ( .A(x[6246]), .B(y[6246]), .Z(n58849) );
  AND U57327 ( .A(n45797), .B(n58849), .Z(n45798) );
  OR U57328 ( .A(n45799), .B(n45798), .Z(n45800) );
  NAND U57329 ( .A(n45801), .B(n45800), .Z(n45802) );
  AND U57330 ( .A(n45803), .B(n45802), .Z(n45804) );
  ANDN U57331 ( .B(n45805), .A(n45804), .Z(n45806) );
  OR U57332 ( .A(n45807), .B(n45806), .Z(n45808) );
  NAND U57333 ( .A(n45809), .B(n45808), .Z(n45810) );
  NAND U57334 ( .A(n45811), .B(n45810), .Z(n45812) );
  AND U57335 ( .A(n45812), .B(n58860), .Z(n45813) );
  NANDN U57336 ( .A(x[6254]), .B(y[6254]), .Z(n58857) );
  AND U57337 ( .A(n45813), .B(n58857), .Z(n45817) );
  AND U57338 ( .A(n45815), .B(n45814), .Z(n45816) );
  NANDN U57339 ( .A(n45817), .B(n45816), .Z(n45818) );
  NAND U57340 ( .A(n45819), .B(n45818), .Z(n45820) );
  NAND U57341 ( .A(n45821), .B(n45820), .Z(n45823) );
  IV U57342 ( .A(n45822), .Z(n51120) );
  AND U57343 ( .A(n45823), .B(n51120), .Z(n45824) );
  NANDN U57344 ( .A(n58864), .B(n45824), .Z(n45825) );
  NAND U57345 ( .A(n45826), .B(n45825), .Z(n45827) );
  NAND U57346 ( .A(n58870), .B(n45827), .Z(n45828) );
  NANDN U57347 ( .A(x[6260]), .B(y[6260]), .Z(n51121) );
  NANDN U57348 ( .A(n45828), .B(n51121), .Z(n45829) );
  AND U57349 ( .A(n45830), .B(n45829), .Z(n45831) );
  OR U57350 ( .A(n45832), .B(n45831), .Z(n45833) );
  NAND U57351 ( .A(n45834), .B(n45833), .Z(n45835) );
  NANDN U57352 ( .A(n45836), .B(n45835), .Z(n45837) );
  NAND U57353 ( .A(n45838), .B(n45837), .Z(n45839) );
  AND U57354 ( .A(n45840), .B(n45839), .Z(n45844) );
  XNOR U57355 ( .A(x[6268]), .B(y[6268]), .Z(n45842) );
  AND U57356 ( .A(n45842), .B(n45841), .Z(n45843) );
  NANDN U57357 ( .A(n45844), .B(n45843), .Z(n45845) );
  NAND U57358 ( .A(n45846), .B(n45845), .Z(n45847) );
  NAND U57359 ( .A(n45848), .B(n45847), .Z(n45849) );
  AND U57360 ( .A(n45849), .B(n58881), .Z(n45850) );
  NANDN U57361 ( .A(x[6270]), .B(y[6270]), .Z(n58879) );
  AND U57362 ( .A(n45850), .B(n58879), .Z(n45854) );
  AND U57363 ( .A(n45852), .B(n45851), .Z(n45853) );
  NANDN U57364 ( .A(n45854), .B(n45853), .Z(n45855) );
  NAND U57365 ( .A(n45856), .B(n45855), .Z(n45857) );
  NAND U57366 ( .A(n45858), .B(n45857), .Z(n45859) );
  AND U57367 ( .A(n45859), .B(n58887), .Z(n45860) );
  NANDN U57368 ( .A(x[6274]), .B(y[6274]), .Z(n51116) );
  AND U57369 ( .A(n45860), .B(n51116), .Z(n45864) );
  AND U57370 ( .A(n45862), .B(n45861), .Z(n45863) );
  NANDN U57371 ( .A(n45864), .B(n45863), .Z(n45865) );
  NAND U57372 ( .A(n45866), .B(n45865), .Z(n45867) );
  AND U57373 ( .A(n45868), .B(n45867), .Z(n45870) );
  NANDN U57374 ( .A(x[6278]), .B(y[6278]), .Z(n58890) );
  AND U57375 ( .A(n58890), .B(n58892), .Z(n45869) );
  NANDN U57376 ( .A(n45870), .B(n45869), .Z(n45871) );
  NAND U57377 ( .A(n45872), .B(n45871), .Z(n45873) );
  OR U57378 ( .A(n45874), .B(n45873), .Z(n45875) );
  NAND U57379 ( .A(n45876), .B(n45875), .Z(n45877) );
  NAND U57380 ( .A(n45878), .B(n45877), .Z(n45879) );
  AND U57381 ( .A(n45879), .B(n58898), .Z(n45880) );
  NANDN U57382 ( .A(x[6282]), .B(y[6282]), .Z(n51114) );
  AND U57383 ( .A(n45880), .B(n51114), .Z(n45884) );
  AND U57384 ( .A(n45882), .B(n45881), .Z(n45883) );
  NANDN U57385 ( .A(n45884), .B(n45883), .Z(n45885) );
  NAND U57386 ( .A(n45886), .B(n45885), .Z(n45887) );
  AND U57387 ( .A(n45888), .B(n45887), .Z(n45889) );
  OR U57388 ( .A(n45890), .B(n45889), .Z(n45891) );
  NAND U57389 ( .A(n45892), .B(n45891), .Z(n45893) );
  NAND U57390 ( .A(n45894), .B(n45893), .Z(n45895) );
  NAND U57391 ( .A(n45896), .B(n45895), .Z(n45897) );
  AND U57392 ( .A(n45897), .B(n58908), .Z(n45898) );
  NANDN U57393 ( .A(x[6290]), .B(y[6290]), .Z(n51112) );
  AND U57394 ( .A(n45898), .B(n51112), .Z(n45899) );
  OR U57395 ( .A(n45900), .B(n45899), .Z(n45901) );
  NAND U57396 ( .A(n45902), .B(n45901), .Z(n45903) );
  NAND U57397 ( .A(n45904), .B(n45903), .Z(n45905) );
  AND U57398 ( .A(n45905), .B(n58914), .Z(n45906) );
  NANDN U57399 ( .A(x[6294]), .B(y[6294]), .Z(n58911) );
  AND U57400 ( .A(n45906), .B(n58911), .Z(n45910) );
  AND U57401 ( .A(n45908), .B(n45907), .Z(n45909) );
  NANDN U57402 ( .A(n45910), .B(n45909), .Z(n45911) );
  NAND U57403 ( .A(n45912), .B(n45911), .Z(n45913) );
  AND U57404 ( .A(n45914), .B(n45913), .Z(n45915) );
  ANDN U57405 ( .B(n58919), .A(n45915), .Z(n45916) );
  NANDN U57406 ( .A(x[6298]), .B(y[6298]), .Z(n51110) );
  AND U57407 ( .A(n45916), .B(n51110), .Z(n45917) );
  OR U57408 ( .A(n45918), .B(n45917), .Z(n45919) );
  NAND U57409 ( .A(n45920), .B(n45919), .Z(n45921) );
  NAND U57410 ( .A(n45922), .B(n45921), .Z(n45923) );
  AND U57411 ( .A(n45923), .B(n58924), .Z(n45924) );
  NANDN U57412 ( .A(x[6302]), .B(y[6302]), .Z(n58922) );
  AND U57413 ( .A(n45924), .B(n58922), .Z(n45928) );
  AND U57414 ( .A(n45926), .B(n45925), .Z(n45927) );
  NANDN U57415 ( .A(n45928), .B(n45927), .Z(n45929) );
  NAND U57416 ( .A(n45930), .B(n45929), .Z(n45931) );
  NAND U57417 ( .A(n45932), .B(n45931), .Z(n45933) );
  AND U57418 ( .A(n45933), .B(n51106), .Z(n45934) );
  NANDN U57419 ( .A(x[6306]), .B(y[6306]), .Z(n51108) );
  AND U57420 ( .A(n45934), .B(n51108), .Z(n45938) );
  AND U57421 ( .A(n45936), .B(n45935), .Z(n45937) );
  NANDN U57422 ( .A(n45938), .B(n45937), .Z(n45939) );
  NAND U57423 ( .A(n45940), .B(n45939), .Z(n45941) );
  NAND U57424 ( .A(n45942), .B(n45941), .Z(n45944) );
  IV U57425 ( .A(n45943), .Z(n58933) );
  AND U57426 ( .A(n45944), .B(n58933), .Z(n45945) );
  NANDN U57427 ( .A(x[6310]), .B(y[6310]), .Z(n58931) );
  AND U57428 ( .A(n45945), .B(n58931), .Z(n45949) );
  AND U57429 ( .A(n45947), .B(n45946), .Z(n45948) );
  NANDN U57430 ( .A(n45949), .B(n45948), .Z(n45950) );
  NAND U57431 ( .A(n45951), .B(n45950), .Z(n45952) );
  NAND U57432 ( .A(n45953), .B(n45952), .Z(n45954) );
  AND U57433 ( .A(n45954), .B(n58938), .Z(n45955) );
  NANDN U57434 ( .A(x[6314]), .B(y[6314]), .Z(n51103) );
  AND U57435 ( .A(n45955), .B(n51103), .Z(n45959) );
  AND U57436 ( .A(n45957), .B(n45956), .Z(n45958) );
  NANDN U57437 ( .A(n45959), .B(n45958), .Z(n45960) );
  NAND U57438 ( .A(n45961), .B(n45960), .Z(n45962) );
  NAND U57439 ( .A(n45963), .B(n45962), .Z(n45964) );
  AND U57440 ( .A(n45964), .B(n58944), .Z(n45965) );
  NANDN U57441 ( .A(x[6318]), .B(y[6318]), .Z(n58942) );
  AND U57442 ( .A(n45965), .B(n58942), .Z(n45969) );
  AND U57443 ( .A(n45967), .B(n45966), .Z(n45968) );
  NANDN U57444 ( .A(n45969), .B(n45968), .Z(n45970) );
  NAND U57445 ( .A(n45971), .B(n45970), .Z(n45972) );
  NAND U57446 ( .A(n45973), .B(n45972), .Z(n45974) );
  AND U57447 ( .A(n45974), .B(n58949), .Z(n45975) );
  NANDN U57448 ( .A(x[6322]), .B(y[6322]), .Z(n51101) );
  AND U57449 ( .A(n45975), .B(n51101), .Z(n45979) );
  AND U57450 ( .A(n45977), .B(n45976), .Z(n45978) );
  NANDN U57451 ( .A(n45979), .B(n45978), .Z(n45980) );
  NAND U57452 ( .A(n45981), .B(n45980), .Z(n45982) );
  AND U57453 ( .A(n45983), .B(n45982), .Z(n45984) );
  ANDN U57454 ( .B(n45985), .A(n45984), .Z(n45986) );
  OR U57455 ( .A(n45987), .B(n45986), .Z(n45988) );
  NAND U57456 ( .A(n45989), .B(n45988), .Z(n45990) );
  AND U57457 ( .A(n45991), .B(n45990), .Z(n45992) );
  OR U57458 ( .A(n45993), .B(n45992), .Z(n45994) );
  NAND U57459 ( .A(n45995), .B(n45994), .Z(n45996) );
  NANDN U57460 ( .A(n45997), .B(n45996), .Z(n45998) );
  ANDN U57461 ( .B(n45999), .A(n45998), .Z(n46000) );
  OR U57462 ( .A(n46001), .B(n46000), .Z(n46002) );
  NAND U57463 ( .A(n46003), .B(n46002), .Z(n46004) );
  NANDN U57464 ( .A(n46005), .B(n46004), .Z(n46006) );
  OR U57465 ( .A(n46007), .B(n46006), .Z(n46008) );
  NAND U57466 ( .A(n46009), .B(n46008), .Z(n46010) );
  AND U57467 ( .A(n46011), .B(n46010), .Z(n46012) );
  OR U57468 ( .A(n46013), .B(n46012), .Z(n46014) );
  NAND U57469 ( .A(n46015), .B(n46014), .Z(n46016) );
  NANDN U57470 ( .A(n46017), .B(n46016), .Z(n46018) );
  NANDN U57471 ( .A(x[6340]), .B(y[6340]), .Z(n51099) );
  NANDN U57472 ( .A(n46018), .B(n51099), .Z(n46019) );
  AND U57473 ( .A(n46020), .B(n46019), .Z(n46021) );
  OR U57474 ( .A(n46022), .B(n46021), .Z(n46023) );
  NAND U57475 ( .A(n46024), .B(n46023), .Z(n46025) );
  NANDN U57476 ( .A(n46026), .B(n46025), .Z(n46028) );
  NANDN U57477 ( .A(n46028), .B(n46027), .Z(n46029) );
  NAND U57478 ( .A(n46030), .B(n46029), .Z(n46031) );
  AND U57479 ( .A(n46032), .B(n46031), .Z(n46036) );
  AND U57480 ( .A(n46034), .B(n46033), .Z(n46035) );
  NANDN U57481 ( .A(n46036), .B(n46035), .Z(n46037) );
  NAND U57482 ( .A(n46038), .B(n46037), .Z(n46039) );
  NAND U57483 ( .A(n46040), .B(n46039), .Z(n46041) );
  AND U57484 ( .A(n46041), .B(n51096), .Z(n46042) );
  NANDN U57485 ( .A(x[6350]), .B(y[6350]), .Z(n58980) );
  AND U57486 ( .A(n46042), .B(n58980), .Z(n46046) );
  AND U57487 ( .A(n46044), .B(n46043), .Z(n46045) );
  NANDN U57488 ( .A(n46046), .B(n46045), .Z(n46047) );
  NAND U57489 ( .A(n46048), .B(n46047), .Z(n46049) );
  NAND U57490 ( .A(n46050), .B(n46049), .Z(n46052) );
  IV U57491 ( .A(n46051), .Z(n58986) );
  AND U57492 ( .A(n46052), .B(n58986), .Z(n46053) );
  NANDN U57493 ( .A(x[6354]), .B(y[6354]), .Z(n58983) );
  AND U57494 ( .A(n46053), .B(n58983), .Z(n46057) );
  AND U57495 ( .A(n46055), .B(n46054), .Z(n46056) );
  NANDN U57496 ( .A(n46057), .B(n46056), .Z(n46058) );
  NAND U57497 ( .A(n46059), .B(n46058), .Z(n46060) );
  NAND U57498 ( .A(n46061), .B(n46060), .Z(n46062) );
  AND U57499 ( .A(n46062), .B(n51094), .Z(n46063) );
  NANDN U57500 ( .A(x[6358]), .B(y[6358]), .Z(n58990) );
  AND U57501 ( .A(n46063), .B(n58990), .Z(n46067) );
  AND U57502 ( .A(n46065), .B(n46064), .Z(n46066) );
  NANDN U57503 ( .A(n46067), .B(n46066), .Z(n46068) );
  NAND U57504 ( .A(n46069), .B(n46068), .Z(n46070) );
  AND U57505 ( .A(n46071), .B(n46070), .Z(n46072) );
  OR U57506 ( .A(n46073), .B(n46072), .Z(n46074) );
  NAND U57507 ( .A(n46075), .B(n46074), .Z(n46076) );
  NANDN U57508 ( .A(n51091), .B(n46076), .Z(n46077) );
  NANDN U57509 ( .A(x[6364]), .B(y[6364]), .Z(n58997) );
  NANDN U57510 ( .A(n46077), .B(n58997), .Z(n46078) );
  AND U57511 ( .A(n46079), .B(n46078), .Z(n46080) );
  ANDN U57512 ( .B(n51092), .A(n46080), .Z(n46081) );
  NAND U57513 ( .A(n46082), .B(n46081), .Z(n46083) );
  NANDN U57514 ( .A(n46084), .B(n46083), .Z(n46085) );
  OR U57515 ( .A(n46086), .B(n46085), .Z(n46087) );
  NAND U57516 ( .A(n46088), .B(n46087), .Z(n46089) );
  NAND U57517 ( .A(n46090), .B(n46089), .Z(n46092) );
  IV U57518 ( .A(n46091), .Z(n51089) );
  AND U57519 ( .A(n46092), .B(n51089), .Z(n46093) );
  NANDN U57520 ( .A(x[6370]), .B(y[6370]), .Z(n59003) );
  AND U57521 ( .A(n46093), .B(n59003), .Z(n46094) );
  OR U57522 ( .A(n46095), .B(n46094), .Z(n46096) );
  NAND U57523 ( .A(n46097), .B(n46096), .Z(n46098) );
  AND U57524 ( .A(n46099), .B(n46098), .Z(n46100) );
  OR U57525 ( .A(n46101), .B(n46100), .Z(n46102) );
  NAND U57526 ( .A(n46103), .B(n46102), .Z(n46104) );
  NANDN U57527 ( .A(n51085), .B(n46104), .Z(n46105) );
  NANDN U57528 ( .A(x[6376]), .B(y[6376]), .Z(n59009) );
  NANDN U57529 ( .A(n46105), .B(n59009), .Z(n46106) );
  NAND U57530 ( .A(n46107), .B(n46106), .Z(n46108) );
  AND U57531 ( .A(n46108), .B(n59012), .Z(n46109) );
  NANDN U57532 ( .A(x[6378]), .B(y[6378]), .Z(n51086) );
  AND U57533 ( .A(n46109), .B(n51086), .Z(n46113) );
  AND U57534 ( .A(n46111), .B(n46110), .Z(n46112) );
  NANDN U57535 ( .A(n46113), .B(n46112), .Z(n46114) );
  NAND U57536 ( .A(n46115), .B(n46114), .Z(n46116) );
  NAND U57537 ( .A(n46117), .B(n46116), .Z(n46118) );
  AND U57538 ( .A(n46118), .B(n59019), .Z(n46119) );
  NANDN U57539 ( .A(x[6382]), .B(y[6382]), .Z(n59017) );
  AND U57540 ( .A(n46119), .B(n59017), .Z(n46123) );
  AND U57541 ( .A(n46121), .B(n46120), .Z(n46122) );
  NANDN U57542 ( .A(n46123), .B(n46122), .Z(n46124) );
  NAND U57543 ( .A(n46125), .B(n46124), .Z(n46126) );
  NAND U57544 ( .A(n46127), .B(n46126), .Z(n46128) );
  AND U57545 ( .A(n46128), .B(n59023), .Z(n46129) );
  NANDN U57546 ( .A(x[6386]), .B(y[6386]), .Z(n51083) );
  AND U57547 ( .A(n46129), .B(n51083), .Z(n46133) );
  AND U57548 ( .A(n46131), .B(n46130), .Z(n46132) );
  NANDN U57549 ( .A(n46133), .B(n46132), .Z(n46134) );
  NAND U57550 ( .A(n46135), .B(n46134), .Z(n46136) );
  NAND U57551 ( .A(n46137), .B(n46136), .Z(n46139) );
  IV U57552 ( .A(n46138), .Z(n59029) );
  AND U57553 ( .A(n46139), .B(n59029), .Z(n46140) );
  NANDN U57554 ( .A(x[6390]), .B(y[6390]), .Z(n59027) );
  AND U57555 ( .A(n46140), .B(n59027), .Z(n46144) );
  AND U57556 ( .A(n46142), .B(n46141), .Z(n46143) );
  NANDN U57557 ( .A(n46144), .B(n46143), .Z(n46145) );
  NAND U57558 ( .A(n46146), .B(n46145), .Z(n46147) );
  NAND U57559 ( .A(n46148), .B(n46147), .Z(n46149) );
  AND U57560 ( .A(n46149), .B(n51078), .Z(n46150) );
  NANDN U57561 ( .A(x[6394]), .B(y[6394]), .Z(n51081) );
  AND U57562 ( .A(n46150), .B(n51081), .Z(n46154) );
  AND U57563 ( .A(n46152), .B(n46151), .Z(n46153) );
  NANDN U57564 ( .A(n46154), .B(n46153), .Z(n46155) );
  NAND U57565 ( .A(n46156), .B(n46155), .Z(n46157) );
  AND U57566 ( .A(n46158), .B(n46157), .Z(n46161) );
  NANDN U57567 ( .A(x[6398]), .B(y[6398]), .Z(n59036) );
  IV U57568 ( .A(n46159), .Z(n59038) );
  AND U57569 ( .A(n59036), .B(n59038), .Z(n46160) );
  NANDN U57570 ( .A(n46161), .B(n46160), .Z(n46162) );
  NANDN U57571 ( .A(n46163), .B(n46162), .Z(n46164) );
  AND U57572 ( .A(n51075), .B(n46164), .Z(n46165) );
  NANDN U57573 ( .A(x[6400]), .B(y[6400]), .Z(n59039) );
  NAND U57574 ( .A(n46165), .B(n59039), .Z(n46166) );
  NAND U57575 ( .A(n46167), .B(n46166), .Z(n46168) );
  AND U57576 ( .A(n46168), .B(n59044), .Z(n46169) );
  NANDN U57577 ( .A(x[6402]), .B(y[6402]), .Z(n51076) );
  AND U57578 ( .A(n46169), .B(n51076), .Z(n46173) );
  AND U57579 ( .A(n46171), .B(n46170), .Z(n46172) );
  NANDN U57580 ( .A(n46173), .B(n46172), .Z(n46174) );
  NAND U57581 ( .A(n46175), .B(n46174), .Z(n46176) );
  NAND U57582 ( .A(n46177), .B(n46176), .Z(n46178) );
  AND U57583 ( .A(n46178), .B(n59050), .Z(n46179) );
  NANDN U57584 ( .A(x[6406]), .B(y[6406]), .Z(n51074) );
  AND U57585 ( .A(n46179), .B(n51074), .Z(n46183) );
  AND U57586 ( .A(n46181), .B(n46180), .Z(n46182) );
  NANDN U57587 ( .A(n46183), .B(n46182), .Z(n46184) );
  NAND U57588 ( .A(n46185), .B(n46184), .Z(n46186) );
  NAND U57589 ( .A(n46187), .B(n46186), .Z(n46188) );
  AND U57590 ( .A(n46188), .B(n59055), .Z(n46189) );
  NANDN U57591 ( .A(x[6410]), .B(y[6410]), .Z(n51073) );
  AND U57592 ( .A(n46189), .B(n51073), .Z(n46190) );
  OR U57593 ( .A(n46191), .B(n46190), .Z(n46192) );
  NAND U57594 ( .A(n46193), .B(n46192), .Z(n46194) );
  NAND U57595 ( .A(n46195), .B(n46194), .Z(n46197) );
  IV U57596 ( .A(n46196), .Z(n59062) );
  AND U57597 ( .A(n46197), .B(n59062), .Z(n46198) );
  NANDN U57598 ( .A(x[6414]), .B(y[6414]), .Z(n59058) );
  AND U57599 ( .A(n46198), .B(n59058), .Z(n46202) );
  AND U57600 ( .A(n46200), .B(n46199), .Z(n46201) );
  NANDN U57601 ( .A(n46202), .B(n46201), .Z(n46203) );
  NAND U57602 ( .A(n46204), .B(n46203), .Z(n46205) );
  AND U57603 ( .A(n46206), .B(n46205), .Z(n46207) );
  ANDN U57604 ( .B(n51071), .A(n46207), .Z(n46208) );
  NAND U57605 ( .A(n59066), .B(n46208), .Z(n46209) );
  NANDN U57606 ( .A(n46210), .B(n46209), .Z(n46211) );
  OR U57607 ( .A(n46212), .B(n46211), .Z(n46213) );
  NAND U57608 ( .A(n46214), .B(n46213), .Z(n46215) );
  NAND U57609 ( .A(n46216), .B(n46215), .Z(n46217) );
  AND U57610 ( .A(n46217), .B(n59071), .Z(n46218) );
  NANDN U57611 ( .A(x[6422]), .B(y[6422]), .Z(n59069) );
  AND U57612 ( .A(n46218), .B(n59069), .Z(n46219) );
  OR U57613 ( .A(n46220), .B(n46219), .Z(n46221) );
  NAND U57614 ( .A(n46222), .B(n46221), .Z(n46223) );
  AND U57615 ( .A(n46224), .B(n46223), .Z(n46225) );
  OR U57616 ( .A(n46226), .B(n46225), .Z(n46227) );
  NAND U57617 ( .A(n46228), .B(n46227), .Z(n46229) );
  NANDN U57618 ( .A(n46230), .B(n46229), .Z(n46231) );
  NAND U57619 ( .A(n46232), .B(n46231), .Z(n46234) );
  IV U57620 ( .A(n46233), .Z(n51065) );
  AND U57621 ( .A(n46234), .B(n51065), .Z(n46236) );
  NANDN U57622 ( .A(x[6430]), .B(y[6430]), .Z(n46235) );
  AND U57623 ( .A(n46236), .B(n46235), .Z(n46237) );
  OR U57624 ( .A(n46238), .B(n46237), .Z(n46239) );
  NAND U57625 ( .A(n46240), .B(n46239), .Z(n46241) );
  NAND U57626 ( .A(n46242), .B(n46241), .Z(n46243) );
  NAND U57627 ( .A(n46244), .B(n46243), .Z(n46245) );
  NAND U57628 ( .A(n46246), .B(n46245), .Z(n46252) );
  NAND U57629 ( .A(n46248), .B(n46247), .Z(n46249) );
  NAND U57630 ( .A(n46250), .B(n46249), .Z(n46251) );
  AND U57631 ( .A(n46252), .B(n46251), .Z(n46253) );
  OR U57632 ( .A(n46254), .B(n46253), .Z(n46255) );
  NAND U57633 ( .A(n46256), .B(n46255), .Z(n46257) );
  NANDN U57634 ( .A(n46258), .B(n46257), .Z(n46259) );
  AND U57635 ( .A(n46259), .B(n59090), .Z(n46260) );
  NANDN U57636 ( .A(x[6440]), .B(y[6440]), .Z(n59088) );
  NAND U57637 ( .A(n46260), .B(n59088), .Z(n46261) );
  AND U57638 ( .A(n46262), .B(n46261), .Z(n46263) );
  ANDN U57639 ( .B(n46264), .A(n46263), .Z(n46265) );
  NAND U57640 ( .A(n59091), .B(n46265), .Z(n46266) );
  NANDN U57641 ( .A(n46267), .B(n46266), .Z(n46268) );
  AND U57642 ( .A(n46269), .B(n46268), .Z(n46270) );
  OR U57643 ( .A(n46271), .B(n46270), .Z(n46272) );
  NAND U57644 ( .A(n46273), .B(n46272), .Z(n46274) );
  NANDN U57645 ( .A(n46275), .B(n46274), .Z(n46277) );
  IV U57646 ( .A(n46276), .Z(n51060) );
  AND U57647 ( .A(n46277), .B(n51060), .Z(n46278) );
  NANDN U57648 ( .A(x[6448]), .B(y[6448]), .Z(n59098) );
  NAND U57649 ( .A(n46278), .B(n59098), .Z(n46279) );
  AND U57650 ( .A(n46280), .B(n46279), .Z(n46281) );
  ANDN U57651 ( .B(n59103), .A(n46281), .Z(n46282) );
  NAND U57652 ( .A(n51061), .B(n46282), .Z(n46283) );
  NANDN U57653 ( .A(n46284), .B(n46283), .Z(n46286) );
  NANDN U57654 ( .A(n46286), .B(n46285), .Z(n46288) );
  AND U57655 ( .A(n46288), .B(n46287), .Z(n46289) );
  NANDN U57656 ( .A(x[6452]), .B(y[6452]), .Z(n59105) );
  AND U57657 ( .A(n46289), .B(n59105), .Z(n46290) );
  OR U57658 ( .A(n46291), .B(n46290), .Z(n46292) );
  NAND U57659 ( .A(n46293), .B(n46292), .Z(n46294) );
  NANDN U57660 ( .A(n46295), .B(n46294), .Z(n46296) );
  NAND U57661 ( .A(n46297), .B(n46296), .Z(n46298) );
  AND U57662 ( .A(n46299), .B(n46298), .Z(n46300) );
  ANDN U57663 ( .B(n59114), .A(n46300), .Z(n46301) );
  NAND U57664 ( .A(n59111), .B(n46301), .Z(n46302) );
  NANDN U57665 ( .A(n46303), .B(n46302), .Z(n46304) );
  AND U57666 ( .A(n46304), .B(n59117), .Z(n46305) );
  NANDN U57667 ( .A(x[6460]), .B(y[6460]), .Z(n59115) );
  NAND U57668 ( .A(n46305), .B(n59115), .Z(n46306) );
  AND U57669 ( .A(n46307), .B(n46306), .Z(n46308) );
  ANDN U57670 ( .B(n51058), .A(n46308), .Z(n46309) );
  NAND U57671 ( .A(n59118), .B(n46309), .Z(n46310) );
  NANDN U57672 ( .A(n46311), .B(n46310), .Z(n46312) );
  AND U57673 ( .A(n46312), .B(n59123), .Z(n46313) );
  NANDN U57674 ( .A(x[6464]), .B(y[6464]), .Z(n51059) );
  NAND U57675 ( .A(n46313), .B(n51059), .Z(n46314) );
  AND U57676 ( .A(n46315), .B(n46314), .Z(n46316) );
  ANDN U57677 ( .B(n59125), .A(n46316), .Z(n46317) );
  NAND U57678 ( .A(n59122), .B(n46317), .Z(n46318) );
  NANDN U57679 ( .A(n46319), .B(n46318), .Z(n46320) );
  AND U57680 ( .A(n46320), .B(n59128), .Z(n46321) );
  NANDN U57681 ( .A(x[6468]), .B(y[6468]), .Z(n59126) );
  NAND U57682 ( .A(n46321), .B(n59126), .Z(n46322) );
  NAND U57683 ( .A(n46323), .B(n46322), .Z(n46325) );
  IV U57684 ( .A(n46324), .Z(n51056) );
  AND U57685 ( .A(n46325), .B(n51056), .Z(n46326) );
  NANDN U57686 ( .A(x[6470]), .B(y[6470]), .Z(n59129) );
  AND U57687 ( .A(n46326), .B(n59129), .Z(n46327) );
  NOR U57688 ( .A(n46328), .B(n46327), .Z(n46330) );
  XNOR U57689 ( .A(x[6472]), .B(y[6472]), .Z(n46329) );
  NAND U57690 ( .A(n46330), .B(n46329), .Z(n46331) );
  AND U57691 ( .A(n46331), .B(n59133), .Z(n46332) );
  NANDN U57692 ( .A(x[6472]), .B(y[6472]), .Z(n51057) );
  NAND U57693 ( .A(n46332), .B(n51057), .Z(n46333) );
  AND U57694 ( .A(n46334), .B(n46333), .Z(n46335) );
  ANDN U57695 ( .B(n59136), .A(n46335), .Z(n46336) );
  NAND U57696 ( .A(n59132), .B(n46336), .Z(n46337) );
  NANDN U57697 ( .A(n46338), .B(n46337), .Z(n46339) );
  AND U57698 ( .A(n46339), .B(n59142), .Z(n46340) );
  NANDN U57699 ( .A(x[6476]), .B(y[6476]), .Z(n59137) );
  AND U57700 ( .A(n46340), .B(n59137), .Z(n46341) );
  OR U57701 ( .A(n46342), .B(n46341), .Z(n46343) );
  NAND U57702 ( .A(n46344), .B(n46343), .Z(n46345) );
  NANDN U57703 ( .A(n46346), .B(n46345), .Z(n46348) );
  OR U57704 ( .A(n46348), .B(n46347), .Z(n46349) );
  AND U57705 ( .A(n59154), .B(n46349), .Z(n46350) );
  NANDN U57706 ( .A(x[6480]), .B(y[6480]), .Z(n51055) );
  NAND U57707 ( .A(n46350), .B(n51055), .Z(n46351) );
  AND U57708 ( .A(n46352), .B(n46351), .Z(n46354) );
  NANDN U57709 ( .A(x[6482]), .B(y[6482]), .Z(n59151) );
  AND U57710 ( .A(n59151), .B(n59158), .Z(n46353) );
  NANDN U57711 ( .A(n46354), .B(n46353), .Z(n46355) );
  NANDN U57712 ( .A(n46356), .B(n46355), .Z(n46357) );
  AND U57713 ( .A(n59164), .B(n46357), .Z(n46358) );
  NANDN U57714 ( .A(x[6484]), .B(y[6484]), .Z(n59159) );
  NAND U57715 ( .A(n46358), .B(n59159), .Z(n46359) );
  AND U57716 ( .A(n46360), .B(n46359), .Z(n46362) );
  NANDN U57717 ( .A(x[6486]), .B(y[6486]), .Z(n59165) );
  AND U57718 ( .A(n59165), .B(n51052), .Z(n46361) );
  NANDN U57719 ( .A(n46362), .B(n46361), .Z(n46363) );
  NANDN U57720 ( .A(n46364), .B(n46363), .Z(n46365) );
  AND U57721 ( .A(n46365), .B(n59175), .Z(n46366) );
  NANDN U57722 ( .A(x[6488]), .B(y[6488]), .Z(n51053) );
  NAND U57723 ( .A(n46366), .B(n51053), .Z(n46367) );
  AND U57724 ( .A(n46368), .B(n46367), .Z(n46370) );
  NANDN U57725 ( .A(x[6490]), .B(y[6490]), .Z(n59173) );
  AND U57726 ( .A(n59177), .B(n59173), .Z(n46369) );
  NANDN U57727 ( .A(n46370), .B(n46369), .Z(n46371) );
  NANDN U57728 ( .A(n46372), .B(n46371), .Z(n46373) );
  AND U57729 ( .A(n59180), .B(n46373), .Z(n46374) );
  NANDN U57730 ( .A(x[6492]), .B(y[6492]), .Z(n59178) );
  NAND U57731 ( .A(n46374), .B(n59178), .Z(n46375) );
  AND U57732 ( .A(n46376), .B(n46375), .Z(n46378) );
  NANDN U57733 ( .A(x[6494]), .B(y[6494]), .Z(n59181) );
  AND U57734 ( .A(n59181), .B(n51050), .Z(n46377) );
  NANDN U57735 ( .A(n46378), .B(n46377), .Z(n46379) );
  NANDN U57736 ( .A(n46380), .B(n46379), .Z(n46381) );
  AND U57737 ( .A(n46381), .B(n59185), .Z(n46382) );
  NANDN U57738 ( .A(x[6496]), .B(y[6496]), .Z(n51051) );
  NAND U57739 ( .A(n46382), .B(n51051), .Z(n46383) );
  AND U57740 ( .A(n46384), .B(n46383), .Z(n46386) );
  NANDN U57741 ( .A(x[6498]), .B(y[6498]), .Z(n59184) );
  AND U57742 ( .A(n59187), .B(n59184), .Z(n46385) );
  NANDN U57743 ( .A(n46386), .B(n46385), .Z(n46387) );
  NANDN U57744 ( .A(n46388), .B(n46387), .Z(n46389) );
  AND U57745 ( .A(n59191), .B(n46389), .Z(n46390) );
  NANDN U57746 ( .A(x[6500]), .B(y[6500]), .Z(n59188) );
  NAND U57747 ( .A(n46390), .B(n59188), .Z(n46391) );
  AND U57748 ( .A(n46392), .B(n46391), .Z(n46394) );
  NANDN U57749 ( .A(x[6502]), .B(y[6502]), .Z(n59192) );
  AND U57750 ( .A(n59192), .B(n51048), .Z(n46393) );
  NANDN U57751 ( .A(n46394), .B(n46393), .Z(n46395) );
  NAND U57752 ( .A(n46396), .B(n46395), .Z(n46397) );
  OR U57753 ( .A(n46398), .B(n46397), .Z(n46399) );
  AND U57754 ( .A(n46399), .B(n59196), .Z(n46400) );
  NANDN U57755 ( .A(x[6504]), .B(y[6504]), .Z(n51049) );
  NAND U57756 ( .A(n46400), .B(n51049), .Z(n46401) );
  AND U57757 ( .A(n46402), .B(n46401), .Z(n46404) );
  NANDN U57758 ( .A(x[6506]), .B(y[6506]), .Z(n59195) );
  AND U57759 ( .A(n59198), .B(n59195), .Z(n46403) );
  NANDN U57760 ( .A(n46404), .B(n46403), .Z(n46405) );
  NANDN U57761 ( .A(n46406), .B(n46405), .Z(n46408) );
  IV U57762 ( .A(n46407), .Z(n59201) );
  AND U57763 ( .A(n46408), .B(n59201), .Z(n46409) );
  NANDN U57764 ( .A(x[6508]), .B(y[6508]), .Z(n59199) );
  NAND U57765 ( .A(n46409), .B(n59199), .Z(n46410) );
  AND U57766 ( .A(n46411), .B(n46410), .Z(n46413) );
  NANDN U57767 ( .A(x[6510]), .B(y[6510]), .Z(n59202) );
  AND U57768 ( .A(n59202), .B(n51046), .Z(n46412) );
  NANDN U57769 ( .A(n46413), .B(n46412), .Z(n46414) );
  NANDN U57770 ( .A(n46415), .B(n46414), .Z(n46416) );
  AND U57771 ( .A(n46416), .B(n59209), .Z(n46417) );
  NANDN U57772 ( .A(x[6512]), .B(y[6512]), .Z(n51047) );
  NAND U57773 ( .A(n46417), .B(n51047), .Z(n46418) );
  NAND U57774 ( .A(n46419), .B(n46418), .Z(n46420) );
  AND U57775 ( .A(n46420), .B(n59210), .Z(n46421) );
  NAND U57776 ( .A(n59207), .B(n46421), .Z(n46422) );
  NANDN U57777 ( .A(n46423), .B(n46422), .Z(n46424) );
  AND U57778 ( .A(n59213), .B(n46424), .Z(n46425) );
  NANDN U57779 ( .A(x[6516]), .B(y[6516]), .Z(n59211) );
  NAND U57780 ( .A(n46425), .B(n59211), .Z(n46426) );
  AND U57781 ( .A(n46427), .B(n46426), .Z(n46429) );
  NANDN U57782 ( .A(x[6518]), .B(y[6518]), .Z(n59214) );
  AND U57783 ( .A(n59214), .B(n51043), .Z(n46428) );
  NANDN U57784 ( .A(n46429), .B(n46428), .Z(n46430) );
  NANDN U57785 ( .A(n46431), .B(n46430), .Z(n46432) );
  AND U57786 ( .A(n46432), .B(n59218), .Z(n46433) );
  NANDN U57787 ( .A(x[6520]), .B(y[6520]), .Z(n51044) );
  NAND U57788 ( .A(n46433), .B(n51044), .Z(n46434) );
  AND U57789 ( .A(n46435), .B(n46434), .Z(n46436) );
  ANDN U57790 ( .B(n59221), .A(n46436), .Z(n46437) );
  NAND U57791 ( .A(n59217), .B(n46437), .Z(n46438) );
  NANDN U57792 ( .A(n46439), .B(n46438), .Z(n46440) );
  AND U57793 ( .A(n46440), .B(n59224), .Z(n46441) );
  NANDN U57794 ( .A(x[6524]), .B(y[6524]), .Z(n59222) );
  NAND U57795 ( .A(n46441), .B(n59222), .Z(n46442) );
  AND U57796 ( .A(n46443), .B(n46442), .Z(n46445) );
  NANDN U57797 ( .A(x[6526]), .B(y[6526]), .Z(n59225) );
  AND U57798 ( .A(n59225), .B(n51041), .Z(n46444) );
  NANDN U57799 ( .A(n46445), .B(n46444), .Z(n46446) );
  NANDN U57800 ( .A(n46447), .B(n46446), .Z(n46448) );
  AND U57801 ( .A(n46449), .B(n46448), .Z(n46450) );
  NANDN U57802 ( .A(x[6528]), .B(y[6528]), .Z(n51042) );
  NAND U57803 ( .A(n46450), .B(n51042), .Z(n46451) );
  AND U57804 ( .A(n46452), .B(n46451), .Z(n46453) );
  OR U57805 ( .A(n46454), .B(n46453), .Z(n46455) );
  NAND U57806 ( .A(n46456), .B(n46455), .Z(n46457) );
  AND U57807 ( .A(n46457), .B(n51039), .Z(n46459) );
  NANDN U57808 ( .A(x[6532]), .B(y[6532]), .Z(n46458) );
  NAND U57809 ( .A(n46459), .B(n46458), .Z(n46460) );
  AND U57810 ( .A(n46461), .B(n46460), .Z(n46462) );
  ANDN U57811 ( .B(n59234), .A(n46462), .Z(n46463) );
  NAND U57812 ( .A(n51040), .B(n46463), .Z(n46464) );
  NANDN U57813 ( .A(n46465), .B(n46464), .Z(n46466) );
  AND U57814 ( .A(n46466), .B(n59236), .Z(n46467) );
  NANDN U57815 ( .A(x[6536]), .B(y[6536]), .Z(n59233) );
  NAND U57816 ( .A(n46467), .B(n59233), .Z(n46468) );
  AND U57817 ( .A(n46469), .B(n46468), .Z(n46470) );
  ANDN U57818 ( .B(n59239), .A(n46470), .Z(n46471) );
  NAND U57819 ( .A(n59237), .B(n46471), .Z(n46472) );
  NANDN U57820 ( .A(n46473), .B(n46472), .Z(n46474) );
  AND U57821 ( .A(n46474), .B(n51036), .Z(n46475) );
  NANDN U57822 ( .A(x[6540]), .B(y[6540]), .Z(n59240) );
  NAND U57823 ( .A(n46475), .B(n59240), .Z(n46476) );
  AND U57824 ( .A(n46477), .B(n46476), .Z(n46478) );
  ANDN U57825 ( .B(n46479), .A(n46478), .Z(n46480) );
  NAND U57826 ( .A(n51037), .B(n46480), .Z(n46481) );
  NANDN U57827 ( .A(n46482), .B(n46481), .Z(n46483) );
  AND U57828 ( .A(n46483), .B(n59245), .Z(n46484) );
  NANDN U57829 ( .A(x[6544]), .B(y[6544]), .Z(n59244) );
  NAND U57830 ( .A(n46484), .B(n59244), .Z(n46485) );
  AND U57831 ( .A(n46486), .B(n46485), .Z(n46487) );
  ANDN U57832 ( .B(n46488), .A(n46487), .Z(n46489) );
  NAND U57833 ( .A(n51034), .B(n46489), .Z(n46490) );
  NANDN U57834 ( .A(n46491), .B(n46490), .Z(n46492) );
  AND U57835 ( .A(n46492), .B(n59251), .Z(n46494) );
  NANDN U57836 ( .A(x[6548]), .B(y[6548]), .Z(n46493) );
  AND U57837 ( .A(n46494), .B(n46493), .Z(n46495) );
  OR U57838 ( .A(n46496), .B(n46495), .Z(n46497) );
  NAND U57839 ( .A(n46498), .B(n46497), .Z(n46499) );
  NANDN U57840 ( .A(n46500), .B(n46499), .Z(n46501) );
  AND U57841 ( .A(n46501), .B(n59256), .Z(n46502) );
  NANDN U57842 ( .A(x[6552]), .B(y[6552]), .Z(n59254) );
  AND U57843 ( .A(n46502), .B(n59254), .Z(n46503) );
  OR U57844 ( .A(n46504), .B(n46503), .Z(n46505) );
  NAND U57845 ( .A(n46506), .B(n46505), .Z(n46507) );
  NANDN U57846 ( .A(n46508), .B(n46507), .Z(n46509) );
  OR U57847 ( .A(n46510), .B(n46509), .Z(n46511) );
  AND U57848 ( .A(n46511), .B(n59261), .Z(n46512) );
  NANDN U57849 ( .A(x[6556]), .B(y[6556]), .Z(n51033) );
  NAND U57850 ( .A(n46512), .B(n51033), .Z(n46513) );
  AND U57851 ( .A(n46514), .B(n46513), .Z(n46516) );
  NANDN U57852 ( .A(x[6558]), .B(y[6558]), .Z(n59260) );
  AND U57853 ( .A(n59264), .B(n59260), .Z(n46515) );
  NANDN U57854 ( .A(n46516), .B(n46515), .Z(n46517) );
  NANDN U57855 ( .A(n46518), .B(n46517), .Z(n46519) );
  AND U57856 ( .A(n46520), .B(n46519), .Z(n46521) );
  NANDN U57857 ( .A(x[6560]), .B(y[6560]), .Z(n59265) );
  NAND U57858 ( .A(n46521), .B(n59265), .Z(n46522) );
  AND U57859 ( .A(n46523), .B(n46522), .Z(n46527) );
  NAND U57860 ( .A(n46525), .B(n46524), .Z(n46526) );
  OR U57861 ( .A(n46527), .B(n46526), .Z(n46528) );
  NAND U57862 ( .A(n46529), .B(n46528), .Z(n46530) );
  AND U57863 ( .A(n46531), .B(n46530), .Z(n46532) );
  OR U57864 ( .A(n46533), .B(n46532), .Z(n46534) );
  NAND U57865 ( .A(n46535), .B(n46534), .Z(n46536) );
  NANDN U57866 ( .A(n46537), .B(n46536), .Z(n46538) );
  AND U57867 ( .A(n46538), .B(n59275), .Z(n46539) );
  NANDN U57868 ( .A(x[6568]), .B(y[6568]), .Z(n51030) );
  NAND U57869 ( .A(n46539), .B(n51030), .Z(n46540) );
  AND U57870 ( .A(n46541), .B(n46540), .Z(n46542) );
  ANDN U57871 ( .B(n59277), .A(n46542), .Z(n46543) );
  NAND U57872 ( .A(n59274), .B(n46543), .Z(n46544) );
  NANDN U57873 ( .A(n46545), .B(n46544), .Z(n46546) );
  AND U57874 ( .A(n46546), .B(n59281), .Z(n46547) );
  NANDN U57875 ( .A(x[6572]), .B(y[6572]), .Z(n59278) );
  AND U57876 ( .A(n46547), .B(n59278), .Z(n46551) );
  AND U57877 ( .A(n46549), .B(n46548), .Z(n46550) );
  NANDN U57878 ( .A(n46551), .B(n46550), .Z(n46553) );
  IV U57879 ( .A(n46552), .Z(n51027) );
  AND U57880 ( .A(n46553), .B(n51027), .Z(n46554) );
  NANDN U57881 ( .A(x[6574]), .B(y[6574]), .Z(n59282) );
  AND U57882 ( .A(n46554), .B(n59282), .Z(n46555) );
  NOR U57883 ( .A(n46556), .B(n46555), .Z(n46558) );
  XNOR U57884 ( .A(x[6576]), .B(y[6576]), .Z(n46557) );
  NAND U57885 ( .A(n46558), .B(n46557), .Z(n46559) );
  AND U57886 ( .A(n46559), .B(n59286), .Z(n46560) );
  NANDN U57887 ( .A(x[6576]), .B(y[6576]), .Z(n51028) );
  NAND U57888 ( .A(n46560), .B(n51028), .Z(n46561) );
  NAND U57889 ( .A(n46562), .B(n46561), .Z(n46564) );
  NANDN U57890 ( .A(x[6578]), .B(y[6578]), .Z(n59285) );
  AND U57891 ( .A(n59288), .B(n59285), .Z(n46563) );
  NAND U57892 ( .A(n46564), .B(n46563), .Z(n46565) );
  NANDN U57893 ( .A(n46566), .B(n46565), .Z(n46567) );
  AND U57894 ( .A(n46567), .B(n59291), .Z(n46568) );
  NANDN U57895 ( .A(x[6580]), .B(y[6580]), .Z(n59289) );
  AND U57896 ( .A(n46568), .B(n59289), .Z(n46569) );
  OR U57897 ( .A(n46570), .B(n46569), .Z(n46571) );
  NAND U57898 ( .A(n46572), .B(n46571), .Z(n46573) );
  NANDN U57899 ( .A(n46574), .B(n46573), .Z(n46576) );
  OR U57900 ( .A(n46576), .B(n46575), .Z(n46577) );
  AND U57901 ( .A(n59298), .B(n46577), .Z(n46578) );
  NANDN U57902 ( .A(x[6584]), .B(y[6584]), .Z(n51026) );
  NAND U57903 ( .A(n46578), .B(n51026), .Z(n46579) );
  AND U57904 ( .A(n46580), .B(n46579), .Z(n46582) );
  NANDN U57905 ( .A(x[6586]), .B(y[6586]), .Z(n59297) );
  AND U57906 ( .A(n59297), .B(n59299), .Z(n46581) );
  NANDN U57907 ( .A(n46582), .B(n46581), .Z(n46583) );
  NANDN U57908 ( .A(n46584), .B(n46583), .Z(n46585) );
  AND U57909 ( .A(n59302), .B(n46585), .Z(n46586) );
  NANDN U57910 ( .A(x[6588]), .B(y[6588]), .Z(n59300) );
  NAND U57911 ( .A(n46586), .B(n59300), .Z(n46587) );
  AND U57912 ( .A(n46588), .B(n46587), .Z(n46590) );
  NANDN U57913 ( .A(x[6590]), .B(y[6590]), .Z(n59303) );
  AND U57914 ( .A(n59303), .B(n51022), .Z(n46589) );
  NANDN U57915 ( .A(n46590), .B(n46589), .Z(n46591) );
  NANDN U57916 ( .A(n46592), .B(n46591), .Z(n46593) );
  AND U57917 ( .A(n46593), .B(n59307), .Z(n46594) );
  NANDN U57918 ( .A(x[6592]), .B(y[6592]), .Z(n51023) );
  NAND U57919 ( .A(n46594), .B(n51023), .Z(n46595) );
  AND U57920 ( .A(n46596), .B(n46595), .Z(n46598) );
  NANDN U57921 ( .A(x[6594]), .B(y[6594]), .Z(n59306) );
  AND U57922 ( .A(n59310), .B(n59306), .Z(n46597) );
  NANDN U57923 ( .A(n46598), .B(n46597), .Z(n46599) );
  NANDN U57924 ( .A(n46600), .B(n46599), .Z(n46601) );
  AND U57925 ( .A(n59313), .B(n46601), .Z(n46602) );
  NANDN U57926 ( .A(x[6596]), .B(y[6596]), .Z(n59311) );
  NAND U57927 ( .A(n46602), .B(n59311), .Z(n46603) );
  AND U57928 ( .A(n46604), .B(n46603), .Z(n46606) );
  NANDN U57929 ( .A(x[6598]), .B(y[6598]), .Z(n59314) );
  AND U57930 ( .A(n59314), .B(n51020), .Z(n46605) );
  NANDN U57931 ( .A(n46606), .B(n46605), .Z(n46607) );
  NANDN U57932 ( .A(n46608), .B(n46607), .Z(n46609) );
  AND U57933 ( .A(n46609), .B(n59318), .Z(n46610) );
  NANDN U57934 ( .A(x[6600]), .B(y[6600]), .Z(n51021) );
  NAND U57935 ( .A(n46610), .B(n51021), .Z(n46611) );
  AND U57936 ( .A(n46612), .B(n46611), .Z(n46614) );
  NANDN U57937 ( .A(x[6602]), .B(y[6602]), .Z(n59317) );
  AND U57938 ( .A(n59320), .B(n59317), .Z(n46613) );
  NANDN U57939 ( .A(n46614), .B(n46613), .Z(n46615) );
  NANDN U57940 ( .A(n46616), .B(n46615), .Z(n46617) );
  AND U57941 ( .A(n59323), .B(n46617), .Z(n46618) );
  NANDN U57942 ( .A(x[6604]), .B(y[6604]), .Z(n59321) );
  NAND U57943 ( .A(n46618), .B(n59321), .Z(n46619) );
  AND U57944 ( .A(n46620), .B(n46619), .Z(n46621) );
  ANDN U57945 ( .B(n59326), .A(n46621), .Z(n46622) );
  NAND U57946 ( .A(n59324), .B(n46622), .Z(n46623) );
  NANDN U57947 ( .A(n46624), .B(n46623), .Z(n46626) );
  OR U57948 ( .A(n46626), .B(n46625), .Z(n46627) );
  NAND U57949 ( .A(n46628), .B(n46627), .Z(n46629) );
  NAND U57950 ( .A(n46630), .B(n46629), .Z(n46631) );
  AND U57951 ( .A(n46631), .B(n59331), .Z(n46632) );
  NANDN U57952 ( .A(x[6610]), .B(y[6610]), .Z(n51019) );
  AND U57953 ( .A(n46632), .B(n51019), .Z(n46636) );
  AND U57954 ( .A(n46634), .B(n46633), .Z(n46635) );
  NANDN U57955 ( .A(n46636), .B(n46635), .Z(n46637) );
  NAND U57956 ( .A(n46638), .B(n46637), .Z(n46639) );
  NAND U57957 ( .A(n46640), .B(n46639), .Z(n46641) );
  AND U57958 ( .A(n46641), .B(n59334), .Z(n46642) );
  NANDN U57959 ( .A(x[6614]), .B(y[6614]), .Z(n51017) );
  AND U57960 ( .A(n46642), .B(n51017), .Z(n46646) );
  AND U57961 ( .A(n46644), .B(n46643), .Z(n46645) );
  NANDN U57962 ( .A(n46646), .B(n46645), .Z(n46647) );
  NAND U57963 ( .A(n46648), .B(n46647), .Z(n46649) );
  AND U57964 ( .A(n46650), .B(n46649), .Z(n46651) );
  OR U57965 ( .A(n46652), .B(n46651), .Z(n46653) );
  NAND U57966 ( .A(n46654), .B(n46653), .Z(n46655) );
  NANDN U57967 ( .A(n46656), .B(n46655), .Z(n46657) );
  AND U57968 ( .A(n46658), .B(n46657), .Z(n46659) );
  OR U57969 ( .A(n46660), .B(n46659), .Z(n46661) );
  NAND U57970 ( .A(n46662), .B(n46661), .Z(n46663) );
  NANDN U57971 ( .A(n46664), .B(n46663), .Z(n46665) );
  NAND U57972 ( .A(n46666), .B(n46665), .Z(n46668) );
  AND U57973 ( .A(n46668), .B(n46667), .Z(n46669) );
  NAND U57974 ( .A(n59348), .B(n46669), .Z(n46670) );
  NAND U57975 ( .A(n46671), .B(n46670), .Z(n46672) );
  NANDN U57976 ( .A(n46673), .B(n46672), .Z(n46674) );
  AND U57977 ( .A(n46675), .B(n46674), .Z(n46676) );
  OR U57978 ( .A(n46677), .B(n46676), .Z(n46678) );
  NAND U57979 ( .A(n46679), .B(n46678), .Z(n46680) );
  NANDN U57980 ( .A(n46681), .B(n46680), .Z(n46682) );
  NAND U57981 ( .A(n46683), .B(n46682), .Z(n46684) );
  AND U57982 ( .A(n46684), .B(n59358), .Z(n46686) );
  NANDN U57983 ( .A(x[6634]), .B(y[6634]), .Z(n46685) );
  NAND U57984 ( .A(n46686), .B(n46685), .Z(n46687) );
  NAND U57985 ( .A(n46688), .B(n46687), .Z(n46689) );
  NANDN U57986 ( .A(x[6636]), .B(y[6636]), .Z(n59359) );
  AND U57987 ( .A(n46689), .B(n59359), .Z(n46690) );
  NANDN U57988 ( .A(n59361), .B(n46690), .Z(n46691) );
  NAND U57989 ( .A(n46692), .B(n46691), .Z(n46693) );
  AND U57990 ( .A(n46693), .B(n51010), .Z(n46694) );
  NANDN U57991 ( .A(x[6638]), .B(y[6638]), .Z(n59362) );
  AND U57992 ( .A(n46694), .B(n59362), .Z(n46698) );
  AND U57993 ( .A(n46696), .B(n46695), .Z(n46697) );
  NANDN U57994 ( .A(n46698), .B(n46697), .Z(n46699) );
  NAND U57995 ( .A(n46700), .B(n46699), .Z(n46701) );
  NAND U57996 ( .A(n46702), .B(n46701), .Z(n46703) );
  AND U57997 ( .A(n46703), .B(n51009), .Z(n46704) );
  NANDN U57998 ( .A(x[6642]), .B(y[6642]), .Z(n59366) );
  AND U57999 ( .A(n46704), .B(n59366), .Z(n46708) );
  AND U58000 ( .A(n46706), .B(n46705), .Z(n46707) );
  NANDN U58001 ( .A(n46708), .B(n46707), .Z(n46709) );
  NAND U58002 ( .A(n46710), .B(n46709), .Z(n46711) );
  NAND U58003 ( .A(n46712), .B(n46711), .Z(n46713) );
  AND U58004 ( .A(n46713), .B(n51007), .Z(n46714) );
  NANDN U58005 ( .A(x[6646]), .B(y[6646]), .Z(n59371) );
  AND U58006 ( .A(n46714), .B(n59371), .Z(n46718) );
  AND U58007 ( .A(n46716), .B(n46715), .Z(n46717) );
  NANDN U58008 ( .A(n46718), .B(n46717), .Z(n46719) );
  NAND U58009 ( .A(n46720), .B(n46719), .Z(n46721) );
  AND U58010 ( .A(n46722), .B(n46721), .Z(n46723) );
  OR U58011 ( .A(n46724), .B(n46723), .Z(n46725) );
  NAND U58012 ( .A(n46726), .B(n46725), .Z(n46727) );
  NANDN U58013 ( .A(n46728), .B(n46727), .Z(n46729) );
  NAND U58014 ( .A(n46730), .B(n46729), .Z(n46731) );
  AND U58015 ( .A(n46732), .B(n46731), .Z(n46736) );
  AND U58016 ( .A(n46734), .B(n46733), .Z(n46735) );
  NANDN U58017 ( .A(n46736), .B(n46735), .Z(n46737) );
  NAND U58018 ( .A(n46738), .B(n46737), .Z(n46739) );
  NAND U58019 ( .A(n46740), .B(n46739), .Z(n46741) );
  AND U58020 ( .A(n46741), .B(n51002), .Z(n46742) );
  NANDN U58021 ( .A(x[6658]), .B(y[6658]), .Z(n59383) );
  AND U58022 ( .A(n46742), .B(n59383), .Z(n46746) );
  AND U58023 ( .A(n46744), .B(n46743), .Z(n46745) );
  NANDN U58024 ( .A(n46746), .B(n46745), .Z(n46747) );
  NAND U58025 ( .A(n46748), .B(n46747), .Z(n46749) );
  NAND U58026 ( .A(n46750), .B(n46749), .Z(n46752) );
  IV U58027 ( .A(n46751), .Z(n51000) );
  AND U58028 ( .A(n46752), .B(n51000), .Z(n46753) );
  NANDN U58029 ( .A(x[6662]), .B(y[6662]), .Z(n59389) );
  AND U58030 ( .A(n46753), .B(n59389), .Z(n46757) );
  AND U58031 ( .A(n46755), .B(n46754), .Z(n46756) );
  NANDN U58032 ( .A(n46757), .B(n46756), .Z(n46758) );
  NAND U58033 ( .A(n46759), .B(n46758), .Z(n46760) );
  NAND U58034 ( .A(n46761), .B(n46760), .Z(n46762) );
  AND U58035 ( .A(n46762), .B(n50998), .Z(n46763) );
  NANDN U58036 ( .A(x[6666]), .B(y[6666]), .Z(n59392) );
  AND U58037 ( .A(n46763), .B(n59392), .Z(n46767) );
  AND U58038 ( .A(n46765), .B(n46764), .Z(n46766) );
  NANDN U58039 ( .A(n46767), .B(n46766), .Z(n46768) );
  NAND U58040 ( .A(n46769), .B(n46768), .Z(n46770) );
  AND U58041 ( .A(n46771), .B(n46770), .Z(n46772) );
  OR U58042 ( .A(n46773), .B(n46772), .Z(n46774) );
  NAND U58043 ( .A(n46775), .B(n46774), .Z(n46776) );
  NANDN U58044 ( .A(n46777), .B(n46776), .Z(n46778) );
  AND U58045 ( .A(n46779), .B(n46778), .Z(n46780) );
  OR U58046 ( .A(n46781), .B(n46780), .Z(n46782) );
  NAND U58047 ( .A(n46783), .B(n46782), .Z(n46784) );
  NANDN U58048 ( .A(n46785), .B(n46784), .Z(n46786) );
  NAND U58049 ( .A(n46787), .B(n46786), .Z(n46788) );
  AND U58050 ( .A(n46788), .B(n50993), .Z(n46789) );
  NANDN U58051 ( .A(x[6678]), .B(y[6678]), .Z(n59405) );
  AND U58052 ( .A(n46789), .B(n59405), .Z(n46790) );
  OR U58053 ( .A(n46791), .B(n46790), .Z(n46792) );
  NAND U58054 ( .A(n46793), .B(n46792), .Z(n46794) );
  NAND U58055 ( .A(n46795), .B(n46794), .Z(n46796) );
  AND U58056 ( .A(n46796), .B(n50992), .Z(n46797) );
  NANDN U58057 ( .A(x[6682]), .B(y[6682]), .Z(n59409) );
  AND U58058 ( .A(n46797), .B(n59409), .Z(n46801) );
  AND U58059 ( .A(n46799), .B(n46798), .Z(n46800) );
  NANDN U58060 ( .A(n46801), .B(n46800), .Z(n46802) );
  NAND U58061 ( .A(n46803), .B(n46802), .Z(n46804) );
  AND U58062 ( .A(n46805), .B(n46804), .Z(n46806) );
  ANDN U58063 ( .B(n50989), .A(n46806), .Z(n46807) );
  NANDN U58064 ( .A(x[6686]), .B(y[6686]), .Z(n59415) );
  AND U58065 ( .A(n46807), .B(n59415), .Z(n46808) );
  OR U58066 ( .A(n46809), .B(n46808), .Z(n46810) );
  NAND U58067 ( .A(n46811), .B(n46810), .Z(n46812) );
  NAND U58068 ( .A(n46813), .B(n46812), .Z(n46814) );
  AND U58069 ( .A(n46814), .B(n59419), .Z(n46815) );
  NANDN U58070 ( .A(x[6690]), .B(y[6690]), .Z(n50988) );
  AND U58071 ( .A(n46815), .B(n50988), .Z(n46819) );
  AND U58072 ( .A(n46817), .B(n46816), .Z(n46818) );
  NANDN U58073 ( .A(n46819), .B(n46818), .Z(n46820) );
  NAND U58074 ( .A(n46821), .B(n46820), .Z(n46822) );
  NAND U58075 ( .A(n46823), .B(n46822), .Z(n46824) );
  AND U58076 ( .A(n46824), .B(n59423), .Z(n46825) );
  NANDN U58077 ( .A(x[6694]), .B(y[6694]), .Z(n50986) );
  AND U58078 ( .A(n46825), .B(n50986), .Z(n46829) );
  AND U58079 ( .A(n46827), .B(n46826), .Z(n46828) );
  NANDN U58080 ( .A(n46829), .B(n46828), .Z(n46830) );
  NAND U58081 ( .A(n46831), .B(n46830), .Z(n46832) );
  NAND U58082 ( .A(n46833), .B(n46832), .Z(n46834) );
  AND U58083 ( .A(n46834), .B(n59429), .Z(n46835) );
  NANDN U58084 ( .A(x[6698]), .B(y[6698]), .Z(n59427) );
  AND U58085 ( .A(n46835), .B(n59427), .Z(n46839) );
  AND U58086 ( .A(n46837), .B(n46836), .Z(n46838) );
  NANDN U58087 ( .A(n46839), .B(n46838), .Z(n46840) );
  NAND U58088 ( .A(n46841), .B(n46840), .Z(n46842) );
  NAND U58089 ( .A(n46843), .B(n46842), .Z(n46844) );
  AND U58090 ( .A(n46844), .B(n59435), .Z(n46845) );
  NANDN U58091 ( .A(x[6702]), .B(y[6702]), .Z(n59433) );
  AND U58092 ( .A(n46845), .B(n59433), .Z(n46849) );
  AND U58093 ( .A(n46847), .B(n46846), .Z(n46848) );
  NANDN U58094 ( .A(n46849), .B(n46848), .Z(n46850) );
  NAND U58095 ( .A(n46851), .B(n46850), .Z(n46852) );
  NAND U58096 ( .A(n46853), .B(n46852), .Z(n46854) );
  AND U58097 ( .A(n46854), .B(n50982), .Z(n46855) );
  NANDN U58098 ( .A(x[6706]), .B(y[6706]), .Z(n59439) );
  AND U58099 ( .A(n46855), .B(n59439), .Z(n46859) );
  AND U58100 ( .A(n46857), .B(n46856), .Z(n46858) );
  NANDN U58101 ( .A(n46859), .B(n46858), .Z(n46860) );
  NAND U58102 ( .A(n46861), .B(n46860), .Z(n46862) );
  NAND U58103 ( .A(n46863), .B(n46862), .Z(n46864) );
  AND U58104 ( .A(n46864), .B(n50981), .Z(n46865) );
  NANDN U58105 ( .A(x[6710]), .B(y[6710]), .Z(n59444) );
  AND U58106 ( .A(n46865), .B(n59444), .Z(n46869) );
  AND U58107 ( .A(n46867), .B(n46866), .Z(n46868) );
  NANDN U58108 ( .A(n46869), .B(n46868), .Z(n46870) );
  NAND U58109 ( .A(n46871), .B(n46870), .Z(n46872) );
  AND U58110 ( .A(n46873), .B(n46872), .Z(n46874) );
  OR U58111 ( .A(n46875), .B(n46874), .Z(n46876) );
  NAND U58112 ( .A(n46877), .B(n46876), .Z(n46878) );
  NANDN U58113 ( .A(n46879), .B(n46878), .Z(n46880) );
  NAND U58114 ( .A(n46881), .B(n46880), .Z(n46882) );
  AND U58115 ( .A(n46883), .B(n46882), .Z(n46887) );
  AND U58116 ( .A(n46885), .B(n46884), .Z(n46886) );
  NANDN U58117 ( .A(n46887), .B(n46886), .Z(n46888) );
  NAND U58118 ( .A(n46889), .B(n46888), .Z(n46890) );
  AND U58119 ( .A(n46891), .B(n46890), .Z(n46893) );
  NANDN U58120 ( .A(x[6722]), .B(y[6722]), .Z(n50977) );
  AND U58121 ( .A(n50977), .B(n59458), .Z(n46892) );
  NANDN U58122 ( .A(n46893), .B(n46892), .Z(n46894) );
  NANDN U58123 ( .A(n46895), .B(n46894), .Z(n46896) );
  AND U58124 ( .A(n59461), .B(n46896), .Z(n46897) );
  NANDN U58125 ( .A(x[6724]), .B(y[6724]), .Z(n59459) );
  NAND U58126 ( .A(n46897), .B(n59459), .Z(n46898) );
  NAND U58127 ( .A(n46899), .B(n46898), .Z(n46900) );
  AND U58128 ( .A(n46900), .B(n59464), .Z(n46901) );
  NANDN U58129 ( .A(x[6726]), .B(y[6726]), .Z(n59462) );
  AND U58130 ( .A(n46901), .B(n59462), .Z(n46905) );
  AND U58131 ( .A(n46903), .B(n46902), .Z(n46904) );
  NANDN U58132 ( .A(n46905), .B(n46904), .Z(n46906) );
  NAND U58133 ( .A(n46907), .B(n46906), .Z(n46908) );
  NAND U58134 ( .A(n46909), .B(n46908), .Z(n46910) );
  AND U58135 ( .A(n46910), .B(n50973), .Z(n46911) );
  NANDN U58136 ( .A(x[6730]), .B(y[6730]), .Z(n59468) );
  AND U58137 ( .A(n46911), .B(n59468), .Z(n46915) );
  AND U58138 ( .A(n46913), .B(n46912), .Z(n46914) );
  NANDN U58139 ( .A(n46915), .B(n46914), .Z(n46916) );
  NAND U58140 ( .A(n46917), .B(n46916), .Z(n46918) );
  NAND U58141 ( .A(n46919), .B(n46918), .Z(n46921) );
  AND U58142 ( .A(n46921), .B(n46920), .Z(n46922) );
  NANDN U58143 ( .A(x[6734]), .B(y[6734]), .Z(n59472) );
  AND U58144 ( .A(n46922), .B(n59472), .Z(n46923) );
  OR U58145 ( .A(n46924), .B(n46923), .Z(n46925) );
  NAND U58146 ( .A(n46926), .B(n46925), .Z(n46927) );
  NAND U58147 ( .A(n46928), .B(n46927), .Z(n46929) );
  AND U58148 ( .A(n46929), .B(n59479), .Z(n46930) );
  NANDN U58149 ( .A(x[6738]), .B(y[6738]), .Z(n59477) );
  AND U58150 ( .A(n46930), .B(n59477), .Z(n46934) );
  AND U58151 ( .A(n46932), .B(n46931), .Z(n46933) );
  NANDN U58152 ( .A(n46934), .B(n46933), .Z(n46935) );
  NAND U58153 ( .A(n46936), .B(n46935), .Z(n46937) );
  AND U58154 ( .A(n46938), .B(n46937), .Z(n46940) );
  NANDN U58155 ( .A(x[6742]), .B(y[6742]), .Z(n50971) );
  AND U58156 ( .A(n59483), .B(n50971), .Z(n46939) );
  NANDN U58157 ( .A(n46940), .B(n46939), .Z(n46941) );
  NAND U58158 ( .A(n46942), .B(n46941), .Z(n46943) );
  OR U58159 ( .A(n46944), .B(n46943), .Z(n46945) );
  NAND U58160 ( .A(n46946), .B(n46945), .Z(n46947) );
  NAND U58161 ( .A(n46948), .B(n46947), .Z(n46949) );
  AND U58162 ( .A(n46949), .B(n59490), .Z(n46950) );
  NANDN U58163 ( .A(x[6746]), .B(y[6746]), .Z(n59487) );
  AND U58164 ( .A(n46950), .B(n59487), .Z(n46954) );
  AND U58165 ( .A(n46952), .B(n46951), .Z(n46953) );
  NANDN U58166 ( .A(n46954), .B(n46953), .Z(n46955) );
  NAND U58167 ( .A(n46956), .B(n46955), .Z(n46957) );
  AND U58168 ( .A(n46958), .B(n46957), .Z(n46959) );
  OR U58169 ( .A(n46960), .B(n46959), .Z(n46961) );
  NAND U58170 ( .A(n46962), .B(n46961), .Z(n46963) );
  NANDN U58171 ( .A(n46964), .B(n46963), .Z(n46965) );
  NAND U58172 ( .A(n46966), .B(n46965), .Z(n46967) );
  AND U58173 ( .A(n46967), .B(n50969), .Z(n46968) );
  NANDN U58174 ( .A(x[6754]), .B(y[6754]), .Z(n59499) );
  AND U58175 ( .A(n46968), .B(n59499), .Z(n46972) );
  AND U58176 ( .A(n46970), .B(n46969), .Z(n46971) );
  NANDN U58177 ( .A(n46972), .B(n46971), .Z(n46973) );
  NAND U58178 ( .A(n46974), .B(n46973), .Z(n46975) );
  NAND U58179 ( .A(n46976), .B(n46975), .Z(n46977) );
  AND U58180 ( .A(n46977), .B(n59507), .Z(n46978) );
  NANDN U58181 ( .A(x[6758]), .B(y[6758]), .Z(n59505) );
  AND U58182 ( .A(n46978), .B(n59505), .Z(n46982) );
  AND U58183 ( .A(n46980), .B(n46979), .Z(n46981) );
  NANDN U58184 ( .A(n46982), .B(n46981), .Z(n46983) );
  NAND U58185 ( .A(n46984), .B(n46983), .Z(n46985) );
  NAND U58186 ( .A(n46986), .B(n46985), .Z(n46987) );
  AND U58187 ( .A(n46987), .B(n59512), .Z(n46988) );
  NANDN U58188 ( .A(x[6762]), .B(y[6762]), .Z(n59510) );
  AND U58189 ( .A(n46988), .B(n59510), .Z(n46992) );
  AND U58190 ( .A(n46990), .B(n46989), .Z(n46991) );
  NANDN U58191 ( .A(n46992), .B(n46991), .Z(n46993) );
  NAND U58192 ( .A(n46994), .B(n46993), .Z(n46995) );
  NAND U58193 ( .A(n46996), .B(n46995), .Z(n46997) );
  AND U58194 ( .A(n46997), .B(n59517), .Z(n46998) );
  NANDN U58195 ( .A(x[6766]), .B(y[6766]), .Z(n50966) );
  AND U58196 ( .A(n46998), .B(n50966), .Z(n47002) );
  AND U58197 ( .A(n47000), .B(n46999), .Z(n47001) );
  NANDN U58198 ( .A(n47002), .B(n47001), .Z(n47003) );
  NAND U58199 ( .A(n47004), .B(n47003), .Z(n47005) );
  AND U58200 ( .A(n47006), .B(n47005), .Z(n47007) );
  ANDN U58201 ( .B(n59521), .A(n47007), .Z(n47008) );
  NAND U58202 ( .A(n50964), .B(n47008), .Z(n47009) );
  NANDN U58203 ( .A(n47010), .B(n47009), .Z(n47011) );
  AND U58204 ( .A(n47011), .B(n59524), .Z(n47012) );
  NANDN U58205 ( .A(x[6772]), .B(y[6772]), .Z(n59522) );
  NAND U58206 ( .A(n47012), .B(n59522), .Z(n47013) );
  NAND U58207 ( .A(n47014), .B(n47013), .Z(n47015) );
  AND U58208 ( .A(n47015), .B(n59527), .Z(n47016) );
  NANDN U58209 ( .A(x[6774]), .B(y[6774]), .Z(n59525) );
  AND U58210 ( .A(n47016), .B(n59525), .Z(n47020) );
  AND U58211 ( .A(n47018), .B(n47017), .Z(n47019) );
  NANDN U58212 ( .A(n47020), .B(n47019), .Z(n47021) );
  NAND U58213 ( .A(n47022), .B(n47021), .Z(n47023) );
  NAND U58214 ( .A(n47024), .B(n47023), .Z(n47025) );
  AND U58215 ( .A(n47025), .B(n50962), .Z(n47026) );
  NANDN U58216 ( .A(x[6778]), .B(y[6778]), .Z(n59531) );
  AND U58217 ( .A(n47026), .B(n59531), .Z(n47030) );
  AND U58218 ( .A(n47028), .B(n47027), .Z(n47029) );
  NANDN U58219 ( .A(n47030), .B(n47029), .Z(n47031) );
  NAND U58220 ( .A(n47032), .B(n47031), .Z(n47033) );
  NAND U58221 ( .A(n47034), .B(n47033), .Z(n47035) );
  AND U58222 ( .A(n47035), .B(n50960), .Z(n47036) );
  NANDN U58223 ( .A(x[6782]), .B(y[6782]), .Z(n59537) );
  AND U58224 ( .A(n47036), .B(n59537), .Z(n47040) );
  AND U58225 ( .A(n47038), .B(n47037), .Z(n47039) );
  NANDN U58226 ( .A(n47040), .B(n47039), .Z(n47041) );
  NAND U58227 ( .A(n47042), .B(n47041), .Z(n47043) );
  NAND U58228 ( .A(n47044), .B(n47043), .Z(n47045) );
  AND U58229 ( .A(n47045), .B(n59543), .Z(n47046) );
  NANDN U58230 ( .A(x[6786]), .B(y[6786]), .Z(n59541) );
  AND U58231 ( .A(n47046), .B(n59541), .Z(n47050) );
  AND U58232 ( .A(n47048), .B(n47047), .Z(n47049) );
  NANDN U58233 ( .A(n47050), .B(n47049), .Z(n47051) );
  NAND U58234 ( .A(n47052), .B(n47051), .Z(n47053) );
  NAND U58235 ( .A(n47054), .B(n47053), .Z(n47055) );
  AND U58236 ( .A(n47055), .B(n59548), .Z(n47056) );
  NANDN U58237 ( .A(x[6790]), .B(y[6790]), .Z(n59546) );
  NAND U58238 ( .A(n47056), .B(n59546), .Z(n47057) );
  NAND U58239 ( .A(n47058), .B(n47057), .Z(n47059) );
  ANDN U58240 ( .B(y[6792]), .A(x[6792]), .Z(n59549) );
  ANDN U58241 ( .B(n47059), .A(n59549), .Z(n47060) );
  NAND U58242 ( .A(n50957), .B(n47060), .Z(n47061) );
  NAND U58243 ( .A(n47062), .B(n47061), .Z(n47063) );
  AND U58244 ( .A(n47063), .B(n59554), .Z(n47064) );
  NANDN U58245 ( .A(x[6794]), .B(y[6794]), .Z(n50956) );
  AND U58246 ( .A(n47064), .B(n50956), .Z(n47068) );
  AND U58247 ( .A(n47066), .B(n47065), .Z(n47067) );
  NANDN U58248 ( .A(n47068), .B(n47067), .Z(n47069) );
  NAND U58249 ( .A(n47070), .B(n47069), .Z(n47071) );
  NAND U58250 ( .A(n47072), .B(n47071), .Z(n47073) );
  AND U58251 ( .A(n47073), .B(n59558), .Z(n47074) );
  NANDN U58252 ( .A(x[6798]), .B(y[6798]), .Z(n50955) );
  AND U58253 ( .A(n47074), .B(n50955), .Z(n47078) );
  AND U58254 ( .A(n47076), .B(n47075), .Z(n47077) );
  NANDN U58255 ( .A(n47078), .B(n47077), .Z(n47079) );
  NAND U58256 ( .A(n47080), .B(n47079), .Z(n47081) );
  NAND U58257 ( .A(n47082), .B(n47081), .Z(n47083) );
  AND U58258 ( .A(n47083), .B(n59565), .Z(n47084) );
  NANDN U58259 ( .A(x[6802]), .B(y[6802]), .Z(n59562) );
  AND U58260 ( .A(n47084), .B(n59562), .Z(n47088) );
  AND U58261 ( .A(n47086), .B(n47085), .Z(n47087) );
  NANDN U58262 ( .A(n47088), .B(n47087), .Z(n47089) );
  NAND U58263 ( .A(n47090), .B(n47089), .Z(n47091) );
  NAND U58264 ( .A(n47092), .B(n47091), .Z(n47093) );
  NAND U58265 ( .A(n47094), .B(n47093), .Z(n47095) );
  NAND U58266 ( .A(n59569), .B(n47095), .Z(n47096) );
  AND U58267 ( .A(n47097), .B(n47096), .Z(n47099) );
  XNOR U58268 ( .A(y[6808]), .B(x[6808]), .Z(n47098) );
  NANDN U58269 ( .A(n47099), .B(n47098), .Z(n47100) );
  NAND U58270 ( .A(n47101), .B(n47100), .Z(n47102) );
  NAND U58271 ( .A(n47103), .B(n47102), .Z(n47104) );
  AND U58272 ( .A(n47104), .B(n59574), .Z(n47105) );
  NANDN U58273 ( .A(x[6810]), .B(y[6810]), .Z(n59572) );
  AND U58274 ( .A(n47105), .B(n59572), .Z(n47109) );
  AND U58275 ( .A(n47107), .B(n47106), .Z(n47108) );
  NANDN U58276 ( .A(n47109), .B(n47108), .Z(n47110) );
  NAND U58277 ( .A(n47111), .B(n47110), .Z(n47112) );
  AND U58278 ( .A(n47113), .B(n47112), .Z(n47114) );
  ANDN U58279 ( .B(n59581), .A(n47114), .Z(n47115) );
  NANDN U58280 ( .A(x[6814]), .B(y[6814]), .Z(n59578) );
  AND U58281 ( .A(n47115), .B(n59578), .Z(n47116) );
  OR U58282 ( .A(n47117), .B(n47116), .Z(n47118) );
  NAND U58283 ( .A(n47119), .B(n47118), .Z(n47120) );
  NAND U58284 ( .A(n47121), .B(n47120), .Z(n47122) );
  AND U58285 ( .A(n47122), .B(n59587), .Z(n47123) );
  NANDN U58286 ( .A(x[6818]), .B(y[6818]), .Z(n59585) );
  AND U58287 ( .A(n47123), .B(n59585), .Z(n47127) );
  AND U58288 ( .A(n47125), .B(n47124), .Z(n47126) );
  NANDN U58289 ( .A(n47127), .B(n47126), .Z(n47128) );
  NAND U58290 ( .A(n47129), .B(n47128), .Z(n47130) );
  NAND U58291 ( .A(n47131), .B(n47130), .Z(n47132) );
  AND U58292 ( .A(n47132), .B(n59591), .Z(n47133) );
  NANDN U58293 ( .A(x[6822]), .B(y[6822]), .Z(n50952) );
  AND U58294 ( .A(n47133), .B(n50952), .Z(n47137) );
  AND U58295 ( .A(n47135), .B(n47134), .Z(n47136) );
  NANDN U58296 ( .A(n47137), .B(n47136), .Z(n47138) );
  NAND U58297 ( .A(n47139), .B(n47138), .Z(n47140) );
  NAND U58298 ( .A(n47141), .B(n47140), .Z(n47142) );
  AND U58299 ( .A(n47142), .B(n59598), .Z(n47143) );
  NANDN U58300 ( .A(x[6826]), .B(y[6826]), .Z(n59595) );
  AND U58301 ( .A(n47143), .B(n59595), .Z(n47147) );
  AND U58302 ( .A(n47145), .B(n47144), .Z(n47146) );
  NANDN U58303 ( .A(n47147), .B(n47146), .Z(n47148) );
  NAND U58304 ( .A(n47149), .B(n47148), .Z(n47150) );
  NAND U58305 ( .A(n47151), .B(n47150), .Z(n47153) );
  AND U58306 ( .A(n47153), .B(n47152), .Z(n47154) );
  NANDN U58307 ( .A(x[6830]), .B(y[6830]), .Z(n59602) );
  AND U58308 ( .A(n47154), .B(n59602), .Z(n47158) );
  AND U58309 ( .A(n47156), .B(n47155), .Z(n47157) );
  NANDN U58310 ( .A(n47158), .B(n47157), .Z(n47159) );
  NAND U58311 ( .A(n47160), .B(n47159), .Z(n47161) );
  NAND U58312 ( .A(n47162), .B(n47161), .Z(n47164) );
  IV U58313 ( .A(n47163), .Z(n50947) );
  AND U58314 ( .A(n47164), .B(n50947), .Z(n47165) );
  NANDN U58315 ( .A(x[6834]), .B(y[6834]), .Z(n59606) );
  AND U58316 ( .A(n47165), .B(n59606), .Z(n47169) );
  AND U58317 ( .A(n47167), .B(n47166), .Z(n47168) );
  NANDN U58318 ( .A(n47169), .B(n47168), .Z(n47170) );
  NAND U58319 ( .A(n47171), .B(n47170), .Z(n47172) );
  NAND U58320 ( .A(n47173), .B(n47172), .Z(n47174) );
  AND U58321 ( .A(n47174), .B(n50946), .Z(n47176) );
  NANDN U58322 ( .A(x[6838]), .B(y[6838]), .Z(n47175) );
  AND U58323 ( .A(n47176), .B(n47175), .Z(n47180) );
  AND U58324 ( .A(n47178), .B(n47177), .Z(n47179) );
  NANDN U58325 ( .A(n47180), .B(n47179), .Z(n47181) );
  NAND U58326 ( .A(n47182), .B(n47181), .Z(n47183) );
  AND U58327 ( .A(n47184), .B(n47183), .Z(n47185) );
  ANDN U58328 ( .B(n47186), .A(n47185), .Z(n47187) );
  OR U58329 ( .A(n47188), .B(n47187), .Z(n47189) );
  NAND U58330 ( .A(n47190), .B(n47189), .Z(n47191) );
  NAND U58331 ( .A(n47192), .B(n47191), .Z(n47193) );
  AND U58332 ( .A(n47193), .B(n59617), .Z(n47194) );
  NANDN U58333 ( .A(x[6846]), .B(y[6846]), .Z(n50941) );
  AND U58334 ( .A(n47194), .B(n50941), .Z(n47198) );
  AND U58335 ( .A(n47196), .B(n47195), .Z(n47197) );
  NANDN U58336 ( .A(n47198), .B(n47197), .Z(n47199) );
  NAND U58337 ( .A(n47200), .B(n47199), .Z(n47201) );
  AND U58338 ( .A(n47202), .B(n47201), .Z(n47204) );
  NANDN U58339 ( .A(x[6850]), .B(y[6850]), .Z(n59621) );
  AND U58340 ( .A(n59621), .B(n59623), .Z(n47203) );
  NANDN U58341 ( .A(n47204), .B(n47203), .Z(n47205) );
  NANDN U58342 ( .A(n47206), .B(n47205), .Z(n47207) );
  AND U58343 ( .A(n47208), .B(n47207), .Z(n47209) );
  NANDN U58344 ( .A(x[6852]), .B(y[6852]), .Z(n59624) );
  NAND U58345 ( .A(n47209), .B(n59624), .Z(n47210) );
  AND U58346 ( .A(n47211), .B(n47210), .Z(n47212) );
  OR U58347 ( .A(n47213), .B(n47212), .Z(n47214) );
  NAND U58348 ( .A(n47215), .B(n47214), .Z(n47216) );
  NANDN U58349 ( .A(n47217), .B(n47216), .Z(n47218) );
  NAND U58350 ( .A(n47219), .B(n47218), .Z(n47220) );
  AND U58351 ( .A(n47220), .B(n50936), .Z(n47221) );
  NANDN U58352 ( .A(x[6858]), .B(y[6858]), .Z(n59631) );
  AND U58353 ( .A(n47221), .B(n59631), .Z(n47225) );
  AND U58354 ( .A(n47223), .B(n47222), .Z(n47224) );
  NANDN U58355 ( .A(n47225), .B(n47224), .Z(n47226) );
  NAND U58356 ( .A(n47227), .B(n47226), .Z(n47228) );
  NAND U58357 ( .A(n47229), .B(n47228), .Z(n47230) );
  AND U58358 ( .A(n47230), .B(n59637), .Z(n47231) );
  NANDN U58359 ( .A(x[6862]), .B(y[6862]), .Z(n59635) );
  AND U58360 ( .A(n47231), .B(n59635), .Z(n47232) );
  OR U58361 ( .A(n47233), .B(n47232), .Z(n47234) );
  NAND U58362 ( .A(n47235), .B(n47234), .Z(n47236) );
  NAND U58363 ( .A(n47237), .B(n47236), .Z(n47238) );
  AND U58364 ( .A(n47238), .B(n59644), .Z(n47239) );
  NANDN U58365 ( .A(x[6866]), .B(y[6866]), .Z(n59642) );
  AND U58366 ( .A(n47239), .B(n59642), .Z(n47243) );
  AND U58367 ( .A(n47241), .B(n47240), .Z(n47242) );
  NANDN U58368 ( .A(n47243), .B(n47242), .Z(n47244) );
  NAND U58369 ( .A(n47245), .B(n47244), .Z(n47246) );
  AND U58370 ( .A(n47247), .B(n47246), .Z(n47248) );
  NOR U58371 ( .A(n50933), .B(n47248), .Z(n47249) );
  NAND U58372 ( .A(n59648), .B(n47249), .Z(n47250) );
  NANDN U58373 ( .A(n47251), .B(n47250), .Z(n47252) );
  OR U58374 ( .A(n47253), .B(n47252), .Z(n47254) );
  NAND U58375 ( .A(n47255), .B(n47254), .Z(n47256) );
  NAND U58376 ( .A(n47257), .B(n47256), .Z(n47258) );
  AND U58377 ( .A(n47258), .B(n59652), .Z(n47259) );
  NANDN U58378 ( .A(x[6874]), .B(y[6874]), .Z(n50932) );
  AND U58379 ( .A(n47259), .B(n50932), .Z(n47260) );
  OR U58380 ( .A(n47261), .B(n47260), .Z(n47262) );
  NAND U58381 ( .A(n47263), .B(n47262), .Z(n47264) );
  NAND U58382 ( .A(n47265), .B(n47264), .Z(n47266) );
  AND U58383 ( .A(n47266), .B(n59659), .Z(n47267) );
  NANDN U58384 ( .A(x[6878]), .B(y[6878]), .Z(n59657) );
  AND U58385 ( .A(n47267), .B(n59657), .Z(n47271) );
  AND U58386 ( .A(n47269), .B(n47268), .Z(n47270) );
  NANDN U58387 ( .A(n47271), .B(n47270), .Z(n47272) );
  NAND U58388 ( .A(n47273), .B(n47272), .Z(n47274) );
  NAND U58389 ( .A(n47275), .B(n47274), .Z(n47277) );
  AND U58390 ( .A(n47277), .B(n47276), .Z(n47278) );
  NANDN U58391 ( .A(x[6882]), .B(y[6882]), .Z(n59663) );
  AND U58392 ( .A(n47278), .B(n59663), .Z(n47282) );
  AND U58393 ( .A(n47280), .B(n47279), .Z(n47281) );
  NANDN U58394 ( .A(n47282), .B(n47281), .Z(n47283) );
  NAND U58395 ( .A(n47284), .B(n47283), .Z(n47285) );
  NAND U58396 ( .A(n47286), .B(n47285), .Z(n47288) );
  IV U58397 ( .A(n47287), .Z(n50927) );
  AND U58398 ( .A(n47288), .B(n50927), .Z(n47289) );
  NANDN U58399 ( .A(x[6886]), .B(y[6886]), .Z(n59667) );
  AND U58400 ( .A(n47289), .B(n59667), .Z(n47293) );
  AND U58401 ( .A(n47291), .B(n47290), .Z(n47292) );
  NANDN U58402 ( .A(n47293), .B(n47292), .Z(n47294) );
  NAND U58403 ( .A(n47295), .B(n47294), .Z(n47296) );
  NAND U58404 ( .A(n47297), .B(n47296), .Z(n47298) );
  AND U58405 ( .A(n47298), .B(n59674), .Z(n47299) );
  NANDN U58406 ( .A(x[6890]), .B(y[6890]), .Z(n59672) );
  AND U58407 ( .A(n47299), .B(n59672), .Z(n47303) );
  AND U58408 ( .A(n47301), .B(n47300), .Z(n47302) );
  NANDN U58409 ( .A(n47303), .B(n47302), .Z(n47304) );
  NAND U58410 ( .A(n47305), .B(n47304), .Z(n47306) );
  NAND U58411 ( .A(n47307), .B(n47306), .Z(n47308) );
  AND U58412 ( .A(n47308), .B(n59679), .Z(n47309) );
  NANDN U58413 ( .A(x[6894]), .B(y[6894]), .Z(n59677) );
  AND U58414 ( .A(n47309), .B(n59677), .Z(n47313) );
  AND U58415 ( .A(n47311), .B(n47310), .Z(n47312) );
  NANDN U58416 ( .A(n47313), .B(n47312), .Z(n47314) );
  NAND U58417 ( .A(n47315), .B(n47314), .Z(n47316) );
  NAND U58418 ( .A(n47317), .B(n47316), .Z(n47318) );
  AND U58419 ( .A(n47318), .B(n59683), .Z(n47319) );
  NANDN U58420 ( .A(x[6898]), .B(y[6898]), .Z(n50924) );
  AND U58421 ( .A(n47319), .B(n50924), .Z(n47323) );
  AND U58422 ( .A(n47321), .B(n47320), .Z(n47322) );
  NANDN U58423 ( .A(n47323), .B(n47322), .Z(n47324) );
  NAND U58424 ( .A(n47325), .B(n47324), .Z(n47326) );
  NAND U58425 ( .A(n47327), .B(n47326), .Z(n47328) );
  AND U58426 ( .A(n47329), .B(n47328), .Z(n47333) );
  AND U58427 ( .A(n47331), .B(n47330), .Z(n47332) );
  NANDN U58428 ( .A(n47333), .B(n47332), .Z(n47334) );
  NAND U58429 ( .A(n47335), .B(n47334), .Z(n47336) );
  NAND U58430 ( .A(n47337), .B(n47336), .Z(n47339) );
  AND U58431 ( .A(n47339), .B(n47338), .Z(n47340) );
  NANDN U58432 ( .A(x[6906]), .B(y[6906]), .Z(n50922) );
  AND U58433 ( .A(n47340), .B(n50922), .Z(n47344) );
  AND U58434 ( .A(n47342), .B(n47341), .Z(n47343) );
  NANDN U58435 ( .A(n47344), .B(n47343), .Z(n47345) );
  NAND U58436 ( .A(n47346), .B(n47345), .Z(n47347) );
  NAND U58437 ( .A(n47348), .B(n47347), .Z(n47349) );
  AND U58438 ( .A(n47349), .B(n59699), .Z(n47350) );
  NANDN U58439 ( .A(x[6910]), .B(y[6910]), .Z(n59697) );
  AND U58440 ( .A(n47350), .B(n59697), .Z(n47354) );
  AND U58441 ( .A(n47352), .B(n47351), .Z(n47353) );
  NANDN U58442 ( .A(n47354), .B(n47353), .Z(n47355) );
  NAND U58443 ( .A(n47356), .B(n47355), .Z(n47357) );
  NAND U58444 ( .A(n47358), .B(n47357), .Z(n47359) );
  AND U58445 ( .A(n47359), .B(n59705), .Z(n47360) );
  NANDN U58446 ( .A(x[6914]), .B(y[6914]), .Z(n50919) );
  AND U58447 ( .A(n47360), .B(n50919), .Z(n47364) );
  AND U58448 ( .A(n47362), .B(n47361), .Z(n47363) );
  NANDN U58449 ( .A(n47364), .B(n47363), .Z(n47365) );
  NAND U58450 ( .A(n47366), .B(n47365), .Z(n47367) );
  NAND U58451 ( .A(n47368), .B(n47367), .Z(n47369) );
  AND U58452 ( .A(n47369), .B(n59711), .Z(n47370) );
  NANDN U58453 ( .A(x[6918]), .B(y[6918]), .Z(n59709) );
  AND U58454 ( .A(n47370), .B(n59709), .Z(n47374) );
  AND U58455 ( .A(n47372), .B(n47371), .Z(n47373) );
  NANDN U58456 ( .A(n47374), .B(n47373), .Z(n47375) );
  NAND U58457 ( .A(n47376), .B(n47375), .Z(n47377) );
  NAND U58458 ( .A(n47378), .B(n47377), .Z(n47379) );
  AND U58459 ( .A(n47379), .B(n50915), .Z(n47380) );
  NANDN U58460 ( .A(x[6922]), .B(y[6922]), .Z(n59715) );
  AND U58461 ( .A(n47380), .B(n59715), .Z(n47384) );
  AND U58462 ( .A(n47382), .B(n47381), .Z(n47383) );
  NANDN U58463 ( .A(n47384), .B(n47383), .Z(n47385) );
  NAND U58464 ( .A(n47386), .B(n47385), .Z(n47387) );
  AND U58465 ( .A(n47388), .B(n47387), .Z(n47390) );
  NANDN U58466 ( .A(x[6926]), .B(y[6926]), .Z(n59720) );
  AND U58467 ( .A(n59720), .B(n50913), .Z(n47389) );
  NANDN U58468 ( .A(n47390), .B(n47389), .Z(n47391) );
  NANDN U58469 ( .A(n47392), .B(n47391), .Z(n47393) );
  AND U58470 ( .A(n59723), .B(n47393), .Z(n47394) );
  NANDN U58471 ( .A(x[6928]), .B(y[6928]), .Z(n50914) );
  NAND U58472 ( .A(n47394), .B(n50914), .Z(n47395) );
  NAND U58473 ( .A(n47396), .B(n47395), .Z(n47397) );
  AND U58474 ( .A(n47397), .B(n59726), .Z(n47398) );
  NANDN U58475 ( .A(x[6930]), .B(y[6930]), .Z(n59724) );
  AND U58476 ( .A(n47398), .B(n59724), .Z(n47402) );
  AND U58477 ( .A(n47400), .B(n47399), .Z(n47401) );
  NANDN U58478 ( .A(n47402), .B(n47401), .Z(n47403) );
  NAND U58479 ( .A(n47404), .B(n47403), .Z(n47405) );
  NAND U58480 ( .A(n47406), .B(n47405), .Z(n47407) );
  AND U58481 ( .A(n47407), .B(n59731), .Z(n47408) );
  NANDN U58482 ( .A(x[6934]), .B(y[6934]), .Z(n59728) );
  AND U58483 ( .A(n47408), .B(n59728), .Z(n47412) );
  AND U58484 ( .A(n47410), .B(n47409), .Z(n47411) );
  NANDN U58485 ( .A(n47412), .B(n47411), .Z(n47413) );
  NAND U58486 ( .A(n47414), .B(n47413), .Z(n47415) );
  NAND U58487 ( .A(n47416), .B(n47415), .Z(n47418) );
  AND U58488 ( .A(n47418), .B(n47417), .Z(n47419) );
  NANDN U58489 ( .A(x[6938]), .B(y[6938]), .Z(n50909) );
  AND U58490 ( .A(n47419), .B(n50909), .Z(n47423) );
  AND U58491 ( .A(n47421), .B(n47420), .Z(n47422) );
  NANDN U58492 ( .A(n47423), .B(n47422), .Z(n47424) );
  NAND U58493 ( .A(n47425), .B(n47424), .Z(n47426) );
  NAND U58494 ( .A(n47427), .B(n47426), .Z(n47428) );
  AND U58495 ( .A(n47428), .B(n59741), .Z(n47429) );
  NANDN U58496 ( .A(x[6942]), .B(y[6942]), .Z(n59738) );
  AND U58497 ( .A(n47429), .B(n59738), .Z(n47433) );
  AND U58498 ( .A(n47431), .B(n47430), .Z(n47432) );
  NANDN U58499 ( .A(n47433), .B(n47432), .Z(n47434) );
  NAND U58500 ( .A(n47435), .B(n47434), .Z(n47436) );
  NAND U58501 ( .A(n47437), .B(n47436), .Z(n47438) );
  AND U58502 ( .A(n47438), .B(n59747), .Z(n47439) );
  NANDN U58503 ( .A(x[6946]), .B(y[6946]), .Z(n59745) );
  AND U58504 ( .A(n47439), .B(n59745), .Z(n47443) );
  AND U58505 ( .A(n47441), .B(n47440), .Z(n47442) );
  NANDN U58506 ( .A(n47443), .B(n47442), .Z(n47444) );
  NAND U58507 ( .A(n47445), .B(n47444), .Z(n47446) );
  NAND U58508 ( .A(n47447), .B(n47446), .Z(n47448) );
  AND U58509 ( .A(n47448), .B(n50907), .Z(n47449) );
  NANDN U58510 ( .A(x[6950]), .B(y[6950]), .Z(n59752) );
  AND U58511 ( .A(n47449), .B(n59752), .Z(n47453) );
  AND U58512 ( .A(n47451), .B(n47450), .Z(n47452) );
  NANDN U58513 ( .A(n47453), .B(n47452), .Z(n47454) );
  NAND U58514 ( .A(n47455), .B(n47454), .Z(n47456) );
  NAND U58515 ( .A(n47457), .B(n47456), .Z(n47459) );
  AND U58516 ( .A(n47459), .B(n47458), .Z(n47460) );
  NANDN U58517 ( .A(x[6954]), .B(y[6954]), .Z(n59756) );
  AND U58518 ( .A(n47460), .B(n59756), .Z(n47464) );
  AND U58519 ( .A(n47462), .B(n47461), .Z(n47463) );
  NANDN U58520 ( .A(n47464), .B(n47463), .Z(n47465) );
  NAND U58521 ( .A(n47466), .B(n47465), .Z(n47467) );
  NAND U58522 ( .A(n47468), .B(n47467), .Z(n47469) );
  AND U58523 ( .A(n47469), .B(n50906), .Z(n47470) );
  NANDN U58524 ( .A(x[6958]), .B(y[6958]), .Z(n59761) );
  AND U58525 ( .A(n47470), .B(n59761), .Z(n47474) );
  AND U58526 ( .A(n47472), .B(n47471), .Z(n47473) );
  NANDN U58527 ( .A(n47474), .B(n47473), .Z(n47475) );
  NAND U58528 ( .A(n47476), .B(n47475), .Z(n47477) );
  NAND U58529 ( .A(n47478), .B(n47477), .Z(n47479) );
  AND U58530 ( .A(n47479), .B(n59765), .Z(n47480) );
  NANDN U58531 ( .A(x[6962]), .B(y[6962]), .Z(n50902) );
  AND U58532 ( .A(n47480), .B(n50902), .Z(n47484) );
  AND U58533 ( .A(n47482), .B(n47481), .Z(n47483) );
  NANDN U58534 ( .A(n47484), .B(n47483), .Z(n47485) );
  NAND U58535 ( .A(n47486), .B(n47485), .Z(n47487) );
  NAND U58536 ( .A(n47488), .B(n47487), .Z(n47489) );
  AND U58537 ( .A(n47489), .B(n59769), .Z(n47490) );
  NANDN U58538 ( .A(x[6966]), .B(y[6966]), .Z(n50901) );
  AND U58539 ( .A(n47490), .B(n50901), .Z(n47494) );
  AND U58540 ( .A(n47492), .B(n47491), .Z(n47493) );
  NANDN U58541 ( .A(n47494), .B(n47493), .Z(n47495) );
  NAND U58542 ( .A(n47496), .B(n47495), .Z(n47497) );
  NAND U58543 ( .A(n47498), .B(n47497), .Z(n47499) );
  AND U58544 ( .A(n47499), .B(n59775), .Z(n47500) );
  NANDN U58545 ( .A(x[6970]), .B(y[6970]), .Z(n59773) );
  AND U58546 ( .A(n47500), .B(n59773), .Z(n47504) );
  AND U58547 ( .A(n47502), .B(n47501), .Z(n47503) );
  NANDN U58548 ( .A(n47504), .B(n47503), .Z(n47505) );
  NAND U58549 ( .A(n47506), .B(n47505), .Z(n47507) );
  AND U58550 ( .A(n47508), .B(n47507), .Z(n47509) );
  ANDN U58551 ( .B(n50898), .A(n47509), .Z(n47510) );
  NAND U58552 ( .A(n59780), .B(n47510), .Z(n47511) );
  NANDN U58553 ( .A(n47512), .B(n47511), .Z(n47513) );
  AND U58554 ( .A(n47513), .B(n59783), .Z(n47514) );
  NANDN U58555 ( .A(x[6976]), .B(y[6976]), .Z(n50899) );
  NAND U58556 ( .A(n47514), .B(n50899), .Z(n47515) );
  NAND U58557 ( .A(n47516), .B(n47515), .Z(n47517) );
  AND U58558 ( .A(n47517), .B(n50897), .Z(n47518) );
  NANDN U58559 ( .A(x[6978]), .B(y[6978]), .Z(n59784) );
  AND U58560 ( .A(n47518), .B(n59784), .Z(n47522) );
  AND U58561 ( .A(n47520), .B(n47519), .Z(n47521) );
  NANDN U58562 ( .A(n47522), .B(n47521), .Z(n47523) );
  NAND U58563 ( .A(n47524), .B(n47523), .Z(n47525) );
  NAND U58564 ( .A(n47526), .B(n47525), .Z(n47527) );
  AND U58565 ( .A(n47527), .B(n59790), .Z(n47528) );
  NANDN U58566 ( .A(x[6982]), .B(y[6982]), .Z(n59788) );
  AND U58567 ( .A(n47528), .B(n59788), .Z(n47532) );
  AND U58568 ( .A(n47530), .B(n47529), .Z(n47531) );
  NANDN U58569 ( .A(n47532), .B(n47531), .Z(n47533) );
  NAND U58570 ( .A(n47534), .B(n47533), .Z(n47535) );
  NAND U58571 ( .A(n47536), .B(n47535), .Z(n47537) );
  AND U58572 ( .A(n47537), .B(n59797), .Z(n47538) );
  NANDN U58573 ( .A(x[6986]), .B(y[6986]), .Z(n59795) );
  AND U58574 ( .A(n47538), .B(n59795), .Z(n47542) );
  AND U58575 ( .A(n47540), .B(n47539), .Z(n47541) );
  NANDN U58576 ( .A(n47542), .B(n47541), .Z(n47543) );
  NAND U58577 ( .A(n47544), .B(n47543), .Z(n47545) );
  NAND U58578 ( .A(n47546), .B(n47545), .Z(n47547) );
  AND U58579 ( .A(n47547), .B(n59801), .Z(n47548) );
  NANDN U58580 ( .A(x[6990]), .B(y[6990]), .Z(n50894) );
  AND U58581 ( .A(n47548), .B(n50894), .Z(n47552) );
  AND U58582 ( .A(n47550), .B(n47549), .Z(n47551) );
  NANDN U58583 ( .A(n47552), .B(n47551), .Z(n47553) );
  NAND U58584 ( .A(n47554), .B(n47553), .Z(n47555) );
  NAND U58585 ( .A(n47556), .B(n47555), .Z(n47557) );
  AND U58586 ( .A(n47557), .B(n59806), .Z(n47558) );
  NANDN U58587 ( .A(x[6994]), .B(y[6994]), .Z(n50892) );
  AND U58588 ( .A(n47558), .B(n50892), .Z(n47559) );
  OR U58589 ( .A(n47560), .B(n47559), .Z(n47561) );
  AND U58590 ( .A(n47562), .B(n47561), .Z(n47563) );
  OR U58591 ( .A(n47564), .B(n47563), .Z(n47565) );
  NAND U58592 ( .A(n47566), .B(n47565), .Z(n47567) );
  NANDN U58593 ( .A(n47568), .B(n47567), .Z(n47570) );
  OR U58594 ( .A(n47570), .B(n47569), .Z(n47571) );
  NAND U58595 ( .A(n47572), .B(n47571), .Z(n47573) );
  NAND U58596 ( .A(n47574), .B(n47573), .Z(n47575) );
  AND U58597 ( .A(n47575), .B(n59815), .Z(n47576) );
  NANDN U58598 ( .A(x[7002]), .B(y[7002]), .Z(n59813) );
  AND U58599 ( .A(n47576), .B(n59813), .Z(n47577) );
  OR U58600 ( .A(n47578), .B(n47577), .Z(n47579) );
  NAND U58601 ( .A(n47580), .B(n47579), .Z(n47581) );
  NAND U58602 ( .A(n47582), .B(n47581), .Z(n47583) );
  AND U58603 ( .A(n47583), .B(n59821), .Z(n47584) );
  NANDN U58604 ( .A(x[7006]), .B(y[7006]), .Z(n50888) );
  AND U58605 ( .A(n47584), .B(n50888), .Z(n47588) );
  AND U58606 ( .A(n47586), .B(n47585), .Z(n47587) );
  NANDN U58607 ( .A(n47588), .B(n47587), .Z(n47589) );
  NAND U58608 ( .A(n47590), .B(n47589), .Z(n47591) );
  NAND U58609 ( .A(n47592), .B(n47591), .Z(n47593) );
  AND U58610 ( .A(n47593), .B(n59828), .Z(n47594) );
  NANDN U58611 ( .A(x[7010]), .B(y[7010]), .Z(n59826) );
  AND U58612 ( .A(n47594), .B(n59826), .Z(n47598) );
  AND U58613 ( .A(n47596), .B(n47595), .Z(n47597) );
  NANDN U58614 ( .A(n47598), .B(n47597), .Z(n47599) );
  NAND U58615 ( .A(n47600), .B(n47599), .Z(n47601) );
  NAND U58616 ( .A(n47602), .B(n47601), .Z(n47603) );
  AND U58617 ( .A(n47603), .B(n50886), .Z(n47604) );
  NANDN U58618 ( .A(x[7014]), .B(y[7014]), .Z(n59832) );
  AND U58619 ( .A(n47604), .B(n59832), .Z(n47608) );
  AND U58620 ( .A(n47606), .B(n47605), .Z(n47607) );
  NANDN U58621 ( .A(n47608), .B(n47607), .Z(n47609) );
  NAND U58622 ( .A(n47610), .B(n47609), .Z(n47611) );
  NAND U58623 ( .A(n47612), .B(n47611), .Z(n47613) );
  AND U58624 ( .A(n47613), .B(n50884), .Z(n47614) );
  NANDN U58625 ( .A(x[7018]), .B(y[7018]), .Z(n59836) );
  AND U58626 ( .A(n47614), .B(n59836), .Z(n47618) );
  AND U58627 ( .A(n47616), .B(n47615), .Z(n47617) );
  NANDN U58628 ( .A(n47618), .B(n47617), .Z(n47619) );
  NAND U58629 ( .A(n47620), .B(n47619), .Z(n47621) );
  NAND U58630 ( .A(n47622), .B(n47621), .Z(n47623) );
  AND U58631 ( .A(n47623), .B(n59842), .Z(n47624) );
  NANDN U58632 ( .A(x[7022]), .B(y[7022]), .Z(n59840) );
  AND U58633 ( .A(n47624), .B(n59840), .Z(n47628) );
  AND U58634 ( .A(n47626), .B(n47625), .Z(n47627) );
  NANDN U58635 ( .A(n47628), .B(n47627), .Z(n47629) );
  NAND U58636 ( .A(n47630), .B(n47629), .Z(n47631) );
  NAND U58637 ( .A(n47632), .B(n47631), .Z(n47633) );
  AND U58638 ( .A(n47633), .B(n59846), .Z(n47634) );
  NANDN U58639 ( .A(x[7026]), .B(y[7026]), .Z(n59844) );
  AND U58640 ( .A(n47634), .B(n59844), .Z(n47638) );
  AND U58641 ( .A(n47636), .B(n47635), .Z(n47637) );
  NANDN U58642 ( .A(n47638), .B(n47637), .Z(n47639) );
  NAND U58643 ( .A(n47640), .B(n47639), .Z(n47641) );
  NAND U58644 ( .A(n47642), .B(n47641), .Z(n47643) );
  AND U58645 ( .A(n47643), .B(n59851), .Z(n47644) );
  NANDN U58646 ( .A(x[7030]), .B(y[7030]), .Z(n50878) );
  AND U58647 ( .A(n47644), .B(n50878), .Z(n47648) );
  AND U58648 ( .A(n47646), .B(n47645), .Z(n47647) );
  NANDN U58649 ( .A(n47648), .B(n47647), .Z(n47649) );
  NAND U58650 ( .A(n47650), .B(n47649), .Z(n47651) );
  NAND U58651 ( .A(n47652), .B(n47651), .Z(n47653) );
  AND U58652 ( .A(n47653), .B(n59854), .Z(n47654) );
  NANDN U58653 ( .A(x[7034]), .B(y[7034]), .Z(n50876) );
  AND U58654 ( .A(n47654), .B(n50876), .Z(n47658) );
  AND U58655 ( .A(n47656), .B(n47655), .Z(n47657) );
  NANDN U58656 ( .A(n47658), .B(n47657), .Z(n47659) );
  NAND U58657 ( .A(n47660), .B(n47659), .Z(n47661) );
  NAND U58658 ( .A(n47662), .B(n47661), .Z(n47664) );
  IV U58659 ( .A(n47663), .Z(n59860) );
  AND U58660 ( .A(n47664), .B(n59860), .Z(n47665) );
  NANDN U58661 ( .A(x[7038]), .B(y[7038]), .Z(n59858) );
  AND U58662 ( .A(n47665), .B(n59858), .Z(n47669) );
  AND U58663 ( .A(n47667), .B(n47666), .Z(n47668) );
  NANDN U58664 ( .A(n47669), .B(n47668), .Z(n47670) );
  NAND U58665 ( .A(n47671), .B(n47670), .Z(n47672) );
  NAND U58666 ( .A(n47673), .B(n47672), .Z(n47674) );
  AND U58667 ( .A(n47674), .B(n50873), .Z(n47676) );
  NANDN U58668 ( .A(x[7042]), .B(y[7042]), .Z(n47675) );
  AND U58669 ( .A(n47676), .B(n47675), .Z(n47680) );
  AND U58670 ( .A(n47678), .B(n47677), .Z(n47679) );
  NANDN U58671 ( .A(n47680), .B(n47679), .Z(n47681) );
  NAND U58672 ( .A(n47682), .B(n47681), .Z(n47683) );
  NAND U58673 ( .A(n47684), .B(n47683), .Z(n47685) );
  AND U58674 ( .A(n47685), .B(n59870), .Z(n47686) );
  NANDN U58675 ( .A(x[7046]), .B(y[7046]), .Z(n59868) );
  NAND U58676 ( .A(n47686), .B(n59868), .Z(n47687) );
  NAND U58677 ( .A(n47688), .B(n47687), .Z(n47689) );
  ANDN U58678 ( .B(y[7048]), .A(x[7048]), .Z(n59871) );
  ANDN U58679 ( .B(n47689), .A(n59871), .Z(n47690) );
  NANDN U58680 ( .A(n59872), .B(n47690), .Z(n47691) );
  NAND U58681 ( .A(n47692), .B(n47691), .Z(n47693) );
  AND U58682 ( .A(n47693), .B(n59875), .Z(n47694) );
  NANDN U58683 ( .A(x[7050]), .B(y[7050]), .Z(n59873) );
  AND U58684 ( .A(n47694), .B(n59873), .Z(n47698) );
  AND U58685 ( .A(n47696), .B(n47695), .Z(n47697) );
  NANDN U58686 ( .A(n47698), .B(n47697), .Z(n47699) );
  NAND U58687 ( .A(n47700), .B(n47699), .Z(n47701) );
  NAND U58688 ( .A(n47702), .B(n47701), .Z(n47703) );
  AND U58689 ( .A(n47703), .B(n59880), .Z(n47704) );
  NAND U58690 ( .A(n59878), .B(n47704), .Z(n47705) );
  NAND U58691 ( .A(n47706), .B(n47705), .Z(n47707) );
  NANDN U58692 ( .A(n47708), .B(n47707), .Z(n47709) );
  NANDN U58693 ( .A(x[7056]), .B(y[7056]), .Z(n59881) );
  NANDN U58694 ( .A(n47709), .B(n59881), .Z(n47710) );
  AND U58695 ( .A(n47711), .B(n47710), .Z(n47712) );
  OR U58696 ( .A(n47713), .B(n47712), .Z(n47714) );
  NAND U58697 ( .A(n47715), .B(n47714), .Z(n47716) );
  NANDN U58698 ( .A(n47717), .B(n47716), .Z(n47718) );
  NAND U58699 ( .A(n47719), .B(n47718), .Z(n47720) );
  AND U58700 ( .A(n47720), .B(n59889), .Z(n47721) );
  NANDN U58701 ( .A(x[7062]), .B(y[7062]), .Z(n50868) );
  AND U58702 ( .A(n47721), .B(n50868), .Z(n47725) );
  AND U58703 ( .A(n47723), .B(n47722), .Z(n47724) );
  NANDN U58704 ( .A(n47725), .B(n47724), .Z(n47726) );
  NAND U58705 ( .A(n47727), .B(n47726), .Z(n47728) );
  NAND U58706 ( .A(n47729), .B(n47728), .Z(n47730) );
  AND U58707 ( .A(n47730), .B(n59896), .Z(n47731) );
  NANDN U58708 ( .A(x[7066]), .B(y[7066]), .Z(n59894) );
  AND U58709 ( .A(n47731), .B(n59894), .Z(n47735) );
  AND U58710 ( .A(n47733), .B(n47732), .Z(n47734) );
  NANDN U58711 ( .A(n47735), .B(n47734), .Z(n47736) );
  NAND U58712 ( .A(n47737), .B(n47736), .Z(n47738) );
  NAND U58713 ( .A(n47739), .B(n47738), .Z(n47740) );
  AND U58714 ( .A(n47740), .B(n50865), .Z(n47741) );
  NANDN U58715 ( .A(x[7070]), .B(y[7070]), .Z(n59900) );
  AND U58716 ( .A(n47741), .B(n59900), .Z(n47745) );
  AND U58717 ( .A(n47743), .B(n47742), .Z(n47744) );
  NANDN U58718 ( .A(n47745), .B(n47744), .Z(n47746) );
  NAND U58719 ( .A(n47747), .B(n47746), .Z(n47748) );
  NAND U58720 ( .A(n47749), .B(n47748), .Z(n47750) );
  AND U58721 ( .A(n47750), .B(n50864), .Z(n47751) );
  NANDN U58722 ( .A(x[7074]), .B(y[7074]), .Z(n59904) );
  AND U58723 ( .A(n47751), .B(n59904), .Z(n47755) );
  AND U58724 ( .A(n47753), .B(n47752), .Z(n47754) );
  NANDN U58725 ( .A(n47755), .B(n47754), .Z(n47756) );
  NAND U58726 ( .A(n47757), .B(n47756), .Z(n47758) );
  AND U58727 ( .A(n47759), .B(n47758), .Z(n47761) );
  NANDN U58728 ( .A(x[7078]), .B(y[7078]), .Z(n59909) );
  AND U58729 ( .A(n59909), .B(n59911), .Z(n47760) );
  NANDN U58730 ( .A(n47761), .B(n47760), .Z(n47762) );
  NANDN U58731 ( .A(n47763), .B(n47762), .Z(n47764) );
  AND U58732 ( .A(n59913), .B(n47764), .Z(n47765) );
  NANDN U58733 ( .A(x[7080]), .B(y[7080]), .Z(n59912) );
  NAND U58734 ( .A(n47765), .B(n59912), .Z(n47766) );
  NAND U58735 ( .A(n47767), .B(n47766), .Z(n47768) );
  AND U58736 ( .A(n47768), .B(n50861), .Z(n47769) );
  NANDN U58737 ( .A(x[7082]), .B(y[7082]), .Z(n59914) );
  AND U58738 ( .A(n47769), .B(n59914), .Z(n47773) );
  AND U58739 ( .A(n47771), .B(n47770), .Z(n47772) );
  NANDN U58740 ( .A(n47773), .B(n47772), .Z(n47774) );
  NAND U58741 ( .A(n47775), .B(n47774), .Z(n47776) );
  NAND U58742 ( .A(n47777), .B(n47776), .Z(n47778) );
  AND U58743 ( .A(n47778), .B(n59920), .Z(n47779) );
  NANDN U58744 ( .A(x[7086]), .B(y[7086]), .Z(n59917) );
  AND U58745 ( .A(n47779), .B(n59917), .Z(n47783) );
  AND U58746 ( .A(n47781), .B(n47780), .Z(n47782) );
  NANDN U58747 ( .A(n47783), .B(n47782), .Z(n47784) );
  NAND U58748 ( .A(n47785), .B(n47784), .Z(n47786) );
  NAND U58749 ( .A(n47787), .B(n47786), .Z(n47788) );
  AND U58750 ( .A(n47788), .B(n59925), .Z(n47789) );
  NANDN U58751 ( .A(x[7090]), .B(y[7090]), .Z(n59924) );
  AND U58752 ( .A(n47789), .B(n59924), .Z(n47790) );
  OR U58753 ( .A(n47791), .B(n47790), .Z(n47792) );
  NAND U58754 ( .A(n47793), .B(n47792), .Z(n47794) );
  NAND U58755 ( .A(n47795), .B(n47794), .Z(n47796) );
  AND U58756 ( .A(n47797), .B(n47796), .Z(n47801) );
  AND U58757 ( .A(n47799), .B(n47798), .Z(n47800) );
  NANDN U58758 ( .A(n47801), .B(n47800), .Z(n47802) );
  NAND U58759 ( .A(n47803), .B(n47802), .Z(n47804) );
  NAND U58760 ( .A(n47805), .B(n47804), .Z(n47806) );
  AND U58761 ( .A(n47806), .B(n50855), .Z(n47807) );
  NANDN U58762 ( .A(x[7098]), .B(y[7098]), .Z(n59932) );
  AND U58763 ( .A(n47807), .B(n59932), .Z(n47811) );
  AND U58764 ( .A(n47809), .B(n47808), .Z(n47810) );
  NANDN U58765 ( .A(n47811), .B(n47810), .Z(n47812) );
  NAND U58766 ( .A(n47813), .B(n47812), .Z(n47814) );
  NAND U58767 ( .A(n47815), .B(n47814), .Z(n47816) );
  AND U58768 ( .A(n47816), .B(n59939), .Z(n47817) );
  NANDN U58769 ( .A(x[7102]), .B(y[7102]), .Z(n59937) );
  AND U58770 ( .A(n47817), .B(n59937), .Z(n47821) );
  AND U58771 ( .A(n47819), .B(n47818), .Z(n47820) );
  NANDN U58772 ( .A(n47821), .B(n47820), .Z(n47822) );
  NAND U58773 ( .A(n47823), .B(n47822), .Z(n47824) );
  NAND U58774 ( .A(n47825), .B(n47824), .Z(n47826) );
  AND U58775 ( .A(n47826), .B(n59944), .Z(n47827) );
  NANDN U58776 ( .A(x[7106]), .B(y[7106]), .Z(n59942) );
  AND U58777 ( .A(n47827), .B(n59942), .Z(n47831) );
  AND U58778 ( .A(n47829), .B(n47828), .Z(n47830) );
  NANDN U58779 ( .A(n47831), .B(n47830), .Z(n47832) );
  NAND U58780 ( .A(n47833), .B(n47832), .Z(n47834) );
  NAND U58781 ( .A(n47835), .B(n47834), .Z(n47836) );
  AND U58782 ( .A(n47836), .B(n59949), .Z(n47837) );
  NANDN U58783 ( .A(x[7110]), .B(y[7110]), .Z(n50850) );
  AND U58784 ( .A(n47837), .B(n50850), .Z(n47841) );
  AND U58785 ( .A(n47839), .B(n47838), .Z(n47840) );
  NANDN U58786 ( .A(n47841), .B(n47840), .Z(n47842) );
  NAND U58787 ( .A(n47843), .B(n47842), .Z(n47844) );
  NAND U58788 ( .A(n47845), .B(n47844), .Z(n47846) );
  AND U58789 ( .A(n47846), .B(n59954), .Z(n47847) );
  NANDN U58790 ( .A(x[7114]), .B(y[7114]), .Z(n59952) );
  AND U58791 ( .A(n47847), .B(n59952), .Z(n47851) );
  AND U58792 ( .A(n47849), .B(n47848), .Z(n47850) );
  NANDN U58793 ( .A(n47851), .B(n47850), .Z(n47852) );
  NAND U58794 ( .A(n47853), .B(n47852), .Z(n47854) );
  NAND U58795 ( .A(n47855), .B(n47854), .Z(n47856) );
  AND U58796 ( .A(n47856), .B(n59960), .Z(n47857) );
  NANDN U58797 ( .A(x[7118]), .B(y[7118]), .Z(n59958) );
  AND U58798 ( .A(n47857), .B(n59958), .Z(n47861) );
  AND U58799 ( .A(n47859), .B(n47858), .Z(n47860) );
  NANDN U58800 ( .A(n47861), .B(n47860), .Z(n47862) );
  NAND U58801 ( .A(n47863), .B(n47862), .Z(n47864) );
  NAND U58802 ( .A(n47865), .B(n47864), .Z(n47866) );
  AND U58803 ( .A(n47866), .B(n50844), .Z(n47867) );
  NANDN U58804 ( .A(x[7122]), .B(y[7122]), .Z(n59964) );
  NAND U58805 ( .A(n47867), .B(n59964), .Z(n47868) );
  NAND U58806 ( .A(n47869), .B(n47868), .Z(n47870) );
  ANDN U58807 ( .B(y[7124]), .A(x[7124]), .Z(n50845) );
  ANDN U58808 ( .B(n47870), .A(n50845), .Z(n47871) );
  NANDN U58809 ( .A(n59968), .B(n47871), .Z(n47872) );
  NAND U58810 ( .A(n47873), .B(n47872), .Z(n47875) );
  IV U58811 ( .A(n47874), .Z(n59972) );
  AND U58812 ( .A(n47875), .B(n59972), .Z(n47876) );
  NANDN U58813 ( .A(x[7126]), .B(y[7126]), .Z(n59969) );
  AND U58814 ( .A(n47876), .B(n59969), .Z(n47880) );
  AND U58815 ( .A(n47878), .B(n47877), .Z(n47879) );
  NANDN U58816 ( .A(n47880), .B(n47879), .Z(n47881) );
  NAND U58817 ( .A(n47882), .B(n47881), .Z(n47883) );
  NAND U58818 ( .A(n47884), .B(n47883), .Z(n47885) );
  AND U58819 ( .A(n47885), .B(n59976), .Z(n47886) );
  NANDN U58820 ( .A(x[7130]), .B(y[7130]), .Z(n59974) );
  AND U58821 ( .A(n47886), .B(n59974), .Z(n47890) );
  AND U58822 ( .A(n47888), .B(n47887), .Z(n47889) );
  NANDN U58823 ( .A(n47890), .B(n47889), .Z(n47891) );
  NAND U58824 ( .A(n47892), .B(n47891), .Z(n47893) );
  NAND U58825 ( .A(n47894), .B(n47893), .Z(n47895) );
  AND U58826 ( .A(n47895), .B(n59982), .Z(n47896) );
  NANDN U58827 ( .A(x[7134]), .B(y[7134]), .Z(n59979) );
  AND U58828 ( .A(n47896), .B(n59979), .Z(n47900) );
  AND U58829 ( .A(n47898), .B(n47897), .Z(n47899) );
  NANDN U58830 ( .A(n47900), .B(n47899), .Z(n47901) );
  NAND U58831 ( .A(n47902), .B(n47901), .Z(n47903) );
  NAND U58832 ( .A(n47904), .B(n47903), .Z(n47905) );
  AND U58833 ( .A(n47905), .B(n59987), .Z(n47906) );
  NANDN U58834 ( .A(x[7138]), .B(y[7138]), .Z(n59985) );
  AND U58835 ( .A(n47906), .B(n59985), .Z(n47910) );
  AND U58836 ( .A(n47908), .B(n47907), .Z(n47909) );
  NANDN U58837 ( .A(n47910), .B(n47909), .Z(n47911) );
  NAND U58838 ( .A(n47912), .B(n47911), .Z(n47913) );
  AND U58839 ( .A(n47914), .B(n47913), .Z(n47915) );
  OR U58840 ( .A(n47916), .B(n47915), .Z(n47917) );
  NAND U58841 ( .A(n47918), .B(n47917), .Z(n47919) );
  NANDN U58842 ( .A(n47920), .B(n47919), .Z(n47921) );
  NAND U58843 ( .A(n47922), .B(n47921), .Z(n47923) );
  AND U58844 ( .A(n47923), .B(n50835), .Z(n47924) );
  NANDN U58845 ( .A(x[7146]), .B(y[7146]), .Z(n50838) );
  AND U58846 ( .A(n47924), .B(n50838), .Z(n47928) );
  AND U58847 ( .A(n47926), .B(n47925), .Z(n47927) );
  NANDN U58848 ( .A(n47928), .B(n47927), .Z(n47929) );
  NAND U58849 ( .A(n47930), .B(n47929), .Z(n47931) );
  NAND U58850 ( .A(n47932), .B(n47931), .Z(n47933) );
  AND U58851 ( .A(n47933), .B(n50833), .Z(n47934) );
  NANDN U58852 ( .A(x[7150]), .B(y[7150]), .Z(n59996) );
  AND U58853 ( .A(n47934), .B(n59996), .Z(n47938) );
  AND U58854 ( .A(n47936), .B(n47935), .Z(n47937) );
  NANDN U58855 ( .A(n47938), .B(n47937), .Z(n47939) );
  NAND U58856 ( .A(n47940), .B(n47939), .Z(n47941) );
  AND U58857 ( .A(n47942), .B(n47941), .Z(n47944) );
  NANDN U58858 ( .A(x[7154]), .B(y[7154]), .Z(n60000) );
  AND U58859 ( .A(n60000), .B(n50830), .Z(n47943) );
  NANDN U58860 ( .A(n47944), .B(n47943), .Z(n47945) );
  NANDN U58861 ( .A(n47946), .B(n47945), .Z(n47947) );
  AND U58862 ( .A(n50827), .B(n47947), .Z(n47948) );
  NANDN U58863 ( .A(x[7156]), .B(y[7156]), .Z(n50831) );
  NAND U58864 ( .A(n47948), .B(n50831), .Z(n47949) );
  NAND U58865 ( .A(n47950), .B(n47949), .Z(n47952) );
  AND U58866 ( .A(n47952), .B(n47951), .Z(n47953) );
  NANDN U58867 ( .A(x[7158]), .B(y[7158]), .Z(n50828) );
  AND U58868 ( .A(n47953), .B(n50828), .Z(n47957) );
  AND U58869 ( .A(n47955), .B(n47954), .Z(n47956) );
  NANDN U58870 ( .A(n47957), .B(n47956), .Z(n47958) );
  NAND U58871 ( .A(n47959), .B(n47958), .Z(n47960) );
  NAND U58872 ( .A(n47961), .B(n47960), .Z(n47962) );
  AND U58873 ( .A(n47962), .B(n60008), .Z(n47963) );
  NANDN U58874 ( .A(x[7162]), .B(y[7162]), .Z(n60006) );
  AND U58875 ( .A(n47963), .B(n60006), .Z(n47967) );
  AND U58876 ( .A(n47965), .B(n47964), .Z(n47966) );
  NANDN U58877 ( .A(n47967), .B(n47966), .Z(n47968) );
  NAND U58878 ( .A(n47969), .B(n47968), .Z(n47970) );
  NAND U58879 ( .A(n47971), .B(n47970), .Z(n47972) );
  AND U58880 ( .A(n47972), .B(n60014), .Z(n47973) );
  NANDN U58881 ( .A(x[7166]), .B(y[7166]), .Z(n60012) );
  AND U58882 ( .A(n47973), .B(n60012), .Z(n47977) );
  AND U58883 ( .A(n47975), .B(n47974), .Z(n47976) );
  NANDN U58884 ( .A(n47977), .B(n47976), .Z(n47978) );
  NAND U58885 ( .A(n47979), .B(n47978), .Z(n47980) );
  NAND U58886 ( .A(n47981), .B(n47980), .Z(n47983) );
  AND U58887 ( .A(n47983), .B(n47982), .Z(n47984) );
  NANDN U58888 ( .A(x[7170]), .B(y[7170]), .Z(n60019) );
  AND U58889 ( .A(n47984), .B(n60019), .Z(n47988) );
  AND U58890 ( .A(n47986), .B(n47985), .Z(n47987) );
  NANDN U58891 ( .A(n47988), .B(n47987), .Z(n47989) );
  NAND U58892 ( .A(n47990), .B(n47989), .Z(n47991) );
  AND U58893 ( .A(n47992), .B(n47991), .Z(n47993) );
  ANDN U58894 ( .B(n50822), .A(n47993), .Z(n47994) );
  NAND U58895 ( .A(n60023), .B(n47994), .Z(n47995) );
  NANDN U58896 ( .A(n47996), .B(n47995), .Z(n47997) );
  OR U58897 ( .A(n47998), .B(n47997), .Z(n47999) );
  NAND U58898 ( .A(n48000), .B(n47999), .Z(n48001) );
  NAND U58899 ( .A(n48002), .B(n48001), .Z(n48003) );
  AND U58900 ( .A(n48003), .B(n60028), .Z(n48004) );
  NANDN U58901 ( .A(x[7178]), .B(y[7178]), .Z(n60026) );
  AND U58902 ( .A(n48004), .B(n60026), .Z(n48005) );
  OR U58903 ( .A(n48006), .B(n48005), .Z(n48007) );
  NAND U58904 ( .A(n48008), .B(n48007), .Z(n48009) );
  NAND U58905 ( .A(n48010), .B(n48009), .Z(n48011) );
  AND U58906 ( .A(n48011), .B(n60035), .Z(n48012) );
  NANDN U58907 ( .A(x[7182]), .B(y[7182]), .Z(n60033) );
  AND U58908 ( .A(n48012), .B(n60033), .Z(n48016) );
  AND U58909 ( .A(n48014), .B(n48013), .Z(n48015) );
  NANDN U58910 ( .A(n48016), .B(n48015), .Z(n48017) );
  NAND U58911 ( .A(n48018), .B(n48017), .Z(n48019) );
  NAND U58912 ( .A(n48020), .B(n48019), .Z(n48021) );
  AND U58913 ( .A(n48021), .B(n60039), .Z(n48022) );
  NANDN U58914 ( .A(x[7186]), .B(y[7186]), .Z(n50819) );
  AND U58915 ( .A(n48022), .B(n50819), .Z(n48026) );
  AND U58916 ( .A(n48024), .B(n48023), .Z(n48025) );
  NANDN U58917 ( .A(n48026), .B(n48025), .Z(n48027) );
  NAND U58918 ( .A(n48028), .B(n48027), .Z(n48029) );
  AND U58919 ( .A(n48030), .B(n48029), .Z(n48031) );
  OR U58920 ( .A(n48032), .B(n48031), .Z(n48033) );
  NAND U58921 ( .A(n48034), .B(n48033), .Z(n48035) );
  NANDN U58922 ( .A(n60046), .B(n48035), .Z(n48037) );
  NANDN U58923 ( .A(n48037), .B(n48036), .Z(n48038) );
  NAND U58924 ( .A(n48039), .B(n48038), .Z(n48040) );
  AND U58925 ( .A(n48040), .B(n50816), .Z(n48041) );
  NANDN U58926 ( .A(x[7194]), .B(y[7194]), .Z(n60047) );
  AND U58927 ( .A(n48041), .B(n60047), .Z(n48045) );
  AND U58928 ( .A(n48043), .B(n48042), .Z(n48044) );
  NANDN U58929 ( .A(n48045), .B(n48044), .Z(n48046) );
  NAND U58930 ( .A(n48047), .B(n48046), .Z(n48048) );
  NAND U58931 ( .A(n48049), .B(n48048), .Z(n48050) );
  AND U58932 ( .A(n48050), .B(n50815), .Z(n48051) );
  NANDN U58933 ( .A(x[7198]), .B(y[7198]), .Z(n60052) );
  AND U58934 ( .A(n48051), .B(n60052), .Z(n48055) );
  AND U58935 ( .A(n48053), .B(n48052), .Z(n48054) );
  NANDN U58936 ( .A(n48055), .B(n48054), .Z(n48056) );
  NAND U58937 ( .A(n48057), .B(n48056), .Z(n48058) );
  AND U58938 ( .A(n48059), .B(n48058), .Z(n48060) );
  OR U58939 ( .A(n48061), .B(n48060), .Z(n48062) );
  NAND U58940 ( .A(n48063), .B(n48062), .Z(n48064) );
  NANDN U58941 ( .A(n48065), .B(n48064), .Z(n48066) );
  NANDN U58942 ( .A(x[7204]), .B(y[7204]), .Z(n50812) );
  NANDN U58943 ( .A(n48066), .B(n50812), .Z(n48067) );
  AND U58944 ( .A(n48068), .B(n48067), .Z(n48069) );
  OR U58945 ( .A(n48070), .B(n48069), .Z(n48071) );
  NAND U58946 ( .A(n48072), .B(n48071), .Z(n48073) );
  NANDN U58947 ( .A(n48074), .B(n48073), .Z(n48075) );
  NANDN U58948 ( .A(n48075), .B(n60064), .Z(n48076) );
  NAND U58949 ( .A(n48077), .B(n48076), .Z(n48078) );
  AND U58950 ( .A(n48078), .B(n60066), .Z(n48079) );
  NANDN U58951 ( .A(x[7210]), .B(y[7210]), .Z(n60063) );
  AND U58952 ( .A(n48079), .B(n60063), .Z(n48083) );
  AND U58953 ( .A(n48081), .B(n48080), .Z(n48082) );
  NANDN U58954 ( .A(n48083), .B(n48082), .Z(n48084) );
  NAND U58955 ( .A(n48085), .B(n48084), .Z(n48086) );
  NAND U58956 ( .A(n48087), .B(n48086), .Z(n48088) );
  AND U58957 ( .A(n48088), .B(n60071), .Z(n48089) );
  NANDN U58958 ( .A(x[7214]), .B(y[7214]), .Z(n60070) );
  AND U58959 ( .A(n48089), .B(n60070), .Z(n48093) );
  AND U58960 ( .A(n48091), .B(n48090), .Z(n48092) );
  NANDN U58961 ( .A(n48093), .B(n48092), .Z(n48094) );
  NAND U58962 ( .A(n48095), .B(n48094), .Z(n48096) );
  NAND U58963 ( .A(n48097), .B(n48096), .Z(n48099) );
  AND U58964 ( .A(n48099), .B(n48098), .Z(n48100) );
  NANDN U58965 ( .A(x[7218]), .B(y[7218]), .Z(n60075) );
  AND U58966 ( .A(n48100), .B(n60075), .Z(n48104) );
  AND U58967 ( .A(n48102), .B(n48101), .Z(n48103) );
  NANDN U58968 ( .A(n48104), .B(n48103), .Z(n48105) );
  NAND U58969 ( .A(n48106), .B(n48105), .Z(n48107) );
  NAND U58970 ( .A(n48108), .B(n48107), .Z(n48109) );
  AND U58971 ( .A(n48109), .B(n50808), .Z(n48110) );
  NANDN U58972 ( .A(x[7222]), .B(y[7222]), .Z(n60080) );
  AND U58973 ( .A(n48110), .B(n60080), .Z(n48114) );
  AND U58974 ( .A(n48112), .B(n48111), .Z(n48113) );
  NANDN U58975 ( .A(n48114), .B(n48113), .Z(n48115) );
  NAND U58976 ( .A(n48116), .B(n48115), .Z(n48117) );
  NAND U58977 ( .A(n48118), .B(n48117), .Z(n48119) );
  AND U58978 ( .A(n48119), .B(n60085), .Z(n48120) );
  NANDN U58979 ( .A(x[7226]), .B(y[7226]), .Z(n60083) );
  AND U58980 ( .A(n48120), .B(n60083), .Z(n48124) );
  AND U58981 ( .A(n48122), .B(n48121), .Z(n48123) );
  NANDN U58982 ( .A(n48124), .B(n48123), .Z(n48125) );
  NAND U58983 ( .A(n48126), .B(n48125), .Z(n48127) );
  AND U58984 ( .A(n48128), .B(n48127), .Z(n48130) );
  NANDN U58985 ( .A(x[7230]), .B(y[7230]), .Z(n60088) );
  AND U58986 ( .A(n60088), .B(n60090), .Z(n48129) );
  NANDN U58987 ( .A(n48130), .B(n48129), .Z(n48131) );
  NAND U58988 ( .A(n48132), .B(n48131), .Z(n48133) );
  OR U58989 ( .A(n48134), .B(n48133), .Z(n48135) );
  NAND U58990 ( .A(n48136), .B(n48135), .Z(n48137) );
  NAND U58991 ( .A(n48138), .B(n48137), .Z(n48139) );
  AND U58992 ( .A(n48139), .B(n60094), .Z(n48140) );
  NANDN U58993 ( .A(x[7234]), .B(y[7234]), .Z(n50803) );
  AND U58994 ( .A(n48140), .B(n50803), .Z(n48141) );
  OR U58995 ( .A(n48142), .B(n48141), .Z(n48143) );
  NAND U58996 ( .A(n48144), .B(n48143), .Z(n48145) );
  NAND U58997 ( .A(n48146), .B(n48145), .Z(n48147) );
  AND U58998 ( .A(n48147), .B(n60098), .Z(n48148) );
  NANDN U58999 ( .A(x[7238]), .B(y[7238]), .Z(n50801) );
  AND U59000 ( .A(n48148), .B(n50801), .Z(n48152) );
  AND U59001 ( .A(n48150), .B(n48149), .Z(n48151) );
  NANDN U59002 ( .A(n48152), .B(n48151), .Z(n48153) );
  NAND U59003 ( .A(n48154), .B(n48153), .Z(n48155) );
  AND U59004 ( .A(n48156), .B(n48155), .Z(n48157) );
  OR U59005 ( .A(n48158), .B(n48157), .Z(n48159) );
  NAND U59006 ( .A(n48160), .B(n48159), .Z(n48161) );
  NANDN U59007 ( .A(n48162), .B(n48161), .Z(n48163) );
  NAND U59008 ( .A(n48164), .B(n48163), .Z(n48165) );
  AND U59009 ( .A(n48165), .B(n50799), .Z(n48167) );
  NANDN U59010 ( .A(x[7246]), .B(y[7246]), .Z(n48166) );
  AND U59011 ( .A(n48167), .B(n48166), .Z(n48171) );
  AND U59012 ( .A(n48169), .B(n48168), .Z(n48170) );
  NANDN U59013 ( .A(n48171), .B(n48170), .Z(n48172) );
  NAND U59014 ( .A(n48173), .B(n48172), .Z(n48174) );
  NAND U59015 ( .A(n48175), .B(n48174), .Z(n48177) );
  IV U59016 ( .A(n48176), .Z(n50795) );
  AND U59017 ( .A(n48177), .B(n50795), .Z(n48178) );
  NANDN U59018 ( .A(x[7250]), .B(y[7250]), .Z(n60112) );
  AND U59019 ( .A(n48178), .B(n60112), .Z(n48182) );
  AND U59020 ( .A(n48180), .B(n48179), .Z(n48181) );
  NANDN U59021 ( .A(n48182), .B(n48181), .Z(n48183) );
  NAND U59022 ( .A(n48184), .B(n48183), .Z(n48185) );
  NAND U59023 ( .A(n48186), .B(n48185), .Z(n48187) );
  AND U59024 ( .A(n48187), .B(n60120), .Z(n48188) );
  NANDN U59025 ( .A(x[7254]), .B(y[7254]), .Z(n60117) );
  AND U59026 ( .A(n48188), .B(n60117), .Z(n48192) );
  AND U59027 ( .A(n48190), .B(n48189), .Z(n48191) );
  NANDN U59028 ( .A(n48192), .B(n48191), .Z(n48193) );
  NAND U59029 ( .A(n48194), .B(n48193), .Z(n48195) );
  NAND U59030 ( .A(n48196), .B(n48195), .Z(n48197) );
  AND U59031 ( .A(n48197), .B(n60125), .Z(n48198) );
  NANDN U59032 ( .A(x[7258]), .B(y[7258]), .Z(n60123) );
  AND U59033 ( .A(n48198), .B(n60123), .Z(n48202) );
  AND U59034 ( .A(n48200), .B(n48199), .Z(n48201) );
  NANDN U59035 ( .A(n48202), .B(n48201), .Z(n48203) );
  NAND U59036 ( .A(n48204), .B(n48203), .Z(n48205) );
  NAND U59037 ( .A(n48206), .B(n48205), .Z(n48207) );
  AND U59038 ( .A(n48207), .B(n60130), .Z(n48208) );
  NANDN U59039 ( .A(n48209), .B(n48208), .Z(n48210) );
  NAND U59040 ( .A(n48211), .B(n48210), .Z(n48212) );
  NANDN U59041 ( .A(n50794), .B(n48212), .Z(n48213) );
  NANDN U59042 ( .A(x[7264]), .B(y[7264]), .Z(n60131) );
  NANDN U59043 ( .A(n48213), .B(n60131), .Z(n48214) );
  NAND U59044 ( .A(n48215), .B(n48214), .Z(n48216) );
  AND U59045 ( .A(n48216), .B(n50791), .Z(n48217) );
  NANDN U59046 ( .A(x[7266]), .B(y[7266]), .Z(n50793) );
  AND U59047 ( .A(n48217), .B(n50793), .Z(n48221) );
  AND U59048 ( .A(n48219), .B(n48218), .Z(n48220) );
  NANDN U59049 ( .A(n48221), .B(n48220), .Z(n48222) );
  NAND U59050 ( .A(n48223), .B(n48222), .Z(n48224) );
  NAND U59051 ( .A(n48225), .B(n48224), .Z(n48226) );
  AND U59052 ( .A(n48226), .B(n50790), .Z(n48227) );
  NANDN U59053 ( .A(x[7270]), .B(y[7270]), .Z(n60138) );
  AND U59054 ( .A(n48227), .B(n60138), .Z(n48231) );
  AND U59055 ( .A(n48229), .B(n48228), .Z(n48230) );
  NANDN U59056 ( .A(n48231), .B(n48230), .Z(n48232) );
  NAND U59057 ( .A(n48233), .B(n48232), .Z(n48234) );
  NAND U59058 ( .A(n48235), .B(n48234), .Z(n48236) );
  AND U59059 ( .A(n48236), .B(n60144), .Z(n48237) );
  NANDN U59060 ( .A(x[7274]), .B(y[7274]), .Z(n60142) );
  AND U59061 ( .A(n48237), .B(n60142), .Z(n48241) );
  AND U59062 ( .A(n48239), .B(n48238), .Z(n48240) );
  NANDN U59063 ( .A(n48241), .B(n48240), .Z(n48242) );
  NAND U59064 ( .A(n48243), .B(n48242), .Z(n48244) );
  NAND U59065 ( .A(n48245), .B(n48244), .Z(n48246) );
  AND U59066 ( .A(n48246), .B(n60150), .Z(n48247) );
  NANDN U59067 ( .A(x[7278]), .B(y[7278]), .Z(n60148) );
  AND U59068 ( .A(n48247), .B(n60148), .Z(n48251) );
  AND U59069 ( .A(n48249), .B(n48248), .Z(n48250) );
  NANDN U59070 ( .A(n48251), .B(n48250), .Z(n48252) );
  NAND U59071 ( .A(n48253), .B(n48252), .Z(n48254) );
  AND U59072 ( .A(n48255), .B(n48254), .Z(n48258) );
  NANDN U59073 ( .A(x[7282]), .B(y[7282]), .Z(n50787) );
  IV U59074 ( .A(n48256), .Z(n60154) );
  AND U59075 ( .A(n50787), .B(n60154), .Z(n48257) );
  NANDN U59076 ( .A(n48258), .B(n48257), .Z(n48259) );
  NANDN U59077 ( .A(n48260), .B(n48259), .Z(n48261) );
  AND U59078 ( .A(n48262), .B(n48261), .Z(n48263) );
  OR U59079 ( .A(n48264), .B(n48263), .Z(n48265) );
  NAND U59080 ( .A(n48266), .B(n48265), .Z(n48267) );
  NANDN U59081 ( .A(n48268), .B(n48267), .Z(n48269) );
  NAND U59082 ( .A(n48270), .B(n48269), .Z(n48271) );
  NAND U59083 ( .A(n48272), .B(n48271), .Z(n48273) );
  AND U59084 ( .A(n48273), .B(n50784), .Z(n48274) );
  NANDN U59085 ( .A(x[7290]), .B(y[7290]), .Z(n60162) );
  AND U59086 ( .A(n48274), .B(n60162), .Z(n48278) );
  AND U59087 ( .A(n48276), .B(n48275), .Z(n48277) );
  NANDN U59088 ( .A(n48278), .B(n48277), .Z(n48279) );
  NAND U59089 ( .A(n48280), .B(n48279), .Z(n48281) );
  AND U59090 ( .A(n48282), .B(n48281), .Z(n48283) );
  OR U59091 ( .A(n48284), .B(n48283), .Z(n48285) );
  NAND U59092 ( .A(n48286), .B(n48285), .Z(n48287) );
  NANDN U59093 ( .A(n48288), .B(n48287), .Z(n48289) );
  NAND U59094 ( .A(n48290), .B(n48289), .Z(n48291) );
  AND U59095 ( .A(n48292), .B(n48291), .Z(n48296) );
  AND U59096 ( .A(n48294), .B(n48293), .Z(n48295) );
  NANDN U59097 ( .A(n48296), .B(n48295), .Z(n48297) );
  NAND U59098 ( .A(n48298), .B(n48297), .Z(n48299) );
  NAND U59099 ( .A(n48300), .B(n48299), .Z(n48301) );
  AND U59100 ( .A(n48301), .B(n60174), .Z(n48302) );
  NANDN U59101 ( .A(x[7302]), .B(y[7302]), .Z(n50778) );
  AND U59102 ( .A(n48302), .B(n50778), .Z(n48306) );
  AND U59103 ( .A(n48304), .B(n48303), .Z(n48305) );
  NANDN U59104 ( .A(n48306), .B(n48305), .Z(n48307) );
  NAND U59105 ( .A(n48308), .B(n48307), .Z(n48309) );
  AND U59106 ( .A(n48310), .B(n48309), .Z(n48311) );
  ANDN U59107 ( .B(n60178), .A(n48311), .Z(n48312) );
  NANDN U59108 ( .A(x[7306]), .B(y[7306]), .Z(n50777) );
  AND U59109 ( .A(n48312), .B(n50777), .Z(n48316) );
  NAND U59110 ( .A(n48314), .B(n48313), .Z(n48315) );
  OR U59111 ( .A(n48316), .B(n48315), .Z(n48317) );
  AND U59112 ( .A(n48318), .B(n48317), .Z(n48319) );
  OR U59113 ( .A(n48320), .B(n48319), .Z(n48321) );
  NAND U59114 ( .A(n48322), .B(n48321), .Z(n48323) );
  NANDN U59115 ( .A(n48324), .B(n48323), .Z(n48325) );
  OR U59116 ( .A(n48326), .B(n48325), .Z(n48327) );
  NAND U59117 ( .A(n48328), .B(n48327), .Z(n48329) );
  NAND U59118 ( .A(n48330), .B(n48329), .Z(n48331) );
  AND U59119 ( .A(n48331), .B(n50774), .Z(n48332) );
  NANDN U59120 ( .A(x[7314]), .B(y[7314]), .Z(n60188) );
  AND U59121 ( .A(n48332), .B(n60188), .Z(n48333) );
  OR U59122 ( .A(n48334), .B(n48333), .Z(n48335) );
  NAND U59123 ( .A(n48336), .B(n48335), .Z(n48337) );
  NAND U59124 ( .A(n48338), .B(n48337), .Z(n48339) );
  AND U59125 ( .A(n48339), .B(n50773), .Z(n48340) );
  NANDN U59126 ( .A(x[7318]), .B(y[7318]), .Z(n60193) );
  AND U59127 ( .A(n48340), .B(n60193), .Z(n48344) );
  AND U59128 ( .A(n48342), .B(n48341), .Z(n48343) );
  NANDN U59129 ( .A(n48344), .B(n48343), .Z(n48345) );
  NAND U59130 ( .A(n48346), .B(n48345), .Z(n48347) );
  NAND U59131 ( .A(n48348), .B(n48347), .Z(n48349) );
  AND U59132 ( .A(n48349), .B(n60199), .Z(n48350) );
  NANDN U59133 ( .A(x[7322]), .B(y[7322]), .Z(n60197) );
  AND U59134 ( .A(n48350), .B(n60197), .Z(n48354) );
  AND U59135 ( .A(n48352), .B(n48351), .Z(n48353) );
  NANDN U59136 ( .A(n48354), .B(n48353), .Z(n48355) );
  NAND U59137 ( .A(n48356), .B(n48355), .Z(n48357) );
  NAND U59138 ( .A(n48358), .B(n48357), .Z(n48359) );
  AND U59139 ( .A(n48359), .B(n60205), .Z(n48360) );
  NANDN U59140 ( .A(x[7326]), .B(y[7326]), .Z(n60203) );
  AND U59141 ( .A(n48360), .B(n60203), .Z(n48364) );
  AND U59142 ( .A(n48362), .B(n48361), .Z(n48363) );
  NANDN U59143 ( .A(n48364), .B(n48363), .Z(n48365) );
  NAND U59144 ( .A(n48366), .B(n48365), .Z(n48367) );
  NAND U59145 ( .A(n48368), .B(n48367), .Z(n48369) );
  AND U59146 ( .A(n48369), .B(n60209), .Z(n48370) );
  NANDN U59147 ( .A(x[7330]), .B(y[7330]), .Z(n50770) );
  AND U59148 ( .A(n48370), .B(n50770), .Z(n48374) );
  AND U59149 ( .A(n48372), .B(n48371), .Z(n48373) );
  NANDN U59150 ( .A(n48374), .B(n48373), .Z(n48375) );
  NAND U59151 ( .A(n48376), .B(n48375), .Z(n48377) );
  NAND U59152 ( .A(n48378), .B(n48377), .Z(n48380) );
  IV U59153 ( .A(n48379), .Z(n60212) );
  AND U59154 ( .A(n48380), .B(n60212), .Z(n48381) );
  NANDN U59155 ( .A(x[7334]), .B(y[7334]), .Z(n50768) );
  AND U59156 ( .A(n48381), .B(n50768), .Z(n48385) );
  AND U59157 ( .A(n48383), .B(n48382), .Z(n48384) );
  NANDN U59158 ( .A(n48385), .B(n48384), .Z(n48386) );
  NAND U59159 ( .A(n48387), .B(n48386), .Z(n48388) );
  AND U59160 ( .A(n48389), .B(n48388), .Z(n48390) );
  ANDN U59161 ( .B(n60219), .A(n48390), .Z(n48391) );
  NAND U59162 ( .A(n60217), .B(n48391), .Z(n48392) );
  NANDN U59163 ( .A(n48393), .B(n48392), .Z(n48394) );
  AND U59164 ( .A(n48394), .B(n60222), .Z(n48395) );
  NANDN U59165 ( .A(x[7340]), .B(y[7340]), .Z(n60220) );
  NAND U59166 ( .A(n48395), .B(n60220), .Z(n48396) );
  NAND U59167 ( .A(n48397), .B(n48396), .Z(n48398) );
  AND U59168 ( .A(n48398), .B(n50764), .Z(n48399) );
  NANDN U59169 ( .A(x[7342]), .B(y[7342]), .Z(n60223) );
  AND U59170 ( .A(n48399), .B(n60223), .Z(n48403) );
  AND U59171 ( .A(n48401), .B(n48400), .Z(n48402) );
  NANDN U59172 ( .A(n48403), .B(n48402), .Z(n48404) );
  NAND U59173 ( .A(n48405), .B(n48404), .Z(n48406) );
  AND U59174 ( .A(n48407), .B(n48406), .Z(n48408) );
  OR U59175 ( .A(n48409), .B(n48408), .Z(n48410) );
  NAND U59176 ( .A(n48411), .B(n48410), .Z(n48412) );
  NANDN U59177 ( .A(n48413), .B(n48412), .Z(n48414) );
  NAND U59178 ( .A(n48415), .B(n48414), .Z(n48416) );
  AND U59179 ( .A(n48416), .B(n60233), .Z(n48417) );
  NANDN U59180 ( .A(x[7350]), .B(y[7350]), .Z(n60231) );
  AND U59181 ( .A(n48417), .B(n60231), .Z(n48421) );
  AND U59182 ( .A(n48419), .B(n48418), .Z(n48420) );
  NANDN U59183 ( .A(n48421), .B(n48420), .Z(n48422) );
  NAND U59184 ( .A(n48423), .B(n48422), .Z(n48424) );
  NAND U59185 ( .A(n48425), .B(n48424), .Z(n48426) );
  AND U59186 ( .A(n48426), .B(n60237), .Z(n48427) );
  NANDN U59187 ( .A(x[7354]), .B(y[7354]), .Z(n50760) );
  AND U59188 ( .A(n48427), .B(n50760), .Z(n48431) );
  AND U59189 ( .A(n48429), .B(n48428), .Z(n48430) );
  NANDN U59190 ( .A(n48431), .B(n48430), .Z(n48432) );
  NAND U59191 ( .A(n48433), .B(n48432), .Z(n48434) );
  AND U59192 ( .A(n48435), .B(n48434), .Z(n48436) );
  ANDN U59193 ( .B(n48437), .A(n48436), .Z(n48438) );
  OR U59194 ( .A(n48439), .B(n48438), .Z(n48440) );
  NAND U59195 ( .A(n48441), .B(n48440), .Z(n48442) );
  NAND U59196 ( .A(n48443), .B(n48442), .Z(n48445) );
  AND U59197 ( .A(n48445), .B(n48444), .Z(n48446) );
  NANDN U59198 ( .A(x[7362]), .B(y[7362]), .Z(n60248) );
  AND U59199 ( .A(n48446), .B(n60248), .Z(n48450) );
  AND U59200 ( .A(n48448), .B(n48447), .Z(n48449) );
  NANDN U59201 ( .A(n48450), .B(n48449), .Z(n48451) );
  NAND U59202 ( .A(n48452), .B(n48451), .Z(n48453) );
  NAND U59203 ( .A(n48454), .B(n48453), .Z(n48455) );
  AND U59204 ( .A(n48455), .B(n50758), .Z(n48456) );
  NANDN U59205 ( .A(x[7366]), .B(y[7366]), .Z(n60252) );
  AND U59206 ( .A(n48456), .B(n60252), .Z(n48460) );
  AND U59207 ( .A(n48458), .B(n48457), .Z(n48459) );
  NANDN U59208 ( .A(n48460), .B(n48459), .Z(n48461) );
  NAND U59209 ( .A(n48462), .B(n48461), .Z(n48463) );
  NAND U59210 ( .A(n48464), .B(n48463), .Z(n48466) );
  IV U59211 ( .A(n48465), .Z(n50755) );
  AND U59212 ( .A(n48466), .B(n50755), .Z(n48467) );
  NANDN U59213 ( .A(x[7370]), .B(y[7370]), .Z(n60256) );
  AND U59214 ( .A(n48467), .B(n60256), .Z(n48471) );
  AND U59215 ( .A(n48469), .B(n48468), .Z(n48470) );
  NANDN U59216 ( .A(n48471), .B(n48470), .Z(n48472) );
  NAND U59217 ( .A(n48473), .B(n48472), .Z(n48474) );
  NAND U59218 ( .A(n48475), .B(n48474), .Z(n48476) );
  AND U59219 ( .A(n48476), .B(n50751), .Z(n48477) );
  NANDN U59220 ( .A(x[7374]), .B(y[7374]), .Z(n50754) );
  AND U59221 ( .A(n48477), .B(n50754), .Z(n48481) );
  AND U59222 ( .A(n48479), .B(n48478), .Z(n48480) );
  NANDN U59223 ( .A(n48481), .B(n48480), .Z(n48482) );
  NAND U59224 ( .A(n48483), .B(n48482), .Z(n48484) );
  AND U59225 ( .A(n48485), .B(n48484), .Z(n48486) );
  OR U59226 ( .A(n48487), .B(n48486), .Z(n48488) );
  NAND U59227 ( .A(n48489), .B(n48488), .Z(n48490) );
  NANDN U59228 ( .A(n48491), .B(n48490), .Z(n48492) );
  NAND U59229 ( .A(n48493), .B(n48492), .Z(n48494) );
  AND U59230 ( .A(n48495), .B(n48494), .Z(n48499) );
  AND U59231 ( .A(n48497), .B(n48496), .Z(n48498) );
  NANDN U59232 ( .A(n48499), .B(n48498), .Z(n48500) );
  NAND U59233 ( .A(n48501), .B(n48500), .Z(n48502) );
  NAND U59234 ( .A(n48503), .B(n48502), .Z(n48504) );
  AND U59235 ( .A(n48504), .B(n50747), .Z(n48505) );
  NANDN U59236 ( .A(x[7386]), .B(y[7386]), .Z(n60273) );
  AND U59237 ( .A(n48505), .B(n60273), .Z(n48509) );
  AND U59238 ( .A(n48507), .B(n48506), .Z(n48508) );
  NANDN U59239 ( .A(n48509), .B(n48508), .Z(n48510) );
  NAND U59240 ( .A(n48511), .B(n48510), .Z(n48512) );
  NAND U59241 ( .A(n48513), .B(n48512), .Z(n48515) );
  AND U59242 ( .A(n48515), .B(n48514), .Z(n48516) );
  NAND U59243 ( .A(n60276), .B(n48516), .Z(n48517) );
  NAND U59244 ( .A(n48518), .B(n48517), .Z(n48519) );
  NANDN U59245 ( .A(n48520), .B(n48519), .Z(n48521) );
  AND U59246 ( .A(n48522), .B(n48521), .Z(n48523) );
  OR U59247 ( .A(n48524), .B(n48523), .Z(n48525) );
  NAND U59248 ( .A(n48526), .B(n48525), .Z(n48527) );
  NANDN U59249 ( .A(n48528), .B(n48527), .Z(n48529) );
  NAND U59250 ( .A(n48530), .B(n48529), .Z(n48531) );
  AND U59251 ( .A(n48531), .B(n60286), .Z(n48532) );
  NANDN U59252 ( .A(x[7398]), .B(y[7398]), .Z(n60284) );
  AND U59253 ( .A(n48532), .B(n60284), .Z(n48536) );
  AND U59254 ( .A(n48534), .B(n48533), .Z(n48535) );
  NANDN U59255 ( .A(n48536), .B(n48535), .Z(n48537) );
  NAND U59256 ( .A(n48538), .B(n48537), .Z(n48539) );
  NAND U59257 ( .A(n48540), .B(n48539), .Z(n48541) );
  AND U59258 ( .A(n48541), .B(n60293), .Z(n48542) );
  NANDN U59259 ( .A(x[7402]), .B(y[7402]), .Z(n60290) );
  AND U59260 ( .A(n48542), .B(n60290), .Z(n48546) );
  AND U59261 ( .A(n48544), .B(n48543), .Z(n48545) );
  NANDN U59262 ( .A(n48546), .B(n48545), .Z(n48547) );
  NAND U59263 ( .A(n48548), .B(n48547), .Z(n48549) );
  NAND U59264 ( .A(n48550), .B(n48549), .Z(n48551) );
  AND U59265 ( .A(n48551), .B(n50741), .Z(n48552) );
  NANDN U59266 ( .A(x[7406]), .B(y[7406]), .Z(n60298) );
  AND U59267 ( .A(n48552), .B(n60298), .Z(n48556) );
  AND U59268 ( .A(n48554), .B(n48553), .Z(n48555) );
  NANDN U59269 ( .A(n48556), .B(n48555), .Z(n48557) );
  NAND U59270 ( .A(n48558), .B(n48557), .Z(n48559) );
  NAND U59271 ( .A(n48560), .B(n48559), .Z(n48561) );
  AND U59272 ( .A(n48561), .B(n60304), .Z(n48562) );
  NANDN U59273 ( .A(x[7410]), .B(y[7410]), .Z(n60302) );
  AND U59274 ( .A(n48562), .B(n60302), .Z(n48566) );
  AND U59275 ( .A(n48564), .B(n48563), .Z(n48565) );
  NANDN U59276 ( .A(n48566), .B(n48565), .Z(n48567) );
  NAND U59277 ( .A(n48568), .B(n48567), .Z(n48569) );
  AND U59278 ( .A(n48570), .B(n48569), .Z(n48572) );
  NANDN U59279 ( .A(x[7414]), .B(y[7414]), .Z(n60308) );
  AND U59280 ( .A(n60308), .B(n60311), .Z(n48571) );
  NANDN U59281 ( .A(n48572), .B(n48571), .Z(n48573) );
  NAND U59282 ( .A(n48574), .B(n48573), .Z(n48575) );
  OR U59283 ( .A(n48576), .B(n48575), .Z(n48577) );
  NAND U59284 ( .A(n48578), .B(n48577), .Z(n48579) );
  NAND U59285 ( .A(n48580), .B(n48579), .Z(n48581) );
  AND U59286 ( .A(n48581), .B(n50738), .Z(n48582) );
  NANDN U59287 ( .A(x[7418]), .B(y[7418]), .Z(n60314) );
  AND U59288 ( .A(n48582), .B(n60314), .Z(n48586) );
  AND U59289 ( .A(n48584), .B(n48583), .Z(n48585) );
  NANDN U59290 ( .A(n48586), .B(n48585), .Z(n48587) );
  NAND U59291 ( .A(n48588), .B(n48587), .Z(n48589) );
  AND U59292 ( .A(n48590), .B(n48589), .Z(n48591) );
  OR U59293 ( .A(n48592), .B(n48591), .Z(n48593) );
  NAND U59294 ( .A(n48594), .B(n48593), .Z(n48595) );
  NANDN U59295 ( .A(n48596), .B(n48595), .Z(n48597) );
  NAND U59296 ( .A(n48598), .B(n48597), .Z(n48600) );
  IV U59297 ( .A(n48599), .Z(n50733) );
  AND U59298 ( .A(n48600), .B(n50733), .Z(n48601) );
  NANDN U59299 ( .A(x[7426]), .B(y[7426]), .Z(n50735) );
  AND U59300 ( .A(n48601), .B(n50735), .Z(n48602) );
  OR U59301 ( .A(n48603), .B(n48602), .Z(n48604) );
  NAND U59302 ( .A(n48605), .B(n48604), .Z(n48606) );
  NAND U59303 ( .A(n48607), .B(n48606), .Z(n48608) );
  AND U59304 ( .A(n48608), .B(n50731), .Z(n48609) );
  NANDN U59305 ( .A(x[7430]), .B(y[7430]), .Z(n60327) );
  AND U59306 ( .A(n48609), .B(n60327), .Z(n48613) );
  AND U59307 ( .A(n48611), .B(n48610), .Z(n48612) );
  NANDN U59308 ( .A(n48613), .B(n48612), .Z(n48614) );
  NAND U59309 ( .A(n48615), .B(n48614), .Z(n48616) );
  AND U59310 ( .A(n48617), .B(n48616), .Z(n48618) );
  ANDN U59311 ( .B(n60333), .A(n48618), .Z(n48619) );
  NANDN U59312 ( .A(x[7434]), .B(y[7434]), .Z(n60331) );
  AND U59313 ( .A(n48619), .B(n60331), .Z(n48620) );
  OR U59314 ( .A(n48621), .B(n48620), .Z(n48622) );
  NAND U59315 ( .A(n48623), .B(n48622), .Z(n48624) );
  NAND U59316 ( .A(n48625), .B(n48624), .Z(n48626) );
  AND U59317 ( .A(n48626), .B(n60340), .Z(n48627) );
  NANDN U59318 ( .A(x[7438]), .B(y[7438]), .Z(n60337) );
  AND U59319 ( .A(n48627), .B(n60337), .Z(n48631) );
  AND U59320 ( .A(n48629), .B(n48628), .Z(n48630) );
  NANDN U59321 ( .A(n48631), .B(n48630), .Z(n48632) );
  NAND U59322 ( .A(n48633), .B(n48632), .Z(n48634) );
  NAND U59323 ( .A(n48635), .B(n48634), .Z(n48636) );
  AND U59324 ( .A(n48636), .B(n60344), .Z(n48637) );
  NANDN U59325 ( .A(x[7442]), .B(y[7442]), .Z(n50728) );
  AND U59326 ( .A(n48637), .B(n50728), .Z(n48641) );
  AND U59327 ( .A(n48639), .B(n48638), .Z(n48640) );
  NANDN U59328 ( .A(n48641), .B(n48640), .Z(n48642) );
  NAND U59329 ( .A(n48643), .B(n48642), .Z(n48644) );
  NAND U59330 ( .A(n48645), .B(n48644), .Z(n48647) );
  IV U59331 ( .A(n48646), .Z(n60347) );
  AND U59332 ( .A(n48647), .B(n60347), .Z(n48648) );
  NANDN U59333 ( .A(x[7446]), .B(y[7446]), .Z(n50727) );
  AND U59334 ( .A(n48648), .B(n50727), .Z(n48652) );
  AND U59335 ( .A(n48650), .B(n48649), .Z(n48651) );
  NANDN U59336 ( .A(n48652), .B(n48651), .Z(n48653) );
  NAND U59337 ( .A(n48654), .B(n48653), .Z(n48655) );
  NAND U59338 ( .A(n48656), .B(n48655), .Z(n48657) );
  AND U59339 ( .A(n48657), .B(n60353), .Z(n48659) );
  NANDN U59340 ( .A(x[7450]), .B(y[7450]), .Z(n48658) );
  AND U59341 ( .A(n48659), .B(n48658), .Z(n48663) );
  AND U59342 ( .A(n48661), .B(n48660), .Z(n48662) );
  NANDN U59343 ( .A(n48663), .B(n48662), .Z(n48664) );
  NAND U59344 ( .A(n48665), .B(n48664), .Z(n48666) );
  NAND U59345 ( .A(n48667), .B(n48666), .Z(n48668) );
  AND U59346 ( .A(n48668), .B(n60360), .Z(n48669) );
  NANDN U59347 ( .A(x[7454]), .B(y[7454]), .Z(n60357) );
  AND U59348 ( .A(n48669), .B(n60357), .Z(n48673) );
  AND U59349 ( .A(n48671), .B(n48670), .Z(n48672) );
  NANDN U59350 ( .A(n48673), .B(n48672), .Z(n48674) );
  NAND U59351 ( .A(n48675), .B(n48674), .Z(n48676) );
  NAND U59352 ( .A(n48677), .B(n48676), .Z(n48678) );
  AND U59353 ( .A(n48678), .B(n60365), .Z(n48679) );
  NANDN U59354 ( .A(x[7458]), .B(y[7458]), .Z(n60363) );
  AND U59355 ( .A(n48679), .B(n60363), .Z(n48683) );
  AND U59356 ( .A(n48681), .B(n48680), .Z(n48682) );
  NANDN U59357 ( .A(n48683), .B(n48682), .Z(n48684) );
  NAND U59358 ( .A(n48685), .B(n48684), .Z(n48686) );
  AND U59359 ( .A(n48687), .B(n48686), .Z(n48688) );
  ANDN U59360 ( .B(n48689), .A(n48688), .Z(n48690) );
  OR U59361 ( .A(n48691), .B(n48690), .Z(n48692) );
  NAND U59362 ( .A(n48693), .B(n48692), .Z(n48694) );
  AND U59363 ( .A(n48695), .B(n48694), .Z(n48696) );
  NOR U59364 ( .A(n48697), .B(n48696), .Z(n48698) );
  NAND U59365 ( .A(n48699), .B(n48698), .Z(n48700) );
  NANDN U59366 ( .A(n48701), .B(n48700), .Z(n48702) );
  OR U59367 ( .A(n48703), .B(n48702), .Z(n48704) );
  NAND U59368 ( .A(n48705), .B(n48704), .Z(n48706) );
  NAND U59369 ( .A(n48707), .B(n48706), .Z(n48709) );
  AND U59370 ( .A(n48709), .B(n48708), .Z(n48710) );
  NANDN U59371 ( .A(x[7470]), .B(y[7470]), .Z(n60378) );
  AND U59372 ( .A(n48710), .B(n60378), .Z(n48714) );
  AND U59373 ( .A(n48712), .B(n48711), .Z(n48713) );
  NANDN U59374 ( .A(n48714), .B(n48713), .Z(n48715) );
  NAND U59375 ( .A(n48716), .B(n48715), .Z(n48717) );
  NAND U59376 ( .A(n48718), .B(n48717), .Z(n48719) );
  AND U59377 ( .A(n48719), .B(n50719), .Z(n48720) );
  NANDN U59378 ( .A(x[7474]), .B(y[7474]), .Z(n60382) );
  AND U59379 ( .A(n48720), .B(n60382), .Z(n48724) );
  AND U59380 ( .A(n48722), .B(n48721), .Z(n48723) );
  NANDN U59381 ( .A(n48724), .B(n48723), .Z(n48725) );
  NAND U59382 ( .A(n48726), .B(n48725), .Z(n48727) );
  AND U59383 ( .A(n48728), .B(n48727), .Z(n48729) );
  OR U59384 ( .A(n48730), .B(n48729), .Z(n48731) );
  NAND U59385 ( .A(n48732), .B(n48731), .Z(n48733) );
  NAND U59386 ( .A(n50713), .B(n48733), .Z(n48734) );
  NANDN U59387 ( .A(x[7480]), .B(y[7480]), .Z(n50716) );
  NANDN U59388 ( .A(n48734), .B(n50716), .Z(n48735) );
  NAND U59389 ( .A(n48736), .B(n48735), .Z(n48738) );
  AND U59390 ( .A(n48738), .B(n48737), .Z(n48739) );
  NANDN U59391 ( .A(n50712), .B(n48739), .Z(n48740) );
  NAND U59392 ( .A(n48741), .B(n48740), .Z(n48742) );
  NANDN U59393 ( .A(n48743), .B(n48742), .Z(n48744) );
  AND U59394 ( .A(n48745), .B(n48744), .Z(n48746) );
  OR U59395 ( .A(n48747), .B(n48746), .Z(n48748) );
  NAND U59396 ( .A(n48749), .B(n48748), .Z(n48750) );
  NANDN U59397 ( .A(n48751), .B(n48750), .Z(n48753) );
  NANDN U59398 ( .A(n48753), .B(n48752), .Z(n48754) );
  AND U59399 ( .A(n48755), .B(n48754), .Z(n48756) );
  OR U59400 ( .A(n48757), .B(n48756), .Z(n48758) );
  NAND U59401 ( .A(n48759), .B(n48758), .Z(n48760) );
  NANDN U59402 ( .A(n48761), .B(n48760), .Z(n48762) );
  AND U59403 ( .A(n48763), .B(n48762), .Z(n48764) );
  OR U59404 ( .A(n48765), .B(n48764), .Z(n48766) );
  NAND U59405 ( .A(n48767), .B(n48766), .Z(n48768) );
  NAND U59406 ( .A(n50711), .B(n48768), .Z(n48770) );
  NANDN U59407 ( .A(n48770), .B(n48769), .Z(n48771) );
  NAND U59408 ( .A(n48772), .B(n48771), .Z(n48773) );
  AND U59409 ( .A(n48773), .B(n60404), .Z(n48774) );
  NANDN U59410 ( .A(x[7498]), .B(y[7498]), .Z(n50710) );
  AND U59411 ( .A(n48774), .B(n50710), .Z(n48778) );
  AND U59412 ( .A(n48776), .B(n48775), .Z(n48777) );
  NANDN U59413 ( .A(n48778), .B(n48777), .Z(n48779) );
  NAND U59414 ( .A(n48780), .B(n48779), .Z(n48781) );
  NAND U59415 ( .A(n48782), .B(n48781), .Z(n48783) );
  AND U59416 ( .A(n48783), .B(n60408), .Z(n48784) );
  NANDN U59417 ( .A(x[7502]), .B(y[7502]), .Z(n50709) );
  AND U59418 ( .A(n48784), .B(n50709), .Z(n48788) );
  AND U59419 ( .A(n48786), .B(n48785), .Z(n48787) );
  NANDN U59420 ( .A(n48788), .B(n48787), .Z(n48789) );
  NAND U59421 ( .A(n48790), .B(n48789), .Z(n48791) );
  NAND U59422 ( .A(n48792), .B(n48791), .Z(n48793) );
  AND U59423 ( .A(n48793), .B(n60414), .Z(n48794) );
  NANDN U59424 ( .A(x[7506]), .B(y[7506]), .Z(n60412) );
  AND U59425 ( .A(n48794), .B(n60412), .Z(n48798) );
  AND U59426 ( .A(n48796), .B(n48795), .Z(n48797) );
  NANDN U59427 ( .A(n48798), .B(n48797), .Z(n48799) );
  NAND U59428 ( .A(n48800), .B(n48799), .Z(n48801) );
  NAND U59429 ( .A(n48802), .B(n48801), .Z(n48804) );
  AND U59430 ( .A(n48804), .B(n48803), .Z(n48805) );
  NANDN U59431 ( .A(x[7510]), .B(y[7510]), .Z(n50706) );
  AND U59432 ( .A(n48805), .B(n50706), .Z(n48809) );
  AND U59433 ( .A(n48807), .B(n48806), .Z(n48808) );
  NANDN U59434 ( .A(n48809), .B(n48808), .Z(n48810) );
  NAND U59435 ( .A(n48811), .B(n48810), .Z(n48812) );
  NAND U59436 ( .A(n48813), .B(n48812), .Z(n48814) );
  AND U59437 ( .A(n48814), .B(n60424), .Z(n48815) );
  NANDN U59438 ( .A(x[7514]), .B(y[7514]), .Z(n60422) );
  AND U59439 ( .A(n48815), .B(n60422), .Z(n48819) );
  AND U59440 ( .A(n48817), .B(n48816), .Z(n48818) );
  NANDN U59441 ( .A(n48819), .B(n48818), .Z(n48820) );
  NAND U59442 ( .A(n48821), .B(n48820), .Z(n48822) );
  NAND U59443 ( .A(n48823), .B(n48822), .Z(n48824) );
  AND U59444 ( .A(n48824), .B(n60429), .Z(n48825) );
  NANDN U59445 ( .A(x[7518]), .B(y[7518]), .Z(n50703) );
  AND U59446 ( .A(n48825), .B(n50703), .Z(n48829) );
  AND U59447 ( .A(n48827), .B(n48826), .Z(n48828) );
  NANDN U59448 ( .A(n48829), .B(n48828), .Z(n48830) );
  NAND U59449 ( .A(n48831), .B(n48830), .Z(n48832) );
  NAND U59450 ( .A(n48833), .B(n48832), .Z(n48834) );
  AND U59451 ( .A(n48834), .B(n60434), .Z(n48835) );
  NANDN U59452 ( .A(x[7522]), .B(y[7522]), .Z(n60432) );
  AND U59453 ( .A(n48835), .B(n60432), .Z(n48839) );
  AND U59454 ( .A(n48837), .B(n48836), .Z(n48838) );
  NANDN U59455 ( .A(n48839), .B(n48838), .Z(n48840) );
  NAND U59456 ( .A(n48841), .B(n48840), .Z(n48842) );
  NAND U59457 ( .A(n48843), .B(n48842), .Z(n48844) );
  AND U59458 ( .A(n48844), .B(n50700), .Z(n48845) );
  NANDN U59459 ( .A(x[7526]), .B(y[7526]), .Z(n60439) );
  AND U59460 ( .A(n48845), .B(n60439), .Z(n48849) );
  AND U59461 ( .A(n48847), .B(n48846), .Z(n48848) );
  NANDN U59462 ( .A(n48849), .B(n48848), .Z(n48850) );
  NAND U59463 ( .A(n48851), .B(n48850), .Z(n48852) );
  NAND U59464 ( .A(n48853), .B(n48852), .Z(n48854) );
  AND U59465 ( .A(n48854), .B(n50699), .Z(n48855) );
  NANDN U59466 ( .A(x[7530]), .B(y[7530]), .Z(n60443) );
  AND U59467 ( .A(n48855), .B(n60443), .Z(n48859) );
  AND U59468 ( .A(n48857), .B(n48856), .Z(n48858) );
  NANDN U59469 ( .A(n48859), .B(n48858), .Z(n48860) );
  NAND U59470 ( .A(n48861), .B(n48860), .Z(n48862) );
  NAND U59471 ( .A(n48863), .B(n48862), .Z(n48864) );
  AND U59472 ( .A(n48864), .B(n60450), .Z(n48865) );
  NANDN U59473 ( .A(x[7534]), .B(y[7534]), .Z(n60447) );
  AND U59474 ( .A(n48865), .B(n60447), .Z(n48869) );
  AND U59475 ( .A(n48867), .B(n48866), .Z(n48868) );
  NANDN U59476 ( .A(n48869), .B(n48868), .Z(n48870) );
  NAND U59477 ( .A(n48871), .B(n48870), .Z(n48872) );
  NAND U59478 ( .A(n48873), .B(n48872), .Z(n48874) );
  AND U59479 ( .A(n48874), .B(n60455), .Z(n48875) );
  NANDN U59480 ( .A(x[7538]), .B(y[7538]), .Z(n60453) );
  AND U59481 ( .A(n48875), .B(n60453), .Z(n48879) );
  AND U59482 ( .A(n48877), .B(n48876), .Z(n48878) );
  NANDN U59483 ( .A(n48879), .B(n48878), .Z(n48880) );
  NAND U59484 ( .A(n48881), .B(n48880), .Z(n48882) );
  NAND U59485 ( .A(n48883), .B(n48882), .Z(n48884) );
  AND U59486 ( .A(n48884), .B(n60459), .Z(n48885) );
  NANDN U59487 ( .A(x[7542]), .B(y[7542]), .Z(n50696) );
  AND U59488 ( .A(n48885), .B(n50696), .Z(n48889) );
  AND U59489 ( .A(n48887), .B(n48886), .Z(n48888) );
  NANDN U59490 ( .A(n48889), .B(n48888), .Z(n48890) );
  NAND U59491 ( .A(n48891), .B(n48890), .Z(n48892) );
  NAND U59492 ( .A(n48893), .B(n48892), .Z(n48894) );
  AND U59493 ( .A(n48894), .B(n60465), .Z(n48895) );
  NANDN U59494 ( .A(x[7546]), .B(y[7546]), .Z(n50694) );
  AND U59495 ( .A(n48895), .B(n50694), .Z(n48899) );
  AND U59496 ( .A(n48897), .B(n48896), .Z(n48898) );
  NANDN U59497 ( .A(n48899), .B(n48898), .Z(n48900) );
  NAND U59498 ( .A(n48901), .B(n48900), .Z(n48902) );
  NAND U59499 ( .A(n48903), .B(n48902), .Z(n48904) );
  AND U59500 ( .A(n48904), .B(n60470), .Z(n48905) );
  NANDN U59501 ( .A(x[7550]), .B(y[7550]), .Z(n60469) );
  AND U59502 ( .A(n48905), .B(n60469), .Z(n48909) );
  AND U59503 ( .A(n48907), .B(n48906), .Z(n48908) );
  NANDN U59504 ( .A(n48909), .B(n48908), .Z(n48910) );
  NAND U59505 ( .A(n48911), .B(n48910), .Z(n48912) );
  NAND U59506 ( .A(n48913), .B(n48912), .Z(n48914) );
  AND U59507 ( .A(n48914), .B(n50691), .Z(n48915) );
  NANDN U59508 ( .A(x[7554]), .B(y[7554]), .Z(n60474) );
  AND U59509 ( .A(n48915), .B(n60474), .Z(n48919) );
  AND U59510 ( .A(n48917), .B(n48916), .Z(n48918) );
  NANDN U59511 ( .A(n48919), .B(n48918), .Z(n48920) );
  NAND U59512 ( .A(n48921), .B(n48920), .Z(n48922) );
  NAND U59513 ( .A(n48923), .B(n48922), .Z(n48924) );
  AND U59514 ( .A(n48924), .B(n50689), .Z(n48925) );
  NANDN U59515 ( .A(x[7558]), .B(y[7558]), .Z(n60478) );
  AND U59516 ( .A(n48925), .B(n60478), .Z(n48929) );
  AND U59517 ( .A(n48927), .B(n48926), .Z(n48928) );
  NANDN U59518 ( .A(n48929), .B(n48928), .Z(n48930) );
  NAND U59519 ( .A(n48931), .B(n48930), .Z(n48932) );
  NAND U59520 ( .A(n48933), .B(n48932), .Z(n48934) );
  AND U59521 ( .A(n48934), .B(n60486), .Z(n48935) );
  NANDN U59522 ( .A(x[7562]), .B(y[7562]), .Z(n60484) );
  AND U59523 ( .A(n48935), .B(n60484), .Z(n48939) );
  AND U59524 ( .A(n48937), .B(n48936), .Z(n48938) );
  NANDN U59525 ( .A(n48939), .B(n48938), .Z(n48940) );
  NAND U59526 ( .A(n48941), .B(n48940), .Z(n48942) );
  NAND U59527 ( .A(n48943), .B(n48942), .Z(n48944) );
  AND U59528 ( .A(n48944), .B(n60492), .Z(n48945) );
  NANDN U59529 ( .A(x[7566]), .B(y[7566]), .Z(n60489) );
  AND U59530 ( .A(n48945), .B(n60489), .Z(n48949) );
  AND U59531 ( .A(n48947), .B(n48946), .Z(n48948) );
  NANDN U59532 ( .A(n48949), .B(n48948), .Z(n48950) );
  NAND U59533 ( .A(n48951), .B(n48950), .Z(n48952) );
  NAND U59534 ( .A(n48953), .B(n48952), .Z(n48954) );
  AND U59535 ( .A(n48954), .B(n60498), .Z(n48955) );
  NANDN U59536 ( .A(x[7570]), .B(y[7570]), .Z(n60494) );
  AND U59537 ( .A(n48955), .B(n60494), .Z(n48959) );
  AND U59538 ( .A(n48957), .B(n48956), .Z(n48958) );
  NANDN U59539 ( .A(n48959), .B(n48958), .Z(n48960) );
  NAND U59540 ( .A(n48961), .B(n48960), .Z(n48962) );
  AND U59541 ( .A(n48963), .B(n48962), .Z(n48964) );
  OR U59542 ( .A(n48965), .B(n48964), .Z(n48966) );
  NAND U59543 ( .A(n48967), .B(n48966), .Z(n48968) );
  NANDN U59544 ( .A(n60504), .B(n48968), .Z(n48969) );
  NANDN U59545 ( .A(x[7576]), .B(y[7576]), .Z(n60502) );
  NANDN U59546 ( .A(n48969), .B(n60502), .Z(n48970) );
  NAND U59547 ( .A(n48971), .B(n48970), .Z(n48973) );
  AND U59548 ( .A(n48973), .B(n48972), .Z(n48974) );
  NANDN U59549 ( .A(n60505), .B(n48974), .Z(n48975) );
  NAND U59550 ( .A(n48976), .B(n48975), .Z(n48977) );
  NANDN U59551 ( .A(n48978), .B(n48977), .Z(n48979) );
  NAND U59552 ( .A(n48980), .B(n48979), .Z(n48981) );
  AND U59553 ( .A(n48981), .B(n50684), .Z(n48982) );
  NANDN U59554 ( .A(x[7582]), .B(y[7582]), .Z(n60511) );
  AND U59555 ( .A(n48982), .B(n60511), .Z(n48986) );
  AND U59556 ( .A(n48984), .B(n48983), .Z(n48985) );
  NANDN U59557 ( .A(n48986), .B(n48985), .Z(n48987) );
  NAND U59558 ( .A(n48988), .B(n48987), .Z(n48989) );
  NAND U59559 ( .A(n48990), .B(n48989), .Z(n48991) );
  AND U59560 ( .A(n48991), .B(n60515), .Z(n48992) );
  NANDN U59561 ( .A(x[7586]), .B(y[7586]), .Z(n50681) );
  AND U59562 ( .A(n48992), .B(n50681), .Z(n48996) );
  AND U59563 ( .A(n48994), .B(n48993), .Z(n48995) );
  NANDN U59564 ( .A(n48996), .B(n48995), .Z(n48997) );
  NAND U59565 ( .A(n48998), .B(n48997), .Z(n48999) );
  NAND U59566 ( .A(n49000), .B(n48999), .Z(n49002) );
  IV U59567 ( .A(n49001), .Z(n60518) );
  AND U59568 ( .A(n49002), .B(n60518), .Z(n49003) );
  NANDN U59569 ( .A(x[7590]), .B(y[7590]), .Z(n50680) );
  AND U59570 ( .A(n49003), .B(n50680), .Z(n49007) );
  AND U59571 ( .A(n49005), .B(n49004), .Z(n49006) );
  NANDN U59572 ( .A(n49007), .B(n49006), .Z(n49008) );
  NAND U59573 ( .A(n49009), .B(n49008), .Z(n49010) );
  NAND U59574 ( .A(n49011), .B(n49010), .Z(n49012) );
  AND U59575 ( .A(n49012), .B(n60525), .Z(n49013) );
  NANDN U59576 ( .A(x[7594]), .B(y[7594]), .Z(n60523) );
  AND U59577 ( .A(n49013), .B(n60523), .Z(n49017) );
  AND U59578 ( .A(n49015), .B(n49014), .Z(n49016) );
  NANDN U59579 ( .A(n49017), .B(n49016), .Z(n49018) );
  NAND U59580 ( .A(n49019), .B(n49018), .Z(n49020) );
  NAND U59581 ( .A(n49021), .B(n49020), .Z(n49022) );
  AND U59582 ( .A(n49022), .B(n50676), .Z(n49023) );
  NANDN U59583 ( .A(x[7598]), .B(y[7598]), .Z(n60529) );
  AND U59584 ( .A(n49023), .B(n60529), .Z(n49027) );
  AND U59585 ( .A(n49025), .B(n49024), .Z(n49026) );
  NANDN U59586 ( .A(n49027), .B(n49026), .Z(n49028) );
  NAND U59587 ( .A(n49029), .B(n49028), .Z(n49030) );
  NAND U59588 ( .A(n49031), .B(n49030), .Z(n49032) );
  AND U59589 ( .A(n49032), .B(n50675), .Z(n49033) );
  NANDN U59590 ( .A(x[7602]), .B(y[7602]), .Z(n60533) );
  AND U59591 ( .A(n49033), .B(n60533), .Z(n49037) );
  AND U59592 ( .A(n49035), .B(n49034), .Z(n49036) );
  NANDN U59593 ( .A(n49037), .B(n49036), .Z(n49038) );
  NAND U59594 ( .A(n49039), .B(n49038), .Z(n49040) );
  NAND U59595 ( .A(n49041), .B(n49040), .Z(n49043) );
  IV U59596 ( .A(n49042), .Z(n60541) );
  AND U59597 ( .A(n49043), .B(n60541), .Z(n49044) );
  NANDN U59598 ( .A(x[7606]), .B(y[7606]), .Z(n60539) );
  AND U59599 ( .A(n49044), .B(n60539), .Z(n49048) );
  AND U59600 ( .A(n49046), .B(n49045), .Z(n49047) );
  NANDN U59601 ( .A(n49048), .B(n49047), .Z(n49049) );
  NAND U59602 ( .A(n49050), .B(n49049), .Z(n49051) );
  NAND U59603 ( .A(n49052), .B(n49051), .Z(n49053) );
  AND U59604 ( .A(n49053), .B(n60546), .Z(n49054) );
  NANDN U59605 ( .A(x[7610]), .B(y[7610]), .Z(n60544) );
  AND U59606 ( .A(n49054), .B(n60544), .Z(n49058) );
  AND U59607 ( .A(n49056), .B(n49055), .Z(n49057) );
  NANDN U59608 ( .A(n49058), .B(n49057), .Z(n49059) );
  NAND U59609 ( .A(n49060), .B(n49059), .Z(n49061) );
  NAND U59610 ( .A(n49062), .B(n49061), .Z(n49063) );
  AND U59611 ( .A(n49063), .B(n60550), .Z(n49064) );
  NANDN U59612 ( .A(x[7614]), .B(y[7614]), .Z(n50672) );
  AND U59613 ( .A(n49064), .B(n50672), .Z(n49068) );
  AND U59614 ( .A(n49066), .B(n49065), .Z(n49067) );
  NANDN U59615 ( .A(n49068), .B(n49067), .Z(n49069) );
  NAND U59616 ( .A(n49070), .B(n49069), .Z(n49071) );
  AND U59617 ( .A(n49072), .B(n49071), .Z(n49073) );
  OR U59618 ( .A(n49074), .B(n49073), .Z(n49075) );
  NAND U59619 ( .A(n49076), .B(n49075), .Z(n49077) );
  NANDN U59620 ( .A(n49078), .B(n49077), .Z(n49079) );
  NAND U59621 ( .A(n49080), .B(n49079), .Z(n49081) );
  AND U59622 ( .A(n49081), .B(n50662), .Z(n49082) );
  NANDN U59623 ( .A(x[7622]), .B(y[7622]), .Z(n50666) );
  AND U59624 ( .A(n49082), .B(n50666), .Z(n49086) );
  AND U59625 ( .A(n49084), .B(n49083), .Z(n49085) );
  NANDN U59626 ( .A(n49086), .B(n49085), .Z(n49087) );
  NAND U59627 ( .A(n49088), .B(n49087), .Z(n49089) );
  AND U59628 ( .A(n49090), .B(n49089), .Z(n49091) );
  ANDN U59629 ( .B(n49092), .A(n49091), .Z(n49093) );
  OR U59630 ( .A(n49094), .B(n49093), .Z(n49095) );
  NAND U59631 ( .A(n49096), .B(n49095), .Z(n49097) );
  NAND U59632 ( .A(n49098), .B(n49097), .Z(n49099) );
  AND U59633 ( .A(n49099), .B(n60565), .Z(n49100) );
  NANDN U59634 ( .A(x[7630]), .B(y[7630]), .Z(n60563) );
  AND U59635 ( .A(n49100), .B(n60563), .Z(n49104) );
  AND U59636 ( .A(n49102), .B(n49101), .Z(n49103) );
  NANDN U59637 ( .A(n49104), .B(n49103), .Z(n49105) );
  NAND U59638 ( .A(n49106), .B(n49105), .Z(n49107) );
  NAND U59639 ( .A(n49108), .B(n49107), .Z(n49109) );
  AND U59640 ( .A(n49109), .B(n60568), .Z(n49110) );
  NANDN U59641 ( .A(n50657), .B(n49110), .Z(n49111) );
  NAND U59642 ( .A(n49112), .B(n49111), .Z(n49113) );
  NANDN U59643 ( .A(n50655), .B(n49113), .Z(n49114) );
  NANDN U59644 ( .A(x[7636]), .B(y[7636]), .Z(n60569) );
  NANDN U59645 ( .A(n49114), .B(n60569), .Z(n49115) );
  NAND U59646 ( .A(n49116), .B(n49115), .Z(n49117) );
  AND U59647 ( .A(n49117), .B(n60572), .Z(n49118) );
  NANDN U59648 ( .A(x[7638]), .B(y[7638]), .Z(n50656) );
  AND U59649 ( .A(n49118), .B(n50656), .Z(n49122) );
  AND U59650 ( .A(n49120), .B(n49119), .Z(n49121) );
  NANDN U59651 ( .A(n49122), .B(n49121), .Z(n49123) );
  NAND U59652 ( .A(n49124), .B(n49123), .Z(n49125) );
  NAND U59653 ( .A(n49126), .B(n49125), .Z(n49128) );
  AND U59654 ( .A(n49128), .B(n49127), .Z(n49129) );
  NANDN U59655 ( .A(x[7642]), .B(y[7642]), .Z(n60577) );
  AND U59656 ( .A(n49129), .B(n60577), .Z(n49133) );
  AND U59657 ( .A(n49131), .B(n49130), .Z(n49132) );
  NANDN U59658 ( .A(n49133), .B(n49132), .Z(n49134) );
  NAND U59659 ( .A(n49135), .B(n49134), .Z(n49136) );
  NAND U59660 ( .A(n49137), .B(n49136), .Z(n49138) );
  AND U59661 ( .A(n49138), .B(n50653), .Z(n49139) );
  NANDN U59662 ( .A(x[7646]), .B(y[7646]), .Z(n60582) );
  AND U59663 ( .A(n49139), .B(n60582), .Z(n49143) );
  AND U59664 ( .A(n49141), .B(n49140), .Z(n49142) );
  NANDN U59665 ( .A(n49143), .B(n49142), .Z(n49144) );
  NAND U59666 ( .A(n49145), .B(n49144), .Z(n49146) );
  NAND U59667 ( .A(n49147), .B(n49146), .Z(n49148) );
  AND U59668 ( .A(n49148), .B(n60590), .Z(n49149) );
  NANDN U59669 ( .A(x[7650]), .B(y[7650]), .Z(n60586) );
  AND U59670 ( .A(n49149), .B(n60586), .Z(n49153) );
  AND U59671 ( .A(n49151), .B(n49150), .Z(n49152) );
  NANDN U59672 ( .A(n49153), .B(n49152), .Z(n49154) );
  NAND U59673 ( .A(n49155), .B(n49154), .Z(n49156) );
  NAND U59674 ( .A(n49157), .B(n49156), .Z(n49158) );
  AND U59675 ( .A(n49158), .B(n60597), .Z(n49159) );
  NANDN U59676 ( .A(x[7654]), .B(y[7654]), .Z(n60595) );
  AND U59677 ( .A(n49159), .B(n60595), .Z(n49163) );
  AND U59678 ( .A(n49161), .B(n49160), .Z(n49162) );
  NANDN U59679 ( .A(n49163), .B(n49162), .Z(n49164) );
  NAND U59680 ( .A(n49165), .B(n49164), .Z(n49166) );
  NAND U59681 ( .A(n49167), .B(n49166), .Z(n49169) );
  IV U59682 ( .A(n49168), .Z(n50649) );
  AND U59683 ( .A(n49169), .B(n50649), .Z(n49170) );
  NANDN U59684 ( .A(x[7658]), .B(y[7658]), .Z(n60600) );
  AND U59685 ( .A(n49170), .B(n60600), .Z(n49174) );
  AND U59686 ( .A(n49172), .B(n49171), .Z(n49173) );
  NANDN U59687 ( .A(n49174), .B(n49173), .Z(n49175) );
  NAND U59688 ( .A(n49176), .B(n49175), .Z(n49177) );
  NAND U59689 ( .A(n49178), .B(n49177), .Z(n49179) );
  AND U59690 ( .A(n49179), .B(n60607), .Z(n49180) );
  NANDN U59691 ( .A(x[7662]), .B(y[7662]), .Z(n60603) );
  AND U59692 ( .A(n49180), .B(n60603), .Z(n49184) );
  AND U59693 ( .A(n49182), .B(n49181), .Z(n49183) );
  NANDN U59694 ( .A(n49184), .B(n49183), .Z(n49185) );
  NAND U59695 ( .A(n49186), .B(n49185), .Z(n49187) );
  NAND U59696 ( .A(n49188), .B(n49187), .Z(n49189) );
  AND U59697 ( .A(n49189), .B(n50645), .Z(n49190) );
  NANDN U59698 ( .A(x[7666]), .B(y[7666]), .Z(n50647) );
  AND U59699 ( .A(n49190), .B(n50647), .Z(n49194) );
  AND U59700 ( .A(n49192), .B(n49191), .Z(n49193) );
  NANDN U59701 ( .A(n49194), .B(n49193), .Z(n49195) );
  NAND U59702 ( .A(n49196), .B(n49195), .Z(n49197) );
  AND U59703 ( .A(n49198), .B(n49197), .Z(n49199) );
  OR U59704 ( .A(n49200), .B(n49199), .Z(n49201) );
  NAND U59705 ( .A(n49202), .B(n49201), .Z(n49203) );
  NANDN U59706 ( .A(n49204), .B(n49203), .Z(n49206) );
  NANDN U59707 ( .A(n49206), .B(n49205), .Z(n49207) );
  NAND U59708 ( .A(n49208), .B(n49207), .Z(n49209) );
  AND U59709 ( .A(n49210), .B(n49209), .Z(n49211) );
  OR U59710 ( .A(n49212), .B(n49211), .Z(n49213) );
  NAND U59711 ( .A(n49214), .B(n49213), .Z(n49215) );
  NAND U59712 ( .A(n49216), .B(n49215), .Z(n49217) );
  AND U59713 ( .A(n49217), .B(n60622), .Z(n49218) );
  NANDN U59714 ( .A(x[7678]), .B(y[7678]), .Z(n50643) );
  AND U59715 ( .A(n49218), .B(n50643), .Z(n49222) );
  AND U59716 ( .A(n49220), .B(n49219), .Z(n49221) );
  NANDN U59717 ( .A(n49222), .B(n49221), .Z(n49223) );
  NAND U59718 ( .A(n49224), .B(n49223), .Z(n49225) );
  AND U59719 ( .A(n49226), .B(n49225), .Z(n49227) );
  OR U59720 ( .A(n49228), .B(n49227), .Z(n49229) );
  NAND U59721 ( .A(n49230), .B(n49229), .Z(n49231) );
  NANDN U59722 ( .A(n49232), .B(n49231), .Z(n49233) );
  NAND U59723 ( .A(n49234), .B(n49233), .Z(n49235) );
  AND U59724 ( .A(n49235), .B(n50634), .Z(n49236) );
  NANDN U59725 ( .A(x[7686]), .B(y[7686]), .Z(n50638) );
  AND U59726 ( .A(n49236), .B(n50638), .Z(n49240) );
  AND U59727 ( .A(n49238), .B(n49237), .Z(n49239) );
  NANDN U59728 ( .A(n49240), .B(n49239), .Z(n49241) );
  NAND U59729 ( .A(n49242), .B(n49241), .Z(n49243) );
  NAND U59730 ( .A(n49244), .B(n49243), .Z(n49246) );
  AND U59731 ( .A(n49246), .B(n49245), .Z(n49247) );
  NANDN U59732 ( .A(x[7690]), .B(y[7690]), .Z(n60630) );
  AND U59733 ( .A(n49247), .B(n60630), .Z(n49251) );
  AND U59734 ( .A(n49249), .B(n49248), .Z(n49250) );
  NANDN U59735 ( .A(n49251), .B(n49250), .Z(n49252) );
  NAND U59736 ( .A(n49253), .B(n49252), .Z(n49254) );
  NAND U59737 ( .A(n49255), .B(n49254), .Z(n49256) );
  AND U59738 ( .A(n49256), .B(n50631), .Z(n49257) );
  NANDN U59739 ( .A(x[7694]), .B(y[7694]), .Z(n60635) );
  AND U59740 ( .A(n49257), .B(n60635), .Z(n49261) );
  AND U59741 ( .A(n49259), .B(n49258), .Z(n49260) );
  NANDN U59742 ( .A(n49261), .B(n49260), .Z(n49262) );
  NAND U59743 ( .A(n49263), .B(n49262), .Z(n49264) );
  NAND U59744 ( .A(n49265), .B(n49264), .Z(n49266) );
  AND U59745 ( .A(n49267), .B(n49266), .Z(n49271) );
  AND U59746 ( .A(n49269), .B(n49268), .Z(n49270) );
  NANDN U59747 ( .A(n49271), .B(n49270), .Z(n49272) );
  NAND U59748 ( .A(n49273), .B(n49272), .Z(n49274) );
  NAND U59749 ( .A(n49275), .B(n49274), .Z(n49276) );
  AND U59750 ( .A(n49276), .B(n60645), .Z(n49277) );
  NANDN U59751 ( .A(x[7702]), .B(y[7702]), .Z(n50629) );
  AND U59752 ( .A(n49277), .B(n50629), .Z(n49281) );
  AND U59753 ( .A(n49279), .B(n49278), .Z(n49280) );
  NANDN U59754 ( .A(n49281), .B(n49280), .Z(n49282) );
  NAND U59755 ( .A(n49283), .B(n49282), .Z(n49284) );
  NAND U59756 ( .A(n49285), .B(n49284), .Z(n49286) );
  AND U59757 ( .A(n49286), .B(n60651), .Z(n49287) );
  NANDN U59758 ( .A(x[7706]), .B(y[7706]), .Z(n60649) );
  AND U59759 ( .A(n49287), .B(n60649), .Z(n49291) );
  AND U59760 ( .A(n49289), .B(n49288), .Z(n49290) );
  NANDN U59761 ( .A(n49291), .B(n49290), .Z(n49292) );
  NAND U59762 ( .A(n49293), .B(n49292), .Z(n49294) );
  NAND U59763 ( .A(n49295), .B(n49294), .Z(n49296) );
  AND U59764 ( .A(n49296), .B(n50624), .Z(n49297) );
  NANDN U59765 ( .A(x[7710]), .B(y[7710]), .Z(n60655) );
  AND U59766 ( .A(n49297), .B(n60655), .Z(n49301) );
  AND U59767 ( .A(n49299), .B(n49298), .Z(n49300) );
  NANDN U59768 ( .A(n49301), .B(n49300), .Z(n49302) );
  NAND U59769 ( .A(n49303), .B(n49302), .Z(n49304) );
  AND U59770 ( .A(n49305), .B(n49304), .Z(n49307) );
  NANDN U59771 ( .A(x[7714]), .B(y[7714]), .Z(n60660) );
  AND U59772 ( .A(n60660), .B(n50622), .Z(n49306) );
  NANDN U59773 ( .A(n49307), .B(n49306), .Z(n49308) );
  NANDN U59774 ( .A(n49309), .B(n49308), .Z(n49310) );
  AND U59775 ( .A(n60663), .B(n49310), .Z(n49311) );
  NANDN U59776 ( .A(x[7716]), .B(y[7716]), .Z(n50623) );
  NAND U59777 ( .A(n49311), .B(n50623), .Z(n49312) );
  NAND U59778 ( .A(n49313), .B(n49312), .Z(n49314) );
  AND U59779 ( .A(n49314), .B(n60666), .Z(n49315) );
  NANDN U59780 ( .A(x[7718]), .B(y[7718]), .Z(n60664) );
  AND U59781 ( .A(n49315), .B(n60664), .Z(n49319) );
  AND U59782 ( .A(n49317), .B(n49316), .Z(n49318) );
  NANDN U59783 ( .A(n49319), .B(n49318), .Z(n49320) );
  NAND U59784 ( .A(n49321), .B(n49320), .Z(n49322) );
  NAND U59785 ( .A(n49323), .B(n49322), .Z(n49324) );
  AND U59786 ( .A(n49324), .B(n60671), .Z(n49325) );
  NANDN U59787 ( .A(x[7722]), .B(y[7722]), .Z(n60669) );
  AND U59788 ( .A(n49325), .B(n60669), .Z(n49329) );
  AND U59789 ( .A(n49327), .B(n49326), .Z(n49328) );
  NANDN U59790 ( .A(n49329), .B(n49328), .Z(n49330) );
  NAND U59791 ( .A(n49331), .B(n49330), .Z(n49332) );
  NAND U59792 ( .A(n49333), .B(n49332), .Z(n49334) );
  AND U59793 ( .A(n49334), .B(n60681), .Z(n49335) );
  NANDN U59794 ( .A(x[7726]), .B(y[7726]), .Z(n50620) );
  AND U59795 ( .A(n49335), .B(n50620), .Z(n49336) );
  OR U59796 ( .A(n49337), .B(n49336), .Z(n49338) );
  NAND U59797 ( .A(n49339), .B(n49338), .Z(n49340) );
  NAND U59798 ( .A(n49341), .B(n49340), .Z(n49342) );
  AND U59799 ( .A(n49342), .B(n60691), .Z(n49343) );
  NANDN U59800 ( .A(x[7730]), .B(y[7730]), .Z(n50618) );
  AND U59801 ( .A(n49343), .B(n50618), .Z(n49347) );
  AND U59802 ( .A(n49345), .B(n49344), .Z(n49346) );
  NANDN U59803 ( .A(n49347), .B(n49346), .Z(n49348) );
  NAND U59804 ( .A(n49349), .B(n49348), .Z(n49350) );
  NAND U59805 ( .A(n49351), .B(n49350), .Z(n49352) );
  AND U59806 ( .A(n49352), .B(n60703), .Z(n49353) );
  NANDN U59807 ( .A(x[7734]), .B(y[7734]), .Z(n60698) );
  AND U59808 ( .A(n49353), .B(n60698), .Z(n49357) );
  AND U59809 ( .A(n49355), .B(n49354), .Z(n49356) );
  NANDN U59810 ( .A(n49357), .B(n49356), .Z(n49358) );
  NAND U59811 ( .A(n49359), .B(n49358), .Z(n49360) );
  NAND U59812 ( .A(n49361), .B(n49360), .Z(n49362) );
  AND U59813 ( .A(n49362), .B(n50615), .Z(n49363) );
  NANDN U59814 ( .A(x[7738]), .B(y[7738]), .Z(n60710) );
  AND U59815 ( .A(n49363), .B(n60710), .Z(n49367) );
  AND U59816 ( .A(n49365), .B(n49364), .Z(n49366) );
  NANDN U59817 ( .A(n49367), .B(n49366), .Z(n49368) );
  NAND U59818 ( .A(n49369), .B(n49368), .Z(n49370) );
  NAND U59819 ( .A(n49371), .B(n49370), .Z(n49372) );
  AND U59820 ( .A(n49372), .B(n50614), .Z(n49373) );
  NANDN U59821 ( .A(x[7742]), .B(y[7742]), .Z(n60714) );
  AND U59822 ( .A(n49373), .B(n60714), .Z(n49377) );
  AND U59823 ( .A(n49375), .B(n49374), .Z(n49376) );
  NANDN U59824 ( .A(n49377), .B(n49376), .Z(n49378) );
  NAND U59825 ( .A(n49379), .B(n49378), .Z(n49380) );
  NAND U59826 ( .A(n49381), .B(n49380), .Z(n49382) );
  AND U59827 ( .A(n49382), .B(n60719), .Z(n49383) );
  NANDN U59828 ( .A(x[7746]), .B(y[7746]), .Z(n60717) );
  AND U59829 ( .A(n49383), .B(n60717), .Z(n49387) );
  AND U59830 ( .A(n49385), .B(n49384), .Z(n49386) );
  NANDN U59831 ( .A(n49387), .B(n49386), .Z(n49388) );
  NAND U59832 ( .A(n49389), .B(n49388), .Z(n49390) );
  NAND U59833 ( .A(n49391), .B(n49390), .Z(n49392) );
  AND U59834 ( .A(n49392), .B(n60725), .Z(n49393) );
  NANDN U59835 ( .A(x[7750]), .B(y[7750]), .Z(n60723) );
  AND U59836 ( .A(n49393), .B(n60723), .Z(n49397) );
  AND U59837 ( .A(n49395), .B(n49394), .Z(n49396) );
  NANDN U59838 ( .A(n49397), .B(n49396), .Z(n49398) );
  NAND U59839 ( .A(n49399), .B(n49398), .Z(n49400) );
  NAND U59840 ( .A(n49401), .B(n49400), .Z(n49402) );
  AND U59841 ( .A(n49402), .B(n60729), .Z(n49403) );
  NANDN U59842 ( .A(x[7754]), .B(y[7754]), .Z(n50610) );
  AND U59843 ( .A(n49403), .B(n50610), .Z(n49407) );
  AND U59844 ( .A(n49405), .B(n49404), .Z(n49406) );
  NANDN U59845 ( .A(n49407), .B(n49406), .Z(n49408) );
  NAND U59846 ( .A(n49409), .B(n49408), .Z(n49410) );
  NAND U59847 ( .A(n49411), .B(n49410), .Z(n49413) );
  IV U59848 ( .A(n49412), .Z(n60732) );
  AND U59849 ( .A(n49413), .B(n60732), .Z(n49414) );
  NANDN U59850 ( .A(x[7758]), .B(y[7758]), .Z(n50608) );
  AND U59851 ( .A(n49414), .B(n50608), .Z(n49418) );
  AND U59852 ( .A(n49416), .B(n49415), .Z(n49417) );
  NANDN U59853 ( .A(n49418), .B(n49417), .Z(n49419) );
  NAND U59854 ( .A(n49420), .B(n49419), .Z(n49421) );
  NAND U59855 ( .A(n49422), .B(n49421), .Z(n49423) );
  AND U59856 ( .A(n49423), .B(n60739), .Z(n49424) );
  NANDN U59857 ( .A(x[7762]), .B(y[7762]), .Z(n60737) );
  AND U59858 ( .A(n49424), .B(n60737), .Z(n49428) );
  AND U59859 ( .A(n49426), .B(n49425), .Z(n49427) );
  NANDN U59860 ( .A(n49428), .B(n49427), .Z(n49429) );
  NAND U59861 ( .A(n49430), .B(n49429), .Z(n49431) );
  AND U59862 ( .A(n49432), .B(n49431), .Z(n49433) );
  OR U59863 ( .A(n49434), .B(n49433), .Z(n49435) );
  NAND U59864 ( .A(n49436), .B(n49435), .Z(n49437) );
  NANDN U59865 ( .A(n49438), .B(n49437), .Z(n49439) );
  NANDN U59866 ( .A(x[7768]), .B(y[7768]), .Z(n50605) );
  NANDN U59867 ( .A(n49439), .B(n50605), .Z(n49440) );
  AND U59868 ( .A(n49441), .B(n49440), .Z(n49442) );
  OR U59869 ( .A(n49443), .B(n49442), .Z(n49444) );
  NAND U59870 ( .A(n49445), .B(n49444), .Z(n49446) );
  NANDN U59871 ( .A(n49447), .B(n49446), .Z(n49448) );
  NANDN U59872 ( .A(n49448), .B(n60748), .Z(n49449) );
  NAND U59873 ( .A(n49450), .B(n49449), .Z(n49451) );
  AND U59874 ( .A(n49451), .B(n60751), .Z(n49452) );
  NANDN U59875 ( .A(x[7774]), .B(y[7774]), .Z(n60749) );
  AND U59876 ( .A(n49452), .B(n60749), .Z(n49456) );
  AND U59877 ( .A(n49454), .B(n49453), .Z(n49455) );
  NANDN U59878 ( .A(n49456), .B(n49455), .Z(n49457) );
  NAND U59879 ( .A(n49458), .B(n49457), .Z(n49459) );
  NAND U59880 ( .A(n49460), .B(n49459), .Z(n49461) );
  AND U59881 ( .A(n49461), .B(n60755), .Z(n49462) );
  NANDN U59882 ( .A(x[7778]), .B(y[7778]), .Z(n50601) );
  AND U59883 ( .A(n49462), .B(n50601), .Z(n49466) );
  AND U59884 ( .A(n49464), .B(n49463), .Z(n49465) );
  NANDN U59885 ( .A(n49466), .B(n49465), .Z(n49467) );
  NAND U59886 ( .A(n49468), .B(n49467), .Z(n49469) );
  NAND U59887 ( .A(n49470), .B(n49469), .Z(n49471) );
  AND U59888 ( .A(n49471), .B(n60760), .Z(n49472) );
  NANDN U59889 ( .A(x[7782]), .B(y[7782]), .Z(n50599) );
  AND U59890 ( .A(n49472), .B(n50599), .Z(n49476) );
  AND U59891 ( .A(n49474), .B(n49473), .Z(n49475) );
  NANDN U59892 ( .A(n49476), .B(n49475), .Z(n49477) );
  NAND U59893 ( .A(n49478), .B(n49477), .Z(n49479) );
  NAND U59894 ( .A(n49480), .B(n49479), .Z(n49482) );
  IV U59895 ( .A(n49481), .Z(n50594) );
  AND U59896 ( .A(n49482), .B(n50594), .Z(n49483) );
  NANDN U59897 ( .A(x[7786]), .B(y[7786]), .Z(n50597) );
  AND U59898 ( .A(n49483), .B(n50597), .Z(n49487) );
  AND U59899 ( .A(n49485), .B(n49484), .Z(n49486) );
  NANDN U59900 ( .A(n49487), .B(n49486), .Z(n49488) );
  NAND U59901 ( .A(n49489), .B(n49488), .Z(n49490) );
  NAND U59902 ( .A(n49491), .B(n49490), .Z(n49492) );
  AND U59903 ( .A(n49492), .B(n50593), .Z(n49493) );
  NANDN U59904 ( .A(x[7790]), .B(y[7790]), .Z(n60766) );
  AND U59905 ( .A(n49493), .B(n60766), .Z(n49497) );
  AND U59906 ( .A(n49495), .B(n49494), .Z(n49496) );
  NANDN U59907 ( .A(n49497), .B(n49496), .Z(n49498) );
  NAND U59908 ( .A(n49499), .B(n49498), .Z(n49500) );
  NAND U59909 ( .A(n49501), .B(n49500), .Z(n49502) );
  AND U59910 ( .A(n49502), .B(n60773), .Z(n49503) );
  NANDN U59911 ( .A(x[7794]), .B(y[7794]), .Z(n60770) );
  AND U59912 ( .A(n49503), .B(n60770), .Z(n49507) );
  AND U59913 ( .A(n49505), .B(n49504), .Z(n49506) );
  NANDN U59914 ( .A(n49507), .B(n49506), .Z(n49508) );
  NAND U59915 ( .A(n49509), .B(n49508), .Z(n49510) );
  NAND U59916 ( .A(n49511), .B(n49510), .Z(n49512) );
  AND U59917 ( .A(n49512), .B(n50590), .Z(n49513) );
  NANDN U59918 ( .A(x[7798]), .B(y[7798]), .Z(n60776) );
  AND U59919 ( .A(n49513), .B(n60776), .Z(n49517) );
  AND U59920 ( .A(n49515), .B(n49514), .Z(n49516) );
  NANDN U59921 ( .A(n49517), .B(n49516), .Z(n49518) );
  NAND U59922 ( .A(n49519), .B(n49518), .Z(n49520) );
  NAND U59923 ( .A(n49521), .B(n49520), .Z(n49522) );
  AND U59924 ( .A(n49522), .B(n60779), .Z(n49523) );
  NANDN U59925 ( .A(x[7802]), .B(y[7802]), .Z(n50586) );
  AND U59926 ( .A(n49523), .B(n50586), .Z(n49527) );
  AND U59927 ( .A(n49525), .B(n49524), .Z(n49526) );
  NANDN U59928 ( .A(n49527), .B(n49526), .Z(n49528) );
  NAND U59929 ( .A(n49529), .B(n49528), .Z(n49530) );
  NAND U59930 ( .A(n49531), .B(n49530), .Z(n49532) );
  AND U59931 ( .A(n49532), .B(n60791), .Z(n49533) );
  NANDN U59932 ( .A(x[7806]), .B(y[7806]), .Z(n60784) );
  AND U59933 ( .A(n49533), .B(n60784), .Z(n49537) );
  AND U59934 ( .A(n49535), .B(n49534), .Z(n49536) );
  NANDN U59935 ( .A(n49537), .B(n49536), .Z(n49538) );
  NAND U59936 ( .A(n49539), .B(n49538), .Z(n49540) );
  NAND U59937 ( .A(n49541), .B(n49540), .Z(n49542) );
  AND U59938 ( .A(n49542), .B(n60803), .Z(n49543) );
  NANDN U59939 ( .A(x[7810]), .B(y[7810]), .Z(n60798) );
  AND U59940 ( .A(n49543), .B(n60798), .Z(n49547) );
  AND U59941 ( .A(n49545), .B(n49544), .Z(n49546) );
  NANDN U59942 ( .A(n49547), .B(n49546), .Z(n49548) );
  NAND U59943 ( .A(n49549), .B(n49548), .Z(n49550) );
  AND U59944 ( .A(n49551), .B(n49550), .Z(n49552) );
  ANDN U59945 ( .B(n50584), .A(n49552), .Z(n49553) );
  NAND U59946 ( .A(n60810), .B(n49553), .Z(n49554) );
  NANDN U59947 ( .A(n49555), .B(n49554), .Z(n49556) );
  AND U59948 ( .A(n49556), .B(n60819), .Z(n49557) );
  NANDN U59949 ( .A(x[7816]), .B(y[7816]), .Z(n50585) );
  NAND U59950 ( .A(n49557), .B(n50585), .Z(n49558) );
  NAND U59951 ( .A(n49559), .B(n49558), .Z(n49560) );
  AND U59952 ( .A(n49560), .B(n50583), .Z(n49561) );
  NANDN U59953 ( .A(x[7818]), .B(y[7818]), .Z(n60820) );
  AND U59954 ( .A(n49561), .B(n60820), .Z(n49565) );
  AND U59955 ( .A(n49563), .B(n49562), .Z(n49564) );
  NANDN U59956 ( .A(n49565), .B(n49564), .Z(n49566) );
  NAND U59957 ( .A(n49567), .B(n49566), .Z(n49568) );
  NAND U59958 ( .A(n49569), .B(n49568), .Z(n49570) );
  AND U59959 ( .A(n49570), .B(n60828), .Z(n49571) );
  NANDN U59960 ( .A(x[7822]), .B(y[7822]), .Z(n60826) );
  AND U59961 ( .A(n49571), .B(n60826), .Z(n49575) );
  AND U59962 ( .A(n49573), .B(n49572), .Z(n49574) );
  NANDN U59963 ( .A(n49575), .B(n49574), .Z(n49576) );
  NAND U59964 ( .A(n49577), .B(n49576), .Z(n49578) );
  NAND U59965 ( .A(n49579), .B(n49578), .Z(n49580) );
  AND U59966 ( .A(n49580), .B(n60833), .Z(n49581) );
  NANDN U59967 ( .A(x[7826]), .B(y[7826]), .Z(n60831) );
  AND U59968 ( .A(n49581), .B(n60831), .Z(n49585) );
  AND U59969 ( .A(n49583), .B(n49582), .Z(n49584) );
  NANDN U59970 ( .A(n49585), .B(n49584), .Z(n49586) );
  NAND U59971 ( .A(n49587), .B(n49586), .Z(n49588) );
  NAND U59972 ( .A(n49589), .B(n49588), .Z(n49590) );
  AND U59973 ( .A(n49590), .B(n60840), .Z(n49591) );
  NANDN U59974 ( .A(x[7830]), .B(y[7830]), .Z(n50579) );
  AND U59975 ( .A(n49591), .B(n50579), .Z(n49595) );
  AND U59976 ( .A(n49593), .B(n49592), .Z(n49594) );
  NANDN U59977 ( .A(n49595), .B(n49594), .Z(n49596) );
  NAND U59978 ( .A(n49597), .B(n49596), .Z(n49598) );
  AND U59979 ( .A(n49599), .B(n49598), .Z(n49600) );
  ANDN U59980 ( .B(n49601), .A(n49600), .Z(n49602) );
  OR U59981 ( .A(n49603), .B(n49602), .Z(n49604) );
  NAND U59982 ( .A(n49605), .B(n49604), .Z(n49606) );
  NAND U59983 ( .A(n49607), .B(n49606), .Z(n49609) );
  AND U59984 ( .A(n49609), .B(n49608), .Z(n49610) );
  NANDN U59985 ( .A(x[7838]), .B(y[7838]), .Z(n60847) );
  AND U59986 ( .A(n49610), .B(n60847), .Z(n49614) );
  AND U59987 ( .A(n49612), .B(n49611), .Z(n49613) );
  NANDN U59988 ( .A(n49614), .B(n49613), .Z(n49615) );
  NAND U59989 ( .A(n49616), .B(n49615), .Z(n49617) );
  NAND U59990 ( .A(n49618), .B(n49617), .Z(n49620) );
  IV U59991 ( .A(n49619), .Z(n50572) );
  AND U59992 ( .A(n49620), .B(n50572), .Z(n49621) );
  NANDN U59993 ( .A(n60851), .B(n49621), .Z(n49622) );
  NAND U59994 ( .A(n49623), .B(n49622), .Z(n49624) );
  NANDN U59995 ( .A(n60856), .B(n49624), .Z(n49625) );
  NANDN U59996 ( .A(x[7844]), .B(y[7844]), .Z(n50573) );
  NANDN U59997 ( .A(n49625), .B(n50573), .Z(n49626) );
  NAND U59998 ( .A(n49627), .B(n49626), .Z(n49628) );
  AND U59999 ( .A(n49628), .B(n60859), .Z(n49629) );
  NANDN U60000 ( .A(x[7846]), .B(y[7846]), .Z(n60857) );
  AND U60001 ( .A(n49629), .B(n60857), .Z(n49633) );
  AND U60002 ( .A(n49631), .B(n49630), .Z(n49632) );
  NANDN U60003 ( .A(n49633), .B(n49632), .Z(n49634) );
  NAND U60004 ( .A(n49635), .B(n49634), .Z(n49636) );
  NAND U60005 ( .A(n49637), .B(n49636), .Z(n49638) );
  AND U60006 ( .A(n49638), .B(n60864), .Z(n49639) );
  NANDN U60007 ( .A(x[7850]), .B(y[7850]), .Z(n60862) );
  AND U60008 ( .A(n49639), .B(n60862), .Z(n49643) );
  AND U60009 ( .A(n49641), .B(n49640), .Z(n49642) );
  NANDN U60010 ( .A(n49643), .B(n49642), .Z(n49644) );
  NAND U60011 ( .A(n49645), .B(n49644), .Z(n49646) );
  NAND U60012 ( .A(n49647), .B(n49646), .Z(n49648) );
  AND U60013 ( .A(n49648), .B(n60870), .Z(n49649) );
  NANDN U60014 ( .A(x[7854]), .B(y[7854]), .Z(n50570) );
  AND U60015 ( .A(n49649), .B(n50570), .Z(n49653) );
  AND U60016 ( .A(n49651), .B(n49650), .Z(n49652) );
  NANDN U60017 ( .A(n49653), .B(n49652), .Z(n49654) );
  NAND U60018 ( .A(n49655), .B(n49654), .Z(n49656) );
  NAND U60019 ( .A(n49657), .B(n49656), .Z(n49658) );
  AND U60020 ( .A(n49658), .B(n60877), .Z(n49659) );
  NANDN U60021 ( .A(x[7858]), .B(y[7858]), .Z(n60873) );
  AND U60022 ( .A(n49659), .B(n60873), .Z(n49660) );
  OR U60023 ( .A(n49661), .B(n49660), .Z(n49662) );
  AND U60024 ( .A(n49663), .B(n49662), .Z(n49664) );
  OR U60025 ( .A(n49665), .B(n49664), .Z(n49666) );
  NAND U60026 ( .A(n49667), .B(n49666), .Z(n49668) );
  NANDN U60027 ( .A(n49669), .B(n49668), .Z(n49670) );
  OR U60028 ( .A(n49671), .B(n49670), .Z(n49672) );
  NAND U60029 ( .A(n49673), .B(n49672), .Z(n49674) );
  AND U60030 ( .A(n49675), .B(n49674), .Z(n49676) );
  OR U60031 ( .A(n49677), .B(n49676), .Z(n49678) );
  NAND U60032 ( .A(n49679), .B(n49678), .Z(n49680) );
  NANDN U60033 ( .A(n49681), .B(n49680), .Z(n49682) );
  NAND U60034 ( .A(n49683), .B(n49682), .Z(n49685) );
  AND U60035 ( .A(n49685), .B(n49684), .Z(n49686) );
  NAND U60036 ( .A(n50565), .B(n49686), .Z(n49687) );
  NAND U60037 ( .A(n49688), .B(n49687), .Z(n49689) );
  NANDN U60038 ( .A(n49690), .B(n49689), .Z(n49691) );
  NAND U60039 ( .A(n49692), .B(n49691), .Z(n49694) );
  AND U60040 ( .A(n49694), .B(n49693), .Z(n49695) );
  NANDN U60041 ( .A(n60890), .B(n49695), .Z(n49696) );
  NAND U60042 ( .A(n49697), .B(n49696), .Z(n49698) );
  NANDN U60043 ( .A(n49699), .B(n49698), .Z(n49700) );
  AND U60044 ( .A(n49701), .B(n49700), .Z(n49702) );
  OR U60045 ( .A(n49703), .B(n49702), .Z(n49704) );
  NAND U60046 ( .A(n49705), .B(n49704), .Z(n49706) );
  NANDN U60047 ( .A(n49707), .B(n49706), .Z(n49708) );
  NAND U60048 ( .A(n49709), .B(n49708), .Z(n49710) );
  AND U60049 ( .A(n49711), .B(n49710), .Z(n49715) );
  AND U60050 ( .A(n49713), .B(n49712), .Z(n49714) );
  NANDN U60051 ( .A(n49715), .B(n49714), .Z(n49716) );
  NAND U60052 ( .A(n49717), .B(n49716), .Z(n49718) );
  NAND U60053 ( .A(n49719), .B(n49718), .Z(n49720) );
  AND U60054 ( .A(n49720), .B(n60905), .Z(n49721) );
  NANDN U60055 ( .A(x[7886]), .B(y[7886]), .Z(n50559) );
  AND U60056 ( .A(n49721), .B(n50559), .Z(n49725) );
  AND U60057 ( .A(n49723), .B(n49722), .Z(n49724) );
  NANDN U60058 ( .A(n49725), .B(n49724), .Z(n49726) );
  NAND U60059 ( .A(n49727), .B(n49726), .Z(n49728) );
  AND U60060 ( .A(n49729), .B(n49728), .Z(n49730) );
  ANDN U60061 ( .B(n60910), .A(n49730), .Z(n49731) );
  NANDN U60062 ( .A(x[7890]), .B(y[7890]), .Z(n50558) );
  AND U60063 ( .A(n49731), .B(n50558), .Z(n49732) );
  OR U60064 ( .A(n49733), .B(n49732), .Z(n49734) );
  NAND U60065 ( .A(n49735), .B(n49734), .Z(n49736) );
  NAND U60066 ( .A(n49737), .B(n49736), .Z(n49739) );
  IV U60067 ( .A(n49738), .Z(n60915) );
  AND U60068 ( .A(n49739), .B(n60915), .Z(n49740) );
  NANDN U60069 ( .A(x[7894]), .B(y[7894]), .Z(n60914) );
  AND U60070 ( .A(n49740), .B(n60914), .Z(n49744) );
  AND U60071 ( .A(n49742), .B(n49741), .Z(n49743) );
  NANDN U60072 ( .A(n49744), .B(n49743), .Z(n49745) );
  NAND U60073 ( .A(n49746), .B(n49745), .Z(n49747) );
  NAND U60074 ( .A(n49748), .B(n49747), .Z(n49749) );
  AND U60075 ( .A(n49749), .B(n50554), .Z(n49750) );
  NANDN U60076 ( .A(x[7898]), .B(y[7898]), .Z(n60919) );
  AND U60077 ( .A(n49750), .B(n60919), .Z(n49754) );
  AND U60078 ( .A(n49752), .B(n49751), .Z(n49753) );
  NANDN U60079 ( .A(n49754), .B(n49753), .Z(n49755) );
  NAND U60080 ( .A(n49756), .B(n49755), .Z(n49757) );
  NAND U60081 ( .A(n49758), .B(n49757), .Z(n49759) );
  AND U60082 ( .A(n49759), .B(n50553), .Z(n49760) );
  NANDN U60083 ( .A(x[7902]), .B(y[7902]), .Z(n60923) );
  AND U60084 ( .A(n49760), .B(n60923), .Z(n49764) );
  AND U60085 ( .A(n49762), .B(n49761), .Z(n49763) );
  NANDN U60086 ( .A(n49764), .B(n49763), .Z(n49765) );
  NAND U60087 ( .A(n49766), .B(n49765), .Z(n49767) );
  NAND U60088 ( .A(n49768), .B(n49767), .Z(n49769) );
  AND U60089 ( .A(n49769), .B(n60931), .Z(n49770) );
  NANDN U60090 ( .A(x[7906]), .B(y[7906]), .Z(n60929) );
  AND U60091 ( .A(n49770), .B(n60929), .Z(n49774) );
  AND U60092 ( .A(n49772), .B(n49771), .Z(n49773) );
  NANDN U60093 ( .A(n49774), .B(n49773), .Z(n49775) );
  NAND U60094 ( .A(n49776), .B(n49775), .Z(n49777) );
  NAND U60095 ( .A(n49778), .B(n49777), .Z(n49779) );
  AND U60096 ( .A(n49779), .B(n60935), .Z(n49780) );
  NANDN U60097 ( .A(x[7910]), .B(y[7910]), .Z(n60933) );
  AND U60098 ( .A(n49780), .B(n60933), .Z(n49784) );
  AND U60099 ( .A(n49782), .B(n49781), .Z(n49783) );
  NANDN U60100 ( .A(n49784), .B(n49783), .Z(n49785) );
  NAND U60101 ( .A(n49786), .B(n49785), .Z(n49787) );
  NAND U60102 ( .A(n49788), .B(n49787), .Z(n49789) );
  AND U60103 ( .A(n49789), .B(n60941), .Z(n49790) );
  NANDN U60104 ( .A(x[7914]), .B(y[7914]), .Z(n50549) );
  AND U60105 ( .A(n49790), .B(n50549), .Z(n49794) );
  AND U60106 ( .A(n49792), .B(n49791), .Z(n49793) );
  NANDN U60107 ( .A(n49794), .B(n49793), .Z(n49795) );
  NAND U60108 ( .A(n49796), .B(n49795), .Z(n49797) );
  NAND U60109 ( .A(n49798), .B(n49797), .Z(n49799) );
  AND U60110 ( .A(n49799), .B(n60945), .Z(n49800) );
  NANDN U60111 ( .A(x[7918]), .B(y[7918]), .Z(n50547) );
  AND U60112 ( .A(n49800), .B(n50547), .Z(n49804) );
  AND U60113 ( .A(n49802), .B(n49801), .Z(n49803) );
  NANDN U60114 ( .A(n49804), .B(n49803), .Z(n49805) );
  NAND U60115 ( .A(n49806), .B(n49805), .Z(n49807) );
  NAND U60116 ( .A(n49808), .B(n49807), .Z(n49810) );
  IV U60117 ( .A(n49809), .Z(n60950) );
  AND U60118 ( .A(n49810), .B(n60950), .Z(n49811) );
  NANDN U60119 ( .A(x[7922]), .B(y[7922]), .Z(n60949) );
  AND U60120 ( .A(n49811), .B(n60949), .Z(n49815) );
  AND U60121 ( .A(n49813), .B(n49812), .Z(n49814) );
  NANDN U60122 ( .A(n49815), .B(n49814), .Z(n49816) );
  NAND U60123 ( .A(n49817), .B(n49816), .Z(n49818) );
  NAND U60124 ( .A(n49819), .B(n49818), .Z(n49820) );
  AND U60125 ( .A(n49820), .B(n50543), .Z(n49821) );
  NANDN U60126 ( .A(x[7926]), .B(y[7926]), .Z(n60955) );
  AND U60127 ( .A(n49821), .B(n60955), .Z(n49825) );
  AND U60128 ( .A(n49823), .B(n49822), .Z(n49824) );
  NANDN U60129 ( .A(n49825), .B(n49824), .Z(n49826) );
  NAND U60130 ( .A(n49827), .B(n49826), .Z(n49828) );
  NAND U60131 ( .A(n49829), .B(n49828), .Z(n49830) );
  AND U60132 ( .A(n49830), .B(n50542), .Z(n49831) );
  NANDN U60133 ( .A(x[7930]), .B(y[7930]), .Z(n60959) );
  AND U60134 ( .A(n49831), .B(n60959), .Z(n49835) );
  AND U60135 ( .A(n49833), .B(n49832), .Z(n49834) );
  NANDN U60136 ( .A(n49835), .B(n49834), .Z(n49836) );
  NAND U60137 ( .A(n49837), .B(n49836), .Z(n49838) );
  NAND U60138 ( .A(n49839), .B(n49838), .Z(n49840) );
  AND U60139 ( .A(n49840), .B(n60965), .Z(n49841) );
  NANDN U60140 ( .A(x[7934]), .B(y[7934]), .Z(n60962) );
  AND U60141 ( .A(n49841), .B(n60962), .Z(n49845) );
  AND U60142 ( .A(n49843), .B(n49842), .Z(n49844) );
  NANDN U60143 ( .A(n49845), .B(n49844), .Z(n49846) );
  NAND U60144 ( .A(n49847), .B(n49846), .Z(n49848) );
  NAND U60145 ( .A(n49849), .B(n49848), .Z(n49850) );
  AND U60146 ( .A(n49850), .B(n60970), .Z(n49851) );
  NANDN U60147 ( .A(x[7938]), .B(y[7938]), .Z(n60968) );
  AND U60148 ( .A(n49851), .B(n60968), .Z(n49855) );
  AND U60149 ( .A(n49853), .B(n49852), .Z(n49854) );
  NANDN U60150 ( .A(n49855), .B(n49854), .Z(n49856) );
  NAND U60151 ( .A(n49857), .B(n49856), .Z(n49858) );
  AND U60152 ( .A(n49859), .B(n49858), .Z(n49860) );
  ANDN U60153 ( .B(n49861), .A(n49860), .Z(n49862) );
  OR U60154 ( .A(n49863), .B(n49862), .Z(n49864) );
  NAND U60155 ( .A(n49865), .B(n49864), .Z(n49866) );
  NAND U60156 ( .A(n49867), .B(n49866), .Z(n49869) );
  IV U60157 ( .A(n49868), .Z(n60977) );
  AND U60158 ( .A(n49869), .B(n60977), .Z(n49870) );
  NANDN U60159 ( .A(x[7946]), .B(y[7946]), .Z(n50536) );
  AND U60160 ( .A(n49870), .B(n50536), .Z(n49874) );
  AND U60161 ( .A(n49872), .B(n49871), .Z(n49873) );
  NANDN U60162 ( .A(n49874), .B(n49873), .Z(n49875) );
  NAND U60163 ( .A(n49876), .B(n49875), .Z(n49877) );
  NAND U60164 ( .A(n49878), .B(n49877), .Z(n49880) );
  IV U60165 ( .A(n49879), .Z(n60982) );
  AND U60166 ( .A(n49880), .B(n60982), .Z(n49881) );
  NANDN U60167 ( .A(n50533), .B(n49881), .Z(n49882) );
  NAND U60168 ( .A(n49883), .B(n49882), .Z(n49884) );
  NANDN U60169 ( .A(n60985), .B(n49884), .Z(n49885) );
  NANDN U60170 ( .A(x[7952]), .B(y[7952]), .Z(n60983) );
  NANDN U60171 ( .A(n49885), .B(n60983), .Z(n49886) );
  NAND U60172 ( .A(n49887), .B(n49886), .Z(n49888) );
  AND U60173 ( .A(n49888), .B(n50530), .Z(n49889) );
  NANDN U60174 ( .A(x[7954]), .B(y[7954]), .Z(n60986) );
  AND U60175 ( .A(n49889), .B(n60986), .Z(n49893) );
  AND U60176 ( .A(n49891), .B(n49890), .Z(n49892) );
  NANDN U60177 ( .A(n49893), .B(n49892), .Z(n49894) );
  NAND U60178 ( .A(n49895), .B(n49894), .Z(n49896) );
  AND U60179 ( .A(n49897), .B(n49896), .Z(n49898) );
  OR U60180 ( .A(n49899), .B(n49898), .Z(n49900) );
  NAND U60181 ( .A(n49901), .B(n49900), .Z(n49902) );
  NANDN U60182 ( .A(n60996), .B(n49902), .Z(n49903) );
  NANDN U60183 ( .A(x[7960]), .B(y[7960]), .Z(n60991) );
  NANDN U60184 ( .A(n49903), .B(n60991), .Z(n49904) );
  NAND U60185 ( .A(n49905), .B(n49904), .Z(n49906) );
  AND U60186 ( .A(n49906), .B(n50529), .Z(n49907) );
  NANDN U60187 ( .A(x[7962]), .B(y[7962]), .Z(n60997) );
  AND U60188 ( .A(n49907), .B(n60997), .Z(n49911) );
  AND U60189 ( .A(n49909), .B(n49908), .Z(n49910) );
  NANDN U60190 ( .A(n49911), .B(n49910), .Z(n49912) );
  NAND U60191 ( .A(n49913), .B(n49912), .Z(n49914) );
  AND U60192 ( .A(n49915), .B(n49914), .Z(n49916) );
  OR U60193 ( .A(n49917), .B(n49916), .Z(n49918) );
  NAND U60194 ( .A(n49919), .B(n49918), .Z(n49920) );
  NANDN U60195 ( .A(n49921), .B(n49920), .Z(n49922) );
  NANDN U60196 ( .A(n49922), .B(n61004), .Z(n49923) );
  NAND U60197 ( .A(n49924), .B(n49923), .Z(n49926) );
  IV U60198 ( .A(n49925), .Z(n61005) );
  AND U60199 ( .A(n49926), .B(n61005), .Z(n49927) );
  NANDN U60200 ( .A(x[7970]), .B(y[7970]), .Z(n61003) );
  AND U60201 ( .A(n49927), .B(n61003), .Z(n49931) );
  AND U60202 ( .A(n49929), .B(n49928), .Z(n49930) );
  NANDN U60203 ( .A(n49931), .B(n49930), .Z(n49932) );
  NAND U60204 ( .A(n49933), .B(n49932), .Z(n49934) );
  NAND U60205 ( .A(n49935), .B(n49934), .Z(n49936) );
  AND U60206 ( .A(n49936), .B(n61012), .Z(n49937) );
  NANDN U60207 ( .A(x[7974]), .B(y[7974]), .Z(n61010) );
  AND U60208 ( .A(n49937), .B(n61010), .Z(n49941) );
  AND U60209 ( .A(n49939), .B(n49938), .Z(n49940) );
  NANDN U60210 ( .A(n49941), .B(n49940), .Z(n49942) );
  NAND U60211 ( .A(n49943), .B(n49942), .Z(n49944) );
  AND U60212 ( .A(n49945), .B(n49944), .Z(n49947) );
  NANDN U60213 ( .A(x[7978]), .B(y[7978]), .Z(n61016) );
  AND U60214 ( .A(n61016), .B(n50524), .Z(n49946) );
  NANDN U60215 ( .A(n49947), .B(n49946), .Z(n49948) );
  NANDN U60216 ( .A(n49949), .B(n49948), .Z(n49950) );
  AND U60217 ( .A(n61019), .B(n49950), .Z(n49951) );
  NANDN U60218 ( .A(x[7980]), .B(y[7980]), .Z(n50525) );
  NAND U60219 ( .A(n49951), .B(n50525), .Z(n49952) );
  NAND U60220 ( .A(n49953), .B(n49952), .Z(n49954) );
  AND U60221 ( .A(n49954), .B(n50523), .Z(n49955) );
  NANDN U60222 ( .A(x[7982]), .B(y[7982]), .Z(n61020) );
  AND U60223 ( .A(n49955), .B(n61020), .Z(n49959) );
  AND U60224 ( .A(n49957), .B(n49956), .Z(n49958) );
  NANDN U60225 ( .A(n49959), .B(n49958), .Z(n49960) );
  NAND U60226 ( .A(n49961), .B(n49960), .Z(n49962) );
  NAND U60227 ( .A(n49963), .B(n49962), .Z(n49964) );
  AND U60228 ( .A(n49964), .B(n61027), .Z(n49965) );
  NANDN U60229 ( .A(x[7986]), .B(y[7986]), .Z(n61025) );
  AND U60230 ( .A(n49965), .B(n61025), .Z(n49969) );
  AND U60231 ( .A(n49967), .B(n49966), .Z(n49968) );
  NANDN U60232 ( .A(n49969), .B(n49968), .Z(n49970) );
  NAND U60233 ( .A(n49971), .B(n49970), .Z(n49972) );
  NAND U60234 ( .A(n49973), .B(n49972), .Z(n49974) );
  AND U60235 ( .A(n49974), .B(n61032), .Z(n49975) );
  NANDN U60236 ( .A(x[7990]), .B(y[7990]), .Z(n61030) );
  AND U60237 ( .A(n49975), .B(n61030), .Z(n49976) );
  OR U60238 ( .A(n49977), .B(n49976), .Z(n49978) );
  NAND U60239 ( .A(n49979), .B(n49978), .Z(n49980) );
  NAND U60240 ( .A(n49981), .B(n49980), .Z(n49982) );
  AND U60241 ( .A(n49982), .B(n61037), .Z(n49983) );
  NANDN U60242 ( .A(x[7994]), .B(y[7994]), .Z(n50519) );
  AND U60243 ( .A(n49983), .B(n50519), .Z(n49987) );
  AND U60244 ( .A(n49985), .B(n49984), .Z(n49986) );
  NANDN U60245 ( .A(n49987), .B(n49986), .Z(n49988) );
  NAND U60246 ( .A(n49989), .B(n49988), .Z(n49990) );
  AND U60247 ( .A(n49991), .B(n49990), .Z(n49992) );
  ANDN U60248 ( .B(n50517), .A(n49992), .Z(n49993) );
  NAND U60249 ( .A(n61042), .B(n49993), .Z(n49994) );
  NANDN U60250 ( .A(n49995), .B(n49994), .Z(n49996) );
  OR U60251 ( .A(n49997), .B(n49996), .Z(n49998) );
  NAND U60252 ( .A(n49999), .B(n49998), .Z(n50000) );
  NAND U60253 ( .A(n50001), .B(n50000), .Z(n50002) );
  AND U60254 ( .A(n50002), .B(n61048), .Z(n50003) );
  NANDN U60255 ( .A(x[8002]), .B(y[8002]), .Z(n61046) );
  AND U60256 ( .A(n50003), .B(n61046), .Z(n50004) );
  OR U60257 ( .A(n50005), .B(n50004), .Z(n50006) );
  NAND U60258 ( .A(n50007), .B(n50006), .Z(n50008) );
  NAND U60259 ( .A(n50009), .B(n50008), .Z(n50010) );
  AND U60260 ( .A(n50010), .B(n50514), .Z(n50011) );
  NANDN U60261 ( .A(x[8006]), .B(y[8006]), .Z(n61052) );
  AND U60262 ( .A(n50011), .B(n61052), .Z(n50015) );
  AND U60263 ( .A(n50013), .B(n50012), .Z(n50014) );
  NANDN U60264 ( .A(n50015), .B(n50014), .Z(n50016) );
  NAND U60265 ( .A(n50017), .B(n50016), .Z(n50018) );
  NAND U60266 ( .A(n50019), .B(n50018), .Z(n50020) );
  AND U60267 ( .A(n50020), .B(n50513), .Z(n50021) );
  NANDN U60268 ( .A(x[8010]), .B(y[8010]), .Z(n61058) );
  AND U60269 ( .A(n50021), .B(n61058), .Z(n50025) );
  AND U60270 ( .A(n50023), .B(n50022), .Z(n50024) );
  NANDN U60271 ( .A(n50025), .B(n50024), .Z(n50026) );
  NAND U60272 ( .A(n50027), .B(n50026), .Z(n50028) );
  NAND U60273 ( .A(n50029), .B(n50028), .Z(n50030) );
  AND U60274 ( .A(n50030), .B(n61064), .Z(n50031) );
  NANDN U60275 ( .A(x[8014]), .B(y[8014]), .Z(n61062) );
  AND U60276 ( .A(n50031), .B(n61062), .Z(n50035) );
  AND U60277 ( .A(n50033), .B(n50032), .Z(n50034) );
  NANDN U60278 ( .A(n50035), .B(n50034), .Z(n50036) );
  NAND U60279 ( .A(n50037), .B(n50036), .Z(n50038) );
  NAND U60280 ( .A(n50039), .B(n50038), .Z(n50040) );
  AND U60281 ( .A(n50040), .B(n61070), .Z(n50041) );
  NANDN U60282 ( .A(x[8018]), .B(y[8018]), .Z(n61067) );
  AND U60283 ( .A(n50041), .B(n61067), .Z(n50045) );
  AND U60284 ( .A(n50043), .B(n50042), .Z(n50044) );
  NANDN U60285 ( .A(n50045), .B(n50044), .Z(n50046) );
  NAND U60286 ( .A(n50047), .B(n50046), .Z(n50048) );
  NAND U60287 ( .A(n50049), .B(n50048), .Z(n50051) );
  IV U60288 ( .A(n50050), .Z(n61074) );
  AND U60289 ( .A(n50051), .B(n61074), .Z(n50052) );
  NANDN U60290 ( .A(x[8022]), .B(y[8022]), .Z(n50510) );
  AND U60291 ( .A(n50052), .B(n50510), .Z(n50056) );
  AND U60292 ( .A(n50054), .B(n50053), .Z(n50055) );
  NANDN U60293 ( .A(n50056), .B(n50055), .Z(n50057) );
  NAND U60294 ( .A(n50058), .B(n50057), .Z(n50059) );
  NAND U60295 ( .A(n50060), .B(n50059), .Z(n50061) );
  AND U60296 ( .A(n50061), .B(n61078), .Z(n50062) );
  NANDN U60297 ( .A(x[8026]), .B(y[8026]), .Z(n50508) );
  AND U60298 ( .A(n50062), .B(n50508), .Z(n50066) );
  AND U60299 ( .A(n50064), .B(n50063), .Z(n50065) );
  NANDN U60300 ( .A(n50066), .B(n50065), .Z(n50067) );
  NAND U60301 ( .A(n50068), .B(n50067), .Z(n50069) );
  NAND U60302 ( .A(n50070), .B(n50069), .Z(n50071) );
  AND U60303 ( .A(n50071), .B(n61084), .Z(n50072) );
  NANDN U60304 ( .A(x[8030]), .B(y[8030]), .Z(n61082) );
  AND U60305 ( .A(n50072), .B(n61082), .Z(n50076) );
  AND U60306 ( .A(n50074), .B(n50073), .Z(n50075) );
  NANDN U60307 ( .A(n50076), .B(n50075), .Z(n50077) );
  NAND U60308 ( .A(n50078), .B(n50077), .Z(n50079) );
  NAND U60309 ( .A(n50080), .B(n50079), .Z(n50081) );
  AND U60310 ( .A(n50081), .B(n50504), .Z(n50082) );
  NANDN U60311 ( .A(x[8034]), .B(y[8034]), .Z(n61088) );
  AND U60312 ( .A(n50082), .B(n61088), .Z(n50086) );
  AND U60313 ( .A(n50084), .B(n50083), .Z(n50085) );
  NANDN U60314 ( .A(n50086), .B(n50085), .Z(n50087) );
  NAND U60315 ( .A(n50088), .B(n50087), .Z(n50089) );
  NAND U60316 ( .A(n50090), .B(n50089), .Z(n50092) );
  IV U60317 ( .A(n50091), .Z(n50502) );
  AND U60318 ( .A(n50092), .B(n50502), .Z(n50093) );
  NANDN U60319 ( .A(x[8038]), .B(y[8038]), .Z(n61092) );
  AND U60320 ( .A(n50093), .B(n61092), .Z(n50097) );
  AND U60321 ( .A(n50095), .B(n50094), .Z(n50096) );
  NANDN U60322 ( .A(n50097), .B(n50096), .Z(n50098) );
  NAND U60323 ( .A(n50099), .B(n50098), .Z(n50100) );
  NAND U60324 ( .A(n50101), .B(n50100), .Z(n50102) );
  AND U60325 ( .A(n50102), .B(n61099), .Z(n50103) );
  NANDN U60326 ( .A(x[8042]), .B(y[8042]), .Z(n61097) );
  AND U60327 ( .A(n50103), .B(n61097), .Z(n50107) );
  AND U60328 ( .A(n50105), .B(n50104), .Z(n50106) );
  NANDN U60329 ( .A(n50107), .B(n50106), .Z(n50108) );
  NAND U60330 ( .A(n50109), .B(n50108), .Z(n50110) );
  NAND U60331 ( .A(n50111), .B(n50110), .Z(n50112) );
  AND U60332 ( .A(n50112), .B(n61103), .Z(n50113) );
  NANDN U60333 ( .A(x[8046]), .B(y[8046]), .Z(n61101) );
  AND U60334 ( .A(n50113), .B(n61101), .Z(n50117) );
  AND U60335 ( .A(n50115), .B(n50114), .Z(n50116) );
  NANDN U60336 ( .A(n50117), .B(n50116), .Z(n50118) );
  NAND U60337 ( .A(n50119), .B(n50118), .Z(n50120) );
  AND U60338 ( .A(n50121), .B(n50120), .Z(n50122) );
  ANDN U60339 ( .B(n61107), .A(n50122), .Z(n50123) );
  NAND U60340 ( .A(n50499), .B(n50123), .Z(n50124) );
  NANDN U60341 ( .A(n50125), .B(n50124), .Z(n50127) );
  AND U60342 ( .A(n50127), .B(n50126), .Z(n50128) );
  NANDN U60343 ( .A(x[8052]), .B(y[8052]), .Z(n61108) );
  NAND U60344 ( .A(n50128), .B(n61108), .Z(n50129) );
  AND U60345 ( .A(n50130), .B(n50129), .Z(n50134) );
  IV U60346 ( .A(n50131), .Z(n61112) );
  AND U60347 ( .A(n50132), .B(n61112), .Z(n50133) );
  NANDN U60348 ( .A(n50134), .B(n50133), .Z(n50135) );
  NANDN U60349 ( .A(n50136), .B(n50135), .Z(n50137) );
  AND U60350 ( .A(n61115), .B(n50137), .Z(n50138) );
  NANDN U60351 ( .A(x[8056]), .B(y[8056]), .Z(n61113) );
  NAND U60352 ( .A(n50138), .B(n61113), .Z(n50139) );
  AND U60353 ( .A(n50140), .B(n50139), .Z(n50141) );
  OR U60354 ( .A(n50142), .B(n50141), .Z(n50143) );
  NAND U60355 ( .A(n50144), .B(n50143), .Z(n50145) );
  NANDN U60356 ( .A(n50146), .B(n50145), .Z(n50147) );
  NAND U60357 ( .A(n50148), .B(n50147), .Z(n50150) );
  IV U60358 ( .A(n50149), .Z(n50492) );
  AND U60359 ( .A(n50150), .B(n50492), .Z(n50151) );
  NANDN U60360 ( .A(x[8062]), .B(y[8062]), .Z(n61119) );
  AND U60361 ( .A(n50151), .B(n61119), .Z(n50155) );
  AND U60362 ( .A(n50153), .B(n50152), .Z(n50154) );
  NANDN U60363 ( .A(n50155), .B(n50154), .Z(n50156) );
  NAND U60364 ( .A(n50157), .B(n50156), .Z(n50158) );
  NAND U60365 ( .A(n50159), .B(n50158), .Z(n50160) );
  AND U60366 ( .A(n50161), .B(n50160), .Z(n50165) );
  AND U60367 ( .A(n50163), .B(n50162), .Z(n50164) );
  NANDN U60368 ( .A(n50165), .B(n50164), .Z(n50166) );
  NAND U60369 ( .A(n50167), .B(n50166), .Z(n50168) );
  NAND U60370 ( .A(n50169), .B(n50168), .Z(n50170) );
  AND U60371 ( .A(n50170), .B(n61127), .Z(n50171) );
  NANDN U60372 ( .A(x[8070]), .B(y[8070]), .Z(n50487) );
  AND U60373 ( .A(n50171), .B(n50487), .Z(n50175) );
  AND U60374 ( .A(n50173), .B(n50172), .Z(n50174) );
  NANDN U60375 ( .A(n50175), .B(n50174), .Z(n50176) );
  NAND U60376 ( .A(n50177), .B(n50176), .Z(n50178) );
  NAND U60377 ( .A(n50179), .B(n50178), .Z(n50180) );
  AND U60378 ( .A(n50180), .B(n61132), .Z(n50181) );
  NANDN U60379 ( .A(x[8074]), .B(y[8074]), .Z(n50486) );
  AND U60380 ( .A(n50181), .B(n50486), .Z(n50182) );
  OR U60381 ( .A(n50183), .B(n50182), .Z(n50184) );
  AND U60382 ( .A(n50185), .B(n50184), .Z(n50186) );
  OR U60383 ( .A(n50187), .B(n50186), .Z(n50188) );
  NAND U60384 ( .A(n50189), .B(n50188), .Z(n50190) );
  NANDN U60385 ( .A(n50191), .B(n50190), .Z(n50192) );
  OR U60386 ( .A(n50193), .B(n50192), .Z(n50194) );
  NAND U60387 ( .A(n50195), .B(n50194), .Z(n50196) );
  NAND U60388 ( .A(n50197), .B(n50196), .Z(n50198) );
  AND U60389 ( .A(n50198), .B(n50481), .Z(n50199) );
  NANDN U60390 ( .A(x[8082]), .B(y[8082]), .Z(n61138) );
  AND U60391 ( .A(n50199), .B(n61138), .Z(n50203) );
  AND U60392 ( .A(n50201), .B(n50200), .Z(n50202) );
  NANDN U60393 ( .A(n50203), .B(n50202), .Z(n50204) );
  NAND U60394 ( .A(n50205), .B(n50204), .Z(n50206) );
  NAND U60395 ( .A(n50207), .B(n50206), .Z(n50208) );
  AND U60396 ( .A(n50208), .B(n61144), .Z(n50209) );
  NANDN U60397 ( .A(x[8086]), .B(y[8086]), .Z(n61141) );
  AND U60398 ( .A(n50209), .B(n61141), .Z(n50213) );
  AND U60399 ( .A(n50211), .B(n50210), .Z(n50212) );
  NANDN U60400 ( .A(n50213), .B(n50212), .Z(n50214) );
  NAND U60401 ( .A(n50215), .B(n50214), .Z(n50216) );
  NAND U60402 ( .A(n50217), .B(n50216), .Z(n50218) );
  AND U60403 ( .A(n50218), .B(n61148), .Z(n50219) );
  NANDN U60404 ( .A(x[8090]), .B(y[8090]), .Z(n50479) );
  AND U60405 ( .A(n50219), .B(n50479), .Z(n50223) );
  AND U60406 ( .A(n50221), .B(n50220), .Z(n50222) );
  NANDN U60407 ( .A(n50223), .B(n50222), .Z(n50224) );
  NAND U60408 ( .A(n50225), .B(n50224), .Z(n50226) );
  NAND U60409 ( .A(n50227), .B(n50226), .Z(n50228) );
  AND U60410 ( .A(n50228), .B(n61152), .Z(n50229) );
  NANDN U60411 ( .A(x[8094]), .B(y[8094]), .Z(n50477) );
  AND U60412 ( .A(n50229), .B(n50477), .Z(n50233) );
  AND U60413 ( .A(n50231), .B(n50230), .Z(n50232) );
  NANDN U60414 ( .A(n50233), .B(n50232), .Z(n50234) );
  NAND U60415 ( .A(n50235), .B(n50234), .Z(n50236) );
  NAND U60416 ( .A(n50237), .B(n50236), .Z(n50238) );
  AND U60417 ( .A(n50238), .B(n61159), .Z(n50239) );
  NANDN U60418 ( .A(x[8098]), .B(y[8098]), .Z(n61156) );
  AND U60419 ( .A(n50239), .B(n61156), .Z(n50243) );
  AND U60420 ( .A(n50241), .B(n50240), .Z(n50242) );
  NANDN U60421 ( .A(n50243), .B(n50242), .Z(n50244) );
  NAND U60422 ( .A(n50245), .B(n50244), .Z(n50246) );
  NAND U60423 ( .A(n50247), .B(n50246), .Z(n50249) );
  IV U60424 ( .A(n50248), .Z(n50473) );
  AND U60425 ( .A(n50249), .B(n50473), .Z(n50250) );
  NANDN U60426 ( .A(x[8102]), .B(y[8102]), .Z(n61162) );
  AND U60427 ( .A(n50250), .B(n61162), .Z(n50254) );
  AND U60428 ( .A(n50252), .B(n50251), .Z(n50253) );
  NANDN U60429 ( .A(n50254), .B(n50253), .Z(n50255) );
  NAND U60430 ( .A(n50256), .B(n50255), .Z(n50257) );
  AND U60431 ( .A(n50258), .B(n50257), .Z(n50259) );
  ANDN U60432 ( .B(n61169), .A(n50259), .Z(n50260) );
  NAND U60433 ( .A(n61166), .B(n50260), .Z(n50261) );
  NANDN U60434 ( .A(n50262), .B(n50261), .Z(n50263) );
  AND U60435 ( .A(n50263), .B(n61171), .Z(n50264) );
  NANDN U60436 ( .A(x[8108]), .B(y[8108]), .Z(n61168) );
  NAND U60437 ( .A(n50264), .B(n61168), .Z(n50265) );
  NAND U60438 ( .A(n50266), .B(n50265), .Z(n50267) );
  AND U60439 ( .A(n50267), .B(n61175), .Z(n50268) );
  NANDN U60440 ( .A(x[8110]), .B(y[8110]), .Z(n61172) );
  AND U60441 ( .A(n50268), .B(n61172), .Z(n50272) );
  AND U60442 ( .A(n50270), .B(n50269), .Z(n50271) );
  NANDN U60443 ( .A(n50272), .B(n50271), .Z(n50273) );
  NAND U60444 ( .A(n50274), .B(n50273), .Z(n50275) );
  NAND U60445 ( .A(n50276), .B(n50275), .Z(n50277) );
  AND U60446 ( .A(n50277), .B(n50470), .Z(n50278) );
  NANDN U60447 ( .A(x[8114]), .B(y[8114]), .Z(n61178) );
  AND U60448 ( .A(n50278), .B(n61178), .Z(n50282) );
  AND U60449 ( .A(n50280), .B(n50279), .Z(n50281) );
  NANDN U60450 ( .A(n50282), .B(n50281), .Z(n50283) );
  NAND U60451 ( .A(n50284), .B(n50283), .Z(n50285) );
  NAND U60452 ( .A(n50286), .B(n50285), .Z(n50288) );
  IV U60453 ( .A(n50287), .Z(n61183) );
  AND U60454 ( .A(n50288), .B(n61183), .Z(n50289) );
  NANDN U60455 ( .A(x[8118]), .B(y[8118]), .Z(n61181) );
  AND U60456 ( .A(n50289), .B(n61181), .Z(n50293) );
  AND U60457 ( .A(n50291), .B(n50290), .Z(n50292) );
  NANDN U60458 ( .A(n50293), .B(n50292), .Z(n50294) );
  NAND U60459 ( .A(n50295), .B(n50294), .Z(n50296) );
  NAND U60460 ( .A(n50297), .B(n50296), .Z(n50298) );
  AND U60461 ( .A(n50298), .B(n50468), .Z(n50299) );
  NANDN U60462 ( .A(x[8122]), .B(y[8122]), .Z(n61188) );
  AND U60463 ( .A(n50299), .B(n61188), .Z(n50303) );
  AND U60464 ( .A(n50301), .B(n50300), .Z(n50302) );
  NANDN U60465 ( .A(n50303), .B(n50302), .Z(n50304) );
  NAND U60466 ( .A(n50305), .B(n50304), .Z(n50306) );
  AND U60467 ( .A(n50307), .B(n50306), .Z(n50308) );
  ANDN U60468 ( .B(n50309), .A(n50308), .Z(n50310) );
  OR U60469 ( .A(n50311), .B(n50310), .Z(n50312) );
  NAND U60470 ( .A(n50313), .B(n50312), .Z(n50314) );
  NAND U60471 ( .A(n50315), .B(n50314), .Z(n50316) );
  AND U60472 ( .A(n50316), .B(n61201), .Z(n50317) );
  NANDN U60473 ( .A(x[8130]), .B(y[8130]), .Z(n61198) );
  AND U60474 ( .A(n50317), .B(n61198), .Z(n50321) );
  AND U60475 ( .A(n50319), .B(n50318), .Z(n50320) );
  NANDN U60476 ( .A(n50321), .B(n50320), .Z(n50322) );
  NAND U60477 ( .A(n50323), .B(n50322), .Z(n50324) );
  NAND U60478 ( .A(n50325), .B(n50324), .Z(n50327) );
  IV U60479 ( .A(n50326), .Z(n61210) );
  AND U60480 ( .A(n50327), .B(n61210), .Z(n50328) );
  NANDN U60481 ( .A(n50465), .B(n50328), .Z(n50329) );
  NAND U60482 ( .A(n50330), .B(n50329), .Z(n50331) );
  NANDN U60483 ( .A(n50463), .B(n50331), .Z(n50332) );
  NANDN U60484 ( .A(x[8136]), .B(y[8136]), .Z(n61212) );
  NANDN U60485 ( .A(n50332), .B(n61212), .Z(n50333) );
  NAND U60486 ( .A(n50334), .B(n50333), .Z(n50335) );
  AND U60487 ( .A(n50335), .B(n61221), .Z(n50336) );
  NANDN U60488 ( .A(x[8138]), .B(y[8138]), .Z(n50464) );
  AND U60489 ( .A(n50336), .B(n50464), .Z(n50340) );
  AND U60490 ( .A(n50338), .B(n50337), .Z(n50339) );
  NANDN U60491 ( .A(n50340), .B(n50339), .Z(n50341) );
  NAND U60492 ( .A(n50342), .B(n50341), .Z(n50343) );
  NAND U60493 ( .A(n50344), .B(n50343), .Z(n50345) );
  AND U60494 ( .A(n50345), .B(n61233), .Z(n50346) );
  NANDN U60495 ( .A(x[8142]), .B(y[8142]), .Z(n61228) );
  AND U60496 ( .A(n50346), .B(n61228), .Z(n50350) );
  AND U60497 ( .A(n50348), .B(n50347), .Z(n50349) );
  NANDN U60498 ( .A(n50350), .B(n50349), .Z(n50351) );
  NAND U60499 ( .A(n50352), .B(n50351), .Z(n50353) );
  NAND U60500 ( .A(n50354), .B(n50353), .Z(n50355) );
  AND U60501 ( .A(n50355), .B(n50461), .Z(n50356) );
  NANDN U60502 ( .A(x[8146]), .B(y[8146]), .Z(n61239) );
  AND U60503 ( .A(n50356), .B(n61239), .Z(n50360) );
  AND U60504 ( .A(n50358), .B(n50357), .Z(n50359) );
  NANDN U60505 ( .A(n50360), .B(n50359), .Z(n50361) );
  NAND U60506 ( .A(n50362), .B(n50361), .Z(n50363) );
  AND U60507 ( .A(n50364), .B(n50363), .Z(n50365) );
  OR U60508 ( .A(n50366), .B(n50365), .Z(n50367) );
  NAND U60509 ( .A(n50368), .B(n50367), .Z(n50369) );
  NANDN U60510 ( .A(n50370), .B(n50369), .Z(n50372) );
  NANDN U60511 ( .A(n50372), .B(n50371), .Z(n50373) );
  AND U60512 ( .A(n50374), .B(n50373), .Z(n50375) );
  OR U60513 ( .A(n50376), .B(n50375), .Z(n50377) );
  NAND U60514 ( .A(n50378), .B(n50377), .Z(n50379) );
  NANDN U60515 ( .A(n50458), .B(n50379), .Z(n50381) );
  NANDN U60516 ( .A(n50381), .B(n50380), .Z(n50382) );
  NAND U60517 ( .A(n50383), .B(n50382), .Z(n50384) );
  AND U60518 ( .A(n50384), .B(n50455), .Z(n50385) );
  NANDN U60519 ( .A(x[8158]), .B(y[8158]), .Z(n50459) );
  AND U60520 ( .A(n50385), .B(n50459), .Z(n50389) );
  AND U60521 ( .A(n50387), .B(n50386), .Z(n50388) );
  NANDN U60522 ( .A(n50389), .B(n50388), .Z(n50390) );
  NAND U60523 ( .A(n50391), .B(n50390), .Z(n50392) );
  NAND U60524 ( .A(n50393), .B(n50392), .Z(n50394) );
  AND U60525 ( .A(n50394), .B(n50452), .Z(n50395) );
  NANDN U60526 ( .A(x[8162]), .B(y[8162]), .Z(n50453) );
  AND U60527 ( .A(n50395), .B(n50453), .Z(n50399) );
  XNOR U60528 ( .A(y[8164]), .B(x[8164]), .Z(n50396) );
  AND U60529 ( .A(n50397), .B(n50396), .Z(n50398) );
  NANDN U60530 ( .A(n50399), .B(n50398), .Z(n50400) );
  NAND U60531 ( .A(n50401), .B(n50400), .Z(n50402) );
  AND U60532 ( .A(n50403), .B(n50402), .Z(n50404) );
  OR U60533 ( .A(n50405), .B(n50404), .Z(n50406) );
  NAND U60534 ( .A(n50407), .B(n50406), .Z(n50408) );
  NANDN U60535 ( .A(n50409), .B(n50408), .Z(n50410) );
  NAND U60536 ( .A(n50411), .B(n50410), .Z(n50412) );
  AND U60537 ( .A(n50412), .B(n61261), .Z(n50413) );
  NANDN U60538 ( .A(x[8170]), .B(y[8170]), .Z(n61259) );
  AND U60539 ( .A(n50413), .B(n61259), .Z(n50414) );
  OR U60540 ( .A(n50415), .B(n50414), .Z(n50416) );
  NAND U60541 ( .A(n50417), .B(n50416), .Z(n50418) );
  NAND U60542 ( .A(n50419), .B(n50418), .Z(n50421) );
  IV U60543 ( .A(n50420), .Z(n61267) );
  AND U60544 ( .A(n50421), .B(n61267), .Z(n50422) );
  NANDN U60545 ( .A(x[8174]), .B(y[8174]), .Z(n61265) );
  AND U60546 ( .A(n50422), .B(n61265), .Z(n50426) );
  AND U60547 ( .A(n50424), .B(n50423), .Z(n50425) );
  NANDN U60548 ( .A(n50426), .B(n50425), .Z(n50427) );
  NAND U60549 ( .A(n50428), .B(n50427), .Z(n50429) );
  NAND U60550 ( .A(n50430), .B(n50429), .Z(n50431) );
  NANDN U60551 ( .A(x[8179]), .B(y[8179]), .Z(n61271) );
  AND U60552 ( .A(n50431), .B(n61271), .Z(n50432) );
  NANDN U60553 ( .A(x[8178]), .B(y[8178]), .Z(n50446) );
  AND U60554 ( .A(n50432), .B(n50446), .Z(n50436) );
  AND U60555 ( .A(n50434), .B(n50433), .Z(n50435) );
  NANDN U60556 ( .A(n50436), .B(n50435), .Z(n50437) );
  NAND U60557 ( .A(n50438), .B(n50437), .Z(n50439) );
  NAND U60558 ( .A(n50440), .B(n50439), .Z(n50441) );
  NAND U60559 ( .A(n50442), .B(n50441), .Z(n61283) );
  NANDN U60560 ( .A(n61283), .B(e), .Z(n5) );
  IV U60561 ( .A(n50455), .Z(n50457) );
  ANDN U60562 ( .B(n50464), .A(n50463), .Z(n61217) );
  NOR U60563 ( .A(n50466), .B(n50465), .Z(n61207) );
  AND U60564 ( .A(n50493), .B(n50492), .Z(n61122) );
  IV U60565 ( .A(n50521), .Z(n61023) );
  ANDN U60566 ( .B(n50549), .A(n50548), .Z(n60939) );
  IV U60567 ( .A(n50562), .Z(n60898) );
  IV U60568 ( .A(n50581), .Z(n50582) );
  AND U60569 ( .A(n50585), .B(n50584), .Z(n60815) );
  AND U60570 ( .A(n50618), .B(n50617), .Z(n60687) );
  ANDN U60571 ( .B(n50620), .A(n50619), .Z(n60677) );
  IV U60572 ( .A(n50624), .Z(n50626) );
  IV U60573 ( .A(n50633), .Z(n50635) );
  IV U60574 ( .A(n50668), .Z(n50669) );
  ANDN U60575 ( .B(n50694), .A(n50693), .Z(n60463) );
  AND U60576 ( .A(n50724), .B(n50723), .Z(n60369) );
  NAND U60577 ( .A(n50735), .B(n50734), .Z(n60323) );
  AND U60578 ( .A(n50796), .B(n50795), .Z(n60114) );
  IV U60579 ( .A(n50820), .Z(n60031) );
  IV U60580 ( .A(n50844), .Z(n50846) );
  IV U60581 ( .A(n50848), .Z(n59948) );
  IV U60582 ( .A(n50853), .Z(n50854) );
  IV U60583 ( .A(n50882), .Z(n50883) );
  IV U60584 ( .A(n50895), .Z(n59792) );
  IV U60585 ( .A(n50915), .Z(n50917) );
  IV U60586 ( .A(n50926), .Z(n59670) );
  ANDN U60587 ( .B(n50962), .A(n50961), .Z(n59534) );
  IV U60588 ( .A(n50973), .Z(n50975) );
  IV U60589 ( .A(n51002), .Z(n51004) );
  AND U60590 ( .A(n51026), .B(n51025), .Z(n59295) );
  AND U60591 ( .A(n51047), .B(n51046), .Z(n59205) );
  AND U60592 ( .A(n51053), .B(n51052), .Z(n59170) );
  ANDN U60593 ( .B(n51055), .A(n51054), .Z(n59148) );
  AND U60594 ( .A(n51061), .B(n51060), .Z(n59101) );
  AND U60595 ( .A(n51090), .B(n51089), .Z(n59006) );
  ANDN U60596 ( .B(n51132), .A(n51131), .Z(n58831) );
  AND U60597 ( .A(n51186), .B(n51185), .Z(n58642) );
  AND U60598 ( .A(n51227), .B(n51226), .Z(n58475) );
  IV U60599 ( .A(n51263), .Z(n51264) );
  AND U60600 ( .A(n51267), .B(n51266), .Z(n58314) );
  AND U60601 ( .A(n51269), .B(n51268), .Z(n58288) );
  AND U60602 ( .A(n51272), .B(n51271), .Z(n58265) );
  IV U60603 ( .A(n51301), .Z(n58177) );
  AND U60604 ( .A(n51325), .B(n51324), .Z(n58091) );
  IV U60605 ( .A(n51332), .Z(n58059) );
  IV U60606 ( .A(n51368), .Z(n57893) );
  AND U60607 ( .A(n51384), .B(n51383), .Z(n57831) );
  IV U60608 ( .A(n51388), .Z(n57816) );
  IV U60609 ( .A(n51391), .Z(n51392) );
  IV U60610 ( .A(n51408), .Z(n57736) );
  IV U60611 ( .A(n51429), .Z(n57668) );
  AND U60612 ( .A(n51458), .B(n51457), .Z(n57565) );
  IV U60613 ( .A(n51470), .Z(n57508) );
  IV U60614 ( .A(n51475), .Z(n57496) );
  IV U60615 ( .A(n51479), .Z(n57483) );
  IV U60616 ( .A(n51506), .Z(n57348) );
  IV U60617 ( .A(n51519), .Z(n57268) );
  IV U60618 ( .A(n51552), .Z(n51553) );
  IV U60619 ( .A(n51561), .Z(n57050) );
  AND U60620 ( .A(n51572), .B(n51571), .Z(n57011) );
  IV U60621 ( .A(n51587), .Z(n56910) );
  IV U60622 ( .A(n51607), .Z(n56753) );
  IV U60623 ( .A(n51617), .Z(n51618) );
  IV U60624 ( .A(n51632), .Z(n56651) );
  AND U60625 ( .A(n51644), .B(n51643), .Z(n56617) );
  IV U60626 ( .A(n51655), .Z(n56583) );
  IV U60627 ( .A(n51672), .Z(n56498) );
  AND U60628 ( .A(n51677), .B(n51676), .Z(n56478) );
  IV U60629 ( .A(n51689), .Z(n56387) );
  AND U60630 ( .A(n51696), .B(n51695), .Z(n56377) );
  IV U60631 ( .A(n51708), .Z(n56335) );
  IV U60632 ( .A(n51733), .Z(n56269) );
  IV U60633 ( .A(n51749), .Z(n56222) );
  IV U60634 ( .A(n51760), .Z(n56183) );
  IV U60635 ( .A(n51763), .Z(n56170) );
  IV U60636 ( .A(n51766), .Z(n56158) );
  IV U60637 ( .A(n51776), .Z(n56118) );
  IV U60638 ( .A(n51827), .Z(n55930) );
  IV U60639 ( .A(n51842), .Z(n55891) );
  IV U60640 ( .A(n51879), .Z(n55761) );
  IV U60641 ( .A(n51906), .Z(n55572) );
  IV U60642 ( .A(n51919), .Z(n55545) );
  IV U60643 ( .A(n51940), .Z(n55475) );
  XNOR U60644 ( .A(x[3192]), .B(y[3192]), .Z(n55447) );
  IV U60645 ( .A(n51966), .Z(n55382) );
  IV U60646 ( .A(n51976), .Z(n55289) );
  IV U60647 ( .A(n52005), .Z(n55070) );
  IV U60648 ( .A(n52022), .Z(n54926) );
  IV U60649 ( .A(n52028), .Z(n54835) );
  IV U60650 ( .A(n52036), .Z(n54829) );
  IV U60651 ( .A(n52074), .Z(n54658) );
  IV U60652 ( .A(n52102), .Z(n54493) );
  ANDN U60653 ( .B(n52150), .A(n52149), .Z(n54222) );
  IV U60654 ( .A(n52158), .Z(n54130) );
  IV U60655 ( .A(n52176), .Z(n54085) );
  IV U60656 ( .A(n52214), .Z(n53867) );
  IV U60657 ( .A(n52231), .Z(n53824) );
  ANDN U60658 ( .B(n52237), .A(n52236), .Z(n53778) );
  IV U60659 ( .A(n52289), .Z(n53437) );
  IV U60660 ( .A(n52319), .Z(n53253) );
  IV U60661 ( .A(n52323), .Z(n53240) );
  IV U60662 ( .A(n52328), .Z(n53209) );
  IV U60663 ( .A(n52345), .Z(n53162) );
  IV U60664 ( .A(n52371), .Z(n52893) );
  IV U60665 ( .A(n52382), .Z(n52875) );
  IV U60666 ( .A(n52389), .Z(n52869) );
  IV U60667 ( .A(n52407), .Z(n52744) );
  NANDN U60668 ( .A(n52528), .B(n52527), .Z(n52529) );
  AND U60669 ( .A(n52530), .B(n52529), .Z(n52531) );
  OR U60670 ( .A(n52532), .B(n52531), .Z(n52533) );
  NAND U60671 ( .A(n52534), .B(n52533), .Z(n52535) );
  NANDN U60672 ( .A(n52536), .B(n52535), .Z(n52537) );
  NAND U60673 ( .A(n52538), .B(n52537), .Z(n52539) );
  NANDN U60674 ( .A(n52540), .B(n52539), .Z(n52541) );
  AND U60675 ( .A(n52542), .B(n52541), .Z(n52543) );
  OR U60676 ( .A(n52544), .B(n52543), .Z(n52545) );
  NAND U60677 ( .A(n52546), .B(n52545), .Z(n52547) );
  NANDN U60678 ( .A(n52548), .B(n52547), .Z(n52549) );
  NAND U60679 ( .A(n52550), .B(n52549), .Z(n52551) );
  NANDN U60680 ( .A(n52552), .B(n52551), .Z(n52553) );
  AND U60681 ( .A(n52554), .B(n52553), .Z(n52555) );
  OR U60682 ( .A(n52556), .B(n52555), .Z(n52557) );
  NAND U60683 ( .A(n52558), .B(n52557), .Z(n52559) );
  NANDN U60684 ( .A(n52560), .B(n52559), .Z(n52561) );
  NAND U60685 ( .A(n52562), .B(n52561), .Z(n52563) );
  NANDN U60686 ( .A(n52564), .B(n52563), .Z(n52565) );
  AND U60687 ( .A(n52566), .B(n52565), .Z(n52567) );
  NANDN U60688 ( .A(n52611), .B(n52610), .Z(n52612) );
  AND U60689 ( .A(n52613), .B(n52612), .Z(n52614) );
  OR U60690 ( .A(n52615), .B(n52614), .Z(n52616) );
  NAND U60691 ( .A(n52617), .B(n52616), .Z(n52618) );
  NANDN U60692 ( .A(n52619), .B(n52618), .Z(n52620) );
  NAND U60693 ( .A(n52621), .B(n52620), .Z(n52622) );
  NANDN U60694 ( .A(n52623), .B(n52622), .Z(n52624) );
  AND U60695 ( .A(n52625), .B(n52624), .Z(n52626) );
  OR U60696 ( .A(n52627), .B(n52626), .Z(n52628) );
  NAND U60697 ( .A(n52629), .B(n52628), .Z(n52630) );
  NANDN U60698 ( .A(n52631), .B(n52630), .Z(n52632) );
  NAND U60699 ( .A(n52633), .B(n52632), .Z(n52634) );
  NANDN U60700 ( .A(n52635), .B(n52634), .Z(n52636) );
  AND U60701 ( .A(n52637), .B(n52636), .Z(n52638) );
  OR U60702 ( .A(n52639), .B(n52638), .Z(n52640) );
  NAND U60703 ( .A(n52641), .B(n52640), .Z(n52642) );
  NANDN U60704 ( .A(n52643), .B(n52642), .Z(n52644) );
  NAND U60705 ( .A(n52645), .B(n52644), .Z(n52646) );
  NANDN U60706 ( .A(n52647), .B(n52646), .Z(n52648) );
  AND U60707 ( .A(n52649), .B(n52648), .Z(n52650) );
  NAND U60708 ( .A(n52688), .B(n52687), .Z(n52689) );
  NANDN U60709 ( .A(n52690), .B(n52689), .Z(n52691) );
  NAND U60710 ( .A(n52692), .B(n52691), .Z(n52693) );
  NANDN U60711 ( .A(n52694), .B(n52693), .Z(n52695) );
  AND U60712 ( .A(n52696), .B(n52695), .Z(n52698) );
  NANDN U60713 ( .A(n52698), .B(n52697), .Z(n52699) );
  NAND U60714 ( .A(n52700), .B(n52699), .Z(n52701) );
  NANDN U60715 ( .A(n52702), .B(n52701), .Z(n52703) );
  NAND U60716 ( .A(n52704), .B(n52703), .Z(n52705) );
  NANDN U60717 ( .A(n52706), .B(n52705), .Z(n52707) );
  AND U60718 ( .A(n52708), .B(n52707), .Z(n52709) );
  OR U60719 ( .A(n52710), .B(n52709), .Z(n52711) );
  NAND U60720 ( .A(n52712), .B(n52711), .Z(n52713) );
  NANDN U60721 ( .A(n52714), .B(n52713), .Z(n52715) );
  NAND U60722 ( .A(n52716), .B(n52715), .Z(n52717) );
  NANDN U60723 ( .A(n52718), .B(n52717), .Z(n52719) );
  AND U60724 ( .A(n52720), .B(n52719), .Z(n52721) );
  OR U60725 ( .A(n52722), .B(n52721), .Z(n52723) );
  NAND U60726 ( .A(n52724), .B(n52723), .Z(n52725) );
  NANDN U60727 ( .A(n52726), .B(n52725), .Z(n52727) );
  NANDN U60728 ( .A(n52766), .B(n52765), .Z(n52767) );
  NANDN U60729 ( .A(n52768), .B(n52767), .Z(n52769) );
  AND U60730 ( .A(n52770), .B(n52769), .Z(n52771) );
  OR U60731 ( .A(n52772), .B(n52771), .Z(n52773) );
  NAND U60732 ( .A(n52774), .B(n52773), .Z(n52775) );
  NANDN U60733 ( .A(n52776), .B(n52775), .Z(n52777) );
  NAND U60734 ( .A(n52778), .B(n52777), .Z(n52779) );
  NANDN U60735 ( .A(n52780), .B(n52779), .Z(n52781) );
  AND U60736 ( .A(n52782), .B(n52781), .Z(n52783) );
  OR U60737 ( .A(n52784), .B(n52783), .Z(n52785) );
  NAND U60738 ( .A(n52786), .B(n52785), .Z(n52787) );
  NANDN U60739 ( .A(n52788), .B(n52787), .Z(n52789) );
  NAND U60740 ( .A(n52790), .B(n52789), .Z(n52791) );
  NANDN U60741 ( .A(n52792), .B(n52791), .Z(n52793) );
  AND U60742 ( .A(n52794), .B(n52793), .Z(n52795) );
  OR U60743 ( .A(n52796), .B(n52795), .Z(n52797) );
  NAND U60744 ( .A(n52798), .B(n52797), .Z(n52799) );
  NANDN U60745 ( .A(n52800), .B(n52799), .Z(n52801) );
  NANDN U60746 ( .A(n52802), .B(n52801), .Z(n52803) );
  NAND U60747 ( .A(n52804), .B(n52803), .Z(n52807) );
  IV U60748 ( .A(n52805), .Z(n52806) );
  AND U60749 ( .A(n52807), .B(n52806), .Z(n52809) );
  NANDN U60750 ( .A(n52809), .B(n52808), .Z(n52810) );
  NAND U60751 ( .A(n52811), .B(n52810), .Z(n52812) );
  NANDN U60752 ( .A(n52813), .B(n52812), .Z(n52814) );
  NAND U60753 ( .A(n52815), .B(n52814), .Z(n52816) );
  NANDN U60754 ( .A(n52817), .B(n52816), .Z(n52818) );
  AND U60755 ( .A(n52819), .B(n52818), .Z(n52820) );
  OR U60756 ( .A(n52821), .B(n52820), .Z(n52822) );
  NAND U60757 ( .A(n52823), .B(n52822), .Z(n52824) );
  NANDN U60758 ( .A(n52825), .B(n52824), .Z(n52826) );
  NAND U60759 ( .A(n52827), .B(n52826), .Z(n52828) );
  NANDN U60760 ( .A(n52829), .B(n52828), .Z(n52830) );
  AND U60761 ( .A(n52831), .B(n52830), .Z(n52832) );
  OR U60762 ( .A(n52833), .B(n52832), .Z(n52834) );
  NAND U60763 ( .A(n52835), .B(n52834), .Z(n52836) );
  NANDN U60764 ( .A(n52837), .B(n52836), .Z(n52838) );
  NAND U60765 ( .A(n52839), .B(n52838), .Z(n52840) );
  NANDN U60766 ( .A(n52841), .B(n52840), .Z(n52842) );
  AND U60767 ( .A(n52843), .B(n52842), .Z(n52844) );
  OR U60768 ( .A(n52845), .B(n52844), .Z(n52846) );
  IV U60769 ( .A(n52901), .Z(n52902) );
  IV U60770 ( .A(n52945), .Z(n52946) );
  IV U60771 ( .A(n53072), .Z(n53073) );
  NANDN U60772 ( .A(n53122), .B(n53121), .Z(n53123) );
  NAND U60773 ( .A(n53124), .B(n53123), .Z(n53125) );
  NANDN U60774 ( .A(n53126), .B(n53125), .Z(n53127) );
  AND U60775 ( .A(n53128), .B(n53127), .Z(n53129) );
  OR U60776 ( .A(n53130), .B(n53129), .Z(n53131) );
  NAND U60777 ( .A(n53132), .B(n53131), .Z(n53133) );
  NANDN U60778 ( .A(n53134), .B(n53133), .Z(n53135) );
  NAND U60779 ( .A(n53136), .B(n53135), .Z(n53137) );
  NANDN U60780 ( .A(n53138), .B(n53137), .Z(n53139) );
  AND U60781 ( .A(n53140), .B(n53139), .Z(n53141) );
  OR U60782 ( .A(n53142), .B(n53141), .Z(n53143) );
  NAND U60783 ( .A(n53144), .B(n53143), .Z(n53145) );
  NANDN U60784 ( .A(n53146), .B(n53145), .Z(n53148) );
  NAND U60785 ( .A(n53148), .B(n53147), .Z(n53149) );
  NANDN U60786 ( .A(n53150), .B(n53149), .Z(n53151) );
  AND U60787 ( .A(n53152), .B(n53151), .Z(n53153) );
  OR U60788 ( .A(n53154), .B(n53153), .Z(n53155) );
  NAND U60789 ( .A(n53156), .B(n53155), .Z(n53157) );
  NANDN U60790 ( .A(n53158), .B(n53157), .Z(n53159) );
  NAND U60791 ( .A(n53160), .B(n53159), .Z(n53161) );
  IV U60792 ( .A(n53169), .Z(n53170) );
  IV U60793 ( .A(n53172), .Z(n53173) );
  IV U60794 ( .A(n53178), .Z(n53179) );
  IV U60795 ( .A(n53272), .Z(n53273) );
  NANDN U60796 ( .A(n53364), .B(n53363), .Z(n53365) );
  NANDN U60797 ( .A(n53366), .B(n53365), .Z(n53367) );
  AND U60798 ( .A(n53368), .B(n53367), .Z(n53369) );
  OR U60799 ( .A(n53370), .B(n53369), .Z(n53371) );
  NAND U60800 ( .A(n53372), .B(n53371), .Z(n53373) );
  NANDN U60801 ( .A(n53374), .B(n53373), .Z(n53375) );
  NAND U60802 ( .A(n53376), .B(n53375), .Z(n53377) );
  NANDN U60803 ( .A(n53378), .B(n53377), .Z(n53379) );
  AND U60804 ( .A(n53380), .B(n53379), .Z(n53381) );
  OR U60805 ( .A(n53382), .B(n53381), .Z(n53383) );
  NAND U60806 ( .A(n53384), .B(n53383), .Z(n53385) );
  NANDN U60807 ( .A(n53386), .B(n53385), .Z(n53387) );
  NAND U60808 ( .A(n53388), .B(n53387), .Z(n53389) );
  NANDN U60809 ( .A(n53390), .B(n53389), .Z(n53391) );
  AND U60810 ( .A(n53392), .B(n53391), .Z(n53393) );
  OR U60811 ( .A(n53394), .B(n53393), .Z(n53395) );
  NAND U60812 ( .A(n53396), .B(n53395), .Z(n53397) );
  NANDN U60813 ( .A(n53398), .B(n53397), .Z(n53399) );
  NAND U60814 ( .A(n53400), .B(n53399), .Z(n53401) );
  NANDN U60815 ( .A(n53402), .B(n53401), .Z(n53403) );
  IV U60816 ( .A(n53430), .Z(n53431) );
  IV U60817 ( .A(n53438), .Z(n53439) );
  IV U60818 ( .A(n53449), .Z(n53450) );
  IV U60819 ( .A(n53480), .Z(n53481) );
  IV U60820 ( .A(n53483), .Z(n53484) );
  NANDN U60821 ( .A(n53635), .B(n53634), .Z(n53636) );
  NAND U60822 ( .A(n53637), .B(n53636), .Z(n53638) );
  NANDN U60823 ( .A(n53639), .B(n53638), .Z(n53640) );
  AND U60824 ( .A(n53641), .B(n53640), .Z(n53643) );
  OR U60825 ( .A(n53643), .B(n53642), .Z(n53644) );
  AND U60826 ( .A(n53645), .B(n53644), .Z(n53646) );
  OR U60827 ( .A(n53647), .B(n53646), .Z(n53648) );
  AND U60828 ( .A(n53649), .B(n53648), .Z(n53651) );
  NANDN U60829 ( .A(n53651), .B(n53650), .Z(n53652) );
  NAND U60830 ( .A(n53653), .B(n53652), .Z(n53654) );
  NANDN U60831 ( .A(n53655), .B(n53654), .Z(n53656) );
  NAND U60832 ( .A(n53657), .B(n53656), .Z(n53658) );
  NANDN U60833 ( .A(n53659), .B(n53658), .Z(n53660) );
  AND U60834 ( .A(n53661), .B(n53660), .Z(n53662) );
  OR U60835 ( .A(n53663), .B(n53662), .Z(n53664) );
  NAND U60836 ( .A(n53665), .B(n53664), .Z(n53666) );
  NANDN U60837 ( .A(n53667), .B(n53666), .Z(n53668) );
  NAND U60838 ( .A(n53669), .B(n53668), .Z(n53670) );
  NANDN U60839 ( .A(n53671), .B(n53670), .Z(n53672) );
  AND U60840 ( .A(n53673), .B(n53672), .Z(n53674) );
  IV U60841 ( .A(n53691), .Z(n53692) );
  OR U60842 ( .A(n53752), .B(n53751), .Z(n53753) );
  NAND U60843 ( .A(n53754), .B(n53753), .Z(n53755) );
  NANDN U60844 ( .A(n53756), .B(n53755), .Z(n53757) );
  NAND U60845 ( .A(n53758), .B(n53757), .Z(n53759) );
  NANDN U60846 ( .A(n53760), .B(n53759), .Z(n53761) );
  AND U60847 ( .A(n53762), .B(n53761), .Z(n53763) );
  OR U60848 ( .A(n53764), .B(n53763), .Z(n53765) );
  NAND U60849 ( .A(n53766), .B(n53765), .Z(n53767) );
  NANDN U60850 ( .A(n53768), .B(n53767), .Z(n53769) );
  NAND U60851 ( .A(n53770), .B(n53769), .Z(n53771) );
  NANDN U60852 ( .A(n53772), .B(n53771), .Z(n53773) );
  AND U60853 ( .A(n53774), .B(n53773), .Z(n53775) );
  OR U60854 ( .A(n53776), .B(n53775), .Z(n53777) );
  AND U60855 ( .A(n53778), .B(n53777), .Z(n53782) );
  AND U60856 ( .A(n53780), .B(n53779), .Z(n53781) );
  NANDN U60857 ( .A(n53782), .B(n53781), .Z(n53784) );
  ANDN U60858 ( .B(n53784), .A(n53783), .Z(n53786) );
  NAND U60859 ( .A(n53786), .B(n53785), .Z(n53787) );
  NANDN U60860 ( .A(n53788), .B(n53787), .Z(n53789) );
  IV U60861 ( .A(n53829), .Z(n53830) );
  IV U60862 ( .A(n53913), .Z(n53914) );
  IV U60863 ( .A(n53916), .Z(n53917) );
  IV U60864 ( .A(n54094), .Z(n54095) );
  IV U60865 ( .A(n54097), .Z(n54098) );
  IV U60866 ( .A(n54114), .Z(n54115) );
  IV U60867 ( .A(n54196), .Z(n54197) );
  NANDN U60868 ( .A(n54212), .B(n54211), .Z(n54213) );
  NANDN U60869 ( .A(n54214), .B(n54213), .Z(n54215) );
  AND U60870 ( .A(n54216), .B(n54215), .Z(n54218) );
  OR U60871 ( .A(n54218), .B(n54217), .Z(n54219) );
  AND U60872 ( .A(n54220), .B(n54219), .Z(n54221) );
  ANDN U60873 ( .B(n54222), .A(n54221), .Z(n54224) );
  NANDN U60874 ( .A(n54224), .B(n54223), .Z(n54225) );
  AND U60875 ( .A(n54226), .B(n54225), .Z(n54228) );
  NANDN U60876 ( .A(n54228), .B(n54227), .Z(n54229) );
  NAND U60877 ( .A(n54230), .B(n54229), .Z(n54231) );
  NANDN U60878 ( .A(n54232), .B(n54231), .Z(n54234) );
  ANDN U60879 ( .B(n54234), .A(n54233), .Z(n54236) );
  NANDN U60880 ( .A(n54236), .B(n54235), .Z(n54237) );
  NANDN U60881 ( .A(n54238), .B(n54237), .Z(n54240) );
  AND U60882 ( .A(n54240), .B(n54239), .Z(n54242) );
  NANDN U60883 ( .A(n54242), .B(n54241), .Z(n54243) );
  AND U60884 ( .A(n54244), .B(n54243), .Z(n54246) );
  NANDN U60885 ( .A(n54246), .B(n54245), .Z(n54247) );
  AND U60886 ( .A(n54248), .B(n54247), .Z(n54249) );
  IV U60887 ( .A(n54302), .Z(n54303) );
  IV U60888 ( .A(n54349), .Z(n54350) );
  IV U60889 ( .A(n54369), .Z(n54370) );
  IV U60890 ( .A(n54372), .Z(n54373) );
  IV U60891 ( .A(n54397), .Z(n54398) );
  IV U60892 ( .A(n54421), .Z(n54422) );
  AND U60893 ( .A(n54469), .B(n54468), .Z(n54470) );
  IV U60894 ( .A(n54548), .Z(n54549) );
  IV U60895 ( .A(n54566), .Z(n54567) );
  IV U60896 ( .A(n54597), .Z(n54598) );
  IV U60897 ( .A(n54600), .Z(n54601) );
  IV U60898 ( .A(n54617), .Z(n54618) );
  IV U60899 ( .A(n54641), .Z(n54642) );
  IV U60900 ( .A(n54817), .Z(n54818) );
  IV U60901 ( .A(n54820), .Z(n54821) );
  IV U60902 ( .A(n54836), .Z(n54837) );
  IV U60903 ( .A(n54868), .Z(n54869) );
  IV U60904 ( .A(n54884), .Z(n54885) );
  OR U60905 ( .A(n54886), .B(n54885), .Z(n54887) );
  AND U60906 ( .A(n54888), .B(n54887), .Z(n54889) );
  OR U60907 ( .A(n54890), .B(n54889), .Z(n54891) );
  NAND U60908 ( .A(n54892), .B(n54891), .Z(n54893) );
  NANDN U60909 ( .A(n54894), .B(n54893), .Z(n54895) );
  NANDN U60910 ( .A(n54896), .B(n54895), .Z(n54897) );
  AND U60911 ( .A(n54898), .B(n54897), .Z(n54899) );
  OR U60912 ( .A(n54900), .B(n54899), .Z(n54901) );
  NAND U60913 ( .A(n54902), .B(n54901), .Z(n54903) );
  NANDN U60914 ( .A(n54904), .B(n54903), .Z(n54905) );
  NANDN U60915 ( .A(n54906), .B(n54905), .Z(n54907) );
  AND U60916 ( .A(n54908), .B(n54907), .Z(n54909) );
  OR U60917 ( .A(n54910), .B(n54909), .Z(n54911) );
  NAND U60918 ( .A(n54912), .B(n54911), .Z(n54913) );
  NANDN U60919 ( .A(n54914), .B(n54913), .Z(n54915) );
  NANDN U60920 ( .A(n54916), .B(n54915), .Z(n54917) );
  AND U60921 ( .A(n54918), .B(n54917), .Z(n54919) );
  OR U60922 ( .A(n54920), .B(n54919), .Z(n54921) );
  NAND U60923 ( .A(n54922), .B(n54921), .Z(n54923) );
  NANDN U60924 ( .A(n54924), .B(n54923), .Z(n54925) );
  NAND U60925 ( .A(n54959), .B(n54958), .Z(n54962) );
  IV U60926 ( .A(n54960), .Z(n54961) );
  OR U60927 ( .A(n54962), .B(n54961), .Z(n54963) );
  NANDN U60928 ( .A(n54964), .B(n54963), .Z(n54965) );
  AND U60929 ( .A(n54966), .B(n54965), .Z(n54967) );
  OR U60930 ( .A(n54968), .B(n54967), .Z(n54969) );
  NAND U60931 ( .A(n54970), .B(n54969), .Z(n54971) );
  NANDN U60932 ( .A(n54972), .B(n54971), .Z(n54973) );
  NANDN U60933 ( .A(n54974), .B(n54973), .Z(n54975) );
  NAND U60934 ( .A(n54976), .B(n54975), .Z(n54977) );
  AND U60935 ( .A(n54978), .B(n54977), .Z(n54979) );
  NANDN U60936 ( .A(n54980), .B(n54979), .Z(n54981) );
  NAND U60937 ( .A(n54982), .B(n54981), .Z(n54983) );
  NANDN U60938 ( .A(n54984), .B(n54983), .Z(n54985) );
  OR U60939 ( .A(n54986), .B(n54985), .Z(n54987) );
  AND U60940 ( .A(n54988), .B(n54987), .Z(n54989) );
  OR U60941 ( .A(n54990), .B(n54989), .Z(n54991) );
  NAND U60942 ( .A(n54992), .B(n54991), .Z(n54993) );
  NANDN U60943 ( .A(n54994), .B(n54993), .Z(n54995) );
  NANDN U60944 ( .A(n54996), .B(n54995), .Z(n54997) );
  AND U60945 ( .A(n54998), .B(n54997), .Z(n55000) );
  IV U60946 ( .A(n55080), .Z(n55081) );
  IV U60947 ( .A(n55098), .Z(n55099) );
  IV U60948 ( .A(n55166), .Z(n55167) );
  IV U60949 ( .A(n55169), .Z(n55170) );
  AND U60950 ( .A(n55176), .B(n55175), .Z(n55177) );
  IV U60951 ( .A(n55212), .Z(n55213) );
  OR U60952 ( .A(n55229), .B(n55228), .Z(n55230) );
  NAND U60953 ( .A(n55231), .B(n55230), .Z(n55232) );
  NANDN U60954 ( .A(n55233), .B(n55232), .Z(n55234) );
  NANDN U60955 ( .A(n55235), .B(n55234), .Z(n55236) );
  AND U60956 ( .A(n55237), .B(n55236), .Z(n55238) );
  OR U60957 ( .A(n55239), .B(n55238), .Z(n55240) );
  NAND U60958 ( .A(n55241), .B(n55240), .Z(n55242) );
  NANDN U60959 ( .A(n55243), .B(n55242), .Z(n55244) );
  NANDN U60960 ( .A(n55245), .B(n55244), .Z(n55246) );
  AND U60961 ( .A(n55247), .B(n55246), .Z(n55248) );
  OR U60962 ( .A(n55249), .B(n55248), .Z(n55250) );
  NAND U60963 ( .A(n55251), .B(n55250), .Z(n55252) );
  NANDN U60964 ( .A(n55253), .B(n55252), .Z(n55254) );
  NANDN U60965 ( .A(n55255), .B(n55254), .Z(n55256) );
  AND U60966 ( .A(n55257), .B(n55256), .Z(n55258) );
  OR U60967 ( .A(n55259), .B(n55258), .Z(n55260) );
  NAND U60968 ( .A(n55261), .B(n55260), .Z(n55262) );
  NANDN U60969 ( .A(n55263), .B(n55262), .Z(n55264) );
  NANDN U60970 ( .A(n55265), .B(n55264), .Z(n55266) );
  AND U60971 ( .A(n55267), .B(n55266), .Z(n55270) );
  IV U60972 ( .A(n55268), .Z(n55269) );
  AND U60973 ( .A(n55322), .B(n55321), .Z(n55323) );
  OR U60974 ( .A(n55324), .B(n55323), .Z(n55325) );
  NAND U60975 ( .A(n55326), .B(n55325), .Z(n55327) );
  NANDN U60976 ( .A(n55328), .B(n55327), .Z(n55329) );
  NANDN U60977 ( .A(n55330), .B(n55329), .Z(n55331) );
  AND U60978 ( .A(n55332), .B(n55331), .Z(n55333) );
  OR U60979 ( .A(n55334), .B(n55333), .Z(n55335) );
  NAND U60980 ( .A(n55336), .B(n55335), .Z(n55337) );
  NANDN U60981 ( .A(n55338), .B(n55337), .Z(n55339) );
  NANDN U60982 ( .A(n55340), .B(n55339), .Z(n55341) );
  AND U60983 ( .A(n55342), .B(n55341), .Z(n55343) );
  OR U60984 ( .A(n55344), .B(n55343), .Z(n55345) );
  NAND U60985 ( .A(n55346), .B(n55345), .Z(n55347) );
  NANDN U60986 ( .A(n55348), .B(n55347), .Z(n55349) );
  NANDN U60987 ( .A(n55350), .B(n55349), .Z(n55351) );
  AND U60988 ( .A(n55352), .B(n55351), .Z(n55353) );
  OR U60989 ( .A(n55354), .B(n55353), .Z(n55355) );
  NAND U60990 ( .A(n55356), .B(n55355), .Z(n55357) );
  NANDN U60991 ( .A(n55358), .B(n55357), .Z(n55359) );
  NANDN U60992 ( .A(n55360), .B(n55359), .Z(n55361) );
  IV U60993 ( .A(n55383), .Z(n55384) );
  IV U60994 ( .A(n55476), .Z(n55477) );
  IV U60995 ( .A(n55488), .Z(n55489) );
  IV U60996 ( .A(n55580), .Z(n55581) );
  IV U60997 ( .A(n55600), .Z(n55601) );
  IV U60998 ( .A(n55612), .Z(n55613) );
  IV U60999 ( .A(n55615), .Z(n55616) );
  IV U61000 ( .A(n55628), .Z(n55629) );
  NANDN U61001 ( .A(n55664), .B(n55663), .Z(n55665) );
  NANDN U61002 ( .A(n55666), .B(n55665), .Z(n55667) );
  AND U61003 ( .A(n55668), .B(n55667), .Z(n55669) );
  OR U61004 ( .A(n55670), .B(n55669), .Z(n55671) );
  NAND U61005 ( .A(n55672), .B(n55671), .Z(n55673) );
  NANDN U61006 ( .A(n55674), .B(n55673), .Z(n55675) );
  NANDN U61007 ( .A(n55676), .B(n55675), .Z(n55677) );
  AND U61008 ( .A(n55678), .B(n55677), .Z(n55679) );
  OR U61009 ( .A(n55680), .B(n55679), .Z(n55681) );
  NAND U61010 ( .A(n55682), .B(n55681), .Z(n55683) );
  NANDN U61011 ( .A(n55684), .B(n55683), .Z(n55685) );
  NANDN U61012 ( .A(n55686), .B(n55685), .Z(n55687) );
  AND U61013 ( .A(n55688), .B(n55687), .Z(n55689) );
  OR U61014 ( .A(n55690), .B(n55689), .Z(n55691) );
  NAND U61015 ( .A(n55692), .B(n55691), .Z(n55693) );
  NANDN U61016 ( .A(n55694), .B(n55693), .Z(n55695) );
  NANDN U61017 ( .A(n55696), .B(n55695), .Z(n55697) );
  AND U61018 ( .A(n55698), .B(n55697), .Z(n55699) );
  OR U61019 ( .A(n55700), .B(n55699), .Z(n55701) );
  NAND U61020 ( .A(n55702), .B(n55701), .Z(n55703) );
  NANDN U61021 ( .A(n55704), .B(n55703), .Z(n55705) );
  NANDN U61022 ( .A(n55706), .B(n55705), .Z(n55707) );
  AND U61023 ( .A(n55708), .B(n55707), .Z(n55709) );
  OR U61024 ( .A(n55710), .B(n55709), .Z(n55711) );
  NAND U61025 ( .A(n55712), .B(n55711), .Z(n55713) );
  NANDN U61026 ( .A(n55714), .B(n55713), .Z(n55718) );
  AND U61027 ( .A(n55716), .B(n55715), .Z(n55717) );
  NAND U61028 ( .A(n55718), .B(n55717), .Z(n55719) );
  AND U61029 ( .A(n55720), .B(n55719), .Z(n55721) );
  OR U61030 ( .A(n55722), .B(n55721), .Z(n55723) );
  NAND U61031 ( .A(n55724), .B(n55723), .Z(n55725) );
  NANDN U61032 ( .A(n55726), .B(n55725), .Z(n55727) );
  NANDN U61033 ( .A(n55728), .B(n55727), .Z(n55729) );
  AND U61034 ( .A(n55730), .B(n55729), .Z(n55731) );
  OR U61035 ( .A(n55732), .B(n55731), .Z(n55733) );
  NAND U61036 ( .A(n55734), .B(n55733), .Z(n55735) );
  NANDN U61037 ( .A(n55736), .B(n55735), .Z(n55737) );
  NANDN U61038 ( .A(n55738), .B(n55737), .Z(n55739) );
  AND U61039 ( .A(n55740), .B(n55739), .Z(n55741) );
  OR U61040 ( .A(n55742), .B(n55741), .Z(n55743) );
  IV U61041 ( .A(n55815), .Z(n55816) );
  IV U61042 ( .A(n55860), .Z(n55861) );
  IV U61043 ( .A(n55877), .Z(n55878) );
  IV U61044 ( .A(n55892), .Z(n55893) );
  IV U61045 ( .A(n55899), .Z(n55900) );
  IV U61046 ( .A(n55931), .Z(n55932) );
  AND U61047 ( .A(n55975), .B(n55974), .Z(n55976) );
  IV U61048 ( .A(n56061), .Z(n56062) );
  IV U61049 ( .A(n56072), .Z(n56073) );
  IV U61050 ( .A(n56081), .Z(n56082) );
  IV U61051 ( .A(n56094), .Z(n56095) );
  IV U61052 ( .A(n56171), .Z(n56172) );
  IV U61053 ( .A(n56207), .Z(n56208) );
  IV U61054 ( .A(n56249), .Z(n56250) );
  IV U61055 ( .A(n56259), .Z(n56260) );
  IV U61056 ( .A(n56271), .Z(n56272) );
  IV U61057 ( .A(n56304), .Z(n56305) );
  IV U61058 ( .A(n56424), .Z(n56425) );
  OR U61059 ( .A(n56446), .B(n56445), .Z(n56447) );
  NAND U61060 ( .A(n56448), .B(n56447), .Z(n56449) );
  NANDN U61061 ( .A(n56450), .B(n56449), .Z(n56451) );
  AND U61062 ( .A(n56452), .B(n56451), .Z(n56454) );
  NANDN U61063 ( .A(n56454), .B(n56453), .Z(n56455) );
  NANDN U61064 ( .A(n56456), .B(n56455), .Z(n56457) );
  AND U61065 ( .A(n56458), .B(n56457), .Z(n56459) );
  OR U61066 ( .A(n56460), .B(n56459), .Z(n56461) );
  NAND U61067 ( .A(n56462), .B(n56461), .Z(n56463) );
  NANDN U61068 ( .A(n56464), .B(n56463), .Z(n56465) );
  NAND U61069 ( .A(n56466), .B(n56465), .Z(n56468) );
  AND U61070 ( .A(n56468), .B(n56467), .Z(n56469) );
  NAND U61071 ( .A(n56470), .B(n56469), .Z(n56471) );
  NANDN U61072 ( .A(n56472), .B(n56471), .Z(n56473) );
  AND U61073 ( .A(n56474), .B(n56473), .Z(n56475) );
  OR U61074 ( .A(n56476), .B(n56475), .Z(n56477) );
  AND U61075 ( .A(n56478), .B(n56477), .Z(n56479) );
  OR U61076 ( .A(n56480), .B(n56479), .Z(n56481) );
  NAND U61077 ( .A(n56482), .B(n56481), .Z(n56483) );
  IV U61078 ( .A(n56526), .Z(n56527) );
  IV U61079 ( .A(n56537), .Z(n56538) );
  IV U61080 ( .A(n56584), .Z(n56585) );
  IV U61081 ( .A(n56591), .Z(n56592) );
  IV U61082 ( .A(n56594), .Z(n56595) );
  IV U61083 ( .A(n56606), .Z(n56607) );
  IV U61084 ( .A(n56618), .Z(n56619) );
  IV U61085 ( .A(n56695), .Z(n56696) );
  IV U61086 ( .A(n56710), .Z(n56711) );
  AND U61087 ( .A(n56766), .B(n56765), .Z(n56770) );
  AND U61088 ( .A(n56768), .B(n56767), .Z(n56769) );
  NANDN U61089 ( .A(n56770), .B(n56769), .Z(n56771) );
  NAND U61090 ( .A(n56772), .B(n56771), .Z(n56773) );
  AND U61091 ( .A(n56774), .B(n56773), .Z(n56776) );
  AND U61092 ( .A(n56776), .B(n56775), .Z(n56778) );
  OR U61093 ( .A(n56778), .B(n56777), .Z(n56779) );
  AND U61094 ( .A(n56780), .B(n56779), .Z(n56781) );
  OR U61095 ( .A(n56782), .B(n56781), .Z(n56783) );
  NAND U61096 ( .A(n56784), .B(n56783), .Z(n56785) );
  NANDN U61097 ( .A(n56786), .B(n56785), .Z(n56787) );
  AND U61098 ( .A(n56788), .B(n56787), .Z(n56790) );
  AND U61099 ( .A(n56790), .B(n56789), .Z(n56792) );
  OR U61100 ( .A(n56792), .B(n56791), .Z(n56793) );
  AND U61101 ( .A(n56794), .B(n56793), .Z(n56795) );
  OR U61102 ( .A(n56796), .B(n56795), .Z(n56797) );
  NAND U61103 ( .A(n56798), .B(n56797), .Z(n56799) );
  NANDN U61104 ( .A(n56800), .B(n56799), .Z(n56801) );
  AND U61105 ( .A(n56802), .B(n56801), .Z(n56803) );
  OR U61106 ( .A(n56804), .B(n56803), .Z(n56805) );
  IV U61107 ( .A(n56870), .Z(n56871) );
  IV U61108 ( .A(n56873), .Z(n56874) );
  IV U61109 ( .A(n56886), .Z(n56887) );
  IV U61110 ( .A(n56894), .Z(n56895) );
  IV U61111 ( .A(n56922), .Z(n56923) );
  IV U61112 ( .A(n56956), .Z(n56957) );
  IV U61113 ( .A(n57051), .Z(n57052) );
  IV U61114 ( .A(n57053), .Z(n57054) );
  IV U61115 ( .A(n57081), .Z(n57082) );
  IV U61116 ( .A(n57108), .Z(n57109) );
  IV U61117 ( .A(n57139), .Z(n57140) );
  IV U61118 ( .A(n57168), .Z(n57169) );
  IV U61119 ( .A(n57171), .Z(n57172) );
  IV U61120 ( .A(n57185), .Z(n57186) );
  IV U61121 ( .A(n57225), .Z(n57226) );
  IV U61122 ( .A(n57281), .Z(n57282) );
  IV U61123 ( .A(n57299), .Z(n57300) );
  IV U61124 ( .A(n57349), .Z(n57350) );
  IV U61125 ( .A(n57434), .Z(n57435) );
  IV U61126 ( .A(n57467), .Z(n57468) );
  IV U61127 ( .A(n57553), .Z(n57554) );
  IV U61128 ( .A(n57572), .Z(n57573) );
  IV U61129 ( .A(n57582), .Z(n57583) );
  ANDN U61130 ( .B(n57643), .A(n57642), .Z(n57644) );
  IV U61131 ( .A(n57646), .Z(n57647) );
  IV U61132 ( .A(n57654), .Z(n57655) );
  IV U61133 ( .A(n57669), .Z(n57670) );
  IV U61134 ( .A(n57709), .Z(n57710) );
  IV U61135 ( .A(n57722), .Z(n57723) );
  IV U61136 ( .A(n57725), .Z(n57727) );
  IV U61137 ( .A(n57747), .Z(n57748) );
  IV U61138 ( .A(n57766), .Z(n57767) );
  IV U61139 ( .A(n57817), .Z(n57818) );
  IV U61140 ( .A(n57942), .Z(n57943) );
  IV U61141 ( .A(n57944), .Z(n57945) );
  IV U61142 ( .A(n57996), .Z(n57998) );
  IV U61143 ( .A(n58074), .Z(n58075) );
  IV U61144 ( .A(n58107), .Z(n58108) );
  IV U61145 ( .A(n58131), .Z(n58132) );
  IV U61146 ( .A(n58234), .Z(n58235) );
  IV U61147 ( .A(n58237), .Z(n58238) );
  AND U61148 ( .A(n58283), .B(n58282), .Z(n58286) );
  IV U61149 ( .A(n58284), .Z(n58285) );
  OR U61150 ( .A(n58286), .B(n58285), .Z(n58287) );
  NAND U61151 ( .A(n58288), .B(n58287), .Z(n58289) );
  AND U61152 ( .A(n58290), .B(n58289), .Z(n58294) );
  AND U61153 ( .A(n58292), .B(n58291), .Z(n58293) );
  NANDN U61154 ( .A(n58294), .B(n58293), .Z(n58295) );
  NANDN U61155 ( .A(n58296), .B(n58295), .Z(n58297) );
  AND U61156 ( .A(n58298), .B(n58297), .Z(n58300) );
  AND U61157 ( .A(n58300), .B(n58299), .Z(n58302) );
  OR U61158 ( .A(n58302), .B(n58301), .Z(n58303) );
  AND U61159 ( .A(n58304), .B(n58303), .Z(n58306) );
  AND U61160 ( .A(n58306), .B(n58305), .Z(n58308) );
  OR U61161 ( .A(n58308), .B(n58307), .Z(n58309) );
  AND U61162 ( .A(n58310), .B(n58309), .Z(n58311) );
  OR U61163 ( .A(n58312), .B(n58311), .Z(n58313) );
  NAND U61164 ( .A(n58314), .B(n58313), .Z(n58315) );
  NANDN U61165 ( .A(n58316), .B(n58315), .Z(n58317) );
  AND U61166 ( .A(n58318), .B(n58317), .Z(n58320) );
  IV U61167 ( .A(n58417), .Z(n58418) );
  IV U61168 ( .A(n58420), .Z(n58421) );
  IV U61169 ( .A(n58436), .Z(n58437) );
  IV U61170 ( .A(n58477), .Z(n58478) );
  IV U61171 ( .A(n58504), .Z(n58505) );
  IV U61172 ( .A(n58522), .Z(n58523) );
  IV U61173 ( .A(n58525), .Z(n58526) );
  IV U61174 ( .A(n58575), .Z(n58576) );
  IV U61175 ( .A(n58578), .Z(n58579) );
  IV U61176 ( .A(n58644), .Z(n58645) );
  AND U61177 ( .A(n58674), .B(n58673), .Z(n58675) );
  NOR U61178 ( .A(n58724), .B(n58723), .Z(n58725) );
  IV U61179 ( .A(n58766), .Z(n58767) );
  IV U61180 ( .A(n58768), .Z(n58769) );
  IV U61181 ( .A(n58866), .Z(n58867) );
  IV U61182 ( .A(n58973), .Z(n58974) );
  IV U61183 ( .A(n58975), .Z(n58976) );
  IV U61184 ( .A(n59014), .Z(n59015) );
  IV U61185 ( .A(n59030), .Z(n59031) );
  IV U61186 ( .A(n59041), .Z(n59042) );
  IV U61187 ( .A(n59060), .Z(n59061) );
  IV U61188 ( .A(n59082), .Z(n59083) );
  IV U61189 ( .A(n59103), .Z(n59104) );
  AND U61190 ( .A(n59136), .B(n59135), .Z(n59138) );
  AND U61191 ( .A(n59138), .B(n59137), .Z(n59140) );
  OR U61192 ( .A(n59140), .B(n59139), .Z(n59141) );
  AND U61193 ( .A(n59142), .B(n59141), .Z(n59144) );
  AND U61194 ( .A(n59144), .B(n59143), .Z(n59146) );
  NANDN U61195 ( .A(n59146), .B(n59145), .Z(n59147) );
  NAND U61196 ( .A(n59148), .B(n59147), .Z(n59149) );
  NAND U61197 ( .A(n59150), .B(n59149), .Z(n59152) );
  AND U61198 ( .A(n59152), .B(n59151), .Z(n59153) );
  NAND U61199 ( .A(n59154), .B(n59153), .Z(n59155) );
  NAND U61200 ( .A(n59156), .B(n59155), .Z(n59157) );
  AND U61201 ( .A(n59158), .B(n59157), .Z(n59160) );
  AND U61202 ( .A(n59160), .B(n59159), .Z(n59162) );
  OR U61203 ( .A(n59162), .B(n59161), .Z(n59163) );
  AND U61204 ( .A(n59164), .B(n59163), .Z(n59166) );
  AND U61205 ( .A(n59166), .B(n59165), .Z(n59167) );
  OR U61206 ( .A(n59168), .B(n59167), .Z(n59169) );
  NAND U61207 ( .A(n59170), .B(n59169), .Z(n59171) );
  IV U61208 ( .A(n59173), .Z(n59174) );
  IV U61209 ( .A(n59207), .Z(n59208) );
  IV U61210 ( .A(n59384), .Z(n59385) );
  IV U61211 ( .A(n59500), .Z(n59501) );
  IV U61212 ( .A(n59549), .Z(n59550) );
  IV U61213 ( .A(n59684), .Z(n59685) );
  IV U61214 ( .A(n59700), .Z(n59701) );
  IV U61215 ( .A(n59732), .Z(n59733) );
  IV U61216 ( .A(n59818), .Z(n59819) );
  IV U61217 ( .A(n59821), .Z(n59823) );
  IV U61218 ( .A(n59933), .Z(n59934) );
  IV U61219 ( .A(n60133), .Z(n60134) );
  IV U61220 ( .A(n60258), .Z(n60259) );
  IV U61221 ( .A(n60294), .Z(n60295) );
  IV U61222 ( .A(n60480), .Z(n60481) );
  IV U61223 ( .A(n60588), .Z(n60589) );
  IV U61224 ( .A(n60590), .Z(n60592) );
  IV U61225 ( .A(n60642), .Z(n60643) );
  AND U61226 ( .A(n60673), .B(n60672), .Z(n60675) );
  NANDN U61227 ( .A(n60675), .B(n60674), .Z(n60676) );
  NAND U61228 ( .A(n60677), .B(n60676), .Z(n60678) );
  NAND U61229 ( .A(n60679), .B(n60678), .Z(n60680) );
  AND U61230 ( .A(n60681), .B(n60680), .Z(n60683) );
  AND U61231 ( .A(n60683), .B(n60682), .Z(n60685) );
  NANDN U61232 ( .A(n60685), .B(n60684), .Z(n60686) );
  NAND U61233 ( .A(n60687), .B(n60686), .Z(n60688) );
  NANDN U61234 ( .A(n60689), .B(n60688), .Z(n60690) );
  AND U61235 ( .A(n60691), .B(n60690), .Z(n60693) );
  NAND U61236 ( .A(n60693), .B(n60692), .Z(n60694) );
  NAND U61237 ( .A(n60695), .B(n60694), .Z(n60697) );
  ANDN U61238 ( .B(n60697), .A(n60696), .Z(n60699) );
  NAND U61239 ( .A(n60699), .B(n60698), .Z(n60700) );
  NAND U61240 ( .A(n60701), .B(n60700), .Z(n60702) );
  AND U61241 ( .A(n60703), .B(n60702), .Z(n60705) );
  NAND U61242 ( .A(n60705), .B(n60704), .Z(n60706) );
  NAND U61243 ( .A(n60707), .B(n60706), .Z(n60709) );
  IV U61244 ( .A(n60781), .Z(n60782) );
  AND U61245 ( .A(n60783), .B(n60782), .Z(n60787) );
  NANDN U61246 ( .A(n60787), .B(n60786), .Z(n60788) );
  NANDN U61247 ( .A(n60789), .B(n60788), .Z(n60790) );
  AND U61248 ( .A(n60791), .B(n60790), .Z(n60793) );
  NAND U61249 ( .A(n60793), .B(n60792), .Z(n60794) );
  NAND U61250 ( .A(n60795), .B(n60794), .Z(n60797) );
  ANDN U61251 ( .B(n60797), .A(n60796), .Z(n60799) );
  NAND U61252 ( .A(n60799), .B(n60798), .Z(n60800) );
  NANDN U61253 ( .A(n60801), .B(n60800), .Z(n60802) );
  AND U61254 ( .A(n60803), .B(n60802), .Z(n60805) );
  NAND U61255 ( .A(n60805), .B(n60804), .Z(n60806) );
  NAND U61256 ( .A(n60807), .B(n60806), .Z(n60809) );
  ANDN U61257 ( .B(n60809), .A(n60808), .Z(n60811) );
  AND U61258 ( .A(n60811), .B(n60810), .Z(n60813) );
  NANDN U61259 ( .A(n60813), .B(n60812), .Z(n60814) );
  NAND U61260 ( .A(n60815), .B(n60814), .Z(n60816) );
  NAND U61261 ( .A(n60817), .B(n60816), .Z(n60818) );
  AND U61262 ( .A(n60819), .B(n60818), .Z(n60821) );
  AND U61263 ( .A(n60821), .B(n60820), .Z(n60822) );
  IV U61264 ( .A(n60838), .Z(n60839) );
  IV U61265 ( .A(n60852), .Z(n60853) );
  IV U61266 ( .A(n60867), .Z(n60868) );
  IV U61267 ( .A(n60882), .Z(n60883) );
  IV U61268 ( .A(n60924), .Z(n60925) );
  IV U61269 ( .A(n61038), .Z(n61039) );
  IV U61270 ( .A(n61109), .Z(n61110) );
  AND U61271 ( .A(n61201), .B(n61200), .Z(n61203) );
  AND U61272 ( .A(n61203), .B(n61202), .Z(n61205) );
  NANDN U61273 ( .A(n61205), .B(n61204), .Z(n61206) );
  NAND U61274 ( .A(n61207), .B(n61206), .Z(n61208) );
  NAND U61275 ( .A(n61209), .B(n61208), .Z(n61211) );
  AND U61276 ( .A(n61211), .B(n61210), .Z(n61213) );
  AND U61277 ( .A(n61213), .B(n61212), .Z(n61215) );
  NANDN U61278 ( .A(n61215), .B(n61214), .Z(n61216) );
  NAND U61279 ( .A(n61217), .B(n61216), .Z(n61218) );
  NANDN U61280 ( .A(n61219), .B(n61218), .Z(n61220) );
  AND U61281 ( .A(n61221), .B(n61220), .Z(n61223) );
  NAND U61282 ( .A(n61223), .B(n61222), .Z(n61224) );
  NAND U61283 ( .A(n61225), .B(n61224), .Z(n61227) );
  ANDN U61284 ( .B(n61227), .A(n61226), .Z(n61229) );
  NAND U61285 ( .A(n61229), .B(n61228), .Z(n61230) );
  NANDN U61286 ( .A(n61231), .B(n61230), .Z(n61232) );
  AND U61287 ( .A(n61233), .B(n61232), .Z(n61235) );
  NAND U61288 ( .A(n61235), .B(n61234), .Z(n61236) );
endmodule

