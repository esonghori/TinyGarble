
module stackMachine_N16 ( clk, rst, x, opcode, o );
  input [15:0] x;
  input [2:0] opcode;
  output [15:0] o;
  input clk, rst;
  wire   \stack[7][15] , \stack[7][14] , \stack[7][13] , \stack[7][12] ,
         \stack[7][11] , \stack[7][10] , \stack[7][9] , \stack[7][8] ,
         \stack[7][7] , \stack[7][6] , \stack[7][5] , \stack[7][4] ,
         \stack[7][3] , \stack[7][2] , \stack[7][1] , \stack[7][0] ,
         \stack[6][15] , \stack[6][14] , \stack[6][13] , \stack[6][12] ,
         \stack[6][11] , \stack[6][10] , \stack[6][9] , \stack[6][8] ,
         \stack[6][7] , \stack[6][6] , \stack[6][5] , \stack[6][4] ,
         \stack[6][3] , \stack[6][2] , \stack[6][1] , \stack[6][0] ,
         \stack[5][15] , \stack[5][14] , \stack[5][13] , \stack[5][12] ,
         \stack[5][11] , \stack[5][10] , \stack[5][9] , \stack[5][8] ,
         \stack[5][7] , \stack[5][6] , \stack[5][5] , \stack[5][4] ,
         \stack[5][3] , \stack[5][2] , \stack[5][1] , \stack[5][0] ,
         \stack[4][15] , \stack[4][14] , \stack[4][13] , \stack[4][12] ,
         \stack[4][11] , \stack[4][10] , \stack[4][9] , \stack[4][8] ,
         \stack[4][7] , \stack[4][6] , \stack[4][5] , \stack[4][4] ,
         \stack[4][3] , \stack[4][2] , \stack[4][1] , \stack[4][0] ,
         \stack[3][15] , \stack[3][14] , \stack[3][13] , \stack[3][12] ,
         \stack[3][11] , \stack[3][10] , \stack[3][9] , \stack[3][8] ,
         \stack[3][7] , \stack[3][6] , \stack[3][5] , \stack[3][4] ,
         \stack[3][3] , \stack[3][2] , \stack[3][1] , \stack[3][0] ,
         \stack[2][15] , \stack[2][14] , \stack[2][13] , \stack[2][12] ,
         \stack[2][11] , \stack[2][10] , \stack[2][9] , \stack[2][8] ,
         \stack[2][7] , \stack[2][6] , \stack[2][5] , \stack[2][4] ,
         \stack[2][3] , \stack[2][2] , \stack[2][1] , \stack[2][0] ,
         \stack[1][15] , \stack[1][14] , \stack[1][13] , \stack[1][12] ,
         \stack[1][11] , \stack[1][10] , \stack[1][9] , \stack[1][8] ,
         \stack[1][7] , \stack[1][6] , \stack[1][5] , \stack[1][4] ,
         \stack[1][3] , \stack[1][2] , \stack[1][1] , \stack[1][0] ,
         \C3/DATA5_0 , \C3/DATA5_1 , \C3/DATA5_2 , \C3/DATA5_3 , \C3/DATA5_4 ,
         \C3/DATA5_5 , \C3/DATA5_6 , \C3/DATA5_7 , \C3/DATA5_8 , \C3/DATA5_9 ,
         \C3/DATA5_10 , \C3/DATA5_11 , \C3/DATA5_12 , \C3/DATA5_13 ,
         \C3/DATA5_14 , \C3/DATA5_15 , n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, \C1/Z_0 , \U1/RSOP_16/C3/Z_15 , \U1/RSOP_16/C3/Z_14 ,
         \U1/RSOP_16/C3/Z_13 , \U1/RSOP_16/C3/Z_12 , \U1/RSOP_16/C3/Z_11 ,
         \U1/RSOP_16/C3/Z_10 , \U1/RSOP_16/C3/Z_9 , \U1/RSOP_16/C3/Z_8 ,
         \U1/RSOP_16/C3/Z_7 , \U1/RSOP_16/C3/Z_6 , \U1/RSOP_16/C3/Z_5 ,
         \U1/RSOP_16/C3/Z_4 , \U1/RSOP_16/C3/Z_3 , \U1/RSOP_16/C3/Z_2 ,
         \U1/RSOP_16/C3/Z_1 , \U1/RSOP_16/C3/Z_0 , \U1/RSOP_16/C2/Z_15 ,
         \U1/RSOP_16/C2/Z_14 , \U1/RSOP_16/C2/Z_13 , \U1/RSOP_16/C2/Z_12 ,
         \U1/RSOP_16/C2/Z_11 , \U1/RSOP_16/C2/Z_10 , \U1/RSOP_16/C2/Z_9 ,
         \U1/RSOP_16/C2/Z_8 , \U1/RSOP_16/C2/Z_7 , \U1/RSOP_16/C2/Z_6 ,
         \U1/RSOP_16/C2/Z_5 , \U1/RSOP_16/C2/Z_4 , \U1/RSOP_16/C2/Z_3 ,
         \U1/RSOP_16/C2/Z_2 , \U1/RSOP_16/C2/Z_1 , \U1/RSOP_16/C2/Z_0 ,
         \DP_OP_25_64_3291/n169 , \DP_OP_25_64_3291/n168 ,
         \DP_OP_25_64_3291/n167 , \DP_OP_25_64_3291/n166 ,
         \DP_OP_25_64_3291/n165 , \DP_OP_25_64_3291/n164 ,
         \DP_OP_25_64_3291/n163 , \DP_OP_25_64_3291/n162 ,
         \DP_OP_25_64_3291/n161 , \DP_OP_25_64_3291/n160 ,
         \DP_OP_25_64_3291/n159 , \DP_OP_25_64_3291/n158 ,
         \DP_OP_25_64_3291/n157 , \DP_OP_25_64_3291/n156 ,
         \DP_OP_25_64_3291/n155 , \DP_OP_25_64_3291/n154 ,
         \DP_OP_25_64_3291/n149 , \DP_OP_25_64_3291/n148 ,
         \DP_OP_25_64_3291/n147 , \DP_OP_25_64_3291/n146 ,
         \DP_OP_25_64_3291/n145 , \DP_OP_25_64_3291/n144 ,
         \DP_OP_25_64_3291/n143 , \DP_OP_25_64_3291/n142 ,
         \DP_OP_25_64_3291/n141 , \DP_OP_25_64_3291/n140 ,
         \DP_OP_25_64_3291/n139 , \DP_OP_25_64_3291/n138 ,
         \DP_OP_25_64_3291/n137 , \DP_OP_25_64_3291/n136 ,
         \DP_OP_25_64_3291/n135 , \DP_OP_25_64_3291/n134 ,
         \DP_OP_25_64_3291/n133 , \DP_OP_25_64_3291/n132 ,
         \DP_OP_25_64_3291/n131 , \DP_OP_25_64_3291/n130 ,
         \DP_OP_25_64_3291/n129 , \DP_OP_25_64_3291/n128 ,
         \DP_OP_25_64_3291/n127 , \DP_OP_25_64_3291/n126 ,
         \DP_OP_25_64_3291/n125 , \DP_OP_25_64_3291/n124 ,
         \DP_OP_25_64_3291/n123 , \DP_OP_25_64_3291/n122 ,
         \DP_OP_25_64_3291/n121 , \DP_OP_25_64_3291/n120 ,
         \DP_OP_25_64_3291/n119 , \DP_OP_25_64_3291/n117 ,
         \DP_OP_25_64_3291/n116 , \DP_OP_25_64_3291/n110 ,
         \DP_OP_25_64_3291/n109 , \DP_OP_25_64_3291/n103 ,
         \DP_OP_25_64_3291/n102 , \DP_OP_25_64_3291/n96 ,
         \DP_OP_25_64_3291/n95 , \DP_OP_25_64_3291/n89 ,
         \DP_OP_25_64_3291/n88 , \DP_OP_25_64_3291/n82 ,
         \DP_OP_25_64_3291/n81 , \DP_OP_25_64_3291/n70 ,
         \DP_OP_25_64_3291/n69 , \DP_OP_25_64_3291/n57 ,
         \DP_OP_25_64_3291/n56 , \DP_OP_25_64_3291/n50 ,
         \DP_OP_25_64_3291/n49 , \DP_OP_25_64_3291/n43 ,
         \DP_OP_25_64_3291/n42 , \DP_OP_25_64_3291/n36 ,
         \DP_OP_25_64_3291/n35 , \DP_OP_25_64_3291/n29 ,
         \DP_OP_25_64_3291/n28 , \DP_OP_25_64_3291/n22 ,
         \DP_OP_25_64_3291/n21 , \DP_OP_25_64_3291/n15 ,
         \DP_OP_25_64_3291/n14 , \DP_OP_25_64_3291/n8 , \DP_OP_25_64_3291/n5 ,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
         n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
         n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
         n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
         n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
         n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
         n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
         n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
         n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
         n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
         n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
         n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
         n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
         n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
         n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
         n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
         n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
         n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
         n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
         n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
         n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
         n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
         n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
         n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
         n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
         n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
         n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
         n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
         n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
         n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
         n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
         n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
         n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
         n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
         n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
         n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
         n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
         n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
         n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
         n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
         n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
         n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
         n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
         n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
         n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
         n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
         n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
         n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
         n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
         n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
         n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
         n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
         n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
         n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
         n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968,
         n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
         n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
         n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998,
         n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008,
         n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018,
         n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028,
         n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
         n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
         n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058,
         n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068,
         n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078,
         n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088,
         n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098,
         n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108,
         n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
         n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
         n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
         n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
         n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
         n2159, n2160;

  DFF \stack_reg[0][0]  ( .D(n680), .CLK(clk), .RST(rst), .Q(o[0]) );
  DFF \stack_reg[1][0]  ( .D(n679), .CLK(clk), .RST(rst), .Q(\stack[1][0] ) );
  DFF \stack_reg[0][1]  ( .D(n678), .CLK(clk), .RST(rst), .Q(o[1]) );
  DFF \stack_reg[1][1]  ( .D(n677), .CLK(clk), .RST(rst), .Q(\stack[1][1] ) );
  DFF \stack_reg[2][1]  ( .D(n676), .CLK(clk), .RST(rst), .Q(\stack[2][1] ) );
  DFF \stack_reg[3][1]  ( .D(n675), .CLK(clk), .RST(rst), .Q(\stack[3][1] ) );
  DFF \stack_reg[4][1]  ( .D(n674), .CLK(clk), .RST(rst), .Q(\stack[4][1] ) );
  DFF \stack_reg[5][1]  ( .D(n673), .CLK(clk), .RST(rst), .Q(\stack[5][1] ) );
  DFF \stack_reg[6][1]  ( .D(n672), .CLK(clk), .RST(rst), .Q(\stack[6][1] ) );
  DFF \stack_reg[7][1]  ( .D(n671), .CLK(clk), .RST(rst), .Q(\stack[7][1] ) );
  DFF \stack_reg[0][2]  ( .D(n670), .CLK(clk), .RST(rst), .Q(o[2]) );
  DFF \stack_reg[1][2]  ( .D(n669), .CLK(clk), .RST(rst), .Q(\stack[1][2] ) );
  DFF \stack_reg[2][2]  ( .D(n668), .CLK(clk), .RST(rst), .Q(\stack[2][2] ) );
  DFF \stack_reg[3][2]  ( .D(n667), .CLK(clk), .RST(rst), .Q(\stack[3][2] ) );
  DFF \stack_reg[4][2]  ( .D(n666), .CLK(clk), .RST(rst), .Q(\stack[4][2] ) );
  DFF \stack_reg[5][2]  ( .D(n665), .CLK(clk), .RST(rst), .Q(\stack[5][2] ) );
  DFF \stack_reg[6][2]  ( .D(n664), .CLK(clk), .RST(rst), .Q(\stack[6][2] ) );
  DFF \stack_reg[7][2]  ( .D(n663), .CLK(clk), .RST(rst), .Q(\stack[7][2] ) );
  DFF \stack_reg[0][3]  ( .D(n662), .CLK(clk), .RST(rst), .Q(o[3]) );
  DFF \stack_reg[1][3]  ( .D(n661), .CLK(clk), .RST(rst), .Q(\stack[1][3] ) );
  DFF \stack_reg[2][3]  ( .D(n660), .CLK(clk), .RST(rst), .Q(\stack[2][3] ) );
  DFF \stack_reg[3][3]  ( .D(n659), .CLK(clk), .RST(rst), .Q(\stack[3][3] ) );
  DFF \stack_reg[4][3]  ( .D(n658), .CLK(clk), .RST(rst), .Q(\stack[4][3] ) );
  DFF \stack_reg[5][3]  ( .D(n657), .CLK(clk), .RST(rst), .Q(\stack[5][3] ) );
  DFF \stack_reg[6][3]  ( .D(n656), .CLK(clk), .RST(rst), .Q(\stack[6][3] ) );
  DFF \stack_reg[7][3]  ( .D(n655), .CLK(clk), .RST(rst), .Q(\stack[7][3] ) );
  DFF \stack_reg[0][4]  ( .D(n654), .CLK(clk), .RST(rst), .Q(o[4]) );
  DFF \stack_reg[1][4]  ( .D(n653), .CLK(clk), .RST(rst), .Q(\stack[1][4] ) );
  DFF \stack_reg[2][4]  ( .D(n652), .CLK(clk), .RST(rst), .Q(\stack[2][4] ) );
  DFF \stack_reg[3][4]  ( .D(n651), .CLK(clk), .RST(rst), .Q(\stack[3][4] ) );
  DFF \stack_reg[4][4]  ( .D(n650), .CLK(clk), .RST(rst), .Q(\stack[4][4] ) );
  DFF \stack_reg[5][4]  ( .D(n649), .CLK(clk), .RST(rst), .Q(\stack[5][4] ) );
  DFF \stack_reg[6][4]  ( .D(n648), .CLK(clk), .RST(rst), .Q(\stack[6][4] ) );
  DFF \stack_reg[7][4]  ( .D(n647), .CLK(clk), .RST(rst), .Q(\stack[7][4] ) );
  DFF \stack_reg[0][5]  ( .D(n646), .CLK(clk), .RST(rst), .Q(o[5]) );
  DFF \stack_reg[1][5]  ( .D(n645), .CLK(clk), .RST(rst), .Q(\stack[1][5] ) );
  DFF \stack_reg[2][5]  ( .D(n644), .CLK(clk), .RST(rst), .Q(\stack[2][5] ) );
  DFF \stack_reg[3][5]  ( .D(n643), .CLK(clk), .RST(rst), .Q(\stack[3][5] ) );
  DFF \stack_reg[4][5]  ( .D(n642), .CLK(clk), .RST(rst), .Q(\stack[4][5] ) );
  DFF \stack_reg[5][5]  ( .D(n641), .CLK(clk), .RST(rst), .Q(\stack[5][5] ) );
  DFF \stack_reg[6][5]  ( .D(n640), .CLK(clk), .RST(rst), .Q(\stack[6][5] ) );
  DFF \stack_reg[7][5]  ( .D(n639), .CLK(clk), .RST(rst), .Q(\stack[7][5] ) );
  DFF \stack_reg[0][6]  ( .D(n638), .CLK(clk), .RST(rst), .Q(o[6]) );
  DFF \stack_reg[1][6]  ( .D(n637), .CLK(clk), .RST(rst), .Q(\stack[1][6] ) );
  DFF \stack_reg[2][6]  ( .D(n636), .CLK(clk), .RST(rst), .Q(\stack[2][6] ) );
  DFF \stack_reg[3][6]  ( .D(n635), .CLK(clk), .RST(rst), .Q(\stack[3][6] ) );
  DFF \stack_reg[4][6]  ( .D(n634), .CLK(clk), .RST(rst), .Q(\stack[4][6] ) );
  DFF \stack_reg[5][6]  ( .D(n633), .CLK(clk), .RST(rst), .Q(\stack[5][6] ) );
  DFF \stack_reg[6][6]  ( .D(n632), .CLK(clk), .RST(rst), .Q(\stack[6][6] ) );
  DFF \stack_reg[7][6]  ( .D(n631), .CLK(clk), .RST(rst), .Q(\stack[7][6] ) );
  DFF \stack_reg[0][7]  ( .D(n630), .CLK(clk), .RST(rst), .Q(o[7]) );
  DFF \stack_reg[1][7]  ( .D(n629), .CLK(clk), .RST(rst), .Q(\stack[1][7] ) );
  DFF \stack_reg[2][7]  ( .D(n628), .CLK(clk), .RST(rst), .Q(\stack[2][7] ) );
  DFF \stack_reg[3][7]  ( .D(n627), .CLK(clk), .RST(rst), .Q(\stack[3][7] ) );
  DFF \stack_reg[4][7]  ( .D(n626), .CLK(clk), .RST(rst), .Q(\stack[4][7] ) );
  DFF \stack_reg[5][7]  ( .D(n625), .CLK(clk), .RST(rst), .Q(\stack[5][7] ) );
  DFF \stack_reg[6][7]  ( .D(n624), .CLK(clk), .RST(rst), .Q(\stack[6][7] ) );
  DFF \stack_reg[7][7]  ( .D(n623), .CLK(clk), .RST(rst), .Q(\stack[7][7] ) );
  DFF \stack_reg[0][8]  ( .D(n622), .CLK(clk), .RST(rst), .Q(o[8]) );
  DFF \stack_reg[1][8]  ( .D(n621), .CLK(clk), .RST(rst), .Q(\stack[1][8] ) );
  DFF \stack_reg[2][8]  ( .D(n620), .CLK(clk), .RST(rst), .Q(\stack[2][8] ) );
  DFF \stack_reg[3][8]  ( .D(n619), .CLK(clk), .RST(rst), .Q(\stack[3][8] ) );
  DFF \stack_reg[4][8]  ( .D(n618), .CLK(clk), .RST(rst), .Q(\stack[4][8] ) );
  DFF \stack_reg[5][8]  ( .D(n617), .CLK(clk), .RST(rst), .Q(\stack[5][8] ) );
  DFF \stack_reg[6][8]  ( .D(n616), .CLK(clk), .RST(rst), .Q(\stack[6][8] ) );
  DFF \stack_reg[7][8]  ( .D(n615), .CLK(clk), .RST(rst), .Q(\stack[7][8] ) );
  DFF \stack_reg[0][9]  ( .D(n614), .CLK(clk), .RST(rst), .Q(o[9]) );
  DFF \stack_reg[1][9]  ( .D(n613), .CLK(clk), .RST(rst), .Q(\stack[1][9] ) );
  DFF \stack_reg[2][9]  ( .D(n612), .CLK(clk), .RST(rst), .Q(\stack[2][9] ) );
  DFF \stack_reg[3][9]  ( .D(n611), .CLK(clk), .RST(rst), .Q(\stack[3][9] ) );
  DFF \stack_reg[4][9]  ( .D(n610), .CLK(clk), .RST(rst), .Q(\stack[4][9] ) );
  DFF \stack_reg[5][9]  ( .D(n609), .CLK(clk), .RST(rst), .Q(\stack[5][9] ) );
  DFF \stack_reg[6][9]  ( .D(n608), .CLK(clk), .RST(rst), .Q(\stack[6][9] ) );
  DFF \stack_reg[7][9]  ( .D(n607), .CLK(clk), .RST(rst), .Q(\stack[7][9] ) );
  DFF \stack_reg[0][10]  ( .D(n606), .CLK(clk), .RST(rst), .Q(o[10]) );
  DFF \stack_reg[1][10]  ( .D(n605), .CLK(clk), .RST(rst), .Q(\stack[1][10] )
         );
  DFF \stack_reg[2][10]  ( .D(n604), .CLK(clk), .RST(rst), .Q(\stack[2][10] )
         );
  DFF \stack_reg[3][10]  ( .D(n603), .CLK(clk), .RST(rst), .Q(\stack[3][10] )
         );
  DFF \stack_reg[4][10]  ( .D(n602), .CLK(clk), .RST(rst), .Q(\stack[4][10] )
         );
  DFF \stack_reg[5][10]  ( .D(n601), .CLK(clk), .RST(rst), .Q(\stack[5][10] )
         );
  DFF \stack_reg[6][10]  ( .D(n600), .CLK(clk), .RST(rst), .Q(\stack[6][10] )
         );
  DFF \stack_reg[7][10]  ( .D(n599), .CLK(clk), .RST(rst), .Q(\stack[7][10] )
         );
  DFF \stack_reg[0][11]  ( .D(n598), .CLK(clk), .RST(rst), .Q(o[11]) );
  DFF \stack_reg[1][11]  ( .D(n597), .CLK(clk), .RST(rst), .Q(\stack[1][11] )
         );
  DFF \stack_reg[2][11]  ( .D(n596), .CLK(clk), .RST(rst), .Q(\stack[2][11] )
         );
  DFF \stack_reg[3][11]  ( .D(n595), .CLK(clk), .RST(rst), .Q(\stack[3][11] )
         );
  DFF \stack_reg[4][11]  ( .D(n594), .CLK(clk), .RST(rst), .Q(\stack[4][11] )
         );
  DFF \stack_reg[5][11]  ( .D(n593), .CLK(clk), .RST(rst), .Q(\stack[5][11] )
         );
  DFF \stack_reg[6][11]  ( .D(n592), .CLK(clk), .RST(rst), .Q(\stack[6][11] )
         );
  DFF \stack_reg[7][11]  ( .D(n591), .CLK(clk), .RST(rst), .Q(\stack[7][11] )
         );
  DFF \stack_reg[0][12]  ( .D(n590), .CLK(clk), .RST(rst), .Q(o[12]) );
  DFF \stack_reg[1][12]  ( .D(n589), .CLK(clk), .RST(rst), .Q(\stack[1][12] )
         );
  DFF \stack_reg[2][12]  ( .D(n588), .CLK(clk), .RST(rst), .Q(\stack[2][12] )
         );
  DFF \stack_reg[3][12]  ( .D(n587), .CLK(clk), .RST(rst), .Q(\stack[3][12] )
         );
  DFF \stack_reg[4][12]  ( .D(n586), .CLK(clk), .RST(rst), .Q(\stack[4][12] )
         );
  DFF \stack_reg[5][12]  ( .D(n585), .CLK(clk), .RST(rst), .Q(\stack[5][12] )
         );
  DFF \stack_reg[6][12]  ( .D(n584), .CLK(clk), .RST(rst), .Q(\stack[6][12] )
         );
  DFF \stack_reg[7][12]  ( .D(n583), .CLK(clk), .RST(rst), .Q(\stack[7][12] )
         );
  DFF \stack_reg[0][13]  ( .D(n582), .CLK(clk), .RST(rst), .Q(o[13]) );
  DFF \stack_reg[1][13]  ( .D(n581), .CLK(clk), .RST(rst), .Q(\stack[1][13] )
         );
  DFF \stack_reg[2][13]  ( .D(n580), .CLK(clk), .RST(rst), .Q(\stack[2][13] )
         );
  DFF \stack_reg[3][13]  ( .D(n579), .CLK(clk), .RST(rst), .Q(\stack[3][13] )
         );
  DFF \stack_reg[4][13]  ( .D(n578), .CLK(clk), .RST(rst), .Q(\stack[4][13] )
         );
  DFF \stack_reg[5][13]  ( .D(n577), .CLK(clk), .RST(rst), .Q(\stack[5][13] )
         );
  DFF \stack_reg[6][13]  ( .D(n576), .CLK(clk), .RST(rst), .Q(\stack[6][13] )
         );
  DFF \stack_reg[7][13]  ( .D(n575), .CLK(clk), .RST(rst), .Q(\stack[7][13] )
         );
  DFF \stack_reg[0][14]  ( .D(n574), .CLK(clk), .RST(rst), .Q(o[14]) );
  DFF \stack_reg[1][14]  ( .D(n573), .CLK(clk), .RST(rst), .Q(\stack[1][14] )
         );
  DFF \stack_reg[2][14]  ( .D(n572), .CLK(clk), .RST(rst), .Q(\stack[2][14] )
         );
  DFF \stack_reg[3][14]  ( .D(n571), .CLK(clk), .RST(rst), .Q(\stack[3][14] )
         );
  DFF \stack_reg[4][14]  ( .D(n570), .CLK(clk), .RST(rst), .Q(\stack[4][14] )
         );
  DFF \stack_reg[5][14]  ( .D(n569), .CLK(clk), .RST(rst), .Q(\stack[5][14] )
         );
  DFF \stack_reg[6][14]  ( .D(n568), .CLK(clk), .RST(rst), .Q(\stack[6][14] )
         );
  DFF \stack_reg[7][14]  ( .D(n567), .CLK(clk), .RST(rst), .Q(\stack[7][14] )
         );
  DFF \stack_reg[0][15]  ( .D(n566), .CLK(clk), .RST(rst), .Q(o[15]) );
  DFF \stack_reg[1][15]  ( .D(n565), .CLK(clk), .RST(rst), .Q(\stack[1][15] )
         );
  DFF \stack_reg[2][15]  ( .D(n564), .CLK(clk), .RST(rst), .Q(\stack[2][15] )
         );
  DFF \stack_reg[3][15]  ( .D(n563), .CLK(clk), .RST(rst), .Q(\stack[3][15] )
         );
  DFF \stack_reg[4][15]  ( .D(n562), .CLK(clk), .RST(rst), .Q(\stack[4][15] )
         );
  DFF \stack_reg[5][15]  ( .D(n561), .CLK(clk), .RST(rst), .Q(\stack[5][15] )
         );
  DFF \stack_reg[6][15]  ( .D(n560), .CLK(clk), .RST(rst), .Q(\stack[6][15] )
         );
  DFF \stack_reg[7][15]  ( .D(n559), .CLK(clk), .RST(rst), .Q(\stack[7][15] )
         );
  DFF \stack_reg[2][0]  ( .D(n558), .CLK(clk), .RST(rst), .Q(\stack[2][0] ) );
  DFF \stack_reg[3][0]  ( .D(n557), .CLK(clk), .RST(rst), .Q(\stack[3][0] ) );
  DFF \stack_reg[4][0]  ( .D(n556), .CLK(clk), .RST(rst), .Q(\stack[4][0] ) );
  DFF \stack_reg[5][0]  ( .D(n555), .CLK(clk), .RST(rst), .Q(\stack[5][0] ) );
  DFF \stack_reg[6][0]  ( .D(n554), .CLK(clk), .RST(rst), .Q(\stack[6][0] ) );
  DFF \stack_reg[7][0]  ( .D(n553), .CLK(clk), .RST(rst), .Q(\stack[7][0] ) );
  XOR \DP_OP_25_64_3291/U80  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_0 ), .Z(
        \DP_OP_25_64_3291/n169 ) );
  XOR \DP_OP_25_64_3291/U79  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_1 ), .Z(
        \DP_OP_25_64_3291/n168 ) );
  XOR \DP_OP_25_64_3291/U78  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_2 ), .Z(
        \DP_OP_25_64_3291/n167 ) );
  XOR \DP_OP_25_64_3291/U77  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_3 ), .Z(
        \DP_OP_25_64_3291/n166 ) );
  XOR \DP_OP_25_64_3291/U76  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_4 ), .Z(
        \DP_OP_25_64_3291/n165 ) );
  XOR \DP_OP_25_64_3291/U75  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_5 ), .Z(
        \DP_OP_25_64_3291/n164 ) );
  XOR \DP_OP_25_64_3291/U74  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_6 ), .Z(
        \DP_OP_25_64_3291/n163 ) );
  XOR \DP_OP_25_64_3291/U73  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_7 ), .Z(
        \DP_OP_25_64_3291/n162 ) );
  XOR \DP_OP_25_64_3291/U72  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_8 ), .Z(
        \DP_OP_25_64_3291/n161 ) );
  XOR \DP_OP_25_64_3291/U71  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_9 ), .Z(
        \DP_OP_25_64_3291/n160 ) );
  XOR \DP_OP_25_64_3291/U70  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_10 ), .Z(
        \DP_OP_25_64_3291/n159 ) );
  XOR \DP_OP_25_64_3291/U69  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_11 ), .Z(
        \DP_OP_25_64_3291/n158 ) );
  XOR \DP_OP_25_64_3291/U68  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_12 ), .Z(
        \DP_OP_25_64_3291/n157 ) );
  XOR \DP_OP_25_64_3291/U67  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_13 ), .Z(
        \DP_OP_25_64_3291/n156 ) );
  XOR \DP_OP_25_64_3291/U66  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_14 ), .Z(
        \DP_OP_25_64_3291/n155 ) );
  XOR \DP_OP_25_64_3291/U65  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_15 ), .Z(
        \DP_OP_25_64_3291/n154 ) );
  XOR \DP_OP_25_64_3291/U62  ( .A(\U1/RSOP_16/C2/Z_0 ), .B(\C1/Z_0 ), .Z(
        \DP_OP_25_64_3291/n134 ) );
  XOR \DP_OP_25_64_3291/U61  ( .A(\DP_OP_25_64_3291/n134 ), .B(
        \DP_OP_25_64_3291/n169 ), .Z(\C3/DATA5_0 ) );
  XOR \DP_OP_25_64_3291/U60  ( .A(\DP_OP_25_64_3291/n168 ), .B(
        \U1/RSOP_16/C2/Z_1 ), .Z(\DP_OP_25_64_3291/n133 ) );
  XOR \DP_OP_25_64_3291/U59  ( .A(\DP_OP_25_64_3291/n149 ), .B(
        \DP_OP_25_64_3291/n133 ), .Z(\C3/DATA5_1 ) );
  XOR \DP_OP_25_64_3291/U58  ( .A(\DP_OP_25_64_3291/n167 ), .B(
        \U1/RSOP_16/C2/Z_2 ), .Z(\DP_OP_25_64_3291/n132 ) );
  XOR \DP_OP_25_64_3291/U57  ( .A(\DP_OP_25_64_3291/n148 ), .B(
        \DP_OP_25_64_3291/n132 ), .Z(\C3/DATA5_2 ) );
  XOR \DP_OP_25_64_3291/U56  ( .A(\DP_OP_25_64_3291/n166 ), .B(
        \U1/RSOP_16/C2/Z_3 ), .Z(\DP_OP_25_64_3291/n131 ) );
  XOR \DP_OP_25_64_3291/U55  ( .A(\DP_OP_25_64_3291/n147 ), .B(
        \DP_OP_25_64_3291/n131 ), .Z(\C3/DATA5_3 ) );
  XOR \DP_OP_25_64_3291/U54  ( .A(\DP_OP_25_64_3291/n165 ), .B(
        \U1/RSOP_16/C2/Z_4 ), .Z(\DP_OP_25_64_3291/n130 ) );
  XOR \DP_OP_25_64_3291/U53  ( .A(\DP_OP_25_64_3291/n146 ), .B(
        \DP_OP_25_64_3291/n130 ), .Z(\C3/DATA5_4 ) );
  XOR \DP_OP_25_64_3291/U52  ( .A(\DP_OP_25_64_3291/n164 ), .B(
        \U1/RSOP_16/C2/Z_5 ), .Z(\DP_OP_25_64_3291/n129 ) );
  XOR \DP_OP_25_64_3291/U51  ( .A(\DP_OP_25_64_3291/n145 ), .B(
        \DP_OP_25_64_3291/n129 ), .Z(\C3/DATA5_5 ) );
  XOR \DP_OP_25_64_3291/U50  ( .A(\DP_OP_25_64_3291/n163 ), .B(
        \U1/RSOP_16/C2/Z_6 ), .Z(\DP_OP_25_64_3291/n128 ) );
  XOR \DP_OP_25_64_3291/U49  ( .A(\DP_OP_25_64_3291/n144 ), .B(
        \DP_OP_25_64_3291/n128 ), .Z(\C3/DATA5_6 ) );
  XOR \DP_OP_25_64_3291/U48  ( .A(\DP_OP_25_64_3291/n162 ), .B(
        \U1/RSOP_16/C2/Z_7 ), .Z(\DP_OP_25_64_3291/n127 ) );
  XOR \DP_OP_25_64_3291/U47  ( .A(\DP_OP_25_64_3291/n143 ), .B(
        \DP_OP_25_64_3291/n127 ), .Z(\C3/DATA5_7 ) );
  XOR \DP_OP_25_64_3291/U46  ( .A(\DP_OP_25_64_3291/n161 ), .B(
        \U1/RSOP_16/C2/Z_8 ), .Z(\DP_OP_25_64_3291/n126 ) );
  XOR \DP_OP_25_64_3291/U45  ( .A(\DP_OP_25_64_3291/n142 ), .B(
        \DP_OP_25_64_3291/n126 ), .Z(\C3/DATA5_8 ) );
  XOR \DP_OP_25_64_3291/U44  ( .A(\DP_OP_25_64_3291/n160 ), .B(
        \U1/RSOP_16/C2/Z_9 ), .Z(\DP_OP_25_64_3291/n125 ) );
  XOR \DP_OP_25_64_3291/U43  ( .A(\DP_OP_25_64_3291/n141 ), .B(
        \DP_OP_25_64_3291/n125 ), .Z(\C3/DATA5_9 ) );
  XOR \DP_OP_25_64_3291/U42  ( .A(\DP_OP_25_64_3291/n159 ), .B(
        \U1/RSOP_16/C2/Z_10 ), .Z(\DP_OP_25_64_3291/n124 ) );
  XOR \DP_OP_25_64_3291/U41  ( .A(\DP_OP_25_64_3291/n140 ), .B(
        \DP_OP_25_64_3291/n124 ), .Z(\C3/DATA5_10 ) );
  XOR \DP_OP_25_64_3291/U40  ( .A(\DP_OP_25_64_3291/n158 ), .B(
        \U1/RSOP_16/C2/Z_11 ), .Z(\DP_OP_25_64_3291/n123 ) );
  XOR \DP_OP_25_64_3291/U30  ( .A(\DP_OP_25_64_3291/n139 ), .B(
        \DP_OP_25_64_3291/n123 ), .Z(\C3/DATA5_11 ) );
  XOR \DP_OP_25_64_3291/U20  ( .A(\DP_OP_25_64_3291/n157 ), .B(
        \U1/RSOP_16/C2/Z_12 ), .Z(\DP_OP_25_64_3291/n122 ) );
  XOR \DP_OP_25_64_3291/U10  ( .A(\DP_OP_25_64_3291/n138 ), .B(
        \DP_OP_25_64_3291/n122 ), .Z(\C3/DATA5_12 ) );
  XOR \DP_OP_25_64_3291/U9  ( .A(\DP_OP_25_64_3291/n156 ), .B(
        \U1/RSOP_16/C2/Z_13 ), .Z(\DP_OP_25_64_3291/n121 ) );
  XOR \DP_OP_25_64_3291/U8  ( .A(\DP_OP_25_64_3291/n137 ), .B(
        \DP_OP_25_64_3291/n121 ), .Z(\C3/DATA5_13 ) );
  XOR \DP_OP_25_64_3291/U7  ( .A(\DP_OP_25_64_3291/n155 ), .B(
        \U1/RSOP_16/C2/Z_14 ), .Z(\DP_OP_25_64_3291/n120 ) );
  XOR \DP_OP_25_64_3291/U6  ( .A(\DP_OP_25_64_3291/n136 ), .B(
        \DP_OP_25_64_3291/n120 ), .Z(\C3/DATA5_14 ) );
  XOR \DP_OP_25_64_3291/U5  ( .A(\DP_OP_25_64_3291/n154 ), .B(
        \U1/RSOP_16/C2/Z_15 ), .Z(\DP_OP_25_64_3291/n119 ) );
  XOR \DP_OP_25_64_3291/U4  ( .A(\DP_OP_25_64_3291/n135 ), .B(
        \DP_OP_25_64_3291/n119 ), .Z(\C3/DATA5_15 ) );
  NAND \DP_OP_25_64_3291/U114  ( .A(\DP_OP_25_64_3291/n155 ), .B(
        \U1/RSOP_16/C2/Z_14 ), .Z(\DP_OP_25_64_3291/n5 ) );
  NAND \DP_OP_25_64_3291/U214  ( .A(\DP_OP_25_64_3291/n136 ), .B(
        \DP_OP_25_64_3291/n120 ), .Z(\DP_OP_25_64_3291/n8 ) );
  NAND \DP_OP_25_64_3291/U314  ( .A(\DP_OP_25_64_3291/n5 ), .B(
        \DP_OP_25_64_3291/n8 ), .Z(\DP_OP_25_64_3291/n135 ) );
  NAND \DP_OP_25_64_3291/U113  ( .A(\DP_OP_25_64_3291/n156 ), .B(
        \U1/RSOP_16/C2/Z_13 ), .Z(\DP_OP_25_64_3291/n14 ) );
  NAND \DP_OP_25_64_3291/U213  ( .A(\DP_OP_25_64_3291/n137 ), .B(
        \DP_OP_25_64_3291/n121 ), .Z(\DP_OP_25_64_3291/n15 ) );
  NAND \DP_OP_25_64_3291/U313  ( .A(\DP_OP_25_64_3291/n14 ), .B(
        \DP_OP_25_64_3291/n15 ), .Z(\DP_OP_25_64_3291/n136 ) );
  NAND \DP_OP_25_64_3291/U112  ( .A(\DP_OP_25_64_3291/n157 ), .B(
        \U1/RSOP_16/C2/Z_12 ), .Z(\DP_OP_25_64_3291/n21 ) );
  NAND \DP_OP_25_64_3291/U212  ( .A(\DP_OP_25_64_3291/n138 ), .B(
        \DP_OP_25_64_3291/n122 ), .Z(\DP_OP_25_64_3291/n22 ) );
  NAND \DP_OP_25_64_3291/U312  ( .A(\DP_OP_25_64_3291/n21 ), .B(
        \DP_OP_25_64_3291/n22 ), .Z(\DP_OP_25_64_3291/n137 ) );
  NAND \DP_OP_25_64_3291/U111  ( .A(\DP_OP_25_64_3291/n158 ), .B(
        \U1/RSOP_16/C2/Z_11 ), .Z(\DP_OP_25_64_3291/n28 ) );
  NAND \DP_OP_25_64_3291/U211  ( .A(\DP_OP_25_64_3291/n139 ), .B(
        \DP_OP_25_64_3291/n123 ), .Z(\DP_OP_25_64_3291/n29 ) );
  NAND \DP_OP_25_64_3291/U311  ( .A(\DP_OP_25_64_3291/n28 ), .B(
        \DP_OP_25_64_3291/n29 ), .Z(\DP_OP_25_64_3291/n138 ) );
  NAND \DP_OP_25_64_3291/U110  ( .A(\DP_OP_25_64_3291/n159 ), .B(
        \U1/RSOP_16/C2/Z_10 ), .Z(\DP_OP_25_64_3291/n35 ) );
  NAND \DP_OP_25_64_3291/U210  ( .A(\DP_OP_25_64_3291/n140 ), .B(
        \DP_OP_25_64_3291/n124 ), .Z(\DP_OP_25_64_3291/n36 ) );
  NAND \DP_OP_25_64_3291/U310  ( .A(\DP_OP_25_64_3291/n35 ), .B(
        \DP_OP_25_64_3291/n36 ), .Z(\DP_OP_25_64_3291/n139 ) );
  NAND \DP_OP_25_64_3291/U19  ( .A(\DP_OP_25_64_3291/n160 ), .B(
        \U1/RSOP_16/C2/Z_9 ), .Z(\DP_OP_25_64_3291/n42 ) );
  NAND \DP_OP_25_64_3291/U29  ( .A(\DP_OP_25_64_3291/n141 ), .B(
        \DP_OP_25_64_3291/n125 ), .Z(\DP_OP_25_64_3291/n43 ) );
  NAND \DP_OP_25_64_3291/U39  ( .A(\DP_OP_25_64_3291/n42 ), .B(
        \DP_OP_25_64_3291/n43 ), .Z(\DP_OP_25_64_3291/n140 ) );
  NAND \DP_OP_25_64_3291/U18  ( .A(\DP_OP_25_64_3291/n161 ), .B(
        \U1/RSOP_16/C2/Z_8 ), .Z(\DP_OP_25_64_3291/n49 ) );
  NAND \DP_OP_25_64_3291/U28  ( .A(\DP_OP_25_64_3291/n142 ), .B(
        \DP_OP_25_64_3291/n126 ), .Z(\DP_OP_25_64_3291/n50 ) );
  NAND \DP_OP_25_64_3291/U38  ( .A(\DP_OP_25_64_3291/n49 ), .B(
        \DP_OP_25_64_3291/n50 ), .Z(\DP_OP_25_64_3291/n141 ) );
  NAND \DP_OP_25_64_3291/U17  ( .A(\DP_OP_25_64_3291/n162 ), .B(
        \U1/RSOP_16/C2/Z_7 ), .Z(\DP_OP_25_64_3291/n56 ) );
  NAND \DP_OP_25_64_3291/U27  ( .A(\DP_OP_25_64_3291/n143 ), .B(
        \DP_OP_25_64_3291/n127 ), .Z(\DP_OP_25_64_3291/n57 ) );
  NAND \DP_OP_25_64_3291/U37  ( .A(\DP_OP_25_64_3291/n56 ), .B(
        \DP_OP_25_64_3291/n57 ), .Z(\DP_OP_25_64_3291/n142 ) );
  NAND \DP_OP_25_64_3291/U16  ( .A(\DP_OP_25_64_3291/n163 ), .B(
        \U1/RSOP_16/C2/Z_6 ), .Z(\DP_OP_25_64_3291/n69 ) );
  NAND \DP_OP_25_64_3291/U26  ( .A(\DP_OP_25_64_3291/n144 ), .B(
        \DP_OP_25_64_3291/n128 ), .Z(\DP_OP_25_64_3291/n70 ) );
  NAND \DP_OP_25_64_3291/U36  ( .A(\DP_OP_25_64_3291/n69 ), .B(
        \DP_OP_25_64_3291/n70 ), .Z(\DP_OP_25_64_3291/n143 ) );
  NAND \DP_OP_25_64_3291/U15  ( .A(\DP_OP_25_64_3291/n164 ), .B(
        \U1/RSOP_16/C2/Z_5 ), .Z(\DP_OP_25_64_3291/n81 ) );
  NAND \DP_OP_25_64_3291/U25  ( .A(\DP_OP_25_64_3291/n145 ), .B(
        \DP_OP_25_64_3291/n129 ), .Z(\DP_OP_25_64_3291/n82 ) );
  NAND \DP_OP_25_64_3291/U35  ( .A(\DP_OP_25_64_3291/n81 ), .B(
        \DP_OP_25_64_3291/n82 ), .Z(\DP_OP_25_64_3291/n144 ) );
  NAND \DP_OP_25_64_3291/U14  ( .A(\DP_OP_25_64_3291/n165 ), .B(
        \U1/RSOP_16/C2/Z_4 ), .Z(\DP_OP_25_64_3291/n88 ) );
  NAND \DP_OP_25_64_3291/U24  ( .A(\DP_OP_25_64_3291/n146 ), .B(
        \DP_OP_25_64_3291/n130 ), .Z(\DP_OP_25_64_3291/n89 ) );
  NAND \DP_OP_25_64_3291/U34  ( .A(\DP_OP_25_64_3291/n88 ), .B(
        \DP_OP_25_64_3291/n89 ), .Z(\DP_OP_25_64_3291/n145 ) );
  NAND \DP_OP_25_64_3291/U13  ( .A(\DP_OP_25_64_3291/n166 ), .B(
        \U1/RSOP_16/C2/Z_3 ), .Z(\DP_OP_25_64_3291/n95 ) );
  NAND \DP_OP_25_64_3291/U23  ( .A(\DP_OP_25_64_3291/n147 ), .B(
        \DP_OP_25_64_3291/n131 ), .Z(\DP_OP_25_64_3291/n96 ) );
  NAND \DP_OP_25_64_3291/U33  ( .A(\DP_OP_25_64_3291/n95 ), .B(
        \DP_OP_25_64_3291/n96 ), .Z(\DP_OP_25_64_3291/n146 ) );
  NAND \DP_OP_25_64_3291/U12  ( .A(\DP_OP_25_64_3291/n167 ), .B(
        \U1/RSOP_16/C2/Z_2 ), .Z(\DP_OP_25_64_3291/n102 ) );
  NAND \DP_OP_25_64_3291/U22  ( .A(\DP_OP_25_64_3291/n148 ), .B(
        \DP_OP_25_64_3291/n132 ), .Z(\DP_OP_25_64_3291/n103 ) );
  NAND \DP_OP_25_64_3291/U32  ( .A(\DP_OP_25_64_3291/n102 ), .B(
        \DP_OP_25_64_3291/n103 ), .Z(\DP_OP_25_64_3291/n147 ) );
  NAND \DP_OP_25_64_3291/U11  ( .A(\DP_OP_25_64_3291/n168 ), .B(
        \U1/RSOP_16/C2/Z_1 ), .Z(\DP_OP_25_64_3291/n109 ) );
  NAND \DP_OP_25_64_3291/U21  ( .A(\DP_OP_25_64_3291/n149 ), .B(
        \DP_OP_25_64_3291/n133 ), .Z(\DP_OP_25_64_3291/n110 ) );
  NAND \DP_OP_25_64_3291/U31  ( .A(\DP_OP_25_64_3291/n109 ), .B(
        \DP_OP_25_64_3291/n110 ), .Z(\DP_OP_25_64_3291/n148 ) );
  NAND \DP_OP_25_64_3291/U1  ( .A(\U1/RSOP_16/C2/Z_0 ), .B(\C1/Z_0 ), .Z(
        \DP_OP_25_64_3291/n116 ) );
  NAND \DP_OP_25_64_3291/U2  ( .A(\DP_OP_25_64_3291/n134 ), .B(
        \DP_OP_25_64_3291/n169 ), .Z(\DP_OP_25_64_3291/n117 ) );
  NAND \DP_OP_25_64_3291/U3  ( .A(\DP_OP_25_64_3291/n116 ), .B(
        \DP_OP_25_64_3291/n117 ), .Z(\DP_OP_25_64_3291/n149 ) );
  NAND U758 ( .A(n1374), .B(n1376), .Z(n757) );
  XOR U759 ( .A(n1374), .B(n1376), .Z(n758) );
  NAND U760 ( .A(n758), .B(n1373), .Z(n759) );
  NAND U761 ( .A(n757), .B(n759), .Z(n1382) );
  NAND U762 ( .A(n1271), .B(n1272), .Z(n760) );
  XOR U763 ( .A(n1271), .B(n1272), .Z(n761) );
  NANDN U764 ( .A(n1270), .B(n761), .Z(n762) );
  NAND U765 ( .A(n760), .B(n762), .Z(n1295) );
  XNOR U766 ( .A(n1011), .B(n1012), .Z(n763) );
  XNOR U767 ( .A(n1010), .B(n763), .Z(n1035) );
  NAND U768 ( .A(n1493), .B(n1491), .Z(n764) );
  XOR U769 ( .A(n1493), .B(n1491), .Z(n765) );
  NANDN U770 ( .A(n1490), .B(n765), .Z(n766) );
  NAND U771 ( .A(n764), .B(n766), .Z(n1496) );
  NAND U772 ( .A(n1473), .B(n1475), .Z(n767) );
  XOR U773 ( .A(n1473), .B(n1475), .Z(n768) );
  NAND U774 ( .A(n768), .B(n1474), .Z(n769) );
  NAND U775 ( .A(n767), .B(n769), .Z(n1478) );
  OR U776 ( .A(n1469), .B(n1472), .Z(n1323) );
  XOR U777 ( .A(n1536), .B(n1537), .Z(n1827) );
  NAND U778 ( .A(n1119), .B(n1116), .Z(n770) );
  XOR U779 ( .A(n1119), .B(n1116), .Z(n771) );
  NANDN U780 ( .A(n1117), .B(n771), .Z(n772) );
  NAND U781 ( .A(n770), .B(n772), .Z(n1145) );
  XOR U782 ( .A(n1108), .B(n1109), .Z(n773) );
  XNOR U783 ( .A(n1107), .B(n773), .Z(n1110) );
  NAND U784 ( .A(n1031), .B(n1034), .Z(n774) );
  XOR U785 ( .A(n1031), .B(n1034), .Z(n775) );
  NAND U786 ( .A(n775), .B(n1032), .Z(n776) );
  NAND U787 ( .A(n774), .B(n776), .Z(n1036) );
  NAND U788 ( .A(n1458), .B(n1460), .Z(n777) );
  XOR U789 ( .A(n1458), .B(n1460), .Z(n778) );
  NAND U790 ( .A(n778), .B(n1457), .Z(n779) );
  NAND U791 ( .A(n777), .B(n779), .Z(n1472) );
  NAND U792 ( .A(n1343), .B(n1344), .Z(n780) );
  XOR U793 ( .A(n1343), .B(n1344), .Z(n781) );
  NANDN U794 ( .A(n1342), .B(n781), .Z(n782) );
  NAND U795 ( .A(n780), .B(n782), .Z(n1356) );
  NAND U796 ( .A(n1573), .B(n1575), .Z(n783) );
  XOR U797 ( .A(n1573), .B(n1575), .Z(n784) );
  NAND U798 ( .A(n784), .B(n1572), .Z(n785) );
  NAND U799 ( .A(n783), .B(n785), .Z(n1578) );
  XOR U800 ( .A(n1520), .B(n1521), .Z(n1904) );
  NAND U801 ( .A(n1338), .B(n1339), .Z(n786) );
  XOR U802 ( .A(n1338), .B(n1339), .Z(n787) );
  NANDN U803 ( .A(n1341), .B(n787), .Z(n788) );
  NAND U804 ( .A(n786), .B(n788), .Z(n1350) );
  NAND U805 ( .A(n1274), .B(n1273), .Z(n789) );
  XOR U806 ( .A(n1274), .B(n1273), .Z(n790) );
  NAND U807 ( .A(n790), .B(n1275), .Z(n791) );
  NAND U808 ( .A(n789), .B(n791), .Z(n1289) );
  NAND U809 ( .A(n1047), .B(n1044), .Z(n792) );
  XOR U810 ( .A(n1047), .B(n1044), .Z(n793) );
  NANDN U811 ( .A(n1045), .B(n793), .Z(n794) );
  NAND U812 ( .A(n792), .B(n794), .Z(n1070) );
  NAND U813 ( .A(n1301), .B(n1303), .Z(n795) );
  XOR U814 ( .A(n1301), .B(n1303), .Z(n796) );
  NAND U815 ( .A(n796), .B(n1302), .Z(n797) );
  NAND U816 ( .A(n795), .B(n797), .Z(n1315) );
  XNOR U817 ( .A(n1478), .B(n1477), .Z(n798) );
  XNOR U818 ( .A(n1479), .B(n798), .Z(n1476) );
  NAND U819 ( .A(n1499), .B(n1497), .Z(n799) );
  XOR U820 ( .A(n1499), .B(n1497), .Z(n800) );
  NAND U821 ( .A(n800), .B(n1496), .Z(n801) );
  NAND U822 ( .A(n799), .B(n801), .Z(n1506) );
  XOR U823 ( .A(n1504), .B(n1505), .Z(n1981) );
  NAND U824 ( .A(n1385), .B(n1383), .Z(n802) );
  XOR U825 ( .A(n1385), .B(n1383), .Z(n803) );
  NAND U826 ( .A(n803), .B(n1382), .Z(n804) );
  NAND U827 ( .A(n802), .B(n804), .Z(n1394) );
  XNOR U828 ( .A(n1171), .B(n1170), .Z(n805) );
  XNOR U829 ( .A(n1173), .B(n805), .Z(n1353) );
  NAND U830 ( .A(n1152), .B(n1150), .Z(n806) );
  XOR U831 ( .A(n1152), .B(n1150), .Z(n807) );
  NAND U832 ( .A(n807), .B(n1149), .Z(n808) );
  NAND U833 ( .A(n806), .B(n808), .Z(n1161) );
  XNOR U834 ( .A(n1036), .B(n1037), .Z(n809) );
  XNOR U835 ( .A(n1035), .B(n809), .Z(n1038) );
  NAND U836 ( .A(n1305), .B(n1307), .Z(n810) );
  XOR U837 ( .A(n1305), .B(n1307), .Z(n811) );
  NAND U838 ( .A(n811), .B(n1306), .Z(n812) );
  NAND U839 ( .A(n810), .B(n812), .Z(n1326) );
  NAND U840 ( .A(n1531), .B(n1529), .Z(n813) );
  XOR U841 ( .A(n1531), .B(n1529), .Z(n814) );
  NAND U842 ( .A(n814), .B(n1528), .Z(n815) );
  NAND U843 ( .A(n813), .B(n815), .Z(n1538) );
  XOR U844 ( .A(n1479), .B(n1477), .Z(n816) );
  NAND U845 ( .A(n816), .B(n1478), .Z(n817) );
  NAND U846 ( .A(n1479), .B(n1477), .Z(n818) );
  AND U847 ( .A(n817), .B(n818), .Z(n1480) );
  XOR U848 ( .A(n1488), .B(n1489), .Z(n2058) );
  NAND U849 ( .A(n1096), .B(n1097), .Z(n819) );
  XOR U850 ( .A(n1096), .B(n1097), .Z(n820) );
  NANDN U851 ( .A(n1098), .B(n820), .Z(n821) );
  NAND U852 ( .A(n819), .B(n821), .Z(n1106) );
  XOR U853 ( .A(n1274), .B(n1275), .Z(n822) );
  XNOR U854 ( .A(n1273), .B(n822), .Z(n1293) );
  XOR U855 ( .A(n1334), .B(n1335), .Z(n1493) );
  AND U856 ( .A(n1164), .B(n1163), .Z(n823) );
  XNOR U857 ( .A(n1115), .B(n1114), .Z(n824) );
  XNOR U858 ( .A(n823), .B(n824), .Z(n825) );
  OR U859 ( .A(n1327), .B(n1328), .Z(n826) );
  NANDN U860 ( .A(n1326), .B(n1324), .Z(n827) );
  AND U861 ( .A(n826), .B(n827), .Z(n828) );
  AND U862 ( .A(n1323), .B(n1322), .Z(n829) );
  XNOR U863 ( .A(n825), .B(n828), .Z(n830) );
  XNOR U864 ( .A(n829), .B(n830), .Z(n831) );
  NAND U865 ( .A(n1329), .B(n1331), .Z(n832) );
  XOR U866 ( .A(n1329), .B(n1331), .Z(n833) );
  NAND U867 ( .A(n1330), .B(n833), .Z(n834) );
  AND U868 ( .A(n832), .B(n834), .Z(n835) );
  XNOR U869 ( .A(n831), .B(n835), .Z(n836) );
  NANDN U870 ( .A(n1581), .B(n1579), .Z(n837) );
  OR U871 ( .A(n1579), .B(n1476), .Z(n838) );
  NAND U872 ( .A(n1578), .B(n838), .Z(n839) );
  NAND U873 ( .A(n837), .B(n839), .Z(n840) );
  XNOR U874 ( .A(n836), .B(n840), .Z(n1481) );
  XOR U875 ( .A(n1482), .B(n1483), .Z(n2096) );
  ANDN U876 ( .B(opcode[1]), .A(opcode[0]), .Z(n841) );
  NANDN U877 ( .A(opcode[2]), .B(n841), .Z(n877) );
  ANDN U878 ( .B(opcode[0]), .A(opcode[1]), .Z(n878) );
  NANDN U879 ( .A(opcode[2]), .B(n878), .Z(n842) );
  NAND U880 ( .A(n877), .B(n842), .Z(n873) );
  AND U881 ( .A(o[15]), .B(n873), .Z(\U1/RSOP_16/C2/Z_15 ) );
  AND U882 ( .A(o[14]), .B(n873), .Z(\U1/RSOP_16/C2/Z_14 ) );
  AND U883 ( .A(o[13]), .B(n873), .Z(\U1/RSOP_16/C2/Z_13 ) );
  AND U884 ( .A(o[12]), .B(n873), .Z(\U1/RSOP_16/C2/Z_12 ) );
  AND U885 ( .A(o[11]), .B(n873), .Z(\U1/RSOP_16/C2/Z_11 ) );
  AND U886 ( .A(o[10]), .B(n873), .Z(\U1/RSOP_16/C2/Z_10 ) );
  AND U887 ( .A(o[9]), .B(n873), .Z(\U1/RSOP_16/C2/Z_9 ) );
  AND U888 ( .A(o[8]), .B(n873), .Z(\U1/RSOP_16/C2/Z_8 ) );
  AND U889 ( .A(o[7]), .B(n873), .Z(\U1/RSOP_16/C2/Z_7 ) );
  AND U890 ( .A(o[6]), .B(n873), .Z(\U1/RSOP_16/C2/Z_6 ) );
  AND U891 ( .A(o[5]), .B(n873), .Z(\U1/RSOP_16/C2/Z_5 ) );
  AND U892 ( .A(o[4]), .B(n873), .Z(\U1/RSOP_16/C2/Z_4 ) );
  AND U893 ( .A(o[3]), .B(n873), .Z(\U1/RSOP_16/C2/Z_3 ) );
  AND U894 ( .A(o[2]), .B(n873), .Z(\U1/RSOP_16/C2/Z_2 ) );
  AND U895 ( .A(o[1]), .B(n873), .Z(\U1/RSOP_16/C2/Z_1 ) );
  AND U896 ( .A(o[0]), .B(n873), .Z(\U1/RSOP_16/C2/Z_0 ) );
  AND U897 ( .A(n878), .B(opcode[2]), .Z(n876) );
  NAND U898 ( .A(n876), .B(o[15]), .Z(n844) );
  NAND U899 ( .A(\stack[1][15] ), .B(n873), .Z(n843) );
  NAND U900 ( .A(n844), .B(n843), .Z(\U1/RSOP_16/C3/Z_15 ) );
  NAND U901 ( .A(n876), .B(o[14]), .Z(n846) );
  NAND U902 ( .A(\stack[1][14] ), .B(n873), .Z(n845) );
  NAND U903 ( .A(n846), .B(n845), .Z(\U1/RSOP_16/C3/Z_14 ) );
  NAND U904 ( .A(n876), .B(o[13]), .Z(n848) );
  NAND U905 ( .A(\stack[1][13] ), .B(n873), .Z(n847) );
  NAND U906 ( .A(n848), .B(n847), .Z(\U1/RSOP_16/C3/Z_13 ) );
  NAND U907 ( .A(n876), .B(o[12]), .Z(n850) );
  NAND U908 ( .A(\stack[1][12] ), .B(n873), .Z(n849) );
  NAND U909 ( .A(n850), .B(n849), .Z(\U1/RSOP_16/C3/Z_12 ) );
  NAND U910 ( .A(n876), .B(o[11]), .Z(n852) );
  NAND U911 ( .A(\stack[1][11] ), .B(n873), .Z(n851) );
  NAND U912 ( .A(n852), .B(n851), .Z(\U1/RSOP_16/C3/Z_11 ) );
  NAND U913 ( .A(n876), .B(o[10]), .Z(n854) );
  NAND U914 ( .A(\stack[1][10] ), .B(n873), .Z(n853) );
  NAND U915 ( .A(n854), .B(n853), .Z(\U1/RSOP_16/C3/Z_10 ) );
  NAND U916 ( .A(n876), .B(o[9]), .Z(n856) );
  NAND U917 ( .A(\stack[1][9] ), .B(n873), .Z(n855) );
  NAND U918 ( .A(n856), .B(n855), .Z(\U1/RSOP_16/C3/Z_9 ) );
  NAND U919 ( .A(n876), .B(o[8]), .Z(n858) );
  NAND U920 ( .A(\stack[1][8] ), .B(n873), .Z(n857) );
  NAND U921 ( .A(n858), .B(n857), .Z(\U1/RSOP_16/C3/Z_8 ) );
  NAND U922 ( .A(n876), .B(o[7]), .Z(n860) );
  NAND U923 ( .A(\stack[1][7] ), .B(n873), .Z(n859) );
  NAND U924 ( .A(n860), .B(n859), .Z(\U1/RSOP_16/C3/Z_7 ) );
  NAND U925 ( .A(n876), .B(o[6]), .Z(n862) );
  NAND U926 ( .A(\stack[1][6] ), .B(n873), .Z(n861) );
  NAND U927 ( .A(n862), .B(n861), .Z(\U1/RSOP_16/C3/Z_6 ) );
  NAND U928 ( .A(n876), .B(o[5]), .Z(n864) );
  NAND U929 ( .A(\stack[1][5] ), .B(n873), .Z(n863) );
  NAND U930 ( .A(n864), .B(n863), .Z(\U1/RSOP_16/C3/Z_5 ) );
  NAND U931 ( .A(n876), .B(o[4]), .Z(n866) );
  NAND U932 ( .A(\stack[1][4] ), .B(n873), .Z(n865) );
  NAND U933 ( .A(n866), .B(n865), .Z(\U1/RSOP_16/C3/Z_4 ) );
  NAND U934 ( .A(n876), .B(o[3]), .Z(n868) );
  NAND U935 ( .A(\stack[1][3] ), .B(n873), .Z(n867) );
  NAND U936 ( .A(n868), .B(n867), .Z(\U1/RSOP_16/C3/Z_3 ) );
  NAND U937 ( .A(n876), .B(o[2]), .Z(n870) );
  NAND U938 ( .A(\stack[1][2] ), .B(n873), .Z(n869) );
  NAND U939 ( .A(n870), .B(n869), .Z(\U1/RSOP_16/C3/Z_2 ) );
  NAND U940 ( .A(n876), .B(o[1]), .Z(n872) );
  NAND U941 ( .A(\stack[1][1] ), .B(n873), .Z(n871) );
  NAND U942 ( .A(n872), .B(n871), .Z(\U1/RSOP_16/C3/Z_1 ) );
  NAND U943 ( .A(n876), .B(o[0]), .Z(n875) );
  NAND U944 ( .A(\stack[1][0] ), .B(n873), .Z(n874) );
  NAND U945 ( .A(n875), .B(n874), .Z(\U1/RSOP_16/C3/Z_0 ) );
  NANDN U946 ( .A(n876), .B(n877), .Z(\C1/Z_0 ) );
  NANDN U947 ( .A(n878), .B(n877), .Z(n894) );
  NAND U948 ( .A(\C3/DATA5_15 ), .B(n894), .Z(n879) );
  ANDN U949 ( .B(n879), .A(n1598), .Z(n1599) );
  NAND U950 ( .A(\C3/DATA5_14 ), .B(n894), .Z(n880) );
  ANDN U951 ( .B(n880), .A(n1630), .Z(n1631) );
  NAND U952 ( .A(\C3/DATA5_13 ), .B(n894), .Z(n881) );
  AND U953 ( .A(n1672), .B(n881), .Z(n1677) );
  NAND U954 ( .A(\C3/DATA5_12 ), .B(n894), .Z(n882) );
  ANDN U955 ( .B(n882), .A(n1707), .Z(n1708) );
  NAND U956 ( .A(\C3/DATA5_11 ), .B(n894), .Z(n883) );
  NAND U957 ( .A(n1743), .B(n883), .Z(n1747) );
  NAND U958 ( .A(\C3/DATA5_10 ), .B(n894), .Z(n884) );
  ANDN U959 ( .B(n884), .A(n1784), .Z(n1785) );
  NAND U960 ( .A(\C3/DATA5_9 ), .B(n894), .Z(n885) );
  AND U961 ( .A(n1826), .B(n885), .Z(n1831) );
  NAND U962 ( .A(\C3/DATA5_8 ), .B(n894), .Z(n886) );
  ANDN U963 ( .B(n886), .A(n1861), .Z(n1862) );
  NAND U964 ( .A(\C3/DATA5_7 ), .B(n894), .Z(n887) );
  AND U965 ( .A(n1899), .B(n887), .Z(n1900) );
  NAND U966 ( .A(\C3/DATA5_6 ), .B(n894), .Z(n888) );
  ANDN U967 ( .B(n888), .A(n1938), .Z(n1939) );
  NAND U968 ( .A(\C3/DATA5_5 ), .B(n894), .Z(n889) );
  AND U969 ( .A(n1976), .B(n889), .Z(n1977) );
  NAND U970 ( .A(\C3/DATA5_4 ), .B(n894), .Z(n890) );
  ANDN U971 ( .B(n890), .A(n2015), .Z(n2016) );
  NAND U972 ( .A(\C3/DATA5_3 ), .B(n894), .Z(n891) );
  AND U973 ( .A(n2053), .B(n891), .Z(n2054) );
  NAND U974 ( .A(\C3/DATA5_2 ), .B(n894), .Z(n892) );
  AND U975 ( .A(n2091), .B(n892), .Z(n2092) );
  NAND U976 ( .A(\C3/DATA5_1 ), .B(n894), .Z(n893) );
  AND U977 ( .A(n2139), .B(n893), .Z(n2140) );
  NAND U978 ( .A(\C3/DATA5_0 ), .B(n894), .Z(n895) );
  NAND U979 ( .A(n2149), .B(n895), .Z(n2160) );
  NOR U980 ( .A(opcode[1]), .B(opcode[0]), .Z(n896) );
  AND U981 ( .A(opcode[2]), .B(n896), .Z(n2150) );
  NAND U982 ( .A(\stack[6][0] ), .B(n2150), .Z(n898) );
  NANDN U983 ( .A(n2150), .B(\stack[7][0] ), .Z(n897) );
  NAND U984 ( .A(n898), .B(n897), .Z(n553) );
  NAND U985 ( .A(\stack[5][0] ), .B(n2150), .Z(n901) );
  NANDN U986 ( .A(opcode[2]), .B(opcode[0]), .Z(n899) );
  ANDN U987 ( .B(n899), .A(opcode[1]), .Z(n2142) );
  NANDN U988 ( .A(n2142), .B(\stack[7][0] ), .Z(n900) );
  AND U989 ( .A(n901), .B(n900), .Z(n903) );
  ANDN U990 ( .B(n2142), .A(n2150), .Z(n2145) );
  NAND U991 ( .A(n2145), .B(\stack[6][0] ), .Z(n902) );
  NAND U992 ( .A(n903), .B(n902), .Z(n554) );
  NAND U993 ( .A(\stack[4][0] ), .B(n2150), .Z(n905) );
  NANDN U994 ( .A(n2142), .B(\stack[6][0] ), .Z(n904) );
  AND U995 ( .A(n905), .B(n904), .Z(n907) );
  NAND U996 ( .A(n2145), .B(\stack[5][0] ), .Z(n906) );
  NAND U997 ( .A(n907), .B(n906), .Z(n555) );
  NAND U998 ( .A(\stack[3][0] ), .B(n2150), .Z(n909) );
  NANDN U999 ( .A(n2142), .B(\stack[5][0] ), .Z(n908) );
  AND U1000 ( .A(n909), .B(n908), .Z(n911) );
  NAND U1001 ( .A(n2145), .B(\stack[4][0] ), .Z(n910) );
  NAND U1002 ( .A(n911), .B(n910), .Z(n556) );
  NAND U1003 ( .A(\stack[2][0] ), .B(n2150), .Z(n913) );
  NANDN U1004 ( .A(n2142), .B(\stack[4][0] ), .Z(n912) );
  AND U1005 ( .A(n913), .B(n912), .Z(n915) );
  NAND U1006 ( .A(n2145), .B(\stack[3][0] ), .Z(n914) );
  NAND U1007 ( .A(n915), .B(n914), .Z(n557) );
  NAND U1008 ( .A(n2150), .B(\stack[1][0] ), .Z(n917) );
  NANDN U1009 ( .A(n2142), .B(\stack[3][0] ), .Z(n916) );
  AND U1010 ( .A(n917), .B(n916), .Z(n919) );
  NAND U1011 ( .A(n2145), .B(\stack[2][0] ), .Z(n918) );
  NAND U1012 ( .A(n919), .B(n918), .Z(n558) );
  NAND U1013 ( .A(\stack[6][15] ), .B(n2150), .Z(n921) );
  NANDN U1014 ( .A(n2150), .B(\stack[7][15] ), .Z(n920) );
  NAND U1015 ( .A(n921), .B(n920), .Z(n559) );
  NAND U1016 ( .A(\stack[5][15] ), .B(n2150), .Z(n923) );
  NANDN U1017 ( .A(n2142), .B(\stack[7][15] ), .Z(n922) );
  AND U1018 ( .A(n923), .B(n922), .Z(n925) );
  NAND U1019 ( .A(n2145), .B(\stack[6][15] ), .Z(n924) );
  NAND U1020 ( .A(n925), .B(n924), .Z(n560) );
  NAND U1021 ( .A(\stack[4][15] ), .B(n2150), .Z(n927) );
  NANDN U1022 ( .A(n2142), .B(\stack[6][15] ), .Z(n926) );
  AND U1023 ( .A(n927), .B(n926), .Z(n929) );
  NAND U1024 ( .A(n2145), .B(\stack[5][15] ), .Z(n928) );
  NAND U1025 ( .A(n929), .B(n928), .Z(n561) );
  NAND U1026 ( .A(\stack[3][15] ), .B(n2150), .Z(n931) );
  NANDN U1027 ( .A(n2142), .B(\stack[5][15] ), .Z(n930) );
  AND U1028 ( .A(n931), .B(n930), .Z(n933) );
  NAND U1029 ( .A(n2145), .B(\stack[4][15] ), .Z(n932) );
  NAND U1030 ( .A(n933), .B(n932), .Z(n562) );
  NAND U1031 ( .A(\stack[2][15] ), .B(n2150), .Z(n935) );
  NANDN U1032 ( .A(n2142), .B(\stack[4][15] ), .Z(n934) );
  AND U1033 ( .A(n935), .B(n934), .Z(n937) );
  NAND U1034 ( .A(n2145), .B(\stack[3][15] ), .Z(n936) );
  NAND U1035 ( .A(n937), .B(n936), .Z(n563) );
  NAND U1036 ( .A(n2150), .B(\stack[1][15] ), .Z(n939) );
  NANDN U1037 ( .A(n2142), .B(\stack[3][15] ), .Z(n938) );
  AND U1038 ( .A(n939), .B(n938), .Z(n941) );
  NAND U1039 ( .A(n2145), .B(\stack[2][15] ), .Z(n940) );
  NAND U1040 ( .A(n941), .B(n940), .Z(n564) );
  NAND U1041 ( .A(n2150), .B(o[15]), .Z(n943) );
  NANDN U1042 ( .A(n2142), .B(\stack[2][15] ), .Z(n942) );
  AND U1043 ( .A(n943), .B(n942), .Z(n945) );
  NAND U1044 ( .A(\stack[1][15] ), .B(n2145), .Z(n944) );
  NAND U1045 ( .A(n945), .B(n944), .Z(n565) );
  AND U1046 ( .A(n2150), .B(x[15]), .Z(n1593) );
  AND U1047 ( .A(opcode[1]), .B(opcode[0]), .Z(n1589) );
  NANDN U1048 ( .A(opcode[2]), .B(n1589), .Z(n2151) );
  AND U1049 ( .A(o[14]), .B(\stack[1][1] ), .Z(n969) );
  AND U1050 ( .A(o[13]), .B(\stack[1][2] ), .Z(n951) );
  AND U1051 ( .A(o[0]), .B(\stack[1][14] ), .Z(n971) );
  AND U1052 ( .A(o[1]), .B(\stack[1][13] ), .Z(n970) );
  AND U1053 ( .A(n971), .B(n970), .Z(n949) );
  AND U1054 ( .A(\stack[1][14] ), .B(o[1]), .Z(n947) );
  NAND U1055 ( .A(\stack[1][0] ), .B(o[15]), .Z(n946) );
  XNOR U1056 ( .A(n947), .B(n946), .Z(n948) );
  XNOR U1057 ( .A(n949), .B(n948), .Z(n950) );
  XNOR U1058 ( .A(n951), .B(n950), .Z(n967) );
  AND U1059 ( .A(\stack[1][12] ), .B(o[3]), .Z(n953) );
  NAND U1060 ( .A(o[0]), .B(\stack[1][15] ), .Z(n952) );
  XNOR U1061 ( .A(n953), .B(n952), .Z(n957) );
  AND U1062 ( .A(o[11]), .B(\stack[1][4] ), .Z(n955) );
  NAND U1063 ( .A(o[12]), .B(\stack[1][3] ), .Z(n954) );
  XNOR U1064 ( .A(n955), .B(n954), .Z(n956) );
  XOR U1065 ( .A(n957), .B(n956), .Z(n965) );
  AND U1066 ( .A(o[8]), .B(\stack[1][7] ), .Z(n959) );
  NAND U1067 ( .A(\stack[1][11] ), .B(o[4]), .Z(n958) );
  XNOR U1068 ( .A(n959), .B(n958), .Z(n963) );
  AND U1069 ( .A(\stack[1][10] ), .B(o[5]), .Z(n961) );
  NAND U1070 ( .A(\stack[1][13] ), .B(o[2]), .Z(n960) );
  XNOR U1071 ( .A(n961), .B(n960), .Z(n962) );
  XNOR U1072 ( .A(n963), .B(n962), .Z(n964) );
  XNOR U1073 ( .A(n965), .B(n964), .Z(n966) );
  XNOR U1074 ( .A(n967), .B(n966), .Z(n968) );
  XNOR U1075 ( .A(n969), .B(n968), .Z(n976) );
  AND U1076 ( .A(o[2]), .B(\stack[1][12] ), .Z(n994) );
  AND U1077 ( .A(o[1]), .B(\stack[1][12] ), .Z(n986) );
  AND U1078 ( .A(o[0]), .B(\stack[1][13] ), .Z(n985) );
  NAND U1079 ( .A(n986), .B(n985), .Z(n992) );
  NANDN U1080 ( .A(n994), .B(n992), .Z(n974) );
  XOR U1081 ( .A(n971), .B(n970), .Z(n991) );
  ANDN U1082 ( .B(n994), .A(n992), .Z(n972) );
  OR U1083 ( .A(n991), .B(n972), .Z(n973) );
  NAND U1084 ( .A(n974), .B(n973), .Z(n975) );
  XNOR U1085 ( .A(n976), .B(n975), .Z(n984) );
  AND U1086 ( .A(\stack[1][8] ), .B(o[7]), .Z(n978) );
  NAND U1087 ( .A(\stack[1][9] ), .B(o[6]), .Z(n977) );
  XNOR U1088 ( .A(n978), .B(n977), .Z(n982) );
  AND U1089 ( .A(o[9]), .B(\stack[1][6] ), .Z(n980) );
  NAND U1090 ( .A(o[10]), .B(\stack[1][5] ), .Z(n979) );
  XNOR U1091 ( .A(n980), .B(n979), .Z(n981) );
  XNOR U1092 ( .A(n982), .B(n981), .Z(n983) );
  XNOR U1093 ( .A(n984), .B(n983), .Z(n999) );
  AND U1094 ( .A(o[0]), .B(\stack[1][12] ), .Z(n1001) );
  AND U1095 ( .A(o[1]), .B(\stack[1][11] ), .Z(n1000) );
  AND U1096 ( .A(n1001), .B(n1000), .Z(n1006) );
  NAND U1097 ( .A(o[2]), .B(\stack[1][11] ), .Z(n1008) );
  NANDN U1098 ( .A(n1006), .B(n1008), .Z(n989) );
  XOR U1099 ( .A(n986), .B(n985), .Z(n1005) );
  ANDN U1100 ( .B(n1006), .A(n1008), .Z(n987) );
  OR U1101 ( .A(n1005), .B(n987), .Z(n988) );
  AND U1102 ( .A(n989), .B(n988), .Z(n1012) );
  AND U1103 ( .A(o[3]), .B(\stack[1][11] ), .Z(n1011) );
  IV U1104 ( .A(n1011), .Z(n990) );
  NANDN U1105 ( .A(n1012), .B(n990), .Z(n997) );
  AND U1106 ( .A(n1012), .B(n1011), .Z(n995) );
  XOR U1107 ( .A(n992), .B(n991), .Z(n993) );
  XNOR U1108 ( .A(n994), .B(n993), .Z(n1010) );
  OR U1109 ( .A(n995), .B(n1010), .Z(n996) );
  NAND U1110 ( .A(n997), .B(n996), .Z(n998) );
  XNOR U1111 ( .A(n999), .B(n998), .Z(n1017) );
  XOR U1112 ( .A(n1001), .B(n1000), .Z(n1026) );
  NAND U1113 ( .A(o[2]), .B(\stack[1][10] ), .Z(n1023) );
  NANDN U1114 ( .A(n1026), .B(n1023), .Z(n1004) );
  AND U1115 ( .A(o[1]), .B(\stack[1][10] ), .Z(n1019) );
  AND U1116 ( .A(o[0]), .B(\stack[1][11] ), .Z(n1018) );
  AND U1117 ( .A(n1019), .B(n1018), .Z(n1024) );
  ANDN U1118 ( .B(n1026), .A(n1023), .Z(n1002) );
  OR U1119 ( .A(n1024), .B(n1002), .Z(n1003) );
  AND U1120 ( .A(n1004), .B(n1003), .Z(n1032) );
  AND U1121 ( .A(o[3]), .B(\stack[1][10] ), .Z(n1031) );
  XNOR U1122 ( .A(n1006), .B(n1005), .Z(n1007) );
  XOR U1123 ( .A(n1008), .B(n1007), .Z(n1034) );
  AND U1124 ( .A(o[4]), .B(\stack[1][10] ), .Z(n1037) );
  IV U1125 ( .A(n1037), .Z(n1009) );
  NANDN U1126 ( .A(n1036), .B(n1009), .Z(n1015) );
  AND U1127 ( .A(n1036), .B(n1037), .Z(n1013) );
  OR U1128 ( .A(n1013), .B(n1035), .Z(n1014) );
  NAND U1129 ( .A(n1015), .B(n1014), .Z(n1016) );
  XNOR U1130 ( .A(n1017), .B(n1016), .Z(n1043) );
  XNOR U1131 ( .A(n1019), .B(n1018), .Z(n1055) );
  NAND U1132 ( .A(o[2]), .B(\stack[1][9] ), .Z(n1059) );
  NAND U1133 ( .A(n1055), .B(n1059), .Z(n1022) );
  AND U1134 ( .A(o[0]), .B(\stack[1][10] ), .Z(n1051) );
  AND U1135 ( .A(o[1]), .B(\stack[1][9] ), .Z(n1050) );
  AND U1136 ( .A(n1051), .B(n1050), .Z(n1057) );
  NOR U1137 ( .A(n1055), .B(n1059), .Z(n1020) );
  OR U1138 ( .A(n1057), .B(n1020), .Z(n1021) );
  AND U1139 ( .A(n1022), .B(n1021), .Z(n1064) );
  XOR U1140 ( .A(n1024), .B(n1023), .Z(n1025) );
  XNOR U1141 ( .A(n1026), .B(n1025), .Z(n1027) );
  IV U1142 ( .A(n1027), .Z(n1067) );
  NANDN U1143 ( .A(n1064), .B(n1067), .Z(n1030) );
  AND U1144 ( .A(o[3]), .B(\stack[1][9] ), .Z(n1065) );
  AND U1145 ( .A(n1064), .B(n1027), .Z(n1028) );
  OR U1146 ( .A(n1065), .B(n1028), .Z(n1029) );
  AND U1147 ( .A(n1030), .B(n1029), .Z(n1044) );
  NAND U1148 ( .A(o[4]), .B(\stack[1][9] ), .Z(n1045) );
  XNOR U1149 ( .A(n1032), .B(n1031), .Z(n1033) );
  XNOR U1150 ( .A(n1034), .B(n1033), .Z(n1047) );
  IV U1151 ( .A(n1038), .Z(n1073) );
  NANDN U1152 ( .A(n1070), .B(n1073), .Z(n1041) );
  AND U1153 ( .A(o[5]), .B(\stack[1][9] ), .Z(n1071) );
  AND U1154 ( .A(n1070), .B(n1038), .Z(n1039) );
  OR U1155 ( .A(n1071), .B(n1039), .Z(n1040) );
  NAND U1156 ( .A(n1041), .B(n1040), .Z(n1042) );
  XNOR U1157 ( .A(n1043), .B(n1042), .Z(n1078) );
  AND U1158 ( .A(o[5]), .B(\stack[1][8] ), .Z(n1049) );
  XOR U1159 ( .A(n1045), .B(n1044), .Z(n1046) );
  XNOR U1160 ( .A(n1047), .B(n1046), .Z(n1048) );
  NAND U1161 ( .A(n1049), .B(n1048), .Z(n1069) );
  XOR U1162 ( .A(n1049), .B(n1048), .Z(n1105) );
  XOR U1163 ( .A(n1051), .B(n1050), .Z(n1087) );
  NAND U1164 ( .A(o[2]), .B(\stack[1][8] ), .Z(n1084) );
  NANDN U1165 ( .A(n1087), .B(n1084), .Z(n1054) );
  AND U1166 ( .A(o[1]), .B(\stack[1][8] ), .Z(n1080) );
  AND U1167 ( .A(o[0]), .B(\stack[1][9] ), .Z(n1079) );
  AND U1168 ( .A(n1080), .B(n1079), .Z(n1085) );
  ANDN U1169 ( .B(n1087), .A(n1084), .Z(n1052) );
  OR U1170 ( .A(n1085), .B(n1052), .Z(n1053) );
  AND U1171 ( .A(n1054), .B(n1053), .Z(n1095) );
  IV U1172 ( .A(n1055), .Z(n1056) );
  XNOR U1173 ( .A(n1057), .B(n1056), .Z(n1058) );
  XNOR U1174 ( .A(n1059), .B(n1058), .Z(n1060) );
  NANDN U1175 ( .A(n1095), .B(n1060), .Z(n1063) );
  AND U1176 ( .A(o[3]), .B(\stack[1][8] ), .Z(n1093) );
  IV U1177 ( .A(n1060), .Z(n1092) );
  AND U1178 ( .A(n1095), .B(n1092), .Z(n1061) );
  OR U1179 ( .A(n1093), .B(n1061), .Z(n1062) );
  AND U1180 ( .A(n1063), .B(n1062), .Z(n1097) );
  NAND U1181 ( .A(o[4]), .B(\stack[1][8] ), .Z(n1098) );
  XNOR U1182 ( .A(n1065), .B(n1064), .Z(n1066) );
  XOR U1183 ( .A(n1067), .B(n1066), .Z(n1096) );
  NAND U1184 ( .A(n1105), .B(n1106), .Z(n1068) );
  NAND U1185 ( .A(n1069), .B(n1068), .Z(n1109) );
  AND U1186 ( .A(o[6]), .B(\stack[1][8] ), .Z(n1108) );
  OR U1187 ( .A(n1109), .B(n1108), .Z(n1076) );
  AND U1188 ( .A(n1109), .B(n1108), .Z(n1074) );
  XNOR U1189 ( .A(n1071), .B(n1070), .Z(n1072) );
  XOR U1190 ( .A(n1073), .B(n1072), .Z(n1107) );
  OR U1191 ( .A(n1074), .B(n1107), .Z(n1075) );
  NAND U1192 ( .A(n1076), .B(n1075), .Z(n1077) );
  XNOR U1193 ( .A(n1078), .B(n1077), .Z(n1115) );
  XNOR U1194 ( .A(n1080), .B(n1079), .Z(n1127) );
  NAND U1195 ( .A(o[2]), .B(\stack[1][7] ), .Z(n1131) );
  NAND U1196 ( .A(n1127), .B(n1131), .Z(n1083) );
  AND U1197 ( .A(o[0]), .B(\stack[1][8] ), .Z(n1123) );
  AND U1198 ( .A(o[1]), .B(\stack[1][7] ), .Z(n1122) );
  AND U1199 ( .A(n1123), .B(n1122), .Z(n1129) );
  NOR U1200 ( .A(n1127), .B(n1131), .Z(n1081) );
  OR U1201 ( .A(n1129), .B(n1081), .Z(n1082) );
  AND U1202 ( .A(n1083), .B(n1082), .Z(n1136) );
  XOR U1203 ( .A(n1085), .B(n1084), .Z(n1086) );
  XNOR U1204 ( .A(n1087), .B(n1086), .Z(n1088) );
  IV U1205 ( .A(n1088), .Z(n1139) );
  NANDN U1206 ( .A(n1136), .B(n1139), .Z(n1091) );
  AND U1207 ( .A(o[3]), .B(\stack[1][7] ), .Z(n1137) );
  AND U1208 ( .A(n1136), .B(n1088), .Z(n1089) );
  OR U1209 ( .A(n1137), .B(n1089), .Z(n1090) );
  AND U1210 ( .A(n1091), .B(n1090), .Z(n1116) );
  NAND U1211 ( .A(o[4]), .B(\stack[1][7] ), .Z(n1117) );
  XNOR U1212 ( .A(n1093), .B(n1092), .Z(n1094) );
  XNOR U1213 ( .A(n1095), .B(n1094), .Z(n1119) );
  IV U1214 ( .A(n1096), .Z(n1100) );
  XOR U1215 ( .A(n1098), .B(n1097), .Z(n1099) );
  XOR U1216 ( .A(n1100), .B(n1099), .Z(n1101) );
  IV U1217 ( .A(n1101), .Z(n1148) );
  NANDN U1218 ( .A(n1145), .B(n1148), .Z(n1104) );
  AND U1219 ( .A(o[5]), .B(\stack[1][7] ), .Z(n1146) );
  AND U1220 ( .A(n1145), .B(n1101), .Z(n1102) );
  OR U1221 ( .A(n1146), .B(n1102), .Z(n1103) );
  AND U1222 ( .A(n1104), .B(n1103), .Z(n1149) );
  AND U1223 ( .A(o[6]), .B(\stack[1][7] ), .Z(n1152) );
  XOR U1224 ( .A(n1106), .B(n1105), .Z(n1150) );
  NANDN U1225 ( .A(n1161), .B(n1110), .Z(n1113) );
  AND U1226 ( .A(o[7]), .B(\stack[1][7] ), .Z(n1159) );
  IV U1227 ( .A(n1110), .Z(n1158) );
  AND U1228 ( .A(n1161), .B(n1158), .Z(n1111) );
  OR U1229 ( .A(n1159), .B(n1111), .Z(n1112) );
  NAND U1230 ( .A(n1113), .B(n1112), .Z(n1114) );
  AND U1231 ( .A(o[5]), .B(\stack[1][6] ), .Z(n1121) );
  XOR U1232 ( .A(n1117), .B(n1116), .Z(n1118) );
  XNOR U1233 ( .A(n1119), .B(n1118), .Z(n1120) );
  NAND U1234 ( .A(n1121), .B(n1120), .Z(n1144) );
  XOR U1235 ( .A(n1121), .B(n1120), .Z(n1250) );
  AND U1236 ( .A(o[2]), .B(\stack[1][6] ), .Z(n1183) );
  XNOR U1237 ( .A(n1123), .B(n1122), .Z(n1186) );
  NANDN U1238 ( .A(n1183), .B(n1186), .Z(n1126) );
  AND U1239 ( .A(o[1]), .B(\stack[1][6] ), .Z(n1179) );
  AND U1240 ( .A(o[0]), .B(\stack[1][7] ), .Z(n1178) );
  AND U1241 ( .A(n1179), .B(n1178), .Z(n1184) );
  ANDN U1242 ( .B(n1183), .A(n1186), .Z(n1124) );
  OR U1243 ( .A(n1184), .B(n1124), .Z(n1125) );
  AND U1244 ( .A(n1126), .B(n1125), .Z(n1212) );
  IV U1245 ( .A(n1127), .Z(n1128) );
  XNOR U1246 ( .A(n1129), .B(n1128), .Z(n1130) );
  XNOR U1247 ( .A(n1131), .B(n1130), .Z(n1132) );
  NANDN U1248 ( .A(n1212), .B(n1132), .Z(n1135) );
  AND U1249 ( .A(o[3]), .B(\stack[1][6] ), .Z(n1210) );
  IV U1250 ( .A(n1132), .Z(n1209) );
  AND U1251 ( .A(n1212), .B(n1209), .Z(n1133) );
  OR U1252 ( .A(n1210), .B(n1133), .Z(n1134) );
  AND U1253 ( .A(n1135), .B(n1134), .Z(n1225) );
  NAND U1254 ( .A(o[4]), .B(\stack[1][6] ), .Z(n1226) );
  ANDN U1255 ( .B(n1225), .A(n1226), .Z(n1140) );
  XNOR U1256 ( .A(n1137), .B(n1136), .Z(n1138) );
  XOR U1257 ( .A(n1139), .B(n1138), .Z(n1224) );
  OR U1258 ( .A(n1140), .B(n1224), .Z(n1142) );
  ANDN U1259 ( .B(n1226), .A(n1225), .Z(n1141) );
  ANDN U1260 ( .B(n1142), .A(n1141), .Z(n1251) );
  NAND U1261 ( .A(n1250), .B(n1251), .Z(n1143) );
  NAND U1262 ( .A(n1144), .B(n1143), .Z(n1275) );
  AND U1263 ( .A(\stack[1][6] ), .B(o[6]), .Z(n1274) );
  XNOR U1264 ( .A(n1146), .B(n1145), .Z(n1147) );
  XOR U1265 ( .A(n1148), .B(n1147), .Z(n1273) );
  XNOR U1266 ( .A(n1150), .B(n1149), .Z(n1151) );
  XOR U1267 ( .A(n1152), .B(n1151), .Z(n1153) );
  NANDN U1268 ( .A(n1289), .B(n1153), .Z(n1156) );
  AND U1269 ( .A(\stack[1][6] ), .B(o[7]), .Z(n1290) );
  IV U1270 ( .A(n1153), .Z(n1292) );
  AND U1271 ( .A(n1289), .B(n1292), .Z(n1154) );
  OR U1272 ( .A(n1290), .B(n1154), .Z(n1155) );
  AND U1273 ( .A(n1156), .B(n1155), .Z(n1308) );
  AND U1274 ( .A(\stack[1][6] ), .B(o[8]), .Z(n1309) );
  IV U1275 ( .A(n1309), .Z(n1157) );
  NANDN U1276 ( .A(n1308), .B(n1157), .Z(n1164) );
  AND U1277 ( .A(n1308), .B(n1309), .Z(n1162) );
  XNOR U1278 ( .A(n1159), .B(n1158), .Z(n1160) );
  XNOR U1279 ( .A(n1161), .B(n1160), .Z(n1311) );
  OR U1280 ( .A(n1162), .B(n1311), .Z(n1163) );
  AND U1281 ( .A(o[2]), .B(\stack[1][3] ), .Z(n1338) );
  AND U1282 ( .A(o[0]), .B(\stack[1][5] ), .Z(n1166) );
  AND U1283 ( .A(o[1]), .B(\stack[1][4] ), .Z(n1165) );
  XNOR U1284 ( .A(n1166), .B(n1165), .Z(n1341) );
  AND U1285 ( .A(o[1]), .B(\stack[1][3] ), .Z(n1333) );
  AND U1286 ( .A(o[0]), .B(\stack[1][4] ), .Z(n1332) );
  AND U1287 ( .A(n1333), .B(n1332), .Z(n1339) );
  NAND U1288 ( .A(o[2]), .B(\stack[1][4] ), .Z(n1170) );
  AND U1289 ( .A(n1166), .B(n1165), .Z(n1173) );
  AND U1290 ( .A(o[1]), .B(\stack[1][5] ), .Z(n1177) );
  AND U1291 ( .A(o[0]), .B(\stack[1][6] ), .Z(n1176) );
  XNOR U1292 ( .A(n1177), .B(n1176), .Z(n1171) );
  OR U1293 ( .A(n1350), .B(n1353), .Z(n1169) );
  AND U1294 ( .A(n1353), .B(n1350), .Z(n1167) );
  AND U1295 ( .A(o[3]), .B(\stack[1][3] ), .Z(n1349) );
  OR U1296 ( .A(n1167), .B(n1349), .Z(n1168) );
  AND U1297 ( .A(n1169), .B(n1168), .Z(n1373) );
  AND U1298 ( .A(\stack[1][3] ), .B(o[4]), .Z(n1374) );
  NAND U1299 ( .A(n1171), .B(n1170), .Z(n1175) );
  NOR U1300 ( .A(n1171), .B(n1170), .Z(n1172) );
  OR U1301 ( .A(n1173), .B(n1172), .Z(n1174) );
  AND U1302 ( .A(n1175), .B(n1174), .Z(n1196) );
  AND U1303 ( .A(o[3]), .B(\stack[1][4] ), .Z(n1198) );
  NAND U1304 ( .A(o[2]), .B(\stack[1][5] ), .Z(n1187) );
  AND U1305 ( .A(n1177), .B(n1176), .Z(n1190) );
  XNOR U1306 ( .A(n1179), .B(n1178), .Z(n1188) );
  IV U1307 ( .A(n1188), .Z(n1180) );
  XNOR U1308 ( .A(n1190), .B(n1180), .Z(n1181) );
  XNOR U1309 ( .A(n1187), .B(n1181), .Z(n1194) );
  IV U1310 ( .A(n1194), .Z(n1195) );
  XNOR U1311 ( .A(n1198), .B(n1195), .Z(n1182) );
  XNOR U1312 ( .A(n1196), .B(n1182), .Z(n1376) );
  XNOR U1313 ( .A(n1184), .B(n1183), .Z(n1185) );
  XNOR U1314 ( .A(n1186), .B(n1185), .Z(n1213) );
  IV U1315 ( .A(n1213), .Z(n1214) );
  AND U1316 ( .A(o[3]), .B(\stack[1][5] ), .Z(n1217) );
  NAND U1317 ( .A(n1188), .B(n1187), .Z(n1192) );
  NOR U1318 ( .A(n1188), .B(n1187), .Z(n1189) );
  OR U1319 ( .A(n1190), .B(n1189), .Z(n1191) );
  AND U1320 ( .A(n1192), .B(n1191), .Z(n1215) );
  XNOR U1321 ( .A(n1217), .B(n1215), .Z(n1193) );
  XNOR U1322 ( .A(n1214), .B(n1193), .Z(n1203) );
  NAND U1323 ( .A(\stack[1][4] ), .B(o[4]), .Z(n1206) );
  NANDN U1324 ( .A(n1196), .B(n1194), .Z(n1200) );
  AND U1325 ( .A(n1196), .B(n1195), .Z(n1197) );
  OR U1326 ( .A(n1198), .B(n1197), .Z(n1199) );
  AND U1327 ( .A(n1200), .B(n1199), .Z(n1205) );
  XOR U1328 ( .A(n1206), .B(n1205), .Z(n1201) );
  XNOR U1329 ( .A(n1203), .B(n1201), .Z(n1385) );
  AND U1330 ( .A(\stack[1][3] ), .B(o[5]), .Z(n1383) );
  AND U1331 ( .A(\stack[1][3] ), .B(o[6]), .Z(n1397) );
  IV U1332 ( .A(n1397), .Z(n1202) );
  NANDN U1333 ( .A(n1394), .B(n1202), .Z(n1223) );
  ANDN U1334 ( .B(n1205), .A(n1206), .Z(n1204) );
  OR U1335 ( .A(n1204), .B(n1203), .Z(n1208) );
  ANDN U1336 ( .B(n1206), .A(n1205), .Z(n1207) );
  ANDN U1337 ( .B(n1208), .A(n1207), .Z(n1238) );
  AND U1338 ( .A(\stack[1][4] ), .B(o[5]), .Z(n1237) );
  XNOR U1339 ( .A(n1210), .B(n1209), .Z(n1211) );
  XNOR U1340 ( .A(n1212), .B(n1211), .Z(n1229) );
  NAND U1341 ( .A(o[4]), .B(\stack[1][5] ), .Z(n1232) );
  NANDN U1342 ( .A(n1215), .B(n1213), .Z(n1219) );
  AND U1343 ( .A(n1215), .B(n1214), .Z(n1216) );
  OR U1344 ( .A(n1217), .B(n1216), .Z(n1218) );
  AND U1345 ( .A(n1219), .B(n1218), .Z(n1231) );
  XOR U1346 ( .A(n1232), .B(n1231), .Z(n1220) );
  XNOR U1347 ( .A(n1229), .B(n1220), .Z(n1236) );
  XOR U1348 ( .A(n1237), .B(n1236), .Z(n1239) );
  XOR U1349 ( .A(n1238), .B(n1239), .Z(n1395) );
  AND U1350 ( .A(n1394), .B(n1397), .Z(n1221) );
  OR U1351 ( .A(n1395), .B(n1221), .Z(n1222) );
  AND U1352 ( .A(n1223), .B(n1222), .Z(n1412) );
  IV U1353 ( .A(n1224), .Z(n1228) );
  XOR U1354 ( .A(n1226), .B(n1225), .Z(n1227) );
  XOR U1355 ( .A(n1228), .B(n1227), .Z(n1254) );
  IV U1356 ( .A(n1254), .Z(n1252) );
  NAND U1357 ( .A(o[5]), .B(\stack[1][5] ), .Z(n1256) );
  ANDN U1358 ( .B(n1231), .A(n1232), .Z(n1230) );
  OR U1359 ( .A(n1230), .B(n1229), .Z(n1234) );
  ANDN U1360 ( .B(n1232), .A(n1231), .Z(n1233) );
  ANDN U1361 ( .B(n1234), .A(n1233), .Z(n1253) );
  XOR U1362 ( .A(n1256), .B(n1253), .Z(n1235) );
  XOR U1363 ( .A(n1252), .B(n1235), .Z(n1262) );
  IV U1364 ( .A(n1262), .Z(n1244) );
  NAND U1365 ( .A(n1237), .B(n1236), .Z(n1241) );
  NAND U1366 ( .A(n1239), .B(n1238), .Z(n1240) );
  NAND U1367 ( .A(n1241), .B(n1240), .Z(n1261) );
  AND U1368 ( .A(\stack[1][4] ), .B(o[6]), .Z(n1260) );
  IV U1369 ( .A(n1260), .Z(n1242) );
  XNOR U1370 ( .A(n1261), .B(n1242), .Z(n1243) );
  XOR U1371 ( .A(n1244), .B(n1243), .Z(n1245) );
  NANDN U1372 ( .A(n1412), .B(n1245), .Z(n1248) );
  AND U1373 ( .A(\stack[1][3] ), .B(o[7]), .Z(n1410) );
  IV U1374 ( .A(n1245), .Z(n1409) );
  AND U1375 ( .A(n1412), .B(n1409), .Z(n1246) );
  OR U1376 ( .A(n1410), .B(n1246), .Z(n1247) );
  AND U1377 ( .A(n1248), .B(n1247), .Z(n1426) );
  AND U1378 ( .A(\stack[1][3] ), .B(o[8]), .Z(n1427) );
  IV U1379 ( .A(n1427), .Z(n1249) );
  NANDN U1380 ( .A(n1426), .B(n1249), .Z(n1269) );
  AND U1381 ( .A(n1426), .B(n1427), .Z(n1267) );
  NAND U1382 ( .A(\stack[1][5] ), .B(o[6]), .Z(n1270) );
  XOR U1383 ( .A(n1251), .B(n1250), .Z(n1272) );
  NANDN U1384 ( .A(n1253), .B(n1252), .Z(n1258) );
  NAND U1385 ( .A(n1254), .B(n1253), .Z(n1255) );
  NAND U1386 ( .A(n1256), .B(n1255), .Z(n1257) );
  AND U1387 ( .A(n1258), .B(n1257), .Z(n1271) );
  XNOR U1388 ( .A(n1272), .B(n1271), .Z(n1259) );
  XNOR U1389 ( .A(n1270), .B(n1259), .Z(n1277) );
  IV U1390 ( .A(n1277), .Z(n1278) );
  AND U1391 ( .A(\stack[1][4] ), .B(o[7]), .Z(n1281) );
  OR U1392 ( .A(n1261), .B(n1260), .Z(n1265) );
  AND U1393 ( .A(n1261), .B(n1260), .Z(n1263) );
  OR U1394 ( .A(n1263), .B(n1262), .Z(n1264) );
  AND U1395 ( .A(n1265), .B(n1264), .Z(n1279) );
  XNOR U1396 ( .A(n1281), .B(n1279), .Z(n1266) );
  XNOR U1397 ( .A(n1278), .B(n1266), .Z(n1429) );
  OR U1398 ( .A(n1267), .B(n1429), .Z(n1268) );
  AND U1399 ( .A(n1269), .B(n1268), .Z(n1444) );
  AND U1400 ( .A(\stack[1][5] ), .B(o[7]), .Z(n1297) );
  IV U1401 ( .A(n1293), .Z(n1294) );
  XNOR U1402 ( .A(n1297), .B(n1294), .Z(n1276) );
  XNOR U1403 ( .A(n1295), .B(n1276), .Z(n1303) );
  AND U1404 ( .A(\stack[1][4] ), .B(o[8]), .Z(n1301) );
  NANDN U1405 ( .A(n1279), .B(n1277), .Z(n1283) );
  AND U1406 ( .A(n1279), .B(n1278), .Z(n1280) );
  OR U1407 ( .A(n1281), .B(n1280), .Z(n1282) );
  AND U1408 ( .A(n1283), .B(n1282), .Z(n1302) );
  XNOR U1409 ( .A(n1301), .B(n1302), .Z(n1284) );
  XNOR U1410 ( .A(n1303), .B(n1284), .Z(n1441) );
  IV U1411 ( .A(n1441), .Z(n1285) );
  NANDN U1412 ( .A(n1444), .B(n1285), .Z(n1288) );
  AND U1413 ( .A(\stack[1][3] ), .B(o[9]), .Z(n1442) );
  AND U1414 ( .A(n1444), .B(n1441), .Z(n1286) );
  OR U1415 ( .A(n1442), .B(n1286), .Z(n1287) );
  AND U1416 ( .A(n1288), .B(n1287), .Z(n1457) );
  AND U1417 ( .A(\stack[1][3] ), .B(o[10]), .Z(n1458) );
  XNOR U1418 ( .A(n1290), .B(n1289), .Z(n1291) );
  XNOR U1419 ( .A(n1292), .B(n1291), .Z(n1307) );
  AND U1420 ( .A(\stack[1][5] ), .B(o[8]), .Z(n1305) );
  NANDN U1421 ( .A(n1295), .B(n1293), .Z(n1299) );
  AND U1422 ( .A(n1295), .B(n1294), .Z(n1296) );
  OR U1423 ( .A(n1297), .B(n1296), .Z(n1298) );
  AND U1424 ( .A(n1299), .B(n1298), .Z(n1306) );
  XNOR U1425 ( .A(n1305), .B(n1306), .Z(n1300) );
  XNOR U1426 ( .A(n1307), .B(n1300), .Z(n1314) );
  AND U1427 ( .A(\stack[1][4] ), .B(o[9]), .Z(n1317) );
  XNOR U1428 ( .A(n1317), .B(n1315), .Z(n1304) );
  XNOR U1429 ( .A(n1314), .B(n1304), .Z(n1460) );
  AND U1430 ( .A(\stack[1][5] ), .B(o[9]), .Z(n1328) );
  XNOR U1431 ( .A(n1309), .B(n1308), .Z(n1310) );
  XNOR U1432 ( .A(n1311), .B(n1310), .Z(n1325) );
  XNOR U1433 ( .A(n1328), .B(n1325), .Z(n1312) );
  XNOR U1434 ( .A(n1326), .B(n1312), .Z(n1331) );
  AND U1435 ( .A(\stack[1][4] ), .B(o[10]), .Z(n1329) );
  IV U1436 ( .A(n1314), .Z(n1313) );
  NANDN U1437 ( .A(n1315), .B(n1313), .Z(n1319) );
  AND U1438 ( .A(n1315), .B(n1314), .Z(n1316) );
  OR U1439 ( .A(n1317), .B(n1316), .Z(n1318) );
  AND U1440 ( .A(n1319), .B(n1318), .Z(n1330) );
  XNOR U1441 ( .A(n1329), .B(n1330), .Z(n1320) );
  XNOR U1442 ( .A(n1331), .B(n1320), .Z(n1469) );
  AND U1443 ( .A(\stack[1][3] ), .B(o[11]), .Z(n1470) );
  AND U1444 ( .A(n1472), .B(n1469), .Z(n1321) );
  OR U1445 ( .A(n1470), .B(n1321), .Z(n1322) );
  IV U1446 ( .A(n1325), .Z(n1324) );
  AND U1447 ( .A(n1326), .B(n1325), .Z(n1327) );
  AND U1448 ( .A(o[0]), .B(\stack[1][3] ), .Z(n1335) );
  AND U1449 ( .A(o[1]), .B(\stack[1][2] ), .Z(n1334) );
  NAND U1450 ( .A(\stack[1][1] ), .B(o[2]), .Z(n1490) );
  AND U1451 ( .A(o[0]), .B(\stack[1][2] ), .Z(n1485) );
  AND U1452 ( .A(o[1]), .B(\stack[1][1] ), .Z(n1484) );
  AND U1453 ( .A(n1485), .B(n1484), .Z(n1491) );
  XNOR U1454 ( .A(n1333), .B(n1332), .Z(n1342) );
  AND U1455 ( .A(n1335), .B(n1334), .Z(n1344) );
  AND U1456 ( .A(o[2]), .B(\stack[1][2] ), .Z(n1343) );
  XNOR U1457 ( .A(n1344), .B(n1343), .Z(n1336) );
  XOR U1458 ( .A(n1342), .B(n1336), .Z(n1499) );
  AND U1459 ( .A(\stack[1][1] ), .B(o[3]), .Z(n1497) );
  AND U1460 ( .A(\stack[1][1] ), .B(o[4]), .Z(n1507) );
  IV U1461 ( .A(n1507), .Z(n1337) );
  NANDN U1462 ( .A(n1506), .B(n1337), .Z(n1348) );
  AND U1463 ( .A(n1506), .B(n1507), .Z(n1346) );
  XNOR U1464 ( .A(n1339), .B(n1338), .Z(n1340) );
  XNOR U1465 ( .A(n1341), .B(n1340), .Z(n1354) );
  IV U1466 ( .A(n1354), .Z(n1355) );
  AND U1467 ( .A(\stack[1][2] ), .B(o[3]), .Z(n1358) );
  XNOR U1468 ( .A(n1358), .B(n1356), .Z(n1345) );
  XNOR U1469 ( .A(n1355), .B(n1345), .Z(n1509) );
  OR U1470 ( .A(n1346), .B(n1509), .Z(n1347) );
  AND U1471 ( .A(n1348), .B(n1347), .Z(n1512) );
  IV U1472 ( .A(n1349), .Z(n1351) );
  XNOR U1473 ( .A(n1351), .B(n1350), .Z(n1352) );
  XOR U1474 ( .A(n1353), .B(n1352), .Z(n1369) );
  AND U1475 ( .A(\stack[1][2] ), .B(o[4]), .Z(n1367) );
  NANDN U1476 ( .A(n1356), .B(n1354), .Z(n1360) );
  AND U1477 ( .A(n1356), .B(n1355), .Z(n1357) );
  OR U1478 ( .A(n1358), .B(n1357), .Z(n1359) );
  AND U1479 ( .A(n1360), .B(n1359), .Z(n1368) );
  XNOR U1480 ( .A(n1367), .B(n1368), .Z(n1361) );
  XNOR U1481 ( .A(n1369), .B(n1361), .Z(n1362) );
  IV U1482 ( .A(n1362), .Z(n1515) );
  NANDN U1483 ( .A(n1512), .B(n1515), .Z(n1365) );
  AND U1484 ( .A(\stack[1][1] ), .B(o[5]), .Z(n1513) );
  AND U1485 ( .A(n1512), .B(n1362), .Z(n1363) );
  OR U1486 ( .A(n1513), .B(n1363), .Z(n1364) );
  AND U1487 ( .A(n1365), .B(n1364), .Z(n1522) );
  AND U1488 ( .A(\stack[1][1] ), .B(o[6]), .Z(n1378) );
  IV U1489 ( .A(n1378), .Z(n1525) );
  NANDN U1490 ( .A(n1522), .B(n1525), .Z(n1381) );
  IV U1491 ( .A(n1367), .Z(n1366) );
  NANDN U1492 ( .A(n1368), .B(n1366), .Z(n1372) );
  AND U1493 ( .A(n1368), .B(n1367), .Z(n1370) );
  OR U1494 ( .A(n1370), .B(n1369), .Z(n1371) );
  AND U1495 ( .A(n1372), .B(n1371), .Z(n1388) );
  AND U1496 ( .A(\stack[1][2] ), .B(o[5]), .Z(n1386) );
  XNOR U1497 ( .A(n1374), .B(n1373), .Z(n1375) );
  XNOR U1498 ( .A(n1376), .B(n1375), .Z(n1387) );
  IV U1499 ( .A(n1387), .Z(n1377) );
  XNOR U1500 ( .A(n1386), .B(n1377), .Z(n1389) );
  XOR U1501 ( .A(n1388), .B(n1389), .Z(n1523) );
  AND U1502 ( .A(n1522), .B(n1378), .Z(n1379) );
  OR U1503 ( .A(n1523), .B(n1379), .Z(n1380) );
  AND U1504 ( .A(n1381), .B(n1380), .Z(n1528) );
  XNOR U1505 ( .A(n1383), .B(n1382), .Z(n1384) );
  XNOR U1506 ( .A(n1385), .B(n1384), .Z(n1401) );
  NAND U1507 ( .A(n1387), .B(n1386), .Z(n1391) );
  NAND U1508 ( .A(n1389), .B(n1388), .Z(n1390) );
  NAND U1509 ( .A(n1391), .B(n1390), .Z(n1399) );
  IV U1510 ( .A(n1399), .Z(n1398) );
  AND U1511 ( .A(\stack[1][2] ), .B(o[6]), .Z(n1400) );
  XNOR U1512 ( .A(n1398), .B(n1400), .Z(n1392) );
  XOR U1513 ( .A(n1401), .B(n1392), .Z(n1531) );
  AND U1514 ( .A(\stack[1][1] ), .B(o[7]), .Z(n1529) );
  AND U1515 ( .A(\stack[1][1] ), .B(o[8]), .Z(n1539) );
  IV U1516 ( .A(n1539), .Z(n1393) );
  NANDN U1517 ( .A(n1538), .B(n1393), .Z(n1408) );
  AND U1518 ( .A(n1538), .B(n1539), .Z(n1406) );
  XNOR U1519 ( .A(n1395), .B(n1394), .Z(n1396) );
  XOR U1520 ( .A(n1397), .B(n1396), .Z(n1413) );
  IV U1521 ( .A(n1413), .Z(n1414) );
  AND U1522 ( .A(\stack[1][2] ), .B(o[7]), .Z(n1417) );
  NANDN U1523 ( .A(n1400), .B(n1398), .Z(n1404) );
  AND U1524 ( .A(n1400), .B(n1399), .Z(n1402) );
  OR U1525 ( .A(n1402), .B(n1401), .Z(n1403) );
  AND U1526 ( .A(n1404), .B(n1403), .Z(n1415) );
  XNOR U1527 ( .A(n1417), .B(n1415), .Z(n1405) );
  XNOR U1528 ( .A(n1414), .B(n1405), .Z(n1541) );
  OR U1529 ( .A(n1406), .B(n1541), .Z(n1407) );
  AND U1530 ( .A(n1408), .B(n1407), .Z(n1544) );
  XNOR U1531 ( .A(n1410), .B(n1409), .Z(n1411) );
  XNOR U1532 ( .A(n1412), .B(n1411), .Z(n1433) );
  AND U1533 ( .A(\stack[1][2] ), .B(o[8]), .Z(n1431) );
  NANDN U1534 ( .A(n1415), .B(n1413), .Z(n1419) );
  AND U1535 ( .A(n1415), .B(n1414), .Z(n1416) );
  OR U1536 ( .A(n1417), .B(n1416), .Z(n1418) );
  AND U1537 ( .A(n1419), .B(n1418), .Z(n1432) );
  XNOR U1538 ( .A(n1431), .B(n1432), .Z(n1420) );
  XNOR U1539 ( .A(n1433), .B(n1420), .Z(n1421) );
  IV U1540 ( .A(n1421), .Z(n1547) );
  NANDN U1541 ( .A(n1544), .B(n1547), .Z(n1424) );
  AND U1542 ( .A(\stack[1][1] ), .B(o[9]), .Z(n1545) );
  AND U1543 ( .A(n1544), .B(n1421), .Z(n1422) );
  OR U1544 ( .A(n1545), .B(n1422), .Z(n1423) );
  AND U1545 ( .A(n1424), .B(n1423), .Z(n1555) );
  AND U1546 ( .A(\stack[1][1] ), .B(o[10]), .Z(n1556) );
  IV U1547 ( .A(n1556), .Z(n1425) );
  NANDN U1548 ( .A(n1555), .B(n1425), .Z(n1440) );
  AND U1549 ( .A(n1555), .B(n1556), .Z(n1438) );
  XNOR U1550 ( .A(n1427), .B(n1426), .Z(n1428) );
  XNOR U1551 ( .A(n1429), .B(n1428), .Z(n1446) );
  AND U1552 ( .A(\stack[1][2] ), .B(o[9]), .Z(n1449) );
  IV U1553 ( .A(n1431), .Z(n1430) );
  NANDN U1554 ( .A(n1432), .B(n1430), .Z(n1436) );
  AND U1555 ( .A(n1432), .B(n1431), .Z(n1434) );
  OR U1556 ( .A(n1434), .B(n1433), .Z(n1435) );
  AND U1557 ( .A(n1436), .B(n1435), .Z(n1447) );
  XNOR U1558 ( .A(n1449), .B(n1447), .Z(n1437) );
  XNOR U1559 ( .A(n1446), .B(n1437), .Z(n1558) );
  OR U1560 ( .A(n1438), .B(n1558), .Z(n1439) );
  AND U1561 ( .A(n1440), .B(n1439), .Z(n1561) );
  XNOR U1562 ( .A(n1442), .B(n1441), .Z(n1443) );
  XNOR U1563 ( .A(n1444), .B(n1443), .Z(n1464) );
  AND U1564 ( .A(\stack[1][2] ), .B(o[10]), .Z(n1462) );
  IV U1565 ( .A(n1446), .Z(n1445) );
  NANDN U1566 ( .A(n1447), .B(n1445), .Z(n1451) );
  AND U1567 ( .A(n1447), .B(n1446), .Z(n1448) );
  OR U1568 ( .A(n1449), .B(n1448), .Z(n1450) );
  AND U1569 ( .A(n1451), .B(n1450), .Z(n1463) );
  XNOR U1570 ( .A(n1462), .B(n1463), .Z(n1452) );
  XNOR U1571 ( .A(n1464), .B(n1452), .Z(n1453) );
  IV U1572 ( .A(n1453), .Z(n1564) );
  NANDN U1573 ( .A(n1561), .B(n1564), .Z(n1456) );
  AND U1574 ( .A(\stack[1][1] ), .B(o[11]), .Z(n1562) );
  AND U1575 ( .A(n1561), .B(n1453), .Z(n1454) );
  OR U1576 ( .A(n1562), .B(n1454), .Z(n1455) );
  AND U1577 ( .A(n1456), .B(n1455), .Z(n1572) );
  AND U1578 ( .A(\stack[1][1] ), .B(o[12]), .Z(n1573) );
  XNOR U1579 ( .A(n1458), .B(n1457), .Z(n1459) );
  XNOR U1580 ( .A(n1460), .B(n1459), .Z(n1473) );
  AND U1581 ( .A(\stack[1][2] ), .B(o[11]), .Z(n1475) );
  IV U1582 ( .A(n1462), .Z(n1461) );
  NANDN U1583 ( .A(n1463), .B(n1461), .Z(n1467) );
  AND U1584 ( .A(n1463), .B(n1462), .Z(n1465) );
  OR U1585 ( .A(n1465), .B(n1464), .Z(n1466) );
  AND U1586 ( .A(n1467), .B(n1466), .Z(n1474) );
  XNOR U1587 ( .A(n1475), .B(n1474), .Z(n1468) );
  XNOR U1588 ( .A(n1473), .B(n1468), .Z(n1575) );
  XNOR U1589 ( .A(n1470), .B(n1469), .Z(n1471) );
  XNOR U1590 ( .A(n1472), .B(n1471), .Z(n1479) );
  AND U1591 ( .A(\stack[1][2] ), .B(o[12]), .Z(n1477) );
  IV U1592 ( .A(n1476), .Z(n1581) );
  AND U1593 ( .A(\stack[1][1] ), .B(o[13]), .Z(n1579) );
  XNOR U1594 ( .A(n1481), .B(n1480), .Z(n1587) );
  AND U1595 ( .A(\stack[1][0] ), .B(o[1]), .Z(n2127) );
  AND U1596 ( .A(o[0]), .B(\stack[1][1] ), .Z(n2131) );
  NAND U1597 ( .A(n2127), .B(n2131), .Z(n1482) );
  NAND U1598 ( .A(\stack[1][0] ), .B(o[2]), .Z(n1483) );
  NAND U1599 ( .A(n1482), .B(n1483), .Z(n1487) );
  XNOR U1600 ( .A(n1485), .B(n1484), .Z(n2097) );
  NAND U1601 ( .A(n2096), .B(n2097), .Z(n1486) );
  NAND U1602 ( .A(n1487), .B(n1486), .Z(n1488) );
  NAND U1603 ( .A(\stack[1][0] ), .B(o[3]), .Z(n1489) );
  NAND U1604 ( .A(n1488), .B(n1489), .Z(n1495) );
  XOR U1605 ( .A(n1491), .B(n1490), .Z(n1492) );
  XOR U1606 ( .A(n1493), .B(n1492), .Z(n2059) );
  NAND U1607 ( .A(n2058), .B(n2059), .Z(n1494) );
  NAND U1608 ( .A(n1495), .B(n1494), .Z(n1502) );
  XNOR U1609 ( .A(n1497), .B(n1496), .Z(n1498) );
  XOR U1610 ( .A(n1499), .B(n1498), .Z(n1501) );
  XOR U1611 ( .A(n1502), .B(n1501), .Z(n2018) );
  NAND U1612 ( .A(o[4]), .B(\stack[1][0] ), .Z(n1500) );
  AND U1613 ( .A(n2018), .B(n1500), .Z(n2014) );
  NAND U1614 ( .A(n1502), .B(n1501), .Z(n1503) );
  NANDN U1615 ( .A(n2014), .B(n1503), .Z(n1504) );
  NAND U1616 ( .A(\stack[1][0] ), .B(o[5]), .Z(n1505) );
  NAND U1617 ( .A(n1504), .B(n1505), .Z(n1511) );
  XNOR U1618 ( .A(n1507), .B(n1506), .Z(n1508) );
  XOR U1619 ( .A(n1509), .B(n1508), .Z(n1982) );
  NAND U1620 ( .A(n1981), .B(n1982), .Z(n1510) );
  NAND U1621 ( .A(n1511), .B(n1510), .Z(n1518) );
  XNOR U1622 ( .A(n1513), .B(n1512), .Z(n1514) );
  XNOR U1623 ( .A(n1515), .B(n1514), .Z(n1517) );
  XOR U1624 ( .A(n1518), .B(n1517), .Z(n1941) );
  NAND U1625 ( .A(o[6]), .B(\stack[1][0] ), .Z(n1516) );
  AND U1626 ( .A(n1941), .B(n1516), .Z(n1937) );
  NAND U1627 ( .A(n1518), .B(n1517), .Z(n1519) );
  NANDN U1628 ( .A(n1937), .B(n1519), .Z(n1520) );
  NAND U1629 ( .A(\stack[1][0] ), .B(o[7]), .Z(n1521) );
  NAND U1630 ( .A(n1520), .B(n1521), .Z(n1527) );
  XNOR U1631 ( .A(n1523), .B(n1522), .Z(n1524) );
  XNOR U1632 ( .A(n1525), .B(n1524), .Z(n1905) );
  NAND U1633 ( .A(n1904), .B(n1905), .Z(n1526) );
  NAND U1634 ( .A(n1527), .B(n1526), .Z(n1534) );
  XNOR U1635 ( .A(n1529), .B(n1528), .Z(n1530) );
  XOR U1636 ( .A(n1531), .B(n1530), .Z(n1533) );
  XOR U1637 ( .A(n1534), .B(n1533), .Z(n1864) );
  NAND U1638 ( .A(o[8]), .B(\stack[1][0] ), .Z(n1532) );
  AND U1639 ( .A(n1864), .B(n1532), .Z(n1860) );
  NAND U1640 ( .A(n1534), .B(n1533), .Z(n1535) );
  NANDN U1641 ( .A(n1860), .B(n1535), .Z(n1536) );
  NAND U1642 ( .A(\stack[1][0] ), .B(o[9]), .Z(n1537) );
  NAND U1643 ( .A(n1536), .B(n1537), .Z(n1543) );
  XNOR U1644 ( .A(n1539), .B(n1538), .Z(n1540) );
  XOR U1645 ( .A(n1541), .B(n1540), .Z(n1828) );
  NAND U1646 ( .A(n1827), .B(n1828), .Z(n1542) );
  NAND U1647 ( .A(n1543), .B(n1542), .Z(n1550) );
  XNOR U1648 ( .A(n1545), .B(n1544), .Z(n1546) );
  XNOR U1649 ( .A(n1547), .B(n1546), .Z(n1549) );
  XOR U1650 ( .A(n1550), .B(n1549), .Z(n1787) );
  NAND U1651 ( .A(o[10]), .B(\stack[1][0] ), .Z(n1548) );
  AND U1652 ( .A(n1787), .B(n1548), .Z(n1783) );
  NAND U1653 ( .A(n1550), .B(n1549), .Z(n1551) );
  NANDN U1654 ( .A(n1783), .B(n1551), .Z(n1552) );
  NAND U1655 ( .A(\stack[1][0] ), .B(o[11]), .Z(n1553) );
  NAND U1656 ( .A(n1552), .B(n1553), .Z(n1560) );
  IV U1657 ( .A(n1552), .Z(n1554) );
  XNOR U1658 ( .A(n1554), .B(n1553), .Z(n1750) );
  XNOR U1659 ( .A(n1556), .B(n1555), .Z(n1557) );
  XOR U1660 ( .A(n1558), .B(n1557), .Z(n1751) );
  NAND U1661 ( .A(n1750), .B(n1751), .Z(n1559) );
  NAND U1662 ( .A(n1560), .B(n1559), .Z(n1567) );
  XNOR U1663 ( .A(n1562), .B(n1561), .Z(n1563) );
  XNOR U1664 ( .A(n1564), .B(n1563), .Z(n1566) );
  XOR U1665 ( .A(n1567), .B(n1566), .Z(n1710) );
  NAND U1666 ( .A(o[12]), .B(\stack[1][0] ), .Z(n1565) );
  AND U1667 ( .A(n1710), .B(n1565), .Z(n1706) );
  NAND U1668 ( .A(n1567), .B(n1566), .Z(n1568) );
  NANDN U1669 ( .A(n1706), .B(n1568), .Z(n1569) );
  NAND U1670 ( .A(\stack[1][0] ), .B(o[13]), .Z(n1570) );
  NAND U1671 ( .A(n1569), .B(n1570), .Z(n1577) );
  IV U1672 ( .A(n1569), .Z(n1571) );
  XNOR U1673 ( .A(n1571), .B(n1570), .Z(n1673) );
  XNOR U1674 ( .A(n1573), .B(n1572), .Z(n1574) );
  XOR U1675 ( .A(n1575), .B(n1574), .Z(n1674) );
  NAND U1676 ( .A(n1673), .B(n1674), .Z(n1576) );
  NAND U1677 ( .A(n1577), .B(n1576), .Z(n1584) );
  XNOR U1678 ( .A(n1579), .B(n1578), .Z(n1580) );
  XNOR U1679 ( .A(n1581), .B(n1580), .Z(n1583) );
  XOR U1680 ( .A(n1584), .B(n1583), .Z(n1633) );
  NAND U1681 ( .A(o[14]), .B(\stack[1][0] ), .Z(n1582) );
  AND U1682 ( .A(n1633), .B(n1582), .Z(n1629) );
  AND U1683 ( .A(n1584), .B(n1583), .Z(n1585) );
  OR U1684 ( .A(n1629), .B(n1585), .Z(n1586) );
  XNOR U1685 ( .A(n1587), .B(n1586), .Z(n1588) );
  NANDN U1686 ( .A(n2151), .B(n1588), .Z(n1591) );
  AND U1687 ( .A(opcode[2]), .B(n1589), .Z(n2154) );
  NAND U1688 ( .A(n2154), .B(\stack[1][15] ), .Z(n1590) );
  AND U1689 ( .A(n1591), .B(n1590), .Z(n1592) );
  NANDN U1690 ( .A(n1593), .B(n1592), .Z(n1600) );
  XNOR U1691 ( .A(opcode[0]), .B(opcode[2]), .Z(n1595) );
  XNOR U1692 ( .A(opcode[2]), .B(opcode[1]), .Z(n1594) );
  NAND U1693 ( .A(n1595), .B(n1594), .Z(n2148) );
  AND U1694 ( .A(opcode[2]), .B(opcode[1]), .Z(n2152) );
  NAND U1695 ( .A(\stack[1][15] ), .B(n2152), .Z(n1596) );
  NAND U1696 ( .A(n2148), .B(n1596), .Z(n1597) );
  AND U1697 ( .A(o[15]), .B(n1597), .Z(n1598) );
  NANDN U1698 ( .A(n1600), .B(n1599), .Z(n566) );
  NAND U1699 ( .A(\stack[6][14] ), .B(n2150), .Z(n1602) );
  NANDN U1700 ( .A(n2150), .B(\stack[7][14] ), .Z(n1601) );
  NAND U1701 ( .A(n1602), .B(n1601), .Z(n567) );
  NAND U1702 ( .A(\stack[5][14] ), .B(n2150), .Z(n1604) );
  NANDN U1703 ( .A(n2142), .B(\stack[7][14] ), .Z(n1603) );
  AND U1704 ( .A(n1604), .B(n1603), .Z(n1606) );
  NAND U1705 ( .A(n2145), .B(\stack[6][14] ), .Z(n1605) );
  NAND U1706 ( .A(n1606), .B(n1605), .Z(n568) );
  NAND U1707 ( .A(\stack[4][14] ), .B(n2150), .Z(n1608) );
  NANDN U1708 ( .A(n2142), .B(\stack[6][14] ), .Z(n1607) );
  AND U1709 ( .A(n1608), .B(n1607), .Z(n1610) );
  NAND U1710 ( .A(n2145), .B(\stack[5][14] ), .Z(n1609) );
  NAND U1711 ( .A(n1610), .B(n1609), .Z(n569) );
  NAND U1712 ( .A(\stack[3][14] ), .B(n2150), .Z(n1612) );
  NANDN U1713 ( .A(n2142), .B(\stack[5][14] ), .Z(n1611) );
  AND U1714 ( .A(n1612), .B(n1611), .Z(n1614) );
  NAND U1715 ( .A(n2145), .B(\stack[4][14] ), .Z(n1613) );
  NAND U1716 ( .A(n1614), .B(n1613), .Z(n570) );
  NAND U1717 ( .A(\stack[2][14] ), .B(n2150), .Z(n1616) );
  NANDN U1718 ( .A(n2142), .B(\stack[4][14] ), .Z(n1615) );
  AND U1719 ( .A(n1616), .B(n1615), .Z(n1618) );
  NAND U1720 ( .A(n2145), .B(\stack[3][14] ), .Z(n1617) );
  NAND U1721 ( .A(n1618), .B(n1617), .Z(n571) );
  NAND U1722 ( .A(n2150), .B(\stack[1][14] ), .Z(n1620) );
  NANDN U1723 ( .A(n2142), .B(\stack[3][14] ), .Z(n1619) );
  AND U1724 ( .A(n1620), .B(n1619), .Z(n1622) );
  NAND U1725 ( .A(n2145), .B(\stack[2][14] ), .Z(n1621) );
  NAND U1726 ( .A(n1622), .B(n1621), .Z(n572) );
  NAND U1727 ( .A(n2150), .B(o[14]), .Z(n1624) );
  NANDN U1728 ( .A(n2142), .B(\stack[2][14] ), .Z(n1623) );
  AND U1729 ( .A(n1624), .B(n1623), .Z(n1626) );
  NAND U1730 ( .A(\stack[1][14] ), .B(n2145), .Z(n1625) );
  NAND U1731 ( .A(n1626), .B(n1625), .Z(n573) );
  NAND U1732 ( .A(x[14]), .B(n2150), .Z(n1628) );
  NAND U1733 ( .A(\stack[1][14] ), .B(n2154), .Z(n1627) );
  NAND U1734 ( .A(n1628), .B(n1627), .Z(n1632) );
  ANDN U1735 ( .B(n1629), .A(n2151), .Z(n1630) );
  NANDN U1736 ( .A(n1632), .B(n1631), .Z(n1639) );
  NANDN U1737 ( .A(n2151), .B(\stack[1][0] ), .Z(n2132) );
  OR U1738 ( .A(n2132), .B(n1633), .Z(n1635) );
  NAND U1739 ( .A(\stack[1][14] ), .B(n2152), .Z(n1634) );
  AND U1740 ( .A(n1635), .B(n1634), .Z(n1636) );
  NAND U1741 ( .A(n2148), .B(n1636), .Z(n1637) );
  NAND U1742 ( .A(o[14]), .B(n1637), .Z(n1638) );
  NANDN U1743 ( .A(n1639), .B(n1638), .Z(n574) );
  NAND U1744 ( .A(\stack[6][13] ), .B(n2150), .Z(n1641) );
  NANDN U1745 ( .A(n2150), .B(\stack[7][13] ), .Z(n1640) );
  NAND U1746 ( .A(n1641), .B(n1640), .Z(n575) );
  NAND U1747 ( .A(\stack[5][13] ), .B(n2150), .Z(n1643) );
  NANDN U1748 ( .A(n2142), .B(\stack[7][13] ), .Z(n1642) );
  AND U1749 ( .A(n1643), .B(n1642), .Z(n1645) );
  NAND U1750 ( .A(n2145), .B(\stack[6][13] ), .Z(n1644) );
  NAND U1751 ( .A(n1645), .B(n1644), .Z(n576) );
  NAND U1752 ( .A(\stack[4][13] ), .B(n2150), .Z(n1647) );
  NANDN U1753 ( .A(n2142), .B(\stack[6][13] ), .Z(n1646) );
  AND U1754 ( .A(n1647), .B(n1646), .Z(n1649) );
  NAND U1755 ( .A(n2145), .B(\stack[5][13] ), .Z(n1648) );
  NAND U1756 ( .A(n1649), .B(n1648), .Z(n577) );
  NAND U1757 ( .A(\stack[3][13] ), .B(n2150), .Z(n1651) );
  NANDN U1758 ( .A(n2142), .B(\stack[5][13] ), .Z(n1650) );
  AND U1759 ( .A(n1651), .B(n1650), .Z(n1653) );
  NAND U1760 ( .A(n2145), .B(\stack[4][13] ), .Z(n1652) );
  NAND U1761 ( .A(n1653), .B(n1652), .Z(n578) );
  NAND U1762 ( .A(\stack[2][13] ), .B(n2150), .Z(n1655) );
  NANDN U1763 ( .A(n2142), .B(\stack[4][13] ), .Z(n1654) );
  AND U1764 ( .A(n1655), .B(n1654), .Z(n1657) );
  NAND U1765 ( .A(n2145), .B(\stack[3][13] ), .Z(n1656) );
  NAND U1766 ( .A(n1657), .B(n1656), .Z(n579) );
  NAND U1767 ( .A(n2150), .B(\stack[1][13] ), .Z(n1659) );
  NANDN U1768 ( .A(n2142), .B(\stack[3][13] ), .Z(n1658) );
  AND U1769 ( .A(n1659), .B(n1658), .Z(n1661) );
  NAND U1770 ( .A(n2145), .B(\stack[2][13] ), .Z(n1660) );
  NAND U1771 ( .A(n1661), .B(n1660), .Z(n580) );
  NAND U1772 ( .A(n2150), .B(o[13]), .Z(n1663) );
  NANDN U1773 ( .A(n2142), .B(\stack[2][13] ), .Z(n1662) );
  AND U1774 ( .A(n1663), .B(n1662), .Z(n1665) );
  NAND U1775 ( .A(\stack[1][13] ), .B(n2145), .Z(n1664) );
  NAND U1776 ( .A(n1665), .B(n1664), .Z(n581) );
  NAND U1777 ( .A(\stack[1][13] ), .B(n2152), .Z(n1666) );
  NAND U1778 ( .A(n2148), .B(n1666), .Z(n1667) );
  NAND U1779 ( .A(o[13]), .B(n1667), .Z(n1671) );
  NAND U1780 ( .A(x[13]), .B(n2150), .Z(n1669) );
  NAND U1781 ( .A(\stack[1][13] ), .B(n2154), .Z(n1668) );
  AND U1782 ( .A(n1669), .B(n1668), .Z(n1670) );
  AND U1783 ( .A(n1671), .B(n1670), .Z(n1672) );
  XNOR U1784 ( .A(n1674), .B(n1673), .Z(n1675) );
  NANDN U1785 ( .A(n2151), .B(n1675), .Z(n1676) );
  NAND U1786 ( .A(n1677), .B(n1676), .Z(n582) );
  NAND U1787 ( .A(\stack[6][12] ), .B(n2150), .Z(n1679) );
  NANDN U1788 ( .A(n2150), .B(\stack[7][12] ), .Z(n1678) );
  NAND U1789 ( .A(n1679), .B(n1678), .Z(n583) );
  NAND U1790 ( .A(\stack[5][12] ), .B(n2150), .Z(n1681) );
  NANDN U1791 ( .A(n2142), .B(\stack[7][12] ), .Z(n1680) );
  AND U1792 ( .A(n1681), .B(n1680), .Z(n1683) );
  NAND U1793 ( .A(n2145), .B(\stack[6][12] ), .Z(n1682) );
  NAND U1794 ( .A(n1683), .B(n1682), .Z(n584) );
  NAND U1795 ( .A(\stack[4][12] ), .B(n2150), .Z(n1685) );
  NANDN U1796 ( .A(n2142), .B(\stack[6][12] ), .Z(n1684) );
  AND U1797 ( .A(n1685), .B(n1684), .Z(n1687) );
  NAND U1798 ( .A(n2145), .B(\stack[5][12] ), .Z(n1686) );
  NAND U1799 ( .A(n1687), .B(n1686), .Z(n585) );
  NAND U1800 ( .A(\stack[3][12] ), .B(n2150), .Z(n1689) );
  NANDN U1801 ( .A(n2142), .B(\stack[5][12] ), .Z(n1688) );
  AND U1802 ( .A(n1689), .B(n1688), .Z(n1691) );
  NAND U1803 ( .A(n2145), .B(\stack[4][12] ), .Z(n1690) );
  NAND U1804 ( .A(n1691), .B(n1690), .Z(n586) );
  NAND U1805 ( .A(\stack[2][12] ), .B(n2150), .Z(n1693) );
  NANDN U1806 ( .A(n2142), .B(\stack[4][12] ), .Z(n1692) );
  AND U1807 ( .A(n1693), .B(n1692), .Z(n1695) );
  NAND U1808 ( .A(n2145), .B(\stack[3][12] ), .Z(n1694) );
  NAND U1809 ( .A(n1695), .B(n1694), .Z(n587) );
  NAND U1810 ( .A(n2150), .B(\stack[1][12] ), .Z(n1697) );
  NANDN U1811 ( .A(n2142), .B(\stack[3][12] ), .Z(n1696) );
  AND U1812 ( .A(n1697), .B(n1696), .Z(n1699) );
  NAND U1813 ( .A(n2145), .B(\stack[2][12] ), .Z(n1698) );
  NAND U1814 ( .A(n1699), .B(n1698), .Z(n588) );
  NAND U1815 ( .A(n2150), .B(o[12]), .Z(n1701) );
  NANDN U1816 ( .A(n2142), .B(\stack[2][12] ), .Z(n1700) );
  AND U1817 ( .A(n1701), .B(n1700), .Z(n1703) );
  NAND U1818 ( .A(\stack[1][12] ), .B(n2145), .Z(n1702) );
  NAND U1819 ( .A(n1703), .B(n1702), .Z(n589) );
  NAND U1820 ( .A(x[12]), .B(n2150), .Z(n1705) );
  NAND U1821 ( .A(\stack[1][12] ), .B(n2154), .Z(n1704) );
  NAND U1822 ( .A(n1705), .B(n1704), .Z(n1709) );
  ANDN U1823 ( .B(n1706), .A(n2151), .Z(n1707) );
  NANDN U1824 ( .A(n1709), .B(n1708), .Z(n1716) );
  OR U1825 ( .A(n2132), .B(n1710), .Z(n1712) );
  NAND U1826 ( .A(\stack[1][12] ), .B(n2152), .Z(n1711) );
  AND U1827 ( .A(n1712), .B(n1711), .Z(n1713) );
  NAND U1828 ( .A(n2148), .B(n1713), .Z(n1714) );
  NAND U1829 ( .A(o[12]), .B(n1714), .Z(n1715) );
  NANDN U1830 ( .A(n1716), .B(n1715), .Z(n590) );
  NAND U1831 ( .A(\stack[6][11] ), .B(n2150), .Z(n1718) );
  NANDN U1832 ( .A(n2150), .B(\stack[7][11] ), .Z(n1717) );
  NAND U1833 ( .A(n1718), .B(n1717), .Z(n591) );
  NAND U1834 ( .A(\stack[5][11] ), .B(n2150), .Z(n1720) );
  NANDN U1835 ( .A(n2142), .B(\stack[7][11] ), .Z(n1719) );
  AND U1836 ( .A(n1720), .B(n1719), .Z(n1722) );
  NAND U1837 ( .A(n2145), .B(\stack[6][11] ), .Z(n1721) );
  NAND U1838 ( .A(n1722), .B(n1721), .Z(n592) );
  NAND U1839 ( .A(\stack[4][11] ), .B(n2150), .Z(n1724) );
  NANDN U1840 ( .A(n2142), .B(\stack[6][11] ), .Z(n1723) );
  AND U1841 ( .A(n1724), .B(n1723), .Z(n1726) );
  NAND U1842 ( .A(n2145), .B(\stack[5][11] ), .Z(n1725) );
  NAND U1843 ( .A(n1726), .B(n1725), .Z(n593) );
  NAND U1844 ( .A(\stack[3][11] ), .B(n2150), .Z(n1728) );
  NANDN U1845 ( .A(n2142), .B(\stack[5][11] ), .Z(n1727) );
  AND U1846 ( .A(n1728), .B(n1727), .Z(n1730) );
  NAND U1847 ( .A(n2145), .B(\stack[4][11] ), .Z(n1729) );
  NAND U1848 ( .A(n1730), .B(n1729), .Z(n594) );
  NAND U1849 ( .A(\stack[2][11] ), .B(n2150), .Z(n1732) );
  NANDN U1850 ( .A(n2142), .B(\stack[4][11] ), .Z(n1731) );
  AND U1851 ( .A(n1732), .B(n1731), .Z(n1734) );
  NAND U1852 ( .A(n2145), .B(\stack[3][11] ), .Z(n1733) );
  NAND U1853 ( .A(n1734), .B(n1733), .Z(n595) );
  NAND U1854 ( .A(n2150), .B(\stack[1][11] ), .Z(n1736) );
  NANDN U1855 ( .A(n2142), .B(\stack[3][11] ), .Z(n1735) );
  AND U1856 ( .A(n1736), .B(n1735), .Z(n1738) );
  NAND U1857 ( .A(n2145), .B(\stack[2][11] ), .Z(n1737) );
  NAND U1858 ( .A(n1738), .B(n1737), .Z(n596) );
  NAND U1859 ( .A(n2150), .B(o[11]), .Z(n1740) );
  NANDN U1860 ( .A(n2142), .B(\stack[2][11] ), .Z(n1739) );
  AND U1861 ( .A(n1740), .B(n1739), .Z(n1742) );
  NAND U1862 ( .A(\stack[1][11] ), .B(n2145), .Z(n1741) );
  NAND U1863 ( .A(n1742), .B(n1741), .Z(n597) );
  NANDN U1864 ( .A(n2148), .B(o[11]), .Z(n1743) );
  NAND U1865 ( .A(o[11]), .B(n2152), .Z(n1744) );
  NANDN U1866 ( .A(n2154), .B(n1744), .Z(n1745) );
  AND U1867 ( .A(\stack[1][11] ), .B(n1745), .Z(n1746) );
  NOR U1868 ( .A(n1747), .B(n1746), .Z(n1749) );
  NAND U1869 ( .A(x[11]), .B(n2150), .Z(n1748) );
  AND U1870 ( .A(n1749), .B(n1748), .Z(n1754) );
  XNOR U1871 ( .A(n1751), .B(n1750), .Z(n1752) );
  NANDN U1872 ( .A(n2151), .B(n1752), .Z(n1753) );
  NAND U1873 ( .A(n1754), .B(n1753), .Z(n598) );
  NAND U1874 ( .A(\stack[6][10] ), .B(n2150), .Z(n1756) );
  NANDN U1875 ( .A(n2150), .B(\stack[7][10] ), .Z(n1755) );
  NAND U1876 ( .A(n1756), .B(n1755), .Z(n599) );
  NAND U1877 ( .A(\stack[5][10] ), .B(n2150), .Z(n1758) );
  NANDN U1878 ( .A(n2142), .B(\stack[7][10] ), .Z(n1757) );
  AND U1879 ( .A(n1758), .B(n1757), .Z(n1760) );
  NAND U1880 ( .A(n2145), .B(\stack[6][10] ), .Z(n1759) );
  NAND U1881 ( .A(n1760), .B(n1759), .Z(n600) );
  NAND U1882 ( .A(\stack[4][10] ), .B(n2150), .Z(n1762) );
  NANDN U1883 ( .A(n2142), .B(\stack[6][10] ), .Z(n1761) );
  AND U1884 ( .A(n1762), .B(n1761), .Z(n1764) );
  NAND U1885 ( .A(n2145), .B(\stack[5][10] ), .Z(n1763) );
  NAND U1886 ( .A(n1764), .B(n1763), .Z(n601) );
  NAND U1887 ( .A(\stack[3][10] ), .B(n2150), .Z(n1766) );
  NANDN U1888 ( .A(n2142), .B(\stack[5][10] ), .Z(n1765) );
  AND U1889 ( .A(n1766), .B(n1765), .Z(n1768) );
  NAND U1890 ( .A(n2145), .B(\stack[4][10] ), .Z(n1767) );
  NAND U1891 ( .A(n1768), .B(n1767), .Z(n602) );
  NAND U1892 ( .A(\stack[2][10] ), .B(n2150), .Z(n1770) );
  NANDN U1893 ( .A(n2142), .B(\stack[4][10] ), .Z(n1769) );
  AND U1894 ( .A(n1770), .B(n1769), .Z(n1772) );
  NAND U1895 ( .A(n2145), .B(\stack[3][10] ), .Z(n1771) );
  NAND U1896 ( .A(n1772), .B(n1771), .Z(n603) );
  NAND U1897 ( .A(n2150), .B(\stack[1][10] ), .Z(n1774) );
  NANDN U1898 ( .A(n2142), .B(\stack[3][10] ), .Z(n1773) );
  AND U1899 ( .A(n1774), .B(n1773), .Z(n1776) );
  NAND U1900 ( .A(n2145), .B(\stack[2][10] ), .Z(n1775) );
  NAND U1901 ( .A(n1776), .B(n1775), .Z(n604) );
  NAND U1902 ( .A(n2150), .B(o[10]), .Z(n1778) );
  NANDN U1903 ( .A(n2142), .B(\stack[2][10] ), .Z(n1777) );
  AND U1904 ( .A(n1778), .B(n1777), .Z(n1780) );
  NAND U1905 ( .A(\stack[1][10] ), .B(n2145), .Z(n1779) );
  NAND U1906 ( .A(n1780), .B(n1779), .Z(n605) );
  NAND U1907 ( .A(x[10]), .B(n2150), .Z(n1782) );
  NAND U1908 ( .A(\stack[1][10] ), .B(n2154), .Z(n1781) );
  NAND U1909 ( .A(n1782), .B(n1781), .Z(n1786) );
  ANDN U1910 ( .B(n1783), .A(n2151), .Z(n1784) );
  NANDN U1911 ( .A(n1786), .B(n1785), .Z(n1793) );
  OR U1912 ( .A(n2132), .B(n1787), .Z(n1789) );
  NAND U1913 ( .A(\stack[1][10] ), .B(n2152), .Z(n1788) );
  AND U1914 ( .A(n1789), .B(n1788), .Z(n1790) );
  NAND U1915 ( .A(n2148), .B(n1790), .Z(n1791) );
  NAND U1916 ( .A(o[10]), .B(n1791), .Z(n1792) );
  NANDN U1917 ( .A(n1793), .B(n1792), .Z(n606) );
  NAND U1918 ( .A(\stack[6][9] ), .B(n2150), .Z(n1795) );
  NANDN U1919 ( .A(n2150), .B(\stack[7][9] ), .Z(n1794) );
  NAND U1920 ( .A(n1795), .B(n1794), .Z(n607) );
  NAND U1921 ( .A(\stack[5][9] ), .B(n2150), .Z(n1797) );
  NANDN U1922 ( .A(n2142), .B(\stack[7][9] ), .Z(n1796) );
  AND U1923 ( .A(n1797), .B(n1796), .Z(n1799) );
  NAND U1924 ( .A(n2145), .B(\stack[6][9] ), .Z(n1798) );
  NAND U1925 ( .A(n1799), .B(n1798), .Z(n608) );
  NAND U1926 ( .A(\stack[4][9] ), .B(n2150), .Z(n1801) );
  NANDN U1927 ( .A(n2142), .B(\stack[6][9] ), .Z(n1800) );
  AND U1928 ( .A(n1801), .B(n1800), .Z(n1803) );
  NAND U1929 ( .A(n2145), .B(\stack[5][9] ), .Z(n1802) );
  NAND U1930 ( .A(n1803), .B(n1802), .Z(n609) );
  NAND U1931 ( .A(\stack[3][9] ), .B(n2150), .Z(n1805) );
  NANDN U1932 ( .A(n2142), .B(\stack[5][9] ), .Z(n1804) );
  AND U1933 ( .A(n1805), .B(n1804), .Z(n1807) );
  NAND U1934 ( .A(n2145), .B(\stack[4][9] ), .Z(n1806) );
  NAND U1935 ( .A(n1807), .B(n1806), .Z(n610) );
  NAND U1936 ( .A(\stack[2][9] ), .B(n2150), .Z(n1809) );
  NANDN U1937 ( .A(n2142), .B(\stack[4][9] ), .Z(n1808) );
  AND U1938 ( .A(n1809), .B(n1808), .Z(n1811) );
  NAND U1939 ( .A(n2145), .B(\stack[3][9] ), .Z(n1810) );
  NAND U1940 ( .A(n1811), .B(n1810), .Z(n611) );
  NAND U1941 ( .A(n2150), .B(\stack[1][9] ), .Z(n1813) );
  NANDN U1942 ( .A(n2142), .B(\stack[3][9] ), .Z(n1812) );
  AND U1943 ( .A(n1813), .B(n1812), .Z(n1815) );
  NAND U1944 ( .A(n2145), .B(\stack[2][9] ), .Z(n1814) );
  NAND U1945 ( .A(n1815), .B(n1814), .Z(n612) );
  NAND U1946 ( .A(n2150), .B(o[9]), .Z(n1817) );
  NANDN U1947 ( .A(n2142), .B(\stack[2][9] ), .Z(n1816) );
  AND U1948 ( .A(n1817), .B(n1816), .Z(n1819) );
  NAND U1949 ( .A(\stack[1][9] ), .B(n2145), .Z(n1818) );
  NAND U1950 ( .A(n1819), .B(n1818), .Z(n613) );
  NAND U1951 ( .A(\stack[1][9] ), .B(n2152), .Z(n1820) );
  NAND U1952 ( .A(n2148), .B(n1820), .Z(n1821) );
  NAND U1953 ( .A(o[9]), .B(n1821), .Z(n1825) );
  NAND U1954 ( .A(x[9]), .B(n2150), .Z(n1823) );
  NAND U1955 ( .A(\stack[1][9] ), .B(n2154), .Z(n1822) );
  AND U1956 ( .A(n1823), .B(n1822), .Z(n1824) );
  AND U1957 ( .A(n1825), .B(n1824), .Z(n1826) );
  XNOR U1958 ( .A(n1828), .B(n1827), .Z(n1829) );
  NANDN U1959 ( .A(n2151), .B(n1829), .Z(n1830) );
  NAND U1960 ( .A(n1831), .B(n1830), .Z(n614) );
  NAND U1961 ( .A(\stack[6][8] ), .B(n2150), .Z(n1833) );
  NANDN U1962 ( .A(n2150), .B(\stack[7][8] ), .Z(n1832) );
  NAND U1963 ( .A(n1833), .B(n1832), .Z(n615) );
  NAND U1964 ( .A(\stack[5][8] ), .B(n2150), .Z(n1835) );
  NANDN U1965 ( .A(n2142), .B(\stack[7][8] ), .Z(n1834) );
  AND U1966 ( .A(n1835), .B(n1834), .Z(n1837) );
  NAND U1967 ( .A(n2145), .B(\stack[6][8] ), .Z(n1836) );
  NAND U1968 ( .A(n1837), .B(n1836), .Z(n616) );
  NAND U1969 ( .A(\stack[4][8] ), .B(n2150), .Z(n1839) );
  NANDN U1970 ( .A(n2142), .B(\stack[6][8] ), .Z(n1838) );
  AND U1971 ( .A(n1839), .B(n1838), .Z(n1841) );
  NAND U1972 ( .A(n2145), .B(\stack[5][8] ), .Z(n1840) );
  NAND U1973 ( .A(n1841), .B(n1840), .Z(n617) );
  NAND U1974 ( .A(\stack[3][8] ), .B(n2150), .Z(n1843) );
  NANDN U1975 ( .A(n2142), .B(\stack[5][8] ), .Z(n1842) );
  AND U1976 ( .A(n1843), .B(n1842), .Z(n1845) );
  NAND U1977 ( .A(n2145), .B(\stack[4][8] ), .Z(n1844) );
  NAND U1978 ( .A(n1845), .B(n1844), .Z(n618) );
  NAND U1979 ( .A(\stack[2][8] ), .B(n2150), .Z(n1847) );
  NANDN U1980 ( .A(n2142), .B(\stack[4][8] ), .Z(n1846) );
  AND U1981 ( .A(n1847), .B(n1846), .Z(n1849) );
  NAND U1982 ( .A(n2145), .B(\stack[3][8] ), .Z(n1848) );
  NAND U1983 ( .A(n1849), .B(n1848), .Z(n619) );
  NAND U1984 ( .A(n2150), .B(\stack[1][8] ), .Z(n1851) );
  NANDN U1985 ( .A(n2142), .B(\stack[3][8] ), .Z(n1850) );
  AND U1986 ( .A(n1851), .B(n1850), .Z(n1853) );
  NAND U1987 ( .A(n2145), .B(\stack[2][8] ), .Z(n1852) );
  NAND U1988 ( .A(n1853), .B(n1852), .Z(n620) );
  NAND U1989 ( .A(n2150), .B(o[8]), .Z(n1855) );
  NANDN U1990 ( .A(n2142), .B(\stack[2][8] ), .Z(n1854) );
  AND U1991 ( .A(n1855), .B(n1854), .Z(n1857) );
  NAND U1992 ( .A(\stack[1][8] ), .B(n2145), .Z(n1856) );
  NAND U1993 ( .A(n1857), .B(n1856), .Z(n621) );
  NAND U1994 ( .A(x[8]), .B(n2150), .Z(n1859) );
  NAND U1995 ( .A(\stack[1][8] ), .B(n2154), .Z(n1858) );
  NAND U1996 ( .A(n1859), .B(n1858), .Z(n1863) );
  ANDN U1997 ( .B(n1860), .A(n2151), .Z(n1861) );
  NANDN U1998 ( .A(n1863), .B(n1862), .Z(n1870) );
  OR U1999 ( .A(n2132), .B(n1864), .Z(n1866) );
  NAND U2000 ( .A(\stack[1][8] ), .B(n2152), .Z(n1865) );
  AND U2001 ( .A(n1866), .B(n1865), .Z(n1867) );
  NAND U2002 ( .A(n2148), .B(n1867), .Z(n1868) );
  NAND U2003 ( .A(o[8]), .B(n1868), .Z(n1869) );
  NANDN U2004 ( .A(n1870), .B(n1869), .Z(n622) );
  NAND U2005 ( .A(\stack[6][7] ), .B(n2150), .Z(n1872) );
  NANDN U2006 ( .A(n2150), .B(\stack[7][7] ), .Z(n1871) );
  NAND U2007 ( .A(n1872), .B(n1871), .Z(n623) );
  NAND U2008 ( .A(\stack[5][7] ), .B(n2150), .Z(n1874) );
  NANDN U2009 ( .A(n2142), .B(\stack[7][7] ), .Z(n1873) );
  AND U2010 ( .A(n1874), .B(n1873), .Z(n1876) );
  NAND U2011 ( .A(n2145), .B(\stack[6][7] ), .Z(n1875) );
  NAND U2012 ( .A(n1876), .B(n1875), .Z(n624) );
  NAND U2013 ( .A(\stack[4][7] ), .B(n2150), .Z(n1878) );
  NANDN U2014 ( .A(n2142), .B(\stack[6][7] ), .Z(n1877) );
  AND U2015 ( .A(n1878), .B(n1877), .Z(n1880) );
  NAND U2016 ( .A(n2145), .B(\stack[5][7] ), .Z(n1879) );
  NAND U2017 ( .A(n1880), .B(n1879), .Z(n625) );
  NAND U2018 ( .A(\stack[3][7] ), .B(n2150), .Z(n1882) );
  NANDN U2019 ( .A(n2142), .B(\stack[5][7] ), .Z(n1881) );
  AND U2020 ( .A(n1882), .B(n1881), .Z(n1884) );
  NAND U2021 ( .A(n2145), .B(\stack[4][7] ), .Z(n1883) );
  NAND U2022 ( .A(n1884), .B(n1883), .Z(n626) );
  NAND U2023 ( .A(\stack[2][7] ), .B(n2150), .Z(n1886) );
  NANDN U2024 ( .A(n2142), .B(\stack[4][7] ), .Z(n1885) );
  AND U2025 ( .A(n1886), .B(n1885), .Z(n1888) );
  NAND U2026 ( .A(n2145), .B(\stack[3][7] ), .Z(n1887) );
  NAND U2027 ( .A(n1888), .B(n1887), .Z(n627) );
  NAND U2028 ( .A(n2150), .B(\stack[1][7] ), .Z(n1890) );
  NANDN U2029 ( .A(n2142), .B(\stack[3][7] ), .Z(n1889) );
  AND U2030 ( .A(n1890), .B(n1889), .Z(n1892) );
  NAND U2031 ( .A(n2145), .B(\stack[2][7] ), .Z(n1891) );
  NAND U2032 ( .A(n1892), .B(n1891), .Z(n628) );
  NAND U2033 ( .A(n2150), .B(o[7]), .Z(n1894) );
  NANDN U2034 ( .A(n2142), .B(\stack[2][7] ), .Z(n1893) );
  AND U2035 ( .A(n1894), .B(n1893), .Z(n1896) );
  NAND U2036 ( .A(\stack[1][7] ), .B(n2145), .Z(n1895) );
  NAND U2037 ( .A(n1896), .B(n1895), .Z(n629) );
  NAND U2038 ( .A(o[7]), .B(n2152), .Z(n1897) );
  NANDN U2039 ( .A(n2154), .B(n1897), .Z(n1898) );
  NAND U2040 ( .A(\stack[1][7] ), .B(n1898), .Z(n1901) );
  NAND U2041 ( .A(x[7]), .B(n2150), .Z(n1899) );
  AND U2042 ( .A(n1901), .B(n1900), .Z(n1903) );
  NANDN U2043 ( .A(n2148), .B(o[7]), .Z(n1902) );
  AND U2044 ( .A(n1903), .B(n1902), .Z(n1908) );
  XNOR U2045 ( .A(n1905), .B(n1904), .Z(n1906) );
  NANDN U2046 ( .A(n2151), .B(n1906), .Z(n1907) );
  NAND U2047 ( .A(n1908), .B(n1907), .Z(n630) );
  NAND U2048 ( .A(\stack[6][6] ), .B(n2150), .Z(n1910) );
  NANDN U2049 ( .A(n2150), .B(\stack[7][6] ), .Z(n1909) );
  NAND U2050 ( .A(n1910), .B(n1909), .Z(n631) );
  NAND U2051 ( .A(\stack[5][6] ), .B(n2150), .Z(n1912) );
  NANDN U2052 ( .A(n2142), .B(\stack[7][6] ), .Z(n1911) );
  AND U2053 ( .A(n1912), .B(n1911), .Z(n1914) );
  NAND U2054 ( .A(n2145), .B(\stack[6][6] ), .Z(n1913) );
  NAND U2055 ( .A(n1914), .B(n1913), .Z(n632) );
  NAND U2056 ( .A(\stack[4][6] ), .B(n2150), .Z(n1916) );
  NANDN U2057 ( .A(n2142), .B(\stack[6][6] ), .Z(n1915) );
  AND U2058 ( .A(n1916), .B(n1915), .Z(n1918) );
  NAND U2059 ( .A(n2145), .B(\stack[5][6] ), .Z(n1917) );
  NAND U2060 ( .A(n1918), .B(n1917), .Z(n633) );
  NAND U2061 ( .A(\stack[3][6] ), .B(n2150), .Z(n1920) );
  NANDN U2062 ( .A(n2142), .B(\stack[5][6] ), .Z(n1919) );
  AND U2063 ( .A(n1920), .B(n1919), .Z(n1922) );
  NAND U2064 ( .A(n2145), .B(\stack[4][6] ), .Z(n1921) );
  NAND U2065 ( .A(n1922), .B(n1921), .Z(n634) );
  NAND U2066 ( .A(\stack[2][6] ), .B(n2150), .Z(n1924) );
  NANDN U2067 ( .A(n2142), .B(\stack[4][6] ), .Z(n1923) );
  AND U2068 ( .A(n1924), .B(n1923), .Z(n1926) );
  NAND U2069 ( .A(n2145), .B(\stack[3][6] ), .Z(n1925) );
  NAND U2070 ( .A(n1926), .B(n1925), .Z(n635) );
  NAND U2071 ( .A(n2150), .B(\stack[1][6] ), .Z(n1928) );
  NANDN U2072 ( .A(n2142), .B(\stack[3][6] ), .Z(n1927) );
  AND U2073 ( .A(n1928), .B(n1927), .Z(n1930) );
  NAND U2074 ( .A(n2145), .B(\stack[2][6] ), .Z(n1929) );
  NAND U2075 ( .A(n1930), .B(n1929), .Z(n636) );
  NAND U2076 ( .A(n2150), .B(o[6]), .Z(n1932) );
  NANDN U2077 ( .A(n2142), .B(\stack[2][6] ), .Z(n1931) );
  AND U2078 ( .A(n1932), .B(n1931), .Z(n1934) );
  NAND U2079 ( .A(\stack[1][6] ), .B(n2145), .Z(n1933) );
  NAND U2080 ( .A(n1934), .B(n1933), .Z(n637) );
  NAND U2081 ( .A(x[6]), .B(n2150), .Z(n1936) );
  NAND U2082 ( .A(\stack[1][6] ), .B(n2154), .Z(n1935) );
  NAND U2083 ( .A(n1936), .B(n1935), .Z(n1940) );
  ANDN U2084 ( .B(n1937), .A(n2151), .Z(n1938) );
  NANDN U2085 ( .A(n1940), .B(n1939), .Z(n1947) );
  OR U2086 ( .A(n2132), .B(n1941), .Z(n1943) );
  NAND U2087 ( .A(\stack[1][6] ), .B(n2152), .Z(n1942) );
  AND U2088 ( .A(n1943), .B(n1942), .Z(n1944) );
  NAND U2089 ( .A(n2148), .B(n1944), .Z(n1945) );
  NAND U2090 ( .A(o[6]), .B(n1945), .Z(n1946) );
  NANDN U2091 ( .A(n1947), .B(n1946), .Z(n638) );
  NAND U2092 ( .A(\stack[6][5] ), .B(n2150), .Z(n1949) );
  NANDN U2093 ( .A(n2150), .B(\stack[7][5] ), .Z(n1948) );
  NAND U2094 ( .A(n1949), .B(n1948), .Z(n639) );
  NAND U2095 ( .A(\stack[5][5] ), .B(n2150), .Z(n1951) );
  NANDN U2096 ( .A(n2142), .B(\stack[7][5] ), .Z(n1950) );
  AND U2097 ( .A(n1951), .B(n1950), .Z(n1953) );
  NAND U2098 ( .A(n2145), .B(\stack[6][5] ), .Z(n1952) );
  NAND U2099 ( .A(n1953), .B(n1952), .Z(n640) );
  NAND U2100 ( .A(\stack[4][5] ), .B(n2150), .Z(n1955) );
  NANDN U2101 ( .A(n2142), .B(\stack[6][5] ), .Z(n1954) );
  AND U2102 ( .A(n1955), .B(n1954), .Z(n1957) );
  NAND U2103 ( .A(n2145), .B(\stack[5][5] ), .Z(n1956) );
  NAND U2104 ( .A(n1957), .B(n1956), .Z(n641) );
  NAND U2105 ( .A(\stack[3][5] ), .B(n2150), .Z(n1959) );
  NANDN U2106 ( .A(n2142), .B(\stack[5][5] ), .Z(n1958) );
  AND U2107 ( .A(n1959), .B(n1958), .Z(n1961) );
  NAND U2108 ( .A(n2145), .B(\stack[4][5] ), .Z(n1960) );
  NAND U2109 ( .A(n1961), .B(n1960), .Z(n642) );
  NAND U2110 ( .A(\stack[2][5] ), .B(n2150), .Z(n1963) );
  NANDN U2111 ( .A(n2142), .B(\stack[4][5] ), .Z(n1962) );
  AND U2112 ( .A(n1963), .B(n1962), .Z(n1965) );
  NAND U2113 ( .A(n2145), .B(\stack[3][5] ), .Z(n1964) );
  NAND U2114 ( .A(n1965), .B(n1964), .Z(n643) );
  NAND U2115 ( .A(n2150), .B(\stack[1][5] ), .Z(n1967) );
  NANDN U2116 ( .A(n2142), .B(\stack[3][5] ), .Z(n1966) );
  AND U2117 ( .A(n1967), .B(n1966), .Z(n1969) );
  NAND U2118 ( .A(n2145), .B(\stack[2][5] ), .Z(n1968) );
  NAND U2119 ( .A(n1969), .B(n1968), .Z(n644) );
  NAND U2120 ( .A(n2150), .B(o[5]), .Z(n1971) );
  NANDN U2121 ( .A(n2142), .B(\stack[2][5] ), .Z(n1970) );
  AND U2122 ( .A(n1971), .B(n1970), .Z(n1973) );
  NAND U2123 ( .A(\stack[1][5] ), .B(n2145), .Z(n1972) );
  NAND U2124 ( .A(n1973), .B(n1972), .Z(n645) );
  NAND U2125 ( .A(o[5]), .B(n2152), .Z(n1974) );
  NANDN U2126 ( .A(n2154), .B(n1974), .Z(n1975) );
  NAND U2127 ( .A(\stack[1][5] ), .B(n1975), .Z(n1978) );
  NAND U2128 ( .A(x[5]), .B(n2150), .Z(n1976) );
  AND U2129 ( .A(n1978), .B(n1977), .Z(n1980) );
  NANDN U2130 ( .A(n2148), .B(o[5]), .Z(n1979) );
  AND U2131 ( .A(n1980), .B(n1979), .Z(n1985) );
  XNOR U2132 ( .A(n1982), .B(n1981), .Z(n1983) );
  NANDN U2133 ( .A(n2151), .B(n1983), .Z(n1984) );
  NAND U2134 ( .A(n1985), .B(n1984), .Z(n646) );
  NAND U2135 ( .A(\stack[6][4] ), .B(n2150), .Z(n1987) );
  NANDN U2136 ( .A(n2150), .B(\stack[7][4] ), .Z(n1986) );
  NAND U2137 ( .A(n1987), .B(n1986), .Z(n647) );
  NAND U2138 ( .A(\stack[5][4] ), .B(n2150), .Z(n1989) );
  NANDN U2139 ( .A(n2142), .B(\stack[7][4] ), .Z(n1988) );
  AND U2140 ( .A(n1989), .B(n1988), .Z(n1991) );
  NAND U2141 ( .A(n2145), .B(\stack[6][4] ), .Z(n1990) );
  NAND U2142 ( .A(n1991), .B(n1990), .Z(n648) );
  NAND U2143 ( .A(\stack[4][4] ), .B(n2150), .Z(n1993) );
  NANDN U2144 ( .A(n2142), .B(\stack[6][4] ), .Z(n1992) );
  AND U2145 ( .A(n1993), .B(n1992), .Z(n1995) );
  NAND U2146 ( .A(n2145), .B(\stack[5][4] ), .Z(n1994) );
  NAND U2147 ( .A(n1995), .B(n1994), .Z(n649) );
  NAND U2148 ( .A(\stack[3][4] ), .B(n2150), .Z(n1997) );
  NANDN U2149 ( .A(n2142), .B(\stack[5][4] ), .Z(n1996) );
  AND U2150 ( .A(n1997), .B(n1996), .Z(n1999) );
  NAND U2151 ( .A(n2145), .B(\stack[4][4] ), .Z(n1998) );
  NAND U2152 ( .A(n1999), .B(n1998), .Z(n650) );
  NAND U2153 ( .A(\stack[2][4] ), .B(n2150), .Z(n2001) );
  NANDN U2154 ( .A(n2142), .B(\stack[4][4] ), .Z(n2000) );
  AND U2155 ( .A(n2001), .B(n2000), .Z(n2003) );
  NAND U2156 ( .A(n2145), .B(\stack[3][4] ), .Z(n2002) );
  NAND U2157 ( .A(n2003), .B(n2002), .Z(n651) );
  NAND U2158 ( .A(n2150), .B(\stack[1][4] ), .Z(n2005) );
  NANDN U2159 ( .A(n2142), .B(\stack[3][4] ), .Z(n2004) );
  AND U2160 ( .A(n2005), .B(n2004), .Z(n2007) );
  NAND U2161 ( .A(n2145), .B(\stack[2][4] ), .Z(n2006) );
  NAND U2162 ( .A(n2007), .B(n2006), .Z(n652) );
  NAND U2163 ( .A(n2150), .B(o[4]), .Z(n2009) );
  NANDN U2164 ( .A(n2142), .B(\stack[2][4] ), .Z(n2008) );
  AND U2165 ( .A(n2009), .B(n2008), .Z(n2011) );
  NAND U2166 ( .A(\stack[1][4] ), .B(n2145), .Z(n2010) );
  NAND U2167 ( .A(n2011), .B(n2010), .Z(n653) );
  NAND U2168 ( .A(x[4]), .B(n2150), .Z(n2013) );
  NAND U2169 ( .A(\stack[1][4] ), .B(n2154), .Z(n2012) );
  NAND U2170 ( .A(n2013), .B(n2012), .Z(n2017) );
  ANDN U2171 ( .B(n2014), .A(n2151), .Z(n2015) );
  NANDN U2172 ( .A(n2017), .B(n2016), .Z(n2024) );
  OR U2173 ( .A(n2132), .B(n2018), .Z(n2020) );
  NAND U2174 ( .A(\stack[1][4] ), .B(n2152), .Z(n2019) );
  AND U2175 ( .A(n2020), .B(n2019), .Z(n2021) );
  NAND U2176 ( .A(n2148), .B(n2021), .Z(n2022) );
  NAND U2177 ( .A(o[4]), .B(n2022), .Z(n2023) );
  NANDN U2178 ( .A(n2024), .B(n2023), .Z(n654) );
  NAND U2179 ( .A(\stack[6][3] ), .B(n2150), .Z(n2026) );
  NANDN U2180 ( .A(n2150), .B(\stack[7][3] ), .Z(n2025) );
  NAND U2181 ( .A(n2026), .B(n2025), .Z(n655) );
  NAND U2182 ( .A(\stack[5][3] ), .B(n2150), .Z(n2028) );
  NANDN U2183 ( .A(n2142), .B(\stack[7][3] ), .Z(n2027) );
  AND U2184 ( .A(n2028), .B(n2027), .Z(n2030) );
  NAND U2185 ( .A(n2145), .B(\stack[6][3] ), .Z(n2029) );
  NAND U2186 ( .A(n2030), .B(n2029), .Z(n656) );
  NAND U2187 ( .A(\stack[4][3] ), .B(n2150), .Z(n2032) );
  NANDN U2188 ( .A(n2142), .B(\stack[6][3] ), .Z(n2031) );
  AND U2189 ( .A(n2032), .B(n2031), .Z(n2034) );
  NAND U2190 ( .A(n2145), .B(\stack[5][3] ), .Z(n2033) );
  NAND U2191 ( .A(n2034), .B(n2033), .Z(n657) );
  NAND U2192 ( .A(\stack[3][3] ), .B(n2150), .Z(n2036) );
  NANDN U2193 ( .A(n2142), .B(\stack[5][3] ), .Z(n2035) );
  AND U2194 ( .A(n2036), .B(n2035), .Z(n2038) );
  NAND U2195 ( .A(n2145), .B(\stack[4][3] ), .Z(n2037) );
  NAND U2196 ( .A(n2038), .B(n2037), .Z(n658) );
  NAND U2197 ( .A(\stack[2][3] ), .B(n2150), .Z(n2040) );
  NANDN U2198 ( .A(n2142), .B(\stack[4][3] ), .Z(n2039) );
  AND U2199 ( .A(n2040), .B(n2039), .Z(n2042) );
  NAND U2200 ( .A(n2145), .B(\stack[3][3] ), .Z(n2041) );
  NAND U2201 ( .A(n2042), .B(n2041), .Z(n659) );
  NAND U2202 ( .A(n2150), .B(\stack[1][3] ), .Z(n2044) );
  NANDN U2203 ( .A(n2142), .B(\stack[3][3] ), .Z(n2043) );
  AND U2204 ( .A(n2044), .B(n2043), .Z(n2046) );
  NAND U2205 ( .A(n2145), .B(\stack[2][3] ), .Z(n2045) );
  NAND U2206 ( .A(n2046), .B(n2045), .Z(n660) );
  NAND U2207 ( .A(n2150), .B(o[3]), .Z(n2048) );
  NANDN U2208 ( .A(n2142), .B(\stack[2][3] ), .Z(n2047) );
  AND U2209 ( .A(n2048), .B(n2047), .Z(n2050) );
  NAND U2210 ( .A(\stack[1][3] ), .B(n2145), .Z(n2049) );
  NAND U2211 ( .A(n2050), .B(n2049), .Z(n661) );
  NAND U2212 ( .A(o[3]), .B(n2152), .Z(n2051) );
  NANDN U2213 ( .A(n2154), .B(n2051), .Z(n2052) );
  NAND U2214 ( .A(\stack[1][3] ), .B(n2052), .Z(n2055) );
  NAND U2215 ( .A(x[3]), .B(n2150), .Z(n2053) );
  AND U2216 ( .A(n2055), .B(n2054), .Z(n2057) );
  NANDN U2217 ( .A(n2148), .B(o[3]), .Z(n2056) );
  AND U2218 ( .A(n2057), .B(n2056), .Z(n2062) );
  XNOR U2219 ( .A(n2059), .B(n2058), .Z(n2060) );
  NANDN U2220 ( .A(n2151), .B(n2060), .Z(n2061) );
  NAND U2221 ( .A(n2062), .B(n2061), .Z(n662) );
  NAND U2222 ( .A(\stack[6][2] ), .B(n2150), .Z(n2064) );
  NANDN U2223 ( .A(n2150), .B(\stack[7][2] ), .Z(n2063) );
  NAND U2224 ( .A(n2064), .B(n2063), .Z(n663) );
  NAND U2225 ( .A(\stack[5][2] ), .B(n2150), .Z(n2066) );
  NANDN U2226 ( .A(n2142), .B(\stack[7][2] ), .Z(n2065) );
  AND U2227 ( .A(n2066), .B(n2065), .Z(n2068) );
  NAND U2228 ( .A(n2145), .B(\stack[6][2] ), .Z(n2067) );
  NAND U2229 ( .A(n2068), .B(n2067), .Z(n664) );
  NAND U2230 ( .A(\stack[4][2] ), .B(n2150), .Z(n2070) );
  NANDN U2231 ( .A(n2142), .B(\stack[6][2] ), .Z(n2069) );
  AND U2232 ( .A(n2070), .B(n2069), .Z(n2072) );
  NAND U2233 ( .A(n2145), .B(\stack[5][2] ), .Z(n2071) );
  NAND U2234 ( .A(n2072), .B(n2071), .Z(n665) );
  NAND U2235 ( .A(\stack[3][2] ), .B(n2150), .Z(n2074) );
  NANDN U2236 ( .A(n2142), .B(\stack[5][2] ), .Z(n2073) );
  AND U2237 ( .A(n2074), .B(n2073), .Z(n2076) );
  NAND U2238 ( .A(n2145), .B(\stack[4][2] ), .Z(n2075) );
  NAND U2239 ( .A(n2076), .B(n2075), .Z(n666) );
  NAND U2240 ( .A(\stack[2][2] ), .B(n2150), .Z(n2078) );
  NANDN U2241 ( .A(n2142), .B(\stack[4][2] ), .Z(n2077) );
  AND U2242 ( .A(n2078), .B(n2077), .Z(n2080) );
  NAND U2243 ( .A(n2145), .B(\stack[3][2] ), .Z(n2079) );
  NAND U2244 ( .A(n2080), .B(n2079), .Z(n667) );
  NAND U2245 ( .A(n2150), .B(\stack[1][2] ), .Z(n2082) );
  NANDN U2246 ( .A(n2142), .B(\stack[3][2] ), .Z(n2081) );
  AND U2247 ( .A(n2082), .B(n2081), .Z(n2084) );
  NAND U2248 ( .A(n2145), .B(\stack[2][2] ), .Z(n2083) );
  NAND U2249 ( .A(n2084), .B(n2083), .Z(n668) );
  NAND U2250 ( .A(n2150), .B(o[2]), .Z(n2086) );
  NANDN U2251 ( .A(n2142), .B(\stack[2][2] ), .Z(n2085) );
  AND U2252 ( .A(n2086), .B(n2085), .Z(n2088) );
  NAND U2253 ( .A(\stack[1][2] ), .B(n2145), .Z(n2087) );
  NAND U2254 ( .A(n2088), .B(n2087), .Z(n669) );
  NAND U2255 ( .A(o[2]), .B(n2152), .Z(n2089) );
  NANDN U2256 ( .A(n2154), .B(n2089), .Z(n2090) );
  NAND U2257 ( .A(\stack[1][2] ), .B(n2090), .Z(n2093) );
  NAND U2258 ( .A(x[2]), .B(n2150), .Z(n2091) );
  AND U2259 ( .A(n2093), .B(n2092), .Z(n2095) );
  NANDN U2260 ( .A(n2148), .B(o[2]), .Z(n2094) );
  AND U2261 ( .A(n2095), .B(n2094), .Z(n2100) );
  XNOR U2262 ( .A(n2097), .B(n2096), .Z(n2098) );
  NANDN U2263 ( .A(n2151), .B(n2098), .Z(n2099) );
  NAND U2264 ( .A(n2100), .B(n2099), .Z(n670) );
  NAND U2265 ( .A(\stack[6][1] ), .B(n2150), .Z(n2102) );
  NANDN U2266 ( .A(n2150), .B(\stack[7][1] ), .Z(n2101) );
  NAND U2267 ( .A(n2102), .B(n2101), .Z(n671) );
  NAND U2268 ( .A(\stack[5][1] ), .B(n2150), .Z(n2104) );
  NANDN U2269 ( .A(n2142), .B(\stack[7][1] ), .Z(n2103) );
  AND U2270 ( .A(n2104), .B(n2103), .Z(n2106) );
  NAND U2271 ( .A(n2145), .B(\stack[6][1] ), .Z(n2105) );
  NAND U2272 ( .A(n2106), .B(n2105), .Z(n672) );
  NAND U2273 ( .A(\stack[4][1] ), .B(n2150), .Z(n2108) );
  NANDN U2274 ( .A(n2142), .B(\stack[6][1] ), .Z(n2107) );
  AND U2275 ( .A(n2108), .B(n2107), .Z(n2110) );
  NAND U2276 ( .A(n2145), .B(\stack[5][1] ), .Z(n2109) );
  NAND U2277 ( .A(n2110), .B(n2109), .Z(n673) );
  NAND U2278 ( .A(\stack[3][1] ), .B(n2150), .Z(n2112) );
  NANDN U2279 ( .A(n2142), .B(\stack[5][1] ), .Z(n2111) );
  AND U2280 ( .A(n2112), .B(n2111), .Z(n2114) );
  NAND U2281 ( .A(n2145), .B(\stack[4][1] ), .Z(n2113) );
  NAND U2282 ( .A(n2114), .B(n2113), .Z(n674) );
  NAND U2283 ( .A(\stack[2][1] ), .B(n2150), .Z(n2116) );
  NANDN U2284 ( .A(n2142), .B(\stack[4][1] ), .Z(n2115) );
  AND U2285 ( .A(n2116), .B(n2115), .Z(n2118) );
  NAND U2286 ( .A(n2145), .B(\stack[3][1] ), .Z(n2117) );
  NAND U2287 ( .A(n2118), .B(n2117), .Z(n675) );
  NAND U2288 ( .A(n2150), .B(\stack[1][1] ), .Z(n2120) );
  NANDN U2289 ( .A(n2142), .B(\stack[3][1] ), .Z(n2119) );
  AND U2290 ( .A(n2120), .B(n2119), .Z(n2122) );
  NAND U2291 ( .A(n2145), .B(\stack[2][1] ), .Z(n2121) );
  NAND U2292 ( .A(n2122), .B(n2121), .Z(n676) );
  NAND U2293 ( .A(n2150), .B(o[1]), .Z(n2124) );
  NANDN U2294 ( .A(n2142), .B(\stack[2][1] ), .Z(n2123) );
  AND U2295 ( .A(n2124), .B(n2123), .Z(n2126) );
  NAND U2296 ( .A(\stack[1][1] ), .B(n2145), .Z(n2125) );
  NAND U2297 ( .A(n2126), .B(n2125), .Z(n677) );
  NAND U2298 ( .A(n2150), .B(x[1]), .Z(n2130) );
  NOR U2299 ( .A(n2151), .B(n2127), .Z(n2128) );
  NAND U2300 ( .A(n2131), .B(n2128), .Z(n2129) );
  AND U2301 ( .A(n2130), .B(n2129), .Z(n2138) );
  OR U2302 ( .A(n2132), .B(n2131), .Z(n2134) );
  NAND U2303 ( .A(\stack[1][1] ), .B(n2152), .Z(n2133) );
  AND U2304 ( .A(n2134), .B(n2133), .Z(n2135) );
  NAND U2305 ( .A(n2135), .B(n2148), .Z(n2136) );
  NAND U2306 ( .A(o[1]), .B(n2136), .Z(n2137) );
  AND U2307 ( .A(n2138), .B(n2137), .Z(n2141) );
  NAND U2308 ( .A(n2154), .B(\stack[1][1] ), .Z(n2139) );
  NAND U2309 ( .A(n2141), .B(n2140), .Z(n678) );
  NAND U2310 ( .A(n2150), .B(o[0]), .Z(n2144) );
  NANDN U2311 ( .A(n2142), .B(\stack[2][0] ), .Z(n2143) );
  AND U2312 ( .A(n2144), .B(n2143), .Z(n2147) );
  NAND U2313 ( .A(\stack[1][0] ), .B(n2145), .Z(n2146) );
  NAND U2314 ( .A(n2147), .B(n2146), .Z(n679) );
  NANDN U2315 ( .A(n2148), .B(o[0]), .Z(n2149) );
  NAND U2316 ( .A(x[0]), .B(n2150), .Z(n2158) );
  NANDN U2317 ( .A(n2152), .B(n2151), .Z(n2153) );
  NAND U2318 ( .A(o[0]), .B(n2153), .Z(n2155) );
  ANDN U2319 ( .B(n2155), .A(n2154), .Z(n2156) );
  NANDN U2320 ( .A(n2156), .B(\stack[1][0] ), .Z(n2157) );
  AND U2321 ( .A(n2158), .B(n2157), .Z(n2159) );
  NANDN U2322 ( .A(n2160), .B(n2159), .Z(n680) );
endmodule

