
module mult_N128_CC64 ( clk, rst, a, b, c );
  input [127:0] a;
  input [1:0] b;
  output [255:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654;
  wire   [255:0] sreg;

  DFF \sreg_reg[253]  ( .D(c[255]), .CLK(clk), .RST(rst), .Q(sreg[253]) );
  DFF \sreg_reg[252]  ( .D(c[254]), .CLK(clk), .RST(rst), .Q(sreg[252]) );
  DFF \sreg_reg[251]  ( .D(c[253]), .CLK(clk), .RST(rst), .Q(sreg[251]) );
  DFF \sreg_reg[250]  ( .D(c[252]), .CLK(clk), .RST(rst), .Q(sreg[250]) );
  DFF \sreg_reg[249]  ( .D(c[251]), .CLK(clk), .RST(rst), .Q(sreg[249]) );
  DFF \sreg_reg[248]  ( .D(c[250]), .CLK(clk), .RST(rst), .Q(sreg[248]) );
  DFF \sreg_reg[247]  ( .D(c[249]), .CLK(clk), .RST(rst), .Q(sreg[247]) );
  DFF \sreg_reg[246]  ( .D(c[248]), .CLK(clk), .RST(rst), .Q(sreg[246]) );
  DFF \sreg_reg[245]  ( .D(c[247]), .CLK(clk), .RST(rst), .Q(sreg[245]) );
  DFF \sreg_reg[244]  ( .D(c[246]), .CLK(clk), .RST(rst), .Q(sreg[244]) );
  DFF \sreg_reg[243]  ( .D(c[245]), .CLK(clk), .RST(rst), .Q(sreg[243]) );
  DFF \sreg_reg[242]  ( .D(c[244]), .CLK(clk), .RST(rst), .Q(sreg[242]) );
  DFF \sreg_reg[241]  ( .D(c[243]), .CLK(clk), .RST(rst), .Q(sreg[241]) );
  DFF \sreg_reg[240]  ( .D(c[242]), .CLK(clk), .RST(rst), .Q(sreg[240]) );
  DFF \sreg_reg[239]  ( .D(c[241]), .CLK(clk), .RST(rst), .Q(sreg[239]) );
  DFF \sreg_reg[238]  ( .D(c[240]), .CLK(clk), .RST(rst), .Q(sreg[238]) );
  DFF \sreg_reg[237]  ( .D(c[239]), .CLK(clk), .RST(rst), .Q(sreg[237]) );
  DFF \sreg_reg[236]  ( .D(c[238]), .CLK(clk), .RST(rst), .Q(sreg[236]) );
  DFF \sreg_reg[235]  ( .D(c[237]), .CLK(clk), .RST(rst), .Q(sreg[235]) );
  DFF \sreg_reg[234]  ( .D(c[236]), .CLK(clk), .RST(rst), .Q(sreg[234]) );
  DFF \sreg_reg[233]  ( .D(c[235]), .CLK(clk), .RST(rst), .Q(sreg[233]) );
  DFF \sreg_reg[232]  ( .D(c[234]), .CLK(clk), .RST(rst), .Q(sreg[232]) );
  DFF \sreg_reg[231]  ( .D(c[233]), .CLK(clk), .RST(rst), .Q(sreg[231]) );
  DFF \sreg_reg[230]  ( .D(c[232]), .CLK(clk), .RST(rst), .Q(sreg[230]) );
  DFF \sreg_reg[229]  ( .D(c[231]), .CLK(clk), .RST(rst), .Q(sreg[229]) );
  DFF \sreg_reg[228]  ( .D(c[230]), .CLK(clk), .RST(rst), .Q(sreg[228]) );
  DFF \sreg_reg[227]  ( .D(c[229]), .CLK(clk), .RST(rst), .Q(sreg[227]) );
  DFF \sreg_reg[226]  ( .D(c[228]), .CLK(clk), .RST(rst), .Q(sreg[226]) );
  DFF \sreg_reg[225]  ( .D(c[227]), .CLK(clk), .RST(rst), .Q(sreg[225]) );
  DFF \sreg_reg[224]  ( .D(c[226]), .CLK(clk), .RST(rst), .Q(sreg[224]) );
  DFF \sreg_reg[223]  ( .D(c[225]), .CLK(clk), .RST(rst), .Q(sreg[223]) );
  DFF \sreg_reg[222]  ( .D(c[224]), .CLK(clk), .RST(rst), .Q(sreg[222]) );
  DFF \sreg_reg[221]  ( .D(c[223]), .CLK(clk), .RST(rst), .Q(sreg[221]) );
  DFF \sreg_reg[220]  ( .D(c[222]), .CLK(clk), .RST(rst), .Q(sreg[220]) );
  DFF \sreg_reg[219]  ( .D(c[221]), .CLK(clk), .RST(rst), .Q(sreg[219]) );
  DFF \sreg_reg[218]  ( .D(c[220]), .CLK(clk), .RST(rst), .Q(sreg[218]) );
  DFF \sreg_reg[217]  ( .D(c[219]), .CLK(clk), .RST(rst), .Q(sreg[217]) );
  DFF \sreg_reg[216]  ( .D(c[218]), .CLK(clk), .RST(rst), .Q(sreg[216]) );
  DFF \sreg_reg[215]  ( .D(c[217]), .CLK(clk), .RST(rst), .Q(sreg[215]) );
  DFF \sreg_reg[214]  ( .D(c[216]), .CLK(clk), .RST(rst), .Q(sreg[214]) );
  DFF \sreg_reg[213]  ( .D(c[215]), .CLK(clk), .RST(rst), .Q(sreg[213]) );
  DFF \sreg_reg[212]  ( .D(c[214]), .CLK(clk), .RST(rst), .Q(sreg[212]) );
  DFF \sreg_reg[211]  ( .D(c[213]), .CLK(clk), .RST(rst), .Q(sreg[211]) );
  DFF \sreg_reg[210]  ( .D(c[212]), .CLK(clk), .RST(rst), .Q(sreg[210]) );
  DFF \sreg_reg[209]  ( .D(c[211]), .CLK(clk), .RST(rst), .Q(sreg[209]) );
  DFF \sreg_reg[208]  ( .D(c[210]), .CLK(clk), .RST(rst), .Q(sreg[208]) );
  DFF \sreg_reg[207]  ( .D(c[209]), .CLK(clk), .RST(rst), .Q(sreg[207]) );
  DFF \sreg_reg[206]  ( .D(c[208]), .CLK(clk), .RST(rst), .Q(sreg[206]) );
  DFF \sreg_reg[205]  ( .D(c[207]), .CLK(clk), .RST(rst), .Q(sreg[205]) );
  DFF \sreg_reg[204]  ( .D(c[206]), .CLK(clk), .RST(rst), .Q(sreg[204]) );
  DFF \sreg_reg[203]  ( .D(c[205]), .CLK(clk), .RST(rst), .Q(sreg[203]) );
  DFF \sreg_reg[202]  ( .D(c[204]), .CLK(clk), .RST(rst), .Q(sreg[202]) );
  DFF \sreg_reg[201]  ( .D(c[203]), .CLK(clk), .RST(rst), .Q(sreg[201]) );
  DFF \sreg_reg[200]  ( .D(c[202]), .CLK(clk), .RST(rst), .Q(sreg[200]) );
  DFF \sreg_reg[199]  ( .D(c[201]), .CLK(clk), .RST(rst), .Q(sreg[199]) );
  DFF \sreg_reg[198]  ( .D(c[200]), .CLK(clk), .RST(rst), .Q(sreg[198]) );
  DFF \sreg_reg[197]  ( .D(c[199]), .CLK(clk), .RST(rst), .Q(sreg[197]) );
  DFF \sreg_reg[196]  ( .D(c[198]), .CLK(clk), .RST(rst), .Q(sreg[196]) );
  DFF \sreg_reg[195]  ( .D(c[197]), .CLK(clk), .RST(rst), .Q(sreg[195]) );
  DFF \sreg_reg[194]  ( .D(c[196]), .CLK(clk), .RST(rst), .Q(sreg[194]) );
  DFF \sreg_reg[193]  ( .D(c[195]), .CLK(clk), .RST(rst), .Q(sreg[193]) );
  DFF \sreg_reg[192]  ( .D(c[194]), .CLK(clk), .RST(rst), .Q(sreg[192]) );
  DFF \sreg_reg[191]  ( .D(c[193]), .CLK(clk), .RST(rst), .Q(sreg[191]) );
  DFF \sreg_reg[190]  ( .D(c[192]), .CLK(clk), .RST(rst), .Q(sreg[190]) );
  DFF \sreg_reg[189]  ( .D(c[191]), .CLK(clk), .RST(rst), .Q(sreg[189]) );
  DFF \sreg_reg[188]  ( .D(c[190]), .CLK(clk), .RST(rst), .Q(sreg[188]) );
  DFF \sreg_reg[187]  ( .D(c[189]), .CLK(clk), .RST(rst), .Q(sreg[187]) );
  DFF \sreg_reg[186]  ( .D(c[188]), .CLK(clk), .RST(rst), .Q(sreg[186]) );
  DFF \sreg_reg[185]  ( .D(c[187]), .CLK(clk), .RST(rst), .Q(sreg[185]) );
  DFF \sreg_reg[184]  ( .D(c[186]), .CLK(clk), .RST(rst), .Q(sreg[184]) );
  DFF \sreg_reg[183]  ( .D(c[185]), .CLK(clk), .RST(rst), .Q(sreg[183]) );
  DFF \sreg_reg[182]  ( .D(c[184]), .CLK(clk), .RST(rst), .Q(sreg[182]) );
  DFF \sreg_reg[181]  ( .D(c[183]), .CLK(clk), .RST(rst), .Q(sreg[181]) );
  DFF \sreg_reg[180]  ( .D(c[182]), .CLK(clk), .RST(rst), .Q(sreg[180]) );
  DFF \sreg_reg[179]  ( .D(c[181]), .CLK(clk), .RST(rst), .Q(sreg[179]) );
  DFF \sreg_reg[178]  ( .D(c[180]), .CLK(clk), .RST(rst), .Q(sreg[178]) );
  DFF \sreg_reg[177]  ( .D(c[179]), .CLK(clk), .RST(rst), .Q(sreg[177]) );
  DFF \sreg_reg[176]  ( .D(c[178]), .CLK(clk), .RST(rst), .Q(sreg[176]) );
  DFF \sreg_reg[175]  ( .D(c[177]), .CLK(clk), .RST(rst), .Q(sreg[175]) );
  DFF \sreg_reg[174]  ( .D(c[176]), .CLK(clk), .RST(rst), .Q(sreg[174]) );
  DFF \sreg_reg[173]  ( .D(c[175]), .CLK(clk), .RST(rst), .Q(sreg[173]) );
  DFF \sreg_reg[172]  ( .D(c[174]), .CLK(clk), .RST(rst), .Q(sreg[172]) );
  DFF \sreg_reg[171]  ( .D(c[173]), .CLK(clk), .RST(rst), .Q(sreg[171]) );
  DFF \sreg_reg[170]  ( .D(c[172]), .CLK(clk), .RST(rst), .Q(sreg[170]) );
  DFF \sreg_reg[169]  ( .D(c[171]), .CLK(clk), .RST(rst), .Q(sreg[169]) );
  DFF \sreg_reg[168]  ( .D(c[170]), .CLK(clk), .RST(rst), .Q(sreg[168]) );
  DFF \sreg_reg[167]  ( .D(c[169]), .CLK(clk), .RST(rst), .Q(sreg[167]) );
  DFF \sreg_reg[166]  ( .D(c[168]), .CLK(clk), .RST(rst), .Q(sreg[166]) );
  DFF \sreg_reg[165]  ( .D(c[167]), .CLK(clk), .RST(rst), .Q(sreg[165]) );
  DFF \sreg_reg[164]  ( .D(c[166]), .CLK(clk), .RST(rst), .Q(sreg[164]) );
  DFF \sreg_reg[163]  ( .D(c[165]), .CLK(clk), .RST(rst), .Q(sreg[163]) );
  DFF \sreg_reg[162]  ( .D(c[164]), .CLK(clk), .RST(rst), .Q(sreg[162]) );
  DFF \sreg_reg[161]  ( .D(c[163]), .CLK(clk), .RST(rst), .Q(sreg[161]) );
  DFF \sreg_reg[160]  ( .D(c[162]), .CLK(clk), .RST(rst), .Q(sreg[160]) );
  DFF \sreg_reg[159]  ( .D(c[161]), .CLK(clk), .RST(rst), .Q(sreg[159]) );
  DFF \sreg_reg[158]  ( .D(c[160]), .CLK(clk), .RST(rst), .Q(sreg[158]) );
  DFF \sreg_reg[157]  ( .D(c[159]), .CLK(clk), .RST(rst), .Q(sreg[157]) );
  DFF \sreg_reg[156]  ( .D(c[158]), .CLK(clk), .RST(rst), .Q(sreg[156]) );
  DFF \sreg_reg[155]  ( .D(c[157]), .CLK(clk), .RST(rst), .Q(sreg[155]) );
  DFF \sreg_reg[154]  ( .D(c[156]), .CLK(clk), .RST(rst), .Q(sreg[154]) );
  DFF \sreg_reg[153]  ( .D(c[155]), .CLK(clk), .RST(rst), .Q(sreg[153]) );
  DFF \sreg_reg[152]  ( .D(c[154]), .CLK(clk), .RST(rst), .Q(sreg[152]) );
  DFF \sreg_reg[151]  ( .D(c[153]), .CLK(clk), .RST(rst), .Q(sreg[151]) );
  DFF \sreg_reg[150]  ( .D(c[152]), .CLK(clk), .RST(rst), .Q(sreg[150]) );
  DFF \sreg_reg[149]  ( .D(c[151]), .CLK(clk), .RST(rst), .Q(sreg[149]) );
  DFF \sreg_reg[148]  ( .D(c[150]), .CLK(clk), .RST(rst), .Q(sreg[148]) );
  DFF \sreg_reg[147]  ( .D(c[149]), .CLK(clk), .RST(rst), .Q(sreg[147]) );
  DFF \sreg_reg[146]  ( .D(c[148]), .CLK(clk), .RST(rst), .Q(sreg[146]) );
  DFF \sreg_reg[145]  ( .D(c[147]), .CLK(clk), .RST(rst), .Q(sreg[145]) );
  DFF \sreg_reg[144]  ( .D(c[146]), .CLK(clk), .RST(rst), .Q(sreg[144]) );
  DFF \sreg_reg[143]  ( .D(c[145]), .CLK(clk), .RST(rst), .Q(sreg[143]) );
  DFF \sreg_reg[142]  ( .D(c[144]), .CLK(clk), .RST(rst), .Q(sreg[142]) );
  DFF \sreg_reg[141]  ( .D(c[143]), .CLK(clk), .RST(rst), .Q(sreg[141]) );
  DFF \sreg_reg[140]  ( .D(c[142]), .CLK(clk), .RST(rst), .Q(sreg[140]) );
  DFF \sreg_reg[139]  ( .D(c[141]), .CLK(clk), .RST(rst), .Q(sreg[139]) );
  DFF \sreg_reg[138]  ( .D(c[140]), .CLK(clk), .RST(rst), .Q(sreg[138]) );
  DFF \sreg_reg[137]  ( .D(c[139]), .CLK(clk), .RST(rst), .Q(sreg[137]) );
  DFF \sreg_reg[136]  ( .D(c[138]), .CLK(clk), .RST(rst), .Q(sreg[136]) );
  DFF \sreg_reg[135]  ( .D(c[137]), .CLK(clk), .RST(rst), .Q(sreg[135]) );
  DFF \sreg_reg[134]  ( .D(c[136]), .CLK(clk), .RST(rst), .Q(sreg[134]) );
  DFF \sreg_reg[133]  ( .D(c[135]), .CLK(clk), .RST(rst), .Q(sreg[133]) );
  DFF \sreg_reg[132]  ( .D(c[134]), .CLK(clk), .RST(rst), .Q(sreg[132]) );
  DFF \sreg_reg[131]  ( .D(c[133]), .CLK(clk), .RST(rst), .Q(sreg[131]) );
  DFF \sreg_reg[130]  ( .D(c[132]), .CLK(clk), .RST(rst), .Q(sreg[130]) );
  DFF \sreg_reg[129]  ( .D(c[131]), .CLK(clk), .RST(rst), .Q(sreg[129]) );
  DFF \sreg_reg[128]  ( .D(c[130]), .CLK(clk), .RST(rst), .Q(sreg[128]) );
  DFF \sreg_reg[127]  ( .D(c[129]), .CLK(clk), .RST(rst), .Q(sreg[127]) );
  DFF \sreg_reg[126]  ( .D(c[128]), .CLK(clk), .RST(rst), .Q(sreg[126]) );
  DFF \sreg_reg[125]  ( .D(c[127]), .CLK(clk), .RST(rst), .Q(c[125]) );
  DFF \sreg_reg[124]  ( .D(c[126]), .CLK(clk), .RST(rst), .Q(c[124]) );
  DFF \sreg_reg[123]  ( .D(c[125]), .CLK(clk), .RST(rst), .Q(c[123]) );
  DFF \sreg_reg[122]  ( .D(c[124]), .CLK(clk), .RST(rst), .Q(c[122]) );
  DFF \sreg_reg[121]  ( .D(c[123]), .CLK(clk), .RST(rst), .Q(c[121]) );
  DFF \sreg_reg[120]  ( .D(c[122]), .CLK(clk), .RST(rst), .Q(c[120]) );
  DFF \sreg_reg[119]  ( .D(c[121]), .CLK(clk), .RST(rst), .Q(c[119]) );
  DFF \sreg_reg[118]  ( .D(c[120]), .CLK(clk), .RST(rst), .Q(c[118]) );
  DFF \sreg_reg[117]  ( .D(c[119]), .CLK(clk), .RST(rst), .Q(c[117]) );
  DFF \sreg_reg[116]  ( .D(c[118]), .CLK(clk), .RST(rst), .Q(c[116]) );
  DFF \sreg_reg[115]  ( .D(c[117]), .CLK(clk), .RST(rst), .Q(c[115]) );
  DFF \sreg_reg[114]  ( .D(c[116]), .CLK(clk), .RST(rst), .Q(c[114]) );
  DFF \sreg_reg[113]  ( .D(c[115]), .CLK(clk), .RST(rst), .Q(c[113]) );
  DFF \sreg_reg[112]  ( .D(c[114]), .CLK(clk), .RST(rst), .Q(c[112]) );
  DFF \sreg_reg[111]  ( .D(c[113]), .CLK(clk), .RST(rst), .Q(c[111]) );
  DFF \sreg_reg[110]  ( .D(c[112]), .CLK(clk), .RST(rst), .Q(c[110]) );
  DFF \sreg_reg[109]  ( .D(c[111]), .CLK(clk), .RST(rst), .Q(c[109]) );
  DFF \sreg_reg[108]  ( .D(c[110]), .CLK(clk), .RST(rst), .Q(c[108]) );
  DFF \sreg_reg[107]  ( .D(c[109]), .CLK(clk), .RST(rst), .Q(c[107]) );
  DFF \sreg_reg[106]  ( .D(c[108]), .CLK(clk), .RST(rst), .Q(c[106]) );
  DFF \sreg_reg[105]  ( .D(c[107]), .CLK(clk), .RST(rst), .Q(c[105]) );
  DFF \sreg_reg[104]  ( .D(c[106]), .CLK(clk), .RST(rst), .Q(c[104]) );
  DFF \sreg_reg[103]  ( .D(c[105]), .CLK(clk), .RST(rst), .Q(c[103]) );
  DFF \sreg_reg[102]  ( .D(c[104]), .CLK(clk), .RST(rst), .Q(c[102]) );
  DFF \sreg_reg[101]  ( .D(c[103]), .CLK(clk), .RST(rst), .Q(c[101]) );
  DFF \sreg_reg[100]  ( .D(c[102]), .CLK(clk), .RST(rst), .Q(c[100]) );
  DFF \sreg_reg[99]  ( .D(c[101]), .CLK(clk), .RST(rst), .Q(c[99]) );
  DFF \sreg_reg[98]  ( .D(c[100]), .CLK(clk), .RST(rst), .Q(c[98]) );
  DFF \sreg_reg[97]  ( .D(c[99]), .CLK(clk), .RST(rst), .Q(c[97]) );
  DFF \sreg_reg[96]  ( .D(c[98]), .CLK(clk), .RST(rst), .Q(c[96]) );
  DFF \sreg_reg[95]  ( .D(c[97]), .CLK(clk), .RST(rst), .Q(c[95]) );
  DFF \sreg_reg[94]  ( .D(c[96]), .CLK(clk), .RST(rst), .Q(c[94]) );
  DFF \sreg_reg[93]  ( .D(c[95]), .CLK(clk), .RST(rst), .Q(c[93]) );
  DFF \sreg_reg[92]  ( .D(c[94]), .CLK(clk), .RST(rst), .Q(c[92]) );
  DFF \sreg_reg[91]  ( .D(c[93]), .CLK(clk), .RST(rst), .Q(c[91]) );
  DFF \sreg_reg[90]  ( .D(c[92]), .CLK(clk), .RST(rst), .Q(c[90]) );
  DFF \sreg_reg[89]  ( .D(c[91]), .CLK(clk), .RST(rst), .Q(c[89]) );
  DFF \sreg_reg[88]  ( .D(c[90]), .CLK(clk), .RST(rst), .Q(c[88]) );
  DFF \sreg_reg[87]  ( .D(c[89]), .CLK(clk), .RST(rst), .Q(c[87]) );
  DFF \sreg_reg[86]  ( .D(c[88]), .CLK(clk), .RST(rst), .Q(c[86]) );
  DFF \sreg_reg[85]  ( .D(c[87]), .CLK(clk), .RST(rst), .Q(c[85]) );
  DFF \sreg_reg[84]  ( .D(c[86]), .CLK(clk), .RST(rst), .Q(c[84]) );
  DFF \sreg_reg[83]  ( .D(c[85]), .CLK(clk), .RST(rst), .Q(c[83]) );
  DFF \sreg_reg[82]  ( .D(c[84]), .CLK(clk), .RST(rst), .Q(c[82]) );
  DFF \sreg_reg[81]  ( .D(c[83]), .CLK(clk), .RST(rst), .Q(c[81]) );
  DFF \sreg_reg[80]  ( .D(c[82]), .CLK(clk), .RST(rst), .Q(c[80]) );
  DFF \sreg_reg[79]  ( .D(c[81]), .CLK(clk), .RST(rst), .Q(c[79]) );
  DFF \sreg_reg[78]  ( .D(c[80]), .CLK(clk), .RST(rst), .Q(c[78]) );
  DFF \sreg_reg[77]  ( .D(c[79]), .CLK(clk), .RST(rst), .Q(c[77]) );
  DFF \sreg_reg[76]  ( .D(c[78]), .CLK(clk), .RST(rst), .Q(c[76]) );
  DFF \sreg_reg[75]  ( .D(c[77]), .CLK(clk), .RST(rst), .Q(c[75]) );
  DFF \sreg_reg[74]  ( .D(c[76]), .CLK(clk), .RST(rst), .Q(c[74]) );
  DFF \sreg_reg[73]  ( .D(c[75]), .CLK(clk), .RST(rst), .Q(c[73]) );
  DFF \sreg_reg[72]  ( .D(c[74]), .CLK(clk), .RST(rst), .Q(c[72]) );
  DFF \sreg_reg[71]  ( .D(c[73]), .CLK(clk), .RST(rst), .Q(c[71]) );
  DFF \sreg_reg[70]  ( .D(c[72]), .CLK(clk), .RST(rst), .Q(c[70]) );
  DFF \sreg_reg[69]  ( .D(c[71]), .CLK(clk), .RST(rst), .Q(c[69]) );
  DFF \sreg_reg[68]  ( .D(c[70]), .CLK(clk), .RST(rst), .Q(c[68]) );
  DFF \sreg_reg[67]  ( .D(c[69]), .CLK(clk), .RST(rst), .Q(c[67]) );
  DFF \sreg_reg[66]  ( .D(c[68]), .CLK(clk), .RST(rst), .Q(c[66]) );
  DFF \sreg_reg[65]  ( .D(c[67]), .CLK(clk), .RST(rst), .Q(c[65]) );
  DFF \sreg_reg[64]  ( .D(c[66]), .CLK(clk), .RST(rst), .Q(c[64]) );
  DFF \sreg_reg[63]  ( .D(c[65]), .CLK(clk), .RST(rst), .Q(c[63]) );
  DFF \sreg_reg[62]  ( .D(c[64]), .CLK(clk), .RST(rst), .Q(c[62]) );
  DFF \sreg_reg[61]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[61]) );
  DFF \sreg_reg[60]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[60]) );
  DFF \sreg_reg[59]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[59]) );
  DFF \sreg_reg[58]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[58]) );
  DFF \sreg_reg[57]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[57]) );
  DFF \sreg_reg[56]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[56]) );
  DFF \sreg_reg[55]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[55]) );
  DFF \sreg_reg[54]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[54]) );
  DFF \sreg_reg[53]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[53]) );
  DFF \sreg_reg[52]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[52]) );
  DFF \sreg_reg[51]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[51]) );
  DFF \sreg_reg[50]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[50]) );
  DFF \sreg_reg[49]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[49]) );
  DFF \sreg_reg[48]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[48]) );
  DFF \sreg_reg[47]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[46]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[45]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[44]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[43]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[42]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[41]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[40]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[39]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[38]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[37]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[36]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[35]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[34]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[33]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[32]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[31]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[30]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[29]  ( .D(c[31]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[28]  ( .D(c[30]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[27]  ( .D(c[29]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[26]  ( .D(c[28]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[25]  ( .D(c[27]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[24]  ( .D(c[26]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[23]  ( .D(c[25]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[22]  ( .D(c[24]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[21]  ( .D(c[23]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[20]  ( .D(c[22]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[19]  ( .D(c[21]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[18]  ( .D(c[20]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[17]  ( .D(c[19]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[16]  ( .D(c[18]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[15]  ( .D(c[17]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[14]  ( .D(c[16]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[13]  ( .D(c[15]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[12]  ( .D(c[14]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[11]  ( .D(c[13]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[10]  ( .D(c[12]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[9]  ( .D(c[11]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[8]  ( .D(c[10]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[7]  ( .D(c[9]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[6]  ( .D(c[8]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[5]  ( .D(c[7]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[4]  ( .D(c[6]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[3]  ( .D(c[5]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[2]  ( .D(c[4]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[1]  ( .D(c[3]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[0]  ( .D(c[2]), .CLK(clk), .RST(rst), .Q(c[0]) );
  NAND U5 ( .A(n1629), .B(n1628), .Z(n1) );
  XOR U6 ( .A(n1628), .B(n1629), .Z(n2) );
  NAND U7 ( .A(n2), .B(n1627), .Z(n3) );
  NAND U8 ( .A(n1), .B(n3), .Z(n1636) );
  NAND U9 ( .A(n796), .B(n795), .Z(n4) );
  XOR U10 ( .A(n795), .B(n796), .Z(n5) );
  NAND U11 ( .A(n5), .B(n794), .Z(n6) );
  NAND U12 ( .A(n4), .B(n6), .Z(n802) );
  NAND U13 ( .A(n817), .B(n815), .Z(n7) );
  XOR U14 ( .A(n815), .B(n817), .Z(n8) );
  NAND U15 ( .A(n8), .B(n816), .Z(n9) );
  NAND U16 ( .A(n7), .B(n9), .Z(n823) );
  NAND U17 ( .A(n838), .B(n837), .Z(n10) );
  XOR U18 ( .A(n837), .B(n838), .Z(n11) );
  NAND U19 ( .A(n11), .B(n836), .Z(n12) );
  NAND U20 ( .A(n10), .B(n12), .Z(n844) );
  NAND U21 ( .A(n859), .B(n858), .Z(n13) );
  XOR U22 ( .A(n858), .B(n859), .Z(n14) );
  NAND U23 ( .A(n14), .B(n857), .Z(n15) );
  NAND U24 ( .A(n13), .B(n15), .Z(n865) );
  NAND U25 ( .A(n880), .B(n879), .Z(n16) );
  XOR U26 ( .A(n879), .B(n880), .Z(n17) );
  NAND U27 ( .A(n17), .B(n878), .Z(n18) );
  NAND U28 ( .A(n16), .B(n18), .Z(n886) );
  NAND U29 ( .A(n901), .B(n899), .Z(n19) );
  XOR U30 ( .A(n899), .B(n901), .Z(n20) );
  NAND U31 ( .A(n20), .B(n900), .Z(n21) );
  NAND U32 ( .A(n19), .B(n21), .Z(n907) );
  NAND U33 ( .A(n922), .B(n921), .Z(n22) );
  XOR U34 ( .A(n921), .B(n922), .Z(n23) );
  NAND U35 ( .A(n23), .B(n920), .Z(n24) );
  NAND U36 ( .A(n22), .B(n24), .Z(n928) );
  NAND U37 ( .A(n943), .B(n942), .Z(n25) );
  XOR U38 ( .A(n942), .B(n943), .Z(n26) );
  NAND U39 ( .A(n26), .B(n941), .Z(n27) );
  NAND U40 ( .A(n25), .B(n27), .Z(n949) );
  NAND U41 ( .A(n964), .B(n963), .Z(n28) );
  XOR U42 ( .A(n963), .B(n964), .Z(n29) );
  NAND U43 ( .A(n29), .B(n962), .Z(n30) );
  NAND U44 ( .A(n28), .B(n30), .Z(n970) );
  NAND U45 ( .A(n985), .B(n984), .Z(n31) );
  XOR U46 ( .A(n984), .B(n985), .Z(n32) );
  NAND U47 ( .A(n32), .B(n983), .Z(n33) );
  NAND U48 ( .A(n31), .B(n33), .Z(n991) );
  NAND U49 ( .A(n1006), .B(n1005), .Z(n34) );
  XOR U50 ( .A(n1005), .B(n1006), .Z(n35) );
  NAND U51 ( .A(n35), .B(n1004), .Z(n36) );
  NAND U52 ( .A(n34), .B(n36), .Z(n1012) );
  NAND U53 ( .A(n1027), .B(n1026), .Z(n37) );
  XOR U54 ( .A(n1026), .B(n1027), .Z(n38) );
  NAND U55 ( .A(n38), .B(n1025), .Z(n39) );
  NAND U56 ( .A(n37), .B(n39), .Z(n1033) );
  NAND U57 ( .A(n1048), .B(n1047), .Z(n40) );
  XOR U58 ( .A(n1047), .B(n1048), .Z(n41) );
  NAND U59 ( .A(n41), .B(n1046), .Z(n42) );
  NAND U60 ( .A(n40), .B(n42), .Z(n1054) );
  NAND U61 ( .A(n1069), .B(n1068), .Z(n43) );
  XOR U62 ( .A(n1068), .B(n1069), .Z(n44) );
  NAND U63 ( .A(n44), .B(n1067), .Z(n45) );
  NAND U64 ( .A(n43), .B(n45), .Z(n1075) );
  NAND U65 ( .A(n1090), .B(n1089), .Z(n46) );
  XOR U66 ( .A(n1089), .B(n1090), .Z(n47) );
  NAND U67 ( .A(n47), .B(n1088), .Z(n48) );
  NAND U68 ( .A(n46), .B(n48), .Z(n1096) );
  NAND U69 ( .A(n1111), .B(n1110), .Z(n49) );
  XOR U70 ( .A(n1110), .B(n1111), .Z(n50) );
  NAND U71 ( .A(n50), .B(n1109), .Z(n51) );
  NAND U72 ( .A(n49), .B(n51), .Z(n1117) );
  NAND U73 ( .A(n1132), .B(n1131), .Z(n52) );
  XOR U74 ( .A(n1131), .B(n1132), .Z(n53) );
  NAND U75 ( .A(n53), .B(n1130), .Z(n54) );
  NAND U76 ( .A(n52), .B(n54), .Z(n1138) );
  NAND U77 ( .A(n1153), .B(n1152), .Z(n55) );
  XOR U78 ( .A(n1152), .B(n1153), .Z(n56) );
  NAND U79 ( .A(n56), .B(n1151), .Z(n57) );
  NAND U80 ( .A(n55), .B(n57), .Z(n1159) );
  NAND U81 ( .A(n1174), .B(n1173), .Z(n58) );
  XOR U82 ( .A(n1173), .B(n1174), .Z(n59) );
  NAND U83 ( .A(n59), .B(n1172), .Z(n60) );
  NAND U84 ( .A(n58), .B(n60), .Z(n1180) );
  NAND U85 ( .A(n1195), .B(n1194), .Z(n61) );
  XOR U86 ( .A(n1194), .B(n1195), .Z(n62) );
  NAND U87 ( .A(n62), .B(n1193), .Z(n63) );
  NAND U88 ( .A(n61), .B(n63), .Z(n1201) );
  NAND U89 ( .A(n1216), .B(n1215), .Z(n64) );
  XOR U90 ( .A(n1215), .B(n1216), .Z(n65) );
  NAND U91 ( .A(n65), .B(n1214), .Z(n66) );
  NAND U92 ( .A(n64), .B(n66), .Z(n1222) );
  NAND U93 ( .A(n1237), .B(n1236), .Z(n67) );
  XOR U94 ( .A(n1236), .B(n1237), .Z(n68) );
  NAND U95 ( .A(n68), .B(n1235), .Z(n69) );
  NAND U96 ( .A(n67), .B(n69), .Z(n1243) );
  NAND U97 ( .A(n1258), .B(n1257), .Z(n70) );
  XOR U98 ( .A(n1257), .B(n1258), .Z(n71) );
  NAND U99 ( .A(n71), .B(n1256), .Z(n72) );
  NAND U100 ( .A(n70), .B(n72), .Z(n1264) );
  NAND U101 ( .A(n1279), .B(n1278), .Z(n73) );
  XOR U102 ( .A(n1278), .B(n1279), .Z(n74) );
  NAND U103 ( .A(n74), .B(n1277), .Z(n75) );
  NAND U104 ( .A(n73), .B(n75), .Z(n1285) );
  NAND U105 ( .A(n1300), .B(n1299), .Z(n76) );
  XOR U106 ( .A(n1299), .B(n1300), .Z(n77) );
  NAND U107 ( .A(n77), .B(n1298), .Z(n78) );
  NAND U108 ( .A(n76), .B(n78), .Z(n1306) );
  NAND U109 ( .A(n1321), .B(n1320), .Z(n79) );
  XOR U110 ( .A(n1320), .B(n1321), .Z(n80) );
  NAND U111 ( .A(n80), .B(n1319), .Z(n81) );
  NAND U112 ( .A(n79), .B(n81), .Z(n1327) );
  NAND U113 ( .A(n1342), .B(n1341), .Z(n82) );
  XOR U114 ( .A(n1341), .B(n1342), .Z(n83) );
  NAND U115 ( .A(n83), .B(n1340), .Z(n84) );
  NAND U116 ( .A(n82), .B(n84), .Z(n1348) );
  NAND U117 ( .A(n1363), .B(n1362), .Z(n85) );
  XOR U118 ( .A(n1362), .B(n1363), .Z(n86) );
  NAND U119 ( .A(n86), .B(n1361), .Z(n87) );
  NAND U120 ( .A(n85), .B(n87), .Z(n1369) );
  NAND U121 ( .A(n1384), .B(n1383), .Z(n88) );
  XOR U122 ( .A(n1383), .B(n1384), .Z(n89) );
  NAND U123 ( .A(n89), .B(n1382), .Z(n90) );
  NAND U124 ( .A(n88), .B(n90), .Z(n1390) );
  NAND U125 ( .A(n1405), .B(n1404), .Z(n91) );
  XOR U126 ( .A(n1404), .B(n1405), .Z(n92) );
  NAND U127 ( .A(n92), .B(n1403), .Z(n93) );
  NAND U128 ( .A(n91), .B(n93), .Z(n1411) );
  NAND U129 ( .A(n1426), .B(n1425), .Z(n94) );
  XOR U130 ( .A(n1425), .B(n1426), .Z(n95) );
  NAND U131 ( .A(n95), .B(n1424), .Z(n96) );
  NAND U132 ( .A(n94), .B(n96), .Z(n1432) );
  NAND U133 ( .A(n1447), .B(n1446), .Z(n97) );
  XOR U134 ( .A(n1446), .B(n1447), .Z(n98) );
  NAND U135 ( .A(n98), .B(n1445), .Z(n99) );
  NAND U136 ( .A(n97), .B(n99), .Z(n1453) );
  NAND U137 ( .A(n1468), .B(n1467), .Z(n100) );
  XOR U138 ( .A(n1467), .B(n1468), .Z(n101) );
  NAND U139 ( .A(n101), .B(n1466), .Z(n102) );
  NAND U140 ( .A(n100), .B(n102), .Z(n1474) );
  NAND U141 ( .A(n1489), .B(n1488), .Z(n103) );
  XOR U142 ( .A(n1488), .B(n1489), .Z(n104) );
  NAND U143 ( .A(n104), .B(n1487), .Z(n105) );
  NAND U144 ( .A(n103), .B(n105), .Z(n1495) );
  NAND U145 ( .A(n1510), .B(n1509), .Z(n106) );
  XOR U146 ( .A(n1509), .B(n1510), .Z(n107) );
  NAND U147 ( .A(n107), .B(n1508), .Z(n108) );
  NAND U148 ( .A(n106), .B(n108), .Z(n1516) );
  NAND U149 ( .A(n1531), .B(n1530), .Z(n109) );
  XOR U150 ( .A(n1530), .B(n1531), .Z(n110) );
  NAND U151 ( .A(n110), .B(n1529), .Z(n111) );
  NAND U152 ( .A(n109), .B(n111), .Z(n1537) );
  NAND U153 ( .A(n1552), .B(n1551), .Z(n112) );
  XOR U154 ( .A(n1551), .B(n1552), .Z(n113) );
  NAND U155 ( .A(n113), .B(n1550), .Z(n114) );
  NAND U156 ( .A(n112), .B(n114), .Z(n1558) );
  NAND U157 ( .A(n1573), .B(n1572), .Z(n115) );
  XOR U158 ( .A(n1572), .B(n1573), .Z(n116) );
  NAND U159 ( .A(n116), .B(n1571), .Z(n117) );
  NAND U160 ( .A(n115), .B(n117), .Z(n1579) );
  NAND U161 ( .A(n1594), .B(n1593), .Z(n118) );
  XOR U162 ( .A(n1593), .B(n1594), .Z(n119) );
  NAND U163 ( .A(n119), .B(n1592), .Z(n120) );
  NAND U164 ( .A(n118), .B(n120), .Z(n1600) );
  NAND U165 ( .A(n1615), .B(n1614), .Z(n121) );
  XOR U166 ( .A(n1614), .B(n1615), .Z(n122) );
  NAND U167 ( .A(n122), .B(n1613), .Z(n123) );
  NAND U168 ( .A(n121), .B(n123), .Z(n1621) );
  XOR U169 ( .A(n1637), .B(n1635), .Z(n124) );
  NAND U170 ( .A(n124), .B(n1636), .Z(n125) );
  NAND U171 ( .A(n1637), .B(n1635), .Z(n126) );
  AND U172 ( .A(n125), .B(n126), .Z(n1646) );
  NAND U173 ( .A(sreg[128]), .B(n764), .Z(n127) );
  XOR U174 ( .A(n764), .B(sreg[128]), .Z(n128) );
  NANDN U175 ( .A(n765), .B(n128), .Z(n129) );
  NAND U176 ( .A(n127), .B(n129), .Z(n777) );
  NAND U177 ( .A(sreg[131]), .B(n791), .Z(n130) );
  XOR U178 ( .A(n791), .B(sreg[131]), .Z(n131) );
  NANDN U179 ( .A(n792), .B(n131), .Z(n132) );
  NAND U180 ( .A(n130), .B(n132), .Z(n798) );
  NAND U181 ( .A(sreg[134]), .B(n813), .Z(n133) );
  XOR U182 ( .A(n813), .B(sreg[134]), .Z(n134) );
  NAND U183 ( .A(n134), .B(n812), .Z(n135) );
  NAND U184 ( .A(n133), .B(n135), .Z(n819) );
  NAND U185 ( .A(sreg[137]), .B(n834), .Z(n136) );
  XOR U186 ( .A(n834), .B(sreg[137]), .Z(n137) );
  NAND U187 ( .A(n137), .B(n833), .Z(n138) );
  NAND U188 ( .A(n136), .B(n138), .Z(n840) );
  NAND U189 ( .A(sreg[140]), .B(n855), .Z(n139) );
  XOR U190 ( .A(n855), .B(sreg[140]), .Z(n140) );
  NAND U191 ( .A(n140), .B(n854), .Z(n141) );
  NAND U192 ( .A(n139), .B(n141), .Z(n861) );
  NAND U193 ( .A(sreg[143]), .B(n875), .Z(n142) );
  XOR U194 ( .A(n875), .B(sreg[143]), .Z(n143) );
  NANDN U195 ( .A(n876), .B(n143), .Z(n144) );
  NAND U196 ( .A(n142), .B(n144), .Z(n882) );
  NAND U197 ( .A(sreg[146]), .B(n897), .Z(n145) );
  XOR U198 ( .A(n897), .B(sreg[146]), .Z(n146) );
  NAND U199 ( .A(n146), .B(n896), .Z(n147) );
  NAND U200 ( .A(n145), .B(n147), .Z(n903) );
  NAND U201 ( .A(sreg[149]), .B(n918), .Z(n148) );
  XOR U202 ( .A(n918), .B(sreg[149]), .Z(n149) );
  NAND U203 ( .A(n149), .B(n917), .Z(n150) );
  NAND U204 ( .A(n148), .B(n150), .Z(n924) );
  NAND U205 ( .A(sreg[152]), .B(n939), .Z(n151) );
  XOR U206 ( .A(n939), .B(sreg[152]), .Z(n152) );
  NAND U207 ( .A(n152), .B(n938), .Z(n153) );
  NAND U208 ( .A(n151), .B(n153), .Z(n945) );
  NAND U209 ( .A(sreg[155]), .B(n960), .Z(n154) );
  XOR U210 ( .A(n960), .B(sreg[155]), .Z(n155) );
  NAND U211 ( .A(n155), .B(n959), .Z(n156) );
  NAND U212 ( .A(n154), .B(n156), .Z(n966) );
  NAND U213 ( .A(sreg[158]), .B(n981), .Z(n157) );
  XOR U214 ( .A(n981), .B(sreg[158]), .Z(n158) );
  NAND U215 ( .A(n158), .B(n980), .Z(n159) );
  NAND U216 ( .A(n157), .B(n159), .Z(n987) );
  NAND U217 ( .A(sreg[161]), .B(n1002), .Z(n160) );
  XOR U218 ( .A(n1002), .B(sreg[161]), .Z(n161) );
  NAND U219 ( .A(n161), .B(n1001), .Z(n162) );
  NAND U220 ( .A(n160), .B(n162), .Z(n1008) );
  NAND U221 ( .A(sreg[164]), .B(n1023), .Z(n163) );
  XOR U222 ( .A(n1023), .B(sreg[164]), .Z(n164) );
  NAND U223 ( .A(n164), .B(n1022), .Z(n165) );
  NAND U224 ( .A(n163), .B(n165), .Z(n1029) );
  NAND U225 ( .A(sreg[167]), .B(n1044), .Z(n166) );
  XOR U226 ( .A(n1044), .B(sreg[167]), .Z(n167) );
  NAND U227 ( .A(n167), .B(n1043), .Z(n168) );
  NAND U228 ( .A(n166), .B(n168), .Z(n1050) );
  NAND U229 ( .A(sreg[170]), .B(n1065), .Z(n169) );
  XOR U230 ( .A(n1065), .B(sreg[170]), .Z(n170) );
  NAND U231 ( .A(n170), .B(n1064), .Z(n171) );
  NAND U232 ( .A(n169), .B(n171), .Z(n1071) );
  NAND U233 ( .A(sreg[173]), .B(n1086), .Z(n172) );
  XOR U234 ( .A(n1086), .B(sreg[173]), .Z(n173) );
  NAND U235 ( .A(n173), .B(n1085), .Z(n174) );
  NAND U236 ( .A(n172), .B(n174), .Z(n1092) );
  NAND U237 ( .A(sreg[176]), .B(n1107), .Z(n175) );
  XOR U238 ( .A(n1107), .B(sreg[176]), .Z(n176) );
  NAND U239 ( .A(n176), .B(n1106), .Z(n177) );
  NAND U240 ( .A(n175), .B(n177), .Z(n1113) );
  NAND U241 ( .A(sreg[179]), .B(n1128), .Z(n178) );
  XOR U242 ( .A(n1128), .B(sreg[179]), .Z(n179) );
  NAND U243 ( .A(n179), .B(n1127), .Z(n180) );
  NAND U244 ( .A(n178), .B(n180), .Z(n1134) );
  NAND U245 ( .A(sreg[182]), .B(n1149), .Z(n181) );
  XOR U246 ( .A(n1149), .B(sreg[182]), .Z(n182) );
  NAND U247 ( .A(n182), .B(n1148), .Z(n183) );
  NAND U248 ( .A(n181), .B(n183), .Z(n1155) );
  NAND U249 ( .A(sreg[185]), .B(n1170), .Z(n184) );
  XOR U250 ( .A(n1170), .B(sreg[185]), .Z(n185) );
  NAND U251 ( .A(n185), .B(n1169), .Z(n186) );
  NAND U252 ( .A(n184), .B(n186), .Z(n1176) );
  NAND U253 ( .A(sreg[188]), .B(n1191), .Z(n187) );
  XOR U254 ( .A(n1191), .B(sreg[188]), .Z(n188) );
  NAND U255 ( .A(n188), .B(n1190), .Z(n189) );
  NAND U256 ( .A(n187), .B(n189), .Z(n1197) );
  NAND U257 ( .A(sreg[191]), .B(n1212), .Z(n190) );
  XOR U258 ( .A(n1212), .B(sreg[191]), .Z(n191) );
  NAND U259 ( .A(n191), .B(n1211), .Z(n192) );
  NAND U260 ( .A(n190), .B(n192), .Z(n1218) );
  NAND U261 ( .A(sreg[194]), .B(n1233), .Z(n193) );
  XOR U262 ( .A(n1233), .B(sreg[194]), .Z(n194) );
  NAND U263 ( .A(n194), .B(n1232), .Z(n195) );
  NAND U264 ( .A(n193), .B(n195), .Z(n1239) );
  NAND U265 ( .A(sreg[197]), .B(n1254), .Z(n196) );
  XOR U266 ( .A(n1254), .B(sreg[197]), .Z(n197) );
  NAND U267 ( .A(n197), .B(n1253), .Z(n198) );
  NAND U268 ( .A(n196), .B(n198), .Z(n1260) );
  NAND U269 ( .A(sreg[200]), .B(n1275), .Z(n199) );
  XOR U270 ( .A(n1275), .B(sreg[200]), .Z(n200) );
  NAND U271 ( .A(n200), .B(n1274), .Z(n201) );
  NAND U272 ( .A(n199), .B(n201), .Z(n1281) );
  NAND U273 ( .A(sreg[203]), .B(n1296), .Z(n202) );
  XOR U274 ( .A(n1296), .B(sreg[203]), .Z(n203) );
  NAND U275 ( .A(n203), .B(n1295), .Z(n204) );
  NAND U276 ( .A(n202), .B(n204), .Z(n1302) );
  NAND U277 ( .A(sreg[206]), .B(n1317), .Z(n205) );
  XOR U278 ( .A(n1317), .B(sreg[206]), .Z(n206) );
  NAND U279 ( .A(n206), .B(n1316), .Z(n207) );
  NAND U280 ( .A(n205), .B(n207), .Z(n1323) );
  NAND U281 ( .A(sreg[209]), .B(n1338), .Z(n208) );
  XOR U282 ( .A(n1338), .B(sreg[209]), .Z(n209) );
  NAND U283 ( .A(n209), .B(n1337), .Z(n210) );
  NAND U284 ( .A(n208), .B(n210), .Z(n1344) );
  NAND U285 ( .A(sreg[212]), .B(n1359), .Z(n211) );
  XOR U286 ( .A(n1359), .B(sreg[212]), .Z(n212) );
  NAND U287 ( .A(n212), .B(n1358), .Z(n213) );
  NAND U288 ( .A(n211), .B(n213), .Z(n1365) );
  NAND U289 ( .A(sreg[215]), .B(n1380), .Z(n214) );
  XOR U290 ( .A(n1380), .B(sreg[215]), .Z(n215) );
  NAND U291 ( .A(n215), .B(n1379), .Z(n216) );
  NAND U292 ( .A(n214), .B(n216), .Z(n1386) );
  NAND U293 ( .A(sreg[218]), .B(n1401), .Z(n217) );
  XOR U294 ( .A(n1401), .B(sreg[218]), .Z(n218) );
  NAND U295 ( .A(n218), .B(n1400), .Z(n219) );
  NAND U296 ( .A(n217), .B(n219), .Z(n1407) );
  NAND U297 ( .A(sreg[221]), .B(n1422), .Z(n220) );
  XOR U298 ( .A(n1422), .B(sreg[221]), .Z(n221) );
  NAND U299 ( .A(n221), .B(n1421), .Z(n222) );
  NAND U300 ( .A(n220), .B(n222), .Z(n1428) );
  NAND U301 ( .A(sreg[224]), .B(n1443), .Z(n223) );
  XOR U302 ( .A(n1443), .B(sreg[224]), .Z(n224) );
  NAND U303 ( .A(n224), .B(n1442), .Z(n225) );
  NAND U304 ( .A(n223), .B(n225), .Z(n1449) );
  NAND U305 ( .A(sreg[227]), .B(n1464), .Z(n226) );
  XOR U306 ( .A(n1464), .B(sreg[227]), .Z(n227) );
  NAND U307 ( .A(n227), .B(n1463), .Z(n228) );
  NAND U308 ( .A(n226), .B(n228), .Z(n1470) );
  NAND U309 ( .A(sreg[230]), .B(n1485), .Z(n229) );
  XOR U310 ( .A(n1485), .B(sreg[230]), .Z(n230) );
  NAND U311 ( .A(n230), .B(n1484), .Z(n231) );
  NAND U312 ( .A(n229), .B(n231), .Z(n1491) );
  NAND U313 ( .A(sreg[233]), .B(n1506), .Z(n232) );
  XOR U314 ( .A(n1506), .B(sreg[233]), .Z(n233) );
  NAND U315 ( .A(n233), .B(n1505), .Z(n234) );
  NAND U316 ( .A(n232), .B(n234), .Z(n1512) );
  NAND U317 ( .A(sreg[236]), .B(n1527), .Z(n235) );
  XOR U318 ( .A(n1527), .B(sreg[236]), .Z(n236) );
  NAND U319 ( .A(n236), .B(n1526), .Z(n237) );
  NAND U320 ( .A(n235), .B(n237), .Z(n1533) );
  NAND U321 ( .A(sreg[239]), .B(n1548), .Z(n238) );
  XOR U322 ( .A(n1548), .B(sreg[239]), .Z(n239) );
  NAND U323 ( .A(n239), .B(n1547), .Z(n240) );
  NAND U324 ( .A(n238), .B(n240), .Z(n1554) );
  NAND U325 ( .A(sreg[242]), .B(n1569), .Z(n241) );
  XOR U326 ( .A(n1569), .B(sreg[242]), .Z(n242) );
  NAND U327 ( .A(n242), .B(n1568), .Z(n243) );
  NAND U328 ( .A(n241), .B(n243), .Z(n1575) );
  NAND U329 ( .A(sreg[245]), .B(n1590), .Z(n244) );
  XOR U330 ( .A(n1590), .B(sreg[245]), .Z(n245) );
  NAND U331 ( .A(n245), .B(n1589), .Z(n246) );
  NAND U332 ( .A(n244), .B(n246), .Z(n1596) );
  NAND U333 ( .A(sreg[248]), .B(n1611), .Z(n247) );
  XOR U334 ( .A(n1611), .B(sreg[248]), .Z(n248) );
  NAND U335 ( .A(n248), .B(n1610), .Z(n249) );
  NAND U336 ( .A(n247), .B(n249), .Z(n1617) );
  NAND U337 ( .A(sreg[251]), .B(n1632), .Z(n250) );
  XOR U338 ( .A(n1632), .B(sreg[251]), .Z(n251) );
  NAND U339 ( .A(n251), .B(n1631), .Z(n252) );
  NAND U340 ( .A(n250), .B(n252), .Z(n1638) );
  NAND U341 ( .A(n782), .B(n781), .Z(n253) );
  XOR U342 ( .A(n781), .B(n782), .Z(n254) );
  NANDN U343 ( .A(n780), .B(n254), .Z(n255) );
  NAND U344 ( .A(n253), .B(n255), .Z(n788) );
  NAND U345 ( .A(n803), .B(n802), .Z(n256) );
  XOR U346 ( .A(n802), .B(n803), .Z(n257) );
  NAND U347 ( .A(n257), .B(n801), .Z(n258) );
  NAND U348 ( .A(n256), .B(n258), .Z(n809) );
  NAND U349 ( .A(n824), .B(n823), .Z(n259) );
  XOR U350 ( .A(n823), .B(n824), .Z(n260) );
  NAND U351 ( .A(n260), .B(n822), .Z(n261) );
  NAND U352 ( .A(n259), .B(n261), .Z(n830) );
  NAND U353 ( .A(n845), .B(n843), .Z(n262) );
  XOR U354 ( .A(n843), .B(n845), .Z(n263) );
  NAND U355 ( .A(n263), .B(n844), .Z(n264) );
  NAND U356 ( .A(n262), .B(n264), .Z(n851) );
  NAND U357 ( .A(n866), .B(n865), .Z(n265) );
  XOR U358 ( .A(n865), .B(n866), .Z(n266) );
  NAND U359 ( .A(n266), .B(n864), .Z(n267) );
  NAND U360 ( .A(n265), .B(n267), .Z(n872) );
  NAND U361 ( .A(n887), .B(n886), .Z(n268) );
  XOR U362 ( .A(n886), .B(n887), .Z(n269) );
  NAND U363 ( .A(n269), .B(n885), .Z(n270) );
  NAND U364 ( .A(n268), .B(n270), .Z(n893) );
  NAND U365 ( .A(n908), .B(n907), .Z(n271) );
  XOR U366 ( .A(n907), .B(n908), .Z(n272) );
  NAND U367 ( .A(n272), .B(n906), .Z(n273) );
  NAND U368 ( .A(n271), .B(n273), .Z(n914) );
  NAND U369 ( .A(n929), .B(n928), .Z(n274) );
  XOR U370 ( .A(n928), .B(n929), .Z(n275) );
  NAND U371 ( .A(n275), .B(n927), .Z(n276) );
  NAND U372 ( .A(n274), .B(n276), .Z(n935) );
  NAND U373 ( .A(n950), .B(n949), .Z(n277) );
  XOR U374 ( .A(n949), .B(n950), .Z(n278) );
  NAND U375 ( .A(n278), .B(n948), .Z(n279) );
  NAND U376 ( .A(n277), .B(n279), .Z(n956) );
  NAND U377 ( .A(n971), .B(n970), .Z(n280) );
  XOR U378 ( .A(n970), .B(n971), .Z(n281) );
  NAND U379 ( .A(n281), .B(n969), .Z(n282) );
  NAND U380 ( .A(n280), .B(n282), .Z(n977) );
  NAND U381 ( .A(n992), .B(n991), .Z(n283) );
  XOR U382 ( .A(n991), .B(n992), .Z(n284) );
  NAND U383 ( .A(n284), .B(n990), .Z(n285) );
  NAND U384 ( .A(n283), .B(n285), .Z(n998) );
  NAND U385 ( .A(n1013), .B(n1012), .Z(n286) );
  XOR U386 ( .A(n1012), .B(n1013), .Z(n287) );
  NAND U387 ( .A(n287), .B(n1011), .Z(n288) );
  NAND U388 ( .A(n286), .B(n288), .Z(n1019) );
  NAND U389 ( .A(n1034), .B(n1033), .Z(n289) );
  XOR U390 ( .A(n1033), .B(n1034), .Z(n290) );
  NAND U391 ( .A(n290), .B(n1032), .Z(n291) );
  NAND U392 ( .A(n289), .B(n291), .Z(n1040) );
  NAND U393 ( .A(n1055), .B(n1054), .Z(n292) );
  XOR U394 ( .A(n1054), .B(n1055), .Z(n293) );
  NAND U395 ( .A(n293), .B(n1053), .Z(n294) );
  NAND U396 ( .A(n292), .B(n294), .Z(n1061) );
  NAND U397 ( .A(n1076), .B(n1075), .Z(n295) );
  XOR U398 ( .A(n1075), .B(n1076), .Z(n296) );
  NAND U399 ( .A(n296), .B(n1074), .Z(n297) );
  NAND U400 ( .A(n295), .B(n297), .Z(n1082) );
  NAND U401 ( .A(n1097), .B(n1096), .Z(n298) );
  XOR U402 ( .A(n1096), .B(n1097), .Z(n299) );
  NAND U403 ( .A(n299), .B(n1095), .Z(n300) );
  NAND U404 ( .A(n298), .B(n300), .Z(n1103) );
  NAND U405 ( .A(n1118), .B(n1117), .Z(n301) );
  XOR U406 ( .A(n1117), .B(n1118), .Z(n302) );
  NAND U407 ( .A(n302), .B(n1116), .Z(n303) );
  NAND U408 ( .A(n301), .B(n303), .Z(n1124) );
  NAND U409 ( .A(n1139), .B(n1138), .Z(n304) );
  XOR U410 ( .A(n1138), .B(n1139), .Z(n305) );
  NAND U411 ( .A(n305), .B(n1137), .Z(n306) );
  NAND U412 ( .A(n304), .B(n306), .Z(n1145) );
  NAND U413 ( .A(n1160), .B(n1159), .Z(n307) );
  XOR U414 ( .A(n1159), .B(n1160), .Z(n308) );
  NAND U415 ( .A(n308), .B(n1158), .Z(n309) );
  NAND U416 ( .A(n307), .B(n309), .Z(n1166) );
  NAND U417 ( .A(n1181), .B(n1180), .Z(n310) );
  XOR U418 ( .A(n1180), .B(n1181), .Z(n311) );
  NAND U419 ( .A(n311), .B(n1179), .Z(n312) );
  NAND U420 ( .A(n310), .B(n312), .Z(n1187) );
  NAND U421 ( .A(n1202), .B(n1201), .Z(n313) );
  XOR U422 ( .A(n1201), .B(n1202), .Z(n314) );
  NAND U423 ( .A(n314), .B(n1200), .Z(n315) );
  NAND U424 ( .A(n313), .B(n315), .Z(n1208) );
  NAND U425 ( .A(n1223), .B(n1222), .Z(n316) );
  XOR U426 ( .A(n1222), .B(n1223), .Z(n317) );
  NAND U427 ( .A(n317), .B(n1221), .Z(n318) );
  NAND U428 ( .A(n316), .B(n318), .Z(n1229) );
  NAND U429 ( .A(n1244), .B(n1243), .Z(n319) );
  XOR U430 ( .A(n1243), .B(n1244), .Z(n320) );
  NAND U431 ( .A(n320), .B(n1242), .Z(n321) );
  NAND U432 ( .A(n319), .B(n321), .Z(n1250) );
  NAND U433 ( .A(n1265), .B(n1264), .Z(n322) );
  XOR U434 ( .A(n1264), .B(n1265), .Z(n323) );
  NAND U435 ( .A(n323), .B(n1263), .Z(n324) );
  NAND U436 ( .A(n322), .B(n324), .Z(n1271) );
  NAND U437 ( .A(n1286), .B(n1285), .Z(n325) );
  XOR U438 ( .A(n1285), .B(n1286), .Z(n326) );
  NAND U439 ( .A(n326), .B(n1284), .Z(n327) );
  NAND U440 ( .A(n325), .B(n327), .Z(n1292) );
  NAND U441 ( .A(n1307), .B(n1306), .Z(n328) );
  XOR U442 ( .A(n1306), .B(n1307), .Z(n329) );
  NAND U443 ( .A(n329), .B(n1305), .Z(n330) );
  NAND U444 ( .A(n328), .B(n330), .Z(n1313) );
  NAND U445 ( .A(n1328), .B(n1327), .Z(n331) );
  XOR U446 ( .A(n1327), .B(n1328), .Z(n332) );
  NAND U447 ( .A(n332), .B(n1326), .Z(n333) );
  NAND U448 ( .A(n331), .B(n333), .Z(n1334) );
  NAND U449 ( .A(n1349), .B(n1348), .Z(n334) );
  XOR U450 ( .A(n1348), .B(n1349), .Z(n335) );
  NAND U451 ( .A(n335), .B(n1347), .Z(n336) );
  NAND U452 ( .A(n334), .B(n336), .Z(n1355) );
  NAND U453 ( .A(n1370), .B(n1369), .Z(n337) );
  XOR U454 ( .A(n1369), .B(n1370), .Z(n338) );
  NAND U455 ( .A(n338), .B(n1368), .Z(n339) );
  NAND U456 ( .A(n337), .B(n339), .Z(n1376) );
  NAND U457 ( .A(n1391), .B(n1390), .Z(n340) );
  XOR U458 ( .A(n1390), .B(n1391), .Z(n341) );
  NAND U459 ( .A(n341), .B(n1389), .Z(n342) );
  NAND U460 ( .A(n340), .B(n342), .Z(n1397) );
  NAND U461 ( .A(n1412), .B(n1411), .Z(n343) );
  XOR U462 ( .A(n1411), .B(n1412), .Z(n344) );
  NAND U463 ( .A(n344), .B(n1410), .Z(n345) );
  NAND U464 ( .A(n343), .B(n345), .Z(n1418) );
  NAND U465 ( .A(n1433), .B(n1432), .Z(n346) );
  XOR U466 ( .A(n1432), .B(n1433), .Z(n347) );
  NAND U467 ( .A(n347), .B(n1431), .Z(n348) );
  NAND U468 ( .A(n346), .B(n348), .Z(n1439) );
  NAND U469 ( .A(n1454), .B(n1453), .Z(n349) );
  XOR U470 ( .A(n1453), .B(n1454), .Z(n350) );
  NAND U471 ( .A(n350), .B(n1452), .Z(n351) );
  NAND U472 ( .A(n349), .B(n351), .Z(n1460) );
  NAND U473 ( .A(n1475), .B(n1474), .Z(n352) );
  XOR U474 ( .A(n1474), .B(n1475), .Z(n353) );
  NAND U475 ( .A(n353), .B(n1473), .Z(n354) );
  NAND U476 ( .A(n352), .B(n354), .Z(n1481) );
  NAND U477 ( .A(n1496), .B(n1495), .Z(n355) );
  XOR U478 ( .A(n1495), .B(n1496), .Z(n356) );
  NAND U479 ( .A(n356), .B(n1494), .Z(n357) );
  NAND U480 ( .A(n355), .B(n357), .Z(n1502) );
  NAND U481 ( .A(n1517), .B(n1516), .Z(n358) );
  XOR U482 ( .A(n1516), .B(n1517), .Z(n359) );
  NAND U483 ( .A(n359), .B(n1515), .Z(n360) );
  NAND U484 ( .A(n358), .B(n360), .Z(n1523) );
  NAND U485 ( .A(n1538), .B(n1537), .Z(n361) );
  XOR U486 ( .A(n1537), .B(n1538), .Z(n362) );
  NAND U487 ( .A(n362), .B(n1536), .Z(n363) );
  NAND U488 ( .A(n361), .B(n363), .Z(n1544) );
  NAND U489 ( .A(n1559), .B(n1558), .Z(n364) );
  XOR U490 ( .A(n1558), .B(n1559), .Z(n365) );
  NAND U491 ( .A(n365), .B(n1557), .Z(n366) );
  NAND U492 ( .A(n364), .B(n366), .Z(n1565) );
  NAND U493 ( .A(n1580), .B(n1579), .Z(n367) );
  XOR U494 ( .A(n1579), .B(n1580), .Z(n368) );
  NAND U495 ( .A(n368), .B(n1578), .Z(n369) );
  NAND U496 ( .A(n367), .B(n369), .Z(n1586) );
  NAND U497 ( .A(n1601), .B(n1600), .Z(n370) );
  XOR U498 ( .A(n1600), .B(n1601), .Z(n371) );
  NAND U499 ( .A(n371), .B(n1599), .Z(n372) );
  NAND U500 ( .A(n370), .B(n372), .Z(n1607) );
  NAND U501 ( .A(n1622), .B(n1621), .Z(n373) );
  XOR U502 ( .A(n1621), .B(n1622), .Z(n374) );
  NAND U503 ( .A(n374), .B(n1620), .Z(n375) );
  NAND U504 ( .A(n373), .B(n375), .Z(n1628) );
  NAND U505 ( .A(sreg[129]), .B(n777), .Z(n376) );
  XOR U506 ( .A(n777), .B(sreg[129]), .Z(n377) );
  NANDN U507 ( .A(n778), .B(n377), .Z(n378) );
  NAND U508 ( .A(n376), .B(n378), .Z(n784) );
  NAND U509 ( .A(sreg[132]), .B(n799), .Z(n379) );
  XOR U510 ( .A(n799), .B(sreg[132]), .Z(n380) );
  NAND U511 ( .A(n380), .B(n798), .Z(n381) );
  NAND U512 ( .A(n379), .B(n381), .Z(n805) );
  NAND U513 ( .A(sreg[135]), .B(n819), .Z(n382) );
  XOR U514 ( .A(n819), .B(sreg[135]), .Z(n383) );
  NANDN U515 ( .A(n820), .B(n383), .Z(n384) );
  NAND U516 ( .A(n382), .B(n384), .Z(n826) );
  NAND U517 ( .A(sreg[138]), .B(n841), .Z(n385) );
  XOR U518 ( .A(n841), .B(sreg[138]), .Z(n386) );
  NAND U519 ( .A(n386), .B(n840), .Z(n387) );
  NAND U520 ( .A(n385), .B(n387), .Z(n847) );
  NAND U521 ( .A(sreg[141]), .B(n862), .Z(n388) );
  XOR U522 ( .A(n862), .B(sreg[141]), .Z(n389) );
  NAND U523 ( .A(n389), .B(n861), .Z(n390) );
  NAND U524 ( .A(n388), .B(n390), .Z(n868) );
  NAND U525 ( .A(sreg[144]), .B(n883), .Z(n391) );
  XOR U526 ( .A(n883), .B(sreg[144]), .Z(n392) );
  NAND U527 ( .A(n392), .B(n882), .Z(n393) );
  NAND U528 ( .A(n391), .B(n393), .Z(n889) );
  NAND U529 ( .A(sreg[147]), .B(n903), .Z(n394) );
  XOR U530 ( .A(n903), .B(sreg[147]), .Z(n395) );
  NANDN U531 ( .A(n904), .B(n395), .Z(n396) );
  NAND U532 ( .A(n394), .B(n396), .Z(n910) );
  NAND U533 ( .A(sreg[150]), .B(n925), .Z(n397) );
  XOR U534 ( .A(n925), .B(sreg[150]), .Z(n398) );
  NAND U535 ( .A(n398), .B(n924), .Z(n399) );
  NAND U536 ( .A(n397), .B(n399), .Z(n931) );
  NAND U537 ( .A(sreg[153]), .B(n946), .Z(n400) );
  XOR U538 ( .A(n946), .B(sreg[153]), .Z(n401) );
  NAND U539 ( .A(n401), .B(n945), .Z(n402) );
  NAND U540 ( .A(n400), .B(n402), .Z(n952) );
  NAND U541 ( .A(sreg[156]), .B(n967), .Z(n403) );
  XOR U542 ( .A(n967), .B(sreg[156]), .Z(n404) );
  NAND U543 ( .A(n404), .B(n966), .Z(n405) );
  NAND U544 ( .A(n403), .B(n405), .Z(n973) );
  NAND U545 ( .A(sreg[159]), .B(n988), .Z(n406) );
  XOR U546 ( .A(n988), .B(sreg[159]), .Z(n407) );
  NAND U547 ( .A(n407), .B(n987), .Z(n408) );
  NAND U548 ( .A(n406), .B(n408), .Z(n994) );
  NAND U549 ( .A(sreg[162]), .B(n1009), .Z(n409) );
  XOR U550 ( .A(n1009), .B(sreg[162]), .Z(n410) );
  NAND U551 ( .A(n410), .B(n1008), .Z(n411) );
  NAND U552 ( .A(n409), .B(n411), .Z(n1015) );
  NAND U553 ( .A(sreg[165]), .B(n1030), .Z(n412) );
  XOR U554 ( .A(n1030), .B(sreg[165]), .Z(n413) );
  NAND U555 ( .A(n413), .B(n1029), .Z(n414) );
  NAND U556 ( .A(n412), .B(n414), .Z(n1036) );
  NAND U557 ( .A(sreg[168]), .B(n1051), .Z(n415) );
  XOR U558 ( .A(n1051), .B(sreg[168]), .Z(n416) );
  NAND U559 ( .A(n416), .B(n1050), .Z(n417) );
  NAND U560 ( .A(n415), .B(n417), .Z(n1057) );
  NAND U561 ( .A(sreg[171]), .B(n1072), .Z(n418) );
  XOR U562 ( .A(n1072), .B(sreg[171]), .Z(n419) );
  NAND U563 ( .A(n419), .B(n1071), .Z(n420) );
  NAND U564 ( .A(n418), .B(n420), .Z(n1078) );
  NAND U565 ( .A(sreg[174]), .B(n1093), .Z(n421) );
  XOR U566 ( .A(n1093), .B(sreg[174]), .Z(n422) );
  NAND U567 ( .A(n422), .B(n1092), .Z(n423) );
  NAND U568 ( .A(n421), .B(n423), .Z(n1099) );
  NAND U569 ( .A(sreg[177]), .B(n1114), .Z(n424) );
  XOR U570 ( .A(n1114), .B(sreg[177]), .Z(n425) );
  NAND U571 ( .A(n425), .B(n1113), .Z(n426) );
  NAND U572 ( .A(n424), .B(n426), .Z(n1120) );
  NAND U573 ( .A(sreg[180]), .B(n1135), .Z(n427) );
  XOR U574 ( .A(n1135), .B(sreg[180]), .Z(n428) );
  NAND U575 ( .A(n428), .B(n1134), .Z(n429) );
  NAND U576 ( .A(n427), .B(n429), .Z(n1141) );
  NAND U577 ( .A(sreg[183]), .B(n1156), .Z(n430) );
  XOR U578 ( .A(n1156), .B(sreg[183]), .Z(n431) );
  NAND U579 ( .A(n431), .B(n1155), .Z(n432) );
  NAND U580 ( .A(n430), .B(n432), .Z(n1162) );
  NAND U581 ( .A(sreg[186]), .B(n1177), .Z(n433) );
  XOR U582 ( .A(n1177), .B(sreg[186]), .Z(n434) );
  NAND U583 ( .A(n434), .B(n1176), .Z(n435) );
  NAND U584 ( .A(n433), .B(n435), .Z(n1183) );
  NAND U585 ( .A(sreg[189]), .B(n1198), .Z(n436) );
  XOR U586 ( .A(n1198), .B(sreg[189]), .Z(n437) );
  NAND U587 ( .A(n437), .B(n1197), .Z(n438) );
  NAND U588 ( .A(n436), .B(n438), .Z(n1204) );
  NAND U589 ( .A(sreg[192]), .B(n1219), .Z(n439) );
  XOR U590 ( .A(n1219), .B(sreg[192]), .Z(n440) );
  NAND U591 ( .A(n440), .B(n1218), .Z(n441) );
  NAND U592 ( .A(n439), .B(n441), .Z(n1225) );
  NAND U593 ( .A(sreg[195]), .B(n1240), .Z(n442) );
  XOR U594 ( .A(n1240), .B(sreg[195]), .Z(n443) );
  NAND U595 ( .A(n443), .B(n1239), .Z(n444) );
  NAND U596 ( .A(n442), .B(n444), .Z(n1246) );
  NAND U597 ( .A(sreg[198]), .B(n1261), .Z(n445) );
  XOR U598 ( .A(n1261), .B(sreg[198]), .Z(n446) );
  NAND U599 ( .A(n446), .B(n1260), .Z(n447) );
  NAND U600 ( .A(n445), .B(n447), .Z(n1267) );
  NAND U601 ( .A(sreg[201]), .B(n1282), .Z(n448) );
  XOR U602 ( .A(n1282), .B(sreg[201]), .Z(n449) );
  NAND U603 ( .A(n449), .B(n1281), .Z(n450) );
  NAND U604 ( .A(n448), .B(n450), .Z(n1288) );
  NAND U605 ( .A(sreg[204]), .B(n1303), .Z(n451) );
  XOR U606 ( .A(n1303), .B(sreg[204]), .Z(n452) );
  NAND U607 ( .A(n452), .B(n1302), .Z(n453) );
  NAND U608 ( .A(n451), .B(n453), .Z(n1309) );
  NAND U609 ( .A(sreg[207]), .B(n1324), .Z(n454) );
  XOR U610 ( .A(n1324), .B(sreg[207]), .Z(n455) );
  NAND U611 ( .A(n455), .B(n1323), .Z(n456) );
  NAND U612 ( .A(n454), .B(n456), .Z(n1330) );
  NAND U613 ( .A(sreg[210]), .B(n1345), .Z(n457) );
  XOR U614 ( .A(n1345), .B(sreg[210]), .Z(n458) );
  NAND U615 ( .A(n458), .B(n1344), .Z(n459) );
  NAND U616 ( .A(n457), .B(n459), .Z(n1351) );
  NAND U617 ( .A(sreg[213]), .B(n1366), .Z(n460) );
  XOR U618 ( .A(n1366), .B(sreg[213]), .Z(n461) );
  NAND U619 ( .A(n461), .B(n1365), .Z(n462) );
  NAND U620 ( .A(n460), .B(n462), .Z(n1372) );
  NAND U621 ( .A(sreg[216]), .B(n1387), .Z(n463) );
  XOR U622 ( .A(n1387), .B(sreg[216]), .Z(n464) );
  NAND U623 ( .A(n464), .B(n1386), .Z(n465) );
  NAND U624 ( .A(n463), .B(n465), .Z(n1393) );
  NAND U625 ( .A(sreg[219]), .B(n1408), .Z(n466) );
  XOR U626 ( .A(n1408), .B(sreg[219]), .Z(n467) );
  NAND U627 ( .A(n467), .B(n1407), .Z(n468) );
  NAND U628 ( .A(n466), .B(n468), .Z(n1414) );
  NAND U629 ( .A(sreg[222]), .B(n1429), .Z(n469) );
  XOR U630 ( .A(n1429), .B(sreg[222]), .Z(n470) );
  NAND U631 ( .A(n470), .B(n1428), .Z(n471) );
  NAND U632 ( .A(n469), .B(n471), .Z(n1435) );
  NAND U633 ( .A(sreg[225]), .B(n1450), .Z(n472) );
  XOR U634 ( .A(n1450), .B(sreg[225]), .Z(n473) );
  NAND U635 ( .A(n473), .B(n1449), .Z(n474) );
  NAND U636 ( .A(n472), .B(n474), .Z(n1456) );
  NAND U637 ( .A(sreg[228]), .B(n1471), .Z(n475) );
  XOR U638 ( .A(n1471), .B(sreg[228]), .Z(n476) );
  NAND U639 ( .A(n476), .B(n1470), .Z(n477) );
  NAND U640 ( .A(n475), .B(n477), .Z(n1477) );
  NAND U641 ( .A(sreg[231]), .B(n1492), .Z(n478) );
  XOR U642 ( .A(n1492), .B(sreg[231]), .Z(n479) );
  NAND U643 ( .A(n479), .B(n1491), .Z(n480) );
  NAND U644 ( .A(n478), .B(n480), .Z(n1498) );
  NAND U645 ( .A(sreg[234]), .B(n1513), .Z(n481) );
  XOR U646 ( .A(n1513), .B(sreg[234]), .Z(n482) );
  NAND U647 ( .A(n482), .B(n1512), .Z(n483) );
  NAND U648 ( .A(n481), .B(n483), .Z(n1519) );
  NAND U649 ( .A(sreg[237]), .B(n1534), .Z(n484) );
  XOR U650 ( .A(n1534), .B(sreg[237]), .Z(n485) );
  NAND U651 ( .A(n485), .B(n1533), .Z(n486) );
  NAND U652 ( .A(n484), .B(n486), .Z(n1540) );
  NAND U653 ( .A(sreg[240]), .B(n1555), .Z(n487) );
  XOR U654 ( .A(n1555), .B(sreg[240]), .Z(n488) );
  NAND U655 ( .A(n488), .B(n1554), .Z(n489) );
  NAND U656 ( .A(n487), .B(n489), .Z(n1561) );
  NAND U657 ( .A(sreg[243]), .B(n1576), .Z(n490) );
  XOR U658 ( .A(n1576), .B(sreg[243]), .Z(n491) );
  NAND U659 ( .A(n491), .B(n1575), .Z(n492) );
  NAND U660 ( .A(n490), .B(n492), .Z(n1582) );
  NAND U661 ( .A(sreg[246]), .B(n1597), .Z(n493) );
  XOR U662 ( .A(n1597), .B(sreg[246]), .Z(n494) );
  NAND U663 ( .A(n494), .B(n1596), .Z(n495) );
  NAND U664 ( .A(n493), .B(n495), .Z(n1603) );
  NAND U665 ( .A(sreg[249]), .B(n1618), .Z(n496) );
  XOR U666 ( .A(n1618), .B(sreg[249]), .Z(n497) );
  NAND U667 ( .A(n497), .B(n1617), .Z(n498) );
  NAND U668 ( .A(n496), .B(n498), .Z(n1624) );
  NAND U669 ( .A(sreg[252]), .B(n1638), .Z(n499) );
  XOR U670 ( .A(n1638), .B(sreg[252]), .Z(n500) );
  NANDN U671 ( .A(n1639), .B(n500), .Z(n501) );
  NAND U672 ( .A(n499), .B(n501), .Z(n1641) );
  NAND U673 ( .A(n789), .B(n787), .Z(n502) );
  XOR U674 ( .A(n787), .B(n789), .Z(n503) );
  NAND U675 ( .A(n503), .B(n788), .Z(n504) );
  NAND U676 ( .A(n502), .B(n504), .Z(n795) );
  NAND U677 ( .A(n810), .B(n809), .Z(n505) );
  XOR U678 ( .A(n809), .B(n810), .Z(n506) );
  NAND U679 ( .A(n506), .B(n808), .Z(n507) );
  NAND U680 ( .A(n505), .B(n507), .Z(n816) );
  NAND U681 ( .A(n831), .B(n830), .Z(n508) );
  XOR U682 ( .A(n830), .B(n831), .Z(n509) );
  NAND U683 ( .A(n509), .B(n829), .Z(n510) );
  NAND U684 ( .A(n508), .B(n510), .Z(n837) );
  NAND U685 ( .A(n852), .B(n851), .Z(n511) );
  XOR U686 ( .A(n851), .B(n852), .Z(n512) );
  NAND U687 ( .A(n512), .B(n850), .Z(n513) );
  NAND U688 ( .A(n511), .B(n513), .Z(n858) );
  NAND U689 ( .A(n873), .B(n871), .Z(n514) );
  XOR U690 ( .A(n871), .B(n873), .Z(n515) );
  NAND U691 ( .A(n515), .B(n872), .Z(n516) );
  NAND U692 ( .A(n514), .B(n516), .Z(n879) );
  NAND U693 ( .A(n894), .B(n893), .Z(n517) );
  XOR U694 ( .A(n893), .B(n894), .Z(n518) );
  NAND U695 ( .A(n518), .B(n892), .Z(n519) );
  NAND U696 ( .A(n517), .B(n519), .Z(n900) );
  NAND U697 ( .A(n915), .B(n914), .Z(n520) );
  XOR U698 ( .A(n914), .B(n915), .Z(n521) );
  NAND U699 ( .A(n521), .B(n913), .Z(n522) );
  NAND U700 ( .A(n520), .B(n522), .Z(n921) );
  NAND U701 ( .A(n936), .B(n935), .Z(n523) );
  XOR U702 ( .A(n935), .B(n936), .Z(n524) );
  NAND U703 ( .A(n524), .B(n934), .Z(n525) );
  NAND U704 ( .A(n523), .B(n525), .Z(n942) );
  NAND U705 ( .A(n957), .B(n956), .Z(n526) );
  XOR U706 ( .A(n956), .B(n957), .Z(n527) );
  NAND U707 ( .A(n527), .B(n955), .Z(n528) );
  NAND U708 ( .A(n526), .B(n528), .Z(n963) );
  NAND U709 ( .A(n978), .B(n977), .Z(n529) );
  XOR U710 ( .A(n977), .B(n978), .Z(n530) );
  NAND U711 ( .A(n530), .B(n976), .Z(n531) );
  NAND U712 ( .A(n529), .B(n531), .Z(n984) );
  NAND U713 ( .A(n999), .B(n998), .Z(n532) );
  XOR U714 ( .A(n998), .B(n999), .Z(n533) );
  NAND U715 ( .A(n533), .B(n997), .Z(n534) );
  NAND U716 ( .A(n532), .B(n534), .Z(n1005) );
  NAND U717 ( .A(n1020), .B(n1019), .Z(n535) );
  XOR U718 ( .A(n1019), .B(n1020), .Z(n536) );
  NAND U719 ( .A(n536), .B(n1018), .Z(n537) );
  NAND U720 ( .A(n535), .B(n537), .Z(n1026) );
  NAND U721 ( .A(n1041), .B(n1040), .Z(n538) );
  XOR U722 ( .A(n1040), .B(n1041), .Z(n539) );
  NAND U723 ( .A(n539), .B(n1039), .Z(n540) );
  NAND U724 ( .A(n538), .B(n540), .Z(n1047) );
  NAND U725 ( .A(n1062), .B(n1061), .Z(n541) );
  XOR U726 ( .A(n1061), .B(n1062), .Z(n542) );
  NAND U727 ( .A(n542), .B(n1060), .Z(n543) );
  NAND U728 ( .A(n541), .B(n543), .Z(n1068) );
  NAND U729 ( .A(n1083), .B(n1082), .Z(n544) );
  XOR U730 ( .A(n1082), .B(n1083), .Z(n545) );
  NAND U731 ( .A(n545), .B(n1081), .Z(n546) );
  NAND U732 ( .A(n544), .B(n546), .Z(n1089) );
  NAND U733 ( .A(n1104), .B(n1103), .Z(n547) );
  XOR U734 ( .A(n1103), .B(n1104), .Z(n548) );
  NAND U735 ( .A(n548), .B(n1102), .Z(n549) );
  NAND U736 ( .A(n547), .B(n549), .Z(n1110) );
  NAND U737 ( .A(n1125), .B(n1124), .Z(n550) );
  XOR U738 ( .A(n1124), .B(n1125), .Z(n551) );
  NAND U739 ( .A(n551), .B(n1123), .Z(n552) );
  NAND U740 ( .A(n550), .B(n552), .Z(n1131) );
  NAND U741 ( .A(n1146), .B(n1145), .Z(n553) );
  XOR U742 ( .A(n1145), .B(n1146), .Z(n554) );
  NAND U743 ( .A(n554), .B(n1144), .Z(n555) );
  NAND U744 ( .A(n553), .B(n555), .Z(n1152) );
  NAND U745 ( .A(n1167), .B(n1166), .Z(n556) );
  XOR U746 ( .A(n1166), .B(n1167), .Z(n557) );
  NAND U747 ( .A(n557), .B(n1165), .Z(n558) );
  NAND U748 ( .A(n556), .B(n558), .Z(n1173) );
  NAND U749 ( .A(n1188), .B(n1187), .Z(n559) );
  XOR U750 ( .A(n1187), .B(n1188), .Z(n560) );
  NAND U751 ( .A(n560), .B(n1186), .Z(n561) );
  NAND U752 ( .A(n559), .B(n561), .Z(n1194) );
  NAND U753 ( .A(n1209), .B(n1208), .Z(n562) );
  XOR U754 ( .A(n1208), .B(n1209), .Z(n563) );
  NAND U755 ( .A(n563), .B(n1207), .Z(n564) );
  NAND U756 ( .A(n562), .B(n564), .Z(n1215) );
  NAND U757 ( .A(n1230), .B(n1229), .Z(n565) );
  XOR U758 ( .A(n1229), .B(n1230), .Z(n566) );
  NAND U759 ( .A(n566), .B(n1228), .Z(n567) );
  NAND U760 ( .A(n565), .B(n567), .Z(n1236) );
  NAND U761 ( .A(n1251), .B(n1250), .Z(n568) );
  XOR U762 ( .A(n1250), .B(n1251), .Z(n569) );
  NAND U763 ( .A(n569), .B(n1249), .Z(n570) );
  NAND U764 ( .A(n568), .B(n570), .Z(n1257) );
  NAND U765 ( .A(n1272), .B(n1271), .Z(n571) );
  XOR U766 ( .A(n1271), .B(n1272), .Z(n572) );
  NAND U767 ( .A(n572), .B(n1270), .Z(n573) );
  NAND U768 ( .A(n571), .B(n573), .Z(n1278) );
  NAND U769 ( .A(n1293), .B(n1292), .Z(n574) );
  XOR U770 ( .A(n1292), .B(n1293), .Z(n575) );
  NAND U771 ( .A(n575), .B(n1291), .Z(n576) );
  NAND U772 ( .A(n574), .B(n576), .Z(n1299) );
  NAND U773 ( .A(n1314), .B(n1313), .Z(n577) );
  XOR U774 ( .A(n1313), .B(n1314), .Z(n578) );
  NAND U775 ( .A(n578), .B(n1312), .Z(n579) );
  NAND U776 ( .A(n577), .B(n579), .Z(n1320) );
  NAND U777 ( .A(n1335), .B(n1334), .Z(n580) );
  XOR U778 ( .A(n1334), .B(n1335), .Z(n581) );
  NAND U779 ( .A(n581), .B(n1333), .Z(n582) );
  NAND U780 ( .A(n580), .B(n582), .Z(n1341) );
  NAND U781 ( .A(n1356), .B(n1355), .Z(n583) );
  XOR U782 ( .A(n1355), .B(n1356), .Z(n584) );
  NAND U783 ( .A(n584), .B(n1354), .Z(n585) );
  NAND U784 ( .A(n583), .B(n585), .Z(n1362) );
  NAND U785 ( .A(n1377), .B(n1376), .Z(n586) );
  XOR U786 ( .A(n1376), .B(n1377), .Z(n587) );
  NAND U787 ( .A(n587), .B(n1375), .Z(n588) );
  NAND U788 ( .A(n586), .B(n588), .Z(n1383) );
  NAND U789 ( .A(n1398), .B(n1397), .Z(n589) );
  XOR U790 ( .A(n1397), .B(n1398), .Z(n590) );
  NAND U791 ( .A(n590), .B(n1396), .Z(n591) );
  NAND U792 ( .A(n589), .B(n591), .Z(n1404) );
  NAND U793 ( .A(n1419), .B(n1418), .Z(n592) );
  XOR U794 ( .A(n1418), .B(n1419), .Z(n593) );
  NAND U795 ( .A(n593), .B(n1417), .Z(n594) );
  NAND U796 ( .A(n592), .B(n594), .Z(n1425) );
  NAND U797 ( .A(n1440), .B(n1439), .Z(n595) );
  XOR U798 ( .A(n1439), .B(n1440), .Z(n596) );
  NAND U799 ( .A(n596), .B(n1438), .Z(n597) );
  NAND U800 ( .A(n595), .B(n597), .Z(n1446) );
  NAND U801 ( .A(n1461), .B(n1460), .Z(n598) );
  XOR U802 ( .A(n1460), .B(n1461), .Z(n599) );
  NAND U803 ( .A(n599), .B(n1459), .Z(n600) );
  NAND U804 ( .A(n598), .B(n600), .Z(n1467) );
  NAND U805 ( .A(n1482), .B(n1481), .Z(n601) );
  XOR U806 ( .A(n1481), .B(n1482), .Z(n602) );
  NAND U807 ( .A(n602), .B(n1480), .Z(n603) );
  NAND U808 ( .A(n601), .B(n603), .Z(n1488) );
  NAND U809 ( .A(n1503), .B(n1502), .Z(n604) );
  XOR U810 ( .A(n1502), .B(n1503), .Z(n605) );
  NAND U811 ( .A(n605), .B(n1501), .Z(n606) );
  NAND U812 ( .A(n604), .B(n606), .Z(n1509) );
  NAND U813 ( .A(n1524), .B(n1523), .Z(n607) );
  XOR U814 ( .A(n1523), .B(n1524), .Z(n608) );
  NAND U815 ( .A(n608), .B(n1522), .Z(n609) );
  NAND U816 ( .A(n607), .B(n609), .Z(n1530) );
  NAND U817 ( .A(n1545), .B(n1544), .Z(n610) );
  XOR U818 ( .A(n1544), .B(n1545), .Z(n611) );
  NAND U819 ( .A(n611), .B(n1543), .Z(n612) );
  NAND U820 ( .A(n610), .B(n612), .Z(n1551) );
  NAND U821 ( .A(n1566), .B(n1565), .Z(n613) );
  XOR U822 ( .A(n1565), .B(n1566), .Z(n614) );
  NAND U823 ( .A(n614), .B(n1564), .Z(n615) );
  NAND U824 ( .A(n613), .B(n615), .Z(n1572) );
  NAND U825 ( .A(n1587), .B(n1586), .Z(n616) );
  XOR U826 ( .A(n1586), .B(n1587), .Z(n617) );
  NAND U827 ( .A(n617), .B(n1585), .Z(n618) );
  NAND U828 ( .A(n616), .B(n618), .Z(n1593) );
  NAND U829 ( .A(n1608), .B(n1607), .Z(n619) );
  XOR U830 ( .A(n1607), .B(n1608), .Z(n620) );
  NAND U831 ( .A(n620), .B(n1606), .Z(n621) );
  NAND U832 ( .A(n619), .B(n621), .Z(n1614) );
  NAND U833 ( .A(sreg[130]), .B(n785), .Z(n622) );
  XOR U834 ( .A(n785), .B(sreg[130]), .Z(n623) );
  NAND U835 ( .A(n623), .B(n784), .Z(n624) );
  NAND U836 ( .A(n622), .B(n624), .Z(n791) );
  NAND U837 ( .A(sreg[133]), .B(n806), .Z(n625) );
  XOR U838 ( .A(n806), .B(sreg[133]), .Z(n626) );
  NAND U839 ( .A(n626), .B(n805), .Z(n627) );
  NAND U840 ( .A(n625), .B(n627), .Z(n812) );
  NAND U841 ( .A(sreg[136]), .B(n827), .Z(n628) );
  XOR U842 ( .A(n827), .B(sreg[136]), .Z(n629) );
  NAND U843 ( .A(n629), .B(n826), .Z(n630) );
  NAND U844 ( .A(n628), .B(n630), .Z(n833) );
  NAND U845 ( .A(sreg[139]), .B(n847), .Z(n631) );
  XOR U846 ( .A(n847), .B(sreg[139]), .Z(n632) );
  NANDN U847 ( .A(n848), .B(n632), .Z(n633) );
  NAND U848 ( .A(n631), .B(n633), .Z(n854) );
  NAND U849 ( .A(sreg[142]), .B(n869), .Z(n634) );
  XOR U850 ( .A(n869), .B(sreg[142]), .Z(n635) );
  NAND U851 ( .A(n635), .B(n868), .Z(n636) );
  NAND U852 ( .A(n634), .B(n636), .Z(n875) );
  NAND U853 ( .A(sreg[145]), .B(n890), .Z(n637) );
  XOR U854 ( .A(n890), .B(sreg[145]), .Z(n638) );
  NAND U855 ( .A(n638), .B(n889), .Z(n639) );
  NAND U856 ( .A(n637), .B(n639), .Z(n896) );
  NAND U857 ( .A(sreg[148]), .B(n911), .Z(n640) );
  XOR U858 ( .A(n911), .B(sreg[148]), .Z(n641) );
  NAND U859 ( .A(n641), .B(n910), .Z(n642) );
  NAND U860 ( .A(n640), .B(n642), .Z(n917) );
  NAND U861 ( .A(sreg[151]), .B(n932), .Z(n643) );
  XOR U862 ( .A(n932), .B(sreg[151]), .Z(n644) );
  NAND U863 ( .A(n644), .B(n931), .Z(n645) );
  NAND U864 ( .A(n643), .B(n645), .Z(n938) );
  NAND U865 ( .A(sreg[154]), .B(n953), .Z(n646) );
  XOR U866 ( .A(n953), .B(sreg[154]), .Z(n647) );
  NAND U867 ( .A(n647), .B(n952), .Z(n648) );
  NAND U868 ( .A(n646), .B(n648), .Z(n959) );
  NAND U869 ( .A(sreg[157]), .B(n974), .Z(n649) );
  XOR U870 ( .A(n974), .B(sreg[157]), .Z(n650) );
  NAND U871 ( .A(n650), .B(n973), .Z(n651) );
  NAND U872 ( .A(n649), .B(n651), .Z(n980) );
  NAND U873 ( .A(sreg[160]), .B(n995), .Z(n652) );
  XOR U874 ( .A(n995), .B(sreg[160]), .Z(n653) );
  NAND U875 ( .A(n653), .B(n994), .Z(n654) );
  NAND U876 ( .A(n652), .B(n654), .Z(n1001) );
  NAND U877 ( .A(sreg[163]), .B(n1016), .Z(n655) );
  XOR U878 ( .A(n1016), .B(sreg[163]), .Z(n656) );
  NAND U879 ( .A(n656), .B(n1015), .Z(n657) );
  NAND U880 ( .A(n655), .B(n657), .Z(n1022) );
  NAND U881 ( .A(sreg[166]), .B(n1037), .Z(n658) );
  XOR U882 ( .A(n1037), .B(sreg[166]), .Z(n659) );
  NAND U883 ( .A(n659), .B(n1036), .Z(n660) );
  NAND U884 ( .A(n658), .B(n660), .Z(n1043) );
  NAND U885 ( .A(sreg[169]), .B(n1058), .Z(n661) );
  XOR U886 ( .A(n1058), .B(sreg[169]), .Z(n662) );
  NAND U887 ( .A(n662), .B(n1057), .Z(n663) );
  NAND U888 ( .A(n661), .B(n663), .Z(n1064) );
  NAND U889 ( .A(sreg[172]), .B(n1079), .Z(n664) );
  XOR U890 ( .A(n1079), .B(sreg[172]), .Z(n665) );
  NAND U891 ( .A(n665), .B(n1078), .Z(n666) );
  NAND U892 ( .A(n664), .B(n666), .Z(n1085) );
  NAND U893 ( .A(sreg[175]), .B(n1100), .Z(n667) );
  XOR U894 ( .A(n1100), .B(sreg[175]), .Z(n668) );
  NAND U895 ( .A(n668), .B(n1099), .Z(n669) );
  NAND U896 ( .A(n667), .B(n669), .Z(n1106) );
  NAND U897 ( .A(sreg[178]), .B(n1121), .Z(n670) );
  XOR U898 ( .A(n1121), .B(sreg[178]), .Z(n671) );
  NAND U899 ( .A(n671), .B(n1120), .Z(n672) );
  NAND U900 ( .A(n670), .B(n672), .Z(n1127) );
  NAND U901 ( .A(sreg[181]), .B(n1142), .Z(n673) );
  XOR U902 ( .A(n1142), .B(sreg[181]), .Z(n674) );
  NAND U903 ( .A(n674), .B(n1141), .Z(n675) );
  NAND U904 ( .A(n673), .B(n675), .Z(n1148) );
  NAND U905 ( .A(sreg[184]), .B(n1163), .Z(n676) );
  XOR U906 ( .A(n1163), .B(sreg[184]), .Z(n677) );
  NAND U907 ( .A(n677), .B(n1162), .Z(n678) );
  NAND U908 ( .A(n676), .B(n678), .Z(n1169) );
  NAND U909 ( .A(sreg[187]), .B(n1184), .Z(n679) );
  XOR U910 ( .A(n1184), .B(sreg[187]), .Z(n680) );
  NAND U911 ( .A(n680), .B(n1183), .Z(n681) );
  NAND U912 ( .A(n679), .B(n681), .Z(n1190) );
  NAND U913 ( .A(sreg[190]), .B(n1205), .Z(n682) );
  XOR U914 ( .A(n1205), .B(sreg[190]), .Z(n683) );
  NAND U915 ( .A(n683), .B(n1204), .Z(n684) );
  NAND U916 ( .A(n682), .B(n684), .Z(n1211) );
  NAND U917 ( .A(sreg[193]), .B(n1226), .Z(n685) );
  XOR U918 ( .A(n1226), .B(sreg[193]), .Z(n686) );
  NAND U919 ( .A(n686), .B(n1225), .Z(n687) );
  NAND U920 ( .A(n685), .B(n687), .Z(n1232) );
  NAND U921 ( .A(sreg[196]), .B(n1247), .Z(n688) );
  XOR U922 ( .A(n1247), .B(sreg[196]), .Z(n689) );
  NAND U923 ( .A(n689), .B(n1246), .Z(n690) );
  NAND U924 ( .A(n688), .B(n690), .Z(n1253) );
  NAND U925 ( .A(sreg[199]), .B(n1268), .Z(n691) );
  XOR U926 ( .A(n1268), .B(sreg[199]), .Z(n692) );
  NAND U927 ( .A(n692), .B(n1267), .Z(n693) );
  NAND U928 ( .A(n691), .B(n693), .Z(n1274) );
  NAND U929 ( .A(sreg[202]), .B(n1289), .Z(n694) );
  XOR U930 ( .A(n1289), .B(sreg[202]), .Z(n695) );
  NAND U931 ( .A(n695), .B(n1288), .Z(n696) );
  NAND U932 ( .A(n694), .B(n696), .Z(n1295) );
  NAND U933 ( .A(sreg[205]), .B(n1310), .Z(n697) );
  XOR U934 ( .A(n1310), .B(sreg[205]), .Z(n698) );
  NAND U935 ( .A(n698), .B(n1309), .Z(n699) );
  NAND U936 ( .A(n697), .B(n699), .Z(n1316) );
  NAND U937 ( .A(sreg[208]), .B(n1331), .Z(n700) );
  XOR U938 ( .A(n1331), .B(sreg[208]), .Z(n701) );
  NAND U939 ( .A(n701), .B(n1330), .Z(n702) );
  NAND U940 ( .A(n700), .B(n702), .Z(n1337) );
  NAND U941 ( .A(sreg[211]), .B(n1352), .Z(n703) );
  XOR U942 ( .A(n1352), .B(sreg[211]), .Z(n704) );
  NAND U943 ( .A(n704), .B(n1351), .Z(n705) );
  NAND U944 ( .A(n703), .B(n705), .Z(n1358) );
  NAND U945 ( .A(sreg[214]), .B(n1373), .Z(n706) );
  XOR U946 ( .A(n1373), .B(sreg[214]), .Z(n707) );
  NAND U947 ( .A(n707), .B(n1372), .Z(n708) );
  NAND U948 ( .A(n706), .B(n708), .Z(n1379) );
  NAND U949 ( .A(sreg[217]), .B(n1394), .Z(n709) );
  XOR U950 ( .A(n1394), .B(sreg[217]), .Z(n710) );
  NAND U951 ( .A(n710), .B(n1393), .Z(n711) );
  NAND U952 ( .A(n709), .B(n711), .Z(n1400) );
  NAND U953 ( .A(sreg[220]), .B(n1415), .Z(n712) );
  XOR U954 ( .A(n1415), .B(sreg[220]), .Z(n713) );
  NAND U955 ( .A(n713), .B(n1414), .Z(n714) );
  NAND U956 ( .A(n712), .B(n714), .Z(n1421) );
  NAND U957 ( .A(sreg[223]), .B(n1436), .Z(n715) );
  XOR U958 ( .A(n1436), .B(sreg[223]), .Z(n716) );
  NAND U959 ( .A(n716), .B(n1435), .Z(n717) );
  NAND U960 ( .A(n715), .B(n717), .Z(n1442) );
  NAND U961 ( .A(sreg[226]), .B(n1457), .Z(n718) );
  XOR U962 ( .A(n1457), .B(sreg[226]), .Z(n719) );
  NAND U963 ( .A(n719), .B(n1456), .Z(n720) );
  NAND U964 ( .A(n718), .B(n720), .Z(n1463) );
  NAND U965 ( .A(sreg[229]), .B(n1478), .Z(n721) );
  XOR U966 ( .A(n1478), .B(sreg[229]), .Z(n722) );
  NAND U967 ( .A(n722), .B(n1477), .Z(n723) );
  NAND U968 ( .A(n721), .B(n723), .Z(n1484) );
  NAND U969 ( .A(sreg[232]), .B(n1499), .Z(n724) );
  XOR U970 ( .A(n1499), .B(sreg[232]), .Z(n725) );
  NAND U971 ( .A(n725), .B(n1498), .Z(n726) );
  NAND U972 ( .A(n724), .B(n726), .Z(n1505) );
  NAND U973 ( .A(sreg[235]), .B(n1520), .Z(n727) );
  XOR U974 ( .A(n1520), .B(sreg[235]), .Z(n728) );
  NAND U975 ( .A(n728), .B(n1519), .Z(n729) );
  NAND U976 ( .A(n727), .B(n729), .Z(n1526) );
  NAND U977 ( .A(sreg[238]), .B(n1541), .Z(n730) );
  XOR U978 ( .A(n1541), .B(sreg[238]), .Z(n731) );
  NAND U979 ( .A(n731), .B(n1540), .Z(n732) );
  NAND U980 ( .A(n730), .B(n732), .Z(n1547) );
  NAND U981 ( .A(sreg[241]), .B(n1562), .Z(n733) );
  XOR U982 ( .A(n1562), .B(sreg[241]), .Z(n734) );
  NAND U983 ( .A(n734), .B(n1561), .Z(n735) );
  NAND U984 ( .A(n733), .B(n735), .Z(n1568) );
  NAND U985 ( .A(sreg[244]), .B(n1583), .Z(n736) );
  XOR U986 ( .A(n1583), .B(sreg[244]), .Z(n737) );
  NAND U987 ( .A(n737), .B(n1582), .Z(n738) );
  NAND U988 ( .A(n736), .B(n738), .Z(n1589) );
  NAND U989 ( .A(sreg[247]), .B(n1604), .Z(n739) );
  XOR U990 ( .A(n1604), .B(sreg[247]), .Z(n740) );
  NAND U991 ( .A(n740), .B(n1603), .Z(n741) );
  NAND U992 ( .A(n739), .B(n741), .Z(n1610) );
  NAND U993 ( .A(sreg[250]), .B(n1625), .Z(n742) );
  XOR U994 ( .A(n1625), .B(sreg[250]), .Z(n743) );
  NAND U995 ( .A(n743), .B(n1624), .Z(n744) );
  NAND U996 ( .A(n742), .B(n744), .Z(n1631) );
  NAND U997 ( .A(sreg[253]), .B(n1642), .Z(n745) );
  XOR U998 ( .A(n1642), .B(sreg[253]), .Z(n746) );
  NAND U999 ( .A(n746), .B(n1641), .Z(n747) );
  NAND U1000 ( .A(n745), .B(n747), .Z(n1652) );
  IV U1001 ( .A(b[1]), .Z(n748) );
  IV U1002 ( .A(b[0]), .Z(n1634) );
  NANDN U1003 ( .A(n1634), .B(a[0]), .Z(n749) );
  XNOR U1004 ( .A(n749), .B(sreg[126]), .Z(c[126]) );
  ANDN U1005 ( .B(a[0]), .A(n748), .Z(n760) );
  ANDN U1006 ( .B(a[1]), .A(n1634), .Z(n773) );
  XNOR U1007 ( .A(n760), .B(n773), .Z(n753) );
  XOR U1008 ( .A(sreg[127]), .B(n753), .Z(n755) );
  NANDN U1009 ( .A(n749), .B(sreg[126]), .Z(n754) );
  XOR U1010 ( .A(n755), .B(n754), .Z(c[127]) );
  IV U1011 ( .A(n773), .Z(n759) );
  ANDN U1012 ( .B(n760), .A(n759), .Z(n770) );
  IV U1013 ( .A(n770), .Z(n767) );
  ANDN U1014 ( .B(a[2]), .A(n1634), .Z(n751) );
  NANDN U1015 ( .A(n748), .B(a[1]), .Z(n750) );
  XNOR U1016 ( .A(n751), .B(n750), .Z(n752) );
  XOR U1017 ( .A(n767), .B(n752), .Z(n765) );
  NANDN U1018 ( .A(n753), .B(sreg[127]), .Z(n757) );
  OR U1019 ( .A(n755), .B(n754), .Z(n756) );
  NAND U1020 ( .A(n757), .B(n756), .Z(n764) );
  XOR U1021 ( .A(n764), .B(sreg[128]), .Z(n758) );
  XNOR U1022 ( .A(n765), .B(n758), .Z(c[128]) );
  NANDN U1023 ( .A(n1634), .B(a[3]), .Z(n771) );
  AND U1024 ( .A(a[2]), .B(b[1]), .Z(n769) );
  XNOR U1025 ( .A(n759), .B(n769), .Z(n762) );
  NANDN U1026 ( .A(n760), .B(n773), .Z(n761) );
  NAND U1027 ( .A(n762), .B(n761), .Z(n763) );
  XNOR U1028 ( .A(n771), .B(n763), .Z(n778) );
  XOR U1029 ( .A(n777), .B(sreg[129]), .Z(n766) );
  XNOR U1030 ( .A(n778), .B(n766), .Z(c[129]) );
  OR U1031 ( .A(n771), .B(n767), .Z(n768) );
  NANDN U1032 ( .A(n769), .B(n768), .Z(n775) );
  ANDN U1033 ( .B(n771), .A(n770), .Z(n772) );
  NANDN U1034 ( .A(n773), .B(n772), .Z(n774) );
  NAND U1035 ( .A(n775), .B(n774), .Z(n780) );
  AND U1036 ( .A(a[3]), .B(b[1]), .Z(n782) );
  ANDN U1037 ( .B(a[4]), .A(n1634), .Z(n781) );
  XNOR U1038 ( .A(n782), .B(n781), .Z(n776) );
  XOR U1039 ( .A(n780), .B(n776), .Z(n785) );
  XOR U1040 ( .A(n784), .B(sreg[130]), .Z(n779) );
  XOR U1041 ( .A(n785), .B(n779), .Z(c[130]) );
  AND U1042 ( .A(a[4]), .B(b[1]), .Z(n789) );
  ANDN U1043 ( .B(a[5]), .A(n1634), .Z(n787) );
  XOR U1044 ( .A(n788), .B(n787), .Z(n783) );
  XNOR U1045 ( .A(n789), .B(n783), .Z(n792) );
  XOR U1046 ( .A(n791), .B(sreg[131]), .Z(n786) );
  XNOR U1047 ( .A(n792), .B(n786), .Z(c[131]) );
  ANDN U1048 ( .B(a[6]), .A(n1634), .Z(n794) );
  AND U1049 ( .A(a[5]), .B(b[1]), .Z(n796) );
  XNOR U1050 ( .A(n796), .B(n795), .Z(n790) );
  XNOR U1051 ( .A(n794), .B(n790), .Z(n799) );
  XOR U1052 ( .A(n798), .B(sreg[132]), .Z(n793) );
  XOR U1053 ( .A(n799), .B(n793), .Z(c[132]) );
  ANDN U1054 ( .B(a[7]), .A(n1634), .Z(n801) );
  AND U1055 ( .A(a[6]), .B(b[1]), .Z(n803) );
  XNOR U1056 ( .A(n803), .B(n802), .Z(n797) );
  XNOR U1057 ( .A(n801), .B(n797), .Z(n806) );
  XOR U1058 ( .A(n805), .B(sreg[133]), .Z(n800) );
  XOR U1059 ( .A(n806), .B(n800), .Z(c[133]) );
  ANDN U1060 ( .B(a[8]), .A(n1634), .Z(n808) );
  AND U1061 ( .A(a[7]), .B(b[1]), .Z(n810) );
  XNOR U1062 ( .A(n810), .B(n809), .Z(n804) );
  XNOR U1063 ( .A(n808), .B(n804), .Z(n813) );
  XOR U1064 ( .A(n812), .B(sreg[134]), .Z(n807) );
  XOR U1065 ( .A(n813), .B(n807), .Z(c[134]) );
  AND U1066 ( .A(a[8]), .B(b[1]), .Z(n817) );
  ANDN U1067 ( .B(a[9]), .A(n1634), .Z(n815) );
  XOR U1068 ( .A(n816), .B(n815), .Z(n811) );
  XNOR U1069 ( .A(n817), .B(n811), .Z(n820) );
  XOR U1070 ( .A(n819), .B(sreg[135]), .Z(n814) );
  XNOR U1071 ( .A(n820), .B(n814), .Z(c[135]) );
  ANDN U1072 ( .B(a[10]), .A(n1634), .Z(n822) );
  AND U1073 ( .A(a[9]), .B(b[1]), .Z(n824) );
  XNOR U1074 ( .A(n824), .B(n823), .Z(n818) );
  XNOR U1075 ( .A(n822), .B(n818), .Z(n827) );
  XOR U1076 ( .A(n826), .B(sreg[136]), .Z(n821) );
  XOR U1077 ( .A(n827), .B(n821), .Z(c[136]) );
  ANDN U1078 ( .B(a[11]), .A(n1634), .Z(n829) );
  AND U1079 ( .A(a[10]), .B(b[1]), .Z(n831) );
  XNOR U1080 ( .A(n831), .B(n830), .Z(n825) );
  XNOR U1081 ( .A(n829), .B(n825), .Z(n834) );
  XOR U1082 ( .A(n833), .B(sreg[137]), .Z(n828) );
  XOR U1083 ( .A(n834), .B(n828), .Z(c[137]) );
  ANDN U1084 ( .B(a[12]), .A(n1634), .Z(n836) );
  AND U1085 ( .A(a[11]), .B(b[1]), .Z(n838) );
  XNOR U1086 ( .A(n838), .B(n837), .Z(n832) );
  XNOR U1087 ( .A(n836), .B(n832), .Z(n841) );
  XOR U1088 ( .A(n840), .B(sreg[138]), .Z(n835) );
  XOR U1089 ( .A(n841), .B(n835), .Z(c[138]) );
  AND U1090 ( .A(a[12]), .B(b[1]), .Z(n845) );
  ANDN U1091 ( .B(a[13]), .A(n1634), .Z(n843) );
  XOR U1092 ( .A(n844), .B(n843), .Z(n839) );
  XNOR U1093 ( .A(n845), .B(n839), .Z(n848) );
  XOR U1094 ( .A(n847), .B(sreg[139]), .Z(n842) );
  XNOR U1095 ( .A(n848), .B(n842), .Z(c[139]) );
  ANDN U1096 ( .B(a[14]), .A(n1634), .Z(n850) );
  AND U1097 ( .A(a[13]), .B(b[1]), .Z(n852) );
  XNOR U1098 ( .A(n852), .B(n851), .Z(n846) );
  XNOR U1099 ( .A(n850), .B(n846), .Z(n855) );
  XOR U1100 ( .A(n854), .B(sreg[140]), .Z(n849) );
  XOR U1101 ( .A(n855), .B(n849), .Z(c[140]) );
  ANDN U1102 ( .B(a[15]), .A(n1634), .Z(n857) );
  AND U1103 ( .A(a[14]), .B(b[1]), .Z(n859) );
  XNOR U1104 ( .A(n859), .B(n858), .Z(n853) );
  XNOR U1105 ( .A(n857), .B(n853), .Z(n862) );
  XOR U1106 ( .A(n861), .B(sreg[141]), .Z(n856) );
  XOR U1107 ( .A(n862), .B(n856), .Z(c[141]) );
  ANDN U1108 ( .B(a[16]), .A(n1634), .Z(n864) );
  AND U1109 ( .A(a[15]), .B(b[1]), .Z(n866) );
  XNOR U1110 ( .A(n866), .B(n865), .Z(n860) );
  XNOR U1111 ( .A(n864), .B(n860), .Z(n869) );
  XOR U1112 ( .A(n868), .B(sreg[142]), .Z(n863) );
  XOR U1113 ( .A(n869), .B(n863), .Z(c[142]) );
  AND U1114 ( .A(a[16]), .B(b[1]), .Z(n873) );
  ANDN U1115 ( .B(a[17]), .A(n1634), .Z(n871) );
  XOR U1116 ( .A(n872), .B(n871), .Z(n867) );
  XNOR U1117 ( .A(n873), .B(n867), .Z(n876) );
  XOR U1118 ( .A(n875), .B(sreg[143]), .Z(n870) );
  XNOR U1119 ( .A(n876), .B(n870), .Z(c[143]) );
  ANDN U1120 ( .B(a[18]), .A(n1634), .Z(n878) );
  AND U1121 ( .A(a[17]), .B(b[1]), .Z(n880) );
  XNOR U1122 ( .A(n880), .B(n879), .Z(n874) );
  XNOR U1123 ( .A(n878), .B(n874), .Z(n883) );
  XOR U1124 ( .A(n882), .B(sreg[144]), .Z(n877) );
  XOR U1125 ( .A(n883), .B(n877), .Z(c[144]) );
  ANDN U1126 ( .B(a[19]), .A(n1634), .Z(n885) );
  AND U1127 ( .A(a[18]), .B(b[1]), .Z(n887) );
  XNOR U1128 ( .A(n887), .B(n886), .Z(n881) );
  XNOR U1129 ( .A(n885), .B(n881), .Z(n890) );
  XOR U1130 ( .A(n889), .B(sreg[145]), .Z(n884) );
  XOR U1131 ( .A(n890), .B(n884), .Z(c[145]) );
  ANDN U1132 ( .B(a[20]), .A(n1634), .Z(n892) );
  AND U1133 ( .A(a[19]), .B(b[1]), .Z(n894) );
  XNOR U1134 ( .A(n894), .B(n893), .Z(n888) );
  XNOR U1135 ( .A(n892), .B(n888), .Z(n897) );
  XOR U1136 ( .A(n896), .B(sreg[146]), .Z(n891) );
  XOR U1137 ( .A(n897), .B(n891), .Z(c[146]) );
  AND U1138 ( .A(a[20]), .B(b[1]), .Z(n901) );
  ANDN U1139 ( .B(a[21]), .A(n1634), .Z(n899) );
  XOR U1140 ( .A(n900), .B(n899), .Z(n895) );
  XNOR U1141 ( .A(n901), .B(n895), .Z(n904) );
  XOR U1142 ( .A(n903), .B(sreg[147]), .Z(n898) );
  XNOR U1143 ( .A(n904), .B(n898), .Z(c[147]) );
  ANDN U1144 ( .B(a[22]), .A(n1634), .Z(n906) );
  AND U1145 ( .A(a[21]), .B(b[1]), .Z(n908) );
  XNOR U1146 ( .A(n908), .B(n907), .Z(n902) );
  XNOR U1147 ( .A(n906), .B(n902), .Z(n911) );
  XOR U1148 ( .A(n910), .B(sreg[148]), .Z(n905) );
  XOR U1149 ( .A(n911), .B(n905), .Z(c[148]) );
  ANDN U1150 ( .B(a[23]), .A(n1634), .Z(n913) );
  AND U1151 ( .A(a[22]), .B(b[1]), .Z(n915) );
  XNOR U1152 ( .A(n914), .B(n915), .Z(n909) );
  XNOR U1153 ( .A(n913), .B(n909), .Z(n918) );
  XOR U1154 ( .A(n917), .B(sreg[149]), .Z(n912) );
  XOR U1155 ( .A(n918), .B(n912), .Z(c[149]) );
  ANDN U1156 ( .B(a[24]), .A(n1634), .Z(n920) );
  AND U1157 ( .A(a[23]), .B(b[1]), .Z(n922) );
  XNOR U1158 ( .A(n922), .B(n921), .Z(n916) );
  XNOR U1159 ( .A(n920), .B(n916), .Z(n925) );
  XOR U1160 ( .A(n924), .B(sreg[150]), .Z(n919) );
  XOR U1161 ( .A(n925), .B(n919), .Z(c[150]) );
  ANDN U1162 ( .B(a[25]), .A(n1634), .Z(n927) );
  AND U1163 ( .A(a[24]), .B(b[1]), .Z(n929) );
  XNOR U1164 ( .A(n928), .B(n929), .Z(n923) );
  XNOR U1165 ( .A(n927), .B(n923), .Z(n932) );
  XOR U1166 ( .A(n931), .B(sreg[151]), .Z(n926) );
  XOR U1167 ( .A(n932), .B(n926), .Z(c[151]) );
  ANDN U1168 ( .B(a[26]), .A(n1634), .Z(n934) );
  AND U1169 ( .A(a[25]), .B(b[1]), .Z(n936) );
  XNOR U1170 ( .A(n936), .B(n935), .Z(n930) );
  XNOR U1171 ( .A(n934), .B(n930), .Z(n939) );
  XOR U1172 ( .A(n938), .B(sreg[152]), .Z(n933) );
  XOR U1173 ( .A(n939), .B(n933), .Z(c[152]) );
  ANDN U1174 ( .B(a[27]), .A(n1634), .Z(n941) );
  AND U1175 ( .A(a[26]), .B(b[1]), .Z(n943) );
  XNOR U1176 ( .A(n943), .B(n942), .Z(n937) );
  XNOR U1177 ( .A(n941), .B(n937), .Z(n946) );
  XOR U1178 ( .A(n945), .B(sreg[153]), .Z(n940) );
  XOR U1179 ( .A(n946), .B(n940), .Z(c[153]) );
  ANDN U1180 ( .B(a[28]), .A(n1634), .Z(n948) );
  AND U1181 ( .A(a[27]), .B(b[1]), .Z(n950) );
  XNOR U1182 ( .A(n950), .B(n949), .Z(n944) );
  XNOR U1183 ( .A(n948), .B(n944), .Z(n953) );
  XOR U1184 ( .A(n952), .B(sreg[154]), .Z(n947) );
  XOR U1185 ( .A(n953), .B(n947), .Z(c[154]) );
  ANDN U1186 ( .B(a[29]), .A(n1634), .Z(n955) );
  AND U1187 ( .A(a[28]), .B(b[1]), .Z(n957) );
  XNOR U1188 ( .A(n957), .B(n956), .Z(n951) );
  XNOR U1189 ( .A(n955), .B(n951), .Z(n960) );
  XOR U1190 ( .A(n959), .B(sreg[155]), .Z(n954) );
  XOR U1191 ( .A(n960), .B(n954), .Z(c[155]) );
  ANDN U1192 ( .B(a[30]), .A(n1634), .Z(n962) );
  AND U1193 ( .A(a[29]), .B(b[1]), .Z(n964) );
  XNOR U1194 ( .A(n964), .B(n963), .Z(n958) );
  XNOR U1195 ( .A(n962), .B(n958), .Z(n967) );
  XOR U1196 ( .A(n966), .B(sreg[156]), .Z(n961) );
  XOR U1197 ( .A(n967), .B(n961), .Z(c[156]) );
  ANDN U1198 ( .B(a[31]), .A(n1634), .Z(n969) );
  AND U1199 ( .A(a[30]), .B(b[1]), .Z(n971) );
  XNOR U1200 ( .A(n971), .B(n970), .Z(n965) );
  XNOR U1201 ( .A(n969), .B(n965), .Z(n974) );
  XOR U1202 ( .A(n973), .B(sreg[157]), .Z(n968) );
  XOR U1203 ( .A(n974), .B(n968), .Z(c[157]) );
  ANDN U1204 ( .B(a[32]), .A(n1634), .Z(n976) );
  AND U1205 ( .A(a[31]), .B(b[1]), .Z(n978) );
  XNOR U1206 ( .A(n978), .B(n977), .Z(n972) );
  XNOR U1207 ( .A(n976), .B(n972), .Z(n981) );
  XOR U1208 ( .A(n980), .B(sreg[158]), .Z(n975) );
  XOR U1209 ( .A(n981), .B(n975), .Z(c[158]) );
  ANDN U1210 ( .B(a[33]), .A(n1634), .Z(n983) );
  AND U1211 ( .A(a[32]), .B(b[1]), .Z(n985) );
  XNOR U1212 ( .A(n985), .B(n984), .Z(n979) );
  XNOR U1213 ( .A(n983), .B(n979), .Z(n988) );
  XOR U1214 ( .A(n987), .B(sreg[159]), .Z(n982) );
  XOR U1215 ( .A(n988), .B(n982), .Z(c[159]) );
  ANDN U1216 ( .B(a[34]), .A(n1634), .Z(n990) );
  AND U1217 ( .A(a[33]), .B(b[1]), .Z(n992) );
  XNOR U1218 ( .A(n992), .B(n991), .Z(n986) );
  XNOR U1219 ( .A(n990), .B(n986), .Z(n995) );
  XOR U1220 ( .A(n994), .B(sreg[160]), .Z(n989) );
  XOR U1221 ( .A(n995), .B(n989), .Z(c[160]) );
  ANDN U1222 ( .B(a[35]), .A(n1634), .Z(n997) );
  AND U1223 ( .A(a[34]), .B(b[1]), .Z(n999) );
  XNOR U1224 ( .A(n999), .B(n998), .Z(n993) );
  XNOR U1225 ( .A(n997), .B(n993), .Z(n1002) );
  XOR U1226 ( .A(n1001), .B(sreg[161]), .Z(n996) );
  XOR U1227 ( .A(n1002), .B(n996), .Z(c[161]) );
  ANDN U1228 ( .B(a[36]), .A(n1634), .Z(n1004) );
  AND U1229 ( .A(a[35]), .B(b[1]), .Z(n1006) );
  XNOR U1230 ( .A(n1006), .B(n1005), .Z(n1000) );
  XNOR U1231 ( .A(n1004), .B(n1000), .Z(n1009) );
  XOR U1232 ( .A(n1008), .B(sreg[162]), .Z(n1003) );
  XOR U1233 ( .A(n1009), .B(n1003), .Z(c[162]) );
  ANDN U1234 ( .B(a[37]), .A(n1634), .Z(n1011) );
  AND U1235 ( .A(a[36]), .B(b[1]), .Z(n1013) );
  XNOR U1236 ( .A(n1013), .B(n1012), .Z(n1007) );
  XNOR U1237 ( .A(n1011), .B(n1007), .Z(n1016) );
  XOR U1238 ( .A(n1015), .B(sreg[163]), .Z(n1010) );
  XOR U1239 ( .A(n1016), .B(n1010), .Z(c[163]) );
  ANDN U1240 ( .B(a[38]), .A(n1634), .Z(n1018) );
  AND U1241 ( .A(a[37]), .B(b[1]), .Z(n1020) );
  XNOR U1242 ( .A(n1020), .B(n1019), .Z(n1014) );
  XNOR U1243 ( .A(n1018), .B(n1014), .Z(n1023) );
  XOR U1244 ( .A(n1022), .B(sreg[164]), .Z(n1017) );
  XOR U1245 ( .A(n1023), .B(n1017), .Z(c[164]) );
  ANDN U1246 ( .B(a[39]), .A(n1634), .Z(n1025) );
  AND U1247 ( .A(a[38]), .B(b[1]), .Z(n1027) );
  XNOR U1248 ( .A(n1027), .B(n1026), .Z(n1021) );
  XNOR U1249 ( .A(n1025), .B(n1021), .Z(n1030) );
  XOR U1250 ( .A(n1029), .B(sreg[165]), .Z(n1024) );
  XOR U1251 ( .A(n1030), .B(n1024), .Z(c[165]) );
  ANDN U1252 ( .B(a[40]), .A(n1634), .Z(n1032) );
  AND U1253 ( .A(a[39]), .B(b[1]), .Z(n1034) );
  XNOR U1254 ( .A(n1034), .B(n1033), .Z(n1028) );
  XNOR U1255 ( .A(n1032), .B(n1028), .Z(n1037) );
  XOR U1256 ( .A(n1036), .B(sreg[166]), .Z(n1031) );
  XOR U1257 ( .A(n1037), .B(n1031), .Z(c[166]) );
  ANDN U1258 ( .B(a[41]), .A(n1634), .Z(n1039) );
  AND U1259 ( .A(a[40]), .B(b[1]), .Z(n1041) );
  XNOR U1260 ( .A(n1041), .B(n1040), .Z(n1035) );
  XNOR U1261 ( .A(n1039), .B(n1035), .Z(n1044) );
  XOR U1262 ( .A(n1043), .B(sreg[167]), .Z(n1038) );
  XOR U1263 ( .A(n1044), .B(n1038), .Z(c[167]) );
  ANDN U1264 ( .B(a[42]), .A(n1634), .Z(n1046) );
  AND U1265 ( .A(a[41]), .B(b[1]), .Z(n1048) );
  XNOR U1266 ( .A(n1048), .B(n1047), .Z(n1042) );
  XNOR U1267 ( .A(n1046), .B(n1042), .Z(n1051) );
  XOR U1268 ( .A(n1050), .B(sreg[168]), .Z(n1045) );
  XOR U1269 ( .A(n1051), .B(n1045), .Z(c[168]) );
  ANDN U1270 ( .B(a[43]), .A(n1634), .Z(n1053) );
  AND U1271 ( .A(a[42]), .B(b[1]), .Z(n1055) );
  XNOR U1272 ( .A(n1055), .B(n1054), .Z(n1049) );
  XNOR U1273 ( .A(n1053), .B(n1049), .Z(n1058) );
  XOR U1274 ( .A(n1057), .B(sreg[169]), .Z(n1052) );
  XOR U1275 ( .A(n1058), .B(n1052), .Z(c[169]) );
  ANDN U1276 ( .B(a[44]), .A(n1634), .Z(n1060) );
  AND U1277 ( .A(a[43]), .B(b[1]), .Z(n1062) );
  XNOR U1278 ( .A(n1062), .B(n1061), .Z(n1056) );
  XNOR U1279 ( .A(n1060), .B(n1056), .Z(n1065) );
  XOR U1280 ( .A(n1064), .B(sreg[170]), .Z(n1059) );
  XOR U1281 ( .A(n1065), .B(n1059), .Z(c[170]) );
  ANDN U1282 ( .B(a[45]), .A(n1634), .Z(n1067) );
  AND U1283 ( .A(a[44]), .B(b[1]), .Z(n1069) );
  XNOR U1284 ( .A(n1069), .B(n1068), .Z(n1063) );
  XNOR U1285 ( .A(n1067), .B(n1063), .Z(n1072) );
  XOR U1286 ( .A(n1071), .B(sreg[171]), .Z(n1066) );
  XOR U1287 ( .A(n1072), .B(n1066), .Z(c[171]) );
  ANDN U1288 ( .B(a[46]), .A(n1634), .Z(n1074) );
  AND U1289 ( .A(a[45]), .B(b[1]), .Z(n1076) );
  XNOR U1290 ( .A(n1076), .B(n1075), .Z(n1070) );
  XNOR U1291 ( .A(n1074), .B(n1070), .Z(n1079) );
  XOR U1292 ( .A(n1078), .B(sreg[172]), .Z(n1073) );
  XOR U1293 ( .A(n1079), .B(n1073), .Z(c[172]) );
  ANDN U1294 ( .B(a[47]), .A(n1634), .Z(n1081) );
  AND U1295 ( .A(a[46]), .B(b[1]), .Z(n1083) );
  XNOR U1296 ( .A(n1083), .B(n1082), .Z(n1077) );
  XNOR U1297 ( .A(n1081), .B(n1077), .Z(n1086) );
  XOR U1298 ( .A(n1085), .B(sreg[173]), .Z(n1080) );
  XOR U1299 ( .A(n1086), .B(n1080), .Z(c[173]) );
  ANDN U1300 ( .B(a[48]), .A(n1634), .Z(n1088) );
  AND U1301 ( .A(a[47]), .B(b[1]), .Z(n1090) );
  XNOR U1302 ( .A(n1090), .B(n1089), .Z(n1084) );
  XNOR U1303 ( .A(n1088), .B(n1084), .Z(n1093) );
  XOR U1304 ( .A(n1092), .B(sreg[174]), .Z(n1087) );
  XOR U1305 ( .A(n1093), .B(n1087), .Z(c[174]) );
  ANDN U1306 ( .B(a[49]), .A(n1634), .Z(n1095) );
  AND U1307 ( .A(a[48]), .B(b[1]), .Z(n1097) );
  XNOR U1308 ( .A(n1097), .B(n1096), .Z(n1091) );
  XNOR U1309 ( .A(n1095), .B(n1091), .Z(n1100) );
  XOR U1310 ( .A(n1099), .B(sreg[175]), .Z(n1094) );
  XOR U1311 ( .A(n1100), .B(n1094), .Z(c[175]) );
  ANDN U1312 ( .B(a[50]), .A(n1634), .Z(n1102) );
  AND U1313 ( .A(a[49]), .B(b[1]), .Z(n1104) );
  XNOR U1314 ( .A(n1104), .B(n1103), .Z(n1098) );
  XNOR U1315 ( .A(n1102), .B(n1098), .Z(n1107) );
  XOR U1316 ( .A(n1106), .B(sreg[176]), .Z(n1101) );
  XOR U1317 ( .A(n1107), .B(n1101), .Z(c[176]) );
  ANDN U1318 ( .B(a[51]), .A(n1634), .Z(n1109) );
  AND U1319 ( .A(a[50]), .B(b[1]), .Z(n1111) );
  XNOR U1320 ( .A(n1111), .B(n1110), .Z(n1105) );
  XNOR U1321 ( .A(n1109), .B(n1105), .Z(n1114) );
  XOR U1322 ( .A(n1113), .B(sreg[177]), .Z(n1108) );
  XOR U1323 ( .A(n1114), .B(n1108), .Z(c[177]) );
  ANDN U1324 ( .B(a[52]), .A(n1634), .Z(n1116) );
  AND U1325 ( .A(a[51]), .B(b[1]), .Z(n1118) );
  XNOR U1326 ( .A(n1118), .B(n1117), .Z(n1112) );
  XNOR U1327 ( .A(n1116), .B(n1112), .Z(n1121) );
  XOR U1328 ( .A(n1120), .B(sreg[178]), .Z(n1115) );
  XOR U1329 ( .A(n1121), .B(n1115), .Z(c[178]) );
  ANDN U1330 ( .B(a[53]), .A(n1634), .Z(n1123) );
  AND U1331 ( .A(a[52]), .B(b[1]), .Z(n1125) );
  XNOR U1332 ( .A(n1125), .B(n1124), .Z(n1119) );
  XNOR U1333 ( .A(n1123), .B(n1119), .Z(n1128) );
  XOR U1334 ( .A(n1127), .B(sreg[179]), .Z(n1122) );
  XOR U1335 ( .A(n1128), .B(n1122), .Z(c[179]) );
  ANDN U1336 ( .B(a[54]), .A(n1634), .Z(n1130) );
  AND U1337 ( .A(a[53]), .B(b[1]), .Z(n1132) );
  XNOR U1338 ( .A(n1132), .B(n1131), .Z(n1126) );
  XNOR U1339 ( .A(n1130), .B(n1126), .Z(n1135) );
  XOR U1340 ( .A(n1134), .B(sreg[180]), .Z(n1129) );
  XOR U1341 ( .A(n1135), .B(n1129), .Z(c[180]) );
  ANDN U1342 ( .B(a[55]), .A(n1634), .Z(n1137) );
  AND U1343 ( .A(a[54]), .B(b[1]), .Z(n1139) );
  XNOR U1344 ( .A(n1139), .B(n1138), .Z(n1133) );
  XNOR U1345 ( .A(n1137), .B(n1133), .Z(n1142) );
  XOR U1346 ( .A(n1141), .B(sreg[181]), .Z(n1136) );
  XOR U1347 ( .A(n1142), .B(n1136), .Z(c[181]) );
  ANDN U1348 ( .B(a[56]), .A(n1634), .Z(n1144) );
  AND U1349 ( .A(a[55]), .B(b[1]), .Z(n1146) );
  XNOR U1350 ( .A(n1146), .B(n1145), .Z(n1140) );
  XNOR U1351 ( .A(n1144), .B(n1140), .Z(n1149) );
  XOR U1352 ( .A(n1148), .B(sreg[182]), .Z(n1143) );
  XOR U1353 ( .A(n1149), .B(n1143), .Z(c[182]) );
  ANDN U1354 ( .B(a[57]), .A(n1634), .Z(n1151) );
  AND U1355 ( .A(a[56]), .B(b[1]), .Z(n1153) );
  XNOR U1356 ( .A(n1153), .B(n1152), .Z(n1147) );
  XNOR U1357 ( .A(n1151), .B(n1147), .Z(n1156) );
  XOR U1358 ( .A(n1155), .B(sreg[183]), .Z(n1150) );
  XOR U1359 ( .A(n1156), .B(n1150), .Z(c[183]) );
  ANDN U1360 ( .B(a[58]), .A(n1634), .Z(n1158) );
  AND U1361 ( .A(a[57]), .B(b[1]), .Z(n1160) );
  XNOR U1362 ( .A(n1160), .B(n1159), .Z(n1154) );
  XNOR U1363 ( .A(n1158), .B(n1154), .Z(n1163) );
  XOR U1364 ( .A(n1162), .B(sreg[184]), .Z(n1157) );
  XOR U1365 ( .A(n1163), .B(n1157), .Z(c[184]) );
  ANDN U1366 ( .B(a[59]), .A(n1634), .Z(n1165) );
  AND U1367 ( .A(a[58]), .B(b[1]), .Z(n1167) );
  XNOR U1368 ( .A(n1167), .B(n1166), .Z(n1161) );
  XNOR U1369 ( .A(n1165), .B(n1161), .Z(n1170) );
  XOR U1370 ( .A(n1169), .B(sreg[185]), .Z(n1164) );
  XOR U1371 ( .A(n1170), .B(n1164), .Z(c[185]) );
  ANDN U1372 ( .B(a[60]), .A(n1634), .Z(n1172) );
  AND U1373 ( .A(a[59]), .B(b[1]), .Z(n1174) );
  XNOR U1374 ( .A(n1174), .B(n1173), .Z(n1168) );
  XNOR U1375 ( .A(n1172), .B(n1168), .Z(n1177) );
  XOR U1376 ( .A(n1176), .B(sreg[186]), .Z(n1171) );
  XOR U1377 ( .A(n1177), .B(n1171), .Z(c[186]) );
  ANDN U1378 ( .B(a[61]), .A(n1634), .Z(n1179) );
  AND U1379 ( .A(a[60]), .B(b[1]), .Z(n1181) );
  XNOR U1380 ( .A(n1181), .B(n1180), .Z(n1175) );
  XNOR U1381 ( .A(n1179), .B(n1175), .Z(n1184) );
  XOR U1382 ( .A(n1183), .B(sreg[187]), .Z(n1178) );
  XOR U1383 ( .A(n1184), .B(n1178), .Z(c[187]) );
  ANDN U1384 ( .B(a[62]), .A(n1634), .Z(n1186) );
  AND U1385 ( .A(a[61]), .B(b[1]), .Z(n1188) );
  XNOR U1386 ( .A(n1188), .B(n1187), .Z(n1182) );
  XNOR U1387 ( .A(n1186), .B(n1182), .Z(n1191) );
  XOR U1388 ( .A(n1190), .B(sreg[188]), .Z(n1185) );
  XOR U1389 ( .A(n1191), .B(n1185), .Z(c[188]) );
  ANDN U1390 ( .B(a[63]), .A(n1634), .Z(n1193) );
  AND U1391 ( .A(a[62]), .B(b[1]), .Z(n1195) );
  XNOR U1392 ( .A(n1195), .B(n1194), .Z(n1189) );
  XNOR U1393 ( .A(n1193), .B(n1189), .Z(n1198) );
  XOR U1394 ( .A(n1197), .B(sreg[189]), .Z(n1192) );
  XOR U1395 ( .A(n1198), .B(n1192), .Z(c[189]) );
  ANDN U1396 ( .B(a[64]), .A(n1634), .Z(n1200) );
  AND U1397 ( .A(a[63]), .B(b[1]), .Z(n1202) );
  XNOR U1398 ( .A(n1202), .B(n1201), .Z(n1196) );
  XNOR U1399 ( .A(n1200), .B(n1196), .Z(n1205) );
  XOR U1400 ( .A(n1204), .B(sreg[190]), .Z(n1199) );
  XOR U1401 ( .A(n1205), .B(n1199), .Z(c[190]) );
  ANDN U1402 ( .B(a[65]), .A(n1634), .Z(n1207) );
  AND U1403 ( .A(a[64]), .B(b[1]), .Z(n1209) );
  XNOR U1404 ( .A(n1209), .B(n1208), .Z(n1203) );
  XNOR U1405 ( .A(n1207), .B(n1203), .Z(n1212) );
  XOR U1406 ( .A(n1211), .B(sreg[191]), .Z(n1206) );
  XOR U1407 ( .A(n1212), .B(n1206), .Z(c[191]) );
  ANDN U1408 ( .B(a[66]), .A(n1634), .Z(n1214) );
  AND U1409 ( .A(a[65]), .B(b[1]), .Z(n1216) );
  XNOR U1410 ( .A(n1216), .B(n1215), .Z(n1210) );
  XNOR U1411 ( .A(n1214), .B(n1210), .Z(n1219) );
  XOR U1412 ( .A(n1218), .B(sreg[192]), .Z(n1213) );
  XOR U1413 ( .A(n1219), .B(n1213), .Z(c[192]) );
  ANDN U1414 ( .B(a[67]), .A(n1634), .Z(n1221) );
  AND U1415 ( .A(a[66]), .B(b[1]), .Z(n1223) );
  XNOR U1416 ( .A(n1223), .B(n1222), .Z(n1217) );
  XNOR U1417 ( .A(n1221), .B(n1217), .Z(n1226) );
  XOR U1418 ( .A(n1225), .B(sreg[193]), .Z(n1220) );
  XOR U1419 ( .A(n1226), .B(n1220), .Z(c[193]) );
  ANDN U1420 ( .B(a[68]), .A(n1634), .Z(n1228) );
  AND U1421 ( .A(a[67]), .B(b[1]), .Z(n1230) );
  XNOR U1422 ( .A(n1230), .B(n1229), .Z(n1224) );
  XNOR U1423 ( .A(n1228), .B(n1224), .Z(n1233) );
  XOR U1424 ( .A(n1232), .B(sreg[194]), .Z(n1227) );
  XOR U1425 ( .A(n1233), .B(n1227), .Z(c[194]) );
  ANDN U1426 ( .B(a[69]), .A(n1634), .Z(n1235) );
  AND U1427 ( .A(a[68]), .B(b[1]), .Z(n1237) );
  XNOR U1428 ( .A(n1237), .B(n1236), .Z(n1231) );
  XNOR U1429 ( .A(n1235), .B(n1231), .Z(n1240) );
  XOR U1430 ( .A(n1239), .B(sreg[195]), .Z(n1234) );
  XOR U1431 ( .A(n1240), .B(n1234), .Z(c[195]) );
  ANDN U1432 ( .B(a[70]), .A(n1634), .Z(n1242) );
  AND U1433 ( .A(a[69]), .B(b[1]), .Z(n1244) );
  XNOR U1434 ( .A(n1244), .B(n1243), .Z(n1238) );
  XNOR U1435 ( .A(n1242), .B(n1238), .Z(n1247) );
  XOR U1436 ( .A(n1246), .B(sreg[196]), .Z(n1241) );
  XOR U1437 ( .A(n1247), .B(n1241), .Z(c[196]) );
  ANDN U1438 ( .B(a[71]), .A(n1634), .Z(n1249) );
  AND U1439 ( .A(a[70]), .B(b[1]), .Z(n1251) );
  XNOR U1440 ( .A(n1251), .B(n1250), .Z(n1245) );
  XNOR U1441 ( .A(n1249), .B(n1245), .Z(n1254) );
  XOR U1442 ( .A(n1253), .B(sreg[197]), .Z(n1248) );
  XOR U1443 ( .A(n1254), .B(n1248), .Z(c[197]) );
  ANDN U1444 ( .B(a[72]), .A(n1634), .Z(n1256) );
  AND U1445 ( .A(a[71]), .B(b[1]), .Z(n1258) );
  XNOR U1446 ( .A(n1258), .B(n1257), .Z(n1252) );
  XNOR U1447 ( .A(n1256), .B(n1252), .Z(n1261) );
  XOR U1448 ( .A(n1260), .B(sreg[198]), .Z(n1255) );
  XOR U1449 ( .A(n1261), .B(n1255), .Z(c[198]) );
  ANDN U1450 ( .B(a[73]), .A(n1634), .Z(n1263) );
  AND U1451 ( .A(a[72]), .B(b[1]), .Z(n1265) );
  XNOR U1452 ( .A(n1265), .B(n1264), .Z(n1259) );
  XNOR U1453 ( .A(n1263), .B(n1259), .Z(n1268) );
  XOR U1454 ( .A(n1267), .B(sreg[199]), .Z(n1262) );
  XOR U1455 ( .A(n1268), .B(n1262), .Z(c[199]) );
  ANDN U1456 ( .B(a[74]), .A(n1634), .Z(n1270) );
  AND U1457 ( .A(a[73]), .B(b[1]), .Z(n1272) );
  XNOR U1458 ( .A(n1272), .B(n1271), .Z(n1266) );
  XNOR U1459 ( .A(n1270), .B(n1266), .Z(n1275) );
  XOR U1460 ( .A(n1274), .B(sreg[200]), .Z(n1269) );
  XOR U1461 ( .A(n1275), .B(n1269), .Z(c[200]) );
  ANDN U1462 ( .B(a[75]), .A(n1634), .Z(n1277) );
  AND U1463 ( .A(a[74]), .B(b[1]), .Z(n1279) );
  XNOR U1464 ( .A(n1279), .B(n1278), .Z(n1273) );
  XNOR U1465 ( .A(n1277), .B(n1273), .Z(n1282) );
  XOR U1466 ( .A(n1281), .B(sreg[201]), .Z(n1276) );
  XOR U1467 ( .A(n1282), .B(n1276), .Z(c[201]) );
  ANDN U1468 ( .B(a[76]), .A(n1634), .Z(n1284) );
  AND U1469 ( .A(a[75]), .B(b[1]), .Z(n1286) );
  XNOR U1470 ( .A(n1286), .B(n1285), .Z(n1280) );
  XNOR U1471 ( .A(n1284), .B(n1280), .Z(n1289) );
  XOR U1472 ( .A(n1288), .B(sreg[202]), .Z(n1283) );
  XOR U1473 ( .A(n1289), .B(n1283), .Z(c[202]) );
  ANDN U1474 ( .B(a[77]), .A(n1634), .Z(n1291) );
  AND U1475 ( .A(a[76]), .B(b[1]), .Z(n1293) );
  XNOR U1476 ( .A(n1293), .B(n1292), .Z(n1287) );
  XNOR U1477 ( .A(n1291), .B(n1287), .Z(n1296) );
  XOR U1478 ( .A(n1295), .B(sreg[203]), .Z(n1290) );
  XOR U1479 ( .A(n1296), .B(n1290), .Z(c[203]) );
  ANDN U1480 ( .B(a[78]), .A(n1634), .Z(n1298) );
  AND U1481 ( .A(a[77]), .B(b[1]), .Z(n1300) );
  XNOR U1482 ( .A(n1300), .B(n1299), .Z(n1294) );
  XNOR U1483 ( .A(n1298), .B(n1294), .Z(n1303) );
  XOR U1484 ( .A(n1302), .B(sreg[204]), .Z(n1297) );
  XOR U1485 ( .A(n1303), .B(n1297), .Z(c[204]) );
  ANDN U1486 ( .B(a[79]), .A(n1634), .Z(n1305) );
  AND U1487 ( .A(a[78]), .B(b[1]), .Z(n1307) );
  XNOR U1488 ( .A(n1307), .B(n1306), .Z(n1301) );
  XNOR U1489 ( .A(n1305), .B(n1301), .Z(n1310) );
  XOR U1490 ( .A(n1309), .B(sreg[205]), .Z(n1304) );
  XOR U1491 ( .A(n1310), .B(n1304), .Z(c[205]) );
  ANDN U1492 ( .B(a[80]), .A(n1634), .Z(n1312) );
  AND U1493 ( .A(a[79]), .B(b[1]), .Z(n1314) );
  XNOR U1494 ( .A(n1314), .B(n1313), .Z(n1308) );
  XNOR U1495 ( .A(n1312), .B(n1308), .Z(n1317) );
  XOR U1496 ( .A(n1316), .B(sreg[206]), .Z(n1311) );
  XOR U1497 ( .A(n1317), .B(n1311), .Z(c[206]) );
  ANDN U1498 ( .B(a[81]), .A(n1634), .Z(n1319) );
  AND U1499 ( .A(a[80]), .B(b[1]), .Z(n1321) );
  XNOR U1500 ( .A(n1321), .B(n1320), .Z(n1315) );
  XNOR U1501 ( .A(n1319), .B(n1315), .Z(n1324) );
  XOR U1502 ( .A(n1323), .B(sreg[207]), .Z(n1318) );
  XOR U1503 ( .A(n1324), .B(n1318), .Z(c[207]) );
  ANDN U1504 ( .B(a[82]), .A(n1634), .Z(n1326) );
  AND U1505 ( .A(a[81]), .B(b[1]), .Z(n1328) );
  XNOR U1506 ( .A(n1328), .B(n1327), .Z(n1322) );
  XNOR U1507 ( .A(n1326), .B(n1322), .Z(n1331) );
  XOR U1508 ( .A(n1330), .B(sreg[208]), .Z(n1325) );
  XOR U1509 ( .A(n1331), .B(n1325), .Z(c[208]) );
  ANDN U1510 ( .B(a[83]), .A(n1634), .Z(n1333) );
  AND U1511 ( .A(a[82]), .B(b[1]), .Z(n1335) );
  XNOR U1512 ( .A(n1335), .B(n1334), .Z(n1329) );
  XNOR U1513 ( .A(n1333), .B(n1329), .Z(n1338) );
  XOR U1514 ( .A(n1337), .B(sreg[209]), .Z(n1332) );
  XOR U1515 ( .A(n1338), .B(n1332), .Z(c[209]) );
  ANDN U1516 ( .B(a[84]), .A(n1634), .Z(n1340) );
  AND U1517 ( .A(a[83]), .B(b[1]), .Z(n1342) );
  XNOR U1518 ( .A(n1342), .B(n1341), .Z(n1336) );
  XNOR U1519 ( .A(n1340), .B(n1336), .Z(n1345) );
  XOR U1520 ( .A(n1344), .B(sreg[210]), .Z(n1339) );
  XOR U1521 ( .A(n1345), .B(n1339), .Z(c[210]) );
  ANDN U1522 ( .B(a[85]), .A(n1634), .Z(n1347) );
  AND U1523 ( .A(a[84]), .B(b[1]), .Z(n1349) );
  XNOR U1524 ( .A(n1349), .B(n1348), .Z(n1343) );
  XNOR U1525 ( .A(n1347), .B(n1343), .Z(n1352) );
  XOR U1526 ( .A(n1351), .B(sreg[211]), .Z(n1346) );
  XOR U1527 ( .A(n1352), .B(n1346), .Z(c[211]) );
  ANDN U1528 ( .B(a[86]), .A(n1634), .Z(n1354) );
  AND U1529 ( .A(a[85]), .B(b[1]), .Z(n1356) );
  XNOR U1530 ( .A(n1356), .B(n1355), .Z(n1350) );
  XNOR U1531 ( .A(n1354), .B(n1350), .Z(n1359) );
  XOR U1532 ( .A(n1358), .B(sreg[212]), .Z(n1353) );
  XOR U1533 ( .A(n1359), .B(n1353), .Z(c[212]) );
  ANDN U1534 ( .B(a[87]), .A(n1634), .Z(n1361) );
  AND U1535 ( .A(a[86]), .B(b[1]), .Z(n1363) );
  XNOR U1536 ( .A(n1363), .B(n1362), .Z(n1357) );
  XNOR U1537 ( .A(n1361), .B(n1357), .Z(n1366) );
  XOR U1538 ( .A(n1365), .B(sreg[213]), .Z(n1360) );
  XOR U1539 ( .A(n1366), .B(n1360), .Z(c[213]) );
  ANDN U1540 ( .B(a[88]), .A(n1634), .Z(n1368) );
  AND U1541 ( .A(a[87]), .B(b[1]), .Z(n1370) );
  XNOR U1542 ( .A(n1370), .B(n1369), .Z(n1364) );
  XNOR U1543 ( .A(n1368), .B(n1364), .Z(n1373) );
  XOR U1544 ( .A(n1372), .B(sreg[214]), .Z(n1367) );
  XOR U1545 ( .A(n1373), .B(n1367), .Z(c[214]) );
  ANDN U1546 ( .B(a[89]), .A(n1634), .Z(n1375) );
  AND U1547 ( .A(a[88]), .B(b[1]), .Z(n1377) );
  XNOR U1548 ( .A(n1377), .B(n1376), .Z(n1371) );
  XNOR U1549 ( .A(n1375), .B(n1371), .Z(n1380) );
  XOR U1550 ( .A(n1379), .B(sreg[215]), .Z(n1374) );
  XOR U1551 ( .A(n1380), .B(n1374), .Z(c[215]) );
  ANDN U1552 ( .B(a[90]), .A(n1634), .Z(n1382) );
  AND U1553 ( .A(a[89]), .B(b[1]), .Z(n1384) );
  XNOR U1554 ( .A(n1384), .B(n1383), .Z(n1378) );
  XNOR U1555 ( .A(n1382), .B(n1378), .Z(n1387) );
  XOR U1556 ( .A(n1386), .B(sreg[216]), .Z(n1381) );
  XOR U1557 ( .A(n1387), .B(n1381), .Z(c[216]) );
  ANDN U1558 ( .B(a[91]), .A(n1634), .Z(n1389) );
  AND U1559 ( .A(a[90]), .B(b[1]), .Z(n1391) );
  XNOR U1560 ( .A(n1391), .B(n1390), .Z(n1385) );
  XNOR U1561 ( .A(n1389), .B(n1385), .Z(n1394) );
  XOR U1562 ( .A(n1393), .B(sreg[217]), .Z(n1388) );
  XOR U1563 ( .A(n1394), .B(n1388), .Z(c[217]) );
  ANDN U1564 ( .B(a[92]), .A(n1634), .Z(n1396) );
  AND U1565 ( .A(a[91]), .B(b[1]), .Z(n1398) );
  XNOR U1566 ( .A(n1398), .B(n1397), .Z(n1392) );
  XNOR U1567 ( .A(n1396), .B(n1392), .Z(n1401) );
  XOR U1568 ( .A(n1400), .B(sreg[218]), .Z(n1395) );
  XOR U1569 ( .A(n1401), .B(n1395), .Z(c[218]) );
  ANDN U1570 ( .B(a[93]), .A(n1634), .Z(n1403) );
  AND U1571 ( .A(a[92]), .B(b[1]), .Z(n1405) );
  XNOR U1572 ( .A(n1405), .B(n1404), .Z(n1399) );
  XNOR U1573 ( .A(n1403), .B(n1399), .Z(n1408) );
  XOR U1574 ( .A(n1407), .B(sreg[219]), .Z(n1402) );
  XOR U1575 ( .A(n1408), .B(n1402), .Z(c[219]) );
  ANDN U1576 ( .B(a[94]), .A(n1634), .Z(n1410) );
  AND U1577 ( .A(a[93]), .B(b[1]), .Z(n1412) );
  XNOR U1578 ( .A(n1412), .B(n1411), .Z(n1406) );
  XNOR U1579 ( .A(n1410), .B(n1406), .Z(n1415) );
  XOR U1580 ( .A(n1414), .B(sreg[220]), .Z(n1409) );
  XOR U1581 ( .A(n1415), .B(n1409), .Z(c[220]) );
  ANDN U1582 ( .B(a[95]), .A(n1634), .Z(n1417) );
  AND U1583 ( .A(a[94]), .B(b[1]), .Z(n1419) );
  XNOR U1584 ( .A(n1419), .B(n1418), .Z(n1413) );
  XNOR U1585 ( .A(n1417), .B(n1413), .Z(n1422) );
  XOR U1586 ( .A(n1421), .B(sreg[221]), .Z(n1416) );
  XOR U1587 ( .A(n1422), .B(n1416), .Z(c[221]) );
  ANDN U1588 ( .B(a[96]), .A(n1634), .Z(n1424) );
  AND U1589 ( .A(a[95]), .B(b[1]), .Z(n1426) );
  XNOR U1590 ( .A(n1426), .B(n1425), .Z(n1420) );
  XNOR U1591 ( .A(n1424), .B(n1420), .Z(n1429) );
  XOR U1592 ( .A(n1428), .B(sreg[222]), .Z(n1423) );
  XOR U1593 ( .A(n1429), .B(n1423), .Z(c[222]) );
  ANDN U1594 ( .B(a[97]), .A(n1634), .Z(n1431) );
  AND U1595 ( .A(a[96]), .B(b[1]), .Z(n1433) );
  XNOR U1596 ( .A(n1433), .B(n1432), .Z(n1427) );
  XNOR U1597 ( .A(n1431), .B(n1427), .Z(n1436) );
  XOR U1598 ( .A(n1435), .B(sreg[223]), .Z(n1430) );
  XOR U1599 ( .A(n1436), .B(n1430), .Z(c[223]) );
  ANDN U1600 ( .B(a[98]), .A(n1634), .Z(n1438) );
  AND U1601 ( .A(a[97]), .B(b[1]), .Z(n1440) );
  XNOR U1602 ( .A(n1440), .B(n1439), .Z(n1434) );
  XNOR U1603 ( .A(n1438), .B(n1434), .Z(n1443) );
  XOR U1604 ( .A(n1442), .B(sreg[224]), .Z(n1437) );
  XOR U1605 ( .A(n1443), .B(n1437), .Z(c[224]) );
  ANDN U1606 ( .B(a[99]), .A(n1634), .Z(n1445) );
  AND U1607 ( .A(a[98]), .B(b[1]), .Z(n1447) );
  XNOR U1608 ( .A(n1447), .B(n1446), .Z(n1441) );
  XNOR U1609 ( .A(n1445), .B(n1441), .Z(n1450) );
  XOR U1610 ( .A(n1449), .B(sreg[225]), .Z(n1444) );
  XOR U1611 ( .A(n1450), .B(n1444), .Z(c[225]) );
  ANDN U1612 ( .B(a[100]), .A(n1634), .Z(n1452) );
  AND U1613 ( .A(a[99]), .B(b[1]), .Z(n1454) );
  XNOR U1614 ( .A(n1454), .B(n1453), .Z(n1448) );
  XNOR U1615 ( .A(n1452), .B(n1448), .Z(n1457) );
  XOR U1616 ( .A(n1456), .B(sreg[226]), .Z(n1451) );
  XOR U1617 ( .A(n1457), .B(n1451), .Z(c[226]) );
  ANDN U1618 ( .B(a[101]), .A(n1634), .Z(n1459) );
  AND U1619 ( .A(a[100]), .B(b[1]), .Z(n1461) );
  XNOR U1620 ( .A(n1461), .B(n1460), .Z(n1455) );
  XNOR U1621 ( .A(n1459), .B(n1455), .Z(n1464) );
  XOR U1622 ( .A(n1463), .B(sreg[227]), .Z(n1458) );
  XOR U1623 ( .A(n1464), .B(n1458), .Z(c[227]) );
  ANDN U1624 ( .B(a[102]), .A(n1634), .Z(n1466) );
  AND U1625 ( .A(a[101]), .B(b[1]), .Z(n1468) );
  XNOR U1626 ( .A(n1468), .B(n1467), .Z(n1462) );
  XNOR U1627 ( .A(n1466), .B(n1462), .Z(n1471) );
  XOR U1628 ( .A(n1470), .B(sreg[228]), .Z(n1465) );
  XOR U1629 ( .A(n1471), .B(n1465), .Z(c[228]) );
  ANDN U1630 ( .B(a[103]), .A(n1634), .Z(n1473) );
  AND U1631 ( .A(a[102]), .B(b[1]), .Z(n1475) );
  XNOR U1632 ( .A(n1475), .B(n1474), .Z(n1469) );
  XNOR U1633 ( .A(n1473), .B(n1469), .Z(n1478) );
  XOR U1634 ( .A(n1477), .B(sreg[229]), .Z(n1472) );
  XOR U1635 ( .A(n1478), .B(n1472), .Z(c[229]) );
  ANDN U1636 ( .B(a[104]), .A(n1634), .Z(n1480) );
  AND U1637 ( .A(a[103]), .B(b[1]), .Z(n1482) );
  XNOR U1638 ( .A(n1482), .B(n1481), .Z(n1476) );
  XNOR U1639 ( .A(n1480), .B(n1476), .Z(n1485) );
  XOR U1640 ( .A(n1484), .B(sreg[230]), .Z(n1479) );
  XOR U1641 ( .A(n1485), .B(n1479), .Z(c[230]) );
  ANDN U1642 ( .B(a[105]), .A(n1634), .Z(n1487) );
  AND U1643 ( .A(a[104]), .B(b[1]), .Z(n1489) );
  XNOR U1644 ( .A(n1489), .B(n1488), .Z(n1483) );
  XNOR U1645 ( .A(n1487), .B(n1483), .Z(n1492) );
  XOR U1646 ( .A(n1491), .B(sreg[231]), .Z(n1486) );
  XOR U1647 ( .A(n1492), .B(n1486), .Z(c[231]) );
  ANDN U1648 ( .B(a[106]), .A(n1634), .Z(n1494) );
  AND U1649 ( .A(a[105]), .B(b[1]), .Z(n1496) );
  XNOR U1650 ( .A(n1496), .B(n1495), .Z(n1490) );
  XNOR U1651 ( .A(n1494), .B(n1490), .Z(n1499) );
  XOR U1652 ( .A(n1498), .B(sreg[232]), .Z(n1493) );
  XOR U1653 ( .A(n1499), .B(n1493), .Z(c[232]) );
  ANDN U1654 ( .B(a[107]), .A(n1634), .Z(n1501) );
  AND U1655 ( .A(a[106]), .B(b[1]), .Z(n1503) );
  XNOR U1656 ( .A(n1503), .B(n1502), .Z(n1497) );
  XNOR U1657 ( .A(n1501), .B(n1497), .Z(n1506) );
  XOR U1658 ( .A(n1505), .B(sreg[233]), .Z(n1500) );
  XOR U1659 ( .A(n1506), .B(n1500), .Z(c[233]) );
  ANDN U1660 ( .B(a[108]), .A(n1634), .Z(n1508) );
  AND U1661 ( .A(a[107]), .B(b[1]), .Z(n1510) );
  XNOR U1662 ( .A(n1510), .B(n1509), .Z(n1504) );
  XNOR U1663 ( .A(n1508), .B(n1504), .Z(n1513) );
  XOR U1664 ( .A(n1512), .B(sreg[234]), .Z(n1507) );
  XOR U1665 ( .A(n1513), .B(n1507), .Z(c[234]) );
  ANDN U1666 ( .B(a[109]), .A(n1634), .Z(n1515) );
  AND U1667 ( .A(a[108]), .B(b[1]), .Z(n1517) );
  XNOR U1668 ( .A(n1517), .B(n1516), .Z(n1511) );
  XNOR U1669 ( .A(n1515), .B(n1511), .Z(n1520) );
  XOR U1670 ( .A(n1519), .B(sreg[235]), .Z(n1514) );
  XOR U1671 ( .A(n1520), .B(n1514), .Z(c[235]) );
  ANDN U1672 ( .B(a[110]), .A(n1634), .Z(n1522) );
  AND U1673 ( .A(a[109]), .B(b[1]), .Z(n1524) );
  XNOR U1674 ( .A(n1524), .B(n1523), .Z(n1518) );
  XNOR U1675 ( .A(n1522), .B(n1518), .Z(n1527) );
  XOR U1676 ( .A(n1526), .B(sreg[236]), .Z(n1521) );
  XOR U1677 ( .A(n1527), .B(n1521), .Z(c[236]) );
  ANDN U1678 ( .B(a[111]), .A(n1634), .Z(n1529) );
  AND U1679 ( .A(a[110]), .B(b[1]), .Z(n1531) );
  XNOR U1680 ( .A(n1531), .B(n1530), .Z(n1525) );
  XNOR U1681 ( .A(n1529), .B(n1525), .Z(n1534) );
  XOR U1682 ( .A(n1533), .B(sreg[237]), .Z(n1528) );
  XOR U1683 ( .A(n1534), .B(n1528), .Z(c[237]) );
  ANDN U1684 ( .B(a[112]), .A(n1634), .Z(n1536) );
  AND U1685 ( .A(a[111]), .B(b[1]), .Z(n1538) );
  XNOR U1686 ( .A(n1538), .B(n1537), .Z(n1532) );
  XNOR U1687 ( .A(n1536), .B(n1532), .Z(n1541) );
  XOR U1688 ( .A(n1540), .B(sreg[238]), .Z(n1535) );
  XOR U1689 ( .A(n1541), .B(n1535), .Z(c[238]) );
  ANDN U1690 ( .B(a[113]), .A(n1634), .Z(n1543) );
  AND U1691 ( .A(a[112]), .B(b[1]), .Z(n1545) );
  XNOR U1692 ( .A(n1545), .B(n1544), .Z(n1539) );
  XNOR U1693 ( .A(n1543), .B(n1539), .Z(n1548) );
  XOR U1694 ( .A(n1547), .B(sreg[239]), .Z(n1542) );
  XOR U1695 ( .A(n1548), .B(n1542), .Z(c[239]) );
  ANDN U1696 ( .B(a[114]), .A(n1634), .Z(n1550) );
  AND U1697 ( .A(a[113]), .B(b[1]), .Z(n1552) );
  XNOR U1698 ( .A(n1552), .B(n1551), .Z(n1546) );
  XNOR U1699 ( .A(n1550), .B(n1546), .Z(n1555) );
  XOR U1700 ( .A(n1554), .B(sreg[240]), .Z(n1549) );
  XOR U1701 ( .A(n1555), .B(n1549), .Z(c[240]) );
  ANDN U1702 ( .B(a[115]), .A(n1634), .Z(n1557) );
  AND U1703 ( .A(a[114]), .B(b[1]), .Z(n1559) );
  XNOR U1704 ( .A(n1559), .B(n1558), .Z(n1553) );
  XNOR U1705 ( .A(n1557), .B(n1553), .Z(n1562) );
  XOR U1706 ( .A(n1561), .B(sreg[241]), .Z(n1556) );
  XOR U1707 ( .A(n1562), .B(n1556), .Z(c[241]) );
  ANDN U1708 ( .B(a[116]), .A(n1634), .Z(n1564) );
  AND U1709 ( .A(a[115]), .B(b[1]), .Z(n1566) );
  XNOR U1710 ( .A(n1566), .B(n1565), .Z(n1560) );
  XNOR U1711 ( .A(n1564), .B(n1560), .Z(n1569) );
  XOR U1712 ( .A(n1568), .B(sreg[242]), .Z(n1563) );
  XOR U1713 ( .A(n1569), .B(n1563), .Z(c[242]) );
  ANDN U1714 ( .B(a[117]), .A(n1634), .Z(n1571) );
  AND U1715 ( .A(a[116]), .B(b[1]), .Z(n1573) );
  XNOR U1716 ( .A(n1573), .B(n1572), .Z(n1567) );
  XNOR U1717 ( .A(n1571), .B(n1567), .Z(n1576) );
  XOR U1718 ( .A(n1575), .B(sreg[243]), .Z(n1570) );
  XOR U1719 ( .A(n1576), .B(n1570), .Z(c[243]) );
  ANDN U1720 ( .B(a[118]), .A(n1634), .Z(n1578) );
  AND U1721 ( .A(a[117]), .B(b[1]), .Z(n1580) );
  XNOR U1722 ( .A(n1580), .B(n1579), .Z(n1574) );
  XNOR U1723 ( .A(n1578), .B(n1574), .Z(n1583) );
  XOR U1724 ( .A(n1582), .B(sreg[244]), .Z(n1577) );
  XOR U1725 ( .A(n1583), .B(n1577), .Z(c[244]) );
  ANDN U1726 ( .B(a[119]), .A(n1634), .Z(n1585) );
  AND U1727 ( .A(a[118]), .B(b[1]), .Z(n1587) );
  XNOR U1728 ( .A(n1587), .B(n1586), .Z(n1581) );
  XNOR U1729 ( .A(n1585), .B(n1581), .Z(n1590) );
  XOR U1730 ( .A(n1589), .B(sreg[245]), .Z(n1584) );
  XOR U1731 ( .A(n1590), .B(n1584), .Z(c[245]) );
  ANDN U1732 ( .B(a[120]), .A(n1634), .Z(n1592) );
  AND U1733 ( .A(a[119]), .B(b[1]), .Z(n1594) );
  XNOR U1734 ( .A(n1594), .B(n1593), .Z(n1588) );
  XNOR U1735 ( .A(n1592), .B(n1588), .Z(n1597) );
  XOR U1736 ( .A(n1596), .B(sreg[246]), .Z(n1591) );
  XOR U1737 ( .A(n1597), .B(n1591), .Z(c[246]) );
  ANDN U1738 ( .B(a[121]), .A(n1634), .Z(n1599) );
  AND U1739 ( .A(a[120]), .B(b[1]), .Z(n1601) );
  XNOR U1740 ( .A(n1601), .B(n1600), .Z(n1595) );
  XNOR U1741 ( .A(n1599), .B(n1595), .Z(n1604) );
  XOR U1742 ( .A(n1603), .B(sreg[247]), .Z(n1598) );
  XOR U1743 ( .A(n1604), .B(n1598), .Z(c[247]) );
  ANDN U1744 ( .B(a[122]), .A(n1634), .Z(n1606) );
  AND U1745 ( .A(a[121]), .B(b[1]), .Z(n1608) );
  XNOR U1746 ( .A(n1608), .B(n1607), .Z(n1602) );
  XNOR U1747 ( .A(n1606), .B(n1602), .Z(n1611) );
  XOR U1748 ( .A(n1610), .B(sreg[248]), .Z(n1605) );
  XOR U1749 ( .A(n1611), .B(n1605), .Z(c[248]) );
  ANDN U1750 ( .B(a[123]), .A(n1634), .Z(n1613) );
  AND U1751 ( .A(a[122]), .B(b[1]), .Z(n1615) );
  XNOR U1752 ( .A(n1615), .B(n1614), .Z(n1609) );
  XNOR U1753 ( .A(n1613), .B(n1609), .Z(n1618) );
  XOR U1754 ( .A(n1617), .B(sreg[249]), .Z(n1612) );
  XOR U1755 ( .A(n1618), .B(n1612), .Z(c[249]) );
  ANDN U1756 ( .B(a[124]), .A(n1634), .Z(n1620) );
  AND U1757 ( .A(a[123]), .B(b[1]), .Z(n1622) );
  XNOR U1758 ( .A(n1622), .B(n1621), .Z(n1616) );
  XNOR U1759 ( .A(n1620), .B(n1616), .Z(n1625) );
  XOR U1760 ( .A(n1624), .B(sreg[250]), .Z(n1619) );
  XOR U1761 ( .A(n1625), .B(n1619), .Z(c[250]) );
  ANDN U1762 ( .B(a[125]), .A(n1634), .Z(n1627) );
  AND U1763 ( .A(a[124]), .B(b[1]), .Z(n1629) );
  XNOR U1764 ( .A(n1629), .B(n1628), .Z(n1623) );
  XNOR U1765 ( .A(n1627), .B(n1623), .Z(n1632) );
  XOR U1766 ( .A(n1631), .B(sreg[251]), .Z(n1626) );
  XOR U1767 ( .A(n1632), .B(n1626), .Z(c[251]) );
  AND U1768 ( .A(a[125]), .B(b[1]), .Z(n1637) );
  AND U1769 ( .A(a[126]), .B(b[0]), .Z(n1635) );
  XNOR U1770 ( .A(n1635), .B(n1636), .Z(n1630) );
  XOR U1771 ( .A(n1637), .B(n1630), .Z(n1639) );
  XOR U1772 ( .A(n1638), .B(sreg[252]), .Z(n1633) );
  XNOR U1773 ( .A(n1639), .B(n1633), .Z(c[252]) );
  NANDN U1774 ( .A(n748), .B(a[126]), .Z(n1644) );
  NANDN U1775 ( .A(n1634), .B(a[127]), .Z(n1643) );
  XOR U1776 ( .A(n1644), .B(n1643), .Z(n1645) );
  XNOR U1777 ( .A(n1645), .B(n1646), .Z(n1642) );
  XOR U1778 ( .A(n1641), .B(sreg[253]), .Z(n1640) );
  XOR U1779 ( .A(n1642), .B(n1640), .Z(c[253]) );
  AND U1780 ( .A(a[127]), .B(b[1]), .Z(n1650) );
  OR U1781 ( .A(n1644), .B(n1643), .Z(n1648) );
  NANDN U1782 ( .A(n1646), .B(n1645), .Z(n1647) );
  AND U1783 ( .A(n1648), .B(n1647), .Z(n1651) );
  XNOR U1784 ( .A(n1652), .B(n1651), .Z(n1649) );
  XOR U1785 ( .A(n1650), .B(n1649), .Z(c[254]) );
  NANDN U1786 ( .A(n1650), .B(n1649), .Z(n1654) );
  NANDN U1787 ( .A(n1652), .B(n1651), .Z(n1653) );
  AND U1788 ( .A(n1654), .B(n1653), .Z(c[255]) );
endmodule

