
module mult_N64_CC64 ( clk, rst, a, b, c );
  input [63:0] a;
  input [0:0] b;
  output [63:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294;
  wire   [63:1] swire;
  wire   [127:64] sreg;

  DFF \sreg_reg[64]  ( .D(swire[1]), .CLK(clk), .RST(rst), .Q(sreg[64]) );
  DFF \sreg_reg[65]  ( .D(swire[2]), .CLK(clk), .RST(rst), .Q(sreg[65]) );
  DFF \sreg_reg[66]  ( .D(swire[3]), .CLK(clk), .RST(rst), .Q(sreg[66]) );
  DFF \sreg_reg[67]  ( .D(swire[4]), .CLK(clk), .RST(rst), .Q(sreg[67]) );
  DFF \sreg_reg[68]  ( .D(swire[5]), .CLK(clk), .RST(rst), .Q(sreg[68]) );
  DFF \sreg_reg[69]  ( .D(swire[6]), .CLK(clk), .RST(rst), .Q(sreg[69]) );
  DFF \sreg_reg[70]  ( .D(swire[7]), .CLK(clk), .RST(rst), .Q(sreg[70]) );
  DFF \sreg_reg[71]  ( .D(swire[8]), .CLK(clk), .RST(rst), .Q(sreg[71]) );
  DFF \sreg_reg[72]  ( .D(swire[9]), .CLK(clk), .RST(rst), .Q(sreg[72]) );
  DFF \sreg_reg[73]  ( .D(swire[10]), .CLK(clk), .RST(rst), .Q(sreg[73]) );
  DFF \sreg_reg[74]  ( .D(swire[11]), .CLK(clk), .RST(rst), .Q(sreg[74]) );
  DFF \sreg_reg[75]  ( .D(swire[12]), .CLK(clk), .RST(rst), .Q(sreg[75]) );
  DFF \sreg_reg[76]  ( .D(swire[13]), .CLK(clk), .RST(rst), .Q(sreg[76]) );
  DFF \sreg_reg[77]  ( .D(swire[14]), .CLK(clk), .RST(rst), .Q(sreg[77]) );
  DFF \sreg_reg[78]  ( .D(swire[15]), .CLK(clk), .RST(rst), .Q(sreg[78]) );
  DFF \sreg_reg[79]  ( .D(swire[16]), .CLK(clk), .RST(rst), .Q(sreg[79]) );
  DFF \sreg_reg[80]  ( .D(swire[17]), .CLK(clk), .RST(rst), .Q(sreg[80]) );
  DFF \sreg_reg[81]  ( .D(swire[18]), .CLK(clk), .RST(rst), .Q(sreg[81]) );
  DFF \sreg_reg[82]  ( .D(swire[19]), .CLK(clk), .RST(rst), .Q(sreg[82]) );
  DFF \sreg_reg[83]  ( .D(swire[20]), .CLK(clk), .RST(rst), .Q(sreg[83]) );
  DFF \sreg_reg[84]  ( .D(swire[21]), .CLK(clk), .RST(rst), .Q(sreg[84]) );
  DFF \sreg_reg[85]  ( .D(swire[22]), .CLK(clk), .RST(rst), .Q(sreg[85]) );
  DFF \sreg_reg[86]  ( .D(swire[23]), .CLK(clk), .RST(rst), .Q(sreg[86]) );
  DFF \sreg_reg[87]  ( .D(swire[24]), .CLK(clk), .RST(rst), .Q(sreg[87]) );
  DFF \sreg_reg[88]  ( .D(swire[25]), .CLK(clk), .RST(rst), .Q(sreg[88]) );
  DFF \sreg_reg[89]  ( .D(swire[26]), .CLK(clk), .RST(rst), .Q(sreg[89]) );
  DFF \sreg_reg[90]  ( .D(swire[27]), .CLK(clk), .RST(rst), .Q(sreg[90]) );
  DFF \sreg_reg[91]  ( .D(swire[28]), .CLK(clk), .RST(rst), .Q(sreg[91]) );
  DFF \sreg_reg[92]  ( .D(swire[29]), .CLK(clk), .RST(rst), .Q(sreg[92]) );
  DFF \sreg_reg[93]  ( .D(swire[30]), .CLK(clk), .RST(rst), .Q(sreg[93]) );
  DFF \sreg_reg[94]  ( .D(swire[31]), .CLK(clk), .RST(rst), .Q(sreg[94]) );
  DFF \sreg_reg[95]  ( .D(swire[32]), .CLK(clk), .RST(rst), .Q(sreg[95]) );
  DFF \sreg_reg[96]  ( .D(swire[33]), .CLK(clk), .RST(rst), .Q(sreg[96]) );
  DFF \sreg_reg[97]  ( .D(swire[34]), .CLK(clk), .RST(rst), .Q(sreg[97]) );
  DFF \sreg_reg[98]  ( .D(swire[35]), .CLK(clk), .RST(rst), .Q(sreg[98]) );
  DFF \sreg_reg[99]  ( .D(swire[36]), .CLK(clk), .RST(rst), .Q(sreg[99]) );
  DFF \sreg_reg[100]  ( .D(swire[37]), .CLK(clk), .RST(rst), .Q(sreg[100]) );
  DFF \sreg_reg[101]  ( .D(swire[38]), .CLK(clk), .RST(rst), .Q(sreg[101]) );
  DFF \sreg_reg[102]  ( .D(swire[39]), .CLK(clk), .RST(rst), .Q(sreg[102]) );
  DFF \sreg_reg[103]  ( .D(swire[40]), .CLK(clk), .RST(rst), .Q(sreg[103]) );
  DFF \sreg_reg[104]  ( .D(swire[41]), .CLK(clk), .RST(rst), .Q(sreg[104]) );
  DFF \sreg_reg[105]  ( .D(swire[42]), .CLK(clk), .RST(rst), .Q(sreg[105]) );
  DFF \sreg_reg[106]  ( .D(swire[43]), .CLK(clk), .RST(rst), .Q(sreg[106]) );
  DFF \sreg_reg[107]  ( .D(swire[44]), .CLK(clk), .RST(rst), .Q(sreg[107]) );
  DFF \sreg_reg[108]  ( .D(swire[45]), .CLK(clk), .RST(rst), .Q(sreg[108]) );
  DFF \sreg_reg[109]  ( .D(swire[46]), .CLK(clk), .RST(rst), .Q(sreg[109]) );
  DFF \sreg_reg[110]  ( .D(swire[47]), .CLK(clk), .RST(rst), .Q(sreg[110]) );
  DFF \sreg_reg[111]  ( .D(swire[48]), .CLK(clk), .RST(rst), .Q(sreg[111]) );
  DFF \sreg_reg[112]  ( .D(swire[49]), .CLK(clk), .RST(rst), .Q(sreg[112]) );
  DFF \sreg_reg[113]  ( .D(swire[50]), .CLK(clk), .RST(rst), .Q(sreg[113]) );
  DFF \sreg_reg[114]  ( .D(swire[51]), .CLK(clk), .RST(rst), .Q(sreg[114]) );
  DFF \sreg_reg[115]  ( .D(swire[52]), .CLK(clk), .RST(rst), .Q(sreg[115]) );
  DFF \sreg_reg[116]  ( .D(swire[53]), .CLK(clk), .RST(rst), .Q(sreg[116]) );
  DFF \sreg_reg[117]  ( .D(swire[54]), .CLK(clk), .RST(rst), .Q(sreg[117]) );
  DFF \sreg_reg[118]  ( .D(swire[55]), .CLK(clk), .RST(rst), .Q(sreg[118]) );
  DFF \sreg_reg[119]  ( .D(swire[56]), .CLK(clk), .RST(rst), .Q(sreg[119]) );
  DFF \sreg_reg[120]  ( .D(swire[57]), .CLK(clk), .RST(rst), .Q(sreg[120]) );
  DFF \sreg_reg[121]  ( .D(swire[58]), .CLK(clk), .RST(rst), .Q(sreg[121]) );
  DFF \sreg_reg[122]  ( .D(swire[59]), .CLK(clk), .RST(rst), .Q(sreg[122]) );
  DFF \sreg_reg[123]  ( .D(swire[60]), .CLK(clk), .RST(rst), .Q(sreg[123]) );
  DFF \sreg_reg[124]  ( .D(swire[61]), .CLK(clk), .RST(rst), .Q(sreg[124]) );
  DFF \sreg_reg[125]  ( .D(swire[62]), .CLK(clk), .RST(rst), .Q(sreg[125]) );
  DFF \sreg_reg[126]  ( .D(swire[63]), .CLK(clk), .RST(rst), .Q(sreg[126]) );
  DFF \sreg_reg[63]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[62]) );
  DFF \sreg_reg[62]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[61]) );
  DFF \sreg_reg[61]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[60]) );
  DFF \sreg_reg[60]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[59]) );
  DFF \sreg_reg[59]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[58]) );
  DFF \sreg_reg[58]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[57]) );
  DFF \sreg_reg[57]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[56]) );
  DFF \sreg_reg[56]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[55]) );
  DFF \sreg_reg[55]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[54]) );
  DFF \sreg_reg[54]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[53]) );
  DFF \sreg_reg[53]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[52]) );
  DFF \sreg_reg[52]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[51]) );
  DFF \sreg_reg[51]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[50]) );
  DFF \sreg_reg[50]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[49]) );
  DFF \sreg_reg[49]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[48]) );
  DFF \sreg_reg[48]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[47]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[46]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[45]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[44]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[43]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[42]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[41]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[40]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[39]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[38]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[37]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[36]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[35]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[34]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[33]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[32]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[31]  ( .D(c[31]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[30]  ( .D(c[30]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[29]  ( .D(c[29]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[28]  ( .D(c[28]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[27]  ( .D(c[27]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[26]  ( .D(c[26]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[25]  ( .D(c[25]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[24]  ( .D(c[24]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[23]  ( .D(c[23]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[22]  ( .D(c[22]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[21]  ( .D(c[21]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[20]  ( .D(c[20]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[19]  ( .D(c[19]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[18]  ( .D(c[18]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[17]  ( .D(c[17]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[16]  ( .D(c[16]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[15]  ( .D(c[15]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[14]  ( .D(c[14]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[13]  ( .D(c[13]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[12]  ( .D(c[12]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[11]  ( .D(c[11]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[10]  ( .D(c[10]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[9]  ( .D(c[9]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[8]  ( .D(c[8]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[7]  ( .D(c[7]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[6]  ( .D(c[6]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[5]  ( .D(c[5]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[4]  ( .D(c[4]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[3]  ( .D(c[3]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[2]  ( .D(c[2]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[1]  ( .D(c[1]), .CLK(clk), .RST(rst), .Q(c[0]) );
  XNOR U4 ( .A(n33), .B(n30), .Z(n31) );
  XNOR U5 ( .A(n48), .B(n45), .Z(n46) );
  XNOR U6 ( .A(n65), .B(n60), .Z(n61) );
  XNOR U7 ( .A(n80), .B(n77), .Z(n78) );
  XNOR U8 ( .A(n95), .B(n92), .Z(n93) );
  XNOR U9 ( .A(n110), .B(n107), .Z(n108) );
  XNOR U10 ( .A(n127), .B(n124), .Z(n125) );
  XNOR U11 ( .A(n142), .B(n139), .Z(n140) );
  XNOR U12 ( .A(n157), .B(n154), .Z(n155) );
  XNOR U13 ( .A(n174), .B(n171), .Z(n172) );
  XNOR U14 ( .A(n189), .B(n186), .Z(n187) );
  XNOR U15 ( .A(n204), .B(n201), .Z(n202) );
  XNOR U16 ( .A(n221), .B(n216), .Z(n217) );
  XNOR U17 ( .A(n236), .B(n233), .Z(n234) );
  XNOR U18 ( .A(n251), .B(n248), .Z(n249) );
  XNOR U19 ( .A(n266), .B(n263), .Z(n264) );
  XNOR U20 ( .A(n275), .B(n274), .Z(n5) );
  XNOR U21 ( .A(n284), .B(n283), .Z(n63) );
  XNOR U22 ( .A(n38), .B(n35), .Z(n36) );
  XNOR U23 ( .A(n53), .B(n50), .Z(n51) );
  XNOR U24 ( .A(n70), .B(n67), .Z(n68) );
  XNOR U25 ( .A(n85), .B(n82), .Z(n83) );
  XNOR U26 ( .A(n100), .B(n97), .Z(n98) );
  XNOR U27 ( .A(n117), .B(n112), .Z(n113) );
  XNOR U28 ( .A(n132), .B(n129), .Z(n130) );
  XNOR U29 ( .A(n147), .B(n144), .Z(n145) );
  XNOR U30 ( .A(n162), .B(n159), .Z(n160) );
  XNOR U31 ( .A(n179), .B(n176), .Z(n177) );
  XNOR U32 ( .A(n194), .B(n191), .Z(n192) );
  XNOR U33 ( .A(n209), .B(n206), .Z(n207) );
  XNOR U34 ( .A(n226), .B(n223), .Z(n224) );
  XNOR U35 ( .A(n241), .B(n238), .Z(n239) );
  XNOR U36 ( .A(n256), .B(n253), .Z(n254) );
  XNOR U37 ( .A(n269), .B(n268), .Z(n2) );
  XNOR U38 ( .A(n278), .B(n277), .Z(n7) );
  XNOR U39 ( .A(n287), .B(n286), .Z(n115) );
  XNOR U40 ( .A(n28), .B(n25), .Z(n26) );
  XNOR U41 ( .A(n43), .B(n40), .Z(n41) );
  XNOR U42 ( .A(n58), .B(n55), .Z(n56) );
  XNOR U43 ( .A(n75), .B(n72), .Z(n73) );
  XNOR U44 ( .A(n90), .B(n87), .Z(n88) );
  XNOR U45 ( .A(n105), .B(n102), .Z(n103) );
  XNOR U46 ( .A(n122), .B(n119), .Z(n120) );
  XNOR U47 ( .A(n137), .B(n134), .Z(n135) );
  XNOR U48 ( .A(n152), .B(n149), .Z(n150) );
  XNOR U49 ( .A(n169), .B(n164), .Z(n165) );
  XNOR U50 ( .A(n184), .B(n181), .Z(n182) );
  XNOR U51 ( .A(n199), .B(n196), .Z(n197) );
  XNOR U52 ( .A(n214), .B(n211), .Z(n212) );
  XNOR U53 ( .A(n231), .B(n228), .Z(n229) );
  XNOR U54 ( .A(n246), .B(n243), .Z(n244) );
  XNOR U55 ( .A(n261), .B(n258), .Z(n259) );
  XNOR U56 ( .A(n272), .B(n271), .Z(n3) );
  XNOR U57 ( .A(n281), .B(n280), .Z(n12) );
  XOR U58 ( .A(n290), .B(n289), .Z(n167) );
  XNOR U59 ( .A(n1), .B(n2), .Z(swire[9]) );
  XNOR U60 ( .A(n3), .B(n4), .Z(swire[8]) );
  XNOR U61 ( .A(n5), .B(n6), .Z(swire[7]) );
  XNOR U62 ( .A(n7), .B(n8), .Z(swire[6]) );
  AND U63 ( .A(a[63]), .B(b[0]), .Z(swire[63]) );
  XOR U64 ( .A(sreg[126]), .B(n9), .Z(swire[62]) );
  AND U65 ( .A(a[62]), .B(b[0]), .Z(n9) );
  XOR U66 ( .A(sreg[125]), .B(n10), .Z(swire[61]) );
  AND U67 ( .A(a[61]), .B(b[0]), .Z(n10) );
  XOR U68 ( .A(sreg[124]), .B(n11), .Z(swire[60]) );
  AND U69 ( .A(a[60]), .B(b[0]), .Z(n11) );
  XNOR U70 ( .A(n12), .B(n13), .Z(swire[5]) );
  XOR U71 ( .A(sreg[123]), .B(n14), .Z(swire[59]) );
  AND U72 ( .A(a[59]), .B(b[0]), .Z(n14) );
  XOR U73 ( .A(n15), .B(n16), .Z(swire[58]) );
  XNOR U74 ( .A(sreg[122]), .B(n17), .Z(n16) );
  XNOR U75 ( .A(n18), .B(n17), .Z(n15) );
  XNOR U76 ( .A(n19), .B(n20), .Z(n17) );
  ANDN U77 ( .B(n21), .A(n22), .Z(n19) );
  AND U78 ( .A(a[58]), .B(b[0]), .Z(n18) );
  XNOR U79 ( .A(n21), .B(n22), .Z(swire[57]) );
  XNOR U80 ( .A(sreg[121]), .B(n20), .Z(n22) );
  XOR U81 ( .A(n23), .B(n20), .Z(n21) );
  XNOR U82 ( .A(n24), .B(n25), .Z(n20) );
  ANDN U83 ( .B(n26), .A(n27), .Z(n24) );
  AND U84 ( .A(a[57]), .B(b[0]), .Z(n23) );
  XNOR U85 ( .A(n26), .B(n27), .Z(swire[56]) );
  XOR U86 ( .A(sreg[120]), .B(n25), .Z(n27) );
  XOR U87 ( .A(n29), .B(n30), .Z(n25) );
  ANDN U88 ( .B(n31), .A(n32), .Z(n29) );
  AND U89 ( .A(a[56]), .B(b[0]), .Z(n28) );
  XNOR U90 ( .A(n31), .B(n32), .Z(swire[55]) );
  XOR U91 ( .A(sreg[119]), .B(n30), .Z(n32) );
  XOR U92 ( .A(n34), .B(n35), .Z(n30) );
  ANDN U93 ( .B(n36), .A(n37), .Z(n34) );
  AND U94 ( .A(a[55]), .B(b[0]), .Z(n33) );
  XNOR U95 ( .A(n36), .B(n37), .Z(swire[54]) );
  XOR U96 ( .A(sreg[118]), .B(n35), .Z(n37) );
  XOR U97 ( .A(n39), .B(n40), .Z(n35) );
  ANDN U98 ( .B(n41), .A(n42), .Z(n39) );
  AND U99 ( .A(a[54]), .B(b[0]), .Z(n38) );
  XNOR U100 ( .A(n41), .B(n42), .Z(swire[53]) );
  XOR U101 ( .A(sreg[117]), .B(n40), .Z(n42) );
  XOR U102 ( .A(n44), .B(n45), .Z(n40) );
  ANDN U103 ( .B(n46), .A(n47), .Z(n44) );
  AND U104 ( .A(a[53]), .B(b[0]), .Z(n43) );
  XNOR U105 ( .A(n46), .B(n47), .Z(swire[52]) );
  XOR U106 ( .A(sreg[116]), .B(n45), .Z(n47) );
  XOR U107 ( .A(n49), .B(n50), .Z(n45) );
  ANDN U108 ( .B(n51), .A(n52), .Z(n49) );
  AND U109 ( .A(a[52]), .B(b[0]), .Z(n48) );
  XNOR U110 ( .A(n51), .B(n52), .Z(swire[51]) );
  XOR U111 ( .A(sreg[115]), .B(n50), .Z(n52) );
  XOR U112 ( .A(n54), .B(n55), .Z(n50) );
  ANDN U113 ( .B(n56), .A(n57), .Z(n54) );
  AND U114 ( .A(a[51]), .B(b[0]), .Z(n53) );
  XNOR U115 ( .A(n56), .B(n57), .Z(swire[50]) );
  XOR U116 ( .A(sreg[114]), .B(n55), .Z(n57) );
  XOR U117 ( .A(n59), .B(n60), .Z(n55) );
  ANDN U118 ( .B(n61), .A(n62), .Z(n59) );
  AND U119 ( .A(a[50]), .B(b[0]), .Z(n58) );
  XNOR U120 ( .A(n63), .B(n64), .Z(swire[4]) );
  XNOR U121 ( .A(n61), .B(n62), .Z(swire[49]) );
  XOR U122 ( .A(sreg[113]), .B(n60), .Z(n62) );
  XOR U123 ( .A(n66), .B(n67), .Z(n60) );
  ANDN U124 ( .B(n68), .A(n69), .Z(n66) );
  AND U125 ( .A(a[49]), .B(b[0]), .Z(n65) );
  XNOR U126 ( .A(n68), .B(n69), .Z(swire[48]) );
  XOR U127 ( .A(sreg[112]), .B(n67), .Z(n69) );
  XOR U128 ( .A(n71), .B(n72), .Z(n67) );
  ANDN U129 ( .B(n73), .A(n74), .Z(n71) );
  AND U130 ( .A(a[48]), .B(b[0]), .Z(n70) );
  XNOR U131 ( .A(n73), .B(n74), .Z(swire[47]) );
  XOR U132 ( .A(sreg[111]), .B(n72), .Z(n74) );
  XOR U133 ( .A(n76), .B(n77), .Z(n72) );
  ANDN U134 ( .B(n78), .A(n79), .Z(n76) );
  AND U135 ( .A(a[47]), .B(b[0]), .Z(n75) );
  XNOR U136 ( .A(n78), .B(n79), .Z(swire[46]) );
  XOR U137 ( .A(sreg[110]), .B(n77), .Z(n79) );
  XOR U138 ( .A(n81), .B(n82), .Z(n77) );
  ANDN U139 ( .B(n83), .A(n84), .Z(n81) );
  AND U140 ( .A(a[46]), .B(b[0]), .Z(n80) );
  XNOR U141 ( .A(n83), .B(n84), .Z(swire[45]) );
  XOR U142 ( .A(sreg[109]), .B(n82), .Z(n84) );
  XOR U143 ( .A(n86), .B(n87), .Z(n82) );
  ANDN U144 ( .B(n88), .A(n89), .Z(n86) );
  AND U145 ( .A(a[45]), .B(b[0]), .Z(n85) );
  XNOR U146 ( .A(n88), .B(n89), .Z(swire[44]) );
  XOR U147 ( .A(sreg[108]), .B(n87), .Z(n89) );
  XOR U148 ( .A(n91), .B(n92), .Z(n87) );
  ANDN U149 ( .B(n93), .A(n94), .Z(n91) );
  AND U150 ( .A(a[44]), .B(b[0]), .Z(n90) );
  XNOR U151 ( .A(n93), .B(n94), .Z(swire[43]) );
  XOR U152 ( .A(sreg[107]), .B(n92), .Z(n94) );
  XOR U153 ( .A(n96), .B(n97), .Z(n92) );
  ANDN U154 ( .B(n98), .A(n99), .Z(n96) );
  AND U155 ( .A(a[43]), .B(b[0]), .Z(n95) );
  XNOR U156 ( .A(n98), .B(n99), .Z(swire[42]) );
  XOR U157 ( .A(sreg[106]), .B(n97), .Z(n99) );
  XOR U158 ( .A(n101), .B(n102), .Z(n97) );
  ANDN U159 ( .B(n103), .A(n104), .Z(n101) );
  AND U160 ( .A(a[42]), .B(b[0]), .Z(n100) );
  XNOR U161 ( .A(n103), .B(n104), .Z(swire[41]) );
  XOR U162 ( .A(sreg[105]), .B(n102), .Z(n104) );
  XOR U163 ( .A(n106), .B(n107), .Z(n102) );
  ANDN U164 ( .B(n108), .A(n109), .Z(n106) );
  AND U165 ( .A(a[41]), .B(b[0]), .Z(n105) );
  XNOR U166 ( .A(n108), .B(n109), .Z(swire[40]) );
  XOR U167 ( .A(sreg[104]), .B(n107), .Z(n109) );
  XOR U168 ( .A(n111), .B(n112), .Z(n107) );
  ANDN U169 ( .B(n113), .A(n114), .Z(n111) );
  AND U170 ( .A(a[40]), .B(b[0]), .Z(n110) );
  XNOR U171 ( .A(n115), .B(n116), .Z(swire[3]) );
  XNOR U172 ( .A(n113), .B(n114), .Z(swire[39]) );
  XOR U173 ( .A(sreg[103]), .B(n112), .Z(n114) );
  XOR U174 ( .A(n118), .B(n119), .Z(n112) );
  ANDN U175 ( .B(n120), .A(n121), .Z(n118) );
  AND U176 ( .A(a[39]), .B(b[0]), .Z(n117) );
  XNOR U177 ( .A(n120), .B(n121), .Z(swire[38]) );
  XOR U178 ( .A(sreg[102]), .B(n119), .Z(n121) );
  XOR U179 ( .A(n123), .B(n124), .Z(n119) );
  ANDN U180 ( .B(n125), .A(n126), .Z(n123) );
  AND U181 ( .A(a[38]), .B(b[0]), .Z(n122) );
  XNOR U182 ( .A(n125), .B(n126), .Z(swire[37]) );
  XOR U183 ( .A(sreg[101]), .B(n124), .Z(n126) );
  XOR U184 ( .A(n128), .B(n129), .Z(n124) );
  ANDN U185 ( .B(n130), .A(n131), .Z(n128) );
  AND U186 ( .A(a[37]), .B(b[0]), .Z(n127) );
  XNOR U187 ( .A(n130), .B(n131), .Z(swire[36]) );
  XOR U188 ( .A(sreg[100]), .B(n129), .Z(n131) );
  XOR U189 ( .A(n133), .B(n134), .Z(n129) );
  ANDN U190 ( .B(n135), .A(n136), .Z(n133) );
  AND U191 ( .A(a[36]), .B(b[0]), .Z(n132) );
  XNOR U192 ( .A(n135), .B(n136), .Z(swire[35]) );
  XOR U193 ( .A(sreg[99]), .B(n134), .Z(n136) );
  XOR U194 ( .A(n138), .B(n139), .Z(n134) );
  ANDN U195 ( .B(n140), .A(n141), .Z(n138) );
  AND U196 ( .A(a[35]), .B(b[0]), .Z(n137) );
  XNOR U197 ( .A(n140), .B(n141), .Z(swire[34]) );
  XOR U198 ( .A(sreg[98]), .B(n139), .Z(n141) );
  XOR U199 ( .A(n143), .B(n144), .Z(n139) );
  ANDN U200 ( .B(n145), .A(n146), .Z(n143) );
  AND U201 ( .A(a[34]), .B(b[0]), .Z(n142) );
  XNOR U202 ( .A(n145), .B(n146), .Z(swire[33]) );
  XOR U203 ( .A(sreg[97]), .B(n144), .Z(n146) );
  XOR U204 ( .A(n148), .B(n149), .Z(n144) );
  ANDN U205 ( .B(n150), .A(n151), .Z(n148) );
  AND U206 ( .A(a[33]), .B(b[0]), .Z(n147) );
  XNOR U207 ( .A(n150), .B(n151), .Z(swire[32]) );
  XOR U208 ( .A(sreg[96]), .B(n149), .Z(n151) );
  XOR U209 ( .A(n153), .B(n154), .Z(n149) );
  ANDN U210 ( .B(n155), .A(n156), .Z(n153) );
  AND U211 ( .A(a[32]), .B(b[0]), .Z(n152) );
  XNOR U212 ( .A(n155), .B(n156), .Z(swire[31]) );
  XOR U213 ( .A(sreg[95]), .B(n154), .Z(n156) );
  XOR U214 ( .A(n158), .B(n159), .Z(n154) );
  ANDN U215 ( .B(n160), .A(n161), .Z(n158) );
  AND U216 ( .A(a[31]), .B(b[0]), .Z(n157) );
  XNOR U217 ( .A(n160), .B(n161), .Z(swire[30]) );
  XOR U218 ( .A(sreg[94]), .B(n159), .Z(n161) );
  XOR U219 ( .A(n163), .B(n164), .Z(n159) );
  ANDN U220 ( .B(n165), .A(n166), .Z(n163) );
  AND U221 ( .A(a[30]), .B(b[0]), .Z(n162) );
  XOR U222 ( .A(n167), .B(n168), .Z(swire[2]) );
  XNOR U223 ( .A(n165), .B(n166), .Z(swire[29]) );
  XOR U224 ( .A(sreg[93]), .B(n164), .Z(n166) );
  XOR U225 ( .A(n170), .B(n171), .Z(n164) );
  ANDN U226 ( .B(n172), .A(n173), .Z(n170) );
  AND U227 ( .A(a[29]), .B(b[0]), .Z(n169) );
  XNOR U228 ( .A(n172), .B(n173), .Z(swire[28]) );
  XOR U229 ( .A(sreg[92]), .B(n171), .Z(n173) );
  XOR U230 ( .A(n175), .B(n176), .Z(n171) );
  ANDN U231 ( .B(n177), .A(n178), .Z(n175) );
  AND U232 ( .A(a[28]), .B(b[0]), .Z(n174) );
  XNOR U233 ( .A(n177), .B(n178), .Z(swire[27]) );
  XOR U234 ( .A(sreg[91]), .B(n176), .Z(n178) );
  XOR U235 ( .A(n180), .B(n181), .Z(n176) );
  ANDN U236 ( .B(n182), .A(n183), .Z(n180) );
  AND U237 ( .A(a[27]), .B(b[0]), .Z(n179) );
  XNOR U238 ( .A(n182), .B(n183), .Z(swire[26]) );
  XOR U239 ( .A(sreg[90]), .B(n181), .Z(n183) );
  XOR U240 ( .A(n185), .B(n186), .Z(n181) );
  ANDN U241 ( .B(n187), .A(n188), .Z(n185) );
  AND U242 ( .A(a[26]), .B(b[0]), .Z(n184) );
  XNOR U243 ( .A(n187), .B(n188), .Z(swire[25]) );
  XOR U244 ( .A(sreg[89]), .B(n186), .Z(n188) );
  XOR U245 ( .A(n190), .B(n191), .Z(n186) );
  ANDN U246 ( .B(n192), .A(n193), .Z(n190) );
  AND U247 ( .A(a[25]), .B(b[0]), .Z(n189) );
  XNOR U248 ( .A(n192), .B(n193), .Z(swire[24]) );
  XOR U249 ( .A(sreg[88]), .B(n191), .Z(n193) );
  XOR U250 ( .A(n195), .B(n196), .Z(n191) );
  ANDN U251 ( .B(n197), .A(n198), .Z(n195) );
  AND U252 ( .A(a[24]), .B(b[0]), .Z(n194) );
  XNOR U253 ( .A(n197), .B(n198), .Z(swire[23]) );
  XOR U254 ( .A(sreg[87]), .B(n196), .Z(n198) );
  XOR U255 ( .A(n200), .B(n201), .Z(n196) );
  ANDN U256 ( .B(n202), .A(n203), .Z(n200) );
  AND U257 ( .A(a[23]), .B(b[0]), .Z(n199) );
  XNOR U258 ( .A(n202), .B(n203), .Z(swire[22]) );
  XOR U259 ( .A(sreg[86]), .B(n201), .Z(n203) );
  XOR U260 ( .A(n205), .B(n206), .Z(n201) );
  ANDN U261 ( .B(n207), .A(n208), .Z(n205) );
  AND U262 ( .A(a[22]), .B(b[0]), .Z(n204) );
  XNOR U263 ( .A(n207), .B(n208), .Z(swire[21]) );
  XOR U264 ( .A(sreg[85]), .B(n206), .Z(n208) );
  XOR U265 ( .A(n210), .B(n211), .Z(n206) );
  ANDN U266 ( .B(n212), .A(n213), .Z(n210) );
  AND U267 ( .A(a[21]), .B(b[0]), .Z(n209) );
  XNOR U268 ( .A(n212), .B(n213), .Z(swire[20]) );
  XOR U269 ( .A(sreg[84]), .B(n211), .Z(n213) );
  XOR U270 ( .A(n215), .B(n216), .Z(n211) );
  ANDN U271 ( .B(n217), .A(n218), .Z(n215) );
  AND U272 ( .A(a[20]), .B(b[0]), .Z(n214) );
  XOR U273 ( .A(n219), .B(n220), .Z(swire[1]) );
  XNOR U274 ( .A(n217), .B(n218), .Z(swire[19]) );
  XOR U275 ( .A(sreg[83]), .B(n216), .Z(n218) );
  XOR U276 ( .A(n222), .B(n223), .Z(n216) );
  ANDN U277 ( .B(n224), .A(n225), .Z(n222) );
  AND U278 ( .A(a[19]), .B(b[0]), .Z(n221) );
  XNOR U279 ( .A(n224), .B(n225), .Z(swire[18]) );
  XOR U280 ( .A(sreg[82]), .B(n223), .Z(n225) );
  XOR U281 ( .A(n227), .B(n228), .Z(n223) );
  ANDN U282 ( .B(n229), .A(n230), .Z(n227) );
  AND U283 ( .A(a[18]), .B(b[0]), .Z(n226) );
  XNOR U284 ( .A(n229), .B(n230), .Z(swire[17]) );
  XOR U285 ( .A(sreg[81]), .B(n228), .Z(n230) );
  XOR U286 ( .A(n232), .B(n233), .Z(n228) );
  ANDN U287 ( .B(n234), .A(n235), .Z(n232) );
  AND U288 ( .A(a[17]), .B(b[0]), .Z(n231) );
  XNOR U289 ( .A(n234), .B(n235), .Z(swire[16]) );
  XOR U290 ( .A(sreg[80]), .B(n233), .Z(n235) );
  XOR U291 ( .A(n237), .B(n238), .Z(n233) );
  ANDN U292 ( .B(n239), .A(n240), .Z(n237) );
  AND U293 ( .A(a[16]), .B(b[0]), .Z(n236) );
  XNOR U294 ( .A(n239), .B(n240), .Z(swire[15]) );
  XOR U295 ( .A(sreg[79]), .B(n238), .Z(n240) );
  XOR U296 ( .A(n242), .B(n243), .Z(n238) );
  ANDN U297 ( .B(n244), .A(n245), .Z(n242) );
  AND U298 ( .A(a[15]), .B(b[0]), .Z(n241) );
  XNOR U299 ( .A(n244), .B(n245), .Z(swire[14]) );
  XOR U300 ( .A(sreg[78]), .B(n243), .Z(n245) );
  XOR U301 ( .A(n247), .B(n248), .Z(n243) );
  ANDN U302 ( .B(n249), .A(n250), .Z(n247) );
  AND U303 ( .A(a[14]), .B(b[0]), .Z(n246) );
  XNOR U304 ( .A(n249), .B(n250), .Z(swire[13]) );
  XOR U305 ( .A(sreg[77]), .B(n248), .Z(n250) );
  XOR U306 ( .A(n252), .B(n253), .Z(n248) );
  ANDN U307 ( .B(n254), .A(n255), .Z(n252) );
  AND U308 ( .A(a[13]), .B(b[0]), .Z(n251) );
  XNOR U309 ( .A(n254), .B(n255), .Z(swire[12]) );
  XOR U310 ( .A(sreg[76]), .B(n253), .Z(n255) );
  XOR U311 ( .A(n257), .B(n258), .Z(n253) );
  ANDN U312 ( .B(n259), .A(n260), .Z(n257) );
  AND U313 ( .A(a[12]), .B(b[0]), .Z(n256) );
  XNOR U314 ( .A(n259), .B(n260), .Z(swire[11]) );
  XOR U315 ( .A(sreg[75]), .B(n258), .Z(n260) );
  XOR U316 ( .A(n262), .B(n263), .Z(n258) );
  ANDN U317 ( .B(n264), .A(n265), .Z(n262) );
  AND U318 ( .A(a[11]), .B(b[0]), .Z(n261) );
  XNOR U319 ( .A(n264), .B(n265), .Z(swire[10]) );
  XOR U320 ( .A(sreg[74]), .B(n263), .Z(n265) );
  XOR U321 ( .A(n267), .B(n268), .Z(n263) );
  ANDN U322 ( .B(n2), .A(n1), .Z(n267) );
  XOR U323 ( .A(sreg[73]), .B(n268), .Z(n1) );
  XOR U324 ( .A(n270), .B(n271), .Z(n268) );
  ANDN U325 ( .B(n3), .A(n4), .Z(n270) );
  XOR U326 ( .A(sreg[72]), .B(n271), .Z(n4) );
  XOR U327 ( .A(n273), .B(n274), .Z(n271) );
  ANDN U328 ( .B(n5), .A(n6), .Z(n273) );
  XOR U329 ( .A(sreg[71]), .B(n274), .Z(n6) );
  XOR U330 ( .A(n276), .B(n277), .Z(n274) );
  ANDN U331 ( .B(n7), .A(n8), .Z(n276) );
  XOR U332 ( .A(sreg[70]), .B(n277), .Z(n8) );
  XOR U333 ( .A(n279), .B(n280), .Z(n277) );
  ANDN U334 ( .B(n12), .A(n13), .Z(n279) );
  XOR U335 ( .A(sreg[69]), .B(n280), .Z(n13) );
  XOR U336 ( .A(n282), .B(n283), .Z(n280) );
  ANDN U337 ( .B(n63), .A(n64), .Z(n282) );
  XOR U338 ( .A(sreg[68]), .B(n283), .Z(n64) );
  XOR U339 ( .A(n285), .B(n286), .Z(n283) );
  ANDN U340 ( .B(n115), .A(n116), .Z(n285) );
  XOR U341 ( .A(sreg[67]), .B(n286), .Z(n116) );
  XOR U342 ( .A(n288), .B(n289), .Z(n286) );
  NOR U343 ( .A(n168), .B(n167), .Z(n288) );
  AND U344 ( .A(a[2]), .B(b[0]), .Z(n290) );
  XOR U345 ( .A(sreg[66]), .B(n289), .Z(n168) );
  XOR U346 ( .A(n291), .B(n292), .Z(n289) );
  NAND U347 ( .A(n219), .B(n220), .Z(n292) );
  XOR U348 ( .A(sreg[65]), .B(n291), .Z(n220) );
  XNOR U349 ( .A(n291), .B(n293), .Z(n219) );
  NAND U350 ( .A(b[0]), .B(a[1]), .Z(n293) );
  ANDN U351 ( .B(sreg[64]), .A(n294), .Z(n291) );
  AND U352 ( .A(a[3]), .B(b[0]), .Z(n287) );
  AND U353 ( .A(a[4]), .B(b[0]), .Z(n284) );
  AND U354 ( .A(a[5]), .B(b[0]), .Z(n281) );
  AND U355 ( .A(a[6]), .B(b[0]), .Z(n278) );
  AND U356 ( .A(a[7]), .B(b[0]), .Z(n275) );
  AND U357 ( .A(a[8]), .B(b[0]), .Z(n272) );
  AND U358 ( .A(a[9]), .B(b[0]), .Z(n269) );
  AND U359 ( .A(a[10]), .B(b[0]), .Z(n266) );
  XNOR U360 ( .A(sreg[64]), .B(n294), .Z(c[63]) );
  NAND U361 ( .A(a[0]), .B(b[0]), .Z(n294) );
endmodule

