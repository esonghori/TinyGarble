
module hamming_N16000_CC640_DW01_add_0 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29;

  XOR U1 ( .A(A[9]), .B(n1), .Z(SUM[9]) );
  XOR U2 ( .A(A[8]), .B(n2), .Z(SUM[8]) );
  XNOR U3 ( .A(A[7]), .B(n3), .Z(SUM[7]) );
  XOR U4 ( .A(A[6]), .B(n4), .Z(SUM[6]) );
  XNOR U5 ( .A(A[5]), .B(n5), .Z(SUM[5]) );
  XOR U6 ( .A(n6), .B(n7), .Z(SUM[4]) );
  XNOR U7 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR U8 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U9 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR U10 ( .A(n10), .B(n11), .Z(SUM[2]) );
  XNOR U11 ( .A(B[2]), .B(A[2]), .Z(n11) );
  XOR U12 ( .A(n12), .B(n13), .Z(SUM[1]) );
  XOR U13 ( .A(B[1]), .B(A[1]), .Z(n13) );
  XOR U14 ( .A(A[13]), .B(n14), .Z(SUM[13]) );
  ANDN U15 ( .B(A[12]), .A(n15), .Z(n14) );
  XNOR U16 ( .A(A[12]), .B(n15), .Z(SUM[12]) );
  NANDN U17 ( .A(n16), .B(A[11]), .Z(n15) );
  XNOR U18 ( .A(A[11]), .B(n16), .Z(SUM[11]) );
  NAND U19 ( .A(n17), .B(A[10]), .Z(n16) );
  XOR U20 ( .A(A[10]), .B(n17), .Z(SUM[10]) );
  AND U21 ( .A(A[9]), .B(n1), .Z(n17) );
  AND U22 ( .A(n2), .B(A[8]), .Z(n1) );
  ANDN U23 ( .B(A[7]), .A(n3), .Z(n2) );
  NAND U24 ( .A(n4), .B(A[6]), .Z(n3) );
  ANDN U25 ( .B(A[5]), .A(n5), .Z(n4) );
  AND U26 ( .A(n18), .B(n19), .Z(n5) );
  NAND U27 ( .A(n20), .B(B[4]), .Z(n19) );
  NANDN U28 ( .A(A[4]), .B(n6), .Z(n20) );
  NANDN U29 ( .A(n6), .B(A[4]), .Z(n18) );
  AND U30 ( .A(n21), .B(n22), .Z(n6) );
  NAND U31 ( .A(n23), .B(B[3]), .Z(n22) );
  NANDN U32 ( .A(A[3]), .B(n8), .Z(n23) );
  NANDN U33 ( .A(n8), .B(A[3]), .Z(n21) );
  AND U34 ( .A(n24), .B(n25), .Z(n8) );
  NAND U35 ( .A(n26), .B(B[2]), .Z(n25) );
  NANDN U36 ( .A(A[2]), .B(n10), .Z(n26) );
  NANDN U37 ( .A(n10), .B(A[2]), .Z(n24) );
  AND U38 ( .A(n27), .B(n28), .Z(n10) );
  NAND U39 ( .A(n29), .B(B[1]), .Z(n28) );
  OR U40 ( .A(n12), .B(A[1]), .Z(n29) );
  NAND U41 ( .A(n12), .B(A[1]), .Z(n27) );
  AND U42 ( .A(B[0]), .B(A[0]), .Z(n12) );
  XOR U43 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC640 ( clk, rst, x, y, o );
  input [24:0] x;
  input [24:0] y;
  output [13:0] o;
  input clk, rst;
  wire   n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190;
  wire   [4:0] olocal;
  wire   [13:0] oglobal;

  DFF \oglobal_reg[0]  ( .D(o[0]), .CLK(clk), .RST(rst), .Q(oglobal[0]) );
  DFF \oglobal_reg[1]  ( .D(o[1]), .CLK(clk), .RST(rst), .Q(oglobal[1]) );
  DFF \oglobal_reg[2]  ( .D(o[2]), .CLK(clk), .RST(rst), .Q(oglobal[2]) );
  DFF \oglobal_reg[3]  ( .D(o[3]), .CLK(clk), .RST(rst), .Q(oglobal[3]) );
  DFF \oglobal_reg[4]  ( .D(o[4]), .CLK(clk), .RST(rst), .Q(oglobal[4]) );
  DFF \oglobal_reg[5]  ( .D(o[5]), .CLK(clk), .RST(rst), .Q(oglobal[5]) );
  DFF \oglobal_reg[6]  ( .D(o[6]), .CLK(clk), .RST(rst), .Q(oglobal[6]) );
  DFF \oglobal_reg[7]  ( .D(o[7]), .CLK(clk), .RST(rst), .Q(oglobal[7]) );
  DFF \oglobal_reg[8]  ( .D(o[8]), .CLK(clk), .RST(rst), .Q(oglobal[8]) );
  DFF \oglobal_reg[9]  ( .D(o[9]), .CLK(clk), .RST(rst), .Q(oglobal[9]) );
  DFF \oglobal_reg[10]  ( .D(o[10]), .CLK(clk), .RST(rst), .Q(oglobal[10]) );
  DFF \oglobal_reg[11]  ( .D(o[11]), .CLK(clk), .RST(rst), .Q(oglobal[11]) );
  DFF \oglobal_reg[12]  ( .D(o[12]), .CLK(clk), .RST(rst), .Q(oglobal[12]) );
  DFF \oglobal_reg[13]  ( .D(o[13]), .CLK(clk), .RST(rst), .Q(oglobal[13]) );
  hamming_N16000_CC640_DW01_add_0 add_97 ( .A(oglobal), .B({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, olocal}), .CI(1'b0), .SUM(o) );
  NAND U61 ( .A(n37), .B(n38), .Z(olocal[4]) );
  NANDN U62 ( .A(n39), .B(n40), .Z(n38) );
  OR U63 ( .A(n41), .B(n42), .Z(n40) );
  NAND U64 ( .A(n41), .B(n42), .Z(n37) );
  XOR U65 ( .A(n41), .B(n43), .Z(olocal[3]) );
  XNOR U66 ( .A(n39), .B(n42), .Z(n43) );
  AND U67 ( .A(n44), .B(n45), .Z(n42) );
  NANDN U68 ( .A(n46), .B(n47), .Z(n45) );
  NANDN U69 ( .A(n48), .B(n49), .Z(n47) );
  NANDN U70 ( .A(n49), .B(n48), .Z(n44) );
  NAND U71 ( .A(n50), .B(n51), .Z(n39) );
  NANDN U72 ( .A(n52), .B(n53), .Z(n51) );
  OR U73 ( .A(n54), .B(n55), .Z(n53) );
  NAND U74 ( .A(n55), .B(n54), .Z(n50) );
  AND U75 ( .A(n56), .B(n57), .Z(n41) );
  NANDN U76 ( .A(n58), .B(n59), .Z(n57) );
  NANDN U77 ( .A(n60), .B(n61), .Z(n59) );
  NANDN U78 ( .A(n61), .B(n60), .Z(n56) );
  XOR U79 ( .A(n55), .B(n62), .Z(olocal[2]) );
  XOR U80 ( .A(n52), .B(n54), .Z(n62) );
  XNOR U81 ( .A(n48), .B(n63), .Z(n54) );
  XNOR U82 ( .A(n46), .B(n49), .Z(n63) );
  NAND U83 ( .A(n64), .B(n65), .Z(n49) );
  NAND U84 ( .A(n66), .B(n67), .Z(n65) );
  NANDN U85 ( .A(n68), .B(n69), .Z(n66) );
  NAND U86 ( .A(n70), .B(n68), .Z(n64) );
  IV U87 ( .A(n69), .Z(n70) );
  NAND U88 ( .A(n71), .B(n72), .Z(n46) );
  NAND U89 ( .A(n73), .B(n74), .Z(n72) );
  NANDN U90 ( .A(n75), .B(n76), .Z(n73) );
  NANDN U91 ( .A(n76), .B(n75), .Z(n71) );
  AND U92 ( .A(n77), .B(n78), .Z(n48) );
  NAND U93 ( .A(n79), .B(n80), .Z(n78) );
  NANDN U94 ( .A(n81), .B(n82), .Z(n79) );
  NAND U95 ( .A(n83), .B(n81), .Z(n77) );
  NAND U96 ( .A(n84), .B(n85), .Z(n52) );
  NANDN U97 ( .A(n86), .B(n87), .Z(n85) );
  OR U98 ( .A(n88), .B(n89), .Z(n87) );
  NAND U99 ( .A(n89), .B(n88), .Z(n84) );
  XNOR U100 ( .A(n60), .B(n90), .Z(n55) );
  XNOR U101 ( .A(n58), .B(n61), .Z(n90) );
  NAND U102 ( .A(n91), .B(n92), .Z(n61) );
  NAND U103 ( .A(n93), .B(n94), .Z(n92) );
  NANDN U104 ( .A(n95), .B(n96), .Z(n93) );
  NAND U105 ( .A(n97), .B(n95), .Z(n91) );
  IV U106 ( .A(n96), .Z(n97) );
  NAND U107 ( .A(n98), .B(n99), .Z(n58) );
  NAND U108 ( .A(n100), .B(n101), .Z(n99) );
  NANDN U109 ( .A(n102), .B(n103), .Z(n100) );
  NAND U110 ( .A(n104), .B(n102), .Z(n98) );
  IV U111 ( .A(n103), .Z(n104) );
  AND U112 ( .A(n105), .B(n106), .Z(n60) );
  NAND U113 ( .A(n107), .B(n108), .Z(n106) );
  NANDN U114 ( .A(n109), .B(n110), .Z(n105) );
  XNOR U115 ( .A(n86), .B(n111), .Z(olocal[1]) );
  XOR U116 ( .A(n88), .B(n89), .Z(n111) );
  XOR U117 ( .A(n101), .B(n112), .Z(n89) );
  XNOR U118 ( .A(n102), .B(n103), .Z(n112) );
  XNOR U119 ( .A(n107), .B(n108), .Z(n103) );
  XNOR U120 ( .A(n110), .B(n109), .Z(n108) );
  AND U121 ( .A(n113), .B(n114), .Z(n109) );
  NANDN U122 ( .A(n115), .B(n116), .Z(n114) );
  NANDN U123 ( .A(n117), .B(n118), .Z(n113) );
  IV U124 ( .A(n119), .Z(n118) );
  NAND U125 ( .A(n120), .B(n121), .Z(n110) );
  NANDN U126 ( .A(n122), .B(n123), .Z(n121) );
  NANDN U127 ( .A(n124), .B(n125), .Z(n120) );
  IV U128 ( .A(n126), .Z(n125) );
  NAND U129 ( .A(n127), .B(n128), .Z(n107) );
  NAND U130 ( .A(n129), .B(n130), .Z(n128) );
  NANDN U131 ( .A(n131), .B(n132), .Z(n127) );
  IV U132 ( .A(n133), .Z(n132) );
  NOR U133 ( .A(n134), .B(n135), .Z(n102) );
  IV U134 ( .A(n136), .Z(n134) );
  XNOR U135 ( .A(n95), .B(n137), .Z(n101) );
  XOR U136 ( .A(n94), .B(n96), .Z(n137) );
  AND U137 ( .A(n138), .B(n139), .Z(n96) );
  NANDN U138 ( .A(n140), .B(n141), .Z(n139) );
  IV U139 ( .A(n142), .Z(n141) );
  OR U140 ( .A(n143), .B(n144), .Z(n138) );
  NAND U141 ( .A(n145), .B(n146), .Z(n94) );
  OR U142 ( .A(n147), .B(n148), .Z(n146) );
  OR U143 ( .A(n149), .B(n150), .Z(n145) );
  ANDN U144 ( .B(n151), .A(n152), .Z(n95) );
  IV U145 ( .A(n153), .Z(n152) );
  ANDN U146 ( .B(n154), .A(n155), .Z(n88) );
  XOR U147 ( .A(n74), .B(n156), .Z(n86) );
  XOR U148 ( .A(n75), .B(n76), .Z(n156) );
  XOR U149 ( .A(n81), .B(n157), .Z(n76) );
  XNOR U150 ( .A(n80), .B(n83), .Z(n157) );
  IV U151 ( .A(n82), .Z(n83) );
  AND U152 ( .A(n158), .B(n159), .Z(n82) );
  OR U153 ( .A(n160), .B(n161), .Z(n159) );
  OR U154 ( .A(n162), .B(n163), .Z(n158) );
  NAND U155 ( .A(n164), .B(n165), .Z(n80) );
  OR U156 ( .A(n166), .B(n167), .Z(n165) );
  OR U157 ( .A(n168), .B(n169), .Z(n164) );
  NOR U158 ( .A(n170), .B(n171), .Z(n81) );
  NOR U159 ( .A(n172), .B(n173), .Z(n75) );
  IV U160 ( .A(n174), .Z(n172) );
  XNOR U161 ( .A(n68), .B(n175), .Z(n74) );
  XOR U162 ( .A(n67), .B(n69), .Z(n175) );
  AND U163 ( .A(n176), .B(n177), .Z(n69) );
  OR U164 ( .A(n178), .B(n179), .Z(n177) );
  OR U165 ( .A(n180), .B(n181), .Z(n176) );
  NAND U166 ( .A(n182), .B(n183), .Z(n67) );
  OR U167 ( .A(n184), .B(n185), .Z(n183) );
  OR U168 ( .A(n186), .B(n187), .Z(n182) );
  NOR U169 ( .A(n188), .B(n189), .Z(n68) );
  IV U170 ( .A(n190), .Z(n188) );
  XNOR U171 ( .A(n155), .B(n154), .Z(olocal[0]) );
  XNOR U172 ( .A(n174), .B(n173), .Z(n154) );
  XOR U173 ( .A(n189), .B(n190), .Z(n173) );
  XOR U174 ( .A(n184), .B(n185), .Z(n190) );
  XNOR U175 ( .A(n186), .B(n187), .Z(n185) );
  XNOR U176 ( .A(y[22]), .B(x[22]), .Z(n187) );
  XNOR U177 ( .A(y[23]), .B(x[23]), .Z(n186) );
  XNOR U178 ( .A(y[21]), .B(x[21]), .Z(n184) );
  XNOR U179 ( .A(n178), .B(n179), .Z(n189) );
  XNOR U180 ( .A(y[18]), .B(x[18]), .Z(n179) );
  XNOR U181 ( .A(n180), .B(n181), .Z(n178) );
  XNOR U182 ( .A(y[19]), .B(x[19]), .Z(n181) );
  XNOR U183 ( .A(y[20]), .B(x[20]), .Z(n180) );
  XOR U184 ( .A(n171), .B(n170), .Z(n174) );
  XNOR U185 ( .A(n166), .B(n167), .Z(n170) );
  XNOR U186 ( .A(y[15]), .B(x[15]), .Z(n167) );
  XNOR U187 ( .A(n168), .B(n169), .Z(n166) );
  XNOR U188 ( .A(y[16]), .B(x[16]), .Z(n169) );
  XNOR U189 ( .A(y[17]), .B(x[17]), .Z(n168) );
  XNOR U190 ( .A(n160), .B(n161), .Z(n171) );
  XNOR U191 ( .A(y[12]), .B(x[12]), .Z(n161) );
  XNOR U192 ( .A(n162), .B(n163), .Z(n160) );
  XNOR U193 ( .A(y[13]), .B(x[13]), .Z(n163) );
  XNOR U194 ( .A(y[14]), .B(x[14]), .Z(n162) );
  XOR U195 ( .A(n135), .B(n136), .Z(n155) );
  XOR U196 ( .A(n153), .B(n151), .Z(n136) );
  XOR U197 ( .A(n147), .B(n148), .Z(n151) );
  XNOR U198 ( .A(n149), .B(n150), .Z(n148) );
  XNOR U199 ( .A(y[10]), .B(x[10]), .Z(n150) );
  XNOR U200 ( .A(y[11]), .B(x[11]), .Z(n149) );
  XNOR U201 ( .A(y[9]), .B(x[9]), .Z(n147) );
  XOR U202 ( .A(n140), .B(n142), .Z(n153) );
  XNOR U203 ( .A(n143), .B(n144), .Z(n142) );
  XNOR U204 ( .A(y[7]), .B(x[7]), .Z(n144) );
  XNOR U205 ( .A(y[8]), .B(x[8]), .Z(n143) );
  XNOR U206 ( .A(y[6]), .B(x[6]), .Z(n140) );
  XNOR U207 ( .A(n130), .B(n129), .Z(n135) );
  XOR U208 ( .A(y[24]), .B(x[24]), .Z(n129) );
  XOR U209 ( .A(n131), .B(n133), .Z(n130) );
  XOR U210 ( .A(n115), .B(n116), .Z(n133) );
  XOR U211 ( .A(n117), .B(n119), .Z(n116) );
  XNOR U212 ( .A(y[1]), .B(x[1]), .Z(n119) );
  XNOR U213 ( .A(y[2]), .B(x[2]), .Z(n117) );
  XNOR U214 ( .A(y[0]), .B(x[0]), .Z(n115) );
  XOR U215 ( .A(n122), .B(n123), .Z(n131) );
  XOR U216 ( .A(n124), .B(n126), .Z(n123) );
  XNOR U217 ( .A(y[4]), .B(x[4]), .Z(n126) );
  XNOR U218 ( .A(y[5]), .B(x[5]), .Z(n124) );
  XNOR U219 ( .A(y[3]), .B(x[3]), .Z(n122) );
endmodule

