
module modmult_N256_CC1024 ( clk, rst, start, x, y, n, o );
  input [255:0] x;
  input [255:0] y;
  input [255:0] n;
  output [255:0] o;
  input clk, rst, start;


endmodule


module modexp_2N_NN_N256_CC524288 ( clk, rst, m, e, n, c );
  input [255:0] m;
  input [255:0] e;
  input [255:0] n;
  output [255:0] c;
  input clk, rst;
  wire   init, mul_pow, first_one, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206;
  wire   [1023:0] start_in;
  wire   [1023:0] start_reg;
  wire   [255:0] ereg;
  wire   [255:0] o;
  wire   [255:0] creg;
  wire   [255:0] x;
  wire   [255:0] y;

  modmult_N256_CC1024 modmult_1 ( .clk(clk), .rst(rst), .start(start_in[0]), 
        .x(x), .y(y), .n(n), .o(o) );
  DFF init_reg ( .D(1'b1), .CLK(clk), .RST(rst), .Q(init) );
  DFF \start_reg_reg[0]  ( .D(start_in[1023]), .CLK(clk), .RST(rst), .Q(
        start_reg[0]) );
  DFF \start_reg_reg[1]  ( .D(start_in[0]), .CLK(clk), .RST(rst), .Q(
        start_reg[1]) );
  DFF \start_reg_reg[2]  ( .D(start_in[1]), .CLK(clk), .RST(rst), .Q(
        start_reg[2]) );
  DFF \start_reg_reg[3]  ( .D(start_in[2]), .CLK(clk), .RST(rst), .Q(
        start_reg[3]) );
  DFF \start_reg_reg[4]  ( .D(start_in[3]), .CLK(clk), .RST(rst), .Q(
        start_reg[4]) );
  DFF \start_reg_reg[5]  ( .D(start_in[4]), .CLK(clk), .RST(rst), .Q(
        start_reg[5]) );
  DFF \start_reg_reg[6]  ( .D(start_in[5]), .CLK(clk), .RST(rst), .Q(
        start_reg[6]) );
  DFF \start_reg_reg[7]  ( .D(start_in[6]), .CLK(clk), .RST(rst), .Q(
        start_reg[7]) );
  DFF \start_reg_reg[8]  ( .D(start_in[7]), .CLK(clk), .RST(rst), .Q(
        start_reg[8]) );
  DFF \start_reg_reg[9]  ( .D(start_in[8]), .CLK(clk), .RST(rst), .Q(
        start_reg[9]) );
  DFF \start_reg_reg[10]  ( .D(start_in[9]), .CLK(clk), .RST(rst), .Q(
        start_reg[10]) );
  DFF \start_reg_reg[11]  ( .D(start_in[10]), .CLK(clk), .RST(rst), .Q(
        start_reg[11]) );
  DFF \start_reg_reg[12]  ( .D(start_in[11]), .CLK(clk), .RST(rst), .Q(
        start_reg[12]) );
  DFF \start_reg_reg[13]  ( .D(start_in[12]), .CLK(clk), .RST(rst), .Q(
        start_reg[13]) );
  DFF \start_reg_reg[14]  ( .D(start_in[13]), .CLK(clk), .RST(rst), .Q(
        start_reg[14]) );
  DFF \start_reg_reg[15]  ( .D(start_in[14]), .CLK(clk), .RST(rst), .Q(
        start_reg[15]) );
  DFF \start_reg_reg[16]  ( .D(start_in[15]), .CLK(clk), .RST(rst), .Q(
        start_reg[16]) );
  DFF \start_reg_reg[17]  ( .D(start_in[16]), .CLK(clk), .RST(rst), .Q(
        start_reg[17]) );
  DFF \start_reg_reg[18]  ( .D(start_in[17]), .CLK(clk), .RST(rst), .Q(
        start_reg[18]) );
  DFF \start_reg_reg[19]  ( .D(start_in[18]), .CLK(clk), .RST(rst), .Q(
        start_reg[19]) );
  DFF \start_reg_reg[20]  ( .D(start_in[19]), .CLK(clk), .RST(rst), .Q(
        start_reg[20]) );
  DFF \start_reg_reg[21]  ( .D(start_in[20]), .CLK(clk), .RST(rst), .Q(
        start_reg[21]) );
  DFF \start_reg_reg[22]  ( .D(start_in[21]), .CLK(clk), .RST(rst), .Q(
        start_reg[22]) );
  DFF \start_reg_reg[23]  ( .D(start_in[22]), .CLK(clk), .RST(rst), .Q(
        start_reg[23]) );
  DFF \start_reg_reg[24]  ( .D(start_in[23]), .CLK(clk), .RST(rst), .Q(
        start_reg[24]) );
  DFF \start_reg_reg[25]  ( .D(start_in[24]), .CLK(clk), .RST(rst), .Q(
        start_reg[25]) );
  DFF \start_reg_reg[26]  ( .D(start_in[25]), .CLK(clk), .RST(rst), .Q(
        start_reg[26]) );
  DFF \start_reg_reg[27]  ( .D(start_in[26]), .CLK(clk), .RST(rst), .Q(
        start_reg[27]) );
  DFF \start_reg_reg[28]  ( .D(start_in[27]), .CLK(clk), .RST(rst), .Q(
        start_reg[28]) );
  DFF \start_reg_reg[29]  ( .D(start_in[28]), .CLK(clk), .RST(rst), .Q(
        start_reg[29]) );
  DFF \start_reg_reg[30]  ( .D(start_in[29]), .CLK(clk), .RST(rst), .Q(
        start_reg[30]) );
  DFF \start_reg_reg[31]  ( .D(start_in[30]), .CLK(clk), .RST(rst), .Q(
        start_reg[31]) );
  DFF \start_reg_reg[32]  ( .D(start_in[31]), .CLK(clk), .RST(rst), .Q(
        start_reg[32]) );
  DFF \start_reg_reg[33]  ( .D(start_in[32]), .CLK(clk), .RST(rst), .Q(
        start_reg[33]) );
  DFF \start_reg_reg[34]  ( .D(start_in[33]), .CLK(clk), .RST(rst), .Q(
        start_reg[34]) );
  DFF \start_reg_reg[35]  ( .D(start_in[34]), .CLK(clk), .RST(rst), .Q(
        start_reg[35]) );
  DFF \start_reg_reg[36]  ( .D(start_in[35]), .CLK(clk), .RST(rst), .Q(
        start_reg[36]) );
  DFF \start_reg_reg[37]  ( .D(start_in[36]), .CLK(clk), .RST(rst), .Q(
        start_reg[37]) );
  DFF \start_reg_reg[38]  ( .D(start_in[37]), .CLK(clk), .RST(rst), .Q(
        start_reg[38]) );
  DFF \start_reg_reg[39]  ( .D(start_in[38]), .CLK(clk), .RST(rst), .Q(
        start_reg[39]) );
  DFF \start_reg_reg[40]  ( .D(start_in[39]), .CLK(clk), .RST(rst), .Q(
        start_reg[40]) );
  DFF \start_reg_reg[41]  ( .D(start_in[40]), .CLK(clk), .RST(rst), .Q(
        start_reg[41]) );
  DFF \start_reg_reg[42]  ( .D(start_in[41]), .CLK(clk), .RST(rst), .Q(
        start_reg[42]) );
  DFF \start_reg_reg[43]  ( .D(start_in[42]), .CLK(clk), .RST(rst), .Q(
        start_reg[43]) );
  DFF \start_reg_reg[44]  ( .D(start_in[43]), .CLK(clk), .RST(rst), .Q(
        start_reg[44]) );
  DFF \start_reg_reg[45]  ( .D(start_in[44]), .CLK(clk), .RST(rst), .Q(
        start_reg[45]) );
  DFF \start_reg_reg[46]  ( .D(start_in[45]), .CLK(clk), .RST(rst), .Q(
        start_reg[46]) );
  DFF \start_reg_reg[47]  ( .D(start_in[46]), .CLK(clk), .RST(rst), .Q(
        start_reg[47]) );
  DFF \start_reg_reg[48]  ( .D(start_in[47]), .CLK(clk), .RST(rst), .Q(
        start_reg[48]) );
  DFF \start_reg_reg[49]  ( .D(start_in[48]), .CLK(clk), .RST(rst), .Q(
        start_reg[49]) );
  DFF \start_reg_reg[50]  ( .D(start_in[49]), .CLK(clk), .RST(rst), .Q(
        start_reg[50]) );
  DFF \start_reg_reg[51]  ( .D(start_in[50]), .CLK(clk), .RST(rst), .Q(
        start_reg[51]) );
  DFF \start_reg_reg[52]  ( .D(start_in[51]), .CLK(clk), .RST(rst), .Q(
        start_reg[52]) );
  DFF \start_reg_reg[53]  ( .D(start_in[52]), .CLK(clk), .RST(rst), .Q(
        start_reg[53]) );
  DFF \start_reg_reg[54]  ( .D(start_in[53]), .CLK(clk), .RST(rst), .Q(
        start_reg[54]) );
  DFF \start_reg_reg[55]  ( .D(start_in[54]), .CLK(clk), .RST(rst), .Q(
        start_reg[55]) );
  DFF \start_reg_reg[56]  ( .D(start_in[55]), .CLK(clk), .RST(rst), .Q(
        start_reg[56]) );
  DFF \start_reg_reg[57]  ( .D(start_in[56]), .CLK(clk), .RST(rst), .Q(
        start_reg[57]) );
  DFF \start_reg_reg[58]  ( .D(start_in[57]), .CLK(clk), .RST(rst), .Q(
        start_reg[58]) );
  DFF \start_reg_reg[59]  ( .D(start_in[58]), .CLK(clk), .RST(rst), .Q(
        start_reg[59]) );
  DFF \start_reg_reg[60]  ( .D(start_in[59]), .CLK(clk), .RST(rst), .Q(
        start_reg[60]) );
  DFF \start_reg_reg[61]  ( .D(start_in[60]), .CLK(clk), .RST(rst), .Q(
        start_reg[61]) );
  DFF \start_reg_reg[62]  ( .D(start_in[61]), .CLK(clk), .RST(rst), .Q(
        start_reg[62]) );
  DFF \start_reg_reg[63]  ( .D(start_in[62]), .CLK(clk), .RST(rst), .Q(
        start_reg[63]) );
  DFF \start_reg_reg[64]  ( .D(start_in[63]), .CLK(clk), .RST(rst), .Q(
        start_reg[64]) );
  DFF \start_reg_reg[65]  ( .D(start_in[64]), .CLK(clk), .RST(rst), .Q(
        start_reg[65]) );
  DFF \start_reg_reg[66]  ( .D(start_in[65]), .CLK(clk), .RST(rst), .Q(
        start_reg[66]) );
  DFF \start_reg_reg[67]  ( .D(start_in[66]), .CLK(clk), .RST(rst), .Q(
        start_reg[67]) );
  DFF \start_reg_reg[68]  ( .D(start_in[67]), .CLK(clk), .RST(rst), .Q(
        start_reg[68]) );
  DFF \start_reg_reg[69]  ( .D(start_in[68]), .CLK(clk), .RST(rst), .Q(
        start_reg[69]) );
  DFF \start_reg_reg[70]  ( .D(start_in[69]), .CLK(clk), .RST(rst), .Q(
        start_reg[70]) );
  DFF \start_reg_reg[71]  ( .D(start_in[70]), .CLK(clk), .RST(rst), .Q(
        start_reg[71]) );
  DFF \start_reg_reg[72]  ( .D(start_in[71]), .CLK(clk), .RST(rst), .Q(
        start_reg[72]) );
  DFF \start_reg_reg[73]  ( .D(start_in[72]), .CLK(clk), .RST(rst), .Q(
        start_reg[73]) );
  DFF \start_reg_reg[74]  ( .D(start_in[73]), .CLK(clk), .RST(rst), .Q(
        start_reg[74]) );
  DFF \start_reg_reg[75]  ( .D(start_in[74]), .CLK(clk), .RST(rst), .Q(
        start_reg[75]) );
  DFF \start_reg_reg[76]  ( .D(start_in[75]), .CLK(clk), .RST(rst), .Q(
        start_reg[76]) );
  DFF \start_reg_reg[77]  ( .D(start_in[76]), .CLK(clk), .RST(rst), .Q(
        start_reg[77]) );
  DFF \start_reg_reg[78]  ( .D(start_in[77]), .CLK(clk), .RST(rst), .Q(
        start_reg[78]) );
  DFF \start_reg_reg[79]  ( .D(start_in[78]), .CLK(clk), .RST(rst), .Q(
        start_reg[79]) );
  DFF \start_reg_reg[80]  ( .D(start_in[79]), .CLK(clk), .RST(rst), .Q(
        start_reg[80]) );
  DFF \start_reg_reg[81]  ( .D(start_in[80]), .CLK(clk), .RST(rst), .Q(
        start_reg[81]) );
  DFF \start_reg_reg[82]  ( .D(start_in[81]), .CLK(clk), .RST(rst), .Q(
        start_reg[82]) );
  DFF \start_reg_reg[83]  ( .D(start_in[82]), .CLK(clk), .RST(rst), .Q(
        start_reg[83]) );
  DFF \start_reg_reg[84]  ( .D(start_in[83]), .CLK(clk), .RST(rst), .Q(
        start_reg[84]) );
  DFF \start_reg_reg[85]  ( .D(start_in[84]), .CLK(clk), .RST(rst), .Q(
        start_reg[85]) );
  DFF \start_reg_reg[86]  ( .D(start_in[85]), .CLK(clk), .RST(rst), .Q(
        start_reg[86]) );
  DFF \start_reg_reg[87]  ( .D(start_in[86]), .CLK(clk), .RST(rst), .Q(
        start_reg[87]) );
  DFF \start_reg_reg[88]  ( .D(start_in[87]), .CLK(clk), .RST(rst), .Q(
        start_reg[88]) );
  DFF \start_reg_reg[89]  ( .D(start_in[88]), .CLK(clk), .RST(rst), .Q(
        start_reg[89]) );
  DFF \start_reg_reg[90]  ( .D(start_in[89]), .CLK(clk), .RST(rst), .Q(
        start_reg[90]) );
  DFF \start_reg_reg[91]  ( .D(start_in[90]), .CLK(clk), .RST(rst), .Q(
        start_reg[91]) );
  DFF \start_reg_reg[92]  ( .D(start_in[91]), .CLK(clk), .RST(rst), .Q(
        start_reg[92]) );
  DFF \start_reg_reg[93]  ( .D(start_in[92]), .CLK(clk), .RST(rst), .Q(
        start_reg[93]) );
  DFF \start_reg_reg[94]  ( .D(start_in[93]), .CLK(clk), .RST(rst), .Q(
        start_reg[94]) );
  DFF \start_reg_reg[95]  ( .D(start_in[94]), .CLK(clk), .RST(rst), .Q(
        start_reg[95]) );
  DFF \start_reg_reg[96]  ( .D(start_in[95]), .CLK(clk), .RST(rst), .Q(
        start_reg[96]) );
  DFF \start_reg_reg[97]  ( .D(start_in[96]), .CLK(clk), .RST(rst), .Q(
        start_reg[97]) );
  DFF \start_reg_reg[98]  ( .D(start_in[97]), .CLK(clk), .RST(rst), .Q(
        start_reg[98]) );
  DFF \start_reg_reg[99]  ( .D(start_in[98]), .CLK(clk), .RST(rst), .Q(
        start_reg[99]) );
  DFF \start_reg_reg[100]  ( .D(start_in[99]), .CLK(clk), .RST(rst), .Q(
        start_reg[100]) );
  DFF \start_reg_reg[101]  ( .D(start_in[100]), .CLK(clk), .RST(rst), .Q(
        start_reg[101]) );
  DFF \start_reg_reg[102]  ( .D(start_in[101]), .CLK(clk), .RST(rst), .Q(
        start_reg[102]) );
  DFF \start_reg_reg[103]  ( .D(start_in[102]), .CLK(clk), .RST(rst), .Q(
        start_reg[103]) );
  DFF \start_reg_reg[104]  ( .D(start_in[103]), .CLK(clk), .RST(rst), .Q(
        start_reg[104]) );
  DFF \start_reg_reg[105]  ( .D(start_in[104]), .CLK(clk), .RST(rst), .Q(
        start_reg[105]) );
  DFF \start_reg_reg[106]  ( .D(start_in[105]), .CLK(clk), .RST(rst), .Q(
        start_reg[106]) );
  DFF \start_reg_reg[107]  ( .D(start_in[106]), .CLK(clk), .RST(rst), .Q(
        start_reg[107]) );
  DFF \start_reg_reg[108]  ( .D(start_in[107]), .CLK(clk), .RST(rst), .Q(
        start_reg[108]) );
  DFF \start_reg_reg[109]  ( .D(start_in[108]), .CLK(clk), .RST(rst), .Q(
        start_reg[109]) );
  DFF \start_reg_reg[110]  ( .D(start_in[109]), .CLK(clk), .RST(rst), .Q(
        start_reg[110]) );
  DFF \start_reg_reg[111]  ( .D(start_in[110]), .CLK(clk), .RST(rst), .Q(
        start_reg[111]) );
  DFF \start_reg_reg[112]  ( .D(start_in[111]), .CLK(clk), .RST(rst), .Q(
        start_reg[112]) );
  DFF \start_reg_reg[113]  ( .D(start_in[112]), .CLK(clk), .RST(rst), .Q(
        start_reg[113]) );
  DFF \start_reg_reg[114]  ( .D(start_in[113]), .CLK(clk), .RST(rst), .Q(
        start_reg[114]) );
  DFF \start_reg_reg[115]  ( .D(start_in[114]), .CLK(clk), .RST(rst), .Q(
        start_reg[115]) );
  DFF \start_reg_reg[116]  ( .D(start_in[115]), .CLK(clk), .RST(rst), .Q(
        start_reg[116]) );
  DFF \start_reg_reg[117]  ( .D(start_in[116]), .CLK(clk), .RST(rst), .Q(
        start_reg[117]) );
  DFF \start_reg_reg[118]  ( .D(start_in[117]), .CLK(clk), .RST(rst), .Q(
        start_reg[118]) );
  DFF \start_reg_reg[119]  ( .D(start_in[118]), .CLK(clk), .RST(rst), .Q(
        start_reg[119]) );
  DFF \start_reg_reg[120]  ( .D(start_in[119]), .CLK(clk), .RST(rst), .Q(
        start_reg[120]) );
  DFF \start_reg_reg[121]  ( .D(start_in[120]), .CLK(clk), .RST(rst), .Q(
        start_reg[121]) );
  DFF \start_reg_reg[122]  ( .D(start_in[121]), .CLK(clk), .RST(rst), .Q(
        start_reg[122]) );
  DFF \start_reg_reg[123]  ( .D(start_in[122]), .CLK(clk), .RST(rst), .Q(
        start_reg[123]) );
  DFF \start_reg_reg[124]  ( .D(start_in[123]), .CLK(clk), .RST(rst), .Q(
        start_reg[124]) );
  DFF \start_reg_reg[125]  ( .D(start_in[124]), .CLK(clk), .RST(rst), .Q(
        start_reg[125]) );
  DFF \start_reg_reg[126]  ( .D(start_in[125]), .CLK(clk), .RST(rst), .Q(
        start_reg[126]) );
  DFF \start_reg_reg[127]  ( .D(start_in[126]), .CLK(clk), .RST(rst), .Q(
        start_reg[127]) );
  DFF \start_reg_reg[128]  ( .D(start_in[127]), .CLK(clk), .RST(rst), .Q(
        start_reg[128]) );
  DFF \start_reg_reg[129]  ( .D(start_in[128]), .CLK(clk), .RST(rst), .Q(
        start_reg[129]) );
  DFF \start_reg_reg[130]  ( .D(start_in[129]), .CLK(clk), .RST(rst), .Q(
        start_reg[130]) );
  DFF \start_reg_reg[131]  ( .D(start_in[130]), .CLK(clk), .RST(rst), .Q(
        start_reg[131]) );
  DFF \start_reg_reg[132]  ( .D(start_in[131]), .CLK(clk), .RST(rst), .Q(
        start_reg[132]) );
  DFF \start_reg_reg[133]  ( .D(start_in[132]), .CLK(clk), .RST(rst), .Q(
        start_reg[133]) );
  DFF \start_reg_reg[134]  ( .D(start_in[133]), .CLK(clk), .RST(rst), .Q(
        start_reg[134]) );
  DFF \start_reg_reg[135]  ( .D(start_in[134]), .CLK(clk), .RST(rst), .Q(
        start_reg[135]) );
  DFF \start_reg_reg[136]  ( .D(start_in[135]), .CLK(clk), .RST(rst), .Q(
        start_reg[136]) );
  DFF \start_reg_reg[137]  ( .D(start_in[136]), .CLK(clk), .RST(rst), .Q(
        start_reg[137]) );
  DFF \start_reg_reg[138]  ( .D(start_in[137]), .CLK(clk), .RST(rst), .Q(
        start_reg[138]) );
  DFF \start_reg_reg[139]  ( .D(start_in[138]), .CLK(clk), .RST(rst), .Q(
        start_reg[139]) );
  DFF \start_reg_reg[140]  ( .D(start_in[139]), .CLK(clk), .RST(rst), .Q(
        start_reg[140]) );
  DFF \start_reg_reg[141]  ( .D(start_in[140]), .CLK(clk), .RST(rst), .Q(
        start_reg[141]) );
  DFF \start_reg_reg[142]  ( .D(start_in[141]), .CLK(clk), .RST(rst), .Q(
        start_reg[142]) );
  DFF \start_reg_reg[143]  ( .D(start_in[142]), .CLK(clk), .RST(rst), .Q(
        start_reg[143]) );
  DFF \start_reg_reg[144]  ( .D(start_in[143]), .CLK(clk), .RST(rst), .Q(
        start_reg[144]) );
  DFF \start_reg_reg[145]  ( .D(start_in[144]), .CLK(clk), .RST(rst), .Q(
        start_reg[145]) );
  DFF \start_reg_reg[146]  ( .D(start_in[145]), .CLK(clk), .RST(rst), .Q(
        start_reg[146]) );
  DFF \start_reg_reg[147]  ( .D(start_in[146]), .CLK(clk), .RST(rst), .Q(
        start_reg[147]) );
  DFF \start_reg_reg[148]  ( .D(start_in[147]), .CLK(clk), .RST(rst), .Q(
        start_reg[148]) );
  DFF \start_reg_reg[149]  ( .D(start_in[148]), .CLK(clk), .RST(rst), .Q(
        start_reg[149]) );
  DFF \start_reg_reg[150]  ( .D(start_in[149]), .CLK(clk), .RST(rst), .Q(
        start_reg[150]) );
  DFF \start_reg_reg[151]  ( .D(start_in[150]), .CLK(clk), .RST(rst), .Q(
        start_reg[151]) );
  DFF \start_reg_reg[152]  ( .D(start_in[151]), .CLK(clk), .RST(rst), .Q(
        start_reg[152]) );
  DFF \start_reg_reg[153]  ( .D(start_in[152]), .CLK(clk), .RST(rst), .Q(
        start_reg[153]) );
  DFF \start_reg_reg[154]  ( .D(start_in[153]), .CLK(clk), .RST(rst), .Q(
        start_reg[154]) );
  DFF \start_reg_reg[155]  ( .D(start_in[154]), .CLK(clk), .RST(rst), .Q(
        start_reg[155]) );
  DFF \start_reg_reg[156]  ( .D(start_in[155]), .CLK(clk), .RST(rst), .Q(
        start_reg[156]) );
  DFF \start_reg_reg[157]  ( .D(start_in[156]), .CLK(clk), .RST(rst), .Q(
        start_reg[157]) );
  DFF \start_reg_reg[158]  ( .D(start_in[157]), .CLK(clk), .RST(rst), .Q(
        start_reg[158]) );
  DFF \start_reg_reg[159]  ( .D(start_in[158]), .CLK(clk), .RST(rst), .Q(
        start_reg[159]) );
  DFF \start_reg_reg[160]  ( .D(start_in[159]), .CLK(clk), .RST(rst), .Q(
        start_reg[160]) );
  DFF \start_reg_reg[161]  ( .D(start_in[160]), .CLK(clk), .RST(rst), .Q(
        start_reg[161]) );
  DFF \start_reg_reg[162]  ( .D(start_in[161]), .CLK(clk), .RST(rst), .Q(
        start_reg[162]) );
  DFF \start_reg_reg[163]  ( .D(start_in[162]), .CLK(clk), .RST(rst), .Q(
        start_reg[163]) );
  DFF \start_reg_reg[164]  ( .D(start_in[163]), .CLK(clk), .RST(rst), .Q(
        start_reg[164]) );
  DFF \start_reg_reg[165]  ( .D(start_in[164]), .CLK(clk), .RST(rst), .Q(
        start_reg[165]) );
  DFF \start_reg_reg[166]  ( .D(start_in[165]), .CLK(clk), .RST(rst), .Q(
        start_reg[166]) );
  DFF \start_reg_reg[167]  ( .D(start_in[166]), .CLK(clk), .RST(rst), .Q(
        start_reg[167]) );
  DFF \start_reg_reg[168]  ( .D(start_in[167]), .CLK(clk), .RST(rst), .Q(
        start_reg[168]) );
  DFF \start_reg_reg[169]  ( .D(start_in[168]), .CLK(clk), .RST(rst), .Q(
        start_reg[169]) );
  DFF \start_reg_reg[170]  ( .D(start_in[169]), .CLK(clk), .RST(rst), .Q(
        start_reg[170]) );
  DFF \start_reg_reg[171]  ( .D(start_in[170]), .CLK(clk), .RST(rst), .Q(
        start_reg[171]) );
  DFF \start_reg_reg[172]  ( .D(start_in[171]), .CLK(clk), .RST(rst), .Q(
        start_reg[172]) );
  DFF \start_reg_reg[173]  ( .D(start_in[172]), .CLK(clk), .RST(rst), .Q(
        start_reg[173]) );
  DFF \start_reg_reg[174]  ( .D(start_in[173]), .CLK(clk), .RST(rst), .Q(
        start_reg[174]) );
  DFF \start_reg_reg[175]  ( .D(start_in[174]), .CLK(clk), .RST(rst), .Q(
        start_reg[175]) );
  DFF \start_reg_reg[176]  ( .D(start_in[175]), .CLK(clk), .RST(rst), .Q(
        start_reg[176]) );
  DFF \start_reg_reg[177]  ( .D(start_in[176]), .CLK(clk), .RST(rst), .Q(
        start_reg[177]) );
  DFF \start_reg_reg[178]  ( .D(start_in[177]), .CLK(clk), .RST(rst), .Q(
        start_reg[178]) );
  DFF \start_reg_reg[179]  ( .D(start_in[178]), .CLK(clk), .RST(rst), .Q(
        start_reg[179]) );
  DFF \start_reg_reg[180]  ( .D(start_in[179]), .CLK(clk), .RST(rst), .Q(
        start_reg[180]) );
  DFF \start_reg_reg[181]  ( .D(start_in[180]), .CLK(clk), .RST(rst), .Q(
        start_reg[181]) );
  DFF \start_reg_reg[182]  ( .D(start_in[181]), .CLK(clk), .RST(rst), .Q(
        start_reg[182]) );
  DFF \start_reg_reg[183]  ( .D(start_in[182]), .CLK(clk), .RST(rst), .Q(
        start_reg[183]) );
  DFF \start_reg_reg[184]  ( .D(start_in[183]), .CLK(clk), .RST(rst), .Q(
        start_reg[184]) );
  DFF \start_reg_reg[185]  ( .D(start_in[184]), .CLK(clk), .RST(rst), .Q(
        start_reg[185]) );
  DFF \start_reg_reg[186]  ( .D(start_in[185]), .CLK(clk), .RST(rst), .Q(
        start_reg[186]) );
  DFF \start_reg_reg[187]  ( .D(start_in[186]), .CLK(clk), .RST(rst), .Q(
        start_reg[187]) );
  DFF \start_reg_reg[188]  ( .D(start_in[187]), .CLK(clk), .RST(rst), .Q(
        start_reg[188]) );
  DFF \start_reg_reg[189]  ( .D(start_in[188]), .CLK(clk), .RST(rst), .Q(
        start_reg[189]) );
  DFF \start_reg_reg[190]  ( .D(start_in[189]), .CLK(clk), .RST(rst), .Q(
        start_reg[190]) );
  DFF \start_reg_reg[191]  ( .D(start_in[190]), .CLK(clk), .RST(rst), .Q(
        start_reg[191]) );
  DFF \start_reg_reg[192]  ( .D(start_in[191]), .CLK(clk), .RST(rst), .Q(
        start_reg[192]) );
  DFF \start_reg_reg[193]  ( .D(start_in[192]), .CLK(clk), .RST(rst), .Q(
        start_reg[193]) );
  DFF \start_reg_reg[194]  ( .D(start_in[193]), .CLK(clk), .RST(rst), .Q(
        start_reg[194]) );
  DFF \start_reg_reg[195]  ( .D(start_in[194]), .CLK(clk), .RST(rst), .Q(
        start_reg[195]) );
  DFF \start_reg_reg[196]  ( .D(start_in[195]), .CLK(clk), .RST(rst), .Q(
        start_reg[196]) );
  DFF \start_reg_reg[197]  ( .D(start_in[196]), .CLK(clk), .RST(rst), .Q(
        start_reg[197]) );
  DFF \start_reg_reg[198]  ( .D(start_in[197]), .CLK(clk), .RST(rst), .Q(
        start_reg[198]) );
  DFF \start_reg_reg[199]  ( .D(start_in[198]), .CLK(clk), .RST(rst), .Q(
        start_reg[199]) );
  DFF \start_reg_reg[200]  ( .D(start_in[199]), .CLK(clk), .RST(rst), .Q(
        start_reg[200]) );
  DFF \start_reg_reg[201]  ( .D(start_in[200]), .CLK(clk), .RST(rst), .Q(
        start_reg[201]) );
  DFF \start_reg_reg[202]  ( .D(start_in[201]), .CLK(clk), .RST(rst), .Q(
        start_reg[202]) );
  DFF \start_reg_reg[203]  ( .D(start_in[202]), .CLK(clk), .RST(rst), .Q(
        start_reg[203]) );
  DFF \start_reg_reg[204]  ( .D(start_in[203]), .CLK(clk), .RST(rst), .Q(
        start_reg[204]) );
  DFF \start_reg_reg[205]  ( .D(start_in[204]), .CLK(clk), .RST(rst), .Q(
        start_reg[205]) );
  DFF \start_reg_reg[206]  ( .D(start_in[205]), .CLK(clk), .RST(rst), .Q(
        start_reg[206]) );
  DFF \start_reg_reg[207]  ( .D(start_in[206]), .CLK(clk), .RST(rst), .Q(
        start_reg[207]) );
  DFF \start_reg_reg[208]  ( .D(start_in[207]), .CLK(clk), .RST(rst), .Q(
        start_reg[208]) );
  DFF \start_reg_reg[209]  ( .D(start_in[208]), .CLK(clk), .RST(rst), .Q(
        start_reg[209]) );
  DFF \start_reg_reg[210]  ( .D(start_in[209]), .CLK(clk), .RST(rst), .Q(
        start_reg[210]) );
  DFF \start_reg_reg[211]  ( .D(start_in[210]), .CLK(clk), .RST(rst), .Q(
        start_reg[211]) );
  DFF \start_reg_reg[212]  ( .D(start_in[211]), .CLK(clk), .RST(rst), .Q(
        start_reg[212]) );
  DFF \start_reg_reg[213]  ( .D(start_in[212]), .CLK(clk), .RST(rst), .Q(
        start_reg[213]) );
  DFF \start_reg_reg[214]  ( .D(start_in[213]), .CLK(clk), .RST(rst), .Q(
        start_reg[214]) );
  DFF \start_reg_reg[215]  ( .D(start_in[214]), .CLK(clk), .RST(rst), .Q(
        start_reg[215]) );
  DFF \start_reg_reg[216]  ( .D(start_in[215]), .CLK(clk), .RST(rst), .Q(
        start_reg[216]) );
  DFF \start_reg_reg[217]  ( .D(start_in[216]), .CLK(clk), .RST(rst), .Q(
        start_reg[217]) );
  DFF \start_reg_reg[218]  ( .D(start_in[217]), .CLK(clk), .RST(rst), .Q(
        start_reg[218]) );
  DFF \start_reg_reg[219]  ( .D(start_in[218]), .CLK(clk), .RST(rst), .Q(
        start_reg[219]) );
  DFF \start_reg_reg[220]  ( .D(start_in[219]), .CLK(clk), .RST(rst), .Q(
        start_reg[220]) );
  DFF \start_reg_reg[221]  ( .D(start_in[220]), .CLK(clk), .RST(rst), .Q(
        start_reg[221]) );
  DFF \start_reg_reg[222]  ( .D(start_in[221]), .CLK(clk), .RST(rst), .Q(
        start_reg[222]) );
  DFF \start_reg_reg[223]  ( .D(start_in[222]), .CLK(clk), .RST(rst), .Q(
        start_reg[223]) );
  DFF \start_reg_reg[224]  ( .D(start_in[223]), .CLK(clk), .RST(rst), .Q(
        start_reg[224]) );
  DFF \start_reg_reg[225]  ( .D(start_in[224]), .CLK(clk), .RST(rst), .Q(
        start_reg[225]) );
  DFF \start_reg_reg[226]  ( .D(start_in[225]), .CLK(clk), .RST(rst), .Q(
        start_reg[226]) );
  DFF \start_reg_reg[227]  ( .D(start_in[226]), .CLK(clk), .RST(rst), .Q(
        start_reg[227]) );
  DFF \start_reg_reg[228]  ( .D(start_in[227]), .CLK(clk), .RST(rst), .Q(
        start_reg[228]) );
  DFF \start_reg_reg[229]  ( .D(start_in[228]), .CLK(clk), .RST(rst), .Q(
        start_reg[229]) );
  DFF \start_reg_reg[230]  ( .D(start_in[229]), .CLK(clk), .RST(rst), .Q(
        start_reg[230]) );
  DFF \start_reg_reg[231]  ( .D(start_in[230]), .CLK(clk), .RST(rst), .Q(
        start_reg[231]) );
  DFF \start_reg_reg[232]  ( .D(start_in[231]), .CLK(clk), .RST(rst), .Q(
        start_reg[232]) );
  DFF \start_reg_reg[233]  ( .D(start_in[232]), .CLK(clk), .RST(rst), .Q(
        start_reg[233]) );
  DFF \start_reg_reg[234]  ( .D(start_in[233]), .CLK(clk), .RST(rst), .Q(
        start_reg[234]) );
  DFF \start_reg_reg[235]  ( .D(start_in[234]), .CLK(clk), .RST(rst), .Q(
        start_reg[235]) );
  DFF \start_reg_reg[236]  ( .D(start_in[235]), .CLK(clk), .RST(rst), .Q(
        start_reg[236]) );
  DFF \start_reg_reg[237]  ( .D(start_in[236]), .CLK(clk), .RST(rst), .Q(
        start_reg[237]) );
  DFF \start_reg_reg[238]  ( .D(start_in[237]), .CLK(clk), .RST(rst), .Q(
        start_reg[238]) );
  DFF \start_reg_reg[239]  ( .D(start_in[238]), .CLK(clk), .RST(rst), .Q(
        start_reg[239]) );
  DFF \start_reg_reg[240]  ( .D(start_in[239]), .CLK(clk), .RST(rst), .Q(
        start_reg[240]) );
  DFF \start_reg_reg[241]  ( .D(start_in[240]), .CLK(clk), .RST(rst), .Q(
        start_reg[241]) );
  DFF \start_reg_reg[242]  ( .D(start_in[241]), .CLK(clk), .RST(rst), .Q(
        start_reg[242]) );
  DFF \start_reg_reg[243]  ( .D(start_in[242]), .CLK(clk), .RST(rst), .Q(
        start_reg[243]) );
  DFF \start_reg_reg[244]  ( .D(start_in[243]), .CLK(clk), .RST(rst), .Q(
        start_reg[244]) );
  DFF \start_reg_reg[245]  ( .D(start_in[244]), .CLK(clk), .RST(rst), .Q(
        start_reg[245]) );
  DFF \start_reg_reg[246]  ( .D(start_in[245]), .CLK(clk), .RST(rst), .Q(
        start_reg[246]) );
  DFF \start_reg_reg[247]  ( .D(start_in[246]), .CLK(clk), .RST(rst), .Q(
        start_reg[247]) );
  DFF \start_reg_reg[248]  ( .D(start_in[247]), .CLK(clk), .RST(rst), .Q(
        start_reg[248]) );
  DFF \start_reg_reg[249]  ( .D(start_in[248]), .CLK(clk), .RST(rst), .Q(
        start_reg[249]) );
  DFF \start_reg_reg[250]  ( .D(start_in[249]), .CLK(clk), .RST(rst), .Q(
        start_reg[250]) );
  DFF \start_reg_reg[251]  ( .D(start_in[250]), .CLK(clk), .RST(rst), .Q(
        start_reg[251]) );
  DFF \start_reg_reg[252]  ( .D(start_in[251]), .CLK(clk), .RST(rst), .Q(
        start_reg[252]) );
  DFF \start_reg_reg[253]  ( .D(start_in[252]), .CLK(clk), .RST(rst), .Q(
        start_reg[253]) );
  DFF \start_reg_reg[254]  ( .D(start_in[253]), .CLK(clk), .RST(rst), .Q(
        start_reg[254]) );
  DFF \start_reg_reg[255]  ( .D(start_in[254]), .CLK(clk), .RST(rst), .Q(
        start_reg[255]) );
  DFF \start_reg_reg[256]  ( .D(start_in[255]), .CLK(clk), .RST(rst), .Q(
        start_reg[256]) );
  DFF \start_reg_reg[257]  ( .D(start_in[256]), .CLK(clk), .RST(rst), .Q(
        start_reg[257]) );
  DFF \start_reg_reg[258]  ( .D(start_in[257]), .CLK(clk), .RST(rst), .Q(
        start_reg[258]) );
  DFF \start_reg_reg[259]  ( .D(start_in[258]), .CLK(clk), .RST(rst), .Q(
        start_reg[259]) );
  DFF \start_reg_reg[260]  ( .D(start_in[259]), .CLK(clk), .RST(rst), .Q(
        start_reg[260]) );
  DFF \start_reg_reg[261]  ( .D(start_in[260]), .CLK(clk), .RST(rst), .Q(
        start_reg[261]) );
  DFF \start_reg_reg[262]  ( .D(start_in[261]), .CLK(clk), .RST(rst), .Q(
        start_reg[262]) );
  DFF \start_reg_reg[263]  ( .D(start_in[262]), .CLK(clk), .RST(rst), .Q(
        start_reg[263]) );
  DFF \start_reg_reg[264]  ( .D(start_in[263]), .CLK(clk), .RST(rst), .Q(
        start_reg[264]) );
  DFF \start_reg_reg[265]  ( .D(start_in[264]), .CLK(clk), .RST(rst), .Q(
        start_reg[265]) );
  DFF \start_reg_reg[266]  ( .D(start_in[265]), .CLK(clk), .RST(rst), .Q(
        start_reg[266]) );
  DFF \start_reg_reg[267]  ( .D(start_in[266]), .CLK(clk), .RST(rst), .Q(
        start_reg[267]) );
  DFF \start_reg_reg[268]  ( .D(start_in[267]), .CLK(clk), .RST(rst), .Q(
        start_reg[268]) );
  DFF \start_reg_reg[269]  ( .D(start_in[268]), .CLK(clk), .RST(rst), .Q(
        start_reg[269]) );
  DFF \start_reg_reg[270]  ( .D(start_in[269]), .CLK(clk), .RST(rst), .Q(
        start_reg[270]) );
  DFF \start_reg_reg[271]  ( .D(start_in[270]), .CLK(clk), .RST(rst), .Q(
        start_reg[271]) );
  DFF \start_reg_reg[272]  ( .D(start_in[271]), .CLK(clk), .RST(rst), .Q(
        start_reg[272]) );
  DFF \start_reg_reg[273]  ( .D(start_in[272]), .CLK(clk), .RST(rst), .Q(
        start_reg[273]) );
  DFF \start_reg_reg[274]  ( .D(start_in[273]), .CLK(clk), .RST(rst), .Q(
        start_reg[274]) );
  DFF \start_reg_reg[275]  ( .D(start_in[274]), .CLK(clk), .RST(rst), .Q(
        start_reg[275]) );
  DFF \start_reg_reg[276]  ( .D(start_in[275]), .CLK(clk), .RST(rst), .Q(
        start_reg[276]) );
  DFF \start_reg_reg[277]  ( .D(start_in[276]), .CLK(clk), .RST(rst), .Q(
        start_reg[277]) );
  DFF \start_reg_reg[278]  ( .D(start_in[277]), .CLK(clk), .RST(rst), .Q(
        start_reg[278]) );
  DFF \start_reg_reg[279]  ( .D(start_in[278]), .CLK(clk), .RST(rst), .Q(
        start_reg[279]) );
  DFF \start_reg_reg[280]  ( .D(start_in[279]), .CLK(clk), .RST(rst), .Q(
        start_reg[280]) );
  DFF \start_reg_reg[281]  ( .D(start_in[280]), .CLK(clk), .RST(rst), .Q(
        start_reg[281]) );
  DFF \start_reg_reg[282]  ( .D(start_in[281]), .CLK(clk), .RST(rst), .Q(
        start_reg[282]) );
  DFF \start_reg_reg[283]  ( .D(start_in[282]), .CLK(clk), .RST(rst), .Q(
        start_reg[283]) );
  DFF \start_reg_reg[284]  ( .D(start_in[283]), .CLK(clk), .RST(rst), .Q(
        start_reg[284]) );
  DFF \start_reg_reg[285]  ( .D(start_in[284]), .CLK(clk), .RST(rst), .Q(
        start_reg[285]) );
  DFF \start_reg_reg[286]  ( .D(start_in[285]), .CLK(clk), .RST(rst), .Q(
        start_reg[286]) );
  DFF \start_reg_reg[287]  ( .D(start_in[286]), .CLK(clk), .RST(rst), .Q(
        start_reg[287]) );
  DFF \start_reg_reg[288]  ( .D(start_in[287]), .CLK(clk), .RST(rst), .Q(
        start_reg[288]) );
  DFF \start_reg_reg[289]  ( .D(start_in[288]), .CLK(clk), .RST(rst), .Q(
        start_reg[289]) );
  DFF \start_reg_reg[290]  ( .D(start_in[289]), .CLK(clk), .RST(rst), .Q(
        start_reg[290]) );
  DFF \start_reg_reg[291]  ( .D(start_in[290]), .CLK(clk), .RST(rst), .Q(
        start_reg[291]) );
  DFF \start_reg_reg[292]  ( .D(start_in[291]), .CLK(clk), .RST(rst), .Q(
        start_reg[292]) );
  DFF \start_reg_reg[293]  ( .D(start_in[292]), .CLK(clk), .RST(rst), .Q(
        start_reg[293]) );
  DFF \start_reg_reg[294]  ( .D(start_in[293]), .CLK(clk), .RST(rst), .Q(
        start_reg[294]) );
  DFF \start_reg_reg[295]  ( .D(start_in[294]), .CLK(clk), .RST(rst), .Q(
        start_reg[295]) );
  DFF \start_reg_reg[296]  ( .D(start_in[295]), .CLK(clk), .RST(rst), .Q(
        start_reg[296]) );
  DFF \start_reg_reg[297]  ( .D(start_in[296]), .CLK(clk), .RST(rst), .Q(
        start_reg[297]) );
  DFF \start_reg_reg[298]  ( .D(start_in[297]), .CLK(clk), .RST(rst), .Q(
        start_reg[298]) );
  DFF \start_reg_reg[299]  ( .D(start_in[298]), .CLK(clk), .RST(rst), .Q(
        start_reg[299]) );
  DFF \start_reg_reg[300]  ( .D(start_in[299]), .CLK(clk), .RST(rst), .Q(
        start_reg[300]) );
  DFF \start_reg_reg[301]  ( .D(start_in[300]), .CLK(clk), .RST(rst), .Q(
        start_reg[301]) );
  DFF \start_reg_reg[302]  ( .D(start_in[301]), .CLK(clk), .RST(rst), .Q(
        start_reg[302]) );
  DFF \start_reg_reg[303]  ( .D(start_in[302]), .CLK(clk), .RST(rst), .Q(
        start_reg[303]) );
  DFF \start_reg_reg[304]  ( .D(start_in[303]), .CLK(clk), .RST(rst), .Q(
        start_reg[304]) );
  DFF \start_reg_reg[305]  ( .D(start_in[304]), .CLK(clk), .RST(rst), .Q(
        start_reg[305]) );
  DFF \start_reg_reg[306]  ( .D(start_in[305]), .CLK(clk), .RST(rst), .Q(
        start_reg[306]) );
  DFF \start_reg_reg[307]  ( .D(start_in[306]), .CLK(clk), .RST(rst), .Q(
        start_reg[307]) );
  DFF \start_reg_reg[308]  ( .D(start_in[307]), .CLK(clk), .RST(rst), .Q(
        start_reg[308]) );
  DFF \start_reg_reg[309]  ( .D(start_in[308]), .CLK(clk), .RST(rst), .Q(
        start_reg[309]) );
  DFF \start_reg_reg[310]  ( .D(start_in[309]), .CLK(clk), .RST(rst), .Q(
        start_reg[310]) );
  DFF \start_reg_reg[311]  ( .D(start_in[310]), .CLK(clk), .RST(rst), .Q(
        start_reg[311]) );
  DFF \start_reg_reg[312]  ( .D(start_in[311]), .CLK(clk), .RST(rst), .Q(
        start_reg[312]) );
  DFF \start_reg_reg[313]  ( .D(start_in[312]), .CLK(clk), .RST(rst), .Q(
        start_reg[313]) );
  DFF \start_reg_reg[314]  ( .D(start_in[313]), .CLK(clk), .RST(rst), .Q(
        start_reg[314]) );
  DFF \start_reg_reg[315]  ( .D(start_in[314]), .CLK(clk), .RST(rst), .Q(
        start_reg[315]) );
  DFF \start_reg_reg[316]  ( .D(start_in[315]), .CLK(clk), .RST(rst), .Q(
        start_reg[316]) );
  DFF \start_reg_reg[317]  ( .D(start_in[316]), .CLK(clk), .RST(rst), .Q(
        start_reg[317]) );
  DFF \start_reg_reg[318]  ( .D(start_in[317]), .CLK(clk), .RST(rst), .Q(
        start_reg[318]) );
  DFF \start_reg_reg[319]  ( .D(start_in[318]), .CLK(clk), .RST(rst), .Q(
        start_reg[319]) );
  DFF \start_reg_reg[320]  ( .D(start_in[319]), .CLK(clk), .RST(rst), .Q(
        start_reg[320]) );
  DFF \start_reg_reg[321]  ( .D(start_in[320]), .CLK(clk), .RST(rst), .Q(
        start_reg[321]) );
  DFF \start_reg_reg[322]  ( .D(start_in[321]), .CLK(clk), .RST(rst), .Q(
        start_reg[322]) );
  DFF \start_reg_reg[323]  ( .D(start_in[322]), .CLK(clk), .RST(rst), .Q(
        start_reg[323]) );
  DFF \start_reg_reg[324]  ( .D(start_in[323]), .CLK(clk), .RST(rst), .Q(
        start_reg[324]) );
  DFF \start_reg_reg[325]  ( .D(start_in[324]), .CLK(clk), .RST(rst), .Q(
        start_reg[325]) );
  DFF \start_reg_reg[326]  ( .D(start_in[325]), .CLK(clk), .RST(rst), .Q(
        start_reg[326]) );
  DFF \start_reg_reg[327]  ( .D(start_in[326]), .CLK(clk), .RST(rst), .Q(
        start_reg[327]) );
  DFF \start_reg_reg[328]  ( .D(start_in[327]), .CLK(clk), .RST(rst), .Q(
        start_reg[328]) );
  DFF \start_reg_reg[329]  ( .D(start_in[328]), .CLK(clk), .RST(rst), .Q(
        start_reg[329]) );
  DFF \start_reg_reg[330]  ( .D(start_in[329]), .CLK(clk), .RST(rst), .Q(
        start_reg[330]) );
  DFF \start_reg_reg[331]  ( .D(start_in[330]), .CLK(clk), .RST(rst), .Q(
        start_reg[331]) );
  DFF \start_reg_reg[332]  ( .D(start_in[331]), .CLK(clk), .RST(rst), .Q(
        start_reg[332]) );
  DFF \start_reg_reg[333]  ( .D(start_in[332]), .CLK(clk), .RST(rst), .Q(
        start_reg[333]) );
  DFF \start_reg_reg[334]  ( .D(start_in[333]), .CLK(clk), .RST(rst), .Q(
        start_reg[334]) );
  DFF \start_reg_reg[335]  ( .D(start_in[334]), .CLK(clk), .RST(rst), .Q(
        start_reg[335]) );
  DFF \start_reg_reg[336]  ( .D(start_in[335]), .CLK(clk), .RST(rst), .Q(
        start_reg[336]) );
  DFF \start_reg_reg[337]  ( .D(start_in[336]), .CLK(clk), .RST(rst), .Q(
        start_reg[337]) );
  DFF \start_reg_reg[338]  ( .D(start_in[337]), .CLK(clk), .RST(rst), .Q(
        start_reg[338]) );
  DFF \start_reg_reg[339]  ( .D(start_in[338]), .CLK(clk), .RST(rst), .Q(
        start_reg[339]) );
  DFF \start_reg_reg[340]  ( .D(start_in[339]), .CLK(clk), .RST(rst), .Q(
        start_reg[340]) );
  DFF \start_reg_reg[341]  ( .D(start_in[340]), .CLK(clk), .RST(rst), .Q(
        start_reg[341]) );
  DFF \start_reg_reg[342]  ( .D(start_in[341]), .CLK(clk), .RST(rst), .Q(
        start_reg[342]) );
  DFF \start_reg_reg[343]  ( .D(start_in[342]), .CLK(clk), .RST(rst), .Q(
        start_reg[343]) );
  DFF \start_reg_reg[344]  ( .D(start_in[343]), .CLK(clk), .RST(rst), .Q(
        start_reg[344]) );
  DFF \start_reg_reg[345]  ( .D(start_in[344]), .CLK(clk), .RST(rst), .Q(
        start_reg[345]) );
  DFF \start_reg_reg[346]  ( .D(start_in[345]), .CLK(clk), .RST(rst), .Q(
        start_reg[346]) );
  DFF \start_reg_reg[347]  ( .D(start_in[346]), .CLK(clk), .RST(rst), .Q(
        start_reg[347]) );
  DFF \start_reg_reg[348]  ( .D(start_in[347]), .CLK(clk), .RST(rst), .Q(
        start_reg[348]) );
  DFF \start_reg_reg[349]  ( .D(start_in[348]), .CLK(clk), .RST(rst), .Q(
        start_reg[349]) );
  DFF \start_reg_reg[350]  ( .D(start_in[349]), .CLK(clk), .RST(rst), .Q(
        start_reg[350]) );
  DFF \start_reg_reg[351]  ( .D(start_in[350]), .CLK(clk), .RST(rst), .Q(
        start_reg[351]) );
  DFF \start_reg_reg[352]  ( .D(start_in[351]), .CLK(clk), .RST(rst), .Q(
        start_reg[352]) );
  DFF \start_reg_reg[353]  ( .D(start_in[352]), .CLK(clk), .RST(rst), .Q(
        start_reg[353]) );
  DFF \start_reg_reg[354]  ( .D(start_in[353]), .CLK(clk), .RST(rst), .Q(
        start_reg[354]) );
  DFF \start_reg_reg[355]  ( .D(start_in[354]), .CLK(clk), .RST(rst), .Q(
        start_reg[355]) );
  DFF \start_reg_reg[356]  ( .D(start_in[355]), .CLK(clk), .RST(rst), .Q(
        start_reg[356]) );
  DFF \start_reg_reg[357]  ( .D(start_in[356]), .CLK(clk), .RST(rst), .Q(
        start_reg[357]) );
  DFF \start_reg_reg[358]  ( .D(start_in[357]), .CLK(clk), .RST(rst), .Q(
        start_reg[358]) );
  DFF \start_reg_reg[359]  ( .D(start_in[358]), .CLK(clk), .RST(rst), .Q(
        start_reg[359]) );
  DFF \start_reg_reg[360]  ( .D(start_in[359]), .CLK(clk), .RST(rst), .Q(
        start_reg[360]) );
  DFF \start_reg_reg[361]  ( .D(start_in[360]), .CLK(clk), .RST(rst), .Q(
        start_reg[361]) );
  DFF \start_reg_reg[362]  ( .D(start_in[361]), .CLK(clk), .RST(rst), .Q(
        start_reg[362]) );
  DFF \start_reg_reg[363]  ( .D(start_in[362]), .CLK(clk), .RST(rst), .Q(
        start_reg[363]) );
  DFF \start_reg_reg[364]  ( .D(start_in[363]), .CLK(clk), .RST(rst), .Q(
        start_reg[364]) );
  DFF \start_reg_reg[365]  ( .D(start_in[364]), .CLK(clk), .RST(rst), .Q(
        start_reg[365]) );
  DFF \start_reg_reg[366]  ( .D(start_in[365]), .CLK(clk), .RST(rst), .Q(
        start_reg[366]) );
  DFF \start_reg_reg[367]  ( .D(start_in[366]), .CLK(clk), .RST(rst), .Q(
        start_reg[367]) );
  DFF \start_reg_reg[368]  ( .D(start_in[367]), .CLK(clk), .RST(rst), .Q(
        start_reg[368]) );
  DFF \start_reg_reg[369]  ( .D(start_in[368]), .CLK(clk), .RST(rst), .Q(
        start_reg[369]) );
  DFF \start_reg_reg[370]  ( .D(start_in[369]), .CLK(clk), .RST(rst), .Q(
        start_reg[370]) );
  DFF \start_reg_reg[371]  ( .D(start_in[370]), .CLK(clk), .RST(rst), .Q(
        start_reg[371]) );
  DFF \start_reg_reg[372]  ( .D(start_in[371]), .CLK(clk), .RST(rst), .Q(
        start_reg[372]) );
  DFF \start_reg_reg[373]  ( .D(start_in[372]), .CLK(clk), .RST(rst), .Q(
        start_reg[373]) );
  DFF \start_reg_reg[374]  ( .D(start_in[373]), .CLK(clk), .RST(rst), .Q(
        start_reg[374]) );
  DFF \start_reg_reg[375]  ( .D(start_in[374]), .CLK(clk), .RST(rst), .Q(
        start_reg[375]) );
  DFF \start_reg_reg[376]  ( .D(start_in[375]), .CLK(clk), .RST(rst), .Q(
        start_reg[376]) );
  DFF \start_reg_reg[377]  ( .D(start_in[376]), .CLK(clk), .RST(rst), .Q(
        start_reg[377]) );
  DFF \start_reg_reg[378]  ( .D(start_in[377]), .CLK(clk), .RST(rst), .Q(
        start_reg[378]) );
  DFF \start_reg_reg[379]  ( .D(start_in[378]), .CLK(clk), .RST(rst), .Q(
        start_reg[379]) );
  DFF \start_reg_reg[380]  ( .D(start_in[379]), .CLK(clk), .RST(rst), .Q(
        start_reg[380]) );
  DFF \start_reg_reg[381]  ( .D(start_in[380]), .CLK(clk), .RST(rst), .Q(
        start_reg[381]) );
  DFF \start_reg_reg[382]  ( .D(start_in[381]), .CLK(clk), .RST(rst), .Q(
        start_reg[382]) );
  DFF \start_reg_reg[383]  ( .D(start_in[382]), .CLK(clk), .RST(rst), .Q(
        start_reg[383]) );
  DFF \start_reg_reg[384]  ( .D(start_in[383]), .CLK(clk), .RST(rst), .Q(
        start_reg[384]) );
  DFF \start_reg_reg[385]  ( .D(start_in[384]), .CLK(clk), .RST(rst), .Q(
        start_reg[385]) );
  DFF \start_reg_reg[386]  ( .D(start_in[385]), .CLK(clk), .RST(rst), .Q(
        start_reg[386]) );
  DFF \start_reg_reg[387]  ( .D(start_in[386]), .CLK(clk), .RST(rst), .Q(
        start_reg[387]) );
  DFF \start_reg_reg[388]  ( .D(start_in[387]), .CLK(clk), .RST(rst), .Q(
        start_reg[388]) );
  DFF \start_reg_reg[389]  ( .D(start_in[388]), .CLK(clk), .RST(rst), .Q(
        start_reg[389]) );
  DFF \start_reg_reg[390]  ( .D(start_in[389]), .CLK(clk), .RST(rst), .Q(
        start_reg[390]) );
  DFF \start_reg_reg[391]  ( .D(start_in[390]), .CLK(clk), .RST(rst), .Q(
        start_reg[391]) );
  DFF \start_reg_reg[392]  ( .D(start_in[391]), .CLK(clk), .RST(rst), .Q(
        start_reg[392]) );
  DFF \start_reg_reg[393]  ( .D(start_in[392]), .CLK(clk), .RST(rst), .Q(
        start_reg[393]) );
  DFF \start_reg_reg[394]  ( .D(start_in[393]), .CLK(clk), .RST(rst), .Q(
        start_reg[394]) );
  DFF \start_reg_reg[395]  ( .D(start_in[394]), .CLK(clk), .RST(rst), .Q(
        start_reg[395]) );
  DFF \start_reg_reg[396]  ( .D(start_in[395]), .CLK(clk), .RST(rst), .Q(
        start_reg[396]) );
  DFF \start_reg_reg[397]  ( .D(start_in[396]), .CLK(clk), .RST(rst), .Q(
        start_reg[397]) );
  DFF \start_reg_reg[398]  ( .D(start_in[397]), .CLK(clk), .RST(rst), .Q(
        start_reg[398]) );
  DFF \start_reg_reg[399]  ( .D(start_in[398]), .CLK(clk), .RST(rst), .Q(
        start_reg[399]) );
  DFF \start_reg_reg[400]  ( .D(start_in[399]), .CLK(clk), .RST(rst), .Q(
        start_reg[400]) );
  DFF \start_reg_reg[401]  ( .D(start_in[400]), .CLK(clk), .RST(rst), .Q(
        start_reg[401]) );
  DFF \start_reg_reg[402]  ( .D(start_in[401]), .CLK(clk), .RST(rst), .Q(
        start_reg[402]) );
  DFF \start_reg_reg[403]  ( .D(start_in[402]), .CLK(clk), .RST(rst), .Q(
        start_reg[403]) );
  DFF \start_reg_reg[404]  ( .D(start_in[403]), .CLK(clk), .RST(rst), .Q(
        start_reg[404]) );
  DFF \start_reg_reg[405]  ( .D(start_in[404]), .CLK(clk), .RST(rst), .Q(
        start_reg[405]) );
  DFF \start_reg_reg[406]  ( .D(start_in[405]), .CLK(clk), .RST(rst), .Q(
        start_reg[406]) );
  DFF \start_reg_reg[407]  ( .D(start_in[406]), .CLK(clk), .RST(rst), .Q(
        start_reg[407]) );
  DFF \start_reg_reg[408]  ( .D(start_in[407]), .CLK(clk), .RST(rst), .Q(
        start_reg[408]) );
  DFF \start_reg_reg[409]  ( .D(start_in[408]), .CLK(clk), .RST(rst), .Q(
        start_reg[409]) );
  DFF \start_reg_reg[410]  ( .D(start_in[409]), .CLK(clk), .RST(rst), .Q(
        start_reg[410]) );
  DFF \start_reg_reg[411]  ( .D(start_in[410]), .CLK(clk), .RST(rst), .Q(
        start_reg[411]) );
  DFF \start_reg_reg[412]  ( .D(start_in[411]), .CLK(clk), .RST(rst), .Q(
        start_reg[412]) );
  DFF \start_reg_reg[413]  ( .D(start_in[412]), .CLK(clk), .RST(rst), .Q(
        start_reg[413]) );
  DFF \start_reg_reg[414]  ( .D(start_in[413]), .CLK(clk), .RST(rst), .Q(
        start_reg[414]) );
  DFF \start_reg_reg[415]  ( .D(start_in[414]), .CLK(clk), .RST(rst), .Q(
        start_reg[415]) );
  DFF \start_reg_reg[416]  ( .D(start_in[415]), .CLK(clk), .RST(rst), .Q(
        start_reg[416]) );
  DFF \start_reg_reg[417]  ( .D(start_in[416]), .CLK(clk), .RST(rst), .Q(
        start_reg[417]) );
  DFF \start_reg_reg[418]  ( .D(start_in[417]), .CLK(clk), .RST(rst), .Q(
        start_reg[418]) );
  DFF \start_reg_reg[419]  ( .D(start_in[418]), .CLK(clk), .RST(rst), .Q(
        start_reg[419]) );
  DFF \start_reg_reg[420]  ( .D(start_in[419]), .CLK(clk), .RST(rst), .Q(
        start_reg[420]) );
  DFF \start_reg_reg[421]  ( .D(start_in[420]), .CLK(clk), .RST(rst), .Q(
        start_reg[421]) );
  DFF \start_reg_reg[422]  ( .D(start_in[421]), .CLK(clk), .RST(rst), .Q(
        start_reg[422]) );
  DFF \start_reg_reg[423]  ( .D(start_in[422]), .CLK(clk), .RST(rst), .Q(
        start_reg[423]) );
  DFF \start_reg_reg[424]  ( .D(start_in[423]), .CLK(clk), .RST(rst), .Q(
        start_reg[424]) );
  DFF \start_reg_reg[425]  ( .D(start_in[424]), .CLK(clk), .RST(rst), .Q(
        start_reg[425]) );
  DFF \start_reg_reg[426]  ( .D(start_in[425]), .CLK(clk), .RST(rst), .Q(
        start_reg[426]) );
  DFF \start_reg_reg[427]  ( .D(start_in[426]), .CLK(clk), .RST(rst), .Q(
        start_reg[427]) );
  DFF \start_reg_reg[428]  ( .D(start_in[427]), .CLK(clk), .RST(rst), .Q(
        start_reg[428]) );
  DFF \start_reg_reg[429]  ( .D(start_in[428]), .CLK(clk), .RST(rst), .Q(
        start_reg[429]) );
  DFF \start_reg_reg[430]  ( .D(start_in[429]), .CLK(clk), .RST(rst), .Q(
        start_reg[430]) );
  DFF \start_reg_reg[431]  ( .D(start_in[430]), .CLK(clk), .RST(rst), .Q(
        start_reg[431]) );
  DFF \start_reg_reg[432]  ( .D(start_in[431]), .CLK(clk), .RST(rst), .Q(
        start_reg[432]) );
  DFF \start_reg_reg[433]  ( .D(start_in[432]), .CLK(clk), .RST(rst), .Q(
        start_reg[433]) );
  DFF \start_reg_reg[434]  ( .D(start_in[433]), .CLK(clk), .RST(rst), .Q(
        start_reg[434]) );
  DFF \start_reg_reg[435]  ( .D(start_in[434]), .CLK(clk), .RST(rst), .Q(
        start_reg[435]) );
  DFF \start_reg_reg[436]  ( .D(start_in[435]), .CLK(clk), .RST(rst), .Q(
        start_reg[436]) );
  DFF \start_reg_reg[437]  ( .D(start_in[436]), .CLK(clk), .RST(rst), .Q(
        start_reg[437]) );
  DFF \start_reg_reg[438]  ( .D(start_in[437]), .CLK(clk), .RST(rst), .Q(
        start_reg[438]) );
  DFF \start_reg_reg[439]  ( .D(start_in[438]), .CLK(clk), .RST(rst), .Q(
        start_reg[439]) );
  DFF \start_reg_reg[440]  ( .D(start_in[439]), .CLK(clk), .RST(rst), .Q(
        start_reg[440]) );
  DFF \start_reg_reg[441]  ( .D(start_in[440]), .CLK(clk), .RST(rst), .Q(
        start_reg[441]) );
  DFF \start_reg_reg[442]  ( .D(start_in[441]), .CLK(clk), .RST(rst), .Q(
        start_reg[442]) );
  DFF \start_reg_reg[443]  ( .D(start_in[442]), .CLK(clk), .RST(rst), .Q(
        start_reg[443]) );
  DFF \start_reg_reg[444]  ( .D(start_in[443]), .CLK(clk), .RST(rst), .Q(
        start_reg[444]) );
  DFF \start_reg_reg[445]  ( .D(start_in[444]), .CLK(clk), .RST(rst), .Q(
        start_reg[445]) );
  DFF \start_reg_reg[446]  ( .D(start_in[445]), .CLK(clk), .RST(rst), .Q(
        start_reg[446]) );
  DFF \start_reg_reg[447]  ( .D(start_in[446]), .CLK(clk), .RST(rst), .Q(
        start_reg[447]) );
  DFF \start_reg_reg[448]  ( .D(start_in[447]), .CLK(clk), .RST(rst), .Q(
        start_reg[448]) );
  DFF \start_reg_reg[449]  ( .D(start_in[448]), .CLK(clk), .RST(rst), .Q(
        start_reg[449]) );
  DFF \start_reg_reg[450]  ( .D(start_in[449]), .CLK(clk), .RST(rst), .Q(
        start_reg[450]) );
  DFF \start_reg_reg[451]  ( .D(start_in[450]), .CLK(clk), .RST(rst), .Q(
        start_reg[451]) );
  DFF \start_reg_reg[452]  ( .D(start_in[451]), .CLK(clk), .RST(rst), .Q(
        start_reg[452]) );
  DFF \start_reg_reg[453]  ( .D(start_in[452]), .CLK(clk), .RST(rst), .Q(
        start_reg[453]) );
  DFF \start_reg_reg[454]  ( .D(start_in[453]), .CLK(clk), .RST(rst), .Q(
        start_reg[454]) );
  DFF \start_reg_reg[455]  ( .D(start_in[454]), .CLK(clk), .RST(rst), .Q(
        start_reg[455]) );
  DFF \start_reg_reg[456]  ( .D(start_in[455]), .CLK(clk), .RST(rst), .Q(
        start_reg[456]) );
  DFF \start_reg_reg[457]  ( .D(start_in[456]), .CLK(clk), .RST(rst), .Q(
        start_reg[457]) );
  DFF \start_reg_reg[458]  ( .D(start_in[457]), .CLK(clk), .RST(rst), .Q(
        start_reg[458]) );
  DFF \start_reg_reg[459]  ( .D(start_in[458]), .CLK(clk), .RST(rst), .Q(
        start_reg[459]) );
  DFF \start_reg_reg[460]  ( .D(start_in[459]), .CLK(clk), .RST(rst), .Q(
        start_reg[460]) );
  DFF \start_reg_reg[461]  ( .D(start_in[460]), .CLK(clk), .RST(rst), .Q(
        start_reg[461]) );
  DFF \start_reg_reg[462]  ( .D(start_in[461]), .CLK(clk), .RST(rst), .Q(
        start_reg[462]) );
  DFF \start_reg_reg[463]  ( .D(start_in[462]), .CLK(clk), .RST(rst), .Q(
        start_reg[463]) );
  DFF \start_reg_reg[464]  ( .D(start_in[463]), .CLK(clk), .RST(rst), .Q(
        start_reg[464]) );
  DFF \start_reg_reg[465]  ( .D(start_in[464]), .CLK(clk), .RST(rst), .Q(
        start_reg[465]) );
  DFF \start_reg_reg[466]  ( .D(start_in[465]), .CLK(clk), .RST(rst), .Q(
        start_reg[466]) );
  DFF \start_reg_reg[467]  ( .D(start_in[466]), .CLK(clk), .RST(rst), .Q(
        start_reg[467]) );
  DFF \start_reg_reg[468]  ( .D(start_in[467]), .CLK(clk), .RST(rst), .Q(
        start_reg[468]) );
  DFF \start_reg_reg[469]  ( .D(start_in[468]), .CLK(clk), .RST(rst), .Q(
        start_reg[469]) );
  DFF \start_reg_reg[470]  ( .D(start_in[469]), .CLK(clk), .RST(rst), .Q(
        start_reg[470]) );
  DFF \start_reg_reg[471]  ( .D(start_in[470]), .CLK(clk), .RST(rst), .Q(
        start_reg[471]) );
  DFF \start_reg_reg[472]  ( .D(start_in[471]), .CLK(clk), .RST(rst), .Q(
        start_reg[472]) );
  DFF \start_reg_reg[473]  ( .D(start_in[472]), .CLK(clk), .RST(rst), .Q(
        start_reg[473]) );
  DFF \start_reg_reg[474]  ( .D(start_in[473]), .CLK(clk), .RST(rst), .Q(
        start_reg[474]) );
  DFF \start_reg_reg[475]  ( .D(start_in[474]), .CLK(clk), .RST(rst), .Q(
        start_reg[475]) );
  DFF \start_reg_reg[476]  ( .D(start_in[475]), .CLK(clk), .RST(rst), .Q(
        start_reg[476]) );
  DFF \start_reg_reg[477]  ( .D(start_in[476]), .CLK(clk), .RST(rst), .Q(
        start_reg[477]) );
  DFF \start_reg_reg[478]  ( .D(start_in[477]), .CLK(clk), .RST(rst), .Q(
        start_reg[478]) );
  DFF \start_reg_reg[479]  ( .D(start_in[478]), .CLK(clk), .RST(rst), .Q(
        start_reg[479]) );
  DFF \start_reg_reg[480]  ( .D(start_in[479]), .CLK(clk), .RST(rst), .Q(
        start_reg[480]) );
  DFF \start_reg_reg[481]  ( .D(start_in[480]), .CLK(clk), .RST(rst), .Q(
        start_reg[481]) );
  DFF \start_reg_reg[482]  ( .D(start_in[481]), .CLK(clk), .RST(rst), .Q(
        start_reg[482]) );
  DFF \start_reg_reg[483]  ( .D(start_in[482]), .CLK(clk), .RST(rst), .Q(
        start_reg[483]) );
  DFF \start_reg_reg[484]  ( .D(start_in[483]), .CLK(clk), .RST(rst), .Q(
        start_reg[484]) );
  DFF \start_reg_reg[485]  ( .D(start_in[484]), .CLK(clk), .RST(rst), .Q(
        start_reg[485]) );
  DFF \start_reg_reg[486]  ( .D(start_in[485]), .CLK(clk), .RST(rst), .Q(
        start_reg[486]) );
  DFF \start_reg_reg[487]  ( .D(start_in[486]), .CLK(clk), .RST(rst), .Q(
        start_reg[487]) );
  DFF \start_reg_reg[488]  ( .D(start_in[487]), .CLK(clk), .RST(rst), .Q(
        start_reg[488]) );
  DFF \start_reg_reg[489]  ( .D(start_in[488]), .CLK(clk), .RST(rst), .Q(
        start_reg[489]) );
  DFF \start_reg_reg[490]  ( .D(start_in[489]), .CLK(clk), .RST(rst), .Q(
        start_reg[490]) );
  DFF \start_reg_reg[491]  ( .D(start_in[490]), .CLK(clk), .RST(rst), .Q(
        start_reg[491]) );
  DFF \start_reg_reg[492]  ( .D(start_in[491]), .CLK(clk), .RST(rst), .Q(
        start_reg[492]) );
  DFF \start_reg_reg[493]  ( .D(start_in[492]), .CLK(clk), .RST(rst), .Q(
        start_reg[493]) );
  DFF \start_reg_reg[494]  ( .D(start_in[493]), .CLK(clk), .RST(rst), .Q(
        start_reg[494]) );
  DFF \start_reg_reg[495]  ( .D(start_in[494]), .CLK(clk), .RST(rst), .Q(
        start_reg[495]) );
  DFF \start_reg_reg[496]  ( .D(start_in[495]), .CLK(clk), .RST(rst), .Q(
        start_reg[496]) );
  DFF \start_reg_reg[497]  ( .D(start_in[496]), .CLK(clk), .RST(rst), .Q(
        start_reg[497]) );
  DFF \start_reg_reg[498]  ( .D(start_in[497]), .CLK(clk), .RST(rst), .Q(
        start_reg[498]) );
  DFF \start_reg_reg[499]  ( .D(start_in[498]), .CLK(clk), .RST(rst), .Q(
        start_reg[499]) );
  DFF \start_reg_reg[500]  ( .D(start_in[499]), .CLK(clk), .RST(rst), .Q(
        start_reg[500]) );
  DFF \start_reg_reg[501]  ( .D(start_in[500]), .CLK(clk), .RST(rst), .Q(
        start_reg[501]) );
  DFF \start_reg_reg[502]  ( .D(start_in[501]), .CLK(clk), .RST(rst), .Q(
        start_reg[502]) );
  DFF \start_reg_reg[503]  ( .D(start_in[502]), .CLK(clk), .RST(rst), .Q(
        start_reg[503]) );
  DFF \start_reg_reg[504]  ( .D(start_in[503]), .CLK(clk), .RST(rst), .Q(
        start_reg[504]) );
  DFF \start_reg_reg[505]  ( .D(start_in[504]), .CLK(clk), .RST(rst), .Q(
        start_reg[505]) );
  DFF \start_reg_reg[506]  ( .D(start_in[505]), .CLK(clk), .RST(rst), .Q(
        start_reg[506]) );
  DFF \start_reg_reg[507]  ( .D(start_in[506]), .CLK(clk), .RST(rst), .Q(
        start_reg[507]) );
  DFF \start_reg_reg[508]  ( .D(start_in[507]), .CLK(clk), .RST(rst), .Q(
        start_reg[508]) );
  DFF \start_reg_reg[509]  ( .D(start_in[508]), .CLK(clk), .RST(rst), .Q(
        start_reg[509]) );
  DFF \start_reg_reg[510]  ( .D(start_in[509]), .CLK(clk), .RST(rst), .Q(
        start_reg[510]) );
  DFF \start_reg_reg[511]  ( .D(start_in[510]), .CLK(clk), .RST(rst), .Q(
        start_reg[511]) );
  DFF \start_reg_reg[512]  ( .D(start_in[511]), .CLK(clk), .RST(rst), .Q(
        start_reg[512]) );
  DFF \start_reg_reg[513]  ( .D(start_in[512]), .CLK(clk), .RST(rst), .Q(
        start_reg[513]) );
  DFF \start_reg_reg[514]  ( .D(start_in[513]), .CLK(clk), .RST(rst), .Q(
        start_reg[514]) );
  DFF \start_reg_reg[515]  ( .D(start_in[514]), .CLK(clk), .RST(rst), .Q(
        start_reg[515]) );
  DFF \start_reg_reg[516]  ( .D(start_in[515]), .CLK(clk), .RST(rst), .Q(
        start_reg[516]) );
  DFF \start_reg_reg[517]  ( .D(start_in[516]), .CLK(clk), .RST(rst), .Q(
        start_reg[517]) );
  DFF \start_reg_reg[518]  ( .D(start_in[517]), .CLK(clk), .RST(rst), .Q(
        start_reg[518]) );
  DFF \start_reg_reg[519]  ( .D(start_in[518]), .CLK(clk), .RST(rst), .Q(
        start_reg[519]) );
  DFF \start_reg_reg[520]  ( .D(start_in[519]), .CLK(clk), .RST(rst), .Q(
        start_reg[520]) );
  DFF \start_reg_reg[521]  ( .D(start_in[520]), .CLK(clk), .RST(rst), .Q(
        start_reg[521]) );
  DFF \start_reg_reg[522]  ( .D(start_in[521]), .CLK(clk), .RST(rst), .Q(
        start_reg[522]) );
  DFF \start_reg_reg[523]  ( .D(start_in[522]), .CLK(clk), .RST(rst), .Q(
        start_reg[523]) );
  DFF \start_reg_reg[524]  ( .D(start_in[523]), .CLK(clk), .RST(rst), .Q(
        start_reg[524]) );
  DFF \start_reg_reg[525]  ( .D(start_in[524]), .CLK(clk), .RST(rst), .Q(
        start_reg[525]) );
  DFF \start_reg_reg[526]  ( .D(start_in[525]), .CLK(clk), .RST(rst), .Q(
        start_reg[526]) );
  DFF \start_reg_reg[527]  ( .D(start_in[526]), .CLK(clk), .RST(rst), .Q(
        start_reg[527]) );
  DFF \start_reg_reg[528]  ( .D(start_in[527]), .CLK(clk), .RST(rst), .Q(
        start_reg[528]) );
  DFF \start_reg_reg[529]  ( .D(start_in[528]), .CLK(clk), .RST(rst), .Q(
        start_reg[529]) );
  DFF \start_reg_reg[530]  ( .D(start_in[529]), .CLK(clk), .RST(rst), .Q(
        start_reg[530]) );
  DFF \start_reg_reg[531]  ( .D(start_in[530]), .CLK(clk), .RST(rst), .Q(
        start_reg[531]) );
  DFF \start_reg_reg[532]  ( .D(start_in[531]), .CLK(clk), .RST(rst), .Q(
        start_reg[532]) );
  DFF \start_reg_reg[533]  ( .D(start_in[532]), .CLK(clk), .RST(rst), .Q(
        start_reg[533]) );
  DFF \start_reg_reg[534]  ( .D(start_in[533]), .CLK(clk), .RST(rst), .Q(
        start_reg[534]) );
  DFF \start_reg_reg[535]  ( .D(start_in[534]), .CLK(clk), .RST(rst), .Q(
        start_reg[535]) );
  DFF \start_reg_reg[536]  ( .D(start_in[535]), .CLK(clk), .RST(rst), .Q(
        start_reg[536]) );
  DFF \start_reg_reg[537]  ( .D(start_in[536]), .CLK(clk), .RST(rst), .Q(
        start_reg[537]) );
  DFF \start_reg_reg[538]  ( .D(start_in[537]), .CLK(clk), .RST(rst), .Q(
        start_reg[538]) );
  DFF \start_reg_reg[539]  ( .D(start_in[538]), .CLK(clk), .RST(rst), .Q(
        start_reg[539]) );
  DFF \start_reg_reg[540]  ( .D(start_in[539]), .CLK(clk), .RST(rst), .Q(
        start_reg[540]) );
  DFF \start_reg_reg[541]  ( .D(start_in[540]), .CLK(clk), .RST(rst), .Q(
        start_reg[541]) );
  DFF \start_reg_reg[542]  ( .D(start_in[541]), .CLK(clk), .RST(rst), .Q(
        start_reg[542]) );
  DFF \start_reg_reg[543]  ( .D(start_in[542]), .CLK(clk), .RST(rst), .Q(
        start_reg[543]) );
  DFF \start_reg_reg[544]  ( .D(start_in[543]), .CLK(clk), .RST(rst), .Q(
        start_reg[544]) );
  DFF \start_reg_reg[545]  ( .D(start_in[544]), .CLK(clk), .RST(rst), .Q(
        start_reg[545]) );
  DFF \start_reg_reg[546]  ( .D(start_in[545]), .CLK(clk), .RST(rst), .Q(
        start_reg[546]) );
  DFF \start_reg_reg[547]  ( .D(start_in[546]), .CLK(clk), .RST(rst), .Q(
        start_reg[547]) );
  DFF \start_reg_reg[548]  ( .D(start_in[547]), .CLK(clk), .RST(rst), .Q(
        start_reg[548]) );
  DFF \start_reg_reg[549]  ( .D(start_in[548]), .CLK(clk), .RST(rst), .Q(
        start_reg[549]) );
  DFF \start_reg_reg[550]  ( .D(start_in[549]), .CLK(clk), .RST(rst), .Q(
        start_reg[550]) );
  DFF \start_reg_reg[551]  ( .D(start_in[550]), .CLK(clk), .RST(rst), .Q(
        start_reg[551]) );
  DFF \start_reg_reg[552]  ( .D(start_in[551]), .CLK(clk), .RST(rst), .Q(
        start_reg[552]) );
  DFF \start_reg_reg[553]  ( .D(start_in[552]), .CLK(clk), .RST(rst), .Q(
        start_reg[553]) );
  DFF \start_reg_reg[554]  ( .D(start_in[553]), .CLK(clk), .RST(rst), .Q(
        start_reg[554]) );
  DFF \start_reg_reg[555]  ( .D(start_in[554]), .CLK(clk), .RST(rst), .Q(
        start_reg[555]) );
  DFF \start_reg_reg[556]  ( .D(start_in[555]), .CLK(clk), .RST(rst), .Q(
        start_reg[556]) );
  DFF \start_reg_reg[557]  ( .D(start_in[556]), .CLK(clk), .RST(rst), .Q(
        start_reg[557]) );
  DFF \start_reg_reg[558]  ( .D(start_in[557]), .CLK(clk), .RST(rst), .Q(
        start_reg[558]) );
  DFF \start_reg_reg[559]  ( .D(start_in[558]), .CLK(clk), .RST(rst), .Q(
        start_reg[559]) );
  DFF \start_reg_reg[560]  ( .D(start_in[559]), .CLK(clk), .RST(rst), .Q(
        start_reg[560]) );
  DFF \start_reg_reg[561]  ( .D(start_in[560]), .CLK(clk), .RST(rst), .Q(
        start_reg[561]) );
  DFF \start_reg_reg[562]  ( .D(start_in[561]), .CLK(clk), .RST(rst), .Q(
        start_reg[562]) );
  DFF \start_reg_reg[563]  ( .D(start_in[562]), .CLK(clk), .RST(rst), .Q(
        start_reg[563]) );
  DFF \start_reg_reg[564]  ( .D(start_in[563]), .CLK(clk), .RST(rst), .Q(
        start_reg[564]) );
  DFF \start_reg_reg[565]  ( .D(start_in[564]), .CLK(clk), .RST(rst), .Q(
        start_reg[565]) );
  DFF \start_reg_reg[566]  ( .D(start_in[565]), .CLK(clk), .RST(rst), .Q(
        start_reg[566]) );
  DFF \start_reg_reg[567]  ( .D(start_in[566]), .CLK(clk), .RST(rst), .Q(
        start_reg[567]) );
  DFF \start_reg_reg[568]  ( .D(start_in[567]), .CLK(clk), .RST(rst), .Q(
        start_reg[568]) );
  DFF \start_reg_reg[569]  ( .D(start_in[568]), .CLK(clk), .RST(rst), .Q(
        start_reg[569]) );
  DFF \start_reg_reg[570]  ( .D(start_in[569]), .CLK(clk), .RST(rst), .Q(
        start_reg[570]) );
  DFF \start_reg_reg[571]  ( .D(start_in[570]), .CLK(clk), .RST(rst), .Q(
        start_reg[571]) );
  DFF \start_reg_reg[572]  ( .D(start_in[571]), .CLK(clk), .RST(rst), .Q(
        start_reg[572]) );
  DFF \start_reg_reg[573]  ( .D(start_in[572]), .CLK(clk), .RST(rst), .Q(
        start_reg[573]) );
  DFF \start_reg_reg[574]  ( .D(start_in[573]), .CLK(clk), .RST(rst), .Q(
        start_reg[574]) );
  DFF \start_reg_reg[575]  ( .D(start_in[574]), .CLK(clk), .RST(rst), .Q(
        start_reg[575]) );
  DFF \start_reg_reg[576]  ( .D(start_in[575]), .CLK(clk), .RST(rst), .Q(
        start_reg[576]) );
  DFF \start_reg_reg[577]  ( .D(start_in[576]), .CLK(clk), .RST(rst), .Q(
        start_reg[577]) );
  DFF \start_reg_reg[578]  ( .D(start_in[577]), .CLK(clk), .RST(rst), .Q(
        start_reg[578]) );
  DFF \start_reg_reg[579]  ( .D(start_in[578]), .CLK(clk), .RST(rst), .Q(
        start_reg[579]) );
  DFF \start_reg_reg[580]  ( .D(start_in[579]), .CLK(clk), .RST(rst), .Q(
        start_reg[580]) );
  DFF \start_reg_reg[581]  ( .D(start_in[580]), .CLK(clk), .RST(rst), .Q(
        start_reg[581]) );
  DFF \start_reg_reg[582]  ( .D(start_in[581]), .CLK(clk), .RST(rst), .Q(
        start_reg[582]) );
  DFF \start_reg_reg[583]  ( .D(start_in[582]), .CLK(clk), .RST(rst), .Q(
        start_reg[583]) );
  DFF \start_reg_reg[584]  ( .D(start_in[583]), .CLK(clk), .RST(rst), .Q(
        start_reg[584]) );
  DFF \start_reg_reg[585]  ( .D(start_in[584]), .CLK(clk), .RST(rst), .Q(
        start_reg[585]) );
  DFF \start_reg_reg[586]  ( .D(start_in[585]), .CLK(clk), .RST(rst), .Q(
        start_reg[586]) );
  DFF \start_reg_reg[587]  ( .D(start_in[586]), .CLK(clk), .RST(rst), .Q(
        start_reg[587]) );
  DFF \start_reg_reg[588]  ( .D(start_in[587]), .CLK(clk), .RST(rst), .Q(
        start_reg[588]) );
  DFF \start_reg_reg[589]  ( .D(start_in[588]), .CLK(clk), .RST(rst), .Q(
        start_reg[589]) );
  DFF \start_reg_reg[590]  ( .D(start_in[589]), .CLK(clk), .RST(rst), .Q(
        start_reg[590]) );
  DFF \start_reg_reg[591]  ( .D(start_in[590]), .CLK(clk), .RST(rst), .Q(
        start_reg[591]) );
  DFF \start_reg_reg[592]  ( .D(start_in[591]), .CLK(clk), .RST(rst), .Q(
        start_reg[592]) );
  DFF \start_reg_reg[593]  ( .D(start_in[592]), .CLK(clk), .RST(rst), .Q(
        start_reg[593]) );
  DFF \start_reg_reg[594]  ( .D(start_in[593]), .CLK(clk), .RST(rst), .Q(
        start_reg[594]) );
  DFF \start_reg_reg[595]  ( .D(start_in[594]), .CLK(clk), .RST(rst), .Q(
        start_reg[595]) );
  DFF \start_reg_reg[596]  ( .D(start_in[595]), .CLK(clk), .RST(rst), .Q(
        start_reg[596]) );
  DFF \start_reg_reg[597]  ( .D(start_in[596]), .CLK(clk), .RST(rst), .Q(
        start_reg[597]) );
  DFF \start_reg_reg[598]  ( .D(start_in[597]), .CLK(clk), .RST(rst), .Q(
        start_reg[598]) );
  DFF \start_reg_reg[599]  ( .D(start_in[598]), .CLK(clk), .RST(rst), .Q(
        start_reg[599]) );
  DFF \start_reg_reg[600]  ( .D(start_in[599]), .CLK(clk), .RST(rst), .Q(
        start_reg[600]) );
  DFF \start_reg_reg[601]  ( .D(start_in[600]), .CLK(clk), .RST(rst), .Q(
        start_reg[601]) );
  DFF \start_reg_reg[602]  ( .D(start_in[601]), .CLK(clk), .RST(rst), .Q(
        start_reg[602]) );
  DFF \start_reg_reg[603]  ( .D(start_in[602]), .CLK(clk), .RST(rst), .Q(
        start_reg[603]) );
  DFF \start_reg_reg[604]  ( .D(start_in[603]), .CLK(clk), .RST(rst), .Q(
        start_reg[604]) );
  DFF \start_reg_reg[605]  ( .D(start_in[604]), .CLK(clk), .RST(rst), .Q(
        start_reg[605]) );
  DFF \start_reg_reg[606]  ( .D(start_in[605]), .CLK(clk), .RST(rst), .Q(
        start_reg[606]) );
  DFF \start_reg_reg[607]  ( .D(start_in[606]), .CLK(clk), .RST(rst), .Q(
        start_reg[607]) );
  DFF \start_reg_reg[608]  ( .D(start_in[607]), .CLK(clk), .RST(rst), .Q(
        start_reg[608]) );
  DFF \start_reg_reg[609]  ( .D(start_in[608]), .CLK(clk), .RST(rst), .Q(
        start_reg[609]) );
  DFF \start_reg_reg[610]  ( .D(start_in[609]), .CLK(clk), .RST(rst), .Q(
        start_reg[610]) );
  DFF \start_reg_reg[611]  ( .D(start_in[610]), .CLK(clk), .RST(rst), .Q(
        start_reg[611]) );
  DFF \start_reg_reg[612]  ( .D(start_in[611]), .CLK(clk), .RST(rst), .Q(
        start_reg[612]) );
  DFF \start_reg_reg[613]  ( .D(start_in[612]), .CLK(clk), .RST(rst), .Q(
        start_reg[613]) );
  DFF \start_reg_reg[614]  ( .D(start_in[613]), .CLK(clk), .RST(rst), .Q(
        start_reg[614]) );
  DFF \start_reg_reg[615]  ( .D(start_in[614]), .CLK(clk), .RST(rst), .Q(
        start_reg[615]) );
  DFF \start_reg_reg[616]  ( .D(start_in[615]), .CLK(clk), .RST(rst), .Q(
        start_reg[616]) );
  DFF \start_reg_reg[617]  ( .D(start_in[616]), .CLK(clk), .RST(rst), .Q(
        start_reg[617]) );
  DFF \start_reg_reg[618]  ( .D(start_in[617]), .CLK(clk), .RST(rst), .Q(
        start_reg[618]) );
  DFF \start_reg_reg[619]  ( .D(start_in[618]), .CLK(clk), .RST(rst), .Q(
        start_reg[619]) );
  DFF \start_reg_reg[620]  ( .D(start_in[619]), .CLK(clk), .RST(rst), .Q(
        start_reg[620]) );
  DFF \start_reg_reg[621]  ( .D(start_in[620]), .CLK(clk), .RST(rst), .Q(
        start_reg[621]) );
  DFF \start_reg_reg[622]  ( .D(start_in[621]), .CLK(clk), .RST(rst), .Q(
        start_reg[622]) );
  DFF \start_reg_reg[623]  ( .D(start_in[622]), .CLK(clk), .RST(rst), .Q(
        start_reg[623]) );
  DFF \start_reg_reg[624]  ( .D(start_in[623]), .CLK(clk), .RST(rst), .Q(
        start_reg[624]) );
  DFF \start_reg_reg[625]  ( .D(start_in[624]), .CLK(clk), .RST(rst), .Q(
        start_reg[625]) );
  DFF \start_reg_reg[626]  ( .D(start_in[625]), .CLK(clk), .RST(rst), .Q(
        start_reg[626]) );
  DFF \start_reg_reg[627]  ( .D(start_in[626]), .CLK(clk), .RST(rst), .Q(
        start_reg[627]) );
  DFF \start_reg_reg[628]  ( .D(start_in[627]), .CLK(clk), .RST(rst), .Q(
        start_reg[628]) );
  DFF \start_reg_reg[629]  ( .D(start_in[628]), .CLK(clk), .RST(rst), .Q(
        start_reg[629]) );
  DFF \start_reg_reg[630]  ( .D(start_in[629]), .CLK(clk), .RST(rst), .Q(
        start_reg[630]) );
  DFF \start_reg_reg[631]  ( .D(start_in[630]), .CLK(clk), .RST(rst), .Q(
        start_reg[631]) );
  DFF \start_reg_reg[632]  ( .D(start_in[631]), .CLK(clk), .RST(rst), .Q(
        start_reg[632]) );
  DFF \start_reg_reg[633]  ( .D(start_in[632]), .CLK(clk), .RST(rst), .Q(
        start_reg[633]) );
  DFF \start_reg_reg[634]  ( .D(start_in[633]), .CLK(clk), .RST(rst), .Q(
        start_reg[634]) );
  DFF \start_reg_reg[635]  ( .D(start_in[634]), .CLK(clk), .RST(rst), .Q(
        start_reg[635]) );
  DFF \start_reg_reg[636]  ( .D(start_in[635]), .CLK(clk), .RST(rst), .Q(
        start_reg[636]) );
  DFF \start_reg_reg[637]  ( .D(start_in[636]), .CLK(clk), .RST(rst), .Q(
        start_reg[637]) );
  DFF \start_reg_reg[638]  ( .D(start_in[637]), .CLK(clk), .RST(rst), .Q(
        start_reg[638]) );
  DFF \start_reg_reg[639]  ( .D(start_in[638]), .CLK(clk), .RST(rst), .Q(
        start_reg[639]) );
  DFF \start_reg_reg[640]  ( .D(start_in[639]), .CLK(clk), .RST(rst), .Q(
        start_reg[640]) );
  DFF \start_reg_reg[641]  ( .D(start_in[640]), .CLK(clk), .RST(rst), .Q(
        start_reg[641]) );
  DFF \start_reg_reg[642]  ( .D(start_in[641]), .CLK(clk), .RST(rst), .Q(
        start_reg[642]) );
  DFF \start_reg_reg[643]  ( .D(start_in[642]), .CLK(clk), .RST(rst), .Q(
        start_reg[643]) );
  DFF \start_reg_reg[644]  ( .D(start_in[643]), .CLK(clk), .RST(rst), .Q(
        start_reg[644]) );
  DFF \start_reg_reg[645]  ( .D(start_in[644]), .CLK(clk), .RST(rst), .Q(
        start_reg[645]) );
  DFF \start_reg_reg[646]  ( .D(start_in[645]), .CLK(clk), .RST(rst), .Q(
        start_reg[646]) );
  DFF \start_reg_reg[647]  ( .D(start_in[646]), .CLK(clk), .RST(rst), .Q(
        start_reg[647]) );
  DFF \start_reg_reg[648]  ( .D(start_in[647]), .CLK(clk), .RST(rst), .Q(
        start_reg[648]) );
  DFF \start_reg_reg[649]  ( .D(start_in[648]), .CLK(clk), .RST(rst), .Q(
        start_reg[649]) );
  DFF \start_reg_reg[650]  ( .D(start_in[649]), .CLK(clk), .RST(rst), .Q(
        start_reg[650]) );
  DFF \start_reg_reg[651]  ( .D(start_in[650]), .CLK(clk), .RST(rst), .Q(
        start_reg[651]) );
  DFF \start_reg_reg[652]  ( .D(start_in[651]), .CLK(clk), .RST(rst), .Q(
        start_reg[652]) );
  DFF \start_reg_reg[653]  ( .D(start_in[652]), .CLK(clk), .RST(rst), .Q(
        start_reg[653]) );
  DFF \start_reg_reg[654]  ( .D(start_in[653]), .CLK(clk), .RST(rst), .Q(
        start_reg[654]) );
  DFF \start_reg_reg[655]  ( .D(start_in[654]), .CLK(clk), .RST(rst), .Q(
        start_reg[655]) );
  DFF \start_reg_reg[656]  ( .D(start_in[655]), .CLK(clk), .RST(rst), .Q(
        start_reg[656]) );
  DFF \start_reg_reg[657]  ( .D(start_in[656]), .CLK(clk), .RST(rst), .Q(
        start_reg[657]) );
  DFF \start_reg_reg[658]  ( .D(start_in[657]), .CLK(clk), .RST(rst), .Q(
        start_reg[658]) );
  DFF \start_reg_reg[659]  ( .D(start_in[658]), .CLK(clk), .RST(rst), .Q(
        start_reg[659]) );
  DFF \start_reg_reg[660]  ( .D(start_in[659]), .CLK(clk), .RST(rst), .Q(
        start_reg[660]) );
  DFF \start_reg_reg[661]  ( .D(start_in[660]), .CLK(clk), .RST(rst), .Q(
        start_reg[661]) );
  DFF \start_reg_reg[662]  ( .D(start_in[661]), .CLK(clk), .RST(rst), .Q(
        start_reg[662]) );
  DFF \start_reg_reg[663]  ( .D(start_in[662]), .CLK(clk), .RST(rst), .Q(
        start_reg[663]) );
  DFF \start_reg_reg[664]  ( .D(start_in[663]), .CLK(clk), .RST(rst), .Q(
        start_reg[664]) );
  DFF \start_reg_reg[665]  ( .D(start_in[664]), .CLK(clk), .RST(rst), .Q(
        start_reg[665]) );
  DFF \start_reg_reg[666]  ( .D(start_in[665]), .CLK(clk), .RST(rst), .Q(
        start_reg[666]) );
  DFF \start_reg_reg[667]  ( .D(start_in[666]), .CLK(clk), .RST(rst), .Q(
        start_reg[667]) );
  DFF \start_reg_reg[668]  ( .D(start_in[667]), .CLK(clk), .RST(rst), .Q(
        start_reg[668]) );
  DFF \start_reg_reg[669]  ( .D(start_in[668]), .CLK(clk), .RST(rst), .Q(
        start_reg[669]) );
  DFF \start_reg_reg[670]  ( .D(start_in[669]), .CLK(clk), .RST(rst), .Q(
        start_reg[670]) );
  DFF \start_reg_reg[671]  ( .D(start_in[670]), .CLK(clk), .RST(rst), .Q(
        start_reg[671]) );
  DFF \start_reg_reg[672]  ( .D(start_in[671]), .CLK(clk), .RST(rst), .Q(
        start_reg[672]) );
  DFF \start_reg_reg[673]  ( .D(start_in[672]), .CLK(clk), .RST(rst), .Q(
        start_reg[673]) );
  DFF \start_reg_reg[674]  ( .D(start_in[673]), .CLK(clk), .RST(rst), .Q(
        start_reg[674]) );
  DFF \start_reg_reg[675]  ( .D(start_in[674]), .CLK(clk), .RST(rst), .Q(
        start_reg[675]) );
  DFF \start_reg_reg[676]  ( .D(start_in[675]), .CLK(clk), .RST(rst), .Q(
        start_reg[676]) );
  DFF \start_reg_reg[677]  ( .D(start_in[676]), .CLK(clk), .RST(rst), .Q(
        start_reg[677]) );
  DFF \start_reg_reg[678]  ( .D(start_in[677]), .CLK(clk), .RST(rst), .Q(
        start_reg[678]) );
  DFF \start_reg_reg[679]  ( .D(start_in[678]), .CLK(clk), .RST(rst), .Q(
        start_reg[679]) );
  DFF \start_reg_reg[680]  ( .D(start_in[679]), .CLK(clk), .RST(rst), .Q(
        start_reg[680]) );
  DFF \start_reg_reg[681]  ( .D(start_in[680]), .CLK(clk), .RST(rst), .Q(
        start_reg[681]) );
  DFF \start_reg_reg[682]  ( .D(start_in[681]), .CLK(clk), .RST(rst), .Q(
        start_reg[682]) );
  DFF \start_reg_reg[683]  ( .D(start_in[682]), .CLK(clk), .RST(rst), .Q(
        start_reg[683]) );
  DFF \start_reg_reg[684]  ( .D(start_in[683]), .CLK(clk), .RST(rst), .Q(
        start_reg[684]) );
  DFF \start_reg_reg[685]  ( .D(start_in[684]), .CLK(clk), .RST(rst), .Q(
        start_reg[685]) );
  DFF \start_reg_reg[686]  ( .D(start_in[685]), .CLK(clk), .RST(rst), .Q(
        start_reg[686]) );
  DFF \start_reg_reg[687]  ( .D(start_in[686]), .CLK(clk), .RST(rst), .Q(
        start_reg[687]) );
  DFF \start_reg_reg[688]  ( .D(start_in[687]), .CLK(clk), .RST(rst), .Q(
        start_reg[688]) );
  DFF \start_reg_reg[689]  ( .D(start_in[688]), .CLK(clk), .RST(rst), .Q(
        start_reg[689]) );
  DFF \start_reg_reg[690]  ( .D(start_in[689]), .CLK(clk), .RST(rst), .Q(
        start_reg[690]) );
  DFF \start_reg_reg[691]  ( .D(start_in[690]), .CLK(clk), .RST(rst), .Q(
        start_reg[691]) );
  DFF \start_reg_reg[692]  ( .D(start_in[691]), .CLK(clk), .RST(rst), .Q(
        start_reg[692]) );
  DFF \start_reg_reg[693]  ( .D(start_in[692]), .CLK(clk), .RST(rst), .Q(
        start_reg[693]) );
  DFF \start_reg_reg[694]  ( .D(start_in[693]), .CLK(clk), .RST(rst), .Q(
        start_reg[694]) );
  DFF \start_reg_reg[695]  ( .D(start_in[694]), .CLK(clk), .RST(rst), .Q(
        start_reg[695]) );
  DFF \start_reg_reg[696]  ( .D(start_in[695]), .CLK(clk), .RST(rst), .Q(
        start_reg[696]) );
  DFF \start_reg_reg[697]  ( .D(start_in[696]), .CLK(clk), .RST(rst), .Q(
        start_reg[697]) );
  DFF \start_reg_reg[698]  ( .D(start_in[697]), .CLK(clk), .RST(rst), .Q(
        start_reg[698]) );
  DFF \start_reg_reg[699]  ( .D(start_in[698]), .CLK(clk), .RST(rst), .Q(
        start_reg[699]) );
  DFF \start_reg_reg[700]  ( .D(start_in[699]), .CLK(clk), .RST(rst), .Q(
        start_reg[700]) );
  DFF \start_reg_reg[701]  ( .D(start_in[700]), .CLK(clk), .RST(rst), .Q(
        start_reg[701]) );
  DFF \start_reg_reg[702]  ( .D(start_in[701]), .CLK(clk), .RST(rst), .Q(
        start_reg[702]) );
  DFF \start_reg_reg[703]  ( .D(start_in[702]), .CLK(clk), .RST(rst), .Q(
        start_reg[703]) );
  DFF \start_reg_reg[704]  ( .D(start_in[703]), .CLK(clk), .RST(rst), .Q(
        start_reg[704]) );
  DFF \start_reg_reg[705]  ( .D(start_in[704]), .CLK(clk), .RST(rst), .Q(
        start_reg[705]) );
  DFF \start_reg_reg[706]  ( .D(start_in[705]), .CLK(clk), .RST(rst), .Q(
        start_reg[706]) );
  DFF \start_reg_reg[707]  ( .D(start_in[706]), .CLK(clk), .RST(rst), .Q(
        start_reg[707]) );
  DFF \start_reg_reg[708]  ( .D(start_in[707]), .CLK(clk), .RST(rst), .Q(
        start_reg[708]) );
  DFF \start_reg_reg[709]  ( .D(start_in[708]), .CLK(clk), .RST(rst), .Q(
        start_reg[709]) );
  DFF \start_reg_reg[710]  ( .D(start_in[709]), .CLK(clk), .RST(rst), .Q(
        start_reg[710]) );
  DFF \start_reg_reg[711]  ( .D(start_in[710]), .CLK(clk), .RST(rst), .Q(
        start_reg[711]) );
  DFF \start_reg_reg[712]  ( .D(start_in[711]), .CLK(clk), .RST(rst), .Q(
        start_reg[712]) );
  DFF \start_reg_reg[713]  ( .D(start_in[712]), .CLK(clk), .RST(rst), .Q(
        start_reg[713]) );
  DFF \start_reg_reg[714]  ( .D(start_in[713]), .CLK(clk), .RST(rst), .Q(
        start_reg[714]) );
  DFF \start_reg_reg[715]  ( .D(start_in[714]), .CLK(clk), .RST(rst), .Q(
        start_reg[715]) );
  DFF \start_reg_reg[716]  ( .D(start_in[715]), .CLK(clk), .RST(rst), .Q(
        start_reg[716]) );
  DFF \start_reg_reg[717]  ( .D(start_in[716]), .CLK(clk), .RST(rst), .Q(
        start_reg[717]) );
  DFF \start_reg_reg[718]  ( .D(start_in[717]), .CLK(clk), .RST(rst), .Q(
        start_reg[718]) );
  DFF \start_reg_reg[719]  ( .D(start_in[718]), .CLK(clk), .RST(rst), .Q(
        start_reg[719]) );
  DFF \start_reg_reg[720]  ( .D(start_in[719]), .CLK(clk), .RST(rst), .Q(
        start_reg[720]) );
  DFF \start_reg_reg[721]  ( .D(start_in[720]), .CLK(clk), .RST(rst), .Q(
        start_reg[721]) );
  DFF \start_reg_reg[722]  ( .D(start_in[721]), .CLK(clk), .RST(rst), .Q(
        start_reg[722]) );
  DFF \start_reg_reg[723]  ( .D(start_in[722]), .CLK(clk), .RST(rst), .Q(
        start_reg[723]) );
  DFF \start_reg_reg[724]  ( .D(start_in[723]), .CLK(clk), .RST(rst), .Q(
        start_reg[724]) );
  DFF \start_reg_reg[725]  ( .D(start_in[724]), .CLK(clk), .RST(rst), .Q(
        start_reg[725]) );
  DFF \start_reg_reg[726]  ( .D(start_in[725]), .CLK(clk), .RST(rst), .Q(
        start_reg[726]) );
  DFF \start_reg_reg[727]  ( .D(start_in[726]), .CLK(clk), .RST(rst), .Q(
        start_reg[727]) );
  DFF \start_reg_reg[728]  ( .D(start_in[727]), .CLK(clk), .RST(rst), .Q(
        start_reg[728]) );
  DFF \start_reg_reg[729]  ( .D(start_in[728]), .CLK(clk), .RST(rst), .Q(
        start_reg[729]) );
  DFF \start_reg_reg[730]  ( .D(start_in[729]), .CLK(clk), .RST(rst), .Q(
        start_reg[730]) );
  DFF \start_reg_reg[731]  ( .D(start_in[730]), .CLK(clk), .RST(rst), .Q(
        start_reg[731]) );
  DFF \start_reg_reg[732]  ( .D(start_in[731]), .CLK(clk), .RST(rst), .Q(
        start_reg[732]) );
  DFF \start_reg_reg[733]  ( .D(start_in[732]), .CLK(clk), .RST(rst), .Q(
        start_reg[733]) );
  DFF \start_reg_reg[734]  ( .D(start_in[733]), .CLK(clk), .RST(rst), .Q(
        start_reg[734]) );
  DFF \start_reg_reg[735]  ( .D(start_in[734]), .CLK(clk), .RST(rst), .Q(
        start_reg[735]) );
  DFF \start_reg_reg[736]  ( .D(start_in[735]), .CLK(clk), .RST(rst), .Q(
        start_reg[736]) );
  DFF \start_reg_reg[737]  ( .D(start_in[736]), .CLK(clk), .RST(rst), .Q(
        start_reg[737]) );
  DFF \start_reg_reg[738]  ( .D(start_in[737]), .CLK(clk), .RST(rst), .Q(
        start_reg[738]) );
  DFF \start_reg_reg[739]  ( .D(start_in[738]), .CLK(clk), .RST(rst), .Q(
        start_reg[739]) );
  DFF \start_reg_reg[740]  ( .D(start_in[739]), .CLK(clk), .RST(rst), .Q(
        start_reg[740]) );
  DFF \start_reg_reg[741]  ( .D(start_in[740]), .CLK(clk), .RST(rst), .Q(
        start_reg[741]) );
  DFF \start_reg_reg[742]  ( .D(start_in[741]), .CLK(clk), .RST(rst), .Q(
        start_reg[742]) );
  DFF \start_reg_reg[743]  ( .D(start_in[742]), .CLK(clk), .RST(rst), .Q(
        start_reg[743]) );
  DFF \start_reg_reg[744]  ( .D(start_in[743]), .CLK(clk), .RST(rst), .Q(
        start_reg[744]) );
  DFF \start_reg_reg[745]  ( .D(start_in[744]), .CLK(clk), .RST(rst), .Q(
        start_reg[745]) );
  DFF \start_reg_reg[746]  ( .D(start_in[745]), .CLK(clk), .RST(rst), .Q(
        start_reg[746]) );
  DFF \start_reg_reg[747]  ( .D(start_in[746]), .CLK(clk), .RST(rst), .Q(
        start_reg[747]) );
  DFF \start_reg_reg[748]  ( .D(start_in[747]), .CLK(clk), .RST(rst), .Q(
        start_reg[748]) );
  DFF \start_reg_reg[749]  ( .D(start_in[748]), .CLK(clk), .RST(rst), .Q(
        start_reg[749]) );
  DFF \start_reg_reg[750]  ( .D(start_in[749]), .CLK(clk), .RST(rst), .Q(
        start_reg[750]) );
  DFF \start_reg_reg[751]  ( .D(start_in[750]), .CLK(clk), .RST(rst), .Q(
        start_reg[751]) );
  DFF \start_reg_reg[752]  ( .D(start_in[751]), .CLK(clk), .RST(rst), .Q(
        start_reg[752]) );
  DFF \start_reg_reg[753]  ( .D(start_in[752]), .CLK(clk), .RST(rst), .Q(
        start_reg[753]) );
  DFF \start_reg_reg[754]  ( .D(start_in[753]), .CLK(clk), .RST(rst), .Q(
        start_reg[754]) );
  DFF \start_reg_reg[755]  ( .D(start_in[754]), .CLK(clk), .RST(rst), .Q(
        start_reg[755]) );
  DFF \start_reg_reg[756]  ( .D(start_in[755]), .CLK(clk), .RST(rst), .Q(
        start_reg[756]) );
  DFF \start_reg_reg[757]  ( .D(start_in[756]), .CLK(clk), .RST(rst), .Q(
        start_reg[757]) );
  DFF \start_reg_reg[758]  ( .D(start_in[757]), .CLK(clk), .RST(rst), .Q(
        start_reg[758]) );
  DFF \start_reg_reg[759]  ( .D(start_in[758]), .CLK(clk), .RST(rst), .Q(
        start_reg[759]) );
  DFF \start_reg_reg[760]  ( .D(start_in[759]), .CLK(clk), .RST(rst), .Q(
        start_reg[760]) );
  DFF \start_reg_reg[761]  ( .D(start_in[760]), .CLK(clk), .RST(rst), .Q(
        start_reg[761]) );
  DFF \start_reg_reg[762]  ( .D(start_in[761]), .CLK(clk), .RST(rst), .Q(
        start_reg[762]) );
  DFF \start_reg_reg[763]  ( .D(start_in[762]), .CLK(clk), .RST(rst), .Q(
        start_reg[763]) );
  DFF \start_reg_reg[764]  ( .D(start_in[763]), .CLK(clk), .RST(rst), .Q(
        start_reg[764]) );
  DFF \start_reg_reg[765]  ( .D(start_in[764]), .CLK(clk), .RST(rst), .Q(
        start_reg[765]) );
  DFF \start_reg_reg[766]  ( .D(start_in[765]), .CLK(clk), .RST(rst), .Q(
        start_reg[766]) );
  DFF \start_reg_reg[767]  ( .D(start_in[766]), .CLK(clk), .RST(rst), .Q(
        start_reg[767]) );
  DFF \start_reg_reg[768]  ( .D(start_in[767]), .CLK(clk), .RST(rst), .Q(
        start_reg[768]) );
  DFF \start_reg_reg[769]  ( .D(start_in[768]), .CLK(clk), .RST(rst), .Q(
        start_reg[769]) );
  DFF \start_reg_reg[770]  ( .D(start_in[769]), .CLK(clk), .RST(rst), .Q(
        start_reg[770]) );
  DFF \start_reg_reg[771]  ( .D(start_in[770]), .CLK(clk), .RST(rst), .Q(
        start_reg[771]) );
  DFF \start_reg_reg[772]  ( .D(start_in[771]), .CLK(clk), .RST(rst), .Q(
        start_reg[772]) );
  DFF \start_reg_reg[773]  ( .D(start_in[772]), .CLK(clk), .RST(rst), .Q(
        start_reg[773]) );
  DFF \start_reg_reg[774]  ( .D(start_in[773]), .CLK(clk), .RST(rst), .Q(
        start_reg[774]) );
  DFF \start_reg_reg[775]  ( .D(start_in[774]), .CLK(clk), .RST(rst), .Q(
        start_reg[775]) );
  DFF \start_reg_reg[776]  ( .D(start_in[775]), .CLK(clk), .RST(rst), .Q(
        start_reg[776]) );
  DFF \start_reg_reg[777]  ( .D(start_in[776]), .CLK(clk), .RST(rst), .Q(
        start_reg[777]) );
  DFF \start_reg_reg[778]  ( .D(start_in[777]), .CLK(clk), .RST(rst), .Q(
        start_reg[778]) );
  DFF \start_reg_reg[779]  ( .D(start_in[778]), .CLK(clk), .RST(rst), .Q(
        start_reg[779]) );
  DFF \start_reg_reg[780]  ( .D(start_in[779]), .CLK(clk), .RST(rst), .Q(
        start_reg[780]) );
  DFF \start_reg_reg[781]  ( .D(start_in[780]), .CLK(clk), .RST(rst), .Q(
        start_reg[781]) );
  DFF \start_reg_reg[782]  ( .D(start_in[781]), .CLK(clk), .RST(rst), .Q(
        start_reg[782]) );
  DFF \start_reg_reg[783]  ( .D(start_in[782]), .CLK(clk), .RST(rst), .Q(
        start_reg[783]) );
  DFF \start_reg_reg[784]  ( .D(start_in[783]), .CLK(clk), .RST(rst), .Q(
        start_reg[784]) );
  DFF \start_reg_reg[785]  ( .D(start_in[784]), .CLK(clk), .RST(rst), .Q(
        start_reg[785]) );
  DFF \start_reg_reg[786]  ( .D(start_in[785]), .CLK(clk), .RST(rst), .Q(
        start_reg[786]) );
  DFF \start_reg_reg[787]  ( .D(start_in[786]), .CLK(clk), .RST(rst), .Q(
        start_reg[787]) );
  DFF \start_reg_reg[788]  ( .D(start_in[787]), .CLK(clk), .RST(rst), .Q(
        start_reg[788]) );
  DFF \start_reg_reg[789]  ( .D(start_in[788]), .CLK(clk), .RST(rst), .Q(
        start_reg[789]) );
  DFF \start_reg_reg[790]  ( .D(start_in[789]), .CLK(clk), .RST(rst), .Q(
        start_reg[790]) );
  DFF \start_reg_reg[791]  ( .D(start_in[790]), .CLK(clk), .RST(rst), .Q(
        start_reg[791]) );
  DFF \start_reg_reg[792]  ( .D(start_in[791]), .CLK(clk), .RST(rst), .Q(
        start_reg[792]) );
  DFF \start_reg_reg[793]  ( .D(start_in[792]), .CLK(clk), .RST(rst), .Q(
        start_reg[793]) );
  DFF \start_reg_reg[794]  ( .D(start_in[793]), .CLK(clk), .RST(rst), .Q(
        start_reg[794]) );
  DFF \start_reg_reg[795]  ( .D(start_in[794]), .CLK(clk), .RST(rst), .Q(
        start_reg[795]) );
  DFF \start_reg_reg[796]  ( .D(start_in[795]), .CLK(clk), .RST(rst), .Q(
        start_reg[796]) );
  DFF \start_reg_reg[797]  ( .D(start_in[796]), .CLK(clk), .RST(rst), .Q(
        start_reg[797]) );
  DFF \start_reg_reg[798]  ( .D(start_in[797]), .CLK(clk), .RST(rst), .Q(
        start_reg[798]) );
  DFF \start_reg_reg[799]  ( .D(start_in[798]), .CLK(clk), .RST(rst), .Q(
        start_reg[799]) );
  DFF \start_reg_reg[800]  ( .D(start_in[799]), .CLK(clk), .RST(rst), .Q(
        start_reg[800]) );
  DFF \start_reg_reg[801]  ( .D(start_in[800]), .CLK(clk), .RST(rst), .Q(
        start_reg[801]) );
  DFF \start_reg_reg[802]  ( .D(start_in[801]), .CLK(clk), .RST(rst), .Q(
        start_reg[802]) );
  DFF \start_reg_reg[803]  ( .D(start_in[802]), .CLK(clk), .RST(rst), .Q(
        start_reg[803]) );
  DFF \start_reg_reg[804]  ( .D(start_in[803]), .CLK(clk), .RST(rst), .Q(
        start_reg[804]) );
  DFF \start_reg_reg[805]  ( .D(start_in[804]), .CLK(clk), .RST(rst), .Q(
        start_reg[805]) );
  DFF \start_reg_reg[806]  ( .D(start_in[805]), .CLK(clk), .RST(rst), .Q(
        start_reg[806]) );
  DFF \start_reg_reg[807]  ( .D(start_in[806]), .CLK(clk), .RST(rst), .Q(
        start_reg[807]) );
  DFF \start_reg_reg[808]  ( .D(start_in[807]), .CLK(clk), .RST(rst), .Q(
        start_reg[808]) );
  DFF \start_reg_reg[809]  ( .D(start_in[808]), .CLK(clk), .RST(rst), .Q(
        start_reg[809]) );
  DFF \start_reg_reg[810]  ( .D(start_in[809]), .CLK(clk), .RST(rst), .Q(
        start_reg[810]) );
  DFF \start_reg_reg[811]  ( .D(start_in[810]), .CLK(clk), .RST(rst), .Q(
        start_reg[811]) );
  DFF \start_reg_reg[812]  ( .D(start_in[811]), .CLK(clk), .RST(rst), .Q(
        start_reg[812]) );
  DFF \start_reg_reg[813]  ( .D(start_in[812]), .CLK(clk), .RST(rst), .Q(
        start_reg[813]) );
  DFF \start_reg_reg[814]  ( .D(start_in[813]), .CLK(clk), .RST(rst), .Q(
        start_reg[814]) );
  DFF \start_reg_reg[815]  ( .D(start_in[814]), .CLK(clk), .RST(rst), .Q(
        start_reg[815]) );
  DFF \start_reg_reg[816]  ( .D(start_in[815]), .CLK(clk), .RST(rst), .Q(
        start_reg[816]) );
  DFF \start_reg_reg[817]  ( .D(start_in[816]), .CLK(clk), .RST(rst), .Q(
        start_reg[817]) );
  DFF \start_reg_reg[818]  ( .D(start_in[817]), .CLK(clk), .RST(rst), .Q(
        start_reg[818]) );
  DFF \start_reg_reg[819]  ( .D(start_in[818]), .CLK(clk), .RST(rst), .Q(
        start_reg[819]) );
  DFF \start_reg_reg[820]  ( .D(start_in[819]), .CLK(clk), .RST(rst), .Q(
        start_reg[820]) );
  DFF \start_reg_reg[821]  ( .D(start_in[820]), .CLK(clk), .RST(rst), .Q(
        start_reg[821]) );
  DFF \start_reg_reg[822]  ( .D(start_in[821]), .CLK(clk), .RST(rst), .Q(
        start_reg[822]) );
  DFF \start_reg_reg[823]  ( .D(start_in[822]), .CLK(clk), .RST(rst), .Q(
        start_reg[823]) );
  DFF \start_reg_reg[824]  ( .D(start_in[823]), .CLK(clk), .RST(rst), .Q(
        start_reg[824]) );
  DFF \start_reg_reg[825]  ( .D(start_in[824]), .CLK(clk), .RST(rst), .Q(
        start_reg[825]) );
  DFF \start_reg_reg[826]  ( .D(start_in[825]), .CLK(clk), .RST(rst), .Q(
        start_reg[826]) );
  DFF \start_reg_reg[827]  ( .D(start_in[826]), .CLK(clk), .RST(rst), .Q(
        start_reg[827]) );
  DFF \start_reg_reg[828]  ( .D(start_in[827]), .CLK(clk), .RST(rst), .Q(
        start_reg[828]) );
  DFF \start_reg_reg[829]  ( .D(start_in[828]), .CLK(clk), .RST(rst), .Q(
        start_reg[829]) );
  DFF \start_reg_reg[830]  ( .D(start_in[829]), .CLK(clk), .RST(rst), .Q(
        start_reg[830]) );
  DFF \start_reg_reg[831]  ( .D(start_in[830]), .CLK(clk), .RST(rst), .Q(
        start_reg[831]) );
  DFF \start_reg_reg[832]  ( .D(start_in[831]), .CLK(clk), .RST(rst), .Q(
        start_reg[832]) );
  DFF \start_reg_reg[833]  ( .D(start_in[832]), .CLK(clk), .RST(rst), .Q(
        start_reg[833]) );
  DFF \start_reg_reg[834]  ( .D(start_in[833]), .CLK(clk), .RST(rst), .Q(
        start_reg[834]) );
  DFF \start_reg_reg[835]  ( .D(start_in[834]), .CLK(clk), .RST(rst), .Q(
        start_reg[835]) );
  DFF \start_reg_reg[836]  ( .D(start_in[835]), .CLK(clk), .RST(rst), .Q(
        start_reg[836]) );
  DFF \start_reg_reg[837]  ( .D(start_in[836]), .CLK(clk), .RST(rst), .Q(
        start_reg[837]) );
  DFF \start_reg_reg[838]  ( .D(start_in[837]), .CLK(clk), .RST(rst), .Q(
        start_reg[838]) );
  DFF \start_reg_reg[839]  ( .D(start_in[838]), .CLK(clk), .RST(rst), .Q(
        start_reg[839]) );
  DFF \start_reg_reg[840]  ( .D(start_in[839]), .CLK(clk), .RST(rst), .Q(
        start_reg[840]) );
  DFF \start_reg_reg[841]  ( .D(start_in[840]), .CLK(clk), .RST(rst), .Q(
        start_reg[841]) );
  DFF \start_reg_reg[842]  ( .D(start_in[841]), .CLK(clk), .RST(rst), .Q(
        start_reg[842]) );
  DFF \start_reg_reg[843]  ( .D(start_in[842]), .CLK(clk), .RST(rst), .Q(
        start_reg[843]) );
  DFF \start_reg_reg[844]  ( .D(start_in[843]), .CLK(clk), .RST(rst), .Q(
        start_reg[844]) );
  DFF \start_reg_reg[845]  ( .D(start_in[844]), .CLK(clk), .RST(rst), .Q(
        start_reg[845]) );
  DFF \start_reg_reg[846]  ( .D(start_in[845]), .CLK(clk), .RST(rst), .Q(
        start_reg[846]) );
  DFF \start_reg_reg[847]  ( .D(start_in[846]), .CLK(clk), .RST(rst), .Q(
        start_reg[847]) );
  DFF \start_reg_reg[848]  ( .D(start_in[847]), .CLK(clk), .RST(rst), .Q(
        start_reg[848]) );
  DFF \start_reg_reg[849]  ( .D(start_in[848]), .CLK(clk), .RST(rst), .Q(
        start_reg[849]) );
  DFF \start_reg_reg[850]  ( .D(start_in[849]), .CLK(clk), .RST(rst), .Q(
        start_reg[850]) );
  DFF \start_reg_reg[851]  ( .D(start_in[850]), .CLK(clk), .RST(rst), .Q(
        start_reg[851]) );
  DFF \start_reg_reg[852]  ( .D(start_in[851]), .CLK(clk), .RST(rst), .Q(
        start_reg[852]) );
  DFF \start_reg_reg[853]  ( .D(start_in[852]), .CLK(clk), .RST(rst), .Q(
        start_reg[853]) );
  DFF \start_reg_reg[854]  ( .D(start_in[853]), .CLK(clk), .RST(rst), .Q(
        start_reg[854]) );
  DFF \start_reg_reg[855]  ( .D(start_in[854]), .CLK(clk), .RST(rst), .Q(
        start_reg[855]) );
  DFF \start_reg_reg[856]  ( .D(start_in[855]), .CLK(clk), .RST(rst), .Q(
        start_reg[856]) );
  DFF \start_reg_reg[857]  ( .D(start_in[856]), .CLK(clk), .RST(rst), .Q(
        start_reg[857]) );
  DFF \start_reg_reg[858]  ( .D(start_in[857]), .CLK(clk), .RST(rst), .Q(
        start_reg[858]) );
  DFF \start_reg_reg[859]  ( .D(start_in[858]), .CLK(clk), .RST(rst), .Q(
        start_reg[859]) );
  DFF \start_reg_reg[860]  ( .D(start_in[859]), .CLK(clk), .RST(rst), .Q(
        start_reg[860]) );
  DFF \start_reg_reg[861]  ( .D(start_in[860]), .CLK(clk), .RST(rst), .Q(
        start_reg[861]) );
  DFF \start_reg_reg[862]  ( .D(start_in[861]), .CLK(clk), .RST(rst), .Q(
        start_reg[862]) );
  DFF \start_reg_reg[863]  ( .D(start_in[862]), .CLK(clk), .RST(rst), .Q(
        start_reg[863]) );
  DFF \start_reg_reg[864]  ( .D(start_in[863]), .CLK(clk), .RST(rst), .Q(
        start_reg[864]) );
  DFF \start_reg_reg[865]  ( .D(start_in[864]), .CLK(clk), .RST(rst), .Q(
        start_reg[865]) );
  DFF \start_reg_reg[866]  ( .D(start_in[865]), .CLK(clk), .RST(rst), .Q(
        start_reg[866]) );
  DFF \start_reg_reg[867]  ( .D(start_in[866]), .CLK(clk), .RST(rst), .Q(
        start_reg[867]) );
  DFF \start_reg_reg[868]  ( .D(start_in[867]), .CLK(clk), .RST(rst), .Q(
        start_reg[868]) );
  DFF \start_reg_reg[869]  ( .D(start_in[868]), .CLK(clk), .RST(rst), .Q(
        start_reg[869]) );
  DFF \start_reg_reg[870]  ( .D(start_in[869]), .CLK(clk), .RST(rst), .Q(
        start_reg[870]) );
  DFF \start_reg_reg[871]  ( .D(start_in[870]), .CLK(clk), .RST(rst), .Q(
        start_reg[871]) );
  DFF \start_reg_reg[872]  ( .D(start_in[871]), .CLK(clk), .RST(rst), .Q(
        start_reg[872]) );
  DFF \start_reg_reg[873]  ( .D(start_in[872]), .CLK(clk), .RST(rst), .Q(
        start_reg[873]) );
  DFF \start_reg_reg[874]  ( .D(start_in[873]), .CLK(clk), .RST(rst), .Q(
        start_reg[874]) );
  DFF \start_reg_reg[875]  ( .D(start_in[874]), .CLK(clk), .RST(rst), .Q(
        start_reg[875]) );
  DFF \start_reg_reg[876]  ( .D(start_in[875]), .CLK(clk), .RST(rst), .Q(
        start_reg[876]) );
  DFF \start_reg_reg[877]  ( .D(start_in[876]), .CLK(clk), .RST(rst), .Q(
        start_reg[877]) );
  DFF \start_reg_reg[878]  ( .D(start_in[877]), .CLK(clk), .RST(rst), .Q(
        start_reg[878]) );
  DFF \start_reg_reg[879]  ( .D(start_in[878]), .CLK(clk), .RST(rst), .Q(
        start_reg[879]) );
  DFF \start_reg_reg[880]  ( .D(start_in[879]), .CLK(clk), .RST(rst), .Q(
        start_reg[880]) );
  DFF \start_reg_reg[881]  ( .D(start_in[880]), .CLK(clk), .RST(rst), .Q(
        start_reg[881]) );
  DFF \start_reg_reg[882]  ( .D(start_in[881]), .CLK(clk), .RST(rst), .Q(
        start_reg[882]) );
  DFF \start_reg_reg[883]  ( .D(start_in[882]), .CLK(clk), .RST(rst), .Q(
        start_reg[883]) );
  DFF \start_reg_reg[884]  ( .D(start_in[883]), .CLK(clk), .RST(rst), .Q(
        start_reg[884]) );
  DFF \start_reg_reg[885]  ( .D(start_in[884]), .CLK(clk), .RST(rst), .Q(
        start_reg[885]) );
  DFF \start_reg_reg[886]  ( .D(start_in[885]), .CLK(clk), .RST(rst), .Q(
        start_reg[886]) );
  DFF \start_reg_reg[887]  ( .D(start_in[886]), .CLK(clk), .RST(rst), .Q(
        start_reg[887]) );
  DFF \start_reg_reg[888]  ( .D(start_in[887]), .CLK(clk), .RST(rst), .Q(
        start_reg[888]) );
  DFF \start_reg_reg[889]  ( .D(start_in[888]), .CLK(clk), .RST(rst), .Q(
        start_reg[889]) );
  DFF \start_reg_reg[890]  ( .D(start_in[889]), .CLK(clk), .RST(rst), .Q(
        start_reg[890]) );
  DFF \start_reg_reg[891]  ( .D(start_in[890]), .CLK(clk), .RST(rst), .Q(
        start_reg[891]) );
  DFF \start_reg_reg[892]  ( .D(start_in[891]), .CLK(clk), .RST(rst), .Q(
        start_reg[892]) );
  DFF \start_reg_reg[893]  ( .D(start_in[892]), .CLK(clk), .RST(rst), .Q(
        start_reg[893]) );
  DFF \start_reg_reg[894]  ( .D(start_in[893]), .CLK(clk), .RST(rst), .Q(
        start_reg[894]) );
  DFF \start_reg_reg[895]  ( .D(start_in[894]), .CLK(clk), .RST(rst), .Q(
        start_reg[895]) );
  DFF \start_reg_reg[896]  ( .D(start_in[895]), .CLK(clk), .RST(rst), .Q(
        start_reg[896]) );
  DFF \start_reg_reg[897]  ( .D(start_in[896]), .CLK(clk), .RST(rst), .Q(
        start_reg[897]) );
  DFF \start_reg_reg[898]  ( .D(start_in[897]), .CLK(clk), .RST(rst), .Q(
        start_reg[898]) );
  DFF \start_reg_reg[899]  ( .D(start_in[898]), .CLK(clk), .RST(rst), .Q(
        start_reg[899]) );
  DFF \start_reg_reg[900]  ( .D(start_in[899]), .CLK(clk), .RST(rst), .Q(
        start_reg[900]) );
  DFF \start_reg_reg[901]  ( .D(start_in[900]), .CLK(clk), .RST(rst), .Q(
        start_reg[901]) );
  DFF \start_reg_reg[902]  ( .D(start_in[901]), .CLK(clk), .RST(rst), .Q(
        start_reg[902]) );
  DFF \start_reg_reg[903]  ( .D(start_in[902]), .CLK(clk), .RST(rst), .Q(
        start_reg[903]) );
  DFF \start_reg_reg[904]  ( .D(start_in[903]), .CLK(clk), .RST(rst), .Q(
        start_reg[904]) );
  DFF \start_reg_reg[905]  ( .D(start_in[904]), .CLK(clk), .RST(rst), .Q(
        start_reg[905]) );
  DFF \start_reg_reg[906]  ( .D(start_in[905]), .CLK(clk), .RST(rst), .Q(
        start_reg[906]) );
  DFF \start_reg_reg[907]  ( .D(start_in[906]), .CLK(clk), .RST(rst), .Q(
        start_reg[907]) );
  DFF \start_reg_reg[908]  ( .D(start_in[907]), .CLK(clk), .RST(rst), .Q(
        start_reg[908]) );
  DFF \start_reg_reg[909]  ( .D(start_in[908]), .CLK(clk), .RST(rst), .Q(
        start_reg[909]) );
  DFF \start_reg_reg[910]  ( .D(start_in[909]), .CLK(clk), .RST(rst), .Q(
        start_reg[910]) );
  DFF \start_reg_reg[911]  ( .D(start_in[910]), .CLK(clk), .RST(rst), .Q(
        start_reg[911]) );
  DFF \start_reg_reg[912]  ( .D(start_in[911]), .CLK(clk), .RST(rst), .Q(
        start_reg[912]) );
  DFF \start_reg_reg[913]  ( .D(start_in[912]), .CLK(clk), .RST(rst), .Q(
        start_reg[913]) );
  DFF \start_reg_reg[914]  ( .D(start_in[913]), .CLK(clk), .RST(rst), .Q(
        start_reg[914]) );
  DFF \start_reg_reg[915]  ( .D(start_in[914]), .CLK(clk), .RST(rst), .Q(
        start_reg[915]) );
  DFF \start_reg_reg[916]  ( .D(start_in[915]), .CLK(clk), .RST(rst), .Q(
        start_reg[916]) );
  DFF \start_reg_reg[917]  ( .D(start_in[916]), .CLK(clk), .RST(rst), .Q(
        start_reg[917]) );
  DFF \start_reg_reg[918]  ( .D(start_in[917]), .CLK(clk), .RST(rst), .Q(
        start_reg[918]) );
  DFF \start_reg_reg[919]  ( .D(start_in[918]), .CLK(clk), .RST(rst), .Q(
        start_reg[919]) );
  DFF \start_reg_reg[920]  ( .D(start_in[919]), .CLK(clk), .RST(rst), .Q(
        start_reg[920]) );
  DFF \start_reg_reg[921]  ( .D(start_in[920]), .CLK(clk), .RST(rst), .Q(
        start_reg[921]) );
  DFF \start_reg_reg[922]  ( .D(start_in[921]), .CLK(clk), .RST(rst), .Q(
        start_reg[922]) );
  DFF \start_reg_reg[923]  ( .D(start_in[922]), .CLK(clk), .RST(rst), .Q(
        start_reg[923]) );
  DFF \start_reg_reg[924]  ( .D(start_in[923]), .CLK(clk), .RST(rst), .Q(
        start_reg[924]) );
  DFF \start_reg_reg[925]  ( .D(start_in[924]), .CLK(clk), .RST(rst), .Q(
        start_reg[925]) );
  DFF \start_reg_reg[926]  ( .D(start_in[925]), .CLK(clk), .RST(rst), .Q(
        start_reg[926]) );
  DFF \start_reg_reg[927]  ( .D(start_in[926]), .CLK(clk), .RST(rst), .Q(
        start_reg[927]) );
  DFF \start_reg_reg[928]  ( .D(start_in[927]), .CLK(clk), .RST(rst), .Q(
        start_reg[928]) );
  DFF \start_reg_reg[929]  ( .D(start_in[928]), .CLK(clk), .RST(rst), .Q(
        start_reg[929]) );
  DFF \start_reg_reg[930]  ( .D(start_in[929]), .CLK(clk), .RST(rst), .Q(
        start_reg[930]) );
  DFF \start_reg_reg[931]  ( .D(start_in[930]), .CLK(clk), .RST(rst), .Q(
        start_reg[931]) );
  DFF \start_reg_reg[932]  ( .D(start_in[931]), .CLK(clk), .RST(rst), .Q(
        start_reg[932]) );
  DFF \start_reg_reg[933]  ( .D(start_in[932]), .CLK(clk), .RST(rst), .Q(
        start_reg[933]) );
  DFF \start_reg_reg[934]  ( .D(start_in[933]), .CLK(clk), .RST(rst), .Q(
        start_reg[934]) );
  DFF \start_reg_reg[935]  ( .D(start_in[934]), .CLK(clk), .RST(rst), .Q(
        start_reg[935]) );
  DFF \start_reg_reg[936]  ( .D(start_in[935]), .CLK(clk), .RST(rst), .Q(
        start_reg[936]) );
  DFF \start_reg_reg[937]  ( .D(start_in[936]), .CLK(clk), .RST(rst), .Q(
        start_reg[937]) );
  DFF \start_reg_reg[938]  ( .D(start_in[937]), .CLK(clk), .RST(rst), .Q(
        start_reg[938]) );
  DFF \start_reg_reg[939]  ( .D(start_in[938]), .CLK(clk), .RST(rst), .Q(
        start_reg[939]) );
  DFF \start_reg_reg[940]  ( .D(start_in[939]), .CLK(clk), .RST(rst), .Q(
        start_reg[940]) );
  DFF \start_reg_reg[941]  ( .D(start_in[940]), .CLK(clk), .RST(rst), .Q(
        start_reg[941]) );
  DFF \start_reg_reg[942]  ( .D(start_in[941]), .CLK(clk), .RST(rst), .Q(
        start_reg[942]) );
  DFF \start_reg_reg[943]  ( .D(start_in[942]), .CLK(clk), .RST(rst), .Q(
        start_reg[943]) );
  DFF \start_reg_reg[944]  ( .D(start_in[943]), .CLK(clk), .RST(rst), .Q(
        start_reg[944]) );
  DFF \start_reg_reg[945]  ( .D(start_in[944]), .CLK(clk), .RST(rst), .Q(
        start_reg[945]) );
  DFF \start_reg_reg[946]  ( .D(start_in[945]), .CLK(clk), .RST(rst), .Q(
        start_reg[946]) );
  DFF \start_reg_reg[947]  ( .D(start_in[946]), .CLK(clk), .RST(rst), .Q(
        start_reg[947]) );
  DFF \start_reg_reg[948]  ( .D(start_in[947]), .CLK(clk), .RST(rst), .Q(
        start_reg[948]) );
  DFF \start_reg_reg[949]  ( .D(start_in[948]), .CLK(clk), .RST(rst), .Q(
        start_reg[949]) );
  DFF \start_reg_reg[950]  ( .D(start_in[949]), .CLK(clk), .RST(rst), .Q(
        start_reg[950]) );
  DFF \start_reg_reg[951]  ( .D(start_in[950]), .CLK(clk), .RST(rst), .Q(
        start_reg[951]) );
  DFF \start_reg_reg[952]  ( .D(start_in[951]), .CLK(clk), .RST(rst), .Q(
        start_reg[952]) );
  DFF \start_reg_reg[953]  ( .D(start_in[952]), .CLK(clk), .RST(rst), .Q(
        start_reg[953]) );
  DFF \start_reg_reg[954]  ( .D(start_in[953]), .CLK(clk), .RST(rst), .Q(
        start_reg[954]) );
  DFF \start_reg_reg[955]  ( .D(start_in[954]), .CLK(clk), .RST(rst), .Q(
        start_reg[955]) );
  DFF \start_reg_reg[956]  ( .D(start_in[955]), .CLK(clk), .RST(rst), .Q(
        start_reg[956]) );
  DFF \start_reg_reg[957]  ( .D(start_in[956]), .CLK(clk), .RST(rst), .Q(
        start_reg[957]) );
  DFF \start_reg_reg[958]  ( .D(start_in[957]), .CLK(clk), .RST(rst), .Q(
        start_reg[958]) );
  DFF \start_reg_reg[959]  ( .D(start_in[958]), .CLK(clk), .RST(rst), .Q(
        start_reg[959]) );
  DFF \start_reg_reg[960]  ( .D(start_in[959]), .CLK(clk), .RST(rst), .Q(
        start_reg[960]) );
  DFF \start_reg_reg[961]  ( .D(start_in[960]), .CLK(clk), .RST(rst), .Q(
        start_reg[961]) );
  DFF \start_reg_reg[962]  ( .D(start_in[961]), .CLK(clk), .RST(rst), .Q(
        start_reg[962]) );
  DFF \start_reg_reg[963]  ( .D(start_in[962]), .CLK(clk), .RST(rst), .Q(
        start_reg[963]) );
  DFF \start_reg_reg[964]  ( .D(start_in[963]), .CLK(clk), .RST(rst), .Q(
        start_reg[964]) );
  DFF \start_reg_reg[965]  ( .D(start_in[964]), .CLK(clk), .RST(rst), .Q(
        start_reg[965]) );
  DFF \start_reg_reg[966]  ( .D(start_in[965]), .CLK(clk), .RST(rst), .Q(
        start_reg[966]) );
  DFF \start_reg_reg[967]  ( .D(start_in[966]), .CLK(clk), .RST(rst), .Q(
        start_reg[967]) );
  DFF \start_reg_reg[968]  ( .D(start_in[967]), .CLK(clk), .RST(rst), .Q(
        start_reg[968]) );
  DFF \start_reg_reg[969]  ( .D(start_in[968]), .CLK(clk), .RST(rst), .Q(
        start_reg[969]) );
  DFF \start_reg_reg[970]  ( .D(start_in[969]), .CLK(clk), .RST(rst), .Q(
        start_reg[970]) );
  DFF \start_reg_reg[971]  ( .D(start_in[970]), .CLK(clk), .RST(rst), .Q(
        start_reg[971]) );
  DFF \start_reg_reg[972]  ( .D(start_in[971]), .CLK(clk), .RST(rst), .Q(
        start_reg[972]) );
  DFF \start_reg_reg[973]  ( .D(start_in[972]), .CLK(clk), .RST(rst), .Q(
        start_reg[973]) );
  DFF \start_reg_reg[974]  ( .D(start_in[973]), .CLK(clk), .RST(rst), .Q(
        start_reg[974]) );
  DFF \start_reg_reg[975]  ( .D(start_in[974]), .CLK(clk), .RST(rst), .Q(
        start_reg[975]) );
  DFF \start_reg_reg[976]  ( .D(start_in[975]), .CLK(clk), .RST(rst), .Q(
        start_reg[976]) );
  DFF \start_reg_reg[977]  ( .D(start_in[976]), .CLK(clk), .RST(rst), .Q(
        start_reg[977]) );
  DFF \start_reg_reg[978]  ( .D(start_in[977]), .CLK(clk), .RST(rst), .Q(
        start_reg[978]) );
  DFF \start_reg_reg[979]  ( .D(start_in[978]), .CLK(clk), .RST(rst), .Q(
        start_reg[979]) );
  DFF \start_reg_reg[980]  ( .D(start_in[979]), .CLK(clk), .RST(rst), .Q(
        start_reg[980]) );
  DFF \start_reg_reg[981]  ( .D(start_in[980]), .CLK(clk), .RST(rst), .Q(
        start_reg[981]) );
  DFF \start_reg_reg[982]  ( .D(start_in[981]), .CLK(clk), .RST(rst), .Q(
        start_reg[982]) );
  DFF \start_reg_reg[983]  ( .D(start_in[982]), .CLK(clk), .RST(rst), .Q(
        start_reg[983]) );
  DFF \start_reg_reg[984]  ( .D(start_in[983]), .CLK(clk), .RST(rst), .Q(
        start_reg[984]) );
  DFF \start_reg_reg[985]  ( .D(start_in[984]), .CLK(clk), .RST(rst), .Q(
        start_reg[985]) );
  DFF \start_reg_reg[986]  ( .D(start_in[985]), .CLK(clk), .RST(rst), .Q(
        start_reg[986]) );
  DFF \start_reg_reg[987]  ( .D(start_in[986]), .CLK(clk), .RST(rst), .Q(
        start_reg[987]) );
  DFF \start_reg_reg[988]  ( .D(start_in[987]), .CLK(clk), .RST(rst), .Q(
        start_reg[988]) );
  DFF \start_reg_reg[989]  ( .D(start_in[988]), .CLK(clk), .RST(rst), .Q(
        start_reg[989]) );
  DFF \start_reg_reg[990]  ( .D(start_in[989]), .CLK(clk), .RST(rst), .Q(
        start_reg[990]) );
  DFF \start_reg_reg[991]  ( .D(start_in[990]), .CLK(clk), .RST(rst), .Q(
        start_reg[991]) );
  DFF \start_reg_reg[992]  ( .D(start_in[991]), .CLK(clk), .RST(rst), .Q(
        start_reg[992]) );
  DFF \start_reg_reg[993]  ( .D(start_in[992]), .CLK(clk), .RST(rst), .Q(
        start_reg[993]) );
  DFF \start_reg_reg[994]  ( .D(start_in[993]), .CLK(clk), .RST(rst), .Q(
        start_reg[994]) );
  DFF \start_reg_reg[995]  ( .D(start_in[994]), .CLK(clk), .RST(rst), .Q(
        start_reg[995]) );
  DFF \start_reg_reg[996]  ( .D(start_in[995]), .CLK(clk), .RST(rst), .Q(
        start_reg[996]) );
  DFF \start_reg_reg[997]  ( .D(start_in[996]), .CLK(clk), .RST(rst), .Q(
        start_reg[997]) );
  DFF \start_reg_reg[998]  ( .D(start_in[997]), .CLK(clk), .RST(rst), .Q(
        start_reg[998]) );
  DFF \start_reg_reg[999]  ( .D(start_in[998]), .CLK(clk), .RST(rst), .Q(
        start_reg[999]) );
  DFF \start_reg_reg[1000]  ( .D(start_in[999]), .CLK(clk), .RST(rst), .Q(
        start_reg[1000]) );
  DFF \start_reg_reg[1001]  ( .D(start_in[1000]), .CLK(clk), .RST(rst), .Q(
        start_reg[1001]) );
  DFF \start_reg_reg[1002]  ( .D(start_in[1001]), .CLK(clk), .RST(rst), .Q(
        start_reg[1002]) );
  DFF \start_reg_reg[1003]  ( .D(start_in[1002]), .CLK(clk), .RST(rst), .Q(
        start_reg[1003]) );
  DFF \start_reg_reg[1004]  ( .D(start_in[1003]), .CLK(clk), .RST(rst), .Q(
        start_reg[1004]) );
  DFF \start_reg_reg[1005]  ( .D(start_in[1004]), .CLK(clk), .RST(rst), .Q(
        start_reg[1005]) );
  DFF \start_reg_reg[1006]  ( .D(start_in[1005]), .CLK(clk), .RST(rst), .Q(
        start_reg[1006]) );
  DFF \start_reg_reg[1007]  ( .D(start_in[1006]), .CLK(clk), .RST(rst), .Q(
        start_reg[1007]) );
  DFF \start_reg_reg[1008]  ( .D(start_in[1007]), .CLK(clk), .RST(rst), .Q(
        start_reg[1008]) );
  DFF \start_reg_reg[1009]  ( .D(start_in[1008]), .CLK(clk), .RST(rst), .Q(
        start_reg[1009]) );
  DFF \start_reg_reg[1010]  ( .D(start_in[1009]), .CLK(clk), .RST(rst), .Q(
        start_reg[1010]) );
  DFF \start_reg_reg[1011]  ( .D(start_in[1010]), .CLK(clk), .RST(rst), .Q(
        start_reg[1011]) );
  DFF \start_reg_reg[1012]  ( .D(start_in[1011]), .CLK(clk), .RST(rst), .Q(
        start_reg[1012]) );
  DFF \start_reg_reg[1013]  ( .D(start_in[1012]), .CLK(clk), .RST(rst), .Q(
        start_reg[1013]) );
  DFF \start_reg_reg[1014]  ( .D(start_in[1013]), .CLK(clk), .RST(rst), .Q(
        start_reg[1014]) );
  DFF \start_reg_reg[1015]  ( .D(start_in[1014]), .CLK(clk), .RST(rst), .Q(
        start_reg[1015]) );
  DFF \start_reg_reg[1016]  ( .D(start_in[1015]), .CLK(clk), .RST(rst), .Q(
        start_reg[1016]) );
  DFF \start_reg_reg[1017]  ( .D(start_in[1016]), .CLK(clk), .RST(rst), .Q(
        start_reg[1017]) );
  DFF \start_reg_reg[1018]  ( .D(start_in[1017]), .CLK(clk), .RST(rst), .Q(
        start_reg[1018]) );
  DFF \start_reg_reg[1019]  ( .D(start_in[1018]), .CLK(clk), .RST(rst), .Q(
        start_reg[1019]) );
  DFF \start_reg_reg[1020]  ( .D(start_in[1019]), .CLK(clk), .RST(rst), .Q(
        start_reg[1020]) );
  DFF \start_reg_reg[1021]  ( .D(start_in[1020]), .CLK(clk), .RST(rst), .Q(
        start_reg[1021]) );
  DFF \start_reg_reg[1022]  ( .D(start_in[1021]), .CLK(clk), .RST(rst), .Q(
        start_reg[1022]) );
  DFF \start_reg_reg[1023]  ( .D(start_in[1022]), .CLK(clk), .RST(rst), .Q(
        start_reg[1023]) );
  DFF mul_pow_reg ( .D(n3860), .CLK(clk), .RST(rst), .Q(mul_pow) );
  DFF \ereg_reg[0]  ( .D(n3859), .CLK(clk), .RST(rst), .Q(ereg[0]) );
  DFF \ereg_reg[1]  ( .D(n3858), .CLK(clk), .RST(rst), .Q(ereg[1]) );
  DFF \ereg_reg[2]  ( .D(n3857), .CLK(clk), .RST(rst), .Q(ereg[2]) );
  DFF \ereg_reg[3]  ( .D(n3856), .CLK(clk), .RST(rst), .Q(ereg[3]) );
  DFF \ereg_reg[4]  ( .D(n3855), .CLK(clk), .RST(rst), .Q(ereg[4]) );
  DFF \ereg_reg[5]  ( .D(n3854), .CLK(clk), .RST(rst), .Q(ereg[5]) );
  DFF \ereg_reg[6]  ( .D(n3853), .CLK(clk), .RST(rst), .Q(ereg[6]) );
  DFF \ereg_reg[7]  ( .D(n3852), .CLK(clk), .RST(rst), .Q(ereg[7]) );
  DFF \ereg_reg[8]  ( .D(n3851), .CLK(clk), .RST(rst), .Q(ereg[8]) );
  DFF \ereg_reg[9]  ( .D(n3850), .CLK(clk), .RST(rst), .Q(ereg[9]) );
  DFF \ereg_reg[10]  ( .D(n3849), .CLK(clk), .RST(rst), .Q(ereg[10]) );
  DFF \ereg_reg[11]  ( .D(n3848), .CLK(clk), .RST(rst), .Q(ereg[11]) );
  DFF \ereg_reg[12]  ( .D(n3847), .CLK(clk), .RST(rst), .Q(ereg[12]) );
  DFF \ereg_reg[13]  ( .D(n3846), .CLK(clk), .RST(rst), .Q(ereg[13]) );
  DFF \ereg_reg[14]  ( .D(n3845), .CLK(clk), .RST(rst), .Q(ereg[14]) );
  DFF \ereg_reg[15]  ( .D(n3844), .CLK(clk), .RST(rst), .Q(ereg[15]) );
  DFF \ereg_reg[16]  ( .D(n3843), .CLK(clk), .RST(rst), .Q(ereg[16]) );
  DFF \ereg_reg[17]  ( .D(n3842), .CLK(clk), .RST(rst), .Q(ereg[17]) );
  DFF \ereg_reg[18]  ( .D(n3841), .CLK(clk), .RST(rst), .Q(ereg[18]) );
  DFF \ereg_reg[19]  ( .D(n3840), .CLK(clk), .RST(rst), .Q(ereg[19]) );
  DFF \ereg_reg[20]  ( .D(n3839), .CLK(clk), .RST(rst), .Q(ereg[20]) );
  DFF \ereg_reg[21]  ( .D(n3838), .CLK(clk), .RST(rst), .Q(ereg[21]) );
  DFF \ereg_reg[22]  ( .D(n3837), .CLK(clk), .RST(rst), .Q(ereg[22]) );
  DFF \ereg_reg[23]  ( .D(n3836), .CLK(clk), .RST(rst), .Q(ereg[23]) );
  DFF \ereg_reg[24]  ( .D(n3835), .CLK(clk), .RST(rst), .Q(ereg[24]) );
  DFF \ereg_reg[25]  ( .D(n3834), .CLK(clk), .RST(rst), .Q(ereg[25]) );
  DFF \ereg_reg[26]  ( .D(n3833), .CLK(clk), .RST(rst), .Q(ereg[26]) );
  DFF \ereg_reg[27]  ( .D(n3832), .CLK(clk), .RST(rst), .Q(ereg[27]) );
  DFF \ereg_reg[28]  ( .D(n3831), .CLK(clk), .RST(rst), .Q(ereg[28]) );
  DFF \ereg_reg[29]  ( .D(n3830), .CLK(clk), .RST(rst), .Q(ereg[29]) );
  DFF \ereg_reg[30]  ( .D(n3829), .CLK(clk), .RST(rst), .Q(ereg[30]) );
  DFF \ereg_reg[31]  ( .D(n3828), .CLK(clk), .RST(rst), .Q(ereg[31]) );
  DFF \ereg_reg[32]  ( .D(n3827), .CLK(clk), .RST(rst), .Q(ereg[32]) );
  DFF \ereg_reg[33]  ( .D(n3826), .CLK(clk), .RST(rst), .Q(ereg[33]) );
  DFF \ereg_reg[34]  ( .D(n3825), .CLK(clk), .RST(rst), .Q(ereg[34]) );
  DFF \ereg_reg[35]  ( .D(n3824), .CLK(clk), .RST(rst), .Q(ereg[35]) );
  DFF \ereg_reg[36]  ( .D(n3823), .CLK(clk), .RST(rst), .Q(ereg[36]) );
  DFF \ereg_reg[37]  ( .D(n3822), .CLK(clk), .RST(rst), .Q(ereg[37]) );
  DFF \ereg_reg[38]  ( .D(n3821), .CLK(clk), .RST(rst), .Q(ereg[38]) );
  DFF \ereg_reg[39]  ( .D(n3820), .CLK(clk), .RST(rst), .Q(ereg[39]) );
  DFF \ereg_reg[40]  ( .D(n3819), .CLK(clk), .RST(rst), .Q(ereg[40]) );
  DFF \ereg_reg[41]  ( .D(n3818), .CLK(clk), .RST(rst), .Q(ereg[41]) );
  DFF \ereg_reg[42]  ( .D(n3817), .CLK(clk), .RST(rst), .Q(ereg[42]) );
  DFF \ereg_reg[43]  ( .D(n3816), .CLK(clk), .RST(rst), .Q(ereg[43]) );
  DFF \ereg_reg[44]  ( .D(n3815), .CLK(clk), .RST(rst), .Q(ereg[44]) );
  DFF \ereg_reg[45]  ( .D(n3814), .CLK(clk), .RST(rst), .Q(ereg[45]) );
  DFF \ereg_reg[46]  ( .D(n3813), .CLK(clk), .RST(rst), .Q(ereg[46]) );
  DFF \ereg_reg[47]  ( .D(n3812), .CLK(clk), .RST(rst), .Q(ereg[47]) );
  DFF \ereg_reg[48]  ( .D(n3811), .CLK(clk), .RST(rst), .Q(ereg[48]) );
  DFF \ereg_reg[49]  ( .D(n3810), .CLK(clk), .RST(rst), .Q(ereg[49]) );
  DFF \ereg_reg[50]  ( .D(n3809), .CLK(clk), .RST(rst), .Q(ereg[50]) );
  DFF \ereg_reg[51]  ( .D(n3808), .CLK(clk), .RST(rst), .Q(ereg[51]) );
  DFF \ereg_reg[52]  ( .D(n3807), .CLK(clk), .RST(rst), .Q(ereg[52]) );
  DFF \ereg_reg[53]  ( .D(n3806), .CLK(clk), .RST(rst), .Q(ereg[53]) );
  DFF \ereg_reg[54]  ( .D(n3805), .CLK(clk), .RST(rst), .Q(ereg[54]) );
  DFF \ereg_reg[55]  ( .D(n3804), .CLK(clk), .RST(rst), .Q(ereg[55]) );
  DFF \ereg_reg[56]  ( .D(n3803), .CLK(clk), .RST(rst), .Q(ereg[56]) );
  DFF \ereg_reg[57]  ( .D(n3802), .CLK(clk), .RST(rst), .Q(ereg[57]) );
  DFF \ereg_reg[58]  ( .D(n3801), .CLK(clk), .RST(rst), .Q(ereg[58]) );
  DFF \ereg_reg[59]  ( .D(n3800), .CLK(clk), .RST(rst), .Q(ereg[59]) );
  DFF \ereg_reg[60]  ( .D(n3799), .CLK(clk), .RST(rst), .Q(ereg[60]) );
  DFF \ereg_reg[61]  ( .D(n3798), .CLK(clk), .RST(rst), .Q(ereg[61]) );
  DFF \ereg_reg[62]  ( .D(n3797), .CLK(clk), .RST(rst), .Q(ereg[62]) );
  DFF \ereg_reg[63]  ( .D(n3796), .CLK(clk), .RST(rst), .Q(ereg[63]) );
  DFF \ereg_reg[64]  ( .D(n3795), .CLK(clk), .RST(rst), .Q(ereg[64]) );
  DFF \ereg_reg[65]  ( .D(n3794), .CLK(clk), .RST(rst), .Q(ereg[65]) );
  DFF \ereg_reg[66]  ( .D(n3793), .CLK(clk), .RST(rst), .Q(ereg[66]) );
  DFF \ereg_reg[67]  ( .D(n3792), .CLK(clk), .RST(rst), .Q(ereg[67]) );
  DFF \ereg_reg[68]  ( .D(n3791), .CLK(clk), .RST(rst), .Q(ereg[68]) );
  DFF \ereg_reg[69]  ( .D(n3790), .CLK(clk), .RST(rst), .Q(ereg[69]) );
  DFF \ereg_reg[70]  ( .D(n3789), .CLK(clk), .RST(rst), .Q(ereg[70]) );
  DFF \ereg_reg[71]  ( .D(n3788), .CLK(clk), .RST(rst), .Q(ereg[71]) );
  DFF \ereg_reg[72]  ( .D(n3787), .CLK(clk), .RST(rst), .Q(ereg[72]) );
  DFF \ereg_reg[73]  ( .D(n3786), .CLK(clk), .RST(rst), .Q(ereg[73]) );
  DFF \ereg_reg[74]  ( .D(n3785), .CLK(clk), .RST(rst), .Q(ereg[74]) );
  DFF \ereg_reg[75]  ( .D(n3784), .CLK(clk), .RST(rst), .Q(ereg[75]) );
  DFF \ereg_reg[76]  ( .D(n3783), .CLK(clk), .RST(rst), .Q(ereg[76]) );
  DFF \ereg_reg[77]  ( .D(n3782), .CLK(clk), .RST(rst), .Q(ereg[77]) );
  DFF \ereg_reg[78]  ( .D(n3781), .CLK(clk), .RST(rst), .Q(ereg[78]) );
  DFF \ereg_reg[79]  ( .D(n3780), .CLK(clk), .RST(rst), .Q(ereg[79]) );
  DFF \ereg_reg[80]  ( .D(n3779), .CLK(clk), .RST(rst), .Q(ereg[80]) );
  DFF \ereg_reg[81]  ( .D(n3778), .CLK(clk), .RST(rst), .Q(ereg[81]) );
  DFF \ereg_reg[82]  ( .D(n3777), .CLK(clk), .RST(rst), .Q(ereg[82]) );
  DFF \ereg_reg[83]  ( .D(n3776), .CLK(clk), .RST(rst), .Q(ereg[83]) );
  DFF \ereg_reg[84]  ( .D(n3775), .CLK(clk), .RST(rst), .Q(ereg[84]) );
  DFF \ereg_reg[85]  ( .D(n3774), .CLK(clk), .RST(rst), .Q(ereg[85]) );
  DFF \ereg_reg[86]  ( .D(n3773), .CLK(clk), .RST(rst), .Q(ereg[86]) );
  DFF \ereg_reg[87]  ( .D(n3772), .CLK(clk), .RST(rst), .Q(ereg[87]) );
  DFF \ereg_reg[88]  ( .D(n3771), .CLK(clk), .RST(rst), .Q(ereg[88]) );
  DFF \ereg_reg[89]  ( .D(n3770), .CLK(clk), .RST(rst), .Q(ereg[89]) );
  DFF \ereg_reg[90]  ( .D(n3769), .CLK(clk), .RST(rst), .Q(ereg[90]) );
  DFF \ereg_reg[91]  ( .D(n3768), .CLK(clk), .RST(rst), .Q(ereg[91]) );
  DFF \ereg_reg[92]  ( .D(n3767), .CLK(clk), .RST(rst), .Q(ereg[92]) );
  DFF \ereg_reg[93]  ( .D(n3766), .CLK(clk), .RST(rst), .Q(ereg[93]) );
  DFF \ereg_reg[94]  ( .D(n3765), .CLK(clk), .RST(rst), .Q(ereg[94]) );
  DFF \ereg_reg[95]  ( .D(n3764), .CLK(clk), .RST(rst), .Q(ereg[95]) );
  DFF \ereg_reg[96]  ( .D(n3763), .CLK(clk), .RST(rst), .Q(ereg[96]) );
  DFF \ereg_reg[97]  ( .D(n3762), .CLK(clk), .RST(rst), .Q(ereg[97]) );
  DFF \ereg_reg[98]  ( .D(n3761), .CLK(clk), .RST(rst), .Q(ereg[98]) );
  DFF \ereg_reg[99]  ( .D(n3760), .CLK(clk), .RST(rst), .Q(ereg[99]) );
  DFF \ereg_reg[100]  ( .D(n3759), .CLK(clk), .RST(rst), .Q(ereg[100]) );
  DFF \ereg_reg[101]  ( .D(n3758), .CLK(clk), .RST(rst), .Q(ereg[101]) );
  DFF \ereg_reg[102]  ( .D(n3757), .CLK(clk), .RST(rst), .Q(ereg[102]) );
  DFF \ereg_reg[103]  ( .D(n3756), .CLK(clk), .RST(rst), .Q(ereg[103]) );
  DFF \ereg_reg[104]  ( .D(n3755), .CLK(clk), .RST(rst), .Q(ereg[104]) );
  DFF \ereg_reg[105]  ( .D(n3754), .CLK(clk), .RST(rst), .Q(ereg[105]) );
  DFF \ereg_reg[106]  ( .D(n3753), .CLK(clk), .RST(rst), .Q(ereg[106]) );
  DFF \ereg_reg[107]  ( .D(n3752), .CLK(clk), .RST(rst), .Q(ereg[107]) );
  DFF \ereg_reg[108]  ( .D(n3751), .CLK(clk), .RST(rst), .Q(ereg[108]) );
  DFF \ereg_reg[109]  ( .D(n3750), .CLK(clk), .RST(rst), .Q(ereg[109]) );
  DFF \ereg_reg[110]  ( .D(n3749), .CLK(clk), .RST(rst), .Q(ereg[110]) );
  DFF \ereg_reg[111]  ( .D(n3748), .CLK(clk), .RST(rst), .Q(ereg[111]) );
  DFF \ereg_reg[112]  ( .D(n3747), .CLK(clk), .RST(rst), .Q(ereg[112]) );
  DFF \ereg_reg[113]  ( .D(n3746), .CLK(clk), .RST(rst), .Q(ereg[113]) );
  DFF \ereg_reg[114]  ( .D(n3745), .CLK(clk), .RST(rst), .Q(ereg[114]) );
  DFF \ereg_reg[115]  ( .D(n3744), .CLK(clk), .RST(rst), .Q(ereg[115]) );
  DFF \ereg_reg[116]  ( .D(n3743), .CLK(clk), .RST(rst), .Q(ereg[116]) );
  DFF \ereg_reg[117]  ( .D(n3742), .CLK(clk), .RST(rst), .Q(ereg[117]) );
  DFF \ereg_reg[118]  ( .D(n3741), .CLK(clk), .RST(rst), .Q(ereg[118]) );
  DFF \ereg_reg[119]  ( .D(n3740), .CLK(clk), .RST(rst), .Q(ereg[119]) );
  DFF \ereg_reg[120]  ( .D(n3739), .CLK(clk), .RST(rst), .Q(ereg[120]) );
  DFF \ereg_reg[121]  ( .D(n3738), .CLK(clk), .RST(rst), .Q(ereg[121]) );
  DFF \ereg_reg[122]  ( .D(n3737), .CLK(clk), .RST(rst), .Q(ereg[122]) );
  DFF \ereg_reg[123]  ( .D(n3736), .CLK(clk), .RST(rst), .Q(ereg[123]) );
  DFF \ereg_reg[124]  ( .D(n3735), .CLK(clk), .RST(rst), .Q(ereg[124]) );
  DFF \ereg_reg[125]  ( .D(n3734), .CLK(clk), .RST(rst), .Q(ereg[125]) );
  DFF \ereg_reg[126]  ( .D(n3733), .CLK(clk), .RST(rst), .Q(ereg[126]) );
  DFF \ereg_reg[127]  ( .D(n3732), .CLK(clk), .RST(rst), .Q(ereg[127]) );
  DFF \ereg_reg[128]  ( .D(n3731), .CLK(clk), .RST(rst), .Q(ereg[128]) );
  DFF \ereg_reg[129]  ( .D(n3730), .CLK(clk), .RST(rst), .Q(ereg[129]) );
  DFF \ereg_reg[130]  ( .D(n3729), .CLK(clk), .RST(rst), .Q(ereg[130]) );
  DFF \ereg_reg[131]  ( .D(n3728), .CLK(clk), .RST(rst), .Q(ereg[131]) );
  DFF \ereg_reg[132]  ( .D(n3727), .CLK(clk), .RST(rst), .Q(ereg[132]) );
  DFF \ereg_reg[133]  ( .D(n3726), .CLK(clk), .RST(rst), .Q(ereg[133]) );
  DFF \ereg_reg[134]  ( .D(n3725), .CLK(clk), .RST(rst), .Q(ereg[134]) );
  DFF \ereg_reg[135]  ( .D(n3724), .CLK(clk), .RST(rst), .Q(ereg[135]) );
  DFF \ereg_reg[136]  ( .D(n3723), .CLK(clk), .RST(rst), .Q(ereg[136]) );
  DFF \ereg_reg[137]  ( .D(n3722), .CLK(clk), .RST(rst), .Q(ereg[137]) );
  DFF \ereg_reg[138]  ( .D(n3721), .CLK(clk), .RST(rst), .Q(ereg[138]) );
  DFF \ereg_reg[139]  ( .D(n3720), .CLK(clk), .RST(rst), .Q(ereg[139]) );
  DFF \ereg_reg[140]  ( .D(n3719), .CLK(clk), .RST(rst), .Q(ereg[140]) );
  DFF \ereg_reg[141]  ( .D(n3718), .CLK(clk), .RST(rst), .Q(ereg[141]) );
  DFF \ereg_reg[142]  ( .D(n3717), .CLK(clk), .RST(rst), .Q(ereg[142]) );
  DFF \ereg_reg[143]  ( .D(n3716), .CLK(clk), .RST(rst), .Q(ereg[143]) );
  DFF \ereg_reg[144]  ( .D(n3715), .CLK(clk), .RST(rst), .Q(ereg[144]) );
  DFF \ereg_reg[145]  ( .D(n3714), .CLK(clk), .RST(rst), .Q(ereg[145]) );
  DFF \ereg_reg[146]  ( .D(n3713), .CLK(clk), .RST(rst), .Q(ereg[146]) );
  DFF \ereg_reg[147]  ( .D(n3712), .CLK(clk), .RST(rst), .Q(ereg[147]) );
  DFF \ereg_reg[148]  ( .D(n3711), .CLK(clk), .RST(rst), .Q(ereg[148]) );
  DFF \ereg_reg[149]  ( .D(n3710), .CLK(clk), .RST(rst), .Q(ereg[149]) );
  DFF \ereg_reg[150]  ( .D(n3709), .CLK(clk), .RST(rst), .Q(ereg[150]) );
  DFF \ereg_reg[151]  ( .D(n3708), .CLK(clk), .RST(rst), .Q(ereg[151]) );
  DFF \ereg_reg[152]  ( .D(n3707), .CLK(clk), .RST(rst), .Q(ereg[152]) );
  DFF \ereg_reg[153]  ( .D(n3706), .CLK(clk), .RST(rst), .Q(ereg[153]) );
  DFF \ereg_reg[154]  ( .D(n3705), .CLK(clk), .RST(rst), .Q(ereg[154]) );
  DFF \ereg_reg[155]  ( .D(n3704), .CLK(clk), .RST(rst), .Q(ereg[155]) );
  DFF \ereg_reg[156]  ( .D(n3703), .CLK(clk), .RST(rst), .Q(ereg[156]) );
  DFF \ereg_reg[157]  ( .D(n3702), .CLK(clk), .RST(rst), .Q(ereg[157]) );
  DFF \ereg_reg[158]  ( .D(n3701), .CLK(clk), .RST(rst), .Q(ereg[158]) );
  DFF \ereg_reg[159]  ( .D(n3700), .CLK(clk), .RST(rst), .Q(ereg[159]) );
  DFF \ereg_reg[160]  ( .D(n3699), .CLK(clk), .RST(rst), .Q(ereg[160]) );
  DFF \ereg_reg[161]  ( .D(n3698), .CLK(clk), .RST(rst), .Q(ereg[161]) );
  DFF \ereg_reg[162]  ( .D(n3697), .CLK(clk), .RST(rst), .Q(ereg[162]) );
  DFF \ereg_reg[163]  ( .D(n3696), .CLK(clk), .RST(rst), .Q(ereg[163]) );
  DFF \ereg_reg[164]  ( .D(n3695), .CLK(clk), .RST(rst), .Q(ereg[164]) );
  DFF \ereg_reg[165]  ( .D(n3694), .CLK(clk), .RST(rst), .Q(ereg[165]) );
  DFF \ereg_reg[166]  ( .D(n3693), .CLK(clk), .RST(rst), .Q(ereg[166]) );
  DFF \ereg_reg[167]  ( .D(n3692), .CLK(clk), .RST(rst), .Q(ereg[167]) );
  DFF \ereg_reg[168]  ( .D(n3691), .CLK(clk), .RST(rst), .Q(ereg[168]) );
  DFF \ereg_reg[169]  ( .D(n3690), .CLK(clk), .RST(rst), .Q(ereg[169]) );
  DFF \ereg_reg[170]  ( .D(n3689), .CLK(clk), .RST(rst), .Q(ereg[170]) );
  DFF \ereg_reg[171]  ( .D(n3688), .CLK(clk), .RST(rst), .Q(ereg[171]) );
  DFF \ereg_reg[172]  ( .D(n3687), .CLK(clk), .RST(rst), .Q(ereg[172]) );
  DFF \ereg_reg[173]  ( .D(n3686), .CLK(clk), .RST(rst), .Q(ereg[173]) );
  DFF \ereg_reg[174]  ( .D(n3685), .CLK(clk), .RST(rst), .Q(ereg[174]) );
  DFF \ereg_reg[175]  ( .D(n3684), .CLK(clk), .RST(rst), .Q(ereg[175]) );
  DFF \ereg_reg[176]  ( .D(n3683), .CLK(clk), .RST(rst), .Q(ereg[176]) );
  DFF \ereg_reg[177]  ( .D(n3682), .CLK(clk), .RST(rst), .Q(ereg[177]) );
  DFF \ereg_reg[178]  ( .D(n3681), .CLK(clk), .RST(rst), .Q(ereg[178]) );
  DFF \ereg_reg[179]  ( .D(n3680), .CLK(clk), .RST(rst), .Q(ereg[179]) );
  DFF \ereg_reg[180]  ( .D(n3679), .CLK(clk), .RST(rst), .Q(ereg[180]) );
  DFF \ereg_reg[181]  ( .D(n3678), .CLK(clk), .RST(rst), .Q(ereg[181]) );
  DFF \ereg_reg[182]  ( .D(n3677), .CLK(clk), .RST(rst), .Q(ereg[182]) );
  DFF \ereg_reg[183]  ( .D(n3676), .CLK(clk), .RST(rst), .Q(ereg[183]) );
  DFF \ereg_reg[184]  ( .D(n3675), .CLK(clk), .RST(rst), .Q(ereg[184]) );
  DFF \ereg_reg[185]  ( .D(n3674), .CLK(clk), .RST(rst), .Q(ereg[185]) );
  DFF \ereg_reg[186]  ( .D(n3673), .CLK(clk), .RST(rst), .Q(ereg[186]) );
  DFF \ereg_reg[187]  ( .D(n3672), .CLK(clk), .RST(rst), .Q(ereg[187]) );
  DFF \ereg_reg[188]  ( .D(n3671), .CLK(clk), .RST(rst), .Q(ereg[188]) );
  DFF \ereg_reg[189]  ( .D(n3670), .CLK(clk), .RST(rst), .Q(ereg[189]) );
  DFF \ereg_reg[190]  ( .D(n3669), .CLK(clk), .RST(rst), .Q(ereg[190]) );
  DFF \ereg_reg[191]  ( .D(n3668), .CLK(clk), .RST(rst), .Q(ereg[191]) );
  DFF \ereg_reg[192]  ( .D(n3667), .CLK(clk), .RST(rst), .Q(ereg[192]) );
  DFF \ereg_reg[193]  ( .D(n3666), .CLK(clk), .RST(rst), .Q(ereg[193]) );
  DFF \ereg_reg[194]  ( .D(n3665), .CLK(clk), .RST(rst), .Q(ereg[194]) );
  DFF \ereg_reg[195]  ( .D(n3664), .CLK(clk), .RST(rst), .Q(ereg[195]) );
  DFF \ereg_reg[196]  ( .D(n3663), .CLK(clk), .RST(rst), .Q(ereg[196]) );
  DFF \ereg_reg[197]  ( .D(n3662), .CLK(clk), .RST(rst), .Q(ereg[197]) );
  DFF \ereg_reg[198]  ( .D(n3661), .CLK(clk), .RST(rst), .Q(ereg[198]) );
  DFF \ereg_reg[199]  ( .D(n3660), .CLK(clk), .RST(rst), .Q(ereg[199]) );
  DFF \ereg_reg[200]  ( .D(n3659), .CLK(clk), .RST(rst), .Q(ereg[200]) );
  DFF \ereg_reg[201]  ( .D(n3658), .CLK(clk), .RST(rst), .Q(ereg[201]) );
  DFF \ereg_reg[202]  ( .D(n3657), .CLK(clk), .RST(rst), .Q(ereg[202]) );
  DFF \ereg_reg[203]  ( .D(n3656), .CLK(clk), .RST(rst), .Q(ereg[203]) );
  DFF \ereg_reg[204]  ( .D(n3655), .CLK(clk), .RST(rst), .Q(ereg[204]) );
  DFF \ereg_reg[205]  ( .D(n3654), .CLK(clk), .RST(rst), .Q(ereg[205]) );
  DFF \ereg_reg[206]  ( .D(n3653), .CLK(clk), .RST(rst), .Q(ereg[206]) );
  DFF \ereg_reg[207]  ( .D(n3652), .CLK(clk), .RST(rst), .Q(ereg[207]) );
  DFF \ereg_reg[208]  ( .D(n3651), .CLK(clk), .RST(rst), .Q(ereg[208]) );
  DFF \ereg_reg[209]  ( .D(n3650), .CLK(clk), .RST(rst), .Q(ereg[209]) );
  DFF \ereg_reg[210]  ( .D(n3649), .CLK(clk), .RST(rst), .Q(ereg[210]) );
  DFF \ereg_reg[211]  ( .D(n3648), .CLK(clk), .RST(rst), .Q(ereg[211]) );
  DFF \ereg_reg[212]  ( .D(n3647), .CLK(clk), .RST(rst), .Q(ereg[212]) );
  DFF \ereg_reg[213]  ( .D(n3646), .CLK(clk), .RST(rst), .Q(ereg[213]) );
  DFF \ereg_reg[214]  ( .D(n3645), .CLK(clk), .RST(rst), .Q(ereg[214]) );
  DFF \ereg_reg[215]  ( .D(n3644), .CLK(clk), .RST(rst), .Q(ereg[215]) );
  DFF \ereg_reg[216]  ( .D(n3643), .CLK(clk), .RST(rst), .Q(ereg[216]) );
  DFF \ereg_reg[217]  ( .D(n3642), .CLK(clk), .RST(rst), .Q(ereg[217]) );
  DFF \ereg_reg[218]  ( .D(n3641), .CLK(clk), .RST(rst), .Q(ereg[218]) );
  DFF \ereg_reg[219]  ( .D(n3640), .CLK(clk), .RST(rst), .Q(ereg[219]) );
  DFF \ereg_reg[220]  ( .D(n3639), .CLK(clk), .RST(rst), .Q(ereg[220]) );
  DFF \ereg_reg[221]  ( .D(n3638), .CLK(clk), .RST(rst), .Q(ereg[221]) );
  DFF \ereg_reg[222]  ( .D(n3637), .CLK(clk), .RST(rst), .Q(ereg[222]) );
  DFF \ereg_reg[223]  ( .D(n3636), .CLK(clk), .RST(rst), .Q(ereg[223]) );
  DFF \ereg_reg[224]  ( .D(n3635), .CLK(clk), .RST(rst), .Q(ereg[224]) );
  DFF \ereg_reg[225]  ( .D(n3634), .CLK(clk), .RST(rst), .Q(ereg[225]) );
  DFF \ereg_reg[226]  ( .D(n3633), .CLK(clk), .RST(rst), .Q(ereg[226]) );
  DFF \ereg_reg[227]  ( .D(n3632), .CLK(clk), .RST(rst), .Q(ereg[227]) );
  DFF \ereg_reg[228]  ( .D(n3631), .CLK(clk), .RST(rst), .Q(ereg[228]) );
  DFF \ereg_reg[229]  ( .D(n3630), .CLK(clk), .RST(rst), .Q(ereg[229]) );
  DFF \ereg_reg[230]  ( .D(n3629), .CLK(clk), .RST(rst), .Q(ereg[230]) );
  DFF \ereg_reg[231]  ( .D(n3628), .CLK(clk), .RST(rst), .Q(ereg[231]) );
  DFF \ereg_reg[232]  ( .D(n3627), .CLK(clk), .RST(rst), .Q(ereg[232]) );
  DFF \ereg_reg[233]  ( .D(n3626), .CLK(clk), .RST(rst), .Q(ereg[233]) );
  DFF \ereg_reg[234]  ( .D(n3625), .CLK(clk), .RST(rst), .Q(ereg[234]) );
  DFF \ereg_reg[235]  ( .D(n3624), .CLK(clk), .RST(rst), .Q(ereg[235]) );
  DFF \ereg_reg[236]  ( .D(n3623), .CLK(clk), .RST(rst), .Q(ereg[236]) );
  DFF \ereg_reg[237]  ( .D(n3622), .CLK(clk), .RST(rst), .Q(ereg[237]) );
  DFF \ereg_reg[238]  ( .D(n3621), .CLK(clk), .RST(rst), .Q(ereg[238]) );
  DFF \ereg_reg[239]  ( .D(n3620), .CLK(clk), .RST(rst), .Q(ereg[239]) );
  DFF \ereg_reg[240]  ( .D(n3619), .CLK(clk), .RST(rst), .Q(ereg[240]) );
  DFF \ereg_reg[241]  ( .D(n3618), .CLK(clk), .RST(rst), .Q(ereg[241]) );
  DFF \ereg_reg[242]  ( .D(n3617), .CLK(clk), .RST(rst), .Q(ereg[242]) );
  DFF \ereg_reg[243]  ( .D(n3616), .CLK(clk), .RST(rst), .Q(ereg[243]) );
  DFF \ereg_reg[244]  ( .D(n3615), .CLK(clk), .RST(rst), .Q(ereg[244]) );
  DFF \ereg_reg[245]  ( .D(n3614), .CLK(clk), .RST(rst), .Q(ereg[245]) );
  DFF \ereg_reg[246]  ( .D(n3613), .CLK(clk), .RST(rst), .Q(ereg[246]) );
  DFF \ereg_reg[247]  ( .D(n3612), .CLK(clk), .RST(rst), .Q(ereg[247]) );
  DFF \ereg_reg[248]  ( .D(n3611), .CLK(clk), .RST(rst), .Q(ereg[248]) );
  DFF \ereg_reg[249]  ( .D(n3610), .CLK(clk), .RST(rst), .Q(ereg[249]) );
  DFF \ereg_reg[250]  ( .D(n3609), .CLK(clk), .RST(rst), .Q(ereg[250]) );
  DFF \ereg_reg[251]  ( .D(n3608), .CLK(clk), .RST(rst), .Q(ereg[251]) );
  DFF \ereg_reg[252]  ( .D(n3607), .CLK(clk), .RST(rst), .Q(ereg[252]) );
  DFF \ereg_reg[253]  ( .D(n3606), .CLK(clk), .RST(rst), .Q(ereg[253]) );
  DFF \ereg_reg[254]  ( .D(n3605), .CLK(clk), .RST(rst), .Q(ereg[254]) );
  DFF \ereg_reg[255]  ( .D(n3604), .CLK(clk), .RST(rst), .Q(ereg[255]) );
  DFF first_one_reg ( .D(n3347), .CLK(clk), .RST(rst), .Q(first_one) );
  DFF \creg_reg[0]  ( .D(n3602), .CLK(clk), .RST(rst), .Q(creg[0]) );
  DFF \creg_reg[1]  ( .D(n3601), .CLK(clk), .RST(rst), .Q(creg[1]) );
  DFF \creg_reg[2]  ( .D(n3600), .CLK(clk), .RST(rst), .Q(creg[2]) );
  DFF \creg_reg[3]  ( .D(n3599), .CLK(clk), .RST(rst), .Q(creg[3]) );
  DFF \creg_reg[4]  ( .D(n3598), .CLK(clk), .RST(rst), .Q(creg[4]) );
  DFF \creg_reg[5]  ( .D(n3597), .CLK(clk), .RST(rst), .Q(creg[5]) );
  DFF \creg_reg[6]  ( .D(n3596), .CLK(clk), .RST(rst), .Q(creg[6]) );
  DFF \creg_reg[7]  ( .D(n3595), .CLK(clk), .RST(rst), .Q(creg[7]) );
  DFF \creg_reg[8]  ( .D(n3594), .CLK(clk), .RST(rst), .Q(creg[8]) );
  DFF \creg_reg[9]  ( .D(n3593), .CLK(clk), .RST(rst), .Q(creg[9]) );
  DFF \creg_reg[10]  ( .D(n3592), .CLK(clk), .RST(rst), .Q(creg[10]) );
  DFF \creg_reg[11]  ( .D(n3591), .CLK(clk), .RST(rst), .Q(creg[11]) );
  DFF \creg_reg[12]  ( .D(n3590), .CLK(clk), .RST(rst), .Q(creg[12]) );
  DFF \creg_reg[13]  ( .D(n3589), .CLK(clk), .RST(rst), .Q(creg[13]) );
  DFF \creg_reg[14]  ( .D(n3588), .CLK(clk), .RST(rst), .Q(creg[14]) );
  DFF \creg_reg[15]  ( .D(n3587), .CLK(clk), .RST(rst), .Q(creg[15]) );
  DFF \creg_reg[16]  ( .D(n3586), .CLK(clk), .RST(rst), .Q(creg[16]) );
  DFF \creg_reg[17]  ( .D(n3585), .CLK(clk), .RST(rst), .Q(creg[17]) );
  DFF \creg_reg[18]  ( .D(n3584), .CLK(clk), .RST(rst), .Q(creg[18]) );
  DFF \creg_reg[19]  ( .D(n3583), .CLK(clk), .RST(rst), .Q(creg[19]) );
  DFF \creg_reg[20]  ( .D(n3582), .CLK(clk), .RST(rst), .Q(creg[20]) );
  DFF \creg_reg[21]  ( .D(n3581), .CLK(clk), .RST(rst), .Q(creg[21]) );
  DFF \creg_reg[22]  ( .D(n3580), .CLK(clk), .RST(rst), .Q(creg[22]) );
  DFF \creg_reg[23]  ( .D(n3579), .CLK(clk), .RST(rst), .Q(creg[23]) );
  DFF \creg_reg[24]  ( .D(n3578), .CLK(clk), .RST(rst), .Q(creg[24]) );
  DFF \creg_reg[25]  ( .D(n3577), .CLK(clk), .RST(rst), .Q(creg[25]) );
  DFF \creg_reg[26]  ( .D(n3576), .CLK(clk), .RST(rst), .Q(creg[26]) );
  DFF \creg_reg[27]  ( .D(n3575), .CLK(clk), .RST(rst), .Q(creg[27]) );
  DFF \creg_reg[28]  ( .D(n3574), .CLK(clk), .RST(rst), .Q(creg[28]) );
  DFF \creg_reg[29]  ( .D(n3573), .CLK(clk), .RST(rst), .Q(creg[29]) );
  DFF \creg_reg[30]  ( .D(n3572), .CLK(clk), .RST(rst), .Q(creg[30]) );
  DFF \creg_reg[31]  ( .D(n3571), .CLK(clk), .RST(rst), .Q(creg[31]) );
  DFF \creg_reg[32]  ( .D(n3570), .CLK(clk), .RST(rst), .Q(creg[32]) );
  DFF \creg_reg[33]  ( .D(n3569), .CLK(clk), .RST(rst), .Q(creg[33]) );
  DFF \creg_reg[34]  ( .D(n3568), .CLK(clk), .RST(rst), .Q(creg[34]) );
  DFF \creg_reg[35]  ( .D(n3567), .CLK(clk), .RST(rst), .Q(creg[35]) );
  DFF \creg_reg[36]  ( .D(n3566), .CLK(clk), .RST(rst), .Q(creg[36]) );
  DFF \creg_reg[37]  ( .D(n3565), .CLK(clk), .RST(rst), .Q(creg[37]) );
  DFF \creg_reg[38]  ( .D(n3564), .CLK(clk), .RST(rst), .Q(creg[38]) );
  DFF \creg_reg[39]  ( .D(n3563), .CLK(clk), .RST(rst), .Q(creg[39]) );
  DFF \creg_reg[40]  ( .D(n3562), .CLK(clk), .RST(rst), .Q(creg[40]) );
  DFF \creg_reg[41]  ( .D(n3561), .CLK(clk), .RST(rst), .Q(creg[41]) );
  DFF \creg_reg[42]  ( .D(n3560), .CLK(clk), .RST(rst), .Q(creg[42]) );
  DFF \creg_reg[43]  ( .D(n3559), .CLK(clk), .RST(rst), .Q(creg[43]) );
  DFF \creg_reg[44]  ( .D(n3558), .CLK(clk), .RST(rst), .Q(creg[44]) );
  DFF \creg_reg[45]  ( .D(n3557), .CLK(clk), .RST(rst), .Q(creg[45]) );
  DFF \creg_reg[46]  ( .D(n3556), .CLK(clk), .RST(rst), .Q(creg[46]) );
  DFF \creg_reg[47]  ( .D(n3555), .CLK(clk), .RST(rst), .Q(creg[47]) );
  DFF \creg_reg[48]  ( .D(n3554), .CLK(clk), .RST(rst), .Q(creg[48]) );
  DFF \creg_reg[49]  ( .D(n3553), .CLK(clk), .RST(rst), .Q(creg[49]) );
  DFF \creg_reg[50]  ( .D(n3552), .CLK(clk), .RST(rst), .Q(creg[50]) );
  DFF \creg_reg[51]  ( .D(n3551), .CLK(clk), .RST(rst), .Q(creg[51]) );
  DFF \creg_reg[52]  ( .D(n3550), .CLK(clk), .RST(rst), .Q(creg[52]) );
  DFF \creg_reg[53]  ( .D(n3549), .CLK(clk), .RST(rst), .Q(creg[53]) );
  DFF \creg_reg[54]  ( .D(n3548), .CLK(clk), .RST(rst), .Q(creg[54]) );
  DFF \creg_reg[55]  ( .D(n3547), .CLK(clk), .RST(rst), .Q(creg[55]) );
  DFF \creg_reg[56]  ( .D(n3546), .CLK(clk), .RST(rst), .Q(creg[56]) );
  DFF \creg_reg[57]  ( .D(n3545), .CLK(clk), .RST(rst), .Q(creg[57]) );
  DFF \creg_reg[58]  ( .D(n3544), .CLK(clk), .RST(rst), .Q(creg[58]) );
  DFF \creg_reg[59]  ( .D(n3543), .CLK(clk), .RST(rst), .Q(creg[59]) );
  DFF \creg_reg[60]  ( .D(n3542), .CLK(clk), .RST(rst), .Q(creg[60]) );
  DFF \creg_reg[61]  ( .D(n3541), .CLK(clk), .RST(rst), .Q(creg[61]) );
  DFF \creg_reg[62]  ( .D(n3540), .CLK(clk), .RST(rst), .Q(creg[62]) );
  DFF \creg_reg[63]  ( .D(n3539), .CLK(clk), .RST(rst), .Q(creg[63]) );
  DFF \creg_reg[64]  ( .D(n3538), .CLK(clk), .RST(rst), .Q(creg[64]) );
  DFF \creg_reg[65]  ( .D(n3537), .CLK(clk), .RST(rst), .Q(creg[65]) );
  DFF \creg_reg[66]  ( .D(n3536), .CLK(clk), .RST(rst), .Q(creg[66]) );
  DFF \creg_reg[67]  ( .D(n3535), .CLK(clk), .RST(rst), .Q(creg[67]) );
  DFF \creg_reg[68]  ( .D(n3534), .CLK(clk), .RST(rst), .Q(creg[68]) );
  DFF \creg_reg[69]  ( .D(n3533), .CLK(clk), .RST(rst), .Q(creg[69]) );
  DFF \creg_reg[70]  ( .D(n3532), .CLK(clk), .RST(rst), .Q(creg[70]) );
  DFF \creg_reg[71]  ( .D(n3531), .CLK(clk), .RST(rst), .Q(creg[71]) );
  DFF \creg_reg[72]  ( .D(n3530), .CLK(clk), .RST(rst), .Q(creg[72]) );
  DFF \creg_reg[73]  ( .D(n3529), .CLK(clk), .RST(rst), .Q(creg[73]) );
  DFF \creg_reg[74]  ( .D(n3528), .CLK(clk), .RST(rst), .Q(creg[74]) );
  DFF \creg_reg[75]  ( .D(n3527), .CLK(clk), .RST(rst), .Q(creg[75]) );
  DFF \creg_reg[76]  ( .D(n3526), .CLK(clk), .RST(rst), .Q(creg[76]) );
  DFF \creg_reg[77]  ( .D(n3525), .CLK(clk), .RST(rst), .Q(creg[77]) );
  DFF \creg_reg[78]  ( .D(n3524), .CLK(clk), .RST(rst), .Q(creg[78]) );
  DFF \creg_reg[79]  ( .D(n3523), .CLK(clk), .RST(rst), .Q(creg[79]) );
  DFF \creg_reg[80]  ( .D(n3522), .CLK(clk), .RST(rst), .Q(creg[80]) );
  DFF \creg_reg[81]  ( .D(n3521), .CLK(clk), .RST(rst), .Q(creg[81]) );
  DFF \creg_reg[82]  ( .D(n3520), .CLK(clk), .RST(rst), .Q(creg[82]) );
  DFF \creg_reg[83]  ( .D(n3519), .CLK(clk), .RST(rst), .Q(creg[83]) );
  DFF \creg_reg[84]  ( .D(n3518), .CLK(clk), .RST(rst), .Q(creg[84]) );
  DFF \creg_reg[85]  ( .D(n3517), .CLK(clk), .RST(rst), .Q(creg[85]) );
  DFF \creg_reg[86]  ( .D(n3516), .CLK(clk), .RST(rst), .Q(creg[86]) );
  DFF \creg_reg[87]  ( .D(n3515), .CLK(clk), .RST(rst), .Q(creg[87]) );
  DFF \creg_reg[88]  ( .D(n3514), .CLK(clk), .RST(rst), .Q(creg[88]) );
  DFF \creg_reg[89]  ( .D(n3513), .CLK(clk), .RST(rst), .Q(creg[89]) );
  DFF \creg_reg[90]  ( .D(n3512), .CLK(clk), .RST(rst), .Q(creg[90]) );
  DFF \creg_reg[91]  ( .D(n3511), .CLK(clk), .RST(rst), .Q(creg[91]) );
  DFF \creg_reg[92]  ( .D(n3510), .CLK(clk), .RST(rst), .Q(creg[92]) );
  DFF \creg_reg[93]  ( .D(n3509), .CLK(clk), .RST(rst), .Q(creg[93]) );
  DFF \creg_reg[94]  ( .D(n3508), .CLK(clk), .RST(rst), .Q(creg[94]) );
  DFF \creg_reg[95]  ( .D(n3507), .CLK(clk), .RST(rst), .Q(creg[95]) );
  DFF \creg_reg[96]  ( .D(n3506), .CLK(clk), .RST(rst), .Q(creg[96]) );
  DFF \creg_reg[97]  ( .D(n3505), .CLK(clk), .RST(rst), .Q(creg[97]) );
  DFF \creg_reg[98]  ( .D(n3504), .CLK(clk), .RST(rst), .Q(creg[98]) );
  DFF \creg_reg[99]  ( .D(n3503), .CLK(clk), .RST(rst), .Q(creg[99]) );
  DFF \creg_reg[100]  ( .D(n3502), .CLK(clk), .RST(rst), .Q(creg[100]) );
  DFF \creg_reg[101]  ( .D(n3501), .CLK(clk), .RST(rst), .Q(creg[101]) );
  DFF \creg_reg[102]  ( .D(n3500), .CLK(clk), .RST(rst), .Q(creg[102]) );
  DFF \creg_reg[103]  ( .D(n3499), .CLK(clk), .RST(rst), .Q(creg[103]) );
  DFF \creg_reg[104]  ( .D(n3498), .CLK(clk), .RST(rst), .Q(creg[104]) );
  DFF \creg_reg[105]  ( .D(n3497), .CLK(clk), .RST(rst), .Q(creg[105]) );
  DFF \creg_reg[106]  ( .D(n3496), .CLK(clk), .RST(rst), .Q(creg[106]) );
  DFF \creg_reg[107]  ( .D(n3495), .CLK(clk), .RST(rst), .Q(creg[107]) );
  DFF \creg_reg[108]  ( .D(n3494), .CLK(clk), .RST(rst), .Q(creg[108]) );
  DFF \creg_reg[109]  ( .D(n3493), .CLK(clk), .RST(rst), .Q(creg[109]) );
  DFF \creg_reg[110]  ( .D(n3492), .CLK(clk), .RST(rst), .Q(creg[110]) );
  DFF \creg_reg[111]  ( .D(n3491), .CLK(clk), .RST(rst), .Q(creg[111]) );
  DFF \creg_reg[112]  ( .D(n3490), .CLK(clk), .RST(rst), .Q(creg[112]) );
  DFF \creg_reg[113]  ( .D(n3489), .CLK(clk), .RST(rst), .Q(creg[113]) );
  DFF \creg_reg[114]  ( .D(n3488), .CLK(clk), .RST(rst), .Q(creg[114]) );
  DFF \creg_reg[115]  ( .D(n3487), .CLK(clk), .RST(rst), .Q(creg[115]) );
  DFF \creg_reg[116]  ( .D(n3486), .CLK(clk), .RST(rst), .Q(creg[116]) );
  DFF \creg_reg[117]  ( .D(n3485), .CLK(clk), .RST(rst), .Q(creg[117]) );
  DFF \creg_reg[118]  ( .D(n3484), .CLK(clk), .RST(rst), .Q(creg[118]) );
  DFF \creg_reg[119]  ( .D(n3483), .CLK(clk), .RST(rst), .Q(creg[119]) );
  DFF \creg_reg[120]  ( .D(n3482), .CLK(clk), .RST(rst), .Q(creg[120]) );
  DFF \creg_reg[121]  ( .D(n3481), .CLK(clk), .RST(rst), .Q(creg[121]) );
  DFF \creg_reg[122]  ( .D(n3480), .CLK(clk), .RST(rst), .Q(creg[122]) );
  DFF \creg_reg[123]  ( .D(n3479), .CLK(clk), .RST(rst), .Q(creg[123]) );
  DFF \creg_reg[124]  ( .D(n3478), .CLK(clk), .RST(rst), .Q(creg[124]) );
  DFF \creg_reg[125]  ( .D(n3477), .CLK(clk), .RST(rst), .Q(creg[125]) );
  DFF \creg_reg[126]  ( .D(n3476), .CLK(clk), .RST(rst), .Q(creg[126]) );
  DFF \creg_reg[127]  ( .D(n3475), .CLK(clk), .RST(rst), .Q(creg[127]) );
  DFF \creg_reg[128]  ( .D(n3474), .CLK(clk), .RST(rst), .Q(creg[128]) );
  DFF \creg_reg[129]  ( .D(n3473), .CLK(clk), .RST(rst), .Q(creg[129]) );
  DFF \creg_reg[130]  ( .D(n3472), .CLK(clk), .RST(rst), .Q(creg[130]) );
  DFF \creg_reg[131]  ( .D(n3471), .CLK(clk), .RST(rst), .Q(creg[131]) );
  DFF \creg_reg[132]  ( .D(n3470), .CLK(clk), .RST(rst), .Q(creg[132]) );
  DFF \creg_reg[133]  ( .D(n3469), .CLK(clk), .RST(rst), .Q(creg[133]) );
  DFF \creg_reg[134]  ( .D(n3468), .CLK(clk), .RST(rst), .Q(creg[134]) );
  DFF \creg_reg[135]  ( .D(n3467), .CLK(clk), .RST(rst), .Q(creg[135]) );
  DFF \creg_reg[136]  ( .D(n3466), .CLK(clk), .RST(rst), .Q(creg[136]) );
  DFF \creg_reg[137]  ( .D(n3465), .CLK(clk), .RST(rst), .Q(creg[137]) );
  DFF \creg_reg[138]  ( .D(n3464), .CLK(clk), .RST(rst), .Q(creg[138]) );
  DFF \creg_reg[139]  ( .D(n3463), .CLK(clk), .RST(rst), .Q(creg[139]) );
  DFF \creg_reg[140]  ( .D(n3462), .CLK(clk), .RST(rst), .Q(creg[140]) );
  DFF \creg_reg[141]  ( .D(n3461), .CLK(clk), .RST(rst), .Q(creg[141]) );
  DFF \creg_reg[142]  ( .D(n3460), .CLK(clk), .RST(rst), .Q(creg[142]) );
  DFF \creg_reg[143]  ( .D(n3459), .CLK(clk), .RST(rst), .Q(creg[143]) );
  DFF \creg_reg[144]  ( .D(n3458), .CLK(clk), .RST(rst), .Q(creg[144]) );
  DFF \creg_reg[145]  ( .D(n3457), .CLK(clk), .RST(rst), .Q(creg[145]) );
  DFF \creg_reg[146]  ( .D(n3456), .CLK(clk), .RST(rst), .Q(creg[146]) );
  DFF \creg_reg[147]  ( .D(n3455), .CLK(clk), .RST(rst), .Q(creg[147]) );
  DFF \creg_reg[148]  ( .D(n3454), .CLK(clk), .RST(rst), .Q(creg[148]) );
  DFF \creg_reg[149]  ( .D(n3453), .CLK(clk), .RST(rst), .Q(creg[149]) );
  DFF \creg_reg[150]  ( .D(n3452), .CLK(clk), .RST(rst), .Q(creg[150]) );
  DFF \creg_reg[151]  ( .D(n3451), .CLK(clk), .RST(rst), .Q(creg[151]) );
  DFF \creg_reg[152]  ( .D(n3450), .CLK(clk), .RST(rst), .Q(creg[152]) );
  DFF \creg_reg[153]  ( .D(n3449), .CLK(clk), .RST(rst), .Q(creg[153]) );
  DFF \creg_reg[154]  ( .D(n3448), .CLK(clk), .RST(rst), .Q(creg[154]) );
  DFF \creg_reg[155]  ( .D(n3447), .CLK(clk), .RST(rst), .Q(creg[155]) );
  DFF \creg_reg[156]  ( .D(n3446), .CLK(clk), .RST(rst), .Q(creg[156]) );
  DFF \creg_reg[157]  ( .D(n3445), .CLK(clk), .RST(rst), .Q(creg[157]) );
  DFF \creg_reg[158]  ( .D(n3444), .CLK(clk), .RST(rst), .Q(creg[158]) );
  DFF \creg_reg[159]  ( .D(n3443), .CLK(clk), .RST(rst), .Q(creg[159]) );
  DFF \creg_reg[160]  ( .D(n3442), .CLK(clk), .RST(rst), .Q(creg[160]) );
  DFF \creg_reg[161]  ( .D(n3441), .CLK(clk), .RST(rst), .Q(creg[161]) );
  DFF \creg_reg[162]  ( .D(n3440), .CLK(clk), .RST(rst), .Q(creg[162]) );
  DFF \creg_reg[163]  ( .D(n3439), .CLK(clk), .RST(rst), .Q(creg[163]) );
  DFF \creg_reg[164]  ( .D(n3438), .CLK(clk), .RST(rst), .Q(creg[164]) );
  DFF \creg_reg[165]  ( .D(n3437), .CLK(clk), .RST(rst), .Q(creg[165]) );
  DFF \creg_reg[166]  ( .D(n3436), .CLK(clk), .RST(rst), .Q(creg[166]) );
  DFF \creg_reg[167]  ( .D(n3435), .CLK(clk), .RST(rst), .Q(creg[167]) );
  DFF \creg_reg[168]  ( .D(n3434), .CLK(clk), .RST(rst), .Q(creg[168]) );
  DFF \creg_reg[169]  ( .D(n3433), .CLK(clk), .RST(rst), .Q(creg[169]) );
  DFF \creg_reg[170]  ( .D(n3432), .CLK(clk), .RST(rst), .Q(creg[170]) );
  DFF \creg_reg[171]  ( .D(n3431), .CLK(clk), .RST(rst), .Q(creg[171]) );
  DFF \creg_reg[172]  ( .D(n3430), .CLK(clk), .RST(rst), .Q(creg[172]) );
  DFF \creg_reg[173]  ( .D(n3429), .CLK(clk), .RST(rst), .Q(creg[173]) );
  DFF \creg_reg[174]  ( .D(n3428), .CLK(clk), .RST(rst), .Q(creg[174]) );
  DFF \creg_reg[175]  ( .D(n3427), .CLK(clk), .RST(rst), .Q(creg[175]) );
  DFF \creg_reg[176]  ( .D(n3426), .CLK(clk), .RST(rst), .Q(creg[176]) );
  DFF \creg_reg[177]  ( .D(n3425), .CLK(clk), .RST(rst), .Q(creg[177]) );
  DFF \creg_reg[178]  ( .D(n3424), .CLK(clk), .RST(rst), .Q(creg[178]) );
  DFF \creg_reg[179]  ( .D(n3423), .CLK(clk), .RST(rst), .Q(creg[179]) );
  DFF \creg_reg[180]  ( .D(n3422), .CLK(clk), .RST(rst), .Q(creg[180]) );
  DFF \creg_reg[181]  ( .D(n3421), .CLK(clk), .RST(rst), .Q(creg[181]) );
  DFF \creg_reg[182]  ( .D(n3420), .CLK(clk), .RST(rst), .Q(creg[182]) );
  DFF \creg_reg[183]  ( .D(n3419), .CLK(clk), .RST(rst), .Q(creg[183]) );
  DFF \creg_reg[184]  ( .D(n3418), .CLK(clk), .RST(rst), .Q(creg[184]) );
  DFF \creg_reg[185]  ( .D(n3417), .CLK(clk), .RST(rst), .Q(creg[185]) );
  DFF \creg_reg[186]  ( .D(n3416), .CLK(clk), .RST(rst), .Q(creg[186]) );
  DFF \creg_reg[187]  ( .D(n3415), .CLK(clk), .RST(rst), .Q(creg[187]) );
  DFF \creg_reg[188]  ( .D(n3414), .CLK(clk), .RST(rst), .Q(creg[188]) );
  DFF \creg_reg[189]  ( .D(n3413), .CLK(clk), .RST(rst), .Q(creg[189]) );
  DFF \creg_reg[190]  ( .D(n3412), .CLK(clk), .RST(rst), .Q(creg[190]) );
  DFF \creg_reg[191]  ( .D(n3411), .CLK(clk), .RST(rst), .Q(creg[191]) );
  DFF \creg_reg[192]  ( .D(n3410), .CLK(clk), .RST(rst), .Q(creg[192]) );
  DFF \creg_reg[193]  ( .D(n3409), .CLK(clk), .RST(rst), .Q(creg[193]) );
  DFF \creg_reg[194]  ( .D(n3408), .CLK(clk), .RST(rst), .Q(creg[194]) );
  DFF \creg_reg[195]  ( .D(n3407), .CLK(clk), .RST(rst), .Q(creg[195]) );
  DFF \creg_reg[196]  ( .D(n3406), .CLK(clk), .RST(rst), .Q(creg[196]) );
  DFF \creg_reg[197]  ( .D(n3405), .CLK(clk), .RST(rst), .Q(creg[197]) );
  DFF \creg_reg[198]  ( .D(n3404), .CLK(clk), .RST(rst), .Q(creg[198]) );
  DFF \creg_reg[199]  ( .D(n3403), .CLK(clk), .RST(rst), .Q(creg[199]) );
  DFF \creg_reg[200]  ( .D(n3402), .CLK(clk), .RST(rst), .Q(creg[200]) );
  DFF \creg_reg[201]  ( .D(n3401), .CLK(clk), .RST(rst), .Q(creg[201]) );
  DFF \creg_reg[202]  ( .D(n3400), .CLK(clk), .RST(rst), .Q(creg[202]) );
  DFF \creg_reg[203]  ( .D(n3399), .CLK(clk), .RST(rst), .Q(creg[203]) );
  DFF \creg_reg[204]  ( .D(n3398), .CLK(clk), .RST(rst), .Q(creg[204]) );
  DFF \creg_reg[205]  ( .D(n3397), .CLK(clk), .RST(rst), .Q(creg[205]) );
  DFF \creg_reg[206]  ( .D(n3396), .CLK(clk), .RST(rst), .Q(creg[206]) );
  DFF \creg_reg[207]  ( .D(n3395), .CLK(clk), .RST(rst), .Q(creg[207]) );
  DFF \creg_reg[208]  ( .D(n3394), .CLK(clk), .RST(rst), .Q(creg[208]) );
  DFF \creg_reg[209]  ( .D(n3393), .CLK(clk), .RST(rst), .Q(creg[209]) );
  DFF \creg_reg[210]  ( .D(n3392), .CLK(clk), .RST(rst), .Q(creg[210]) );
  DFF \creg_reg[211]  ( .D(n3391), .CLK(clk), .RST(rst), .Q(creg[211]) );
  DFF \creg_reg[212]  ( .D(n3390), .CLK(clk), .RST(rst), .Q(creg[212]) );
  DFF \creg_reg[213]  ( .D(n3389), .CLK(clk), .RST(rst), .Q(creg[213]) );
  DFF \creg_reg[214]  ( .D(n3388), .CLK(clk), .RST(rst), .Q(creg[214]) );
  DFF \creg_reg[215]  ( .D(n3387), .CLK(clk), .RST(rst), .Q(creg[215]) );
  DFF \creg_reg[216]  ( .D(n3386), .CLK(clk), .RST(rst), .Q(creg[216]) );
  DFF \creg_reg[217]  ( .D(n3385), .CLK(clk), .RST(rst), .Q(creg[217]) );
  DFF \creg_reg[218]  ( .D(n3384), .CLK(clk), .RST(rst), .Q(creg[218]) );
  DFF \creg_reg[219]  ( .D(n3383), .CLK(clk), .RST(rst), .Q(creg[219]) );
  DFF \creg_reg[220]  ( .D(n3382), .CLK(clk), .RST(rst), .Q(creg[220]) );
  DFF \creg_reg[221]  ( .D(n3381), .CLK(clk), .RST(rst), .Q(creg[221]) );
  DFF \creg_reg[222]  ( .D(n3380), .CLK(clk), .RST(rst), .Q(creg[222]) );
  DFF \creg_reg[223]  ( .D(n3379), .CLK(clk), .RST(rst), .Q(creg[223]) );
  DFF \creg_reg[224]  ( .D(n3378), .CLK(clk), .RST(rst), .Q(creg[224]) );
  DFF \creg_reg[225]  ( .D(n3377), .CLK(clk), .RST(rst), .Q(creg[225]) );
  DFF \creg_reg[226]  ( .D(n3376), .CLK(clk), .RST(rst), .Q(creg[226]) );
  DFF \creg_reg[227]  ( .D(n3375), .CLK(clk), .RST(rst), .Q(creg[227]) );
  DFF \creg_reg[228]  ( .D(n3374), .CLK(clk), .RST(rst), .Q(creg[228]) );
  DFF \creg_reg[229]  ( .D(n3373), .CLK(clk), .RST(rst), .Q(creg[229]) );
  DFF \creg_reg[230]  ( .D(n3372), .CLK(clk), .RST(rst), .Q(creg[230]) );
  DFF \creg_reg[231]  ( .D(n3371), .CLK(clk), .RST(rst), .Q(creg[231]) );
  DFF \creg_reg[232]  ( .D(n3370), .CLK(clk), .RST(rst), .Q(creg[232]) );
  DFF \creg_reg[233]  ( .D(n3369), .CLK(clk), .RST(rst), .Q(creg[233]) );
  DFF \creg_reg[234]  ( .D(n3368), .CLK(clk), .RST(rst), .Q(creg[234]) );
  DFF \creg_reg[235]  ( .D(n3367), .CLK(clk), .RST(rst), .Q(creg[235]) );
  DFF \creg_reg[236]  ( .D(n3366), .CLK(clk), .RST(rst), .Q(creg[236]) );
  DFF \creg_reg[237]  ( .D(n3365), .CLK(clk), .RST(rst), .Q(creg[237]) );
  DFF \creg_reg[238]  ( .D(n3364), .CLK(clk), .RST(rst), .Q(creg[238]) );
  DFF \creg_reg[239]  ( .D(n3363), .CLK(clk), .RST(rst), .Q(creg[239]) );
  DFF \creg_reg[240]  ( .D(n3362), .CLK(clk), .RST(rst), .Q(creg[240]) );
  DFF \creg_reg[241]  ( .D(n3361), .CLK(clk), .RST(rst), .Q(creg[241]) );
  DFF \creg_reg[242]  ( .D(n3360), .CLK(clk), .RST(rst), .Q(creg[242]) );
  DFF \creg_reg[243]  ( .D(n3359), .CLK(clk), .RST(rst), .Q(creg[243]) );
  DFF \creg_reg[244]  ( .D(n3358), .CLK(clk), .RST(rst), .Q(creg[244]) );
  DFF \creg_reg[245]  ( .D(n3357), .CLK(clk), .RST(rst), .Q(creg[245]) );
  DFF \creg_reg[246]  ( .D(n3356), .CLK(clk), .RST(rst), .Q(creg[246]) );
  DFF \creg_reg[247]  ( .D(n3355), .CLK(clk), .RST(rst), .Q(creg[247]) );
  DFF \creg_reg[248]  ( .D(n3354), .CLK(clk), .RST(rst), .Q(creg[248]) );
  DFF \creg_reg[249]  ( .D(n3353), .CLK(clk), .RST(rst), .Q(creg[249]) );
  DFF \creg_reg[250]  ( .D(n3352), .CLK(clk), .RST(rst), .Q(creg[250]) );
  DFF \creg_reg[251]  ( .D(n3351), .CLK(clk), .RST(rst), .Q(creg[251]) );
  DFF \creg_reg[252]  ( .D(n3350), .CLK(clk), .RST(rst), .Q(creg[252]) );
  DFF \creg_reg[253]  ( .D(n3349), .CLK(clk), .RST(rst), .Q(creg[253]) );
  DFF \creg_reg[254]  ( .D(n3348), .CLK(clk), .RST(rst), .Q(creg[254]) );
  DFF \creg_reg[255]  ( .D(n3603), .CLK(clk), .RST(rst), .Q(creg[255]) );
  NAND U5655 ( .A(n3861), .B(n3862), .Z(y[9]) );
  NANDN U5656 ( .A(n3863), .B(m[9]), .Z(n3862) );
  NANDN U5657 ( .A(n3864), .B(creg[9]), .Z(n3861) );
  NAND U5658 ( .A(n3865), .B(n3866), .Z(y[99]) );
  NANDN U5659 ( .A(n3863), .B(m[99]), .Z(n3866) );
  NANDN U5660 ( .A(n3864), .B(creg[99]), .Z(n3865) );
  NAND U5661 ( .A(n3867), .B(n3868), .Z(y[98]) );
  NANDN U5662 ( .A(n3863), .B(m[98]), .Z(n3868) );
  NANDN U5663 ( .A(n3864), .B(creg[98]), .Z(n3867) );
  NAND U5664 ( .A(n3869), .B(n3870), .Z(y[97]) );
  NANDN U5665 ( .A(n3863), .B(m[97]), .Z(n3870) );
  NANDN U5666 ( .A(n3864), .B(creg[97]), .Z(n3869) );
  NAND U5667 ( .A(n3871), .B(n3872), .Z(y[96]) );
  NANDN U5668 ( .A(n3863), .B(m[96]), .Z(n3872) );
  NANDN U5669 ( .A(n3864), .B(creg[96]), .Z(n3871) );
  NAND U5670 ( .A(n3873), .B(n3874), .Z(y[95]) );
  NANDN U5671 ( .A(n3863), .B(m[95]), .Z(n3874) );
  NANDN U5672 ( .A(n3864), .B(creg[95]), .Z(n3873) );
  NAND U5673 ( .A(n3875), .B(n3876), .Z(y[94]) );
  NANDN U5674 ( .A(n3863), .B(m[94]), .Z(n3876) );
  NANDN U5675 ( .A(n3864), .B(creg[94]), .Z(n3875) );
  NAND U5676 ( .A(n3877), .B(n3878), .Z(y[93]) );
  NANDN U5677 ( .A(n3863), .B(m[93]), .Z(n3878) );
  NANDN U5678 ( .A(n3864), .B(creg[93]), .Z(n3877) );
  NAND U5679 ( .A(n3879), .B(n3880), .Z(y[92]) );
  NANDN U5680 ( .A(n3863), .B(m[92]), .Z(n3880) );
  NANDN U5681 ( .A(n3864), .B(creg[92]), .Z(n3879) );
  NAND U5682 ( .A(n3881), .B(n3882), .Z(y[91]) );
  NANDN U5683 ( .A(n3863), .B(m[91]), .Z(n3882) );
  NANDN U5684 ( .A(n3864), .B(creg[91]), .Z(n3881) );
  NAND U5685 ( .A(n3883), .B(n3884), .Z(y[90]) );
  NANDN U5686 ( .A(n3863), .B(m[90]), .Z(n3884) );
  NANDN U5687 ( .A(n3864), .B(creg[90]), .Z(n3883) );
  NAND U5688 ( .A(n3885), .B(n3886), .Z(y[8]) );
  NANDN U5689 ( .A(n3863), .B(m[8]), .Z(n3886) );
  NANDN U5690 ( .A(n3864), .B(creg[8]), .Z(n3885) );
  NAND U5691 ( .A(n3887), .B(n3888), .Z(y[89]) );
  NANDN U5692 ( .A(n3863), .B(m[89]), .Z(n3888) );
  NANDN U5693 ( .A(n3864), .B(creg[89]), .Z(n3887) );
  NAND U5694 ( .A(n3889), .B(n3890), .Z(y[88]) );
  NANDN U5695 ( .A(n3863), .B(m[88]), .Z(n3890) );
  NANDN U5696 ( .A(n3864), .B(creg[88]), .Z(n3889) );
  NAND U5697 ( .A(n3891), .B(n3892), .Z(y[87]) );
  NANDN U5698 ( .A(n3863), .B(m[87]), .Z(n3892) );
  NANDN U5699 ( .A(n3864), .B(creg[87]), .Z(n3891) );
  NAND U5700 ( .A(n3893), .B(n3894), .Z(y[86]) );
  NANDN U5701 ( .A(n3863), .B(m[86]), .Z(n3894) );
  NANDN U5702 ( .A(n3864), .B(creg[86]), .Z(n3893) );
  NAND U5703 ( .A(n3895), .B(n3896), .Z(y[85]) );
  NANDN U5704 ( .A(n3863), .B(m[85]), .Z(n3896) );
  NANDN U5705 ( .A(n3864), .B(creg[85]), .Z(n3895) );
  NAND U5706 ( .A(n3897), .B(n3898), .Z(y[84]) );
  NANDN U5707 ( .A(n3863), .B(m[84]), .Z(n3898) );
  NANDN U5708 ( .A(n3864), .B(creg[84]), .Z(n3897) );
  NAND U5709 ( .A(n3899), .B(n3900), .Z(y[83]) );
  NANDN U5710 ( .A(n3863), .B(m[83]), .Z(n3900) );
  NANDN U5711 ( .A(n3864), .B(creg[83]), .Z(n3899) );
  NAND U5712 ( .A(n3901), .B(n3902), .Z(y[82]) );
  NANDN U5713 ( .A(n3863), .B(m[82]), .Z(n3902) );
  NANDN U5714 ( .A(n3864), .B(creg[82]), .Z(n3901) );
  NAND U5715 ( .A(n3903), .B(n3904), .Z(y[81]) );
  NANDN U5716 ( .A(n3863), .B(m[81]), .Z(n3904) );
  NANDN U5717 ( .A(n3864), .B(creg[81]), .Z(n3903) );
  NAND U5718 ( .A(n3905), .B(n3906), .Z(y[80]) );
  NANDN U5719 ( .A(n3863), .B(m[80]), .Z(n3906) );
  NANDN U5720 ( .A(n3864), .B(creg[80]), .Z(n3905) );
  NAND U5721 ( .A(n3907), .B(n3908), .Z(y[7]) );
  NANDN U5722 ( .A(n3863), .B(m[7]), .Z(n3908) );
  NANDN U5723 ( .A(n3864), .B(creg[7]), .Z(n3907) );
  NAND U5724 ( .A(n3909), .B(n3910), .Z(y[79]) );
  NANDN U5725 ( .A(n3863), .B(m[79]), .Z(n3910) );
  NANDN U5726 ( .A(n3864), .B(creg[79]), .Z(n3909) );
  NAND U5727 ( .A(n3911), .B(n3912), .Z(y[78]) );
  NANDN U5728 ( .A(n3863), .B(m[78]), .Z(n3912) );
  NANDN U5729 ( .A(n3864), .B(creg[78]), .Z(n3911) );
  NAND U5730 ( .A(n3913), .B(n3914), .Z(y[77]) );
  NANDN U5731 ( .A(n3863), .B(m[77]), .Z(n3914) );
  NANDN U5732 ( .A(n3864), .B(creg[77]), .Z(n3913) );
  NAND U5733 ( .A(n3915), .B(n3916), .Z(y[76]) );
  NANDN U5734 ( .A(n3863), .B(m[76]), .Z(n3916) );
  NANDN U5735 ( .A(n3864), .B(creg[76]), .Z(n3915) );
  NAND U5736 ( .A(n3917), .B(n3918), .Z(y[75]) );
  NANDN U5737 ( .A(n3863), .B(m[75]), .Z(n3918) );
  NANDN U5738 ( .A(n3864), .B(creg[75]), .Z(n3917) );
  NAND U5739 ( .A(n3919), .B(n3920), .Z(y[74]) );
  NANDN U5740 ( .A(n3863), .B(m[74]), .Z(n3920) );
  NANDN U5741 ( .A(n3864), .B(creg[74]), .Z(n3919) );
  NAND U5742 ( .A(n3921), .B(n3922), .Z(y[73]) );
  NANDN U5743 ( .A(n3863), .B(m[73]), .Z(n3922) );
  NANDN U5744 ( .A(n3864), .B(creg[73]), .Z(n3921) );
  NAND U5745 ( .A(n3923), .B(n3924), .Z(y[72]) );
  NANDN U5746 ( .A(n3863), .B(m[72]), .Z(n3924) );
  NANDN U5747 ( .A(n3864), .B(creg[72]), .Z(n3923) );
  NAND U5748 ( .A(n3925), .B(n3926), .Z(y[71]) );
  NANDN U5749 ( .A(n3863), .B(m[71]), .Z(n3926) );
  NANDN U5750 ( .A(n3864), .B(creg[71]), .Z(n3925) );
  NAND U5751 ( .A(n3927), .B(n3928), .Z(y[70]) );
  NANDN U5752 ( .A(n3863), .B(m[70]), .Z(n3928) );
  NANDN U5753 ( .A(n3864), .B(creg[70]), .Z(n3927) );
  NAND U5754 ( .A(n3929), .B(n3930), .Z(y[6]) );
  NANDN U5755 ( .A(n3863), .B(m[6]), .Z(n3930) );
  NANDN U5756 ( .A(n3864), .B(creg[6]), .Z(n3929) );
  NAND U5757 ( .A(n3931), .B(n3932), .Z(y[69]) );
  NANDN U5758 ( .A(n3863), .B(m[69]), .Z(n3932) );
  NANDN U5759 ( .A(n3864), .B(creg[69]), .Z(n3931) );
  NAND U5760 ( .A(n3933), .B(n3934), .Z(y[68]) );
  NANDN U5761 ( .A(n3863), .B(m[68]), .Z(n3934) );
  NANDN U5762 ( .A(n3864), .B(creg[68]), .Z(n3933) );
  NAND U5763 ( .A(n3935), .B(n3936), .Z(y[67]) );
  NANDN U5764 ( .A(n3863), .B(m[67]), .Z(n3936) );
  NANDN U5765 ( .A(n3864), .B(creg[67]), .Z(n3935) );
  NAND U5766 ( .A(n3937), .B(n3938), .Z(y[66]) );
  NANDN U5767 ( .A(n3863), .B(m[66]), .Z(n3938) );
  NANDN U5768 ( .A(n3864), .B(creg[66]), .Z(n3937) );
  NAND U5769 ( .A(n3939), .B(n3940), .Z(y[65]) );
  NANDN U5770 ( .A(n3863), .B(m[65]), .Z(n3940) );
  NANDN U5771 ( .A(n3864), .B(creg[65]), .Z(n3939) );
  NAND U5772 ( .A(n3941), .B(n3942), .Z(y[64]) );
  NANDN U5773 ( .A(n3863), .B(m[64]), .Z(n3942) );
  NANDN U5774 ( .A(n3864), .B(creg[64]), .Z(n3941) );
  NAND U5775 ( .A(n3943), .B(n3944), .Z(y[63]) );
  NANDN U5776 ( .A(n3863), .B(m[63]), .Z(n3944) );
  NANDN U5777 ( .A(n3864), .B(creg[63]), .Z(n3943) );
  NAND U5778 ( .A(n3945), .B(n3946), .Z(y[62]) );
  NANDN U5779 ( .A(n3863), .B(m[62]), .Z(n3946) );
  NANDN U5780 ( .A(n3864), .B(creg[62]), .Z(n3945) );
  NAND U5781 ( .A(n3947), .B(n3948), .Z(y[61]) );
  NANDN U5782 ( .A(n3863), .B(m[61]), .Z(n3948) );
  NANDN U5783 ( .A(n3864), .B(creg[61]), .Z(n3947) );
  NAND U5784 ( .A(n3949), .B(n3950), .Z(y[60]) );
  NANDN U5785 ( .A(n3863), .B(m[60]), .Z(n3950) );
  NANDN U5786 ( .A(n3864), .B(creg[60]), .Z(n3949) );
  NAND U5787 ( .A(n3951), .B(n3952), .Z(y[5]) );
  NANDN U5788 ( .A(n3863), .B(m[5]), .Z(n3952) );
  NANDN U5789 ( .A(n3864), .B(creg[5]), .Z(n3951) );
  NAND U5790 ( .A(n3953), .B(n3954), .Z(y[59]) );
  NANDN U5791 ( .A(n3863), .B(m[59]), .Z(n3954) );
  NANDN U5792 ( .A(n3864), .B(creg[59]), .Z(n3953) );
  NAND U5793 ( .A(n3955), .B(n3956), .Z(y[58]) );
  NANDN U5794 ( .A(n3863), .B(m[58]), .Z(n3956) );
  NANDN U5795 ( .A(n3864), .B(creg[58]), .Z(n3955) );
  NAND U5796 ( .A(n3957), .B(n3958), .Z(y[57]) );
  NANDN U5797 ( .A(n3863), .B(m[57]), .Z(n3958) );
  NANDN U5798 ( .A(n3864), .B(creg[57]), .Z(n3957) );
  NAND U5799 ( .A(n3959), .B(n3960), .Z(y[56]) );
  NANDN U5800 ( .A(n3863), .B(m[56]), .Z(n3960) );
  NANDN U5801 ( .A(n3864), .B(creg[56]), .Z(n3959) );
  NAND U5802 ( .A(n3961), .B(n3962), .Z(y[55]) );
  NANDN U5803 ( .A(n3863), .B(m[55]), .Z(n3962) );
  NANDN U5804 ( .A(n3864), .B(creg[55]), .Z(n3961) );
  NAND U5805 ( .A(n3963), .B(n3964), .Z(y[54]) );
  NANDN U5806 ( .A(n3863), .B(m[54]), .Z(n3964) );
  NANDN U5807 ( .A(n3864), .B(creg[54]), .Z(n3963) );
  NAND U5808 ( .A(n3965), .B(n3966), .Z(y[53]) );
  NANDN U5809 ( .A(n3863), .B(m[53]), .Z(n3966) );
  NANDN U5810 ( .A(n3864), .B(creg[53]), .Z(n3965) );
  NAND U5811 ( .A(n3967), .B(n3968), .Z(y[52]) );
  NANDN U5812 ( .A(n3863), .B(m[52]), .Z(n3968) );
  NANDN U5813 ( .A(n3864), .B(creg[52]), .Z(n3967) );
  NAND U5814 ( .A(n3969), .B(n3970), .Z(y[51]) );
  NANDN U5815 ( .A(n3863), .B(m[51]), .Z(n3970) );
  NANDN U5816 ( .A(n3864), .B(creg[51]), .Z(n3969) );
  NAND U5817 ( .A(n3971), .B(n3972), .Z(y[50]) );
  NANDN U5818 ( .A(n3863), .B(m[50]), .Z(n3972) );
  NANDN U5819 ( .A(n3864), .B(creg[50]), .Z(n3971) );
  NAND U5820 ( .A(n3973), .B(n3974), .Z(y[4]) );
  NANDN U5821 ( .A(n3863), .B(m[4]), .Z(n3974) );
  NANDN U5822 ( .A(n3864), .B(creg[4]), .Z(n3973) );
  NAND U5823 ( .A(n3975), .B(n3976), .Z(y[49]) );
  NANDN U5824 ( .A(n3863), .B(m[49]), .Z(n3976) );
  NANDN U5825 ( .A(n3864), .B(creg[49]), .Z(n3975) );
  NAND U5826 ( .A(n3977), .B(n3978), .Z(y[48]) );
  NANDN U5827 ( .A(n3863), .B(m[48]), .Z(n3978) );
  NANDN U5828 ( .A(n3864), .B(creg[48]), .Z(n3977) );
  NAND U5829 ( .A(n3979), .B(n3980), .Z(y[47]) );
  NANDN U5830 ( .A(n3863), .B(m[47]), .Z(n3980) );
  NANDN U5831 ( .A(n3864), .B(creg[47]), .Z(n3979) );
  NAND U5832 ( .A(n3981), .B(n3982), .Z(y[46]) );
  NANDN U5833 ( .A(n3863), .B(m[46]), .Z(n3982) );
  NANDN U5834 ( .A(n3864), .B(creg[46]), .Z(n3981) );
  NAND U5835 ( .A(n3983), .B(n3984), .Z(y[45]) );
  NANDN U5836 ( .A(n3863), .B(m[45]), .Z(n3984) );
  NANDN U5837 ( .A(n3864), .B(creg[45]), .Z(n3983) );
  NAND U5838 ( .A(n3985), .B(n3986), .Z(y[44]) );
  NANDN U5839 ( .A(n3863), .B(m[44]), .Z(n3986) );
  NANDN U5840 ( .A(n3864), .B(creg[44]), .Z(n3985) );
  NAND U5841 ( .A(n3987), .B(n3988), .Z(y[43]) );
  NANDN U5842 ( .A(n3863), .B(m[43]), .Z(n3988) );
  NANDN U5843 ( .A(n3864), .B(creg[43]), .Z(n3987) );
  NAND U5844 ( .A(n3989), .B(n3990), .Z(y[42]) );
  NANDN U5845 ( .A(n3863), .B(m[42]), .Z(n3990) );
  NANDN U5846 ( .A(n3864), .B(creg[42]), .Z(n3989) );
  NAND U5847 ( .A(n3991), .B(n3992), .Z(y[41]) );
  NANDN U5848 ( .A(n3863), .B(m[41]), .Z(n3992) );
  NANDN U5849 ( .A(n3864), .B(creg[41]), .Z(n3991) );
  NAND U5850 ( .A(n3993), .B(n3994), .Z(y[40]) );
  NANDN U5851 ( .A(n3863), .B(m[40]), .Z(n3994) );
  NANDN U5852 ( .A(n3864), .B(creg[40]), .Z(n3993) );
  NAND U5853 ( .A(n3995), .B(n3996), .Z(y[3]) );
  NANDN U5854 ( .A(n3863), .B(m[3]), .Z(n3996) );
  NANDN U5855 ( .A(n3864), .B(creg[3]), .Z(n3995) );
  NAND U5856 ( .A(n3997), .B(n3998), .Z(y[39]) );
  NANDN U5857 ( .A(n3863), .B(m[39]), .Z(n3998) );
  NANDN U5858 ( .A(n3864), .B(creg[39]), .Z(n3997) );
  NAND U5859 ( .A(n3999), .B(n4000), .Z(y[38]) );
  NANDN U5860 ( .A(n3863), .B(m[38]), .Z(n4000) );
  NANDN U5861 ( .A(n3864), .B(creg[38]), .Z(n3999) );
  NAND U5862 ( .A(n4001), .B(n4002), .Z(y[37]) );
  NANDN U5863 ( .A(n3863), .B(m[37]), .Z(n4002) );
  NANDN U5864 ( .A(n3864), .B(creg[37]), .Z(n4001) );
  NAND U5865 ( .A(n4003), .B(n4004), .Z(y[36]) );
  NANDN U5866 ( .A(n3863), .B(m[36]), .Z(n4004) );
  NANDN U5867 ( .A(n3864), .B(creg[36]), .Z(n4003) );
  NAND U5868 ( .A(n4005), .B(n4006), .Z(y[35]) );
  NANDN U5869 ( .A(n3863), .B(m[35]), .Z(n4006) );
  NANDN U5870 ( .A(n3864), .B(creg[35]), .Z(n4005) );
  NAND U5871 ( .A(n4007), .B(n4008), .Z(y[34]) );
  NANDN U5872 ( .A(n3863), .B(m[34]), .Z(n4008) );
  NANDN U5873 ( .A(n3864), .B(creg[34]), .Z(n4007) );
  NAND U5874 ( .A(n4009), .B(n4010), .Z(y[33]) );
  NANDN U5875 ( .A(n3863), .B(m[33]), .Z(n4010) );
  NANDN U5876 ( .A(n3864), .B(creg[33]), .Z(n4009) );
  NAND U5877 ( .A(n4011), .B(n4012), .Z(y[32]) );
  NANDN U5878 ( .A(n3863), .B(m[32]), .Z(n4012) );
  NANDN U5879 ( .A(n3864), .B(creg[32]), .Z(n4011) );
  NAND U5880 ( .A(n4013), .B(n4014), .Z(y[31]) );
  NANDN U5881 ( .A(n3863), .B(m[31]), .Z(n4014) );
  NANDN U5882 ( .A(n3864), .B(creg[31]), .Z(n4013) );
  NAND U5883 ( .A(n4015), .B(n4016), .Z(y[30]) );
  NANDN U5884 ( .A(n3863), .B(m[30]), .Z(n4016) );
  NANDN U5885 ( .A(n3864), .B(creg[30]), .Z(n4015) );
  NAND U5886 ( .A(n4017), .B(n4018), .Z(y[2]) );
  NANDN U5887 ( .A(n3863), .B(m[2]), .Z(n4018) );
  NANDN U5888 ( .A(n3864), .B(creg[2]), .Z(n4017) );
  NAND U5889 ( .A(n4019), .B(n4020), .Z(y[29]) );
  NANDN U5890 ( .A(n3863), .B(m[29]), .Z(n4020) );
  NANDN U5891 ( .A(n3864), .B(creg[29]), .Z(n4019) );
  NAND U5892 ( .A(n4021), .B(n4022), .Z(y[28]) );
  NANDN U5893 ( .A(n3863), .B(m[28]), .Z(n4022) );
  NANDN U5894 ( .A(n3864), .B(creg[28]), .Z(n4021) );
  NAND U5895 ( .A(n4023), .B(n4024), .Z(y[27]) );
  NANDN U5896 ( .A(n3863), .B(m[27]), .Z(n4024) );
  NANDN U5897 ( .A(n3864), .B(creg[27]), .Z(n4023) );
  NAND U5898 ( .A(n4025), .B(n4026), .Z(y[26]) );
  NANDN U5899 ( .A(n3863), .B(m[26]), .Z(n4026) );
  NANDN U5900 ( .A(n3864), .B(creg[26]), .Z(n4025) );
  NAND U5901 ( .A(n4027), .B(n4028), .Z(y[25]) );
  NANDN U5902 ( .A(n3863), .B(m[25]), .Z(n4028) );
  NANDN U5903 ( .A(n3864), .B(creg[25]), .Z(n4027) );
  NAND U5904 ( .A(n4029), .B(n4030), .Z(y[255]) );
  NANDN U5905 ( .A(n3863), .B(m[255]), .Z(n4030) );
  NANDN U5906 ( .A(n3864), .B(creg[255]), .Z(n4029) );
  NAND U5907 ( .A(n4031), .B(n4032), .Z(y[254]) );
  NANDN U5908 ( .A(n3863), .B(m[254]), .Z(n4032) );
  NANDN U5909 ( .A(n3864), .B(creg[254]), .Z(n4031) );
  NAND U5910 ( .A(n4033), .B(n4034), .Z(y[253]) );
  NANDN U5911 ( .A(n3863), .B(m[253]), .Z(n4034) );
  NANDN U5912 ( .A(n3864), .B(creg[253]), .Z(n4033) );
  NAND U5913 ( .A(n4035), .B(n4036), .Z(y[252]) );
  NANDN U5914 ( .A(n3863), .B(m[252]), .Z(n4036) );
  NANDN U5915 ( .A(n3864), .B(creg[252]), .Z(n4035) );
  NAND U5916 ( .A(n4037), .B(n4038), .Z(y[251]) );
  NANDN U5917 ( .A(n3863), .B(m[251]), .Z(n4038) );
  NANDN U5918 ( .A(n3864), .B(creg[251]), .Z(n4037) );
  NAND U5919 ( .A(n4039), .B(n4040), .Z(y[250]) );
  NANDN U5920 ( .A(n3863), .B(m[250]), .Z(n4040) );
  NANDN U5921 ( .A(n3864), .B(creg[250]), .Z(n4039) );
  NAND U5922 ( .A(n4041), .B(n4042), .Z(y[24]) );
  NANDN U5923 ( .A(n3863), .B(m[24]), .Z(n4042) );
  NANDN U5924 ( .A(n3864), .B(creg[24]), .Z(n4041) );
  NAND U5925 ( .A(n4043), .B(n4044), .Z(y[249]) );
  NANDN U5926 ( .A(n3863), .B(m[249]), .Z(n4044) );
  NANDN U5927 ( .A(n3864), .B(creg[249]), .Z(n4043) );
  NAND U5928 ( .A(n4045), .B(n4046), .Z(y[248]) );
  NANDN U5929 ( .A(n3863), .B(m[248]), .Z(n4046) );
  NANDN U5930 ( .A(n3864), .B(creg[248]), .Z(n4045) );
  NAND U5931 ( .A(n4047), .B(n4048), .Z(y[247]) );
  NANDN U5932 ( .A(n3863), .B(m[247]), .Z(n4048) );
  NANDN U5933 ( .A(n3864), .B(creg[247]), .Z(n4047) );
  NAND U5934 ( .A(n4049), .B(n4050), .Z(y[246]) );
  NANDN U5935 ( .A(n3863), .B(m[246]), .Z(n4050) );
  NANDN U5936 ( .A(n3864), .B(creg[246]), .Z(n4049) );
  NAND U5937 ( .A(n4051), .B(n4052), .Z(y[245]) );
  NANDN U5938 ( .A(n3863), .B(m[245]), .Z(n4052) );
  NANDN U5939 ( .A(n3864), .B(creg[245]), .Z(n4051) );
  NAND U5940 ( .A(n4053), .B(n4054), .Z(y[244]) );
  NANDN U5941 ( .A(n3863), .B(m[244]), .Z(n4054) );
  NANDN U5942 ( .A(n3864), .B(creg[244]), .Z(n4053) );
  NAND U5943 ( .A(n4055), .B(n4056), .Z(y[243]) );
  NANDN U5944 ( .A(n3863), .B(m[243]), .Z(n4056) );
  NANDN U5945 ( .A(n3864), .B(creg[243]), .Z(n4055) );
  NAND U5946 ( .A(n4057), .B(n4058), .Z(y[242]) );
  NANDN U5947 ( .A(n3863), .B(m[242]), .Z(n4058) );
  NANDN U5948 ( .A(n3864), .B(creg[242]), .Z(n4057) );
  NAND U5949 ( .A(n4059), .B(n4060), .Z(y[241]) );
  NANDN U5950 ( .A(n3863), .B(m[241]), .Z(n4060) );
  NANDN U5951 ( .A(n3864), .B(creg[241]), .Z(n4059) );
  NAND U5952 ( .A(n4061), .B(n4062), .Z(y[240]) );
  NANDN U5953 ( .A(n3863), .B(m[240]), .Z(n4062) );
  NANDN U5954 ( .A(n3864), .B(creg[240]), .Z(n4061) );
  NAND U5955 ( .A(n4063), .B(n4064), .Z(y[23]) );
  NANDN U5956 ( .A(n3863), .B(m[23]), .Z(n4064) );
  NANDN U5957 ( .A(n3864), .B(creg[23]), .Z(n4063) );
  NAND U5958 ( .A(n4065), .B(n4066), .Z(y[239]) );
  NANDN U5959 ( .A(n3863), .B(m[239]), .Z(n4066) );
  NANDN U5960 ( .A(n3864), .B(creg[239]), .Z(n4065) );
  NAND U5961 ( .A(n4067), .B(n4068), .Z(y[238]) );
  NANDN U5962 ( .A(n3863), .B(m[238]), .Z(n4068) );
  NANDN U5963 ( .A(n3864), .B(creg[238]), .Z(n4067) );
  NAND U5964 ( .A(n4069), .B(n4070), .Z(y[237]) );
  NANDN U5965 ( .A(n3863), .B(m[237]), .Z(n4070) );
  NANDN U5966 ( .A(n3864), .B(creg[237]), .Z(n4069) );
  NAND U5967 ( .A(n4071), .B(n4072), .Z(y[236]) );
  NANDN U5968 ( .A(n3863), .B(m[236]), .Z(n4072) );
  NANDN U5969 ( .A(n3864), .B(creg[236]), .Z(n4071) );
  NAND U5970 ( .A(n4073), .B(n4074), .Z(y[235]) );
  NANDN U5971 ( .A(n3863), .B(m[235]), .Z(n4074) );
  NANDN U5972 ( .A(n3864), .B(creg[235]), .Z(n4073) );
  NAND U5973 ( .A(n4075), .B(n4076), .Z(y[234]) );
  NANDN U5974 ( .A(n3863), .B(m[234]), .Z(n4076) );
  NANDN U5975 ( .A(n3864), .B(creg[234]), .Z(n4075) );
  NAND U5976 ( .A(n4077), .B(n4078), .Z(y[233]) );
  NANDN U5977 ( .A(n3863), .B(m[233]), .Z(n4078) );
  NANDN U5978 ( .A(n3864), .B(creg[233]), .Z(n4077) );
  NAND U5979 ( .A(n4079), .B(n4080), .Z(y[232]) );
  NANDN U5980 ( .A(n3863), .B(m[232]), .Z(n4080) );
  NANDN U5981 ( .A(n3864), .B(creg[232]), .Z(n4079) );
  NAND U5982 ( .A(n4081), .B(n4082), .Z(y[231]) );
  NANDN U5983 ( .A(n3863), .B(m[231]), .Z(n4082) );
  NANDN U5984 ( .A(n3864), .B(creg[231]), .Z(n4081) );
  NAND U5985 ( .A(n4083), .B(n4084), .Z(y[230]) );
  NANDN U5986 ( .A(n3863), .B(m[230]), .Z(n4084) );
  NANDN U5987 ( .A(n3864), .B(creg[230]), .Z(n4083) );
  NAND U5988 ( .A(n4085), .B(n4086), .Z(y[22]) );
  NANDN U5989 ( .A(n3863), .B(m[22]), .Z(n4086) );
  NANDN U5990 ( .A(n3864), .B(creg[22]), .Z(n4085) );
  NAND U5991 ( .A(n4087), .B(n4088), .Z(y[229]) );
  NANDN U5992 ( .A(n3863), .B(m[229]), .Z(n4088) );
  NANDN U5993 ( .A(n3864), .B(creg[229]), .Z(n4087) );
  NAND U5994 ( .A(n4089), .B(n4090), .Z(y[228]) );
  NANDN U5995 ( .A(n3863), .B(m[228]), .Z(n4090) );
  NANDN U5996 ( .A(n3864), .B(creg[228]), .Z(n4089) );
  NAND U5997 ( .A(n4091), .B(n4092), .Z(y[227]) );
  NANDN U5998 ( .A(n3863), .B(m[227]), .Z(n4092) );
  NANDN U5999 ( .A(n3864), .B(creg[227]), .Z(n4091) );
  NAND U6000 ( .A(n4093), .B(n4094), .Z(y[226]) );
  NANDN U6001 ( .A(n3863), .B(m[226]), .Z(n4094) );
  NANDN U6002 ( .A(n3864), .B(creg[226]), .Z(n4093) );
  NAND U6003 ( .A(n4095), .B(n4096), .Z(y[225]) );
  NANDN U6004 ( .A(n3863), .B(m[225]), .Z(n4096) );
  NANDN U6005 ( .A(n3864), .B(creg[225]), .Z(n4095) );
  NAND U6006 ( .A(n4097), .B(n4098), .Z(y[224]) );
  NANDN U6007 ( .A(n3863), .B(m[224]), .Z(n4098) );
  NANDN U6008 ( .A(n3864), .B(creg[224]), .Z(n4097) );
  NAND U6009 ( .A(n4099), .B(n4100), .Z(y[223]) );
  NANDN U6010 ( .A(n3863), .B(m[223]), .Z(n4100) );
  NANDN U6011 ( .A(n3864), .B(creg[223]), .Z(n4099) );
  NAND U6012 ( .A(n4101), .B(n4102), .Z(y[222]) );
  NANDN U6013 ( .A(n3863), .B(m[222]), .Z(n4102) );
  NANDN U6014 ( .A(n3864), .B(creg[222]), .Z(n4101) );
  NAND U6015 ( .A(n4103), .B(n4104), .Z(y[221]) );
  NANDN U6016 ( .A(n3863), .B(m[221]), .Z(n4104) );
  NANDN U6017 ( .A(n3864), .B(creg[221]), .Z(n4103) );
  NAND U6018 ( .A(n4105), .B(n4106), .Z(y[220]) );
  NANDN U6019 ( .A(n3863), .B(m[220]), .Z(n4106) );
  NANDN U6020 ( .A(n3864), .B(creg[220]), .Z(n4105) );
  NAND U6021 ( .A(n4107), .B(n4108), .Z(y[21]) );
  NANDN U6022 ( .A(n3863), .B(m[21]), .Z(n4108) );
  NANDN U6023 ( .A(n3864), .B(creg[21]), .Z(n4107) );
  NAND U6024 ( .A(n4109), .B(n4110), .Z(y[219]) );
  NANDN U6025 ( .A(n3863), .B(m[219]), .Z(n4110) );
  NANDN U6026 ( .A(n3864), .B(creg[219]), .Z(n4109) );
  NAND U6027 ( .A(n4111), .B(n4112), .Z(y[218]) );
  NANDN U6028 ( .A(n3863), .B(m[218]), .Z(n4112) );
  NANDN U6029 ( .A(n3864), .B(creg[218]), .Z(n4111) );
  NAND U6030 ( .A(n4113), .B(n4114), .Z(y[217]) );
  NANDN U6031 ( .A(n3863), .B(m[217]), .Z(n4114) );
  NANDN U6032 ( .A(n3864), .B(creg[217]), .Z(n4113) );
  NAND U6033 ( .A(n4115), .B(n4116), .Z(y[216]) );
  NANDN U6034 ( .A(n3863), .B(m[216]), .Z(n4116) );
  NANDN U6035 ( .A(n3864), .B(creg[216]), .Z(n4115) );
  NAND U6036 ( .A(n4117), .B(n4118), .Z(y[215]) );
  NANDN U6037 ( .A(n3863), .B(m[215]), .Z(n4118) );
  NANDN U6038 ( .A(n3864), .B(creg[215]), .Z(n4117) );
  NAND U6039 ( .A(n4119), .B(n4120), .Z(y[214]) );
  NANDN U6040 ( .A(n3863), .B(m[214]), .Z(n4120) );
  NANDN U6041 ( .A(n3864), .B(creg[214]), .Z(n4119) );
  NAND U6042 ( .A(n4121), .B(n4122), .Z(y[213]) );
  NANDN U6043 ( .A(n3863), .B(m[213]), .Z(n4122) );
  NANDN U6044 ( .A(n3864), .B(creg[213]), .Z(n4121) );
  NAND U6045 ( .A(n4123), .B(n4124), .Z(y[212]) );
  NANDN U6046 ( .A(n3863), .B(m[212]), .Z(n4124) );
  NANDN U6047 ( .A(n3864), .B(creg[212]), .Z(n4123) );
  NAND U6048 ( .A(n4125), .B(n4126), .Z(y[211]) );
  NANDN U6049 ( .A(n3863), .B(m[211]), .Z(n4126) );
  NANDN U6050 ( .A(n3864), .B(creg[211]), .Z(n4125) );
  NAND U6051 ( .A(n4127), .B(n4128), .Z(y[210]) );
  NANDN U6052 ( .A(n3863), .B(m[210]), .Z(n4128) );
  NANDN U6053 ( .A(n3864), .B(creg[210]), .Z(n4127) );
  NAND U6054 ( .A(n4129), .B(n4130), .Z(y[20]) );
  NANDN U6055 ( .A(n3863), .B(m[20]), .Z(n4130) );
  NANDN U6056 ( .A(n3864), .B(creg[20]), .Z(n4129) );
  NAND U6057 ( .A(n4131), .B(n4132), .Z(y[209]) );
  NANDN U6058 ( .A(n3863), .B(m[209]), .Z(n4132) );
  NANDN U6059 ( .A(n3864), .B(creg[209]), .Z(n4131) );
  NAND U6060 ( .A(n4133), .B(n4134), .Z(y[208]) );
  NANDN U6061 ( .A(n3863), .B(m[208]), .Z(n4134) );
  NANDN U6062 ( .A(n3864), .B(creg[208]), .Z(n4133) );
  NAND U6063 ( .A(n4135), .B(n4136), .Z(y[207]) );
  NANDN U6064 ( .A(n3863), .B(m[207]), .Z(n4136) );
  NANDN U6065 ( .A(n3864), .B(creg[207]), .Z(n4135) );
  NAND U6066 ( .A(n4137), .B(n4138), .Z(y[206]) );
  NANDN U6067 ( .A(n3863), .B(m[206]), .Z(n4138) );
  NANDN U6068 ( .A(n3864), .B(creg[206]), .Z(n4137) );
  NAND U6069 ( .A(n4139), .B(n4140), .Z(y[205]) );
  NANDN U6070 ( .A(n3863), .B(m[205]), .Z(n4140) );
  NANDN U6071 ( .A(n3864), .B(creg[205]), .Z(n4139) );
  NAND U6072 ( .A(n4141), .B(n4142), .Z(y[204]) );
  NANDN U6073 ( .A(n3863), .B(m[204]), .Z(n4142) );
  NANDN U6074 ( .A(n3864), .B(creg[204]), .Z(n4141) );
  NAND U6075 ( .A(n4143), .B(n4144), .Z(y[203]) );
  NANDN U6076 ( .A(n3863), .B(m[203]), .Z(n4144) );
  NANDN U6077 ( .A(n3864), .B(creg[203]), .Z(n4143) );
  NAND U6078 ( .A(n4145), .B(n4146), .Z(y[202]) );
  NANDN U6079 ( .A(n3863), .B(m[202]), .Z(n4146) );
  NANDN U6080 ( .A(n3864), .B(creg[202]), .Z(n4145) );
  NAND U6081 ( .A(n4147), .B(n4148), .Z(y[201]) );
  NANDN U6082 ( .A(n3863), .B(m[201]), .Z(n4148) );
  NANDN U6083 ( .A(n3864), .B(creg[201]), .Z(n4147) );
  NAND U6084 ( .A(n4149), .B(n4150), .Z(y[200]) );
  NANDN U6085 ( .A(n3863), .B(m[200]), .Z(n4150) );
  NANDN U6086 ( .A(n3864), .B(creg[200]), .Z(n4149) );
  NAND U6087 ( .A(n4151), .B(n4152), .Z(y[1]) );
  NANDN U6088 ( .A(n3863), .B(m[1]), .Z(n4152) );
  NANDN U6089 ( .A(n3864), .B(creg[1]), .Z(n4151) );
  NAND U6090 ( .A(n4153), .B(n4154), .Z(y[19]) );
  NANDN U6091 ( .A(n3863), .B(m[19]), .Z(n4154) );
  NANDN U6092 ( .A(n3864), .B(creg[19]), .Z(n4153) );
  NAND U6093 ( .A(n4155), .B(n4156), .Z(y[199]) );
  NANDN U6094 ( .A(n3863), .B(m[199]), .Z(n4156) );
  NANDN U6095 ( .A(n3864), .B(creg[199]), .Z(n4155) );
  NAND U6096 ( .A(n4157), .B(n4158), .Z(y[198]) );
  NANDN U6097 ( .A(n3863), .B(m[198]), .Z(n4158) );
  NANDN U6098 ( .A(n3864), .B(creg[198]), .Z(n4157) );
  NAND U6099 ( .A(n4159), .B(n4160), .Z(y[197]) );
  NANDN U6100 ( .A(n3863), .B(m[197]), .Z(n4160) );
  NANDN U6101 ( .A(n3864), .B(creg[197]), .Z(n4159) );
  NAND U6102 ( .A(n4161), .B(n4162), .Z(y[196]) );
  NANDN U6103 ( .A(n3863), .B(m[196]), .Z(n4162) );
  NANDN U6104 ( .A(n3864), .B(creg[196]), .Z(n4161) );
  NAND U6105 ( .A(n4163), .B(n4164), .Z(y[195]) );
  NANDN U6106 ( .A(n3863), .B(m[195]), .Z(n4164) );
  NANDN U6107 ( .A(n3864), .B(creg[195]), .Z(n4163) );
  NAND U6108 ( .A(n4165), .B(n4166), .Z(y[194]) );
  NANDN U6109 ( .A(n3863), .B(m[194]), .Z(n4166) );
  NANDN U6110 ( .A(n3864), .B(creg[194]), .Z(n4165) );
  NAND U6111 ( .A(n4167), .B(n4168), .Z(y[193]) );
  NANDN U6112 ( .A(n3863), .B(m[193]), .Z(n4168) );
  NANDN U6113 ( .A(n3864), .B(creg[193]), .Z(n4167) );
  NAND U6114 ( .A(n4169), .B(n4170), .Z(y[192]) );
  NANDN U6115 ( .A(n3863), .B(m[192]), .Z(n4170) );
  NANDN U6116 ( .A(n3864), .B(creg[192]), .Z(n4169) );
  NAND U6117 ( .A(n4171), .B(n4172), .Z(y[191]) );
  NANDN U6118 ( .A(n3863), .B(m[191]), .Z(n4172) );
  NANDN U6119 ( .A(n3864), .B(creg[191]), .Z(n4171) );
  NAND U6120 ( .A(n4173), .B(n4174), .Z(y[190]) );
  NANDN U6121 ( .A(n3863), .B(m[190]), .Z(n4174) );
  NANDN U6122 ( .A(n3864), .B(creg[190]), .Z(n4173) );
  NAND U6123 ( .A(n4175), .B(n4176), .Z(y[18]) );
  NANDN U6124 ( .A(n3863), .B(m[18]), .Z(n4176) );
  NANDN U6125 ( .A(n3864), .B(creg[18]), .Z(n4175) );
  NAND U6126 ( .A(n4177), .B(n4178), .Z(y[189]) );
  NANDN U6127 ( .A(n3863), .B(m[189]), .Z(n4178) );
  NANDN U6128 ( .A(n3864), .B(creg[189]), .Z(n4177) );
  NAND U6129 ( .A(n4179), .B(n4180), .Z(y[188]) );
  NANDN U6130 ( .A(n3863), .B(m[188]), .Z(n4180) );
  NANDN U6131 ( .A(n3864), .B(creg[188]), .Z(n4179) );
  NAND U6132 ( .A(n4181), .B(n4182), .Z(y[187]) );
  NANDN U6133 ( .A(n3863), .B(m[187]), .Z(n4182) );
  NANDN U6134 ( .A(n3864), .B(creg[187]), .Z(n4181) );
  NAND U6135 ( .A(n4183), .B(n4184), .Z(y[186]) );
  NANDN U6136 ( .A(n3863), .B(m[186]), .Z(n4184) );
  NANDN U6137 ( .A(n3864), .B(creg[186]), .Z(n4183) );
  NAND U6138 ( .A(n4185), .B(n4186), .Z(y[185]) );
  NANDN U6139 ( .A(n3863), .B(m[185]), .Z(n4186) );
  NANDN U6140 ( .A(n3864), .B(creg[185]), .Z(n4185) );
  NAND U6141 ( .A(n4187), .B(n4188), .Z(y[184]) );
  NANDN U6142 ( .A(n3863), .B(m[184]), .Z(n4188) );
  NANDN U6143 ( .A(n3864), .B(creg[184]), .Z(n4187) );
  NAND U6144 ( .A(n4189), .B(n4190), .Z(y[183]) );
  NANDN U6145 ( .A(n3863), .B(m[183]), .Z(n4190) );
  NANDN U6146 ( .A(n3864), .B(creg[183]), .Z(n4189) );
  NAND U6147 ( .A(n4191), .B(n4192), .Z(y[182]) );
  NANDN U6148 ( .A(n3863), .B(m[182]), .Z(n4192) );
  NANDN U6149 ( .A(n3864), .B(creg[182]), .Z(n4191) );
  NAND U6150 ( .A(n4193), .B(n4194), .Z(y[181]) );
  NANDN U6151 ( .A(n3863), .B(m[181]), .Z(n4194) );
  NANDN U6152 ( .A(n3864), .B(creg[181]), .Z(n4193) );
  NAND U6153 ( .A(n4195), .B(n4196), .Z(y[180]) );
  NANDN U6154 ( .A(n3863), .B(m[180]), .Z(n4196) );
  NANDN U6155 ( .A(n3864), .B(creg[180]), .Z(n4195) );
  NAND U6156 ( .A(n4197), .B(n4198), .Z(y[17]) );
  NANDN U6157 ( .A(n3863), .B(m[17]), .Z(n4198) );
  NANDN U6158 ( .A(n3864), .B(creg[17]), .Z(n4197) );
  NAND U6159 ( .A(n4199), .B(n4200), .Z(y[179]) );
  NANDN U6160 ( .A(n3863), .B(m[179]), .Z(n4200) );
  NANDN U6161 ( .A(n3864), .B(creg[179]), .Z(n4199) );
  NAND U6162 ( .A(n4201), .B(n4202), .Z(y[178]) );
  NANDN U6163 ( .A(n3863), .B(m[178]), .Z(n4202) );
  NANDN U6164 ( .A(n3864), .B(creg[178]), .Z(n4201) );
  NAND U6165 ( .A(n4203), .B(n4204), .Z(y[177]) );
  NANDN U6166 ( .A(n3863), .B(m[177]), .Z(n4204) );
  NANDN U6167 ( .A(n3864), .B(creg[177]), .Z(n4203) );
  NAND U6168 ( .A(n4205), .B(n4206), .Z(y[176]) );
  NANDN U6169 ( .A(n3863), .B(m[176]), .Z(n4206) );
  NANDN U6170 ( .A(n3864), .B(creg[176]), .Z(n4205) );
  NAND U6171 ( .A(n4207), .B(n4208), .Z(y[175]) );
  NANDN U6172 ( .A(n3863), .B(m[175]), .Z(n4208) );
  NANDN U6173 ( .A(n3864), .B(creg[175]), .Z(n4207) );
  NAND U6174 ( .A(n4209), .B(n4210), .Z(y[174]) );
  NANDN U6175 ( .A(n3863), .B(m[174]), .Z(n4210) );
  NANDN U6176 ( .A(n3864), .B(creg[174]), .Z(n4209) );
  NAND U6177 ( .A(n4211), .B(n4212), .Z(y[173]) );
  NANDN U6178 ( .A(n3863), .B(m[173]), .Z(n4212) );
  NANDN U6179 ( .A(n3864), .B(creg[173]), .Z(n4211) );
  NAND U6180 ( .A(n4213), .B(n4214), .Z(y[172]) );
  NANDN U6181 ( .A(n3863), .B(m[172]), .Z(n4214) );
  NANDN U6182 ( .A(n3864), .B(creg[172]), .Z(n4213) );
  NAND U6183 ( .A(n4215), .B(n4216), .Z(y[171]) );
  NANDN U6184 ( .A(n3863), .B(m[171]), .Z(n4216) );
  NANDN U6185 ( .A(n3864), .B(creg[171]), .Z(n4215) );
  NAND U6186 ( .A(n4217), .B(n4218), .Z(y[170]) );
  NANDN U6187 ( .A(n3863), .B(m[170]), .Z(n4218) );
  NANDN U6188 ( .A(n3864), .B(creg[170]), .Z(n4217) );
  NAND U6189 ( .A(n4219), .B(n4220), .Z(y[16]) );
  NANDN U6190 ( .A(n3863), .B(m[16]), .Z(n4220) );
  NANDN U6191 ( .A(n3864), .B(creg[16]), .Z(n4219) );
  NAND U6192 ( .A(n4221), .B(n4222), .Z(y[169]) );
  NANDN U6193 ( .A(n3863), .B(m[169]), .Z(n4222) );
  NANDN U6194 ( .A(n3864), .B(creg[169]), .Z(n4221) );
  NAND U6195 ( .A(n4223), .B(n4224), .Z(y[168]) );
  NANDN U6196 ( .A(n3863), .B(m[168]), .Z(n4224) );
  NANDN U6197 ( .A(n3864), .B(creg[168]), .Z(n4223) );
  NAND U6198 ( .A(n4225), .B(n4226), .Z(y[167]) );
  NANDN U6199 ( .A(n3863), .B(m[167]), .Z(n4226) );
  NANDN U6200 ( .A(n3864), .B(creg[167]), .Z(n4225) );
  NAND U6201 ( .A(n4227), .B(n4228), .Z(y[166]) );
  NANDN U6202 ( .A(n3863), .B(m[166]), .Z(n4228) );
  NANDN U6203 ( .A(n3864), .B(creg[166]), .Z(n4227) );
  NAND U6204 ( .A(n4229), .B(n4230), .Z(y[165]) );
  NANDN U6205 ( .A(n3863), .B(m[165]), .Z(n4230) );
  NANDN U6206 ( .A(n3864), .B(creg[165]), .Z(n4229) );
  NAND U6207 ( .A(n4231), .B(n4232), .Z(y[164]) );
  NANDN U6208 ( .A(n3863), .B(m[164]), .Z(n4232) );
  NANDN U6209 ( .A(n3864), .B(creg[164]), .Z(n4231) );
  NAND U6210 ( .A(n4233), .B(n4234), .Z(y[163]) );
  NANDN U6211 ( .A(n3863), .B(m[163]), .Z(n4234) );
  NANDN U6212 ( .A(n3864), .B(creg[163]), .Z(n4233) );
  NAND U6213 ( .A(n4235), .B(n4236), .Z(y[162]) );
  NANDN U6214 ( .A(n3863), .B(m[162]), .Z(n4236) );
  NANDN U6215 ( .A(n3864), .B(creg[162]), .Z(n4235) );
  NAND U6216 ( .A(n4237), .B(n4238), .Z(y[161]) );
  NANDN U6217 ( .A(n3863), .B(m[161]), .Z(n4238) );
  NANDN U6218 ( .A(n3864), .B(creg[161]), .Z(n4237) );
  NAND U6219 ( .A(n4239), .B(n4240), .Z(y[160]) );
  NANDN U6220 ( .A(n3863), .B(m[160]), .Z(n4240) );
  NANDN U6221 ( .A(n3864), .B(creg[160]), .Z(n4239) );
  NAND U6222 ( .A(n4241), .B(n4242), .Z(y[15]) );
  NANDN U6223 ( .A(n3863), .B(m[15]), .Z(n4242) );
  NANDN U6224 ( .A(n3864), .B(creg[15]), .Z(n4241) );
  NAND U6225 ( .A(n4243), .B(n4244), .Z(y[159]) );
  NANDN U6226 ( .A(n3863), .B(m[159]), .Z(n4244) );
  NANDN U6227 ( .A(n3864), .B(creg[159]), .Z(n4243) );
  NAND U6228 ( .A(n4245), .B(n4246), .Z(y[158]) );
  NANDN U6229 ( .A(n3863), .B(m[158]), .Z(n4246) );
  NANDN U6230 ( .A(n3864), .B(creg[158]), .Z(n4245) );
  NAND U6231 ( .A(n4247), .B(n4248), .Z(y[157]) );
  NANDN U6232 ( .A(n3863), .B(m[157]), .Z(n4248) );
  NANDN U6233 ( .A(n3864), .B(creg[157]), .Z(n4247) );
  NAND U6234 ( .A(n4249), .B(n4250), .Z(y[156]) );
  NANDN U6235 ( .A(n3863), .B(m[156]), .Z(n4250) );
  NANDN U6236 ( .A(n3864), .B(creg[156]), .Z(n4249) );
  NAND U6237 ( .A(n4251), .B(n4252), .Z(y[155]) );
  NANDN U6238 ( .A(n3863), .B(m[155]), .Z(n4252) );
  NANDN U6239 ( .A(n3864), .B(creg[155]), .Z(n4251) );
  NAND U6240 ( .A(n4253), .B(n4254), .Z(y[154]) );
  NANDN U6241 ( .A(n3863), .B(m[154]), .Z(n4254) );
  NANDN U6242 ( .A(n3864), .B(creg[154]), .Z(n4253) );
  NAND U6243 ( .A(n4255), .B(n4256), .Z(y[153]) );
  NANDN U6244 ( .A(n3863), .B(m[153]), .Z(n4256) );
  NANDN U6245 ( .A(n3864), .B(creg[153]), .Z(n4255) );
  NAND U6246 ( .A(n4257), .B(n4258), .Z(y[152]) );
  NANDN U6247 ( .A(n3863), .B(m[152]), .Z(n4258) );
  NANDN U6248 ( .A(n3864), .B(creg[152]), .Z(n4257) );
  NAND U6249 ( .A(n4259), .B(n4260), .Z(y[151]) );
  NANDN U6250 ( .A(n3863), .B(m[151]), .Z(n4260) );
  NANDN U6251 ( .A(n3864), .B(creg[151]), .Z(n4259) );
  NAND U6252 ( .A(n4261), .B(n4262), .Z(y[150]) );
  NANDN U6253 ( .A(n3863), .B(m[150]), .Z(n4262) );
  NANDN U6254 ( .A(n3864), .B(creg[150]), .Z(n4261) );
  NAND U6255 ( .A(n4263), .B(n4264), .Z(y[14]) );
  NANDN U6256 ( .A(n3863), .B(m[14]), .Z(n4264) );
  NANDN U6257 ( .A(n3864), .B(creg[14]), .Z(n4263) );
  NAND U6258 ( .A(n4265), .B(n4266), .Z(y[149]) );
  NANDN U6259 ( .A(n3863), .B(m[149]), .Z(n4266) );
  NANDN U6260 ( .A(n3864), .B(creg[149]), .Z(n4265) );
  NAND U6261 ( .A(n4267), .B(n4268), .Z(y[148]) );
  NANDN U6262 ( .A(n3863), .B(m[148]), .Z(n4268) );
  NANDN U6263 ( .A(n3864), .B(creg[148]), .Z(n4267) );
  NAND U6264 ( .A(n4269), .B(n4270), .Z(y[147]) );
  NANDN U6265 ( .A(n3863), .B(m[147]), .Z(n4270) );
  NANDN U6266 ( .A(n3864), .B(creg[147]), .Z(n4269) );
  NAND U6267 ( .A(n4271), .B(n4272), .Z(y[146]) );
  NANDN U6268 ( .A(n3863), .B(m[146]), .Z(n4272) );
  NANDN U6269 ( .A(n3864), .B(creg[146]), .Z(n4271) );
  NAND U6270 ( .A(n4273), .B(n4274), .Z(y[145]) );
  NANDN U6271 ( .A(n3863), .B(m[145]), .Z(n4274) );
  NANDN U6272 ( .A(n3864), .B(creg[145]), .Z(n4273) );
  NAND U6273 ( .A(n4275), .B(n4276), .Z(y[144]) );
  NANDN U6274 ( .A(n3863), .B(m[144]), .Z(n4276) );
  NANDN U6275 ( .A(n3864), .B(creg[144]), .Z(n4275) );
  NAND U6276 ( .A(n4277), .B(n4278), .Z(y[143]) );
  NANDN U6277 ( .A(n3863), .B(m[143]), .Z(n4278) );
  NANDN U6278 ( .A(n3864), .B(creg[143]), .Z(n4277) );
  NAND U6279 ( .A(n4279), .B(n4280), .Z(y[142]) );
  NANDN U6280 ( .A(n3863), .B(m[142]), .Z(n4280) );
  NANDN U6281 ( .A(n3864), .B(creg[142]), .Z(n4279) );
  NAND U6282 ( .A(n4281), .B(n4282), .Z(y[141]) );
  NANDN U6283 ( .A(n3863), .B(m[141]), .Z(n4282) );
  NANDN U6284 ( .A(n3864), .B(creg[141]), .Z(n4281) );
  NAND U6285 ( .A(n4283), .B(n4284), .Z(y[140]) );
  NANDN U6286 ( .A(n3863), .B(m[140]), .Z(n4284) );
  NANDN U6287 ( .A(n3864), .B(creg[140]), .Z(n4283) );
  NAND U6288 ( .A(n4285), .B(n4286), .Z(y[13]) );
  NANDN U6289 ( .A(n3863), .B(m[13]), .Z(n4286) );
  NANDN U6290 ( .A(n3864), .B(creg[13]), .Z(n4285) );
  NAND U6291 ( .A(n4287), .B(n4288), .Z(y[139]) );
  NANDN U6292 ( .A(n3863), .B(m[139]), .Z(n4288) );
  NANDN U6293 ( .A(n3864), .B(creg[139]), .Z(n4287) );
  NAND U6294 ( .A(n4289), .B(n4290), .Z(y[138]) );
  NANDN U6295 ( .A(n3863), .B(m[138]), .Z(n4290) );
  NANDN U6296 ( .A(n3864), .B(creg[138]), .Z(n4289) );
  NAND U6297 ( .A(n4291), .B(n4292), .Z(y[137]) );
  NANDN U6298 ( .A(n3863), .B(m[137]), .Z(n4292) );
  NANDN U6299 ( .A(n3864), .B(creg[137]), .Z(n4291) );
  NAND U6300 ( .A(n4293), .B(n4294), .Z(y[136]) );
  NANDN U6301 ( .A(n3863), .B(m[136]), .Z(n4294) );
  NANDN U6302 ( .A(n3864), .B(creg[136]), .Z(n4293) );
  NAND U6303 ( .A(n4295), .B(n4296), .Z(y[135]) );
  NANDN U6304 ( .A(n3863), .B(m[135]), .Z(n4296) );
  NANDN U6305 ( .A(n3864), .B(creg[135]), .Z(n4295) );
  NAND U6306 ( .A(n4297), .B(n4298), .Z(y[134]) );
  NANDN U6307 ( .A(n3863), .B(m[134]), .Z(n4298) );
  NANDN U6308 ( .A(n3864), .B(creg[134]), .Z(n4297) );
  NAND U6309 ( .A(n4299), .B(n4300), .Z(y[133]) );
  NANDN U6310 ( .A(n3863), .B(m[133]), .Z(n4300) );
  NANDN U6311 ( .A(n3864), .B(creg[133]), .Z(n4299) );
  NAND U6312 ( .A(n4301), .B(n4302), .Z(y[132]) );
  NANDN U6313 ( .A(n3863), .B(m[132]), .Z(n4302) );
  NANDN U6314 ( .A(n3864), .B(creg[132]), .Z(n4301) );
  NAND U6315 ( .A(n4303), .B(n4304), .Z(y[131]) );
  NANDN U6316 ( .A(n3863), .B(m[131]), .Z(n4304) );
  NANDN U6317 ( .A(n3864), .B(creg[131]), .Z(n4303) );
  NAND U6318 ( .A(n4305), .B(n4306), .Z(y[130]) );
  NANDN U6319 ( .A(n3863), .B(m[130]), .Z(n4306) );
  NANDN U6320 ( .A(n3864), .B(creg[130]), .Z(n4305) );
  NAND U6321 ( .A(n4307), .B(n4308), .Z(y[12]) );
  NANDN U6322 ( .A(n3863), .B(m[12]), .Z(n4308) );
  NANDN U6323 ( .A(n3864), .B(creg[12]), .Z(n4307) );
  NAND U6324 ( .A(n4309), .B(n4310), .Z(y[129]) );
  NANDN U6325 ( .A(n3863), .B(m[129]), .Z(n4310) );
  NANDN U6326 ( .A(n3864), .B(creg[129]), .Z(n4309) );
  NAND U6327 ( .A(n4311), .B(n4312), .Z(y[128]) );
  NANDN U6328 ( .A(n3863), .B(m[128]), .Z(n4312) );
  NANDN U6329 ( .A(n3864), .B(creg[128]), .Z(n4311) );
  NAND U6330 ( .A(n4313), .B(n4314), .Z(y[127]) );
  NANDN U6331 ( .A(n3863), .B(m[127]), .Z(n4314) );
  NANDN U6332 ( .A(n3864), .B(creg[127]), .Z(n4313) );
  NAND U6333 ( .A(n4315), .B(n4316), .Z(y[126]) );
  NANDN U6334 ( .A(n3863), .B(m[126]), .Z(n4316) );
  NANDN U6335 ( .A(n3864), .B(creg[126]), .Z(n4315) );
  NAND U6336 ( .A(n4317), .B(n4318), .Z(y[125]) );
  NANDN U6337 ( .A(n3863), .B(m[125]), .Z(n4318) );
  NANDN U6338 ( .A(n3864), .B(creg[125]), .Z(n4317) );
  NAND U6339 ( .A(n4319), .B(n4320), .Z(y[124]) );
  NANDN U6340 ( .A(n3863), .B(m[124]), .Z(n4320) );
  NANDN U6341 ( .A(n3864), .B(creg[124]), .Z(n4319) );
  NAND U6342 ( .A(n4321), .B(n4322), .Z(y[123]) );
  NANDN U6343 ( .A(n3863), .B(m[123]), .Z(n4322) );
  NANDN U6344 ( .A(n3864), .B(creg[123]), .Z(n4321) );
  NAND U6345 ( .A(n4323), .B(n4324), .Z(y[122]) );
  NANDN U6346 ( .A(n3863), .B(m[122]), .Z(n4324) );
  NANDN U6347 ( .A(n3864), .B(creg[122]), .Z(n4323) );
  NAND U6348 ( .A(n4325), .B(n4326), .Z(y[121]) );
  NANDN U6349 ( .A(n3863), .B(m[121]), .Z(n4326) );
  NANDN U6350 ( .A(n3864), .B(creg[121]), .Z(n4325) );
  NAND U6351 ( .A(n4327), .B(n4328), .Z(y[120]) );
  NANDN U6352 ( .A(n3863), .B(m[120]), .Z(n4328) );
  NANDN U6353 ( .A(n3864), .B(creg[120]), .Z(n4327) );
  NAND U6354 ( .A(n4329), .B(n4330), .Z(y[11]) );
  NANDN U6355 ( .A(n3863), .B(m[11]), .Z(n4330) );
  NANDN U6356 ( .A(n3864), .B(creg[11]), .Z(n4329) );
  NAND U6357 ( .A(n4331), .B(n4332), .Z(y[119]) );
  NANDN U6358 ( .A(n3863), .B(m[119]), .Z(n4332) );
  NANDN U6359 ( .A(n3864), .B(creg[119]), .Z(n4331) );
  NAND U6360 ( .A(n4333), .B(n4334), .Z(y[118]) );
  NANDN U6361 ( .A(n3863), .B(m[118]), .Z(n4334) );
  NANDN U6362 ( .A(n3864), .B(creg[118]), .Z(n4333) );
  NAND U6363 ( .A(n4335), .B(n4336), .Z(y[117]) );
  NANDN U6364 ( .A(n3863), .B(m[117]), .Z(n4336) );
  NANDN U6365 ( .A(n3864), .B(creg[117]), .Z(n4335) );
  NAND U6366 ( .A(n4337), .B(n4338), .Z(y[116]) );
  NANDN U6367 ( .A(n3863), .B(m[116]), .Z(n4338) );
  NANDN U6368 ( .A(n3864), .B(creg[116]), .Z(n4337) );
  NAND U6369 ( .A(n4339), .B(n4340), .Z(y[115]) );
  NANDN U6370 ( .A(n3863), .B(m[115]), .Z(n4340) );
  NANDN U6371 ( .A(n3864), .B(creg[115]), .Z(n4339) );
  NAND U6372 ( .A(n4341), .B(n4342), .Z(y[114]) );
  NANDN U6373 ( .A(n3863), .B(m[114]), .Z(n4342) );
  NANDN U6374 ( .A(n3864), .B(creg[114]), .Z(n4341) );
  NAND U6375 ( .A(n4343), .B(n4344), .Z(y[113]) );
  NANDN U6376 ( .A(n3863), .B(m[113]), .Z(n4344) );
  NANDN U6377 ( .A(n3864), .B(creg[113]), .Z(n4343) );
  NAND U6378 ( .A(n4345), .B(n4346), .Z(y[112]) );
  NANDN U6379 ( .A(n3863), .B(m[112]), .Z(n4346) );
  NANDN U6380 ( .A(n3864), .B(creg[112]), .Z(n4345) );
  NAND U6381 ( .A(n4347), .B(n4348), .Z(y[111]) );
  NANDN U6382 ( .A(n3863), .B(m[111]), .Z(n4348) );
  NANDN U6383 ( .A(n3864), .B(creg[111]), .Z(n4347) );
  NAND U6384 ( .A(n4349), .B(n4350), .Z(y[110]) );
  NANDN U6385 ( .A(n3863), .B(m[110]), .Z(n4350) );
  NANDN U6386 ( .A(n3864), .B(creg[110]), .Z(n4349) );
  NAND U6387 ( .A(n4351), .B(n4352), .Z(y[10]) );
  NANDN U6388 ( .A(n3863), .B(m[10]), .Z(n4352) );
  NANDN U6389 ( .A(n3864), .B(creg[10]), .Z(n4351) );
  NAND U6390 ( .A(n4353), .B(n4354), .Z(y[109]) );
  NANDN U6391 ( .A(n3863), .B(m[109]), .Z(n4354) );
  NANDN U6392 ( .A(n3864), .B(creg[109]), .Z(n4353) );
  NAND U6393 ( .A(n4355), .B(n4356), .Z(y[108]) );
  NANDN U6394 ( .A(n3863), .B(m[108]), .Z(n4356) );
  NANDN U6395 ( .A(n3864), .B(creg[108]), .Z(n4355) );
  NAND U6396 ( .A(n4357), .B(n4358), .Z(y[107]) );
  NANDN U6397 ( .A(n3863), .B(m[107]), .Z(n4358) );
  NANDN U6398 ( .A(n3864), .B(creg[107]), .Z(n4357) );
  NAND U6399 ( .A(n4359), .B(n4360), .Z(y[106]) );
  NANDN U6400 ( .A(n3863), .B(m[106]), .Z(n4360) );
  NANDN U6401 ( .A(n3864), .B(creg[106]), .Z(n4359) );
  NAND U6402 ( .A(n4361), .B(n4362), .Z(y[105]) );
  NANDN U6403 ( .A(n3863), .B(m[105]), .Z(n4362) );
  NANDN U6404 ( .A(n3864), .B(creg[105]), .Z(n4361) );
  NAND U6405 ( .A(n4363), .B(n4364), .Z(y[104]) );
  NANDN U6406 ( .A(n3863), .B(m[104]), .Z(n4364) );
  NANDN U6407 ( .A(n3864), .B(creg[104]), .Z(n4363) );
  NAND U6408 ( .A(n4365), .B(n4366), .Z(y[103]) );
  NANDN U6409 ( .A(n3863), .B(m[103]), .Z(n4366) );
  NANDN U6410 ( .A(n3864), .B(creg[103]), .Z(n4365) );
  NAND U6411 ( .A(n4367), .B(n4368), .Z(y[102]) );
  NANDN U6412 ( .A(n3863), .B(m[102]), .Z(n4368) );
  NANDN U6413 ( .A(n3864), .B(creg[102]), .Z(n4367) );
  NAND U6414 ( .A(n4369), .B(n4370), .Z(y[101]) );
  NANDN U6415 ( .A(n3863), .B(m[101]), .Z(n4370) );
  NANDN U6416 ( .A(n3864), .B(creg[101]), .Z(n4369) );
  NAND U6417 ( .A(n4371), .B(n4372), .Z(y[100]) );
  NANDN U6418 ( .A(n3863), .B(m[100]), .Z(n4372) );
  NANDN U6419 ( .A(n3864), .B(creg[100]), .Z(n4371) );
  NAND U6420 ( .A(n4373), .B(n4374), .Z(y[0]) );
  NANDN U6421 ( .A(n3863), .B(m[0]), .Z(n4374) );
  NANDN U6422 ( .A(n3864), .B(creg[0]), .Z(n4373) );
  NAND U6423 ( .A(n4375), .B(n4376), .Z(x[9]) );
  NANDN U6424 ( .A(n4377), .B(creg[9]), .Z(n4375) );
  NAND U6425 ( .A(n4378), .B(n4379), .Z(x[99]) );
  NANDN U6426 ( .A(n4377), .B(creg[99]), .Z(n4378) );
  NAND U6427 ( .A(n4380), .B(n4381), .Z(x[98]) );
  NANDN U6428 ( .A(n4377), .B(creg[98]), .Z(n4380) );
  NAND U6429 ( .A(n4382), .B(n4383), .Z(x[97]) );
  NANDN U6430 ( .A(n4377), .B(creg[97]), .Z(n4382) );
  NAND U6431 ( .A(n4384), .B(n4385), .Z(x[96]) );
  NANDN U6432 ( .A(n4377), .B(creg[96]), .Z(n4384) );
  NAND U6433 ( .A(n4386), .B(n4387), .Z(x[95]) );
  NANDN U6434 ( .A(n4377), .B(creg[95]), .Z(n4386) );
  NAND U6435 ( .A(n4388), .B(n4389), .Z(x[94]) );
  NANDN U6436 ( .A(n4377), .B(creg[94]), .Z(n4388) );
  NAND U6437 ( .A(n4390), .B(n4391), .Z(x[93]) );
  NANDN U6438 ( .A(n4377), .B(creg[93]), .Z(n4390) );
  NAND U6439 ( .A(n4392), .B(n4393), .Z(x[92]) );
  NANDN U6440 ( .A(n4377), .B(creg[92]), .Z(n4392) );
  NAND U6441 ( .A(n4394), .B(n4395), .Z(x[91]) );
  NANDN U6442 ( .A(n4377), .B(creg[91]), .Z(n4394) );
  NAND U6443 ( .A(n4396), .B(n4397), .Z(x[90]) );
  NANDN U6444 ( .A(n4377), .B(creg[90]), .Z(n4396) );
  NAND U6445 ( .A(n4398), .B(n4399), .Z(x[8]) );
  NANDN U6446 ( .A(n4377), .B(creg[8]), .Z(n4398) );
  NAND U6447 ( .A(n4400), .B(n4401), .Z(x[89]) );
  NANDN U6448 ( .A(n4377), .B(creg[89]), .Z(n4400) );
  NAND U6449 ( .A(n4402), .B(n4403), .Z(x[88]) );
  NANDN U6450 ( .A(n4377), .B(creg[88]), .Z(n4402) );
  NAND U6451 ( .A(n4404), .B(n4405), .Z(x[87]) );
  NANDN U6452 ( .A(n4377), .B(creg[87]), .Z(n4404) );
  NAND U6453 ( .A(n4406), .B(n4407), .Z(x[86]) );
  NANDN U6454 ( .A(n4377), .B(creg[86]), .Z(n4406) );
  NAND U6455 ( .A(n4408), .B(n4409), .Z(x[85]) );
  NANDN U6456 ( .A(n4377), .B(creg[85]), .Z(n4408) );
  NAND U6457 ( .A(n4410), .B(n4411), .Z(x[84]) );
  NANDN U6458 ( .A(n4377), .B(creg[84]), .Z(n4410) );
  NAND U6459 ( .A(n4412), .B(n4413), .Z(x[83]) );
  NANDN U6460 ( .A(n4377), .B(creg[83]), .Z(n4412) );
  NAND U6461 ( .A(n4414), .B(n4415), .Z(x[82]) );
  NANDN U6462 ( .A(n4377), .B(creg[82]), .Z(n4414) );
  NAND U6463 ( .A(n4416), .B(n4417), .Z(x[81]) );
  NANDN U6464 ( .A(n4377), .B(creg[81]), .Z(n4416) );
  NAND U6465 ( .A(n4418), .B(n4419), .Z(x[80]) );
  NANDN U6466 ( .A(n4377), .B(creg[80]), .Z(n4418) );
  NAND U6467 ( .A(n4420), .B(n4421), .Z(x[7]) );
  NANDN U6468 ( .A(n4377), .B(creg[7]), .Z(n4420) );
  NAND U6469 ( .A(n4422), .B(n4423), .Z(x[79]) );
  NANDN U6470 ( .A(n4377), .B(creg[79]), .Z(n4422) );
  NAND U6471 ( .A(n4424), .B(n4425), .Z(x[78]) );
  NANDN U6472 ( .A(n4377), .B(creg[78]), .Z(n4424) );
  NAND U6473 ( .A(n4426), .B(n4427), .Z(x[77]) );
  NANDN U6474 ( .A(n4377), .B(creg[77]), .Z(n4426) );
  NAND U6475 ( .A(n4428), .B(n4429), .Z(x[76]) );
  NANDN U6476 ( .A(n4377), .B(creg[76]), .Z(n4428) );
  NAND U6477 ( .A(n4430), .B(n4431), .Z(x[75]) );
  NANDN U6478 ( .A(n4377), .B(creg[75]), .Z(n4430) );
  NAND U6479 ( .A(n4432), .B(n4433), .Z(x[74]) );
  NANDN U6480 ( .A(n4377), .B(creg[74]), .Z(n4432) );
  NAND U6481 ( .A(n4434), .B(n4435), .Z(x[73]) );
  NANDN U6482 ( .A(n4377), .B(creg[73]), .Z(n4434) );
  NAND U6483 ( .A(n4436), .B(n4437), .Z(x[72]) );
  NANDN U6484 ( .A(n4377), .B(creg[72]), .Z(n4436) );
  NAND U6485 ( .A(n4438), .B(n4439), .Z(x[71]) );
  NANDN U6486 ( .A(n4377), .B(creg[71]), .Z(n4438) );
  NAND U6487 ( .A(n4440), .B(n4441), .Z(x[70]) );
  NANDN U6488 ( .A(n4377), .B(creg[70]), .Z(n4440) );
  NAND U6489 ( .A(n4442), .B(n4443), .Z(x[6]) );
  NANDN U6490 ( .A(n4377), .B(creg[6]), .Z(n4442) );
  NAND U6491 ( .A(n4444), .B(n4445), .Z(x[69]) );
  NANDN U6492 ( .A(n4377), .B(creg[69]), .Z(n4444) );
  NAND U6493 ( .A(n4446), .B(n4447), .Z(x[68]) );
  NANDN U6494 ( .A(n4377), .B(creg[68]), .Z(n4446) );
  NAND U6495 ( .A(n4448), .B(n4449), .Z(x[67]) );
  NANDN U6496 ( .A(n4377), .B(creg[67]), .Z(n4448) );
  NAND U6497 ( .A(n4450), .B(n4451), .Z(x[66]) );
  NANDN U6498 ( .A(n4377), .B(creg[66]), .Z(n4450) );
  NAND U6499 ( .A(n4452), .B(n4453), .Z(x[65]) );
  NANDN U6500 ( .A(n4377), .B(creg[65]), .Z(n4452) );
  NAND U6501 ( .A(n4454), .B(n4455), .Z(x[64]) );
  NANDN U6502 ( .A(n4377), .B(creg[64]), .Z(n4454) );
  NAND U6503 ( .A(n4456), .B(n4457), .Z(x[63]) );
  NANDN U6504 ( .A(n4377), .B(creg[63]), .Z(n4456) );
  NAND U6505 ( .A(n4458), .B(n4459), .Z(x[62]) );
  NANDN U6506 ( .A(n4377), .B(creg[62]), .Z(n4458) );
  NAND U6507 ( .A(n4460), .B(n4461), .Z(x[61]) );
  NANDN U6508 ( .A(n4377), .B(creg[61]), .Z(n4460) );
  NAND U6509 ( .A(n4462), .B(n4463), .Z(x[60]) );
  NANDN U6510 ( .A(n4377), .B(creg[60]), .Z(n4462) );
  NAND U6511 ( .A(n4464), .B(n4465), .Z(x[5]) );
  NANDN U6512 ( .A(n4377), .B(creg[5]), .Z(n4464) );
  NAND U6513 ( .A(n4466), .B(n4467), .Z(x[59]) );
  NANDN U6514 ( .A(n4377), .B(creg[59]), .Z(n4466) );
  NAND U6515 ( .A(n4468), .B(n4469), .Z(x[58]) );
  NANDN U6516 ( .A(n4377), .B(creg[58]), .Z(n4468) );
  NAND U6517 ( .A(n4470), .B(n4471), .Z(x[57]) );
  NANDN U6518 ( .A(n4377), .B(creg[57]), .Z(n4470) );
  NAND U6519 ( .A(n4472), .B(n4473), .Z(x[56]) );
  NANDN U6520 ( .A(n4377), .B(creg[56]), .Z(n4472) );
  NAND U6521 ( .A(n4474), .B(n4475), .Z(x[55]) );
  NANDN U6522 ( .A(n4377), .B(creg[55]), .Z(n4474) );
  NAND U6523 ( .A(n4476), .B(n4477), .Z(x[54]) );
  NANDN U6524 ( .A(n4377), .B(creg[54]), .Z(n4476) );
  NAND U6525 ( .A(n4478), .B(n4479), .Z(x[53]) );
  NANDN U6526 ( .A(n4377), .B(creg[53]), .Z(n4478) );
  NAND U6527 ( .A(n4480), .B(n4481), .Z(x[52]) );
  NANDN U6528 ( .A(n4377), .B(creg[52]), .Z(n4480) );
  NAND U6529 ( .A(n4482), .B(n4483), .Z(x[51]) );
  NANDN U6530 ( .A(n4377), .B(creg[51]), .Z(n4482) );
  NAND U6531 ( .A(n4484), .B(n4485), .Z(x[50]) );
  NANDN U6532 ( .A(n4377), .B(creg[50]), .Z(n4484) );
  NAND U6533 ( .A(n4486), .B(n4487), .Z(x[4]) );
  NANDN U6534 ( .A(n4377), .B(creg[4]), .Z(n4486) );
  NAND U6535 ( .A(n4488), .B(n4489), .Z(x[49]) );
  NANDN U6536 ( .A(n4377), .B(creg[49]), .Z(n4488) );
  NAND U6537 ( .A(n4490), .B(n4491), .Z(x[48]) );
  NANDN U6538 ( .A(n4377), .B(creg[48]), .Z(n4490) );
  NAND U6539 ( .A(n4492), .B(n4493), .Z(x[47]) );
  NANDN U6540 ( .A(n4377), .B(creg[47]), .Z(n4492) );
  NAND U6541 ( .A(n4494), .B(n4495), .Z(x[46]) );
  NANDN U6542 ( .A(n4377), .B(creg[46]), .Z(n4494) );
  NAND U6543 ( .A(n4496), .B(n4497), .Z(x[45]) );
  NANDN U6544 ( .A(n4377), .B(creg[45]), .Z(n4496) );
  NAND U6545 ( .A(n4498), .B(n4499), .Z(x[44]) );
  NANDN U6546 ( .A(n4377), .B(creg[44]), .Z(n4498) );
  NAND U6547 ( .A(n4500), .B(n4501), .Z(x[43]) );
  NANDN U6548 ( .A(n4377), .B(creg[43]), .Z(n4500) );
  NAND U6549 ( .A(n4502), .B(n4503), .Z(x[42]) );
  NANDN U6550 ( .A(n4377), .B(creg[42]), .Z(n4502) );
  NAND U6551 ( .A(n4504), .B(n4505), .Z(x[41]) );
  NANDN U6552 ( .A(n4377), .B(creg[41]), .Z(n4504) );
  NAND U6553 ( .A(n4506), .B(n4507), .Z(x[40]) );
  NANDN U6554 ( .A(n4377), .B(creg[40]), .Z(n4506) );
  NAND U6555 ( .A(n4508), .B(n4509), .Z(x[3]) );
  NANDN U6556 ( .A(n4377), .B(creg[3]), .Z(n4508) );
  NAND U6557 ( .A(n4510), .B(n4511), .Z(x[39]) );
  NANDN U6558 ( .A(n4377), .B(creg[39]), .Z(n4510) );
  NAND U6559 ( .A(n4512), .B(n4513), .Z(x[38]) );
  NANDN U6560 ( .A(n4377), .B(creg[38]), .Z(n4512) );
  NAND U6561 ( .A(n4514), .B(n4515), .Z(x[37]) );
  NANDN U6562 ( .A(n4377), .B(creg[37]), .Z(n4514) );
  NAND U6563 ( .A(n4516), .B(n4517), .Z(x[36]) );
  NANDN U6564 ( .A(n4377), .B(creg[36]), .Z(n4516) );
  NAND U6565 ( .A(n4518), .B(n4519), .Z(x[35]) );
  NANDN U6566 ( .A(n4377), .B(creg[35]), .Z(n4518) );
  NAND U6567 ( .A(n4520), .B(n4521), .Z(x[34]) );
  NANDN U6568 ( .A(n4377), .B(creg[34]), .Z(n4520) );
  NAND U6569 ( .A(n4522), .B(n4523), .Z(x[33]) );
  NANDN U6570 ( .A(n4377), .B(creg[33]), .Z(n4522) );
  NAND U6571 ( .A(n4524), .B(n4525), .Z(x[32]) );
  NANDN U6572 ( .A(n4377), .B(creg[32]), .Z(n4524) );
  NAND U6573 ( .A(n4526), .B(n4527), .Z(x[31]) );
  NANDN U6574 ( .A(n4377), .B(creg[31]), .Z(n4526) );
  NAND U6575 ( .A(n4528), .B(n4529), .Z(x[30]) );
  NANDN U6576 ( .A(n4377), .B(creg[30]), .Z(n4528) );
  NAND U6577 ( .A(n4530), .B(n4531), .Z(x[2]) );
  NANDN U6578 ( .A(n4377), .B(creg[2]), .Z(n4530) );
  NAND U6579 ( .A(n4532), .B(n4533), .Z(x[29]) );
  NANDN U6580 ( .A(n4377), .B(creg[29]), .Z(n4532) );
  NAND U6581 ( .A(n4534), .B(n4535), .Z(x[28]) );
  NANDN U6582 ( .A(n4377), .B(creg[28]), .Z(n4534) );
  NAND U6583 ( .A(n4536), .B(n4537), .Z(x[27]) );
  NANDN U6584 ( .A(n4377), .B(creg[27]), .Z(n4536) );
  NAND U6585 ( .A(n4538), .B(n4539), .Z(x[26]) );
  NANDN U6586 ( .A(n4377), .B(creg[26]), .Z(n4538) );
  NAND U6587 ( .A(n4540), .B(n4541), .Z(x[25]) );
  NANDN U6588 ( .A(n4377), .B(creg[25]), .Z(n4540) );
  NAND U6589 ( .A(n4542), .B(n4543), .Z(x[255]) );
  NANDN U6590 ( .A(n4377), .B(creg[255]), .Z(n4542) );
  NAND U6591 ( .A(n4544), .B(n4545), .Z(x[254]) );
  NANDN U6592 ( .A(n4377), .B(creg[254]), .Z(n4544) );
  NAND U6593 ( .A(n4546), .B(n4547), .Z(x[253]) );
  NANDN U6594 ( .A(n4377), .B(creg[253]), .Z(n4546) );
  NAND U6595 ( .A(n4548), .B(n4549), .Z(x[252]) );
  NANDN U6596 ( .A(n4377), .B(creg[252]), .Z(n4548) );
  NAND U6597 ( .A(n4550), .B(n4551), .Z(x[251]) );
  NANDN U6598 ( .A(n4377), .B(creg[251]), .Z(n4550) );
  NAND U6599 ( .A(n4552), .B(n4553), .Z(x[250]) );
  NANDN U6600 ( .A(n4377), .B(creg[250]), .Z(n4552) );
  NAND U6601 ( .A(n4554), .B(n4555), .Z(x[24]) );
  NANDN U6602 ( .A(n4377), .B(creg[24]), .Z(n4554) );
  NAND U6603 ( .A(n4556), .B(n4557), .Z(x[249]) );
  NANDN U6604 ( .A(n4377), .B(creg[249]), .Z(n4556) );
  NAND U6605 ( .A(n4558), .B(n4559), .Z(x[248]) );
  NANDN U6606 ( .A(n4377), .B(creg[248]), .Z(n4558) );
  NAND U6607 ( .A(n4560), .B(n4561), .Z(x[247]) );
  NANDN U6608 ( .A(n4377), .B(creg[247]), .Z(n4560) );
  NAND U6609 ( .A(n4562), .B(n4563), .Z(x[246]) );
  NANDN U6610 ( .A(n4377), .B(creg[246]), .Z(n4562) );
  NAND U6611 ( .A(n4564), .B(n4565), .Z(x[245]) );
  NANDN U6612 ( .A(n4377), .B(creg[245]), .Z(n4564) );
  NAND U6613 ( .A(n4566), .B(n4567), .Z(x[244]) );
  NANDN U6614 ( .A(n4377), .B(creg[244]), .Z(n4566) );
  NAND U6615 ( .A(n4568), .B(n4569), .Z(x[243]) );
  NANDN U6616 ( .A(n4377), .B(creg[243]), .Z(n4568) );
  NAND U6617 ( .A(n4570), .B(n4571), .Z(x[242]) );
  NANDN U6618 ( .A(n4377), .B(creg[242]), .Z(n4570) );
  NAND U6619 ( .A(n4572), .B(n4573), .Z(x[241]) );
  NANDN U6620 ( .A(n4377), .B(creg[241]), .Z(n4572) );
  NAND U6621 ( .A(n4574), .B(n4575), .Z(x[240]) );
  NANDN U6622 ( .A(n4377), .B(creg[240]), .Z(n4574) );
  NAND U6623 ( .A(n4576), .B(n4577), .Z(x[23]) );
  NANDN U6624 ( .A(n4377), .B(creg[23]), .Z(n4576) );
  NAND U6625 ( .A(n4578), .B(n4579), .Z(x[239]) );
  NANDN U6626 ( .A(n4377), .B(creg[239]), .Z(n4578) );
  NAND U6627 ( .A(n4580), .B(n4581), .Z(x[238]) );
  NANDN U6628 ( .A(n4377), .B(creg[238]), .Z(n4580) );
  NAND U6629 ( .A(n4582), .B(n4583), .Z(x[237]) );
  NANDN U6630 ( .A(n4377), .B(creg[237]), .Z(n4582) );
  NAND U6631 ( .A(n4584), .B(n4585), .Z(x[236]) );
  NANDN U6632 ( .A(n4377), .B(creg[236]), .Z(n4584) );
  NAND U6633 ( .A(n4586), .B(n4587), .Z(x[235]) );
  NANDN U6634 ( .A(n4377), .B(creg[235]), .Z(n4586) );
  NAND U6635 ( .A(n4588), .B(n4589), .Z(x[234]) );
  NANDN U6636 ( .A(n4377), .B(creg[234]), .Z(n4588) );
  NAND U6637 ( .A(n4590), .B(n4591), .Z(x[233]) );
  NANDN U6638 ( .A(n4377), .B(creg[233]), .Z(n4590) );
  NAND U6639 ( .A(n4592), .B(n4593), .Z(x[232]) );
  NANDN U6640 ( .A(n4377), .B(creg[232]), .Z(n4592) );
  NAND U6641 ( .A(n4594), .B(n4595), .Z(x[231]) );
  NANDN U6642 ( .A(n4377), .B(creg[231]), .Z(n4594) );
  NAND U6643 ( .A(n4596), .B(n4597), .Z(x[230]) );
  NANDN U6644 ( .A(n4377), .B(creg[230]), .Z(n4596) );
  NAND U6645 ( .A(n4598), .B(n4599), .Z(x[22]) );
  NANDN U6646 ( .A(n4377), .B(creg[22]), .Z(n4598) );
  NAND U6647 ( .A(n4600), .B(n4601), .Z(x[229]) );
  NANDN U6648 ( .A(n4377), .B(creg[229]), .Z(n4600) );
  NAND U6649 ( .A(n4602), .B(n4603), .Z(x[228]) );
  NANDN U6650 ( .A(n4377), .B(creg[228]), .Z(n4602) );
  NAND U6651 ( .A(n4604), .B(n4605), .Z(x[227]) );
  NANDN U6652 ( .A(n4377), .B(creg[227]), .Z(n4604) );
  NAND U6653 ( .A(n4606), .B(n4607), .Z(x[226]) );
  NANDN U6654 ( .A(n4377), .B(creg[226]), .Z(n4606) );
  NAND U6655 ( .A(n4608), .B(n4609), .Z(x[225]) );
  NANDN U6656 ( .A(n4377), .B(creg[225]), .Z(n4608) );
  NAND U6657 ( .A(n4610), .B(n4611), .Z(x[224]) );
  NANDN U6658 ( .A(n4377), .B(creg[224]), .Z(n4610) );
  NAND U6659 ( .A(n4612), .B(n4613), .Z(x[223]) );
  NANDN U6660 ( .A(n4377), .B(creg[223]), .Z(n4612) );
  NAND U6661 ( .A(n4614), .B(n4615), .Z(x[222]) );
  NANDN U6662 ( .A(n4377), .B(creg[222]), .Z(n4614) );
  NAND U6663 ( .A(n4616), .B(n4617), .Z(x[221]) );
  NANDN U6664 ( .A(n4377), .B(creg[221]), .Z(n4616) );
  NAND U6665 ( .A(n4618), .B(n4619), .Z(x[220]) );
  NANDN U6666 ( .A(n4377), .B(creg[220]), .Z(n4618) );
  NAND U6667 ( .A(n4620), .B(n4621), .Z(x[21]) );
  NANDN U6668 ( .A(n4377), .B(creg[21]), .Z(n4620) );
  NAND U6669 ( .A(n4622), .B(n4623), .Z(x[219]) );
  NANDN U6670 ( .A(n4377), .B(creg[219]), .Z(n4622) );
  NAND U6671 ( .A(n4624), .B(n4625), .Z(x[218]) );
  NANDN U6672 ( .A(n4377), .B(creg[218]), .Z(n4624) );
  NAND U6673 ( .A(n4626), .B(n4627), .Z(x[217]) );
  NANDN U6674 ( .A(n4377), .B(creg[217]), .Z(n4626) );
  NAND U6675 ( .A(n4628), .B(n4629), .Z(x[216]) );
  NANDN U6676 ( .A(n4377), .B(creg[216]), .Z(n4628) );
  NAND U6677 ( .A(n4630), .B(n4631), .Z(x[215]) );
  NANDN U6678 ( .A(n4377), .B(creg[215]), .Z(n4630) );
  NAND U6679 ( .A(n4632), .B(n4633), .Z(x[214]) );
  NANDN U6680 ( .A(n4377), .B(creg[214]), .Z(n4632) );
  NAND U6681 ( .A(n4634), .B(n4635), .Z(x[213]) );
  NANDN U6682 ( .A(n4377), .B(creg[213]), .Z(n4634) );
  NAND U6683 ( .A(n4636), .B(n4637), .Z(x[212]) );
  NANDN U6684 ( .A(n4377), .B(creg[212]), .Z(n4636) );
  NAND U6685 ( .A(n4638), .B(n4639), .Z(x[211]) );
  NANDN U6686 ( .A(n4377), .B(creg[211]), .Z(n4638) );
  NAND U6687 ( .A(n4640), .B(n4641), .Z(x[210]) );
  NANDN U6688 ( .A(n4377), .B(creg[210]), .Z(n4640) );
  NAND U6689 ( .A(n4642), .B(n4643), .Z(x[20]) );
  NANDN U6690 ( .A(n4377), .B(creg[20]), .Z(n4642) );
  NAND U6691 ( .A(n4644), .B(n4645), .Z(x[209]) );
  NANDN U6692 ( .A(n4377), .B(creg[209]), .Z(n4644) );
  NAND U6693 ( .A(n4646), .B(n4647), .Z(x[208]) );
  NANDN U6694 ( .A(n4377), .B(creg[208]), .Z(n4646) );
  NAND U6695 ( .A(n4648), .B(n4649), .Z(x[207]) );
  NANDN U6696 ( .A(n4377), .B(creg[207]), .Z(n4648) );
  NAND U6697 ( .A(n4650), .B(n4651), .Z(x[206]) );
  NANDN U6698 ( .A(n4377), .B(creg[206]), .Z(n4650) );
  NAND U6699 ( .A(n4652), .B(n4653), .Z(x[205]) );
  NANDN U6700 ( .A(n4377), .B(creg[205]), .Z(n4652) );
  NAND U6701 ( .A(n4654), .B(n4655), .Z(x[204]) );
  NANDN U6702 ( .A(n4377), .B(creg[204]), .Z(n4654) );
  NAND U6703 ( .A(n4656), .B(n4657), .Z(x[203]) );
  NANDN U6704 ( .A(n4377), .B(creg[203]), .Z(n4656) );
  NAND U6705 ( .A(n4658), .B(n4659), .Z(x[202]) );
  NANDN U6706 ( .A(n4377), .B(creg[202]), .Z(n4658) );
  NAND U6707 ( .A(n4660), .B(n4661), .Z(x[201]) );
  NANDN U6708 ( .A(n4377), .B(creg[201]), .Z(n4660) );
  NAND U6709 ( .A(n4662), .B(n4663), .Z(x[200]) );
  NANDN U6710 ( .A(n4377), .B(creg[200]), .Z(n4662) );
  NAND U6711 ( .A(n4664), .B(n4665), .Z(x[1]) );
  NANDN U6712 ( .A(n4377), .B(creg[1]), .Z(n4664) );
  NAND U6713 ( .A(n4666), .B(n4667), .Z(x[19]) );
  NANDN U6714 ( .A(n4377), .B(creg[19]), .Z(n4666) );
  NAND U6715 ( .A(n4668), .B(n4669), .Z(x[199]) );
  NANDN U6716 ( .A(n4377), .B(creg[199]), .Z(n4668) );
  NAND U6717 ( .A(n4670), .B(n4671), .Z(x[198]) );
  NANDN U6718 ( .A(n4377), .B(creg[198]), .Z(n4670) );
  NAND U6719 ( .A(n4672), .B(n4673), .Z(x[197]) );
  NANDN U6720 ( .A(n4377), .B(creg[197]), .Z(n4672) );
  NAND U6721 ( .A(n4674), .B(n4675), .Z(x[196]) );
  NANDN U6722 ( .A(n4377), .B(creg[196]), .Z(n4674) );
  NAND U6723 ( .A(n4676), .B(n4677), .Z(x[195]) );
  NANDN U6724 ( .A(n4377), .B(creg[195]), .Z(n4676) );
  NAND U6725 ( .A(n4678), .B(n4679), .Z(x[194]) );
  NANDN U6726 ( .A(n4377), .B(creg[194]), .Z(n4678) );
  NAND U6727 ( .A(n4680), .B(n4681), .Z(x[193]) );
  NANDN U6728 ( .A(n4377), .B(creg[193]), .Z(n4680) );
  NAND U6729 ( .A(n4682), .B(n4683), .Z(x[192]) );
  NANDN U6730 ( .A(n4377), .B(creg[192]), .Z(n4682) );
  NAND U6731 ( .A(n4684), .B(n4685), .Z(x[191]) );
  NANDN U6732 ( .A(n4377), .B(creg[191]), .Z(n4684) );
  NAND U6733 ( .A(n4686), .B(n4687), .Z(x[190]) );
  NANDN U6734 ( .A(n4377), .B(creg[190]), .Z(n4686) );
  NAND U6735 ( .A(n4688), .B(n4689), .Z(x[18]) );
  NANDN U6736 ( .A(n4377), .B(creg[18]), .Z(n4688) );
  NAND U6737 ( .A(n4690), .B(n4691), .Z(x[189]) );
  NANDN U6738 ( .A(n4377), .B(creg[189]), .Z(n4690) );
  NAND U6739 ( .A(n4692), .B(n4693), .Z(x[188]) );
  NANDN U6740 ( .A(n4377), .B(creg[188]), .Z(n4692) );
  NAND U6741 ( .A(n4694), .B(n4695), .Z(x[187]) );
  NANDN U6742 ( .A(n4377), .B(creg[187]), .Z(n4694) );
  NAND U6743 ( .A(n4696), .B(n4697), .Z(x[186]) );
  NANDN U6744 ( .A(n4377), .B(creg[186]), .Z(n4696) );
  NAND U6745 ( .A(n4698), .B(n4699), .Z(x[185]) );
  NANDN U6746 ( .A(n4377), .B(creg[185]), .Z(n4698) );
  NAND U6747 ( .A(n4700), .B(n4701), .Z(x[184]) );
  NANDN U6748 ( .A(n4377), .B(creg[184]), .Z(n4700) );
  NAND U6749 ( .A(n4702), .B(n4703), .Z(x[183]) );
  NANDN U6750 ( .A(n4377), .B(creg[183]), .Z(n4702) );
  NAND U6751 ( .A(n4704), .B(n4705), .Z(x[182]) );
  NANDN U6752 ( .A(n4377), .B(creg[182]), .Z(n4704) );
  NAND U6753 ( .A(n4706), .B(n4707), .Z(x[181]) );
  NANDN U6754 ( .A(n4377), .B(creg[181]), .Z(n4706) );
  NAND U6755 ( .A(n4708), .B(n4709), .Z(x[180]) );
  NANDN U6756 ( .A(n4377), .B(creg[180]), .Z(n4708) );
  NAND U6757 ( .A(n4710), .B(n4711), .Z(x[17]) );
  NANDN U6758 ( .A(n4377), .B(creg[17]), .Z(n4710) );
  NAND U6759 ( .A(n4712), .B(n4713), .Z(x[179]) );
  NANDN U6760 ( .A(n4377), .B(creg[179]), .Z(n4712) );
  NAND U6761 ( .A(n4714), .B(n4715), .Z(x[178]) );
  NANDN U6762 ( .A(n4377), .B(creg[178]), .Z(n4714) );
  NAND U6763 ( .A(n4716), .B(n4717), .Z(x[177]) );
  NANDN U6764 ( .A(n4377), .B(creg[177]), .Z(n4716) );
  NAND U6765 ( .A(n4718), .B(n4719), .Z(x[176]) );
  NANDN U6766 ( .A(n4377), .B(creg[176]), .Z(n4718) );
  NAND U6767 ( .A(n4720), .B(n4721), .Z(x[175]) );
  NANDN U6768 ( .A(n4377), .B(creg[175]), .Z(n4720) );
  NAND U6769 ( .A(n4722), .B(n4723), .Z(x[174]) );
  NANDN U6770 ( .A(n4377), .B(creg[174]), .Z(n4722) );
  NAND U6771 ( .A(n4724), .B(n4725), .Z(x[173]) );
  NANDN U6772 ( .A(n4377), .B(creg[173]), .Z(n4724) );
  NAND U6773 ( .A(n4726), .B(n4727), .Z(x[172]) );
  NANDN U6774 ( .A(n4377), .B(creg[172]), .Z(n4726) );
  NAND U6775 ( .A(n4728), .B(n4729), .Z(x[171]) );
  NANDN U6776 ( .A(n4377), .B(creg[171]), .Z(n4728) );
  NAND U6777 ( .A(n4730), .B(n4731), .Z(x[170]) );
  NANDN U6778 ( .A(n4377), .B(creg[170]), .Z(n4730) );
  NAND U6779 ( .A(n4732), .B(n4733), .Z(x[16]) );
  NANDN U6780 ( .A(n4377), .B(creg[16]), .Z(n4732) );
  NAND U6781 ( .A(n4734), .B(n4735), .Z(x[169]) );
  NANDN U6782 ( .A(n4377), .B(creg[169]), .Z(n4734) );
  NAND U6783 ( .A(n4736), .B(n4737), .Z(x[168]) );
  NANDN U6784 ( .A(n4377), .B(creg[168]), .Z(n4736) );
  NAND U6785 ( .A(n4738), .B(n4739), .Z(x[167]) );
  NANDN U6786 ( .A(n4377), .B(creg[167]), .Z(n4738) );
  NAND U6787 ( .A(n4740), .B(n4741), .Z(x[166]) );
  NANDN U6788 ( .A(n4377), .B(creg[166]), .Z(n4740) );
  NAND U6789 ( .A(n4742), .B(n4743), .Z(x[165]) );
  NANDN U6790 ( .A(n4377), .B(creg[165]), .Z(n4742) );
  NAND U6791 ( .A(n4744), .B(n4745), .Z(x[164]) );
  NANDN U6792 ( .A(n4377), .B(creg[164]), .Z(n4744) );
  NAND U6793 ( .A(n4746), .B(n4747), .Z(x[163]) );
  NANDN U6794 ( .A(n4377), .B(creg[163]), .Z(n4746) );
  NAND U6795 ( .A(n4748), .B(n4749), .Z(x[162]) );
  NANDN U6796 ( .A(n4377), .B(creg[162]), .Z(n4748) );
  NAND U6797 ( .A(n4750), .B(n4751), .Z(x[161]) );
  NANDN U6798 ( .A(n4377), .B(creg[161]), .Z(n4750) );
  NAND U6799 ( .A(n4752), .B(n4753), .Z(x[160]) );
  NANDN U6800 ( .A(n4377), .B(creg[160]), .Z(n4752) );
  NAND U6801 ( .A(n4754), .B(n4755), .Z(x[15]) );
  NANDN U6802 ( .A(n4377), .B(creg[15]), .Z(n4754) );
  NAND U6803 ( .A(n4756), .B(n4757), .Z(x[159]) );
  NANDN U6804 ( .A(n4377), .B(creg[159]), .Z(n4756) );
  NAND U6805 ( .A(n4758), .B(n4759), .Z(x[158]) );
  NANDN U6806 ( .A(n4377), .B(creg[158]), .Z(n4758) );
  NAND U6807 ( .A(n4760), .B(n4761), .Z(x[157]) );
  NANDN U6808 ( .A(n4377), .B(creg[157]), .Z(n4760) );
  NAND U6809 ( .A(n4762), .B(n4763), .Z(x[156]) );
  NANDN U6810 ( .A(n4377), .B(creg[156]), .Z(n4762) );
  NAND U6811 ( .A(n4764), .B(n4765), .Z(x[155]) );
  NANDN U6812 ( .A(n4377), .B(creg[155]), .Z(n4764) );
  NAND U6813 ( .A(n4766), .B(n4767), .Z(x[154]) );
  NANDN U6814 ( .A(n4377), .B(creg[154]), .Z(n4766) );
  NAND U6815 ( .A(n4768), .B(n4769), .Z(x[153]) );
  NANDN U6816 ( .A(n4377), .B(creg[153]), .Z(n4768) );
  NAND U6817 ( .A(n4770), .B(n4771), .Z(x[152]) );
  NANDN U6818 ( .A(n4377), .B(creg[152]), .Z(n4770) );
  NAND U6819 ( .A(n4772), .B(n4773), .Z(x[151]) );
  NANDN U6820 ( .A(n4377), .B(creg[151]), .Z(n4772) );
  NAND U6821 ( .A(n4774), .B(n4775), .Z(x[150]) );
  NANDN U6822 ( .A(n4377), .B(creg[150]), .Z(n4774) );
  NAND U6823 ( .A(n4776), .B(n4777), .Z(x[14]) );
  NANDN U6824 ( .A(n4377), .B(creg[14]), .Z(n4776) );
  NAND U6825 ( .A(n4778), .B(n4779), .Z(x[149]) );
  NANDN U6826 ( .A(n4377), .B(creg[149]), .Z(n4778) );
  NAND U6827 ( .A(n4780), .B(n4781), .Z(x[148]) );
  NANDN U6828 ( .A(n4377), .B(creg[148]), .Z(n4780) );
  NAND U6829 ( .A(n4782), .B(n4783), .Z(x[147]) );
  NANDN U6830 ( .A(n4377), .B(creg[147]), .Z(n4782) );
  NAND U6831 ( .A(n4784), .B(n4785), .Z(x[146]) );
  NANDN U6832 ( .A(n4377), .B(creg[146]), .Z(n4784) );
  NAND U6833 ( .A(n4786), .B(n4787), .Z(x[145]) );
  NANDN U6834 ( .A(n4377), .B(creg[145]), .Z(n4786) );
  NAND U6835 ( .A(n4788), .B(n4789), .Z(x[144]) );
  NANDN U6836 ( .A(n4377), .B(creg[144]), .Z(n4788) );
  NAND U6837 ( .A(n4790), .B(n4791), .Z(x[143]) );
  NANDN U6838 ( .A(n4377), .B(creg[143]), .Z(n4790) );
  NAND U6839 ( .A(n4792), .B(n4793), .Z(x[142]) );
  NANDN U6840 ( .A(n4377), .B(creg[142]), .Z(n4792) );
  NAND U6841 ( .A(n4794), .B(n4795), .Z(x[141]) );
  NANDN U6842 ( .A(n4377), .B(creg[141]), .Z(n4794) );
  NAND U6843 ( .A(n4796), .B(n4797), .Z(x[140]) );
  NANDN U6844 ( .A(n4377), .B(creg[140]), .Z(n4796) );
  NAND U6845 ( .A(n4798), .B(n4799), .Z(x[13]) );
  NANDN U6846 ( .A(n4377), .B(creg[13]), .Z(n4798) );
  NAND U6847 ( .A(n4800), .B(n4801), .Z(x[139]) );
  NANDN U6848 ( .A(n4377), .B(creg[139]), .Z(n4800) );
  NAND U6849 ( .A(n4802), .B(n4803), .Z(x[138]) );
  NANDN U6850 ( .A(n4377), .B(creg[138]), .Z(n4802) );
  NAND U6851 ( .A(n4804), .B(n4805), .Z(x[137]) );
  NANDN U6852 ( .A(n4377), .B(creg[137]), .Z(n4804) );
  NAND U6853 ( .A(n4806), .B(n4807), .Z(x[136]) );
  NANDN U6854 ( .A(n4377), .B(creg[136]), .Z(n4806) );
  NAND U6855 ( .A(n4808), .B(n4809), .Z(x[135]) );
  NANDN U6856 ( .A(n4377), .B(creg[135]), .Z(n4808) );
  NAND U6857 ( .A(n4810), .B(n4811), .Z(x[134]) );
  NANDN U6858 ( .A(n4377), .B(creg[134]), .Z(n4810) );
  NAND U6859 ( .A(n4812), .B(n4813), .Z(x[133]) );
  NANDN U6860 ( .A(n4377), .B(creg[133]), .Z(n4812) );
  NAND U6861 ( .A(n4814), .B(n4815), .Z(x[132]) );
  NANDN U6862 ( .A(n4377), .B(creg[132]), .Z(n4814) );
  NAND U6863 ( .A(n4816), .B(n4817), .Z(x[131]) );
  NANDN U6864 ( .A(n4377), .B(creg[131]), .Z(n4816) );
  NAND U6865 ( .A(n4818), .B(n4819), .Z(x[130]) );
  NANDN U6866 ( .A(n4377), .B(creg[130]), .Z(n4818) );
  NAND U6867 ( .A(n4820), .B(n4821), .Z(x[12]) );
  NANDN U6868 ( .A(n4377), .B(creg[12]), .Z(n4820) );
  NAND U6869 ( .A(n4822), .B(n4823), .Z(x[129]) );
  NANDN U6870 ( .A(n4377), .B(creg[129]), .Z(n4822) );
  NAND U6871 ( .A(n4824), .B(n4825), .Z(x[128]) );
  NANDN U6872 ( .A(n4377), .B(creg[128]), .Z(n4824) );
  NAND U6873 ( .A(n4826), .B(n4827), .Z(x[127]) );
  NANDN U6874 ( .A(n4377), .B(creg[127]), .Z(n4826) );
  NAND U6875 ( .A(n4828), .B(n4829), .Z(x[126]) );
  NANDN U6876 ( .A(n4377), .B(creg[126]), .Z(n4828) );
  NAND U6877 ( .A(n4830), .B(n4831), .Z(x[125]) );
  NANDN U6878 ( .A(n4377), .B(creg[125]), .Z(n4830) );
  NAND U6879 ( .A(n4832), .B(n4833), .Z(x[124]) );
  NANDN U6880 ( .A(n4377), .B(creg[124]), .Z(n4832) );
  NAND U6881 ( .A(n4834), .B(n4835), .Z(x[123]) );
  NANDN U6882 ( .A(n4377), .B(creg[123]), .Z(n4834) );
  NAND U6883 ( .A(n4836), .B(n4837), .Z(x[122]) );
  NANDN U6884 ( .A(n4377), .B(creg[122]), .Z(n4836) );
  NAND U6885 ( .A(n4838), .B(n4839), .Z(x[121]) );
  NANDN U6886 ( .A(n4377), .B(creg[121]), .Z(n4838) );
  NAND U6887 ( .A(n4840), .B(n4841), .Z(x[120]) );
  NANDN U6888 ( .A(n4377), .B(creg[120]), .Z(n4840) );
  NAND U6889 ( .A(n4842), .B(n4843), .Z(x[11]) );
  NANDN U6890 ( .A(n4377), .B(creg[11]), .Z(n4842) );
  NAND U6891 ( .A(n4844), .B(n4845), .Z(x[119]) );
  NANDN U6892 ( .A(n4377), .B(creg[119]), .Z(n4844) );
  NAND U6893 ( .A(n4846), .B(n4847), .Z(x[118]) );
  NANDN U6894 ( .A(n4377), .B(creg[118]), .Z(n4846) );
  NAND U6895 ( .A(n4848), .B(n4849), .Z(x[117]) );
  NANDN U6896 ( .A(n4377), .B(creg[117]), .Z(n4848) );
  NAND U6897 ( .A(n4850), .B(n4851), .Z(x[116]) );
  NANDN U6898 ( .A(n4377), .B(creg[116]), .Z(n4850) );
  NAND U6899 ( .A(n4852), .B(n4853), .Z(x[115]) );
  NANDN U6900 ( .A(n4377), .B(creg[115]), .Z(n4852) );
  NAND U6901 ( .A(n4854), .B(n4855), .Z(x[114]) );
  NANDN U6902 ( .A(n4377), .B(creg[114]), .Z(n4854) );
  NAND U6903 ( .A(n4856), .B(n4857), .Z(x[113]) );
  NANDN U6904 ( .A(n4377), .B(creg[113]), .Z(n4856) );
  NAND U6905 ( .A(n4858), .B(n4859), .Z(x[112]) );
  NANDN U6906 ( .A(n4377), .B(creg[112]), .Z(n4858) );
  NAND U6907 ( .A(n4860), .B(n4861), .Z(x[111]) );
  NANDN U6908 ( .A(n4377), .B(creg[111]), .Z(n4860) );
  NAND U6909 ( .A(n4862), .B(n4863), .Z(x[110]) );
  NANDN U6910 ( .A(n4377), .B(creg[110]), .Z(n4862) );
  NAND U6911 ( .A(n4864), .B(n4865), .Z(x[10]) );
  NANDN U6912 ( .A(n4377), .B(creg[10]), .Z(n4864) );
  NAND U6913 ( .A(n4866), .B(n4867), .Z(x[109]) );
  NANDN U6914 ( .A(n4377), .B(creg[109]), .Z(n4866) );
  NAND U6915 ( .A(n4868), .B(n4869), .Z(x[108]) );
  NANDN U6916 ( .A(n4377), .B(creg[108]), .Z(n4868) );
  NAND U6917 ( .A(n4870), .B(n4871), .Z(x[107]) );
  NANDN U6918 ( .A(n4377), .B(creg[107]), .Z(n4870) );
  NAND U6919 ( .A(n4872), .B(n4873), .Z(x[106]) );
  NANDN U6920 ( .A(n4377), .B(creg[106]), .Z(n4872) );
  NAND U6921 ( .A(n4874), .B(n4875), .Z(x[105]) );
  NANDN U6922 ( .A(n4377), .B(creg[105]), .Z(n4874) );
  NAND U6923 ( .A(n4876), .B(n4877), .Z(x[104]) );
  NANDN U6924 ( .A(n4377), .B(creg[104]), .Z(n4876) );
  NAND U6925 ( .A(n4878), .B(n4879), .Z(x[103]) );
  NANDN U6926 ( .A(n4377), .B(creg[103]), .Z(n4878) );
  NAND U6927 ( .A(n4880), .B(n4881), .Z(x[102]) );
  NANDN U6928 ( .A(n4377), .B(creg[102]), .Z(n4880) );
  NAND U6929 ( .A(n4882), .B(n4883), .Z(x[101]) );
  NANDN U6930 ( .A(n4377), .B(creg[101]), .Z(n4882) );
  NAND U6931 ( .A(n4884), .B(n4885), .Z(x[100]) );
  NANDN U6932 ( .A(n4377), .B(creg[100]), .Z(n4884) );
  NAND U6933 ( .A(n4886), .B(n4887), .Z(x[0]) );
  NANDN U6934 ( .A(n4377), .B(creg[0]), .Z(n4886) );
  ANDN U6935 ( .B(start_reg[9]), .A(n4377), .Z(start_in[9]) );
  ANDN U6936 ( .B(start_reg[99]), .A(n4377), .Z(start_in[99]) );
  ANDN U6937 ( .B(start_reg[999]), .A(n4377), .Z(start_in[999]) );
  ANDN U6938 ( .B(start_reg[998]), .A(n4377), .Z(start_in[998]) );
  ANDN U6939 ( .B(start_reg[997]), .A(n4377), .Z(start_in[997]) );
  ANDN U6940 ( .B(start_reg[996]), .A(n4377), .Z(start_in[996]) );
  ANDN U6941 ( .B(start_reg[995]), .A(n4377), .Z(start_in[995]) );
  ANDN U6942 ( .B(start_reg[994]), .A(n4377), .Z(start_in[994]) );
  ANDN U6943 ( .B(start_reg[993]), .A(n4377), .Z(start_in[993]) );
  ANDN U6944 ( .B(start_reg[992]), .A(n4377), .Z(start_in[992]) );
  ANDN U6945 ( .B(start_reg[991]), .A(n4377), .Z(start_in[991]) );
  ANDN U6946 ( .B(start_reg[990]), .A(n4377), .Z(start_in[990]) );
  ANDN U6947 ( .B(start_reg[98]), .A(n4377), .Z(start_in[98]) );
  ANDN U6948 ( .B(start_reg[989]), .A(n4377), .Z(start_in[989]) );
  ANDN U6949 ( .B(start_reg[988]), .A(n4377), .Z(start_in[988]) );
  ANDN U6950 ( .B(start_reg[987]), .A(n4377), .Z(start_in[987]) );
  ANDN U6951 ( .B(start_reg[986]), .A(n4377), .Z(start_in[986]) );
  ANDN U6952 ( .B(start_reg[985]), .A(n4377), .Z(start_in[985]) );
  ANDN U6953 ( .B(start_reg[984]), .A(n4377), .Z(start_in[984]) );
  ANDN U6954 ( .B(start_reg[983]), .A(n4377), .Z(start_in[983]) );
  ANDN U6955 ( .B(start_reg[982]), .A(n4377), .Z(start_in[982]) );
  ANDN U6956 ( .B(start_reg[981]), .A(n4377), .Z(start_in[981]) );
  ANDN U6957 ( .B(start_reg[980]), .A(n4377), .Z(start_in[980]) );
  ANDN U6958 ( .B(start_reg[97]), .A(n4377), .Z(start_in[97]) );
  ANDN U6959 ( .B(start_reg[979]), .A(n4377), .Z(start_in[979]) );
  ANDN U6960 ( .B(start_reg[978]), .A(n4377), .Z(start_in[978]) );
  ANDN U6961 ( .B(start_reg[977]), .A(n4377), .Z(start_in[977]) );
  ANDN U6962 ( .B(start_reg[976]), .A(n4377), .Z(start_in[976]) );
  ANDN U6963 ( .B(start_reg[975]), .A(n4377), .Z(start_in[975]) );
  ANDN U6964 ( .B(start_reg[974]), .A(n4377), .Z(start_in[974]) );
  ANDN U6965 ( .B(start_reg[973]), .A(n4377), .Z(start_in[973]) );
  ANDN U6966 ( .B(start_reg[972]), .A(n4377), .Z(start_in[972]) );
  ANDN U6967 ( .B(start_reg[971]), .A(n4377), .Z(start_in[971]) );
  ANDN U6968 ( .B(start_reg[970]), .A(n4377), .Z(start_in[970]) );
  ANDN U6969 ( .B(start_reg[96]), .A(n4377), .Z(start_in[96]) );
  ANDN U6970 ( .B(start_reg[969]), .A(n4377), .Z(start_in[969]) );
  ANDN U6971 ( .B(start_reg[968]), .A(n4377), .Z(start_in[968]) );
  ANDN U6972 ( .B(start_reg[967]), .A(n4377), .Z(start_in[967]) );
  ANDN U6973 ( .B(start_reg[966]), .A(n4377), .Z(start_in[966]) );
  ANDN U6974 ( .B(start_reg[965]), .A(n4377), .Z(start_in[965]) );
  ANDN U6975 ( .B(start_reg[964]), .A(n4377), .Z(start_in[964]) );
  ANDN U6976 ( .B(start_reg[963]), .A(n4377), .Z(start_in[963]) );
  ANDN U6977 ( .B(start_reg[962]), .A(n4377), .Z(start_in[962]) );
  ANDN U6978 ( .B(start_reg[961]), .A(n4377), .Z(start_in[961]) );
  ANDN U6979 ( .B(start_reg[960]), .A(n4377), .Z(start_in[960]) );
  ANDN U6980 ( .B(start_reg[95]), .A(n4377), .Z(start_in[95]) );
  ANDN U6981 ( .B(start_reg[959]), .A(n4377), .Z(start_in[959]) );
  ANDN U6982 ( .B(start_reg[958]), .A(n4377), .Z(start_in[958]) );
  ANDN U6983 ( .B(start_reg[957]), .A(n4377), .Z(start_in[957]) );
  ANDN U6984 ( .B(start_reg[956]), .A(n4377), .Z(start_in[956]) );
  ANDN U6985 ( .B(start_reg[955]), .A(n4377), .Z(start_in[955]) );
  ANDN U6986 ( .B(start_reg[954]), .A(n4377), .Z(start_in[954]) );
  ANDN U6987 ( .B(start_reg[953]), .A(n4377), .Z(start_in[953]) );
  ANDN U6988 ( .B(start_reg[952]), .A(n4377), .Z(start_in[952]) );
  ANDN U6989 ( .B(start_reg[951]), .A(n4377), .Z(start_in[951]) );
  ANDN U6990 ( .B(start_reg[950]), .A(n4377), .Z(start_in[950]) );
  ANDN U6991 ( .B(start_reg[94]), .A(n4377), .Z(start_in[94]) );
  ANDN U6992 ( .B(start_reg[949]), .A(n4377), .Z(start_in[949]) );
  ANDN U6993 ( .B(start_reg[948]), .A(n4377), .Z(start_in[948]) );
  ANDN U6994 ( .B(start_reg[947]), .A(n4377), .Z(start_in[947]) );
  ANDN U6995 ( .B(start_reg[946]), .A(n4377), .Z(start_in[946]) );
  ANDN U6996 ( .B(start_reg[945]), .A(n4377), .Z(start_in[945]) );
  ANDN U6997 ( .B(start_reg[944]), .A(n4377), .Z(start_in[944]) );
  ANDN U6998 ( .B(start_reg[943]), .A(n4377), .Z(start_in[943]) );
  ANDN U6999 ( .B(start_reg[942]), .A(n4377), .Z(start_in[942]) );
  ANDN U7000 ( .B(start_reg[941]), .A(n4377), .Z(start_in[941]) );
  ANDN U7001 ( .B(start_reg[940]), .A(n4377), .Z(start_in[940]) );
  ANDN U7002 ( .B(start_reg[93]), .A(n4377), .Z(start_in[93]) );
  ANDN U7003 ( .B(start_reg[939]), .A(n4377), .Z(start_in[939]) );
  ANDN U7004 ( .B(start_reg[938]), .A(n4377), .Z(start_in[938]) );
  ANDN U7005 ( .B(start_reg[937]), .A(n4377), .Z(start_in[937]) );
  ANDN U7006 ( .B(start_reg[936]), .A(n4377), .Z(start_in[936]) );
  ANDN U7007 ( .B(start_reg[935]), .A(n4377), .Z(start_in[935]) );
  ANDN U7008 ( .B(start_reg[934]), .A(n4377), .Z(start_in[934]) );
  ANDN U7009 ( .B(start_reg[933]), .A(n4377), .Z(start_in[933]) );
  ANDN U7010 ( .B(start_reg[932]), .A(n4377), .Z(start_in[932]) );
  ANDN U7011 ( .B(start_reg[931]), .A(n4377), .Z(start_in[931]) );
  ANDN U7012 ( .B(start_reg[930]), .A(n4377), .Z(start_in[930]) );
  ANDN U7013 ( .B(start_reg[92]), .A(n4377), .Z(start_in[92]) );
  ANDN U7014 ( .B(start_reg[929]), .A(n4377), .Z(start_in[929]) );
  ANDN U7015 ( .B(start_reg[928]), .A(n4377), .Z(start_in[928]) );
  ANDN U7016 ( .B(start_reg[927]), .A(n4377), .Z(start_in[927]) );
  ANDN U7017 ( .B(start_reg[926]), .A(n4377), .Z(start_in[926]) );
  ANDN U7018 ( .B(start_reg[925]), .A(n4377), .Z(start_in[925]) );
  ANDN U7019 ( .B(start_reg[924]), .A(n4377), .Z(start_in[924]) );
  ANDN U7020 ( .B(start_reg[923]), .A(n4377), .Z(start_in[923]) );
  ANDN U7021 ( .B(start_reg[922]), .A(n4377), .Z(start_in[922]) );
  ANDN U7022 ( .B(start_reg[921]), .A(n4377), .Z(start_in[921]) );
  ANDN U7023 ( .B(start_reg[920]), .A(n4377), .Z(start_in[920]) );
  ANDN U7024 ( .B(start_reg[91]), .A(n4377), .Z(start_in[91]) );
  ANDN U7025 ( .B(start_reg[919]), .A(n4377), .Z(start_in[919]) );
  ANDN U7026 ( .B(start_reg[918]), .A(n4377), .Z(start_in[918]) );
  ANDN U7027 ( .B(start_reg[917]), .A(n4377), .Z(start_in[917]) );
  ANDN U7028 ( .B(start_reg[916]), .A(n4377), .Z(start_in[916]) );
  ANDN U7029 ( .B(start_reg[915]), .A(n4377), .Z(start_in[915]) );
  ANDN U7030 ( .B(start_reg[914]), .A(n4377), .Z(start_in[914]) );
  ANDN U7031 ( .B(start_reg[913]), .A(n4377), .Z(start_in[913]) );
  ANDN U7032 ( .B(start_reg[912]), .A(n4377), .Z(start_in[912]) );
  ANDN U7033 ( .B(start_reg[911]), .A(n4377), .Z(start_in[911]) );
  ANDN U7034 ( .B(start_reg[910]), .A(n4377), .Z(start_in[910]) );
  ANDN U7035 ( .B(start_reg[90]), .A(n4377), .Z(start_in[90]) );
  ANDN U7036 ( .B(start_reg[909]), .A(n4377), .Z(start_in[909]) );
  ANDN U7037 ( .B(start_reg[908]), .A(n4377), .Z(start_in[908]) );
  ANDN U7038 ( .B(start_reg[907]), .A(n4377), .Z(start_in[907]) );
  ANDN U7039 ( .B(start_reg[906]), .A(n4377), .Z(start_in[906]) );
  ANDN U7040 ( .B(start_reg[905]), .A(n4377), .Z(start_in[905]) );
  ANDN U7041 ( .B(start_reg[904]), .A(n4377), .Z(start_in[904]) );
  ANDN U7042 ( .B(start_reg[903]), .A(n4377), .Z(start_in[903]) );
  ANDN U7043 ( .B(start_reg[902]), .A(n4377), .Z(start_in[902]) );
  ANDN U7044 ( .B(start_reg[901]), .A(n4377), .Z(start_in[901]) );
  ANDN U7045 ( .B(start_reg[900]), .A(n4377), .Z(start_in[900]) );
  ANDN U7046 ( .B(start_reg[8]), .A(n4377), .Z(start_in[8]) );
  ANDN U7047 ( .B(start_reg[89]), .A(n4377), .Z(start_in[89]) );
  ANDN U7048 ( .B(start_reg[899]), .A(n4377), .Z(start_in[899]) );
  ANDN U7049 ( .B(start_reg[898]), .A(n4377), .Z(start_in[898]) );
  ANDN U7050 ( .B(start_reg[897]), .A(n4377), .Z(start_in[897]) );
  ANDN U7051 ( .B(start_reg[896]), .A(n4377), .Z(start_in[896]) );
  ANDN U7052 ( .B(start_reg[895]), .A(n4377), .Z(start_in[895]) );
  ANDN U7053 ( .B(start_reg[894]), .A(n4377), .Z(start_in[894]) );
  ANDN U7054 ( .B(start_reg[893]), .A(n4377), .Z(start_in[893]) );
  ANDN U7055 ( .B(start_reg[892]), .A(n4377), .Z(start_in[892]) );
  ANDN U7056 ( .B(start_reg[891]), .A(n4377), .Z(start_in[891]) );
  ANDN U7057 ( .B(start_reg[890]), .A(n4377), .Z(start_in[890]) );
  ANDN U7058 ( .B(start_reg[88]), .A(n4377), .Z(start_in[88]) );
  ANDN U7059 ( .B(start_reg[889]), .A(n4377), .Z(start_in[889]) );
  ANDN U7060 ( .B(start_reg[888]), .A(n4377), .Z(start_in[888]) );
  ANDN U7061 ( .B(start_reg[887]), .A(n4377), .Z(start_in[887]) );
  ANDN U7062 ( .B(start_reg[886]), .A(n4377), .Z(start_in[886]) );
  ANDN U7063 ( .B(start_reg[885]), .A(n4377), .Z(start_in[885]) );
  ANDN U7064 ( .B(start_reg[884]), .A(n4377), .Z(start_in[884]) );
  ANDN U7065 ( .B(start_reg[883]), .A(n4377), .Z(start_in[883]) );
  ANDN U7066 ( .B(start_reg[882]), .A(n4377), .Z(start_in[882]) );
  ANDN U7067 ( .B(start_reg[881]), .A(n4377), .Z(start_in[881]) );
  ANDN U7068 ( .B(start_reg[880]), .A(n4377), .Z(start_in[880]) );
  ANDN U7069 ( .B(start_reg[87]), .A(n4377), .Z(start_in[87]) );
  ANDN U7070 ( .B(start_reg[879]), .A(n4377), .Z(start_in[879]) );
  ANDN U7071 ( .B(start_reg[878]), .A(n4377), .Z(start_in[878]) );
  ANDN U7072 ( .B(start_reg[877]), .A(n4377), .Z(start_in[877]) );
  ANDN U7073 ( .B(start_reg[876]), .A(n4377), .Z(start_in[876]) );
  ANDN U7074 ( .B(start_reg[875]), .A(n4377), .Z(start_in[875]) );
  ANDN U7075 ( .B(start_reg[874]), .A(n4377), .Z(start_in[874]) );
  ANDN U7076 ( .B(start_reg[873]), .A(n4377), .Z(start_in[873]) );
  ANDN U7077 ( .B(start_reg[872]), .A(n4377), .Z(start_in[872]) );
  ANDN U7078 ( .B(start_reg[871]), .A(n4377), .Z(start_in[871]) );
  ANDN U7079 ( .B(start_reg[870]), .A(n4377), .Z(start_in[870]) );
  ANDN U7080 ( .B(start_reg[86]), .A(n4377), .Z(start_in[86]) );
  ANDN U7081 ( .B(start_reg[869]), .A(n4377), .Z(start_in[869]) );
  ANDN U7082 ( .B(start_reg[868]), .A(n4377), .Z(start_in[868]) );
  ANDN U7083 ( .B(start_reg[867]), .A(n4377), .Z(start_in[867]) );
  ANDN U7084 ( .B(start_reg[866]), .A(n4377), .Z(start_in[866]) );
  ANDN U7085 ( .B(start_reg[865]), .A(n4377), .Z(start_in[865]) );
  ANDN U7086 ( .B(start_reg[864]), .A(n4377), .Z(start_in[864]) );
  ANDN U7087 ( .B(start_reg[863]), .A(n4377), .Z(start_in[863]) );
  ANDN U7088 ( .B(start_reg[862]), .A(n4377), .Z(start_in[862]) );
  ANDN U7089 ( .B(start_reg[861]), .A(n4377), .Z(start_in[861]) );
  ANDN U7090 ( .B(start_reg[860]), .A(n4377), .Z(start_in[860]) );
  ANDN U7091 ( .B(start_reg[85]), .A(n4377), .Z(start_in[85]) );
  ANDN U7092 ( .B(start_reg[859]), .A(n4377), .Z(start_in[859]) );
  ANDN U7093 ( .B(start_reg[858]), .A(n4377), .Z(start_in[858]) );
  ANDN U7094 ( .B(start_reg[857]), .A(n4377), .Z(start_in[857]) );
  ANDN U7095 ( .B(start_reg[856]), .A(n4377), .Z(start_in[856]) );
  ANDN U7096 ( .B(start_reg[855]), .A(n4377), .Z(start_in[855]) );
  ANDN U7097 ( .B(start_reg[854]), .A(n4377), .Z(start_in[854]) );
  ANDN U7098 ( .B(start_reg[853]), .A(n4377), .Z(start_in[853]) );
  ANDN U7099 ( .B(start_reg[852]), .A(n4377), .Z(start_in[852]) );
  ANDN U7100 ( .B(start_reg[851]), .A(n4377), .Z(start_in[851]) );
  ANDN U7101 ( .B(start_reg[850]), .A(n4377), .Z(start_in[850]) );
  ANDN U7102 ( .B(start_reg[84]), .A(n4377), .Z(start_in[84]) );
  ANDN U7103 ( .B(start_reg[849]), .A(n4377), .Z(start_in[849]) );
  ANDN U7104 ( .B(start_reg[848]), .A(n4377), .Z(start_in[848]) );
  ANDN U7105 ( .B(start_reg[847]), .A(n4377), .Z(start_in[847]) );
  ANDN U7106 ( .B(start_reg[846]), .A(n4377), .Z(start_in[846]) );
  ANDN U7107 ( .B(start_reg[845]), .A(n4377), .Z(start_in[845]) );
  ANDN U7108 ( .B(start_reg[844]), .A(n4377), .Z(start_in[844]) );
  ANDN U7109 ( .B(start_reg[843]), .A(n4377), .Z(start_in[843]) );
  ANDN U7110 ( .B(start_reg[842]), .A(n4377), .Z(start_in[842]) );
  ANDN U7111 ( .B(start_reg[841]), .A(n4377), .Z(start_in[841]) );
  ANDN U7112 ( .B(start_reg[840]), .A(n4377), .Z(start_in[840]) );
  ANDN U7113 ( .B(start_reg[83]), .A(n4377), .Z(start_in[83]) );
  ANDN U7114 ( .B(start_reg[839]), .A(n4377), .Z(start_in[839]) );
  ANDN U7115 ( .B(start_reg[838]), .A(n4377), .Z(start_in[838]) );
  ANDN U7116 ( .B(start_reg[837]), .A(n4377), .Z(start_in[837]) );
  ANDN U7117 ( .B(start_reg[836]), .A(n4377), .Z(start_in[836]) );
  ANDN U7118 ( .B(start_reg[835]), .A(n4377), .Z(start_in[835]) );
  ANDN U7119 ( .B(start_reg[834]), .A(n4377), .Z(start_in[834]) );
  ANDN U7120 ( .B(start_reg[833]), .A(n4377), .Z(start_in[833]) );
  ANDN U7121 ( .B(start_reg[832]), .A(n4377), .Z(start_in[832]) );
  ANDN U7122 ( .B(start_reg[831]), .A(n4377), .Z(start_in[831]) );
  ANDN U7123 ( .B(start_reg[830]), .A(n4377), .Z(start_in[830]) );
  ANDN U7124 ( .B(start_reg[82]), .A(n4377), .Z(start_in[82]) );
  ANDN U7125 ( .B(start_reg[829]), .A(n4377), .Z(start_in[829]) );
  ANDN U7126 ( .B(start_reg[828]), .A(n4377), .Z(start_in[828]) );
  ANDN U7127 ( .B(start_reg[827]), .A(n4377), .Z(start_in[827]) );
  ANDN U7128 ( .B(start_reg[826]), .A(n4377), .Z(start_in[826]) );
  ANDN U7129 ( .B(start_reg[825]), .A(n4377), .Z(start_in[825]) );
  ANDN U7130 ( .B(start_reg[824]), .A(n4377), .Z(start_in[824]) );
  ANDN U7131 ( .B(start_reg[823]), .A(n4377), .Z(start_in[823]) );
  ANDN U7132 ( .B(start_reg[822]), .A(n4377), .Z(start_in[822]) );
  ANDN U7133 ( .B(start_reg[821]), .A(n4377), .Z(start_in[821]) );
  ANDN U7134 ( .B(start_reg[820]), .A(n4377), .Z(start_in[820]) );
  ANDN U7135 ( .B(start_reg[81]), .A(n4377), .Z(start_in[81]) );
  ANDN U7136 ( .B(start_reg[819]), .A(n4377), .Z(start_in[819]) );
  ANDN U7137 ( .B(start_reg[818]), .A(n4377), .Z(start_in[818]) );
  ANDN U7138 ( .B(start_reg[817]), .A(n4377), .Z(start_in[817]) );
  ANDN U7139 ( .B(start_reg[816]), .A(n4377), .Z(start_in[816]) );
  ANDN U7140 ( .B(start_reg[815]), .A(n4377), .Z(start_in[815]) );
  ANDN U7141 ( .B(start_reg[814]), .A(n4377), .Z(start_in[814]) );
  ANDN U7142 ( .B(start_reg[813]), .A(n4377), .Z(start_in[813]) );
  ANDN U7143 ( .B(start_reg[812]), .A(n4377), .Z(start_in[812]) );
  ANDN U7144 ( .B(start_reg[811]), .A(n4377), .Z(start_in[811]) );
  ANDN U7145 ( .B(start_reg[810]), .A(n4377), .Z(start_in[810]) );
  ANDN U7146 ( .B(start_reg[80]), .A(n4377), .Z(start_in[80]) );
  ANDN U7147 ( .B(start_reg[809]), .A(n4377), .Z(start_in[809]) );
  ANDN U7148 ( .B(start_reg[808]), .A(n4377), .Z(start_in[808]) );
  ANDN U7149 ( .B(start_reg[807]), .A(n4377), .Z(start_in[807]) );
  ANDN U7150 ( .B(start_reg[806]), .A(n4377), .Z(start_in[806]) );
  ANDN U7151 ( .B(start_reg[805]), .A(n4377), .Z(start_in[805]) );
  ANDN U7152 ( .B(start_reg[804]), .A(n4377), .Z(start_in[804]) );
  ANDN U7153 ( .B(start_reg[803]), .A(n4377), .Z(start_in[803]) );
  ANDN U7154 ( .B(start_reg[802]), .A(n4377), .Z(start_in[802]) );
  ANDN U7155 ( .B(start_reg[801]), .A(n4377), .Z(start_in[801]) );
  ANDN U7156 ( .B(start_reg[800]), .A(n4377), .Z(start_in[800]) );
  ANDN U7157 ( .B(start_reg[7]), .A(n4377), .Z(start_in[7]) );
  ANDN U7158 ( .B(start_reg[79]), .A(n4377), .Z(start_in[79]) );
  ANDN U7159 ( .B(start_reg[799]), .A(n4377), .Z(start_in[799]) );
  ANDN U7160 ( .B(start_reg[798]), .A(n4377), .Z(start_in[798]) );
  ANDN U7161 ( .B(start_reg[797]), .A(n4377), .Z(start_in[797]) );
  ANDN U7162 ( .B(start_reg[796]), .A(n4377), .Z(start_in[796]) );
  ANDN U7163 ( .B(start_reg[795]), .A(n4377), .Z(start_in[795]) );
  ANDN U7164 ( .B(start_reg[794]), .A(n4377), .Z(start_in[794]) );
  ANDN U7165 ( .B(start_reg[793]), .A(n4377), .Z(start_in[793]) );
  ANDN U7166 ( .B(start_reg[792]), .A(n4377), .Z(start_in[792]) );
  ANDN U7167 ( .B(start_reg[791]), .A(n4377), .Z(start_in[791]) );
  ANDN U7168 ( .B(start_reg[790]), .A(n4377), .Z(start_in[790]) );
  ANDN U7169 ( .B(start_reg[78]), .A(n4377), .Z(start_in[78]) );
  ANDN U7170 ( .B(start_reg[789]), .A(n4377), .Z(start_in[789]) );
  ANDN U7171 ( .B(start_reg[788]), .A(n4377), .Z(start_in[788]) );
  ANDN U7172 ( .B(start_reg[787]), .A(n4377), .Z(start_in[787]) );
  ANDN U7173 ( .B(start_reg[786]), .A(n4377), .Z(start_in[786]) );
  ANDN U7174 ( .B(start_reg[785]), .A(n4377), .Z(start_in[785]) );
  ANDN U7175 ( .B(start_reg[784]), .A(n4377), .Z(start_in[784]) );
  ANDN U7176 ( .B(start_reg[783]), .A(n4377), .Z(start_in[783]) );
  ANDN U7177 ( .B(start_reg[782]), .A(n4377), .Z(start_in[782]) );
  ANDN U7178 ( .B(start_reg[781]), .A(n4377), .Z(start_in[781]) );
  ANDN U7179 ( .B(start_reg[780]), .A(n4377), .Z(start_in[780]) );
  ANDN U7180 ( .B(start_reg[77]), .A(n4377), .Z(start_in[77]) );
  ANDN U7181 ( .B(start_reg[779]), .A(n4377), .Z(start_in[779]) );
  ANDN U7182 ( .B(start_reg[778]), .A(n4377), .Z(start_in[778]) );
  ANDN U7183 ( .B(start_reg[777]), .A(n4377), .Z(start_in[777]) );
  ANDN U7184 ( .B(start_reg[776]), .A(n4377), .Z(start_in[776]) );
  ANDN U7185 ( .B(start_reg[775]), .A(n4377), .Z(start_in[775]) );
  ANDN U7186 ( .B(start_reg[774]), .A(n4377), .Z(start_in[774]) );
  ANDN U7187 ( .B(start_reg[773]), .A(n4377), .Z(start_in[773]) );
  ANDN U7188 ( .B(start_reg[772]), .A(n4377), .Z(start_in[772]) );
  ANDN U7189 ( .B(start_reg[771]), .A(n4377), .Z(start_in[771]) );
  ANDN U7190 ( .B(start_reg[770]), .A(n4377), .Z(start_in[770]) );
  ANDN U7191 ( .B(start_reg[76]), .A(n4377), .Z(start_in[76]) );
  ANDN U7192 ( .B(start_reg[769]), .A(n4377), .Z(start_in[769]) );
  ANDN U7193 ( .B(start_reg[768]), .A(n4377), .Z(start_in[768]) );
  ANDN U7194 ( .B(start_reg[767]), .A(n4377), .Z(start_in[767]) );
  ANDN U7195 ( .B(start_reg[766]), .A(n4377), .Z(start_in[766]) );
  ANDN U7196 ( .B(start_reg[765]), .A(n4377), .Z(start_in[765]) );
  ANDN U7197 ( .B(start_reg[764]), .A(n4377), .Z(start_in[764]) );
  ANDN U7198 ( .B(start_reg[763]), .A(n4377), .Z(start_in[763]) );
  ANDN U7199 ( .B(start_reg[762]), .A(n4377), .Z(start_in[762]) );
  ANDN U7200 ( .B(start_reg[761]), .A(n4377), .Z(start_in[761]) );
  ANDN U7201 ( .B(start_reg[760]), .A(n4377), .Z(start_in[760]) );
  ANDN U7202 ( .B(start_reg[75]), .A(n4377), .Z(start_in[75]) );
  ANDN U7203 ( .B(start_reg[759]), .A(n4377), .Z(start_in[759]) );
  ANDN U7204 ( .B(start_reg[758]), .A(n4377), .Z(start_in[758]) );
  ANDN U7205 ( .B(start_reg[757]), .A(n4377), .Z(start_in[757]) );
  ANDN U7206 ( .B(start_reg[756]), .A(n4377), .Z(start_in[756]) );
  ANDN U7207 ( .B(start_reg[755]), .A(n4377), .Z(start_in[755]) );
  ANDN U7208 ( .B(start_reg[754]), .A(n4377), .Z(start_in[754]) );
  ANDN U7209 ( .B(start_reg[753]), .A(n4377), .Z(start_in[753]) );
  ANDN U7210 ( .B(start_reg[752]), .A(n4377), .Z(start_in[752]) );
  ANDN U7211 ( .B(start_reg[751]), .A(n4377), .Z(start_in[751]) );
  ANDN U7212 ( .B(start_reg[750]), .A(n4377), .Z(start_in[750]) );
  ANDN U7213 ( .B(start_reg[74]), .A(n4377), .Z(start_in[74]) );
  ANDN U7214 ( .B(start_reg[749]), .A(n4377), .Z(start_in[749]) );
  ANDN U7215 ( .B(start_reg[748]), .A(n4377), .Z(start_in[748]) );
  ANDN U7216 ( .B(start_reg[747]), .A(n4377), .Z(start_in[747]) );
  ANDN U7217 ( .B(start_reg[746]), .A(n4377), .Z(start_in[746]) );
  ANDN U7218 ( .B(start_reg[745]), .A(n4377), .Z(start_in[745]) );
  ANDN U7219 ( .B(start_reg[744]), .A(n4377), .Z(start_in[744]) );
  ANDN U7220 ( .B(start_reg[743]), .A(n4377), .Z(start_in[743]) );
  ANDN U7221 ( .B(start_reg[742]), .A(n4377), .Z(start_in[742]) );
  ANDN U7222 ( .B(start_reg[741]), .A(n4377), .Z(start_in[741]) );
  ANDN U7223 ( .B(start_reg[740]), .A(n4377), .Z(start_in[740]) );
  ANDN U7224 ( .B(start_reg[73]), .A(n4377), .Z(start_in[73]) );
  ANDN U7225 ( .B(start_reg[739]), .A(n4377), .Z(start_in[739]) );
  ANDN U7226 ( .B(start_reg[738]), .A(n4377), .Z(start_in[738]) );
  ANDN U7227 ( .B(start_reg[737]), .A(n4377), .Z(start_in[737]) );
  ANDN U7228 ( .B(start_reg[736]), .A(n4377), .Z(start_in[736]) );
  ANDN U7229 ( .B(start_reg[735]), .A(n4377), .Z(start_in[735]) );
  ANDN U7230 ( .B(start_reg[734]), .A(n4377), .Z(start_in[734]) );
  ANDN U7231 ( .B(start_reg[733]), .A(n4377), .Z(start_in[733]) );
  ANDN U7232 ( .B(start_reg[732]), .A(n4377), .Z(start_in[732]) );
  ANDN U7233 ( .B(start_reg[731]), .A(n4377), .Z(start_in[731]) );
  ANDN U7234 ( .B(start_reg[730]), .A(n4377), .Z(start_in[730]) );
  ANDN U7235 ( .B(start_reg[72]), .A(n4377), .Z(start_in[72]) );
  ANDN U7236 ( .B(start_reg[729]), .A(n4377), .Z(start_in[729]) );
  ANDN U7237 ( .B(start_reg[728]), .A(n4377), .Z(start_in[728]) );
  ANDN U7238 ( .B(start_reg[727]), .A(n4377), .Z(start_in[727]) );
  ANDN U7239 ( .B(start_reg[726]), .A(n4377), .Z(start_in[726]) );
  ANDN U7240 ( .B(start_reg[725]), .A(n4377), .Z(start_in[725]) );
  ANDN U7241 ( .B(start_reg[724]), .A(n4377), .Z(start_in[724]) );
  ANDN U7242 ( .B(start_reg[723]), .A(n4377), .Z(start_in[723]) );
  ANDN U7243 ( .B(start_reg[722]), .A(n4377), .Z(start_in[722]) );
  ANDN U7244 ( .B(start_reg[721]), .A(n4377), .Z(start_in[721]) );
  ANDN U7245 ( .B(start_reg[720]), .A(n4377), .Z(start_in[720]) );
  ANDN U7246 ( .B(start_reg[71]), .A(n4377), .Z(start_in[71]) );
  ANDN U7247 ( .B(start_reg[719]), .A(n4377), .Z(start_in[719]) );
  ANDN U7248 ( .B(start_reg[718]), .A(n4377), .Z(start_in[718]) );
  ANDN U7249 ( .B(start_reg[717]), .A(n4377), .Z(start_in[717]) );
  ANDN U7250 ( .B(start_reg[716]), .A(n4377), .Z(start_in[716]) );
  ANDN U7251 ( .B(start_reg[715]), .A(n4377), .Z(start_in[715]) );
  ANDN U7252 ( .B(start_reg[714]), .A(n4377), .Z(start_in[714]) );
  ANDN U7253 ( .B(start_reg[713]), .A(n4377), .Z(start_in[713]) );
  ANDN U7254 ( .B(start_reg[712]), .A(n4377), .Z(start_in[712]) );
  ANDN U7255 ( .B(start_reg[711]), .A(n4377), .Z(start_in[711]) );
  ANDN U7256 ( .B(start_reg[710]), .A(n4377), .Z(start_in[710]) );
  ANDN U7257 ( .B(start_reg[70]), .A(n4377), .Z(start_in[70]) );
  ANDN U7258 ( .B(start_reg[709]), .A(n4377), .Z(start_in[709]) );
  ANDN U7259 ( .B(start_reg[708]), .A(n4377), .Z(start_in[708]) );
  ANDN U7260 ( .B(start_reg[707]), .A(n4377), .Z(start_in[707]) );
  ANDN U7261 ( .B(start_reg[706]), .A(n4377), .Z(start_in[706]) );
  ANDN U7262 ( .B(start_reg[705]), .A(n4377), .Z(start_in[705]) );
  ANDN U7263 ( .B(start_reg[704]), .A(n4377), .Z(start_in[704]) );
  ANDN U7264 ( .B(start_reg[703]), .A(n4377), .Z(start_in[703]) );
  ANDN U7265 ( .B(start_reg[702]), .A(n4377), .Z(start_in[702]) );
  ANDN U7266 ( .B(start_reg[701]), .A(n4377), .Z(start_in[701]) );
  ANDN U7267 ( .B(start_reg[700]), .A(n4377), .Z(start_in[700]) );
  ANDN U7268 ( .B(start_reg[6]), .A(n4377), .Z(start_in[6]) );
  ANDN U7269 ( .B(start_reg[69]), .A(n4377), .Z(start_in[69]) );
  ANDN U7270 ( .B(start_reg[699]), .A(n4377), .Z(start_in[699]) );
  ANDN U7271 ( .B(start_reg[698]), .A(n4377), .Z(start_in[698]) );
  ANDN U7272 ( .B(start_reg[697]), .A(n4377), .Z(start_in[697]) );
  ANDN U7273 ( .B(start_reg[696]), .A(n4377), .Z(start_in[696]) );
  ANDN U7274 ( .B(start_reg[695]), .A(n4377), .Z(start_in[695]) );
  ANDN U7275 ( .B(start_reg[694]), .A(n4377), .Z(start_in[694]) );
  ANDN U7276 ( .B(start_reg[693]), .A(n4377), .Z(start_in[693]) );
  ANDN U7277 ( .B(start_reg[692]), .A(n4377), .Z(start_in[692]) );
  ANDN U7278 ( .B(start_reg[691]), .A(n4377), .Z(start_in[691]) );
  ANDN U7279 ( .B(start_reg[690]), .A(n4377), .Z(start_in[690]) );
  ANDN U7280 ( .B(start_reg[68]), .A(n4377), .Z(start_in[68]) );
  ANDN U7281 ( .B(start_reg[689]), .A(n4377), .Z(start_in[689]) );
  ANDN U7282 ( .B(start_reg[688]), .A(n4377), .Z(start_in[688]) );
  ANDN U7283 ( .B(start_reg[687]), .A(n4377), .Z(start_in[687]) );
  ANDN U7284 ( .B(start_reg[686]), .A(n4377), .Z(start_in[686]) );
  ANDN U7285 ( .B(start_reg[685]), .A(n4377), .Z(start_in[685]) );
  ANDN U7286 ( .B(start_reg[684]), .A(n4377), .Z(start_in[684]) );
  ANDN U7287 ( .B(start_reg[683]), .A(n4377), .Z(start_in[683]) );
  ANDN U7288 ( .B(start_reg[682]), .A(n4377), .Z(start_in[682]) );
  ANDN U7289 ( .B(start_reg[681]), .A(n4377), .Z(start_in[681]) );
  ANDN U7290 ( .B(start_reg[680]), .A(n4377), .Z(start_in[680]) );
  ANDN U7291 ( .B(start_reg[67]), .A(n4377), .Z(start_in[67]) );
  ANDN U7292 ( .B(start_reg[679]), .A(n4377), .Z(start_in[679]) );
  ANDN U7293 ( .B(start_reg[678]), .A(n4377), .Z(start_in[678]) );
  ANDN U7294 ( .B(start_reg[677]), .A(n4377), .Z(start_in[677]) );
  ANDN U7295 ( .B(start_reg[676]), .A(n4377), .Z(start_in[676]) );
  ANDN U7296 ( .B(start_reg[675]), .A(n4377), .Z(start_in[675]) );
  ANDN U7297 ( .B(start_reg[674]), .A(n4377), .Z(start_in[674]) );
  ANDN U7298 ( .B(start_reg[673]), .A(n4377), .Z(start_in[673]) );
  ANDN U7299 ( .B(start_reg[672]), .A(n4377), .Z(start_in[672]) );
  ANDN U7300 ( .B(start_reg[671]), .A(n4377), .Z(start_in[671]) );
  ANDN U7301 ( .B(start_reg[670]), .A(n4377), .Z(start_in[670]) );
  ANDN U7302 ( .B(start_reg[66]), .A(n4377), .Z(start_in[66]) );
  ANDN U7303 ( .B(start_reg[669]), .A(n4377), .Z(start_in[669]) );
  ANDN U7304 ( .B(start_reg[668]), .A(n4377), .Z(start_in[668]) );
  ANDN U7305 ( .B(start_reg[667]), .A(n4377), .Z(start_in[667]) );
  ANDN U7306 ( .B(start_reg[666]), .A(n4377), .Z(start_in[666]) );
  ANDN U7307 ( .B(start_reg[665]), .A(n4377), .Z(start_in[665]) );
  ANDN U7308 ( .B(start_reg[664]), .A(n4377), .Z(start_in[664]) );
  ANDN U7309 ( .B(start_reg[663]), .A(n4377), .Z(start_in[663]) );
  ANDN U7310 ( .B(start_reg[662]), .A(n4377), .Z(start_in[662]) );
  ANDN U7311 ( .B(start_reg[661]), .A(n4377), .Z(start_in[661]) );
  ANDN U7312 ( .B(start_reg[660]), .A(n4377), .Z(start_in[660]) );
  ANDN U7313 ( .B(start_reg[65]), .A(n4377), .Z(start_in[65]) );
  ANDN U7314 ( .B(start_reg[659]), .A(n4377), .Z(start_in[659]) );
  ANDN U7315 ( .B(start_reg[658]), .A(n4377), .Z(start_in[658]) );
  ANDN U7316 ( .B(start_reg[657]), .A(n4377), .Z(start_in[657]) );
  ANDN U7317 ( .B(start_reg[656]), .A(n4377), .Z(start_in[656]) );
  ANDN U7318 ( .B(start_reg[655]), .A(n4377), .Z(start_in[655]) );
  ANDN U7319 ( .B(start_reg[654]), .A(n4377), .Z(start_in[654]) );
  ANDN U7320 ( .B(start_reg[653]), .A(n4377), .Z(start_in[653]) );
  ANDN U7321 ( .B(start_reg[652]), .A(n4377), .Z(start_in[652]) );
  ANDN U7322 ( .B(start_reg[651]), .A(n4377), .Z(start_in[651]) );
  ANDN U7323 ( .B(start_reg[650]), .A(n4377), .Z(start_in[650]) );
  ANDN U7324 ( .B(start_reg[64]), .A(n4377), .Z(start_in[64]) );
  ANDN U7325 ( .B(start_reg[649]), .A(n4377), .Z(start_in[649]) );
  ANDN U7326 ( .B(start_reg[648]), .A(n4377), .Z(start_in[648]) );
  ANDN U7327 ( .B(start_reg[647]), .A(n4377), .Z(start_in[647]) );
  ANDN U7328 ( .B(start_reg[646]), .A(n4377), .Z(start_in[646]) );
  ANDN U7329 ( .B(start_reg[645]), .A(n4377), .Z(start_in[645]) );
  ANDN U7330 ( .B(start_reg[644]), .A(n4377), .Z(start_in[644]) );
  ANDN U7331 ( .B(start_reg[643]), .A(n4377), .Z(start_in[643]) );
  ANDN U7332 ( .B(start_reg[642]), .A(n4377), .Z(start_in[642]) );
  ANDN U7333 ( .B(start_reg[641]), .A(n4377), .Z(start_in[641]) );
  ANDN U7334 ( .B(start_reg[640]), .A(n4377), .Z(start_in[640]) );
  ANDN U7335 ( .B(start_reg[63]), .A(n4377), .Z(start_in[63]) );
  ANDN U7336 ( .B(start_reg[639]), .A(n4377), .Z(start_in[639]) );
  ANDN U7337 ( .B(start_reg[638]), .A(n4377), .Z(start_in[638]) );
  ANDN U7338 ( .B(start_reg[637]), .A(n4377), .Z(start_in[637]) );
  ANDN U7339 ( .B(start_reg[636]), .A(n4377), .Z(start_in[636]) );
  ANDN U7340 ( .B(start_reg[635]), .A(n4377), .Z(start_in[635]) );
  ANDN U7341 ( .B(start_reg[634]), .A(n4377), .Z(start_in[634]) );
  ANDN U7342 ( .B(start_reg[633]), .A(n4377), .Z(start_in[633]) );
  ANDN U7343 ( .B(start_reg[632]), .A(n4377), .Z(start_in[632]) );
  ANDN U7344 ( .B(start_reg[631]), .A(n4377), .Z(start_in[631]) );
  ANDN U7345 ( .B(start_reg[630]), .A(n4377), .Z(start_in[630]) );
  ANDN U7346 ( .B(start_reg[62]), .A(n4377), .Z(start_in[62]) );
  ANDN U7347 ( .B(start_reg[629]), .A(n4377), .Z(start_in[629]) );
  ANDN U7348 ( .B(start_reg[628]), .A(n4377), .Z(start_in[628]) );
  ANDN U7349 ( .B(start_reg[627]), .A(n4377), .Z(start_in[627]) );
  ANDN U7350 ( .B(start_reg[626]), .A(n4377), .Z(start_in[626]) );
  ANDN U7351 ( .B(start_reg[625]), .A(n4377), .Z(start_in[625]) );
  ANDN U7352 ( .B(start_reg[624]), .A(n4377), .Z(start_in[624]) );
  ANDN U7353 ( .B(start_reg[623]), .A(n4377), .Z(start_in[623]) );
  ANDN U7354 ( .B(start_reg[622]), .A(n4377), .Z(start_in[622]) );
  ANDN U7355 ( .B(start_reg[621]), .A(n4377), .Z(start_in[621]) );
  ANDN U7356 ( .B(start_reg[620]), .A(n4377), .Z(start_in[620]) );
  ANDN U7357 ( .B(start_reg[61]), .A(n4377), .Z(start_in[61]) );
  ANDN U7358 ( .B(start_reg[619]), .A(n4377), .Z(start_in[619]) );
  ANDN U7359 ( .B(start_reg[618]), .A(n4377), .Z(start_in[618]) );
  ANDN U7360 ( .B(start_reg[617]), .A(n4377), .Z(start_in[617]) );
  ANDN U7361 ( .B(start_reg[616]), .A(n4377), .Z(start_in[616]) );
  ANDN U7362 ( .B(start_reg[615]), .A(n4377), .Z(start_in[615]) );
  ANDN U7363 ( .B(start_reg[614]), .A(n4377), .Z(start_in[614]) );
  ANDN U7364 ( .B(start_reg[613]), .A(n4377), .Z(start_in[613]) );
  ANDN U7365 ( .B(start_reg[612]), .A(n4377), .Z(start_in[612]) );
  ANDN U7366 ( .B(start_reg[611]), .A(n4377), .Z(start_in[611]) );
  ANDN U7367 ( .B(start_reg[610]), .A(n4377), .Z(start_in[610]) );
  ANDN U7368 ( .B(start_reg[60]), .A(n4377), .Z(start_in[60]) );
  ANDN U7369 ( .B(start_reg[609]), .A(n4377), .Z(start_in[609]) );
  ANDN U7370 ( .B(start_reg[608]), .A(n4377), .Z(start_in[608]) );
  ANDN U7371 ( .B(start_reg[607]), .A(n4377), .Z(start_in[607]) );
  ANDN U7372 ( .B(start_reg[606]), .A(n4377), .Z(start_in[606]) );
  ANDN U7373 ( .B(start_reg[605]), .A(n4377), .Z(start_in[605]) );
  ANDN U7374 ( .B(start_reg[604]), .A(n4377), .Z(start_in[604]) );
  ANDN U7375 ( .B(start_reg[603]), .A(n4377), .Z(start_in[603]) );
  ANDN U7376 ( .B(start_reg[602]), .A(n4377), .Z(start_in[602]) );
  ANDN U7377 ( .B(start_reg[601]), .A(n4377), .Z(start_in[601]) );
  ANDN U7378 ( .B(start_reg[600]), .A(n4377), .Z(start_in[600]) );
  ANDN U7379 ( .B(start_reg[5]), .A(n4377), .Z(start_in[5]) );
  ANDN U7380 ( .B(start_reg[59]), .A(n4377), .Z(start_in[59]) );
  ANDN U7381 ( .B(start_reg[599]), .A(n4377), .Z(start_in[599]) );
  ANDN U7382 ( .B(start_reg[598]), .A(n4377), .Z(start_in[598]) );
  ANDN U7383 ( .B(start_reg[597]), .A(n4377), .Z(start_in[597]) );
  ANDN U7384 ( .B(start_reg[596]), .A(n4377), .Z(start_in[596]) );
  ANDN U7385 ( .B(start_reg[595]), .A(n4377), .Z(start_in[595]) );
  ANDN U7386 ( .B(start_reg[594]), .A(n4377), .Z(start_in[594]) );
  ANDN U7387 ( .B(start_reg[593]), .A(n4377), .Z(start_in[593]) );
  ANDN U7388 ( .B(start_reg[592]), .A(n4377), .Z(start_in[592]) );
  ANDN U7389 ( .B(start_reg[591]), .A(n4377), .Z(start_in[591]) );
  ANDN U7390 ( .B(start_reg[590]), .A(n4377), .Z(start_in[590]) );
  ANDN U7391 ( .B(start_reg[58]), .A(n4377), .Z(start_in[58]) );
  ANDN U7392 ( .B(start_reg[589]), .A(n4377), .Z(start_in[589]) );
  ANDN U7393 ( .B(start_reg[588]), .A(n4377), .Z(start_in[588]) );
  ANDN U7394 ( .B(start_reg[587]), .A(n4377), .Z(start_in[587]) );
  ANDN U7395 ( .B(start_reg[586]), .A(n4377), .Z(start_in[586]) );
  ANDN U7396 ( .B(start_reg[585]), .A(n4377), .Z(start_in[585]) );
  ANDN U7397 ( .B(start_reg[584]), .A(n4377), .Z(start_in[584]) );
  ANDN U7398 ( .B(start_reg[583]), .A(n4377), .Z(start_in[583]) );
  ANDN U7399 ( .B(start_reg[582]), .A(n4377), .Z(start_in[582]) );
  ANDN U7400 ( .B(start_reg[581]), .A(n4377), .Z(start_in[581]) );
  ANDN U7401 ( .B(start_reg[580]), .A(n4377), .Z(start_in[580]) );
  ANDN U7402 ( .B(start_reg[57]), .A(n4377), .Z(start_in[57]) );
  ANDN U7403 ( .B(start_reg[579]), .A(n4377), .Z(start_in[579]) );
  ANDN U7404 ( .B(start_reg[578]), .A(n4377), .Z(start_in[578]) );
  ANDN U7405 ( .B(start_reg[577]), .A(n4377), .Z(start_in[577]) );
  ANDN U7406 ( .B(start_reg[576]), .A(n4377), .Z(start_in[576]) );
  ANDN U7407 ( .B(start_reg[575]), .A(n4377), .Z(start_in[575]) );
  ANDN U7408 ( .B(start_reg[574]), .A(n4377), .Z(start_in[574]) );
  ANDN U7409 ( .B(start_reg[573]), .A(n4377), .Z(start_in[573]) );
  ANDN U7410 ( .B(start_reg[572]), .A(n4377), .Z(start_in[572]) );
  ANDN U7411 ( .B(start_reg[571]), .A(n4377), .Z(start_in[571]) );
  ANDN U7412 ( .B(start_reg[570]), .A(n4377), .Z(start_in[570]) );
  ANDN U7413 ( .B(start_reg[56]), .A(n4377), .Z(start_in[56]) );
  ANDN U7414 ( .B(start_reg[569]), .A(n4377), .Z(start_in[569]) );
  ANDN U7415 ( .B(start_reg[568]), .A(n4377), .Z(start_in[568]) );
  ANDN U7416 ( .B(start_reg[567]), .A(n4377), .Z(start_in[567]) );
  ANDN U7417 ( .B(start_reg[566]), .A(n4377), .Z(start_in[566]) );
  ANDN U7418 ( .B(start_reg[565]), .A(n4377), .Z(start_in[565]) );
  ANDN U7419 ( .B(start_reg[564]), .A(n4377), .Z(start_in[564]) );
  ANDN U7420 ( .B(start_reg[563]), .A(n4377), .Z(start_in[563]) );
  ANDN U7421 ( .B(start_reg[562]), .A(n4377), .Z(start_in[562]) );
  ANDN U7422 ( .B(start_reg[561]), .A(n4377), .Z(start_in[561]) );
  ANDN U7423 ( .B(start_reg[560]), .A(n4377), .Z(start_in[560]) );
  ANDN U7424 ( .B(start_reg[55]), .A(n4377), .Z(start_in[55]) );
  ANDN U7425 ( .B(start_reg[559]), .A(n4377), .Z(start_in[559]) );
  ANDN U7426 ( .B(start_reg[558]), .A(n4377), .Z(start_in[558]) );
  ANDN U7427 ( .B(start_reg[557]), .A(n4377), .Z(start_in[557]) );
  ANDN U7428 ( .B(start_reg[556]), .A(n4377), .Z(start_in[556]) );
  ANDN U7429 ( .B(start_reg[555]), .A(n4377), .Z(start_in[555]) );
  ANDN U7430 ( .B(start_reg[554]), .A(n4377), .Z(start_in[554]) );
  ANDN U7431 ( .B(start_reg[553]), .A(n4377), .Z(start_in[553]) );
  ANDN U7432 ( .B(start_reg[552]), .A(n4377), .Z(start_in[552]) );
  ANDN U7433 ( .B(start_reg[551]), .A(n4377), .Z(start_in[551]) );
  ANDN U7434 ( .B(start_reg[550]), .A(n4377), .Z(start_in[550]) );
  ANDN U7435 ( .B(start_reg[54]), .A(n4377), .Z(start_in[54]) );
  ANDN U7436 ( .B(start_reg[549]), .A(n4377), .Z(start_in[549]) );
  ANDN U7437 ( .B(start_reg[548]), .A(n4377), .Z(start_in[548]) );
  ANDN U7438 ( .B(start_reg[547]), .A(n4377), .Z(start_in[547]) );
  ANDN U7439 ( .B(start_reg[546]), .A(n4377), .Z(start_in[546]) );
  ANDN U7440 ( .B(start_reg[545]), .A(n4377), .Z(start_in[545]) );
  ANDN U7441 ( .B(start_reg[544]), .A(n4377), .Z(start_in[544]) );
  ANDN U7442 ( .B(start_reg[543]), .A(n4377), .Z(start_in[543]) );
  ANDN U7443 ( .B(start_reg[542]), .A(n4377), .Z(start_in[542]) );
  ANDN U7444 ( .B(start_reg[541]), .A(n4377), .Z(start_in[541]) );
  ANDN U7445 ( .B(start_reg[540]), .A(n4377), .Z(start_in[540]) );
  ANDN U7446 ( .B(start_reg[53]), .A(n4377), .Z(start_in[53]) );
  ANDN U7447 ( .B(start_reg[539]), .A(n4377), .Z(start_in[539]) );
  ANDN U7448 ( .B(start_reg[538]), .A(n4377), .Z(start_in[538]) );
  ANDN U7449 ( .B(start_reg[537]), .A(n4377), .Z(start_in[537]) );
  ANDN U7450 ( .B(start_reg[536]), .A(n4377), .Z(start_in[536]) );
  ANDN U7451 ( .B(start_reg[535]), .A(n4377), .Z(start_in[535]) );
  ANDN U7452 ( .B(start_reg[534]), .A(n4377), .Z(start_in[534]) );
  ANDN U7453 ( .B(start_reg[533]), .A(n4377), .Z(start_in[533]) );
  ANDN U7454 ( .B(start_reg[532]), .A(n4377), .Z(start_in[532]) );
  ANDN U7455 ( .B(start_reg[531]), .A(n4377), .Z(start_in[531]) );
  ANDN U7456 ( .B(start_reg[530]), .A(n4377), .Z(start_in[530]) );
  ANDN U7457 ( .B(start_reg[52]), .A(n4377), .Z(start_in[52]) );
  ANDN U7458 ( .B(start_reg[529]), .A(n4377), .Z(start_in[529]) );
  ANDN U7459 ( .B(start_reg[528]), .A(n4377), .Z(start_in[528]) );
  ANDN U7460 ( .B(start_reg[527]), .A(n4377), .Z(start_in[527]) );
  ANDN U7461 ( .B(start_reg[526]), .A(n4377), .Z(start_in[526]) );
  ANDN U7462 ( .B(start_reg[525]), .A(n4377), .Z(start_in[525]) );
  ANDN U7463 ( .B(start_reg[524]), .A(n4377), .Z(start_in[524]) );
  ANDN U7464 ( .B(start_reg[523]), .A(n4377), .Z(start_in[523]) );
  ANDN U7465 ( .B(start_reg[522]), .A(n4377), .Z(start_in[522]) );
  ANDN U7466 ( .B(start_reg[521]), .A(n4377), .Z(start_in[521]) );
  ANDN U7467 ( .B(start_reg[520]), .A(n4377), .Z(start_in[520]) );
  ANDN U7468 ( .B(start_reg[51]), .A(n4377), .Z(start_in[51]) );
  ANDN U7469 ( .B(start_reg[519]), .A(n4377), .Z(start_in[519]) );
  ANDN U7470 ( .B(start_reg[518]), .A(n4377), .Z(start_in[518]) );
  ANDN U7471 ( .B(start_reg[517]), .A(n4377), .Z(start_in[517]) );
  ANDN U7472 ( .B(start_reg[516]), .A(n4377), .Z(start_in[516]) );
  ANDN U7473 ( .B(start_reg[515]), .A(n4377), .Z(start_in[515]) );
  ANDN U7474 ( .B(start_reg[514]), .A(n4377), .Z(start_in[514]) );
  ANDN U7475 ( .B(start_reg[513]), .A(n4377), .Z(start_in[513]) );
  ANDN U7476 ( .B(start_reg[512]), .A(n4377), .Z(start_in[512]) );
  ANDN U7477 ( .B(start_reg[511]), .A(n4377), .Z(start_in[511]) );
  ANDN U7478 ( .B(start_reg[510]), .A(n4377), .Z(start_in[510]) );
  ANDN U7479 ( .B(start_reg[50]), .A(n4377), .Z(start_in[50]) );
  ANDN U7480 ( .B(start_reg[509]), .A(n4377), .Z(start_in[509]) );
  ANDN U7481 ( .B(start_reg[508]), .A(n4377), .Z(start_in[508]) );
  ANDN U7482 ( .B(start_reg[507]), .A(n4377), .Z(start_in[507]) );
  ANDN U7483 ( .B(start_reg[506]), .A(n4377), .Z(start_in[506]) );
  ANDN U7484 ( .B(start_reg[505]), .A(n4377), .Z(start_in[505]) );
  ANDN U7485 ( .B(start_reg[504]), .A(n4377), .Z(start_in[504]) );
  ANDN U7486 ( .B(start_reg[503]), .A(n4377), .Z(start_in[503]) );
  ANDN U7487 ( .B(start_reg[502]), .A(n4377), .Z(start_in[502]) );
  ANDN U7488 ( .B(start_reg[501]), .A(n4377), .Z(start_in[501]) );
  ANDN U7489 ( .B(start_reg[500]), .A(n4377), .Z(start_in[500]) );
  ANDN U7490 ( .B(start_reg[4]), .A(n4377), .Z(start_in[4]) );
  ANDN U7491 ( .B(start_reg[49]), .A(n4377), .Z(start_in[49]) );
  ANDN U7492 ( .B(start_reg[499]), .A(n4377), .Z(start_in[499]) );
  ANDN U7493 ( .B(start_reg[498]), .A(n4377), .Z(start_in[498]) );
  ANDN U7494 ( .B(start_reg[497]), .A(n4377), .Z(start_in[497]) );
  ANDN U7495 ( .B(start_reg[496]), .A(n4377), .Z(start_in[496]) );
  ANDN U7496 ( .B(start_reg[495]), .A(n4377), .Z(start_in[495]) );
  ANDN U7497 ( .B(start_reg[494]), .A(n4377), .Z(start_in[494]) );
  ANDN U7498 ( .B(start_reg[493]), .A(n4377), .Z(start_in[493]) );
  ANDN U7499 ( .B(start_reg[492]), .A(n4377), .Z(start_in[492]) );
  ANDN U7500 ( .B(start_reg[491]), .A(n4377), .Z(start_in[491]) );
  ANDN U7501 ( .B(start_reg[490]), .A(n4377), .Z(start_in[490]) );
  ANDN U7502 ( .B(start_reg[48]), .A(n4377), .Z(start_in[48]) );
  ANDN U7503 ( .B(start_reg[489]), .A(n4377), .Z(start_in[489]) );
  ANDN U7504 ( .B(start_reg[488]), .A(n4377), .Z(start_in[488]) );
  ANDN U7505 ( .B(start_reg[487]), .A(n4377), .Z(start_in[487]) );
  ANDN U7506 ( .B(start_reg[486]), .A(n4377), .Z(start_in[486]) );
  ANDN U7507 ( .B(start_reg[485]), .A(n4377), .Z(start_in[485]) );
  ANDN U7508 ( .B(start_reg[484]), .A(n4377), .Z(start_in[484]) );
  ANDN U7509 ( .B(start_reg[483]), .A(n4377), .Z(start_in[483]) );
  ANDN U7510 ( .B(start_reg[482]), .A(n4377), .Z(start_in[482]) );
  ANDN U7511 ( .B(start_reg[481]), .A(n4377), .Z(start_in[481]) );
  ANDN U7512 ( .B(start_reg[480]), .A(n4377), .Z(start_in[480]) );
  ANDN U7513 ( .B(start_reg[47]), .A(n4377), .Z(start_in[47]) );
  ANDN U7514 ( .B(start_reg[479]), .A(n4377), .Z(start_in[479]) );
  ANDN U7515 ( .B(start_reg[478]), .A(n4377), .Z(start_in[478]) );
  ANDN U7516 ( .B(start_reg[477]), .A(n4377), .Z(start_in[477]) );
  ANDN U7517 ( .B(start_reg[476]), .A(n4377), .Z(start_in[476]) );
  ANDN U7518 ( .B(start_reg[475]), .A(n4377), .Z(start_in[475]) );
  ANDN U7519 ( .B(start_reg[474]), .A(n4377), .Z(start_in[474]) );
  ANDN U7520 ( .B(start_reg[473]), .A(n4377), .Z(start_in[473]) );
  ANDN U7521 ( .B(start_reg[472]), .A(n4377), .Z(start_in[472]) );
  ANDN U7522 ( .B(start_reg[471]), .A(n4377), .Z(start_in[471]) );
  ANDN U7523 ( .B(start_reg[470]), .A(n4377), .Z(start_in[470]) );
  ANDN U7524 ( .B(start_reg[46]), .A(n4377), .Z(start_in[46]) );
  ANDN U7525 ( .B(start_reg[469]), .A(n4377), .Z(start_in[469]) );
  ANDN U7526 ( .B(start_reg[468]), .A(n4377), .Z(start_in[468]) );
  ANDN U7527 ( .B(start_reg[467]), .A(n4377), .Z(start_in[467]) );
  ANDN U7528 ( .B(start_reg[466]), .A(n4377), .Z(start_in[466]) );
  ANDN U7529 ( .B(start_reg[465]), .A(n4377), .Z(start_in[465]) );
  ANDN U7530 ( .B(start_reg[464]), .A(n4377), .Z(start_in[464]) );
  ANDN U7531 ( .B(start_reg[463]), .A(n4377), .Z(start_in[463]) );
  ANDN U7532 ( .B(start_reg[462]), .A(n4377), .Z(start_in[462]) );
  ANDN U7533 ( .B(start_reg[461]), .A(n4377), .Z(start_in[461]) );
  ANDN U7534 ( .B(start_reg[460]), .A(n4377), .Z(start_in[460]) );
  ANDN U7535 ( .B(start_reg[45]), .A(n4377), .Z(start_in[45]) );
  ANDN U7536 ( .B(start_reg[459]), .A(n4377), .Z(start_in[459]) );
  ANDN U7537 ( .B(start_reg[458]), .A(n4377), .Z(start_in[458]) );
  ANDN U7538 ( .B(start_reg[457]), .A(n4377), .Z(start_in[457]) );
  ANDN U7539 ( .B(start_reg[456]), .A(n4377), .Z(start_in[456]) );
  ANDN U7540 ( .B(start_reg[455]), .A(n4377), .Z(start_in[455]) );
  ANDN U7541 ( .B(start_reg[454]), .A(n4377), .Z(start_in[454]) );
  ANDN U7542 ( .B(start_reg[453]), .A(n4377), .Z(start_in[453]) );
  ANDN U7543 ( .B(start_reg[452]), .A(n4377), .Z(start_in[452]) );
  ANDN U7544 ( .B(start_reg[451]), .A(n4377), .Z(start_in[451]) );
  ANDN U7545 ( .B(start_reg[450]), .A(n4377), .Z(start_in[450]) );
  ANDN U7546 ( .B(start_reg[44]), .A(n4377), .Z(start_in[44]) );
  ANDN U7547 ( .B(start_reg[449]), .A(n4377), .Z(start_in[449]) );
  ANDN U7548 ( .B(start_reg[448]), .A(n4377), .Z(start_in[448]) );
  ANDN U7549 ( .B(start_reg[447]), .A(n4377), .Z(start_in[447]) );
  ANDN U7550 ( .B(start_reg[446]), .A(n4377), .Z(start_in[446]) );
  ANDN U7551 ( .B(start_reg[445]), .A(n4377), .Z(start_in[445]) );
  ANDN U7552 ( .B(start_reg[444]), .A(n4377), .Z(start_in[444]) );
  ANDN U7553 ( .B(start_reg[443]), .A(n4377), .Z(start_in[443]) );
  ANDN U7554 ( .B(start_reg[442]), .A(n4377), .Z(start_in[442]) );
  ANDN U7555 ( .B(start_reg[441]), .A(n4377), .Z(start_in[441]) );
  ANDN U7556 ( .B(start_reg[440]), .A(n4377), .Z(start_in[440]) );
  ANDN U7557 ( .B(start_reg[43]), .A(n4377), .Z(start_in[43]) );
  ANDN U7558 ( .B(start_reg[439]), .A(n4377), .Z(start_in[439]) );
  ANDN U7559 ( .B(start_reg[438]), .A(n4377), .Z(start_in[438]) );
  ANDN U7560 ( .B(start_reg[437]), .A(n4377), .Z(start_in[437]) );
  ANDN U7561 ( .B(start_reg[436]), .A(n4377), .Z(start_in[436]) );
  ANDN U7562 ( .B(start_reg[435]), .A(n4377), .Z(start_in[435]) );
  ANDN U7563 ( .B(start_reg[434]), .A(n4377), .Z(start_in[434]) );
  ANDN U7564 ( .B(start_reg[433]), .A(n4377), .Z(start_in[433]) );
  ANDN U7565 ( .B(start_reg[432]), .A(n4377), .Z(start_in[432]) );
  ANDN U7566 ( .B(start_reg[431]), .A(n4377), .Z(start_in[431]) );
  ANDN U7567 ( .B(start_reg[430]), .A(n4377), .Z(start_in[430]) );
  ANDN U7568 ( .B(start_reg[42]), .A(n4377), .Z(start_in[42]) );
  ANDN U7569 ( .B(start_reg[429]), .A(n4377), .Z(start_in[429]) );
  ANDN U7570 ( .B(start_reg[428]), .A(n4377), .Z(start_in[428]) );
  ANDN U7571 ( .B(start_reg[427]), .A(n4377), .Z(start_in[427]) );
  ANDN U7572 ( .B(start_reg[426]), .A(n4377), .Z(start_in[426]) );
  ANDN U7573 ( .B(start_reg[425]), .A(n4377), .Z(start_in[425]) );
  ANDN U7574 ( .B(start_reg[424]), .A(n4377), .Z(start_in[424]) );
  ANDN U7575 ( .B(start_reg[423]), .A(n4377), .Z(start_in[423]) );
  ANDN U7576 ( .B(start_reg[422]), .A(n4377), .Z(start_in[422]) );
  ANDN U7577 ( .B(start_reg[421]), .A(n4377), .Z(start_in[421]) );
  ANDN U7578 ( .B(start_reg[420]), .A(n4377), .Z(start_in[420]) );
  ANDN U7579 ( .B(start_reg[41]), .A(n4377), .Z(start_in[41]) );
  ANDN U7580 ( .B(start_reg[419]), .A(n4377), .Z(start_in[419]) );
  ANDN U7581 ( .B(start_reg[418]), .A(n4377), .Z(start_in[418]) );
  ANDN U7582 ( .B(start_reg[417]), .A(n4377), .Z(start_in[417]) );
  ANDN U7583 ( .B(start_reg[416]), .A(n4377), .Z(start_in[416]) );
  ANDN U7584 ( .B(start_reg[415]), .A(n4377), .Z(start_in[415]) );
  ANDN U7585 ( .B(start_reg[414]), .A(n4377), .Z(start_in[414]) );
  ANDN U7586 ( .B(start_reg[413]), .A(n4377), .Z(start_in[413]) );
  ANDN U7587 ( .B(start_reg[412]), .A(n4377), .Z(start_in[412]) );
  ANDN U7588 ( .B(start_reg[411]), .A(n4377), .Z(start_in[411]) );
  ANDN U7589 ( .B(start_reg[410]), .A(n4377), .Z(start_in[410]) );
  ANDN U7590 ( .B(start_reg[40]), .A(n4377), .Z(start_in[40]) );
  ANDN U7591 ( .B(start_reg[409]), .A(n4377), .Z(start_in[409]) );
  ANDN U7592 ( .B(start_reg[408]), .A(n4377), .Z(start_in[408]) );
  ANDN U7593 ( .B(start_reg[407]), .A(n4377), .Z(start_in[407]) );
  ANDN U7594 ( .B(start_reg[406]), .A(n4377), .Z(start_in[406]) );
  ANDN U7595 ( .B(start_reg[405]), .A(n4377), .Z(start_in[405]) );
  ANDN U7596 ( .B(start_reg[404]), .A(n4377), .Z(start_in[404]) );
  ANDN U7597 ( .B(start_reg[403]), .A(n4377), .Z(start_in[403]) );
  ANDN U7598 ( .B(start_reg[402]), .A(n4377), .Z(start_in[402]) );
  ANDN U7599 ( .B(start_reg[401]), .A(n4377), .Z(start_in[401]) );
  ANDN U7600 ( .B(start_reg[400]), .A(n4377), .Z(start_in[400]) );
  ANDN U7601 ( .B(start_reg[3]), .A(n4377), .Z(start_in[3]) );
  ANDN U7602 ( .B(start_reg[39]), .A(n4377), .Z(start_in[39]) );
  ANDN U7603 ( .B(start_reg[399]), .A(n4377), .Z(start_in[399]) );
  ANDN U7604 ( .B(start_reg[398]), .A(n4377), .Z(start_in[398]) );
  ANDN U7605 ( .B(start_reg[397]), .A(n4377), .Z(start_in[397]) );
  ANDN U7606 ( .B(start_reg[396]), .A(n4377), .Z(start_in[396]) );
  ANDN U7607 ( .B(start_reg[395]), .A(n4377), .Z(start_in[395]) );
  ANDN U7608 ( .B(start_reg[394]), .A(n4377), .Z(start_in[394]) );
  ANDN U7609 ( .B(start_reg[393]), .A(n4377), .Z(start_in[393]) );
  ANDN U7610 ( .B(start_reg[392]), .A(n4377), .Z(start_in[392]) );
  ANDN U7611 ( .B(start_reg[391]), .A(n4377), .Z(start_in[391]) );
  ANDN U7612 ( .B(start_reg[390]), .A(n4377), .Z(start_in[390]) );
  ANDN U7613 ( .B(start_reg[38]), .A(n4377), .Z(start_in[38]) );
  ANDN U7614 ( .B(start_reg[389]), .A(n4377), .Z(start_in[389]) );
  ANDN U7615 ( .B(start_reg[388]), .A(n4377), .Z(start_in[388]) );
  ANDN U7616 ( .B(start_reg[387]), .A(n4377), .Z(start_in[387]) );
  ANDN U7617 ( .B(start_reg[386]), .A(n4377), .Z(start_in[386]) );
  ANDN U7618 ( .B(start_reg[385]), .A(n4377), .Z(start_in[385]) );
  ANDN U7619 ( .B(start_reg[384]), .A(n4377), .Z(start_in[384]) );
  ANDN U7620 ( .B(start_reg[383]), .A(n4377), .Z(start_in[383]) );
  ANDN U7621 ( .B(start_reg[382]), .A(n4377), .Z(start_in[382]) );
  ANDN U7622 ( .B(start_reg[381]), .A(n4377), .Z(start_in[381]) );
  ANDN U7623 ( .B(start_reg[380]), .A(n4377), .Z(start_in[380]) );
  ANDN U7624 ( .B(start_reg[37]), .A(n4377), .Z(start_in[37]) );
  ANDN U7625 ( .B(start_reg[379]), .A(n4377), .Z(start_in[379]) );
  ANDN U7626 ( .B(start_reg[378]), .A(n4377), .Z(start_in[378]) );
  ANDN U7627 ( .B(start_reg[377]), .A(n4377), .Z(start_in[377]) );
  ANDN U7628 ( .B(start_reg[376]), .A(n4377), .Z(start_in[376]) );
  ANDN U7629 ( .B(start_reg[375]), .A(n4377), .Z(start_in[375]) );
  ANDN U7630 ( .B(start_reg[374]), .A(n4377), .Z(start_in[374]) );
  ANDN U7631 ( .B(start_reg[373]), .A(n4377), .Z(start_in[373]) );
  ANDN U7632 ( .B(start_reg[372]), .A(n4377), .Z(start_in[372]) );
  ANDN U7633 ( .B(start_reg[371]), .A(n4377), .Z(start_in[371]) );
  ANDN U7634 ( .B(start_reg[370]), .A(n4377), .Z(start_in[370]) );
  ANDN U7635 ( .B(start_reg[36]), .A(n4377), .Z(start_in[36]) );
  ANDN U7636 ( .B(start_reg[369]), .A(n4377), .Z(start_in[369]) );
  ANDN U7637 ( .B(start_reg[368]), .A(n4377), .Z(start_in[368]) );
  ANDN U7638 ( .B(start_reg[367]), .A(n4377), .Z(start_in[367]) );
  ANDN U7639 ( .B(start_reg[366]), .A(n4377), .Z(start_in[366]) );
  ANDN U7640 ( .B(start_reg[365]), .A(n4377), .Z(start_in[365]) );
  ANDN U7641 ( .B(start_reg[364]), .A(n4377), .Z(start_in[364]) );
  ANDN U7642 ( .B(start_reg[363]), .A(n4377), .Z(start_in[363]) );
  ANDN U7643 ( .B(start_reg[362]), .A(n4377), .Z(start_in[362]) );
  ANDN U7644 ( .B(start_reg[361]), .A(n4377), .Z(start_in[361]) );
  ANDN U7645 ( .B(start_reg[360]), .A(n4377), .Z(start_in[360]) );
  ANDN U7646 ( .B(start_reg[35]), .A(n4377), .Z(start_in[35]) );
  ANDN U7647 ( .B(start_reg[359]), .A(n4377), .Z(start_in[359]) );
  ANDN U7648 ( .B(start_reg[358]), .A(n4377), .Z(start_in[358]) );
  ANDN U7649 ( .B(start_reg[357]), .A(n4377), .Z(start_in[357]) );
  ANDN U7650 ( .B(start_reg[356]), .A(n4377), .Z(start_in[356]) );
  ANDN U7651 ( .B(start_reg[355]), .A(n4377), .Z(start_in[355]) );
  ANDN U7652 ( .B(start_reg[354]), .A(n4377), .Z(start_in[354]) );
  ANDN U7653 ( .B(start_reg[353]), .A(n4377), .Z(start_in[353]) );
  ANDN U7654 ( .B(start_reg[352]), .A(n4377), .Z(start_in[352]) );
  ANDN U7655 ( .B(start_reg[351]), .A(n4377), .Z(start_in[351]) );
  ANDN U7656 ( .B(start_reg[350]), .A(n4377), .Z(start_in[350]) );
  ANDN U7657 ( .B(start_reg[34]), .A(n4377), .Z(start_in[34]) );
  ANDN U7658 ( .B(start_reg[349]), .A(n4377), .Z(start_in[349]) );
  ANDN U7659 ( .B(start_reg[348]), .A(n4377), .Z(start_in[348]) );
  ANDN U7660 ( .B(start_reg[347]), .A(n4377), .Z(start_in[347]) );
  ANDN U7661 ( .B(start_reg[346]), .A(n4377), .Z(start_in[346]) );
  ANDN U7662 ( .B(start_reg[345]), .A(n4377), .Z(start_in[345]) );
  ANDN U7663 ( .B(start_reg[344]), .A(n4377), .Z(start_in[344]) );
  ANDN U7664 ( .B(start_reg[343]), .A(n4377), .Z(start_in[343]) );
  ANDN U7665 ( .B(start_reg[342]), .A(n4377), .Z(start_in[342]) );
  ANDN U7666 ( .B(start_reg[341]), .A(n4377), .Z(start_in[341]) );
  ANDN U7667 ( .B(start_reg[340]), .A(n4377), .Z(start_in[340]) );
  ANDN U7668 ( .B(start_reg[33]), .A(n4377), .Z(start_in[33]) );
  ANDN U7669 ( .B(start_reg[339]), .A(n4377), .Z(start_in[339]) );
  ANDN U7670 ( .B(start_reg[338]), .A(n4377), .Z(start_in[338]) );
  ANDN U7671 ( .B(start_reg[337]), .A(n4377), .Z(start_in[337]) );
  ANDN U7672 ( .B(start_reg[336]), .A(n4377), .Z(start_in[336]) );
  ANDN U7673 ( .B(start_reg[335]), .A(n4377), .Z(start_in[335]) );
  ANDN U7674 ( .B(start_reg[334]), .A(n4377), .Z(start_in[334]) );
  ANDN U7675 ( .B(start_reg[333]), .A(n4377), .Z(start_in[333]) );
  ANDN U7676 ( .B(start_reg[332]), .A(n4377), .Z(start_in[332]) );
  ANDN U7677 ( .B(start_reg[331]), .A(n4377), .Z(start_in[331]) );
  ANDN U7678 ( .B(start_reg[330]), .A(n4377), .Z(start_in[330]) );
  ANDN U7679 ( .B(start_reg[32]), .A(n4377), .Z(start_in[32]) );
  ANDN U7680 ( .B(start_reg[329]), .A(n4377), .Z(start_in[329]) );
  ANDN U7681 ( .B(start_reg[328]), .A(n4377), .Z(start_in[328]) );
  ANDN U7682 ( .B(start_reg[327]), .A(n4377), .Z(start_in[327]) );
  ANDN U7683 ( .B(start_reg[326]), .A(n4377), .Z(start_in[326]) );
  ANDN U7684 ( .B(start_reg[325]), .A(n4377), .Z(start_in[325]) );
  ANDN U7685 ( .B(start_reg[324]), .A(n4377), .Z(start_in[324]) );
  ANDN U7686 ( .B(start_reg[323]), .A(n4377), .Z(start_in[323]) );
  ANDN U7687 ( .B(start_reg[322]), .A(n4377), .Z(start_in[322]) );
  ANDN U7688 ( .B(start_reg[321]), .A(n4377), .Z(start_in[321]) );
  ANDN U7689 ( .B(start_reg[320]), .A(n4377), .Z(start_in[320]) );
  ANDN U7690 ( .B(start_reg[31]), .A(n4377), .Z(start_in[31]) );
  ANDN U7691 ( .B(start_reg[319]), .A(n4377), .Z(start_in[319]) );
  ANDN U7692 ( .B(start_reg[318]), .A(n4377), .Z(start_in[318]) );
  ANDN U7693 ( .B(start_reg[317]), .A(n4377), .Z(start_in[317]) );
  ANDN U7694 ( .B(start_reg[316]), .A(n4377), .Z(start_in[316]) );
  ANDN U7695 ( .B(start_reg[315]), .A(n4377), .Z(start_in[315]) );
  ANDN U7696 ( .B(start_reg[314]), .A(n4377), .Z(start_in[314]) );
  ANDN U7697 ( .B(start_reg[313]), .A(n4377), .Z(start_in[313]) );
  ANDN U7698 ( .B(start_reg[312]), .A(n4377), .Z(start_in[312]) );
  ANDN U7699 ( .B(start_reg[311]), .A(n4377), .Z(start_in[311]) );
  ANDN U7700 ( .B(start_reg[310]), .A(n4377), .Z(start_in[310]) );
  ANDN U7701 ( .B(start_reg[30]), .A(n4377), .Z(start_in[30]) );
  ANDN U7702 ( .B(start_reg[309]), .A(n4377), .Z(start_in[309]) );
  ANDN U7703 ( .B(start_reg[308]), .A(n4377), .Z(start_in[308]) );
  ANDN U7704 ( .B(start_reg[307]), .A(n4377), .Z(start_in[307]) );
  ANDN U7705 ( .B(start_reg[306]), .A(n4377), .Z(start_in[306]) );
  ANDN U7706 ( .B(start_reg[305]), .A(n4377), .Z(start_in[305]) );
  ANDN U7707 ( .B(start_reg[304]), .A(n4377), .Z(start_in[304]) );
  ANDN U7708 ( .B(start_reg[303]), .A(n4377), .Z(start_in[303]) );
  ANDN U7709 ( .B(start_reg[302]), .A(n4377), .Z(start_in[302]) );
  ANDN U7710 ( .B(start_reg[301]), .A(n4377), .Z(start_in[301]) );
  ANDN U7711 ( .B(start_reg[300]), .A(n4377), .Z(start_in[300]) );
  ANDN U7712 ( .B(start_reg[2]), .A(n4377), .Z(start_in[2]) );
  ANDN U7713 ( .B(start_reg[29]), .A(n4377), .Z(start_in[29]) );
  ANDN U7714 ( .B(start_reg[299]), .A(n4377), .Z(start_in[299]) );
  ANDN U7715 ( .B(start_reg[298]), .A(n4377), .Z(start_in[298]) );
  ANDN U7716 ( .B(start_reg[297]), .A(n4377), .Z(start_in[297]) );
  ANDN U7717 ( .B(start_reg[296]), .A(n4377), .Z(start_in[296]) );
  ANDN U7718 ( .B(start_reg[295]), .A(n4377), .Z(start_in[295]) );
  ANDN U7719 ( .B(start_reg[294]), .A(n4377), .Z(start_in[294]) );
  ANDN U7720 ( .B(start_reg[293]), .A(n4377), .Z(start_in[293]) );
  ANDN U7721 ( .B(start_reg[292]), .A(n4377), .Z(start_in[292]) );
  ANDN U7722 ( .B(start_reg[291]), .A(n4377), .Z(start_in[291]) );
  ANDN U7723 ( .B(start_reg[290]), .A(n4377), .Z(start_in[290]) );
  ANDN U7724 ( .B(start_reg[28]), .A(n4377), .Z(start_in[28]) );
  ANDN U7725 ( .B(start_reg[289]), .A(n4377), .Z(start_in[289]) );
  ANDN U7726 ( .B(start_reg[288]), .A(n4377), .Z(start_in[288]) );
  ANDN U7727 ( .B(start_reg[287]), .A(n4377), .Z(start_in[287]) );
  ANDN U7728 ( .B(start_reg[286]), .A(n4377), .Z(start_in[286]) );
  ANDN U7729 ( .B(start_reg[285]), .A(n4377), .Z(start_in[285]) );
  ANDN U7730 ( .B(start_reg[284]), .A(n4377), .Z(start_in[284]) );
  ANDN U7731 ( .B(start_reg[283]), .A(n4377), .Z(start_in[283]) );
  ANDN U7732 ( .B(start_reg[282]), .A(n4377), .Z(start_in[282]) );
  ANDN U7733 ( .B(start_reg[281]), .A(n4377), .Z(start_in[281]) );
  ANDN U7734 ( .B(start_reg[280]), .A(n4377), .Z(start_in[280]) );
  ANDN U7735 ( .B(start_reg[27]), .A(n4377), .Z(start_in[27]) );
  ANDN U7736 ( .B(start_reg[279]), .A(n4377), .Z(start_in[279]) );
  ANDN U7737 ( .B(start_reg[278]), .A(n4377), .Z(start_in[278]) );
  ANDN U7738 ( .B(start_reg[277]), .A(n4377), .Z(start_in[277]) );
  ANDN U7739 ( .B(start_reg[276]), .A(n4377), .Z(start_in[276]) );
  ANDN U7740 ( .B(start_reg[275]), .A(n4377), .Z(start_in[275]) );
  ANDN U7741 ( .B(start_reg[274]), .A(n4377), .Z(start_in[274]) );
  ANDN U7742 ( .B(start_reg[273]), .A(n4377), .Z(start_in[273]) );
  ANDN U7743 ( .B(start_reg[272]), .A(n4377), .Z(start_in[272]) );
  ANDN U7744 ( .B(start_reg[271]), .A(n4377), .Z(start_in[271]) );
  ANDN U7745 ( .B(start_reg[270]), .A(n4377), .Z(start_in[270]) );
  ANDN U7746 ( .B(start_reg[26]), .A(n4377), .Z(start_in[26]) );
  ANDN U7747 ( .B(start_reg[269]), .A(n4377), .Z(start_in[269]) );
  ANDN U7748 ( .B(start_reg[268]), .A(n4377), .Z(start_in[268]) );
  ANDN U7749 ( .B(start_reg[267]), .A(n4377), .Z(start_in[267]) );
  ANDN U7750 ( .B(start_reg[266]), .A(n4377), .Z(start_in[266]) );
  ANDN U7751 ( .B(start_reg[265]), .A(n4377), .Z(start_in[265]) );
  ANDN U7752 ( .B(start_reg[264]), .A(n4377), .Z(start_in[264]) );
  ANDN U7753 ( .B(start_reg[263]), .A(n4377), .Z(start_in[263]) );
  ANDN U7754 ( .B(start_reg[262]), .A(n4377), .Z(start_in[262]) );
  ANDN U7755 ( .B(start_reg[261]), .A(n4377), .Z(start_in[261]) );
  ANDN U7756 ( .B(start_reg[260]), .A(n4377), .Z(start_in[260]) );
  ANDN U7757 ( .B(start_reg[25]), .A(n4377), .Z(start_in[25]) );
  ANDN U7758 ( .B(start_reg[259]), .A(n4377), .Z(start_in[259]) );
  ANDN U7759 ( .B(start_reg[258]), .A(n4377), .Z(start_in[258]) );
  ANDN U7760 ( .B(start_reg[257]), .A(n4377), .Z(start_in[257]) );
  ANDN U7761 ( .B(start_reg[256]), .A(n4377), .Z(start_in[256]) );
  ANDN U7762 ( .B(start_reg[255]), .A(n4377), .Z(start_in[255]) );
  ANDN U7763 ( .B(start_reg[254]), .A(n4377), .Z(start_in[254]) );
  ANDN U7764 ( .B(start_reg[253]), .A(n4377), .Z(start_in[253]) );
  ANDN U7765 ( .B(start_reg[252]), .A(n4377), .Z(start_in[252]) );
  ANDN U7766 ( .B(start_reg[251]), .A(n4377), .Z(start_in[251]) );
  ANDN U7767 ( .B(start_reg[250]), .A(n4377), .Z(start_in[250]) );
  ANDN U7768 ( .B(start_reg[24]), .A(n4377), .Z(start_in[24]) );
  ANDN U7769 ( .B(start_reg[249]), .A(n4377), .Z(start_in[249]) );
  ANDN U7770 ( .B(start_reg[248]), .A(n4377), .Z(start_in[248]) );
  ANDN U7771 ( .B(start_reg[247]), .A(n4377), .Z(start_in[247]) );
  ANDN U7772 ( .B(start_reg[246]), .A(n4377), .Z(start_in[246]) );
  ANDN U7773 ( .B(start_reg[245]), .A(n4377), .Z(start_in[245]) );
  ANDN U7774 ( .B(start_reg[244]), .A(n4377), .Z(start_in[244]) );
  ANDN U7775 ( .B(start_reg[243]), .A(n4377), .Z(start_in[243]) );
  ANDN U7776 ( .B(start_reg[242]), .A(n4377), .Z(start_in[242]) );
  ANDN U7777 ( .B(start_reg[241]), .A(n4377), .Z(start_in[241]) );
  ANDN U7778 ( .B(start_reg[240]), .A(n4377), .Z(start_in[240]) );
  ANDN U7779 ( .B(start_reg[23]), .A(n4377), .Z(start_in[23]) );
  ANDN U7780 ( .B(start_reg[239]), .A(n4377), .Z(start_in[239]) );
  ANDN U7781 ( .B(start_reg[238]), .A(n4377), .Z(start_in[238]) );
  ANDN U7782 ( .B(start_reg[237]), .A(n4377), .Z(start_in[237]) );
  ANDN U7783 ( .B(start_reg[236]), .A(n4377), .Z(start_in[236]) );
  ANDN U7784 ( .B(start_reg[235]), .A(n4377), .Z(start_in[235]) );
  ANDN U7785 ( .B(start_reg[234]), .A(n4377), .Z(start_in[234]) );
  ANDN U7786 ( .B(start_reg[233]), .A(n4377), .Z(start_in[233]) );
  ANDN U7787 ( .B(start_reg[232]), .A(n4377), .Z(start_in[232]) );
  ANDN U7788 ( .B(start_reg[231]), .A(n4377), .Z(start_in[231]) );
  ANDN U7789 ( .B(start_reg[230]), .A(n4377), .Z(start_in[230]) );
  ANDN U7790 ( .B(start_reg[22]), .A(n4377), .Z(start_in[22]) );
  ANDN U7791 ( .B(start_reg[229]), .A(n4377), .Z(start_in[229]) );
  ANDN U7792 ( .B(start_reg[228]), .A(n4377), .Z(start_in[228]) );
  ANDN U7793 ( .B(start_reg[227]), .A(n4377), .Z(start_in[227]) );
  ANDN U7794 ( .B(start_reg[226]), .A(n4377), .Z(start_in[226]) );
  ANDN U7795 ( .B(start_reg[225]), .A(n4377), .Z(start_in[225]) );
  ANDN U7796 ( .B(start_reg[224]), .A(n4377), .Z(start_in[224]) );
  ANDN U7797 ( .B(start_reg[223]), .A(n4377), .Z(start_in[223]) );
  ANDN U7798 ( .B(start_reg[222]), .A(n4377), .Z(start_in[222]) );
  ANDN U7799 ( .B(start_reg[221]), .A(n4377), .Z(start_in[221]) );
  ANDN U7800 ( .B(start_reg[220]), .A(n4377), .Z(start_in[220]) );
  ANDN U7801 ( .B(start_reg[21]), .A(n4377), .Z(start_in[21]) );
  ANDN U7802 ( .B(start_reg[219]), .A(n4377), .Z(start_in[219]) );
  ANDN U7803 ( .B(start_reg[218]), .A(n4377), .Z(start_in[218]) );
  ANDN U7804 ( .B(start_reg[217]), .A(n4377), .Z(start_in[217]) );
  ANDN U7805 ( .B(start_reg[216]), .A(n4377), .Z(start_in[216]) );
  ANDN U7806 ( .B(start_reg[215]), .A(n4377), .Z(start_in[215]) );
  ANDN U7807 ( .B(start_reg[214]), .A(n4377), .Z(start_in[214]) );
  ANDN U7808 ( .B(start_reg[213]), .A(n4377), .Z(start_in[213]) );
  ANDN U7809 ( .B(start_reg[212]), .A(n4377), .Z(start_in[212]) );
  ANDN U7810 ( .B(start_reg[211]), .A(n4377), .Z(start_in[211]) );
  ANDN U7811 ( .B(start_reg[210]), .A(n4377), .Z(start_in[210]) );
  ANDN U7812 ( .B(start_reg[20]), .A(n4377), .Z(start_in[20]) );
  ANDN U7813 ( .B(start_reg[209]), .A(n4377), .Z(start_in[209]) );
  ANDN U7814 ( .B(start_reg[208]), .A(n4377), .Z(start_in[208]) );
  ANDN U7815 ( .B(start_reg[207]), .A(n4377), .Z(start_in[207]) );
  ANDN U7816 ( .B(start_reg[206]), .A(n4377), .Z(start_in[206]) );
  ANDN U7817 ( .B(start_reg[205]), .A(n4377), .Z(start_in[205]) );
  ANDN U7818 ( .B(start_reg[204]), .A(n4377), .Z(start_in[204]) );
  ANDN U7819 ( .B(start_reg[203]), .A(n4377), .Z(start_in[203]) );
  ANDN U7820 ( .B(start_reg[202]), .A(n4377), .Z(start_in[202]) );
  ANDN U7821 ( .B(start_reg[201]), .A(n4377), .Z(start_in[201]) );
  ANDN U7822 ( .B(start_reg[200]), .A(n4377), .Z(start_in[200]) );
  ANDN U7823 ( .B(start_reg[1]), .A(n4377), .Z(start_in[1]) );
  ANDN U7824 ( .B(start_reg[19]), .A(n4377), .Z(start_in[19]) );
  ANDN U7825 ( .B(start_reg[199]), .A(n4377), .Z(start_in[199]) );
  ANDN U7826 ( .B(start_reg[198]), .A(n4377), .Z(start_in[198]) );
  ANDN U7827 ( .B(start_reg[197]), .A(n4377), .Z(start_in[197]) );
  ANDN U7828 ( .B(start_reg[196]), .A(n4377), .Z(start_in[196]) );
  ANDN U7829 ( .B(start_reg[195]), .A(n4377), .Z(start_in[195]) );
  ANDN U7830 ( .B(start_reg[194]), .A(n4377), .Z(start_in[194]) );
  ANDN U7831 ( .B(start_reg[193]), .A(n4377), .Z(start_in[193]) );
  ANDN U7832 ( .B(start_reg[192]), .A(n4377), .Z(start_in[192]) );
  ANDN U7833 ( .B(start_reg[191]), .A(n4377), .Z(start_in[191]) );
  ANDN U7834 ( .B(start_reg[190]), .A(n4377), .Z(start_in[190]) );
  ANDN U7835 ( .B(start_reg[18]), .A(n4377), .Z(start_in[18]) );
  ANDN U7836 ( .B(start_reg[189]), .A(n4377), .Z(start_in[189]) );
  ANDN U7837 ( .B(start_reg[188]), .A(n4377), .Z(start_in[188]) );
  ANDN U7838 ( .B(start_reg[187]), .A(n4377), .Z(start_in[187]) );
  ANDN U7839 ( .B(start_reg[186]), .A(n4377), .Z(start_in[186]) );
  ANDN U7840 ( .B(start_reg[185]), .A(n4377), .Z(start_in[185]) );
  ANDN U7841 ( .B(start_reg[184]), .A(n4377), .Z(start_in[184]) );
  ANDN U7842 ( .B(start_reg[183]), .A(n4377), .Z(start_in[183]) );
  ANDN U7843 ( .B(start_reg[182]), .A(n4377), .Z(start_in[182]) );
  ANDN U7844 ( .B(start_reg[181]), .A(n4377), .Z(start_in[181]) );
  ANDN U7845 ( .B(start_reg[180]), .A(n4377), .Z(start_in[180]) );
  ANDN U7846 ( .B(start_reg[17]), .A(n4377), .Z(start_in[17]) );
  ANDN U7847 ( .B(start_reg[179]), .A(n4377), .Z(start_in[179]) );
  ANDN U7848 ( .B(start_reg[178]), .A(n4377), .Z(start_in[178]) );
  ANDN U7849 ( .B(start_reg[177]), .A(n4377), .Z(start_in[177]) );
  ANDN U7850 ( .B(start_reg[176]), .A(n4377), .Z(start_in[176]) );
  ANDN U7851 ( .B(start_reg[175]), .A(n4377), .Z(start_in[175]) );
  ANDN U7852 ( .B(start_reg[174]), .A(n4377), .Z(start_in[174]) );
  ANDN U7853 ( .B(start_reg[173]), .A(n4377), .Z(start_in[173]) );
  ANDN U7854 ( .B(start_reg[172]), .A(n4377), .Z(start_in[172]) );
  ANDN U7855 ( .B(start_reg[171]), .A(n4377), .Z(start_in[171]) );
  ANDN U7856 ( .B(start_reg[170]), .A(n4377), .Z(start_in[170]) );
  ANDN U7857 ( .B(start_reg[16]), .A(n4377), .Z(start_in[16]) );
  ANDN U7858 ( .B(start_reg[169]), .A(n4377), .Z(start_in[169]) );
  ANDN U7859 ( .B(start_reg[168]), .A(n4377), .Z(start_in[168]) );
  ANDN U7860 ( .B(start_reg[167]), .A(n4377), .Z(start_in[167]) );
  ANDN U7861 ( .B(start_reg[166]), .A(n4377), .Z(start_in[166]) );
  ANDN U7862 ( .B(start_reg[165]), .A(n4377), .Z(start_in[165]) );
  ANDN U7863 ( .B(start_reg[164]), .A(n4377), .Z(start_in[164]) );
  ANDN U7864 ( .B(start_reg[163]), .A(n4377), .Z(start_in[163]) );
  ANDN U7865 ( .B(start_reg[162]), .A(n4377), .Z(start_in[162]) );
  ANDN U7866 ( .B(start_reg[161]), .A(n4377), .Z(start_in[161]) );
  ANDN U7867 ( .B(start_reg[160]), .A(n4377), .Z(start_in[160]) );
  ANDN U7868 ( .B(start_reg[15]), .A(n4377), .Z(start_in[15]) );
  ANDN U7869 ( .B(start_reg[159]), .A(n4377), .Z(start_in[159]) );
  ANDN U7870 ( .B(start_reg[158]), .A(n4377), .Z(start_in[158]) );
  ANDN U7871 ( .B(start_reg[157]), .A(n4377), .Z(start_in[157]) );
  ANDN U7872 ( .B(start_reg[156]), .A(n4377), .Z(start_in[156]) );
  ANDN U7873 ( .B(start_reg[155]), .A(n4377), .Z(start_in[155]) );
  ANDN U7874 ( .B(start_reg[154]), .A(n4377), .Z(start_in[154]) );
  ANDN U7875 ( .B(start_reg[153]), .A(n4377), .Z(start_in[153]) );
  ANDN U7876 ( .B(start_reg[152]), .A(n4377), .Z(start_in[152]) );
  ANDN U7877 ( .B(start_reg[151]), .A(n4377), .Z(start_in[151]) );
  ANDN U7878 ( .B(start_reg[150]), .A(n4377), .Z(start_in[150]) );
  ANDN U7879 ( .B(start_reg[14]), .A(n4377), .Z(start_in[14]) );
  ANDN U7880 ( .B(start_reg[149]), .A(n4377), .Z(start_in[149]) );
  ANDN U7881 ( .B(start_reg[148]), .A(n4377), .Z(start_in[148]) );
  ANDN U7882 ( .B(start_reg[147]), .A(n4377), .Z(start_in[147]) );
  ANDN U7883 ( .B(start_reg[146]), .A(n4377), .Z(start_in[146]) );
  ANDN U7884 ( .B(start_reg[145]), .A(n4377), .Z(start_in[145]) );
  ANDN U7885 ( .B(start_reg[144]), .A(n4377), .Z(start_in[144]) );
  ANDN U7886 ( .B(start_reg[143]), .A(n4377), .Z(start_in[143]) );
  ANDN U7887 ( .B(start_reg[142]), .A(n4377), .Z(start_in[142]) );
  ANDN U7888 ( .B(start_reg[141]), .A(n4377), .Z(start_in[141]) );
  ANDN U7889 ( .B(start_reg[140]), .A(n4377), .Z(start_in[140]) );
  ANDN U7890 ( .B(start_reg[13]), .A(n4377), .Z(start_in[13]) );
  ANDN U7891 ( .B(start_reg[139]), .A(n4377), .Z(start_in[139]) );
  ANDN U7892 ( .B(start_reg[138]), .A(n4377), .Z(start_in[138]) );
  ANDN U7893 ( .B(start_reg[137]), .A(n4377), .Z(start_in[137]) );
  ANDN U7894 ( .B(start_reg[136]), .A(n4377), .Z(start_in[136]) );
  ANDN U7895 ( .B(start_reg[135]), .A(n4377), .Z(start_in[135]) );
  ANDN U7896 ( .B(start_reg[134]), .A(n4377), .Z(start_in[134]) );
  ANDN U7897 ( .B(start_reg[133]), .A(n4377), .Z(start_in[133]) );
  ANDN U7898 ( .B(start_reg[132]), .A(n4377), .Z(start_in[132]) );
  ANDN U7899 ( .B(start_reg[131]), .A(n4377), .Z(start_in[131]) );
  ANDN U7900 ( .B(start_reg[130]), .A(n4377), .Z(start_in[130]) );
  ANDN U7901 ( .B(start_reg[12]), .A(n4377), .Z(start_in[12]) );
  ANDN U7902 ( .B(start_reg[129]), .A(n4377), .Z(start_in[129]) );
  ANDN U7903 ( .B(start_reg[128]), .A(n4377), .Z(start_in[128]) );
  ANDN U7904 ( .B(start_reg[127]), .A(n4377), .Z(start_in[127]) );
  ANDN U7905 ( .B(start_reg[126]), .A(n4377), .Z(start_in[126]) );
  ANDN U7906 ( .B(start_reg[125]), .A(n4377), .Z(start_in[125]) );
  ANDN U7907 ( .B(start_reg[124]), .A(n4377), .Z(start_in[124]) );
  ANDN U7908 ( .B(start_reg[123]), .A(n4377), .Z(start_in[123]) );
  ANDN U7909 ( .B(start_reg[122]), .A(n4377), .Z(start_in[122]) );
  ANDN U7910 ( .B(start_reg[121]), .A(n4377), .Z(start_in[121]) );
  ANDN U7911 ( .B(start_reg[120]), .A(n4377), .Z(start_in[120]) );
  ANDN U7912 ( .B(start_reg[11]), .A(n4377), .Z(start_in[11]) );
  ANDN U7913 ( .B(start_reg[119]), .A(n4377), .Z(start_in[119]) );
  ANDN U7914 ( .B(start_reg[118]), .A(n4377), .Z(start_in[118]) );
  ANDN U7915 ( .B(start_reg[117]), .A(n4377), .Z(start_in[117]) );
  ANDN U7916 ( .B(start_reg[116]), .A(n4377), .Z(start_in[116]) );
  ANDN U7917 ( .B(start_reg[115]), .A(n4377), .Z(start_in[115]) );
  ANDN U7918 ( .B(start_reg[114]), .A(n4377), .Z(start_in[114]) );
  ANDN U7919 ( .B(start_reg[113]), .A(n4377), .Z(start_in[113]) );
  ANDN U7920 ( .B(start_reg[112]), .A(n4377), .Z(start_in[112]) );
  ANDN U7921 ( .B(start_reg[111]), .A(n4377), .Z(start_in[111]) );
  ANDN U7922 ( .B(start_reg[110]), .A(n4377), .Z(start_in[110]) );
  ANDN U7923 ( .B(start_reg[10]), .A(n4377), .Z(start_in[10]) );
  ANDN U7924 ( .B(start_reg[109]), .A(n4377), .Z(start_in[109]) );
  ANDN U7925 ( .B(start_reg[108]), .A(n4377), .Z(start_in[108]) );
  ANDN U7926 ( .B(start_reg[107]), .A(n4377), .Z(start_in[107]) );
  ANDN U7927 ( .B(start_reg[106]), .A(n4377), .Z(start_in[106]) );
  ANDN U7928 ( .B(start_reg[105]), .A(n4377), .Z(start_in[105]) );
  ANDN U7929 ( .B(start_reg[104]), .A(n4377), .Z(start_in[104]) );
  ANDN U7930 ( .B(start_reg[103]), .A(n4377), .Z(start_in[103]) );
  ANDN U7931 ( .B(start_reg[102]), .A(n4377), .Z(start_in[102]) );
  ANDN U7932 ( .B(start_reg[1022]), .A(n4377), .Z(start_in[1022]) );
  ANDN U7933 ( .B(start_reg[1021]), .A(n4377), .Z(start_in[1021]) );
  ANDN U7934 ( .B(start_reg[1020]), .A(n4377), .Z(start_in[1020]) );
  ANDN U7935 ( .B(start_reg[101]), .A(n4377), .Z(start_in[101]) );
  ANDN U7936 ( .B(start_reg[1019]), .A(n4377), .Z(start_in[1019]) );
  ANDN U7937 ( .B(start_reg[1018]), .A(n4377), .Z(start_in[1018]) );
  ANDN U7938 ( .B(start_reg[1017]), .A(n4377), .Z(start_in[1017]) );
  ANDN U7939 ( .B(start_reg[1016]), .A(n4377), .Z(start_in[1016]) );
  ANDN U7940 ( .B(start_reg[1015]), .A(n4377), .Z(start_in[1015]) );
  ANDN U7941 ( .B(start_reg[1014]), .A(n4377), .Z(start_in[1014]) );
  ANDN U7942 ( .B(start_reg[1013]), .A(n4377), .Z(start_in[1013]) );
  ANDN U7943 ( .B(start_reg[1012]), .A(n4377), .Z(start_in[1012]) );
  ANDN U7944 ( .B(start_reg[1011]), .A(n4377), .Z(start_in[1011]) );
  ANDN U7945 ( .B(start_reg[1010]), .A(n4377), .Z(start_in[1010]) );
  ANDN U7946 ( .B(start_reg[100]), .A(n4377), .Z(start_in[100]) );
  ANDN U7947 ( .B(start_reg[1009]), .A(n4377), .Z(start_in[1009]) );
  ANDN U7948 ( .B(start_reg[1008]), .A(n4377), .Z(start_in[1008]) );
  ANDN U7949 ( .B(start_reg[1007]), .A(n4377), .Z(start_in[1007]) );
  ANDN U7950 ( .B(start_reg[1006]), .A(n4377), .Z(start_in[1006]) );
  ANDN U7951 ( .B(start_reg[1005]), .A(n4377), .Z(start_in[1005]) );
  ANDN U7952 ( .B(start_reg[1004]), .A(n4377), .Z(start_in[1004]) );
  ANDN U7953 ( .B(start_reg[1003]), .A(n4377), .Z(start_in[1003]) );
  ANDN U7954 ( .B(start_reg[1002]), .A(n4377), .Z(start_in[1002]) );
  ANDN U7955 ( .B(start_reg[1001]), .A(n4377), .Z(start_in[1001]) );
  ANDN U7956 ( .B(start_reg[1000]), .A(n4377), .Z(start_in[1000]) );
  OR U7957 ( .A(start_reg[0]), .B(n4377), .Z(start_in[0]) );
  NAND U7958 ( .A(n4888), .B(n4889), .Z(n3860) );
  NANDN U7959 ( .A(n3864), .B(start_reg[1023]), .Z(n4889) );
  IV U7960 ( .A(n3863), .Z(n3864) );
  NANDN U7961 ( .A(start_in[1023]), .B(mul_pow), .Z(n4888) );
  NAND U7962 ( .A(n4890), .B(n4891), .Z(n3859) );
  NAND U7963 ( .A(n4892), .B(ereg[0]), .Z(n4891) );
  NANDN U7964 ( .A(init), .B(e[0]), .Z(n4890) );
  NAND U7965 ( .A(n4893), .B(n4894), .Z(n3858) );
  NANDN U7966 ( .A(init), .B(e[1]), .Z(n4894) );
  AND U7967 ( .A(n4895), .B(n4896), .Z(n4893) );
  NAND U7968 ( .A(ereg[0]), .B(n4897), .Z(n4896) );
  NAND U7969 ( .A(n4892), .B(ereg[1]), .Z(n4895) );
  NAND U7970 ( .A(n4898), .B(n4899), .Z(n3857) );
  NANDN U7971 ( .A(init), .B(e[2]), .Z(n4899) );
  AND U7972 ( .A(n4900), .B(n4901), .Z(n4898) );
  NAND U7973 ( .A(n4897), .B(ereg[1]), .Z(n4901) );
  NAND U7974 ( .A(n4892), .B(ereg[2]), .Z(n4900) );
  NAND U7975 ( .A(n4902), .B(n4903), .Z(n3856) );
  NANDN U7976 ( .A(init), .B(e[3]), .Z(n4903) );
  AND U7977 ( .A(n4904), .B(n4905), .Z(n4902) );
  NAND U7978 ( .A(n4897), .B(ereg[2]), .Z(n4905) );
  NAND U7979 ( .A(n4892), .B(ereg[3]), .Z(n4904) );
  NAND U7980 ( .A(n4906), .B(n4907), .Z(n3855) );
  NANDN U7981 ( .A(init), .B(e[4]), .Z(n4907) );
  AND U7982 ( .A(n4908), .B(n4909), .Z(n4906) );
  NAND U7983 ( .A(n4897), .B(ereg[3]), .Z(n4909) );
  NAND U7984 ( .A(n4892), .B(ereg[4]), .Z(n4908) );
  NAND U7985 ( .A(n4910), .B(n4911), .Z(n3854) );
  NANDN U7986 ( .A(init), .B(e[5]), .Z(n4911) );
  AND U7987 ( .A(n4912), .B(n4913), .Z(n4910) );
  NAND U7988 ( .A(n4897), .B(ereg[4]), .Z(n4913) );
  NAND U7989 ( .A(n4892), .B(ereg[5]), .Z(n4912) );
  NAND U7990 ( .A(n4914), .B(n4915), .Z(n3853) );
  NANDN U7991 ( .A(init), .B(e[6]), .Z(n4915) );
  AND U7992 ( .A(n4916), .B(n4917), .Z(n4914) );
  NAND U7993 ( .A(n4897), .B(ereg[5]), .Z(n4917) );
  NAND U7994 ( .A(n4892), .B(ereg[6]), .Z(n4916) );
  NAND U7995 ( .A(n4918), .B(n4919), .Z(n3852) );
  NANDN U7996 ( .A(init), .B(e[7]), .Z(n4919) );
  AND U7997 ( .A(n4920), .B(n4921), .Z(n4918) );
  NAND U7998 ( .A(n4897), .B(ereg[6]), .Z(n4921) );
  NAND U7999 ( .A(n4892), .B(ereg[7]), .Z(n4920) );
  NAND U8000 ( .A(n4922), .B(n4923), .Z(n3851) );
  NANDN U8001 ( .A(init), .B(e[8]), .Z(n4923) );
  AND U8002 ( .A(n4924), .B(n4925), .Z(n4922) );
  NAND U8003 ( .A(n4897), .B(ereg[7]), .Z(n4925) );
  NAND U8004 ( .A(n4892), .B(ereg[8]), .Z(n4924) );
  NAND U8005 ( .A(n4926), .B(n4927), .Z(n3850) );
  NANDN U8006 ( .A(init), .B(e[9]), .Z(n4927) );
  AND U8007 ( .A(n4928), .B(n4929), .Z(n4926) );
  NAND U8008 ( .A(n4897), .B(ereg[8]), .Z(n4929) );
  NAND U8009 ( .A(n4892), .B(ereg[9]), .Z(n4928) );
  NAND U8010 ( .A(n4930), .B(n4931), .Z(n3849) );
  NANDN U8011 ( .A(init), .B(e[10]), .Z(n4931) );
  AND U8012 ( .A(n4932), .B(n4933), .Z(n4930) );
  NAND U8013 ( .A(n4897), .B(ereg[9]), .Z(n4933) );
  NAND U8014 ( .A(n4892), .B(ereg[10]), .Z(n4932) );
  NAND U8015 ( .A(n4934), .B(n4935), .Z(n3848) );
  NANDN U8016 ( .A(init), .B(e[11]), .Z(n4935) );
  AND U8017 ( .A(n4936), .B(n4937), .Z(n4934) );
  NAND U8018 ( .A(n4897), .B(ereg[10]), .Z(n4937) );
  NAND U8019 ( .A(n4892), .B(ereg[11]), .Z(n4936) );
  NAND U8020 ( .A(n4938), .B(n4939), .Z(n3847) );
  NANDN U8021 ( .A(init), .B(e[12]), .Z(n4939) );
  AND U8022 ( .A(n4940), .B(n4941), .Z(n4938) );
  NAND U8023 ( .A(n4897), .B(ereg[11]), .Z(n4941) );
  NAND U8024 ( .A(n4892), .B(ereg[12]), .Z(n4940) );
  NAND U8025 ( .A(n4942), .B(n4943), .Z(n3846) );
  NANDN U8026 ( .A(init), .B(e[13]), .Z(n4943) );
  AND U8027 ( .A(n4944), .B(n4945), .Z(n4942) );
  NAND U8028 ( .A(n4897), .B(ereg[12]), .Z(n4945) );
  NAND U8029 ( .A(n4892), .B(ereg[13]), .Z(n4944) );
  NAND U8030 ( .A(n4946), .B(n4947), .Z(n3845) );
  NANDN U8031 ( .A(init), .B(e[14]), .Z(n4947) );
  AND U8032 ( .A(n4948), .B(n4949), .Z(n4946) );
  NAND U8033 ( .A(n4897), .B(ereg[13]), .Z(n4949) );
  NAND U8034 ( .A(n4892), .B(ereg[14]), .Z(n4948) );
  NAND U8035 ( .A(n4950), .B(n4951), .Z(n3844) );
  NANDN U8036 ( .A(init), .B(e[15]), .Z(n4951) );
  AND U8037 ( .A(n4952), .B(n4953), .Z(n4950) );
  NAND U8038 ( .A(n4897), .B(ereg[14]), .Z(n4953) );
  NAND U8039 ( .A(n4892), .B(ereg[15]), .Z(n4952) );
  NAND U8040 ( .A(n4954), .B(n4955), .Z(n3843) );
  NANDN U8041 ( .A(init), .B(e[16]), .Z(n4955) );
  AND U8042 ( .A(n4956), .B(n4957), .Z(n4954) );
  NAND U8043 ( .A(n4897), .B(ereg[15]), .Z(n4957) );
  NAND U8044 ( .A(n4892), .B(ereg[16]), .Z(n4956) );
  NAND U8045 ( .A(n4958), .B(n4959), .Z(n3842) );
  NANDN U8046 ( .A(init), .B(e[17]), .Z(n4959) );
  AND U8047 ( .A(n4960), .B(n4961), .Z(n4958) );
  NAND U8048 ( .A(n4897), .B(ereg[16]), .Z(n4961) );
  NAND U8049 ( .A(n4892), .B(ereg[17]), .Z(n4960) );
  NAND U8050 ( .A(n4962), .B(n4963), .Z(n3841) );
  NANDN U8051 ( .A(init), .B(e[18]), .Z(n4963) );
  AND U8052 ( .A(n4964), .B(n4965), .Z(n4962) );
  NAND U8053 ( .A(n4897), .B(ereg[17]), .Z(n4965) );
  NAND U8054 ( .A(n4892), .B(ereg[18]), .Z(n4964) );
  NAND U8055 ( .A(n4966), .B(n4967), .Z(n3840) );
  NANDN U8056 ( .A(init), .B(e[19]), .Z(n4967) );
  AND U8057 ( .A(n4968), .B(n4969), .Z(n4966) );
  NAND U8058 ( .A(n4897), .B(ereg[18]), .Z(n4969) );
  NAND U8059 ( .A(n4892), .B(ereg[19]), .Z(n4968) );
  NAND U8060 ( .A(n4970), .B(n4971), .Z(n3839) );
  NANDN U8061 ( .A(init), .B(e[20]), .Z(n4971) );
  AND U8062 ( .A(n4972), .B(n4973), .Z(n4970) );
  NAND U8063 ( .A(n4897), .B(ereg[19]), .Z(n4973) );
  NAND U8064 ( .A(n4892), .B(ereg[20]), .Z(n4972) );
  NAND U8065 ( .A(n4974), .B(n4975), .Z(n3838) );
  NANDN U8066 ( .A(init), .B(e[21]), .Z(n4975) );
  AND U8067 ( .A(n4976), .B(n4977), .Z(n4974) );
  NAND U8068 ( .A(n4897), .B(ereg[20]), .Z(n4977) );
  NAND U8069 ( .A(n4892), .B(ereg[21]), .Z(n4976) );
  NAND U8070 ( .A(n4978), .B(n4979), .Z(n3837) );
  NANDN U8071 ( .A(init), .B(e[22]), .Z(n4979) );
  AND U8072 ( .A(n4980), .B(n4981), .Z(n4978) );
  NAND U8073 ( .A(n4897), .B(ereg[21]), .Z(n4981) );
  NAND U8074 ( .A(n4892), .B(ereg[22]), .Z(n4980) );
  NAND U8075 ( .A(n4982), .B(n4983), .Z(n3836) );
  NANDN U8076 ( .A(init), .B(e[23]), .Z(n4983) );
  AND U8077 ( .A(n4984), .B(n4985), .Z(n4982) );
  NAND U8078 ( .A(n4897), .B(ereg[22]), .Z(n4985) );
  NAND U8079 ( .A(n4892), .B(ereg[23]), .Z(n4984) );
  NAND U8080 ( .A(n4986), .B(n4987), .Z(n3835) );
  NANDN U8081 ( .A(init), .B(e[24]), .Z(n4987) );
  AND U8082 ( .A(n4988), .B(n4989), .Z(n4986) );
  NAND U8083 ( .A(n4897), .B(ereg[23]), .Z(n4989) );
  NAND U8084 ( .A(n4892), .B(ereg[24]), .Z(n4988) );
  NAND U8085 ( .A(n4990), .B(n4991), .Z(n3834) );
  NANDN U8086 ( .A(init), .B(e[25]), .Z(n4991) );
  AND U8087 ( .A(n4992), .B(n4993), .Z(n4990) );
  NAND U8088 ( .A(n4897), .B(ereg[24]), .Z(n4993) );
  NAND U8089 ( .A(n4892), .B(ereg[25]), .Z(n4992) );
  NAND U8090 ( .A(n4994), .B(n4995), .Z(n3833) );
  NANDN U8091 ( .A(init), .B(e[26]), .Z(n4995) );
  AND U8092 ( .A(n4996), .B(n4997), .Z(n4994) );
  NAND U8093 ( .A(n4897), .B(ereg[25]), .Z(n4997) );
  NAND U8094 ( .A(n4892), .B(ereg[26]), .Z(n4996) );
  NAND U8095 ( .A(n4998), .B(n4999), .Z(n3832) );
  NANDN U8096 ( .A(init), .B(e[27]), .Z(n4999) );
  AND U8097 ( .A(n5000), .B(n5001), .Z(n4998) );
  NAND U8098 ( .A(n4897), .B(ereg[26]), .Z(n5001) );
  NAND U8099 ( .A(n4892), .B(ereg[27]), .Z(n5000) );
  NAND U8100 ( .A(n5002), .B(n5003), .Z(n3831) );
  NANDN U8101 ( .A(init), .B(e[28]), .Z(n5003) );
  AND U8102 ( .A(n5004), .B(n5005), .Z(n5002) );
  NAND U8103 ( .A(n4897), .B(ereg[27]), .Z(n5005) );
  NAND U8104 ( .A(n4892), .B(ereg[28]), .Z(n5004) );
  NAND U8105 ( .A(n5006), .B(n5007), .Z(n3830) );
  NANDN U8106 ( .A(init), .B(e[29]), .Z(n5007) );
  AND U8107 ( .A(n5008), .B(n5009), .Z(n5006) );
  NAND U8108 ( .A(n4897), .B(ereg[28]), .Z(n5009) );
  NAND U8109 ( .A(n4892), .B(ereg[29]), .Z(n5008) );
  NAND U8110 ( .A(n5010), .B(n5011), .Z(n3829) );
  NANDN U8111 ( .A(init), .B(e[30]), .Z(n5011) );
  AND U8112 ( .A(n5012), .B(n5013), .Z(n5010) );
  NAND U8113 ( .A(n4897), .B(ereg[29]), .Z(n5013) );
  NAND U8114 ( .A(n4892), .B(ereg[30]), .Z(n5012) );
  NAND U8115 ( .A(n5014), .B(n5015), .Z(n3828) );
  NANDN U8116 ( .A(init), .B(e[31]), .Z(n5015) );
  AND U8117 ( .A(n5016), .B(n5017), .Z(n5014) );
  NAND U8118 ( .A(n4897), .B(ereg[30]), .Z(n5017) );
  NAND U8119 ( .A(n4892), .B(ereg[31]), .Z(n5016) );
  NAND U8120 ( .A(n5018), .B(n5019), .Z(n3827) );
  NANDN U8121 ( .A(init), .B(e[32]), .Z(n5019) );
  AND U8122 ( .A(n5020), .B(n5021), .Z(n5018) );
  NAND U8123 ( .A(n4897), .B(ereg[31]), .Z(n5021) );
  NAND U8124 ( .A(n4892), .B(ereg[32]), .Z(n5020) );
  NAND U8125 ( .A(n5022), .B(n5023), .Z(n3826) );
  NANDN U8126 ( .A(init), .B(e[33]), .Z(n5023) );
  AND U8127 ( .A(n5024), .B(n5025), .Z(n5022) );
  NAND U8128 ( .A(n4897), .B(ereg[32]), .Z(n5025) );
  NAND U8129 ( .A(n4892), .B(ereg[33]), .Z(n5024) );
  NAND U8130 ( .A(n5026), .B(n5027), .Z(n3825) );
  NANDN U8131 ( .A(init), .B(e[34]), .Z(n5027) );
  AND U8132 ( .A(n5028), .B(n5029), .Z(n5026) );
  NAND U8133 ( .A(n4897), .B(ereg[33]), .Z(n5029) );
  NAND U8134 ( .A(n4892), .B(ereg[34]), .Z(n5028) );
  NAND U8135 ( .A(n5030), .B(n5031), .Z(n3824) );
  NANDN U8136 ( .A(init), .B(e[35]), .Z(n5031) );
  AND U8137 ( .A(n5032), .B(n5033), .Z(n5030) );
  NAND U8138 ( .A(n4897), .B(ereg[34]), .Z(n5033) );
  NAND U8139 ( .A(n4892), .B(ereg[35]), .Z(n5032) );
  NAND U8140 ( .A(n5034), .B(n5035), .Z(n3823) );
  NANDN U8141 ( .A(init), .B(e[36]), .Z(n5035) );
  AND U8142 ( .A(n5036), .B(n5037), .Z(n5034) );
  NAND U8143 ( .A(n4897), .B(ereg[35]), .Z(n5037) );
  NAND U8144 ( .A(n4892), .B(ereg[36]), .Z(n5036) );
  NAND U8145 ( .A(n5038), .B(n5039), .Z(n3822) );
  NANDN U8146 ( .A(init), .B(e[37]), .Z(n5039) );
  AND U8147 ( .A(n5040), .B(n5041), .Z(n5038) );
  NAND U8148 ( .A(n4897), .B(ereg[36]), .Z(n5041) );
  NAND U8149 ( .A(n4892), .B(ereg[37]), .Z(n5040) );
  NAND U8150 ( .A(n5042), .B(n5043), .Z(n3821) );
  NANDN U8151 ( .A(init), .B(e[38]), .Z(n5043) );
  AND U8152 ( .A(n5044), .B(n5045), .Z(n5042) );
  NAND U8153 ( .A(n4897), .B(ereg[37]), .Z(n5045) );
  NAND U8154 ( .A(n4892), .B(ereg[38]), .Z(n5044) );
  NAND U8155 ( .A(n5046), .B(n5047), .Z(n3820) );
  NANDN U8156 ( .A(init), .B(e[39]), .Z(n5047) );
  AND U8157 ( .A(n5048), .B(n5049), .Z(n5046) );
  NAND U8158 ( .A(n4897), .B(ereg[38]), .Z(n5049) );
  NAND U8159 ( .A(n4892), .B(ereg[39]), .Z(n5048) );
  NAND U8160 ( .A(n5050), .B(n5051), .Z(n3819) );
  NANDN U8161 ( .A(init), .B(e[40]), .Z(n5051) );
  AND U8162 ( .A(n5052), .B(n5053), .Z(n5050) );
  NAND U8163 ( .A(n4897), .B(ereg[39]), .Z(n5053) );
  NAND U8164 ( .A(n4892), .B(ereg[40]), .Z(n5052) );
  NAND U8165 ( .A(n5054), .B(n5055), .Z(n3818) );
  NANDN U8166 ( .A(init), .B(e[41]), .Z(n5055) );
  AND U8167 ( .A(n5056), .B(n5057), .Z(n5054) );
  NAND U8168 ( .A(n4897), .B(ereg[40]), .Z(n5057) );
  NAND U8169 ( .A(n4892), .B(ereg[41]), .Z(n5056) );
  NAND U8170 ( .A(n5058), .B(n5059), .Z(n3817) );
  NANDN U8171 ( .A(init), .B(e[42]), .Z(n5059) );
  AND U8172 ( .A(n5060), .B(n5061), .Z(n5058) );
  NAND U8173 ( .A(n4897), .B(ereg[41]), .Z(n5061) );
  NAND U8174 ( .A(n4892), .B(ereg[42]), .Z(n5060) );
  NAND U8175 ( .A(n5062), .B(n5063), .Z(n3816) );
  NANDN U8176 ( .A(init), .B(e[43]), .Z(n5063) );
  AND U8177 ( .A(n5064), .B(n5065), .Z(n5062) );
  NAND U8178 ( .A(n4897), .B(ereg[42]), .Z(n5065) );
  NAND U8179 ( .A(n4892), .B(ereg[43]), .Z(n5064) );
  NAND U8180 ( .A(n5066), .B(n5067), .Z(n3815) );
  NANDN U8181 ( .A(init), .B(e[44]), .Z(n5067) );
  AND U8182 ( .A(n5068), .B(n5069), .Z(n5066) );
  NAND U8183 ( .A(n4897), .B(ereg[43]), .Z(n5069) );
  NAND U8184 ( .A(n4892), .B(ereg[44]), .Z(n5068) );
  NAND U8185 ( .A(n5070), .B(n5071), .Z(n3814) );
  NANDN U8186 ( .A(init), .B(e[45]), .Z(n5071) );
  AND U8187 ( .A(n5072), .B(n5073), .Z(n5070) );
  NAND U8188 ( .A(n4897), .B(ereg[44]), .Z(n5073) );
  NAND U8189 ( .A(n4892), .B(ereg[45]), .Z(n5072) );
  NAND U8190 ( .A(n5074), .B(n5075), .Z(n3813) );
  NANDN U8191 ( .A(init), .B(e[46]), .Z(n5075) );
  AND U8192 ( .A(n5076), .B(n5077), .Z(n5074) );
  NAND U8193 ( .A(n4897), .B(ereg[45]), .Z(n5077) );
  NAND U8194 ( .A(n4892), .B(ereg[46]), .Z(n5076) );
  NAND U8195 ( .A(n5078), .B(n5079), .Z(n3812) );
  NANDN U8196 ( .A(init), .B(e[47]), .Z(n5079) );
  AND U8197 ( .A(n5080), .B(n5081), .Z(n5078) );
  NAND U8198 ( .A(n4897), .B(ereg[46]), .Z(n5081) );
  NAND U8199 ( .A(n4892), .B(ereg[47]), .Z(n5080) );
  NAND U8200 ( .A(n5082), .B(n5083), .Z(n3811) );
  NANDN U8201 ( .A(init), .B(e[48]), .Z(n5083) );
  AND U8202 ( .A(n5084), .B(n5085), .Z(n5082) );
  NAND U8203 ( .A(n4897), .B(ereg[47]), .Z(n5085) );
  NAND U8204 ( .A(n4892), .B(ereg[48]), .Z(n5084) );
  NAND U8205 ( .A(n5086), .B(n5087), .Z(n3810) );
  NANDN U8206 ( .A(init), .B(e[49]), .Z(n5087) );
  AND U8207 ( .A(n5088), .B(n5089), .Z(n5086) );
  NAND U8208 ( .A(n4897), .B(ereg[48]), .Z(n5089) );
  NAND U8209 ( .A(n4892), .B(ereg[49]), .Z(n5088) );
  NAND U8210 ( .A(n5090), .B(n5091), .Z(n3809) );
  NANDN U8211 ( .A(init), .B(e[50]), .Z(n5091) );
  AND U8212 ( .A(n5092), .B(n5093), .Z(n5090) );
  NAND U8213 ( .A(n4897), .B(ereg[49]), .Z(n5093) );
  NAND U8214 ( .A(n4892), .B(ereg[50]), .Z(n5092) );
  NAND U8215 ( .A(n5094), .B(n5095), .Z(n3808) );
  NANDN U8216 ( .A(init), .B(e[51]), .Z(n5095) );
  AND U8217 ( .A(n5096), .B(n5097), .Z(n5094) );
  NAND U8218 ( .A(n4897), .B(ereg[50]), .Z(n5097) );
  NAND U8219 ( .A(n4892), .B(ereg[51]), .Z(n5096) );
  NAND U8220 ( .A(n5098), .B(n5099), .Z(n3807) );
  NANDN U8221 ( .A(init), .B(e[52]), .Z(n5099) );
  AND U8222 ( .A(n5100), .B(n5101), .Z(n5098) );
  NAND U8223 ( .A(n4897), .B(ereg[51]), .Z(n5101) );
  NAND U8224 ( .A(n4892), .B(ereg[52]), .Z(n5100) );
  NAND U8225 ( .A(n5102), .B(n5103), .Z(n3806) );
  NANDN U8226 ( .A(init), .B(e[53]), .Z(n5103) );
  AND U8227 ( .A(n5104), .B(n5105), .Z(n5102) );
  NAND U8228 ( .A(n4897), .B(ereg[52]), .Z(n5105) );
  NAND U8229 ( .A(n4892), .B(ereg[53]), .Z(n5104) );
  NAND U8230 ( .A(n5106), .B(n5107), .Z(n3805) );
  NANDN U8231 ( .A(init), .B(e[54]), .Z(n5107) );
  AND U8232 ( .A(n5108), .B(n5109), .Z(n5106) );
  NAND U8233 ( .A(n4897), .B(ereg[53]), .Z(n5109) );
  NAND U8234 ( .A(n4892), .B(ereg[54]), .Z(n5108) );
  NAND U8235 ( .A(n5110), .B(n5111), .Z(n3804) );
  NANDN U8236 ( .A(init), .B(e[55]), .Z(n5111) );
  AND U8237 ( .A(n5112), .B(n5113), .Z(n5110) );
  NAND U8238 ( .A(n4897), .B(ereg[54]), .Z(n5113) );
  NAND U8239 ( .A(n4892), .B(ereg[55]), .Z(n5112) );
  NAND U8240 ( .A(n5114), .B(n5115), .Z(n3803) );
  NANDN U8241 ( .A(init), .B(e[56]), .Z(n5115) );
  AND U8242 ( .A(n5116), .B(n5117), .Z(n5114) );
  NAND U8243 ( .A(n4897), .B(ereg[55]), .Z(n5117) );
  NAND U8244 ( .A(n4892), .B(ereg[56]), .Z(n5116) );
  NAND U8245 ( .A(n5118), .B(n5119), .Z(n3802) );
  NANDN U8246 ( .A(init), .B(e[57]), .Z(n5119) );
  AND U8247 ( .A(n5120), .B(n5121), .Z(n5118) );
  NAND U8248 ( .A(n4897), .B(ereg[56]), .Z(n5121) );
  NAND U8249 ( .A(n4892), .B(ereg[57]), .Z(n5120) );
  NAND U8250 ( .A(n5122), .B(n5123), .Z(n3801) );
  NANDN U8251 ( .A(init), .B(e[58]), .Z(n5123) );
  AND U8252 ( .A(n5124), .B(n5125), .Z(n5122) );
  NAND U8253 ( .A(n4897), .B(ereg[57]), .Z(n5125) );
  NAND U8254 ( .A(n4892), .B(ereg[58]), .Z(n5124) );
  NAND U8255 ( .A(n5126), .B(n5127), .Z(n3800) );
  NANDN U8256 ( .A(init), .B(e[59]), .Z(n5127) );
  AND U8257 ( .A(n5128), .B(n5129), .Z(n5126) );
  NAND U8258 ( .A(n4897), .B(ereg[58]), .Z(n5129) );
  NAND U8259 ( .A(n4892), .B(ereg[59]), .Z(n5128) );
  NAND U8260 ( .A(n5130), .B(n5131), .Z(n3799) );
  NANDN U8261 ( .A(init), .B(e[60]), .Z(n5131) );
  AND U8262 ( .A(n5132), .B(n5133), .Z(n5130) );
  NAND U8263 ( .A(n4897), .B(ereg[59]), .Z(n5133) );
  NAND U8264 ( .A(n4892), .B(ereg[60]), .Z(n5132) );
  NAND U8265 ( .A(n5134), .B(n5135), .Z(n3798) );
  NANDN U8266 ( .A(init), .B(e[61]), .Z(n5135) );
  AND U8267 ( .A(n5136), .B(n5137), .Z(n5134) );
  NAND U8268 ( .A(n4897), .B(ereg[60]), .Z(n5137) );
  NAND U8269 ( .A(n4892), .B(ereg[61]), .Z(n5136) );
  NAND U8270 ( .A(n5138), .B(n5139), .Z(n3797) );
  NANDN U8271 ( .A(init), .B(e[62]), .Z(n5139) );
  AND U8272 ( .A(n5140), .B(n5141), .Z(n5138) );
  NAND U8273 ( .A(n4897), .B(ereg[61]), .Z(n5141) );
  NAND U8274 ( .A(n4892), .B(ereg[62]), .Z(n5140) );
  NAND U8275 ( .A(n5142), .B(n5143), .Z(n3796) );
  NANDN U8276 ( .A(init), .B(e[63]), .Z(n5143) );
  AND U8277 ( .A(n5144), .B(n5145), .Z(n5142) );
  NAND U8278 ( .A(n4897), .B(ereg[62]), .Z(n5145) );
  NAND U8279 ( .A(n4892), .B(ereg[63]), .Z(n5144) );
  NAND U8280 ( .A(n5146), .B(n5147), .Z(n3795) );
  NANDN U8281 ( .A(init), .B(e[64]), .Z(n5147) );
  AND U8282 ( .A(n5148), .B(n5149), .Z(n5146) );
  NAND U8283 ( .A(n4897), .B(ereg[63]), .Z(n5149) );
  NAND U8284 ( .A(n4892), .B(ereg[64]), .Z(n5148) );
  NAND U8285 ( .A(n5150), .B(n5151), .Z(n3794) );
  NANDN U8286 ( .A(init), .B(e[65]), .Z(n5151) );
  AND U8287 ( .A(n5152), .B(n5153), .Z(n5150) );
  NAND U8288 ( .A(n4897), .B(ereg[64]), .Z(n5153) );
  NAND U8289 ( .A(n4892), .B(ereg[65]), .Z(n5152) );
  NAND U8290 ( .A(n5154), .B(n5155), .Z(n3793) );
  NANDN U8291 ( .A(init), .B(e[66]), .Z(n5155) );
  AND U8292 ( .A(n5156), .B(n5157), .Z(n5154) );
  NAND U8293 ( .A(n4897), .B(ereg[65]), .Z(n5157) );
  NAND U8294 ( .A(n4892), .B(ereg[66]), .Z(n5156) );
  NAND U8295 ( .A(n5158), .B(n5159), .Z(n3792) );
  NANDN U8296 ( .A(init), .B(e[67]), .Z(n5159) );
  AND U8297 ( .A(n5160), .B(n5161), .Z(n5158) );
  NAND U8298 ( .A(n4897), .B(ereg[66]), .Z(n5161) );
  NAND U8299 ( .A(n4892), .B(ereg[67]), .Z(n5160) );
  NAND U8300 ( .A(n5162), .B(n5163), .Z(n3791) );
  NANDN U8301 ( .A(init), .B(e[68]), .Z(n5163) );
  AND U8302 ( .A(n5164), .B(n5165), .Z(n5162) );
  NAND U8303 ( .A(n4897), .B(ereg[67]), .Z(n5165) );
  NAND U8304 ( .A(n4892), .B(ereg[68]), .Z(n5164) );
  NAND U8305 ( .A(n5166), .B(n5167), .Z(n3790) );
  NANDN U8306 ( .A(init), .B(e[69]), .Z(n5167) );
  AND U8307 ( .A(n5168), .B(n5169), .Z(n5166) );
  NAND U8308 ( .A(n4897), .B(ereg[68]), .Z(n5169) );
  NAND U8309 ( .A(n4892), .B(ereg[69]), .Z(n5168) );
  NAND U8310 ( .A(n5170), .B(n5171), .Z(n3789) );
  NANDN U8311 ( .A(init), .B(e[70]), .Z(n5171) );
  AND U8312 ( .A(n5172), .B(n5173), .Z(n5170) );
  NAND U8313 ( .A(n4897), .B(ereg[69]), .Z(n5173) );
  NAND U8314 ( .A(n4892), .B(ereg[70]), .Z(n5172) );
  NAND U8315 ( .A(n5174), .B(n5175), .Z(n3788) );
  NANDN U8316 ( .A(init), .B(e[71]), .Z(n5175) );
  AND U8317 ( .A(n5176), .B(n5177), .Z(n5174) );
  NAND U8318 ( .A(n4897), .B(ereg[70]), .Z(n5177) );
  NAND U8319 ( .A(n4892), .B(ereg[71]), .Z(n5176) );
  NAND U8320 ( .A(n5178), .B(n5179), .Z(n3787) );
  NANDN U8321 ( .A(init), .B(e[72]), .Z(n5179) );
  AND U8322 ( .A(n5180), .B(n5181), .Z(n5178) );
  NAND U8323 ( .A(n4897), .B(ereg[71]), .Z(n5181) );
  NAND U8324 ( .A(n4892), .B(ereg[72]), .Z(n5180) );
  NAND U8325 ( .A(n5182), .B(n5183), .Z(n3786) );
  NANDN U8326 ( .A(init), .B(e[73]), .Z(n5183) );
  AND U8327 ( .A(n5184), .B(n5185), .Z(n5182) );
  NAND U8328 ( .A(n4897), .B(ereg[72]), .Z(n5185) );
  NAND U8329 ( .A(n4892), .B(ereg[73]), .Z(n5184) );
  NAND U8330 ( .A(n5186), .B(n5187), .Z(n3785) );
  NANDN U8331 ( .A(init), .B(e[74]), .Z(n5187) );
  AND U8332 ( .A(n5188), .B(n5189), .Z(n5186) );
  NAND U8333 ( .A(n4897), .B(ereg[73]), .Z(n5189) );
  NAND U8334 ( .A(n4892), .B(ereg[74]), .Z(n5188) );
  NAND U8335 ( .A(n5190), .B(n5191), .Z(n3784) );
  NANDN U8336 ( .A(init), .B(e[75]), .Z(n5191) );
  AND U8337 ( .A(n5192), .B(n5193), .Z(n5190) );
  NAND U8338 ( .A(n4897), .B(ereg[74]), .Z(n5193) );
  NAND U8339 ( .A(n4892), .B(ereg[75]), .Z(n5192) );
  NAND U8340 ( .A(n5194), .B(n5195), .Z(n3783) );
  NANDN U8341 ( .A(init), .B(e[76]), .Z(n5195) );
  AND U8342 ( .A(n5196), .B(n5197), .Z(n5194) );
  NAND U8343 ( .A(n4897), .B(ereg[75]), .Z(n5197) );
  NAND U8344 ( .A(n4892), .B(ereg[76]), .Z(n5196) );
  NAND U8345 ( .A(n5198), .B(n5199), .Z(n3782) );
  NANDN U8346 ( .A(init), .B(e[77]), .Z(n5199) );
  AND U8347 ( .A(n5200), .B(n5201), .Z(n5198) );
  NAND U8348 ( .A(n4897), .B(ereg[76]), .Z(n5201) );
  NAND U8349 ( .A(n4892), .B(ereg[77]), .Z(n5200) );
  NAND U8350 ( .A(n5202), .B(n5203), .Z(n3781) );
  NANDN U8351 ( .A(init), .B(e[78]), .Z(n5203) );
  AND U8352 ( .A(n5204), .B(n5205), .Z(n5202) );
  NAND U8353 ( .A(n4897), .B(ereg[77]), .Z(n5205) );
  NAND U8354 ( .A(n4892), .B(ereg[78]), .Z(n5204) );
  NAND U8355 ( .A(n5206), .B(n5207), .Z(n3780) );
  NANDN U8356 ( .A(init), .B(e[79]), .Z(n5207) );
  AND U8357 ( .A(n5208), .B(n5209), .Z(n5206) );
  NAND U8358 ( .A(n4897), .B(ereg[78]), .Z(n5209) );
  NAND U8359 ( .A(n4892), .B(ereg[79]), .Z(n5208) );
  NAND U8360 ( .A(n5210), .B(n5211), .Z(n3779) );
  NANDN U8361 ( .A(init), .B(e[80]), .Z(n5211) );
  AND U8362 ( .A(n5212), .B(n5213), .Z(n5210) );
  NAND U8363 ( .A(n4897), .B(ereg[79]), .Z(n5213) );
  NAND U8364 ( .A(n4892), .B(ereg[80]), .Z(n5212) );
  NAND U8365 ( .A(n5214), .B(n5215), .Z(n3778) );
  NANDN U8366 ( .A(init), .B(e[81]), .Z(n5215) );
  AND U8367 ( .A(n5216), .B(n5217), .Z(n5214) );
  NAND U8368 ( .A(n4897), .B(ereg[80]), .Z(n5217) );
  NAND U8369 ( .A(n4892), .B(ereg[81]), .Z(n5216) );
  NAND U8370 ( .A(n5218), .B(n5219), .Z(n3777) );
  NANDN U8371 ( .A(init), .B(e[82]), .Z(n5219) );
  AND U8372 ( .A(n5220), .B(n5221), .Z(n5218) );
  NAND U8373 ( .A(n4897), .B(ereg[81]), .Z(n5221) );
  NAND U8374 ( .A(n4892), .B(ereg[82]), .Z(n5220) );
  NAND U8375 ( .A(n5222), .B(n5223), .Z(n3776) );
  NANDN U8376 ( .A(init), .B(e[83]), .Z(n5223) );
  AND U8377 ( .A(n5224), .B(n5225), .Z(n5222) );
  NAND U8378 ( .A(n4897), .B(ereg[82]), .Z(n5225) );
  NAND U8379 ( .A(n4892), .B(ereg[83]), .Z(n5224) );
  NAND U8380 ( .A(n5226), .B(n5227), .Z(n3775) );
  NANDN U8381 ( .A(init), .B(e[84]), .Z(n5227) );
  AND U8382 ( .A(n5228), .B(n5229), .Z(n5226) );
  NAND U8383 ( .A(n4897), .B(ereg[83]), .Z(n5229) );
  NAND U8384 ( .A(n4892), .B(ereg[84]), .Z(n5228) );
  NAND U8385 ( .A(n5230), .B(n5231), .Z(n3774) );
  NANDN U8386 ( .A(init), .B(e[85]), .Z(n5231) );
  AND U8387 ( .A(n5232), .B(n5233), .Z(n5230) );
  NAND U8388 ( .A(n4897), .B(ereg[84]), .Z(n5233) );
  NAND U8389 ( .A(n4892), .B(ereg[85]), .Z(n5232) );
  NAND U8390 ( .A(n5234), .B(n5235), .Z(n3773) );
  NANDN U8391 ( .A(init), .B(e[86]), .Z(n5235) );
  AND U8392 ( .A(n5236), .B(n5237), .Z(n5234) );
  NAND U8393 ( .A(n4897), .B(ereg[85]), .Z(n5237) );
  NAND U8394 ( .A(n4892), .B(ereg[86]), .Z(n5236) );
  NAND U8395 ( .A(n5238), .B(n5239), .Z(n3772) );
  NANDN U8396 ( .A(init), .B(e[87]), .Z(n5239) );
  AND U8397 ( .A(n5240), .B(n5241), .Z(n5238) );
  NAND U8398 ( .A(n4897), .B(ereg[86]), .Z(n5241) );
  NAND U8399 ( .A(n4892), .B(ereg[87]), .Z(n5240) );
  NAND U8400 ( .A(n5242), .B(n5243), .Z(n3771) );
  NANDN U8401 ( .A(init), .B(e[88]), .Z(n5243) );
  AND U8402 ( .A(n5244), .B(n5245), .Z(n5242) );
  NAND U8403 ( .A(n4897), .B(ereg[87]), .Z(n5245) );
  NAND U8404 ( .A(n4892), .B(ereg[88]), .Z(n5244) );
  NAND U8405 ( .A(n5246), .B(n5247), .Z(n3770) );
  NANDN U8406 ( .A(init), .B(e[89]), .Z(n5247) );
  AND U8407 ( .A(n5248), .B(n5249), .Z(n5246) );
  NAND U8408 ( .A(n4897), .B(ereg[88]), .Z(n5249) );
  NAND U8409 ( .A(n4892), .B(ereg[89]), .Z(n5248) );
  NAND U8410 ( .A(n5250), .B(n5251), .Z(n3769) );
  NANDN U8411 ( .A(init), .B(e[90]), .Z(n5251) );
  AND U8412 ( .A(n5252), .B(n5253), .Z(n5250) );
  NAND U8413 ( .A(n4897), .B(ereg[89]), .Z(n5253) );
  NAND U8414 ( .A(n4892), .B(ereg[90]), .Z(n5252) );
  NAND U8415 ( .A(n5254), .B(n5255), .Z(n3768) );
  NANDN U8416 ( .A(init), .B(e[91]), .Z(n5255) );
  AND U8417 ( .A(n5256), .B(n5257), .Z(n5254) );
  NAND U8418 ( .A(n4897), .B(ereg[90]), .Z(n5257) );
  NAND U8419 ( .A(n4892), .B(ereg[91]), .Z(n5256) );
  NAND U8420 ( .A(n5258), .B(n5259), .Z(n3767) );
  NANDN U8421 ( .A(init), .B(e[92]), .Z(n5259) );
  AND U8422 ( .A(n5260), .B(n5261), .Z(n5258) );
  NAND U8423 ( .A(n4897), .B(ereg[91]), .Z(n5261) );
  NAND U8424 ( .A(n4892), .B(ereg[92]), .Z(n5260) );
  NAND U8425 ( .A(n5262), .B(n5263), .Z(n3766) );
  NANDN U8426 ( .A(init), .B(e[93]), .Z(n5263) );
  AND U8427 ( .A(n5264), .B(n5265), .Z(n5262) );
  NAND U8428 ( .A(n4897), .B(ereg[92]), .Z(n5265) );
  NAND U8429 ( .A(n4892), .B(ereg[93]), .Z(n5264) );
  NAND U8430 ( .A(n5266), .B(n5267), .Z(n3765) );
  NANDN U8431 ( .A(init), .B(e[94]), .Z(n5267) );
  AND U8432 ( .A(n5268), .B(n5269), .Z(n5266) );
  NAND U8433 ( .A(n4897), .B(ereg[93]), .Z(n5269) );
  NAND U8434 ( .A(n4892), .B(ereg[94]), .Z(n5268) );
  NAND U8435 ( .A(n5270), .B(n5271), .Z(n3764) );
  NANDN U8436 ( .A(init), .B(e[95]), .Z(n5271) );
  AND U8437 ( .A(n5272), .B(n5273), .Z(n5270) );
  NAND U8438 ( .A(n4897), .B(ereg[94]), .Z(n5273) );
  NAND U8439 ( .A(n4892), .B(ereg[95]), .Z(n5272) );
  NAND U8440 ( .A(n5274), .B(n5275), .Z(n3763) );
  NANDN U8441 ( .A(init), .B(e[96]), .Z(n5275) );
  AND U8442 ( .A(n5276), .B(n5277), .Z(n5274) );
  NAND U8443 ( .A(n4897), .B(ereg[95]), .Z(n5277) );
  NAND U8444 ( .A(n4892), .B(ereg[96]), .Z(n5276) );
  NAND U8445 ( .A(n5278), .B(n5279), .Z(n3762) );
  NANDN U8446 ( .A(init), .B(e[97]), .Z(n5279) );
  AND U8447 ( .A(n5280), .B(n5281), .Z(n5278) );
  NAND U8448 ( .A(n4897), .B(ereg[96]), .Z(n5281) );
  NAND U8449 ( .A(n4892), .B(ereg[97]), .Z(n5280) );
  NAND U8450 ( .A(n5282), .B(n5283), .Z(n3761) );
  NANDN U8451 ( .A(init), .B(e[98]), .Z(n5283) );
  AND U8452 ( .A(n5284), .B(n5285), .Z(n5282) );
  NAND U8453 ( .A(n4897), .B(ereg[97]), .Z(n5285) );
  NAND U8454 ( .A(n4892), .B(ereg[98]), .Z(n5284) );
  NAND U8455 ( .A(n5286), .B(n5287), .Z(n3760) );
  NANDN U8456 ( .A(init), .B(e[99]), .Z(n5287) );
  AND U8457 ( .A(n5288), .B(n5289), .Z(n5286) );
  NAND U8458 ( .A(n4897), .B(ereg[98]), .Z(n5289) );
  NAND U8459 ( .A(n4892), .B(ereg[99]), .Z(n5288) );
  NAND U8460 ( .A(n5290), .B(n5291), .Z(n3759) );
  NANDN U8461 ( .A(init), .B(e[100]), .Z(n5291) );
  AND U8462 ( .A(n5292), .B(n5293), .Z(n5290) );
  NAND U8463 ( .A(n4897), .B(ereg[99]), .Z(n5293) );
  NAND U8464 ( .A(n4892), .B(ereg[100]), .Z(n5292) );
  NAND U8465 ( .A(n5294), .B(n5295), .Z(n3758) );
  NANDN U8466 ( .A(init), .B(e[101]), .Z(n5295) );
  AND U8467 ( .A(n5296), .B(n5297), .Z(n5294) );
  NAND U8468 ( .A(n4897), .B(ereg[100]), .Z(n5297) );
  NAND U8469 ( .A(n4892), .B(ereg[101]), .Z(n5296) );
  NAND U8470 ( .A(n5298), .B(n5299), .Z(n3757) );
  NANDN U8471 ( .A(init), .B(e[102]), .Z(n5299) );
  AND U8472 ( .A(n5300), .B(n5301), .Z(n5298) );
  NAND U8473 ( .A(n4897), .B(ereg[101]), .Z(n5301) );
  NAND U8474 ( .A(n4892), .B(ereg[102]), .Z(n5300) );
  NAND U8475 ( .A(n5302), .B(n5303), .Z(n3756) );
  NANDN U8476 ( .A(init), .B(e[103]), .Z(n5303) );
  AND U8477 ( .A(n5304), .B(n5305), .Z(n5302) );
  NAND U8478 ( .A(n4897), .B(ereg[102]), .Z(n5305) );
  NAND U8479 ( .A(n4892), .B(ereg[103]), .Z(n5304) );
  NAND U8480 ( .A(n5306), .B(n5307), .Z(n3755) );
  NANDN U8481 ( .A(init), .B(e[104]), .Z(n5307) );
  AND U8482 ( .A(n5308), .B(n5309), .Z(n5306) );
  NAND U8483 ( .A(n4897), .B(ereg[103]), .Z(n5309) );
  NAND U8484 ( .A(n4892), .B(ereg[104]), .Z(n5308) );
  NAND U8485 ( .A(n5310), .B(n5311), .Z(n3754) );
  NANDN U8486 ( .A(init), .B(e[105]), .Z(n5311) );
  AND U8487 ( .A(n5312), .B(n5313), .Z(n5310) );
  NAND U8488 ( .A(n4897), .B(ereg[104]), .Z(n5313) );
  NAND U8489 ( .A(n4892), .B(ereg[105]), .Z(n5312) );
  NAND U8490 ( .A(n5314), .B(n5315), .Z(n3753) );
  NANDN U8491 ( .A(init), .B(e[106]), .Z(n5315) );
  AND U8492 ( .A(n5316), .B(n5317), .Z(n5314) );
  NAND U8493 ( .A(n4897), .B(ereg[105]), .Z(n5317) );
  NAND U8494 ( .A(n4892), .B(ereg[106]), .Z(n5316) );
  NAND U8495 ( .A(n5318), .B(n5319), .Z(n3752) );
  NANDN U8496 ( .A(init), .B(e[107]), .Z(n5319) );
  AND U8497 ( .A(n5320), .B(n5321), .Z(n5318) );
  NAND U8498 ( .A(n4897), .B(ereg[106]), .Z(n5321) );
  NAND U8499 ( .A(n4892), .B(ereg[107]), .Z(n5320) );
  NAND U8500 ( .A(n5322), .B(n5323), .Z(n3751) );
  NANDN U8501 ( .A(init), .B(e[108]), .Z(n5323) );
  AND U8502 ( .A(n5324), .B(n5325), .Z(n5322) );
  NAND U8503 ( .A(n4897), .B(ereg[107]), .Z(n5325) );
  NAND U8504 ( .A(n4892), .B(ereg[108]), .Z(n5324) );
  NAND U8505 ( .A(n5326), .B(n5327), .Z(n3750) );
  NANDN U8506 ( .A(init), .B(e[109]), .Z(n5327) );
  AND U8507 ( .A(n5328), .B(n5329), .Z(n5326) );
  NAND U8508 ( .A(n4897), .B(ereg[108]), .Z(n5329) );
  NAND U8509 ( .A(n4892), .B(ereg[109]), .Z(n5328) );
  NAND U8510 ( .A(n5330), .B(n5331), .Z(n3749) );
  NANDN U8511 ( .A(init), .B(e[110]), .Z(n5331) );
  AND U8512 ( .A(n5332), .B(n5333), .Z(n5330) );
  NAND U8513 ( .A(n4897), .B(ereg[109]), .Z(n5333) );
  NAND U8514 ( .A(n4892), .B(ereg[110]), .Z(n5332) );
  NAND U8515 ( .A(n5334), .B(n5335), .Z(n3748) );
  NANDN U8516 ( .A(init), .B(e[111]), .Z(n5335) );
  AND U8517 ( .A(n5336), .B(n5337), .Z(n5334) );
  NAND U8518 ( .A(n4897), .B(ereg[110]), .Z(n5337) );
  NAND U8519 ( .A(n4892), .B(ereg[111]), .Z(n5336) );
  NAND U8520 ( .A(n5338), .B(n5339), .Z(n3747) );
  NANDN U8521 ( .A(init), .B(e[112]), .Z(n5339) );
  AND U8522 ( .A(n5340), .B(n5341), .Z(n5338) );
  NAND U8523 ( .A(n4897), .B(ereg[111]), .Z(n5341) );
  NAND U8524 ( .A(n4892), .B(ereg[112]), .Z(n5340) );
  NAND U8525 ( .A(n5342), .B(n5343), .Z(n3746) );
  NANDN U8526 ( .A(init), .B(e[113]), .Z(n5343) );
  AND U8527 ( .A(n5344), .B(n5345), .Z(n5342) );
  NAND U8528 ( .A(n4897), .B(ereg[112]), .Z(n5345) );
  NAND U8529 ( .A(n4892), .B(ereg[113]), .Z(n5344) );
  NAND U8530 ( .A(n5346), .B(n5347), .Z(n3745) );
  NANDN U8531 ( .A(init), .B(e[114]), .Z(n5347) );
  AND U8532 ( .A(n5348), .B(n5349), .Z(n5346) );
  NAND U8533 ( .A(n4897), .B(ereg[113]), .Z(n5349) );
  NAND U8534 ( .A(n4892), .B(ereg[114]), .Z(n5348) );
  NAND U8535 ( .A(n5350), .B(n5351), .Z(n3744) );
  NANDN U8536 ( .A(init), .B(e[115]), .Z(n5351) );
  AND U8537 ( .A(n5352), .B(n5353), .Z(n5350) );
  NAND U8538 ( .A(n4897), .B(ereg[114]), .Z(n5353) );
  NAND U8539 ( .A(n4892), .B(ereg[115]), .Z(n5352) );
  NAND U8540 ( .A(n5354), .B(n5355), .Z(n3743) );
  NANDN U8541 ( .A(init), .B(e[116]), .Z(n5355) );
  AND U8542 ( .A(n5356), .B(n5357), .Z(n5354) );
  NAND U8543 ( .A(n4897), .B(ereg[115]), .Z(n5357) );
  NAND U8544 ( .A(n4892), .B(ereg[116]), .Z(n5356) );
  NAND U8545 ( .A(n5358), .B(n5359), .Z(n3742) );
  NANDN U8546 ( .A(init), .B(e[117]), .Z(n5359) );
  AND U8547 ( .A(n5360), .B(n5361), .Z(n5358) );
  NAND U8548 ( .A(n4897), .B(ereg[116]), .Z(n5361) );
  NAND U8549 ( .A(n4892), .B(ereg[117]), .Z(n5360) );
  NAND U8550 ( .A(n5362), .B(n5363), .Z(n3741) );
  NANDN U8551 ( .A(init), .B(e[118]), .Z(n5363) );
  AND U8552 ( .A(n5364), .B(n5365), .Z(n5362) );
  NAND U8553 ( .A(n4897), .B(ereg[117]), .Z(n5365) );
  NAND U8554 ( .A(n4892), .B(ereg[118]), .Z(n5364) );
  NAND U8555 ( .A(n5366), .B(n5367), .Z(n3740) );
  NANDN U8556 ( .A(init), .B(e[119]), .Z(n5367) );
  AND U8557 ( .A(n5368), .B(n5369), .Z(n5366) );
  NAND U8558 ( .A(n4897), .B(ereg[118]), .Z(n5369) );
  NAND U8559 ( .A(n4892), .B(ereg[119]), .Z(n5368) );
  NAND U8560 ( .A(n5370), .B(n5371), .Z(n3739) );
  NANDN U8561 ( .A(init), .B(e[120]), .Z(n5371) );
  AND U8562 ( .A(n5372), .B(n5373), .Z(n5370) );
  NAND U8563 ( .A(n4897), .B(ereg[119]), .Z(n5373) );
  NAND U8564 ( .A(n4892), .B(ereg[120]), .Z(n5372) );
  NAND U8565 ( .A(n5374), .B(n5375), .Z(n3738) );
  NANDN U8566 ( .A(init), .B(e[121]), .Z(n5375) );
  AND U8567 ( .A(n5376), .B(n5377), .Z(n5374) );
  NAND U8568 ( .A(n4897), .B(ereg[120]), .Z(n5377) );
  NAND U8569 ( .A(n4892), .B(ereg[121]), .Z(n5376) );
  NAND U8570 ( .A(n5378), .B(n5379), .Z(n3737) );
  NANDN U8571 ( .A(init), .B(e[122]), .Z(n5379) );
  AND U8572 ( .A(n5380), .B(n5381), .Z(n5378) );
  NAND U8573 ( .A(n4897), .B(ereg[121]), .Z(n5381) );
  NAND U8574 ( .A(n4892), .B(ereg[122]), .Z(n5380) );
  NAND U8575 ( .A(n5382), .B(n5383), .Z(n3736) );
  NANDN U8576 ( .A(init), .B(e[123]), .Z(n5383) );
  AND U8577 ( .A(n5384), .B(n5385), .Z(n5382) );
  NAND U8578 ( .A(n4897), .B(ereg[122]), .Z(n5385) );
  NAND U8579 ( .A(n4892), .B(ereg[123]), .Z(n5384) );
  NAND U8580 ( .A(n5386), .B(n5387), .Z(n3735) );
  NANDN U8581 ( .A(init), .B(e[124]), .Z(n5387) );
  AND U8582 ( .A(n5388), .B(n5389), .Z(n5386) );
  NAND U8583 ( .A(n4897), .B(ereg[123]), .Z(n5389) );
  NAND U8584 ( .A(n4892), .B(ereg[124]), .Z(n5388) );
  NAND U8585 ( .A(n5390), .B(n5391), .Z(n3734) );
  NANDN U8586 ( .A(init), .B(e[125]), .Z(n5391) );
  AND U8587 ( .A(n5392), .B(n5393), .Z(n5390) );
  NAND U8588 ( .A(n4897), .B(ereg[124]), .Z(n5393) );
  NAND U8589 ( .A(n4892), .B(ereg[125]), .Z(n5392) );
  NAND U8590 ( .A(n5394), .B(n5395), .Z(n3733) );
  NANDN U8591 ( .A(init), .B(e[126]), .Z(n5395) );
  AND U8592 ( .A(n5396), .B(n5397), .Z(n5394) );
  NAND U8593 ( .A(n4897), .B(ereg[125]), .Z(n5397) );
  NAND U8594 ( .A(n4892), .B(ereg[126]), .Z(n5396) );
  NAND U8595 ( .A(n5398), .B(n5399), .Z(n3732) );
  NANDN U8596 ( .A(init), .B(e[127]), .Z(n5399) );
  AND U8597 ( .A(n5400), .B(n5401), .Z(n5398) );
  NAND U8598 ( .A(n4897), .B(ereg[126]), .Z(n5401) );
  NAND U8599 ( .A(n4892), .B(ereg[127]), .Z(n5400) );
  NAND U8600 ( .A(n5402), .B(n5403), .Z(n3731) );
  NANDN U8601 ( .A(init), .B(e[128]), .Z(n5403) );
  AND U8602 ( .A(n5404), .B(n5405), .Z(n5402) );
  NAND U8603 ( .A(n4897), .B(ereg[127]), .Z(n5405) );
  NAND U8604 ( .A(n4892), .B(ereg[128]), .Z(n5404) );
  NAND U8605 ( .A(n5406), .B(n5407), .Z(n3730) );
  NANDN U8606 ( .A(init), .B(e[129]), .Z(n5407) );
  AND U8607 ( .A(n5408), .B(n5409), .Z(n5406) );
  NAND U8608 ( .A(n4897), .B(ereg[128]), .Z(n5409) );
  NAND U8609 ( .A(n4892), .B(ereg[129]), .Z(n5408) );
  NAND U8610 ( .A(n5410), .B(n5411), .Z(n3729) );
  NANDN U8611 ( .A(init), .B(e[130]), .Z(n5411) );
  AND U8612 ( .A(n5412), .B(n5413), .Z(n5410) );
  NAND U8613 ( .A(n4897), .B(ereg[129]), .Z(n5413) );
  NAND U8614 ( .A(n4892), .B(ereg[130]), .Z(n5412) );
  NAND U8615 ( .A(n5414), .B(n5415), .Z(n3728) );
  NANDN U8616 ( .A(init), .B(e[131]), .Z(n5415) );
  AND U8617 ( .A(n5416), .B(n5417), .Z(n5414) );
  NAND U8618 ( .A(n4897), .B(ereg[130]), .Z(n5417) );
  NAND U8619 ( .A(n4892), .B(ereg[131]), .Z(n5416) );
  NAND U8620 ( .A(n5418), .B(n5419), .Z(n3727) );
  NANDN U8621 ( .A(init), .B(e[132]), .Z(n5419) );
  AND U8622 ( .A(n5420), .B(n5421), .Z(n5418) );
  NAND U8623 ( .A(n4897), .B(ereg[131]), .Z(n5421) );
  NAND U8624 ( .A(n4892), .B(ereg[132]), .Z(n5420) );
  NAND U8625 ( .A(n5422), .B(n5423), .Z(n3726) );
  NANDN U8626 ( .A(init), .B(e[133]), .Z(n5423) );
  AND U8627 ( .A(n5424), .B(n5425), .Z(n5422) );
  NAND U8628 ( .A(n4897), .B(ereg[132]), .Z(n5425) );
  NAND U8629 ( .A(n4892), .B(ereg[133]), .Z(n5424) );
  NAND U8630 ( .A(n5426), .B(n5427), .Z(n3725) );
  NANDN U8631 ( .A(init), .B(e[134]), .Z(n5427) );
  AND U8632 ( .A(n5428), .B(n5429), .Z(n5426) );
  NAND U8633 ( .A(n4897), .B(ereg[133]), .Z(n5429) );
  NAND U8634 ( .A(n4892), .B(ereg[134]), .Z(n5428) );
  NAND U8635 ( .A(n5430), .B(n5431), .Z(n3724) );
  NANDN U8636 ( .A(init), .B(e[135]), .Z(n5431) );
  AND U8637 ( .A(n5432), .B(n5433), .Z(n5430) );
  NAND U8638 ( .A(n4897), .B(ereg[134]), .Z(n5433) );
  NAND U8639 ( .A(n4892), .B(ereg[135]), .Z(n5432) );
  NAND U8640 ( .A(n5434), .B(n5435), .Z(n3723) );
  NANDN U8641 ( .A(init), .B(e[136]), .Z(n5435) );
  AND U8642 ( .A(n5436), .B(n5437), .Z(n5434) );
  NAND U8643 ( .A(n4897), .B(ereg[135]), .Z(n5437) );
  NAND U8644 ( .A(n4892), .B(ereg[136]), .Z(n5436) );
  NAND U8645 ( .A(n5438), .B(n5439), .Z(n3722) );
  NANDN U8646 ( .A(init), .B(e[137]), .Z(n5439) );
  AND U8647 ( .A(n5440), .B(n5441), .Z(n5438) );
  NAND U8648 ( .A(n4897), .B(ereg[136]), .Z(n5441) );
  NAND U8649 ( .A(n4892), .B(ereg[137]), .Z(n5440) );
  NAND U8650 ( .A(n5442), .B(n5443), .Z(n3721) );
  NANDN U8651 ( .A(init), .B(e[138]), .Z(n5443) );
  AND U8652 ( .A(n5444), .B(n5445), .Z(n5442) );
  NAND U8653 ( .A(n4897), .B(ereg[137]), .Z(n5445) );
  NAND U8654 ( .A(n4892), .B(ereg[138]), .Z(n5444) );
  NAND U8655 ( .A(n5446), .B(n5447), .Z(n3720) );
  NANDN U8656 ( .A(init), .B(e[139]), .Z(n5447) );
  AND U8657 ( .A(n5448), .B(n5449), .Z(n5446) );
  NAND U8658 ( .A(n4897), .B(ereg[138]), .Z(n5449) );
  NAND U8659 ( .A(n4892), .B(ereg[139]), .Z(n5448) );
  NAND U8660 ( .A(n5450), .B(n5451), .Z(n3719) );
  NANDN U8661 ( .A(init), .B(e[140]), .Z(n5451) );
  AND U8662 ( .A(n5452), .B(n5453), .Z(n5450) );
  NAND U8663 ( .A(n4897), .B(ereg[139]), .Z(n5453) );
  NAND U8664 ( .A(n4892), .B(ereg[140]), .Z(n5452) );
  NAND U8665 ( .A(n5454), .B(n5455), .Z(n3718) );
  NANDN U8666 ( .A(init), .B(e[141]), .Z(n5455) );
  AND U8667 ( .A(n5456), .B(n5457), .Z(n5454) );
  NAND U8668 ( .A(n4897), .B(ereg[140]), .Z(n5457) );
  NAND U8669 ( .A(n4892), .B(ereg[141]), .Z(n5456) );
  NAND U8670 ( .A(n5458), .B(n5459), .Z(n3717) );
  NANDN U8671 ( .A(init), .B(e[142]), .Z(n5459) );
  AND U8672 ( .A(n5460), .B(n5461), .Z(n5458) );
  NAND U8673 ( .A(n4897), .B(ereg[141]), .Z(n5461) );
  NAND U8674 ( .A(n4892), .B(ereg[142]), .Z(n5460) );
  NAND U8675 ( .A(n5462), .B(n5463), .Z(n3716) );
  NANDN U8676 ( .A(init), .B(e[143]), .Z(n5463) );
  AND U8677 ( .A(n5464), .B(n5465), .Z(n5462) );
  NAND U8678 ( .A(n4897), .B(ereg[142]), .Z(n5465) );
  NAND U8679 ( .A(n4892), .B(ereg[143]), .Z(n5464) );
  NAND U8680 ( .A(n5466), .B(n5467), .Z(n3715) );
  NANDN U8681 ( .A(init), .B(e[144]), .Z(n5467) );
  AND U8682 ( .A(n5468), .B(n5469), .Z(n5466) );
  NAND U8683 ( .A(n4897), .B(ereg[143]), .Z(n5469) );
  NAND U8684 ( .A(n4892), .B(ereg[144]), .Z(n5468) );
  NAND U8685 ( .A(n5470), .B(n5471), .Z(n3714) );
  NANDN U8686 ( .A(init), .B(e[145]), .Z(n5471) );
  AND U8687 ( .A(n5472), .B(n5473), .Z(n5470) );
  NAND U8688 ( .A(n4897), .B(ereg[144]), .Z(n5473) );
  NAND U8689 ( .A(n4892), .B(ereg[145]), .Z(n5472) );
  NAND U8690 ( .A(n5474), .B(n5475), .Z(n3713) );
  NANDN U8691 ( .A(init), .B(e[146]), .Z(n5475) );
  AND U8692 ( .A(n5476), .B(n5477), .Z(n5474) );
  NAND U8693 ( .A(n4897), .B(ereg[145]), .Z(n5477) );
  NAND U8694 ( .A(n4892), .B(ereg[146]), .Z(n5476) );
  NAND U8695 ( .A(n5478), .B(n5479), .Z(n3712) );
  NANDN U8696 ( .A(init), .B(e[147]), .Z(n5479) );
  AND U8697 ( .A(n5480), .B(n5481), .Z(n5478) );
  NAND U8698 ( .A(n4897), .B(ereg[146]), .Z(n5481) );
  NAND U8699 ( .A(n4892), .B(ereg[147]), .Z(n5480) );
  NAND U8700 ( .A(n5482), .B(n5483), .Z(n3711) );
  NANDN U8701 ( .A(init), .B(e[148]), .Z(n5483) );
  AND U8702 ( .A(n5484), .B(n5485), .Z(n5482) );
  NAND U8703 ( .A(n4897), .B(ereg[147]), .Z(n5485) );
  NAND U8704 ( .A(n4892), .B(ereg[148]), .Z(n5484) );
  NAND U8705 ( .A(n5486), .B(n5487), .Z(n3710) );
  NANDN U8706 ( .A(init), .B(e[149]), .Z(n5487) );
  AND U8707 ( .A(n5488), .B(n5489), .Z(n5486) );
  NAND U8708 ( .A(n4897), .B(ereg[148]), .Z(n5489) );
  NAND U8709 ( .A(n4892), .B(ereg[149]), .Z(n5488) );
  NAND U8710 ( .A(n5490), .B(n5491), .Z(n3709) );
  NANDN U8711 ( .A(init), .B(e[150]), .Z(n5491) );
  AND U8712 ( .A(n5492), .B(n5493), .Z(n5490) );
  NAND U8713 ( .A(n4897), .B(ereg[149]), .Z(n5493) );
  NAND U8714 ( .A(n4892), .B(ereg[150]), .Z(n5492) );
  NAND U8715 ( .A(n5494), .B(n5495), .Z(n3708) );
  NANDN U8716 ( .A(init), .B(e[151]), .Z(n5495) );
  AND U8717 ( .A(n5496), .B(n5497), .Z(n5494) );
  NAND U8718 ( .A(n4897), .B(ereg[150]), .Z(n5497) );
  NAND U8719 ( .A(n4892), .B(ereg[151]), .Z(n5496) );
  NAND U8720 ( .A(n5498), .B(n5499), .Z(n3707) );
  NANDN U8721 ( .A(init), .B(e[152]), .Z(n5499) );
  AND U8722 ( .A(n5500), .B(n5501), .Z(n5498) );
  NAND U8723 ( .A(n4897), .B(ereg[151]), .Z(n5501) );
  NAND U8724 ( .A(n4892), .B(ereg[152]), .Z(n5500) );
  NAND U8725 ( .A(n5502), .B(n5503), .Z(n3706) );
  NANDN U8726 ( .A(init), .B(e[153]), .Z(n5503) );
  AND U8727 ( .A(n5504), .B(n5505), .Z(n5502) );
  NAND U8728 ( .A(n4897), .B(ereg[152]), .Z(n5505) );
  NAND U8729 ( .A(n4892), .B(ereg[153]), .Z(n5504) );
  NAND U8730 ( .A(n5506), .B(n5507), .Z(n3705) );
  NANDN U8731 ( .A(init), .B(e[154]), .Z(n5507) );
  AND U8732 ( .A(n5508), .B(n5509), .Z(n5506) );
  NAND U8733 ( .A(n4897), .B(ereg[153]), .Z(n5509) );
  NAND U8734 ( .A(n4892), .B(ereg[154]), .Z(n5508) );
  NAND U8735 ( .A(n5510), .B(n5511), .Z(n3704) );
  NANDN U8736 ( .A(init), .B(e[155]), .Z(n5511) );
  AND U8737 ( .A(n5512), .B(n5513), .Z(n5510) );
  NAND U8738 ( .A(n4897), .B(ereg[154]), .Z(n5513) );
  NAND U8739 ( .A(n4892), .B(ereg[155]), .Z(n5512) );
  NAND U8740 ( .A(n5514), .B(n5515), .Z(n3703) );
  NANDN U8741 ( .A(init), .B(e[156]), .Z(n5515) );
  AND U8742 ( .A(n5516), .B(n5517), .Z(n5514) );
  NAND U8743 ( .A(n4897), .B(ereg[155]), .Z(n5517) );
  NAND U8744 ( .A(n4892), .B(ereg[156]), .Z(n5516) );
  NAND U8745 ( .A(n5518), .B(n5519), .Z(n3702) );
  NANDN U8746 ( .A(init), .B(e[157]), .Z(n5519) );
  AND U8747 ( .A(n5520), .B(n5521), .Z(n5518) );
  NAND U8748 ( .A(n4897), .B(ereg[156]), .Z(n5521) );
  NAND U8749 ( .A(n4892), .B(ereg[157]), .Z(n5520) );
  NAND U8750 ( .A(n5522), .B(n5523), .Z(n3701) );
  NANDN U8751 ( .A(init), .B(e[158]), .Z(n5523) );
  AND U8752 ( .A(n5524), .B(n5525), .Z(n5522) );
  NAND U8753 ( .A(n4897), .B(ereg[157]), .Z(n5525) );
  NAND U8754 ( .A(n4892), .B(ereg[158]), .Z(n5524) );
  NAND U8755 ( .A(n5526), .B(n5527), .Z(n3700) );
  NANDN U8756 ( .A(init), .B(e[159]), .Z(n5527) );
  AND U8757 ( .A(n5528), .B(n5529), .Z(n5526) );
  NAND U8758 ( .A(n4897), .B(ereg[158]), .Z(n5529) );
  NAND U8759 ( .A(n4892), .B(ereg[159]), .Z(n5528) );
  NAND U8760 ( .A(n5530), .B(n5531), .Z(n3699) );
  NANDN U8761 ( .A(init), .B(e[160]), .Z(n5531) );
  AND U8762 ( .A(n5532), .B(n5533), .Z(n5530) );
  NAND U8763 ( .A(n4897), .B(ereg[159]), .Z(n5533) );
  NAND U8764 ( .A(n4892), .B(ereg[160]), .Z(n5532) );
  NAND U8765 ( .A(n5534), .B(n5535), .Z(n3698) );
  NANDN U8766 ( .A(init), .B(e[161]), .Z(n5535) );
  AND U8767 ( .A(n5536), .B(n5537), .Z(n5534) );
  NAND U8768 ( .A(n4897), .B(ereg[160]), .Z(n5537) );
  NAND U8769 ( .A(n4892), .B(ereg[161]), .Z(n5536) );
  NAND U8770 ( .A(n5538), .B(n5539), .Z(n3697) );
  NANDN U8771 ( .A(init), .B(e[162]), .Z(n5539) );
  AND U8772 ( .A(n5540), .B(n5541), .Z(n5538) );
  NAND U8773 ( .A(n4897), .B(ereg[161]), .Z(n5541) );
  NAND U8774 ( .A(n4892), .B(ereg[162]), .Z(n5540) );
  NAND U8775 ( .A(n5542), .B(n5543), .Z(n3696) );
  NANDN U8776 ( .A(init), .B(e[163]), .Z(n5543) );
  AND U8777 ( .A(n5544), .B(n5545), .Z(n5542) );
  NAND U8778 ( .A(n4897), .B(ereg[162]), .Z(n5545) );
  NAND U8779 ( .A(n4892), .B(ereg[163]), .Z(n5544) );
  NAND U8780 ( .A(n5546), .B(n5547), .Z(n3695) );
  NANDN U8781 ( .A(init), .B(e[164]), .Z(n5547) );
  AND U8782 ( .A(n5548), .B(n5549), .Z(n5546) );
  NAND U8783 ( .A(n4897), .B(ereg[163]), .Z(n5549) );
  NAND U8784 ( .A(n4892), .B(ereg[164]), .Z(n5548) );
  NAND U8785 ( .A(n5550), .B(n5551), .Z(n3694) );
  NANDN U8786 ( .A(init), .B(e[165]), .Z(n5551) );
  AND U8787 ( .A(n5552), .B(n5553), .Z(n5550) );
  NAND U8788 ( .A(n4897), .B(ereg[164]), .Z(n5553) );
  NAND U8789 ( .A(n4892), .B(ereg[165]), .Z(n5552) );
  NAND U8790 ( .A(n5554), .B(n5555), .Z(n3693) );
  NANDN U8791 ( .A(init), .B(e[166]), .Z(n5555) );
  AND U8792 ( .A(n5556), .B(n5557), .Z(n5554) );
  NAND U8793 ( .A(n4897), .B(ereg[165]), .Z(n5557) );
  NAND U8794 ( .A(n4892), .B(ereg[166]), .Z(n5556) );
  NAND U8795 ( .A(n5558), .B(n5559), .Z(n3692) );
  NANDN U8796 ( .A(init), .B(e[167]), .Z(n5559) );
  AND U8797 ( .A(n5560), .B(n5561), .Z(n5558) );
  NAND U8798 ( .A(n4897), .B(ereg[166]), .Z(n5561) );
  NAND U8799 ( .A(n4892), .B(ereg[167]), .Z(n5560) );
  NAND U8800 ( .A(n5562), .B(n5563), .Z(n3691) );
  NANDN U8801 ( .A(init), .B(e[168]), .Z(n5563) );
  AND U8802 ( .A(n5564), .B(n5565), .Z(n5562) );
  NAND U8803 ( .A(n4897), .B(ereg[167]), .Z(n5565) );
  NAND U8804 ( .A(n4892), .B(ereg[168]), .Z(n5564) );
  NAND U8805 ( .A(n5566), .B(n5567), .Z(n3690) );
  NANDN U8806 ( .A(init), .B(e[169]), .Z(n5567) );
  AND U8807 ( .A(n5568), .B(n5569), .Z(n5566) );
  NAND U8808 ( .A(n4897), .B(ereg[168]), .Z(n5569) );
  NAND U8809 ( .A(n4892), .B(ereg[169]), .Z(n5568) );
  NAND U8810 ( .A(n5570), .B(n5571), .Z(n3689) );
  NANDN U8811 ( .A(init), .B(e[170]), .Z(n5571) );
  AND U8812 ( .A(n5572), .B(n5573), .Z(n5570) );
  NAND U8813 ( .A(n4897), .B(ereg[169]), .Z(n5573) );
  NAND U8814 ( .A(n4892), .B(ereg[170]), .Z(n5572) );
  NAND U8815 ( .A(n5574), .B(n5575), .Z(n3688) );
  NANDN U8816 ( .A(init), .B(e[171]), .Z(n5575) );
  AND U8817 ( .A(n5576), .B(n5577), .Z(n5574) );
  NAND U8818 ( .A(n4897), .B(ereg[170]), .Z(n5577) );
  NAND U8819 ( .A(n4892), .B(ereg[171]), .Z(n5576) );
  NAND U8820 ( .A(n5578), .B(n5579), .Z(n3687) );
  NANDN U8821 ( .A(init), .B(e[172]), .Z(n5579) );
  AND U8822 ( .A(n5580), .B(n5581), .Z(n5578) );
  NAND U8823 ( .A(n4897), .B(ereg[171]), .Z(n5581) );
  NAND U8824 ( .A(n4892), .B(ereg[172]), .Z(n5580) );
  NAND U8825 ( .A(n5582), .B(n5583), .Z(n3686) );
  NANDN U8826 ( .A(init), .B(e[173]), .Z(n5583) );
  AND U8827 ( .A(n5584), .B(n5585), .Z(n5582) );
  NAND U8828 ( .A(n4897), .B(ereg[172]), .Z(n5585) );
  NAND U8829 ( .A(n4892), .B(ereg[173]), .Z(n5584) );
  NAND U8830 ( .A(n5586), .B(n5587), .Z(n3685) );
  NANDN U8831 ( .A(init), .B(e[174]), .Z(n5587) );
  AND U8832 ( .A(n5588), .B(n5589), .Z(n5586) );
  NAND U8833 ( .A(n4897), .B(ereg[173]), .Z(n5589) );
  NAND U8834 ( .A(n4892), .B(ereg[174]), .Z(n5588) );
  NAND U8835 ( .A(n5590), .B(n5591), .Z(n3684) );
  NANDN U8836 ( .A(init), .B(e[175]), .Z(n5591) );
  AND U8837 ( .A(n5592), .B(n5593), .Z(n5590) );
  NAND U8838 ( .A(n4897), .B(ereg[174]), .Z(n5593) );
  NAND U8839 ( .A(n4892), .B(ereg[175]), .Z(n5592) );
  NAND U8840 ( .A(n5594), .B(n5595), .Z(n3683) );
  NANDN U8841 ( .A(init), .B(e[176]), .Z(n5595) );
  AND U8842 ( .A(n5596), .B(n5597), .Z(n5594) );
  NAND U8843 ( .A(n4897), .B(ereg[175]), .Z(n5597) );
  NAND U8844 ( .A(n4892), .B(ereg[176]), .Z(n5596) );
  NAND U8845 ( .A(n5598), .B(n5599), .Z(n3682) );
  NANDN U8846 ( .A(init), .B(e[177]), .Z(n5599) );
  AND U8847 ( .A(n5600), .B(n5601), .Z(n5598) );
  NAND U8848 ( .A(n4897), .B(ereg[176]), .Z(n5601) );
  NAND U8849 ( .A(n4892), .B(ereg[177]), .Z(n5600) );
  NAND U8850 ( .A(n5602), .B(n5603), .Z(n3681) );
  NANDN U8851 ( .A(init), .B(e[178]), .Z(n5603) );
  AND U8852 ( .A(n5604), .B(n5605), .Z(n5602) );
  NAND U8853 ( .A(n4897), .B(ereg[177]), .Z(n5605) );
  NAND U8854 ( .A(n4892), .B(ereg[178]), .Z(n5604) );
  NAND U8855 ( .A(n5606), .B(n5607), .Z(n3680) );
  NANDN U8856 ( .A(init), .B(e[179]), .Z(n5607) );
  AND U8857 ( .A(n5608), .B(n5609), .Z(n5606) );
  NAND U8858 ( .A(n4897), .B(ereg[178]), .Z(n5609) );
  NAND U8859 ( .A(n4892), .B(ereg[179]), .Z(n5608) );
  NAND U8860 ( .A(n5610), .B(n5611), .Z(n3679) );
  NANDN U8861 ( .A(init), .B(e[180]), .Z(n5611) );
  AND U8862 ( .A(n5612), .B(n5613), .Z(n5610) );
  NAND U8863 ( .A(n4897), .B(ereg[179]), .Z(n5613) );
  NAND U8864 ( .A(n4892), .B(ereg[180]), .Z(n5612) );
  NAND U8865 ( .A(n5614), .B(n5615), .Z(n3678) );
  NANDN U8866 ( .A(init), .B(e[181]), .Z(n5615) );
  AND U8867 ( .A(n5616), .B(n5617), .Z(n5614) );
  NAND U8868 ( .A(n4897), .B(ereg[180]), .Z(n5617) );
  NAND U8869 ( .A(n4892), .B(ereg[181]), .Z(n5616) );
  NAND U8870 ( .A(n5618), .B(n5619), .Z(n3677) );
  NANDN U8871 ( .A(init), .B(e[182]), .Z(n5619) );
  AND U8872 ( .A(n5620), .B(n5621), .Z(n5618) );
  NAND U8873 ( .A(n4897), .B(ereg[181]), .Z(n5621) );
  NAND U8874 ( .A(n4892), .B(ereg[182]), .Z(n5620) );
  NAND U8875 ( .A(n5622), .B(n5623), .Z(n3676) );
  NANDN U8876 ( .A(init), .B(e[183]), .Z(n5623) );
  AND U8877 ( .A(n5624), .B(n5625), .Z(n5622) );
  NAND U8878 ( .A(n4897), .B(ereg[182]), .Z(n5625) );
  NAND U8879 ( .A(n4892), .B(ereg[183]), .Z(n5624) );
  NAND U8880 ( .A(n5626), .B(n5627), .Z(n3675) );
  NANDN U8881 ( .A(init), .B(e[184]), .Z(n5627) );
  AND U8882 ( .A(n5628), .B(n5629), .Z(n5626) );
  NAND U8883 ( .A(n4897), .B(ereg[183]), .Z(n5629) );
  NAND U8884 ( .A(n4892), .B(ereg[184]), .Z(n5628) );
  NAND U8885 ( .A(n5630), .B(n5631), .Z(n3674) );
  NANDN U8886 ( .A(init), .B(e[185]), .Z(n5631) );
  AND U8887 ( .A(n5632), .B(n5633), .Z(n5630) );
  NAND U8888 ( .A(n4897), .B(ereg[184]), .Z(n5633) );
  NAND U8889 ( .A(n4892), .B(ereg[185]), .Z(n5632) );
  NAND U8890 ( .A(n5634), .B(n5635), .Z(n3673) );
  NANDN U8891 ( .A(init), .B(e[186]), .Z(n5635) );
  AND U8892 ( .A(n5636), .B(n5637), .Z(n5634) );
  NAND U8893 ( .A(n4897), .B(ereg[185]), .Z(n5637) );
  NAND U8894 ( .A(n4892), .B(ereg[186]), .Z(n5636) );
  NAND U8895 ( .A(n5638), .B(n5639), .Z(n3672) );
  NANDN U8896 ( .A(init), .B(e[187]), .Z(n5639) );
  AND U8897 ( .A(n5640), .B(n5641), .Z(n5638) );
  NAND U8898 ( .A(n4897), .B(ereg[186]), .Z(n5641) );
  NAND U8899 ( .A(n4892), .B(ereg[187]), .Z(n5640) );
  NAND U8900 ( .A(n5642), .B(n5643), .Z(n3671) );
  NANDN U8901 ( .A(init), .B(e[188]), .Z(n5643) );
  AND U8902 ( .A(n5644), .B(n5645), .Z(n5642) );
  NAND U8903 ( .A(n4897), .B(ereg[187]), .Z(n5645) );
  NAND U8904 ( .A(n4892), .B(ereg[188]), .Z(n5644) );
  NAND U8905 ( .A(n5646), .B(n5647), .Z(n3670) );
  NANDN U8906 ( .A(init), .B(e[189]), .Z(n5647) );
  AND U8907 ( .A(n5648), .B(n5649), .Z(n5646) );
  NAND U8908 ( .A(n4897), .B(ereg[188]), .Z(n5649) );
  NAND U8909 ( .A(n4892), .B(ereg[189]), .Z(n5648) );
  NAND U8910 ( .A(n5650), .B(n5651), .Z(n3669) );
  NANDN U8911 ( .A(init), .B(e[190]), .Z(n5651) );
  AND U8912 ( .A(n5652), .B(n5653), .Z(n5650) );
  NAND U8913 ( .A(n4897), .B(ereg[189]), .Z(n5653) );
  NAND U8914 ( .A(n4892), .B(ereg[190]), .Z(n5652) );
  NAND U8915 ( .A(n5654), .B(n5655), .Z(n3668) );
  NANDN U8916 ( .A(init), .B(e[191]), .Z(n5655) );
  AND U8917 ( .A(n5656), .B(n5657), .Z(n5654) );
  NAND U8918 ( .A(n4897), .B(ereg[190]), .Z(n5657) );
  NAND U8919 ( .A(n4892), .B(ereg[191]), .Z(n5656) );
  NAND U8920 ( .A(n5658), .B(n5659), .Z(n3667) );
  NANDN U8921 ( .A(init), .B(e[192]), .Z(n5659) );
  AND U8922 ( .A(n5660), .B(n5661), .Z(n5658) );
  NAND U8923 ( .A(n4897), .B(ereg[191]), .Z(n5661) );
  NAND U8924 ( .A(n4892), .B(ereg[192]), .Z(n5660) );
  NAND U8925 ( .A(n5662), .B(n5663), .Z(n3666) );
  NANDN U8926 ( .A(init), .B(e[193]), .Z(n5663) );
  AND U8927 ( .A(n5664), .B(n5665), .Z(n5662) );
  NAND U8928 ( .A(n4897), .B(ereg[192]), .Z(n5665) );
  NAND U8929 ( .A(n4892), .B(ereg[193]), .Z(n5664) );
  NAND U8930 ( .A(n5666), .B(n5667), .Z(n3665) );
  NANDN U8931 ( .A(init), .B(e[194]), .Z(n5667) );
  AND U8932 ( .A(n5668), .B(n5669), .Z(n5666) );
  NAND U8933 ( .A(n4897), .B(ereg[193]), .Z(n5669) );
  NAND U8934 ( .A(n4892), .B(ereg[194]), .Z(n5668) );
  NAND U8935 ( .A(n5670), .B(n5671), .Z(n3664) );
  NANDN U8936 ( .A(init), .B(e[195]), .Z(n5671) );
  AND U8937 ( .A(n5672), .B(n5673), .Z(n5670) );
  NAND U8938 ( .A(n4897), .B(ereg[194]), .Z(n5673) );
  NAND U8939 ( .A(n4892), .B(ereg[195]), .Z(n5672) );
  NAND U8940 ( .A(n5674), .B(n5675), .Z(n3663) );
  NANDN U8941 ( .A(init), .B(e[196]), .Z(n5675) );
  AND U8942 ( .A(n5676), .B(n5677), .Z(n5674) );
  NAND U8943 ( .A(n4897), .B(ereg[195]), .Z(n5677) );
  NAND U8944 ( .A(n4892), .B(ereg[196]), .Z(n5676) );
  NAND U8945 ( .A(n5678), .B(n5679), .Z(n3662) );
  NANDN U8946 ( .A(init), .B(e[197]), .Z(n5679) );
  AND U8947 ( .A(n5680), .B(n5681), .Z(n5678) );
  NAND U8948 ( .A(n4897), .B(ereg[196]), .Z(n5681) );
  NAND U8949 ( .A(n4892), .B(ereg[197]), .Z(n5680) );
  NAND U8950 ( .A(n5682), .B(n5683), .Z(n3661) );
  NANDN U8951 ( .A(init), .B(e[198]), .Z(n5683) );
  AND U8952 ( .A(n5684), .B(n5685), .Z(n5682) );
  NAND U8953 ( .A(n4897), .B(ereg[197]), .Z(n5685) );
  NAND U8954 ( .A(n4892), .B(ereg[198]), .Z(n5684) );
  NAND U8955 ( .A(n5686), .B(n5687), .Z(n3660) );
  NANDN U8956 ( .A(init), .B(e[199]), .Z(n5687) );
  AND U8957 ( .A(n5688), .B(n5689), .Z(n5686) );
  NAND U8958 ( .A(n4897), .B(ereg[198]), .Z(n5689) );
  NAND U8959 ( .A(n4892), .B(ereg[199]), .Z(n5688) );
  NAND U8960 ( .A(n5690), .B(n5691), .Z(n3659) );
  NANDN U8961 ( .A(init), .B(e[200]), .Z(n5691) );
  AND U8962 ( .A(n5692), .B(n5693), .Z(n5690) );
  NAND U8963 ( .A(n4897), .B(ereg[199]), .Z(n5693) );
  NAND U8964 ( .A(n4892), .B(ereg[200]), .Z(n5692) );
  NAND U8965 ( .A(n5694), .B(n5695), .Z(n3658) );
  NANDN U8966 ( .A(init), .B(e[201]), .Z(n5695) );
  AND U8967 ( .A(n5696), .B(n5697), .Z(n5694) );
  NAND U8968 ( .A(n4897), .B(ereg[200]), .Z(n5697) );
  NAND U8969 ( .A(n4892), .B(ereg[201]), .Z(n5696) );
  NAND U8970 ( .A(n5698), .B(n5699), .Z(n3657) );
  NANDN U8971 ( .A(init), .B(e[202]), .Z(n5699) );
  AND U8972 ( .A(n5700), .B(n5701), .Z(n5698) );
  NAND U8973 ( .A(n4897), .B(ereg[201]), .Z(n5701) );
  NAND U8974 ( .A(n4892), .B(ereg[202]), .Z(n5700) );
  NAND U8975 ( .A(n5702), .B(n5703), .Z(n3656) );
  NANDN U8976 ( .A(init), .B(e[203]), .Z(n5703) );
  AND U8977 ( .A(n5704), .B(n5705), .Z(n5702) );
  NAND U8978 ( .A(n4897), .B(ereg[202]), .Z(n5705) );
  NAND U8979 ( .A(n4892), .B(ereg[203]), .Z(n5704) );
  NAND U8980 ( .A(n5706), .B(n5707), .Z(n3655) );
  NANDN U8981 ( .A(init), .B(e[204]), .Z(n5707) );
  AND U8982 ( .A(n5708), .B(n5709), .Z(n5706) );
  NAND U8983 ( .A(n4897), .B(ereg[203]), .Z(n5709) );
  NAND U8984 ( .A(n4892), .B(ereg[204]), .Z(n5708) );
  NAND U8985 ( .A(n5710), .B(n5711), .Z(n3654) );
  NANDN U8986 ( .A(init), .B(e[205]), .Z(n5711) );
  AND U8987 ( .A(n5712), .B(n5713), .Z(n5710) );
  NAND U8988 ( .A(n4897), .B(ereg[204]), .Z(n5713) );
  NAND U8989 ( .A(n4892), .B(ereg[205]), .Z(n5712) );
  NAND U8990 ( .A(n5714), .B(n5715), .Z(n3653) );
  NANDN U8991 ( .A(init), .B(e[206]), .Z(n5715) );
  AND U8992 ( .A(n5716), .B(n5717), .Z(n5714) );
  NAND U8993 ( .A(n4897), .B(ereg[205]), .Z(n5717) );
  NAND U8994 ( .A(n4892), .B(ereg[206]), .Z(n5716) );
  NAND U8995 ( .A(n5718), .B(n5719), .Z(n3652) );
  NANDN U8996 ( .A(init), .B(e[207]), .Z(n5719) );
  AND U8997 ( .A(n5720), .B(n5721), .Z(n5718) );
  NAND U8998 ( .A(n4897), .B(ereg[206]), .Z(n5721) );
  NAND U8999 ( .A(n4892), .B(ereg[207]), .Z(n5720) );
  NAND U9000 ( .A(n5722), .B(n5723), .Z(n3651) );
  NANDN U9001 ( .A(init), .B(e[208]), .Z(n5723) );
  AND U9002 ( .A(n5724), .B(n5725), .Z(n5722) );
  NAND U9003 ( .A(n4897), .B(ereg[207]), .Z(n5725) );
  NAND U9004 ( .A(n4892), .B(ereg[208]), .Z(n5724) );
  NAND U9005 ( .A(n5726), .B(n5727), .Z(n3650) );
  NANDN U9006 ( .A(init), .B(e[209]), .Z(n5727) );
  AND U9007 ( .A(n5728), .B(n5729), .Z(n5726) );
  NAND U9008 ( .A(n4897), .B(ereg[208]), .Z(n5729) );
  NAND U9009 ( .A(n4892), .B(ereg[209]), .Z(n5728) );
  NAND U9010 ( .A(n5730), .B(n5731), .Z(n3649) );
  NANDN U9011 ( .A(init), .B(e[210]), .Z(n5731) );
  AND U9012 ( .A(n5732), .B(n5733), .Z(n5730) );
  NAND U9013 ( .A(n4897), .B(ereg[209]), .Z(n5733) );
  NAND U9014 ( .A(n4892), .B(ereg[210]), .Z(n5732) );
  NAND U9015 ( .A(n5734), .B(n5735), .Z(n3648) );
  NANDN U9016 ( .A(init), .B(e[211]), .Z(n5735) );
  AND U9017 ( .A(n5736), .B(n5737), .Z(n5734) );
  NAND U9018 ( .A(n4897), .B(ereg[210]), .Z(n5737) );
  NAND U9019 ( .A(n4892), .B(ereg[211]), .Z(n5736) );
  NAND U9020 ( .A(n5738), .B(n5739), .Z(n3647) );
  NANDN U9021 ( .A(init), .B(e[212]), .Z(n5739) );
  AND U9022 ( .A(n5740), .B(n5741), .Z(n5738) );
  NAND U9023 ( .A(n4897), .B(ereg[211]), .Z(n5741) );
  NAND U9024 ( .A(n4892), .B(ereg[212]), .Z(n5740) );
  NAND U9025 ( .A(n5742), .B(n5743), .Z(n3646) );
  NANDN U9026 ( .A(init), .B(e[213]), .Z(n5743) );
  AND U9027 ( .A(n5744), .B(n5745), .Z(n5742) );
  NAND U9028 ( .A(n4897), .B(ereg[212]), .Z(n5745) );
  NAND U9029 ( .A(n4892), .B(ereg[213]), .Z(n5744) );
  NAND U9030 ( .A(n5746), .B(n5747), .Z(n3645) );
  NANDN U9031 ( .A(init), .B(e[214]), .Z(n5747) );
  AND U9032 ( .A(n5748), .B(n5749), .Z(n5746) );
  NAND U9033 ( .A(n4897), .B(ereg[213]), .Z(n5749) );
  NAND U9034 ( .A(n4892), .B(ereg[214]), .Z(n5748) );
  NAND U9035 ( .A(n5750), .B(n5751), .Z(n3644) );
  NANDN U9036 ( .A(init), .B(e[215]), .Z(n5751) );
  AND U9037 ( .A(n5752), .B(n5753), .Z(n5750) );
  NAND U9038 ( .A(n4897), .B(ereg[214]), .Z(n5753) );
  NAND U9039 ( .A(n4892), .B(ereg[215]), .Z(n5752) );
  NAND U9040 ( .A(n5754), .B(n5755), .Z(n3643) );
  NANDN U9041 ( .A(init), .B(e[216]), .Z(n5755) );
  AND U9042 ( .A(n5756), .B(n5757), .Z(n5754) );
  NAND U9043 ( .A(n4897), .B(ereg[215]), .Z(n5757) );
  NAND U9044 ( .A(n4892), .B(ereg[216]), .Z(n5756) );
  NAND U9045 ( .A(n5758), .B(n5759), .Z(n3642) );
  NANDN U9046 ( .A(init), .B(e[217]), .Z(n5759) );
  AND U9047 ( .A(n5760), .B(n5761), .Z(n5758) );
  NAND U9048 ( .A(n4897), .B(ereg[216]), .Z(n5761) );
  NAND U9049 ( .A(n4892), .B(ereg[217]), .Z(n5760) );
  NAND U9050 ( .A(n5762), .B(n5763), .Z(n3641) );
  NANDN U9051 ( .A(init), .B(e[218]), .Z(n5763) );
  AND U9052 ( .A(n5764), .B(n5765), .Z(n5762) );
  NAND U9053 ( .A(n4897), .B(ereg[217]), .Z(n5765) );
  NAND U9054 ( .A(n4892), .B(ereg[218]), .Z(n5764) );
  NAND U9055 ( .A(n5766), .B(n5767), .Z(n3640) );
  NANDN U9056 ( .A(init), .B(e[219]), .Z(n5767) );
  AND U9057 ( .A(n5768), .B(n5769), .Z(n5766) );
  NAND U9058 ( .A(n4897), .B(ereg[218]), .Z(n5769) );
  NAND U9059 ( .A(n4892), .B(ereg[219]), .Z(n5768) );
  NAND U9060 ( .A(n5770), .B(n5771), .Z(n3639) );
  NANDN U9061 ( .A(init), .B(e[220]), .Z(n5771) );
  AND U9062 ( .A(n5772), .B(n5773), .Z(n5770) );
  NAND U9063 ( .A(n4897), .B(ereg[219]), .Z(n5773) );
  NAND U9064 ( .A(n4892), .B(ereg[220]), .Z(n5772) );
  NAND U9065 ( .A(n5774), .B(n5775), .Z(n3638) );
  NANDN U9066 ( .A(init), .B(e[221]), .Z(n5775) );
  AND U9067 ( .A(n5776), .B(n5777), .Z(n5774) );
  NAND U9068 ( .A(n4897), .B(ereg[220]), .Z(n5777) );
  NAND U9069 ( .A(n4892), .B(ereg[221]), .Z(n5776) );
  NAND U9070 ( .A(n5778), .B(n5779), .Z(n3637) );
  NANDN U9071 ( .A(init), .B(e[222]), .Z(n5779) );
  AND U9072 ( .A(n5780), .B(n5781), .Z(n5778) );
  NAND U9073 ( .A(n4897), .B(ereg[221]), .Z(n5781) );
  NAND U9074 ( .A(n4892), .B(ereg[222]), .Z(n5780) );
  NAND U9075 ( .A(n5782), .B(n5783), .Z(n3636) );
  NANDN U9076 ( .A(init), .B(e[223]), .Z(n5783) );
  AND U9077 ( .A(n5784), .B(n5785), .Z(n5782) );
  NAND U9078 ( .A(n4897), .B(ereg[222]), .Z(n5785) );
  NAND U9079 ( .A(n4892), .B(ereg[223]), .Z(n5784) );
  NAND U9080 ( .A(n5786), .B(n5787), .Z(n3635) );
  NANDN U9081 ( .A(init), .B(e[224]), .Z(n5787) );
  AND U9082 ( .A(n5788), .B(n5789), .Z(n5786) );
  NAND U9083 ( .A(n4897), .B(ereg[223]), .Z(n5789) );
  NAND U9084 ( .A(n4892), .B(ereg[224]), .Z(n5788) );
  NAND U9085 ( .A(n5790), .B(n5791), .Z(n3634) );
  NANDN U9086 ( .A(init), .B(e[225]), .Z(n5791) );
  AND U9087 ( .A(n5792), .B(n5793), .Z(n5790) );
  NAND U9088 ( .A(n4897), .B(ereg[224]), .Z(n5793) );
  NAND U9089 ( .A(n4892), .B(ereg[225]), .Z(n5792) );
  NAND U9090 ( .A(n5794), .B(n5795), .Z(n3633) );
  NANDN U9091 ( .A(init), .B(e[226]), .Z(n5795) );
  AND U9092 ( .A(n5796), .B(n5797), .Z(n5794) );
  NAND U9093 ( .A(n4897), .B(ereg[225]), .Z(n5797) );
  NAND U9094 ( .A(n4892), .B(ereg[226]), .Z(n5796) );
  NAND U9095 ( .A(n5798), .B(n5799), .Z(n3632) );
  NANDN U9096 ( .A(init), .B(e[227]), .Z(n5799) );
  AND U9097 ( .A(n5800), .B(n5801), .Z(n5798) );
  NAND U9098 ( .A(n4897), .B(ereg[226]), .Z(n5801) );
  NAND U9099 ( .A(n4892), .B(ereg[227]), .Z(n5800) );
  NAND U9100 ( .A(n5802), .B(n5803), .Z(n3631) );
  NANDN U9101 ( .A(init), .B(e[228]), .Z(n5803) );
  AND U9102 ( .A(n5804), .B(n5805), .Z(n5802) );
  NAND U9103 ( .A(n4897), .B(ereg[227]), .Z(n5805) );
  NAND U9104 ( .A(n4892), .B(ereg[228]), .Z(n5804) );
  NAND U9105 ( .A(n5806), .B(n5807), .Z(n3630) );
  NANDN U9106 ( .A(init), .B(e[229]), .Z(n5807) );
  AND U9107 ( .A(n5808), .B(n5809), .Z(n5806) );
  NAND U9108 ( .A(n4897), .B(ereg[228]), .Z(n5809) );
  NAND U9109 ( .A(n4892), .B(ereg[229]), .Z(n5808) );
  NAND U9110 ( .A(n5810), .B(n5811), .Z(n3629) );
  NANDN U9111 ( .A(init), .B(e[230]), .Z(n5811) );
  AND U9112 ( .A(n5812), .B(n5813), .Z(n5810) );
  NAND U9113 ( .A(n4897), .B(ereg[229]), .Z(n5813) );
  NAND U9114 ( .A(n4892), .B(ereg[230]), .Z(n5812) );
  NAND U9115 ( .A(n5814), .B(n5815), .Z(n3628) );
  NANDN U9116 ( .A(init), .B(e[231]), .Z(n5815) );
  AND U9117 ( .A(n5816), .B(n5817), .Z(n5814) );
  NAND U9118 ( .A(n4897), .B(ereg[230]), .Z(n5817) );
  NAND U9119 ( .A(n4892), .B(ereg[231]), .Z(n5816) );
  NAND U9120 ( .A(n5818), .B(n5819), .Z(n3627) );
  NANDN U9121 ( .A(init), .B(e[232]), .Z(n5819) );
  AND U9122 ( .A(n5820), .B(n5821), .Z(n5818) );
  NAND U9123 ( .A(n4897), .B(ereg[231]), .Z(n5821) );
  NAND U9124 ( .A(n4892), .B(ereg[232]), .Z(n5820) );
  NAND U9125 ( .A(n5822), .B(n5823), .Z(n3626) );
  NANDN U9126 ( .A(init), .B(e[233]), .Z(n5823) );
  AND U9127 ( .A(n5824), .B(n5825), .Z(n5822) );
  NAND U9128 ( .A(n4897), .B(ereg[232]), .Z(n5825) );
  NAND U9129 ( .A(n4892), .B(ereg[233]), .Z(n5824) );
  NAND U9130 ( .A(n5826), .B(n5827), .Z(n3625) );
  NANDN U9131 ( .A(init), .B(e[234]), .Z(n5827) );
  AND U9132 ( .A(n5828), .B(n5829), .Z(n5826) );
  NAND U9133 ( .A(n4897), .B(ereg[233]), .Z(n5829) );
  NAND U9134 ( .A(n4892), .B(ereg[234]), .Z(n5828) );
  NAND U9135 ( .A(n5830), .B(n5831), .Z(n3624) );
  NANDN U9136 ( .A(init), .B(e[235]), .Z(n5831) );
  AND U9137 ( .A(n5832), .B(n5833), .Z(n5830) );
  NAND U9138 ( .A(n4897), .B(ereg[234]), .Z(n5833) );
  NAND U9139 ( .A(n4892), .B(ereg[235]), .Z(n5832) );
  NAND U9140 ( .A(n5834), .B(n5835), .Z(n3623) );
  NANDN U9141 ( .A(init), .B(e[236]), .Z(n5835) );
  AND U9142 ( .A(n5836), .B(n5837), .Z(n5834) );
  NAND U9143 ( .A(n4897), .B(ereg[235]), .Z(n5837) );
  NAND U9144 ( .A(n4892), .B(ereg[236]), .Z(n5836) );
  NAND U9145 ( .A(n5838), .B(n5839), .Z(n3622) );
  NANDN U9146 ( .A(init), .B(e[237]), .Z(n5839) );
  AND U9147 ( .A(n5840), .B(n5841), .Z(n5838) );
  NAND U9148 ( .A(n4897), .B(ereg[236]), .Z(n5841) );
  NAND U9149 ( .A(n4892), .B(ereg[237]), .Z(n5840) );
  NAND U9150 ( .A(n5842), .B(n5843), .Z(n3621) );
  NANDN U9151 ( .A(init), .B(e[238]), .Z(n5843) );
  AND U9152 ( .A(n5844), .B(n5845), .Z(n5842) );
  NAND U9153 ( .A(n4897), .B(ereg[237]), .Z(n5845) );
  NAND U9154 ( .A(n4892), .B(ereg[238]), .Z(n5844) );
  NAND U9155 ( .A(n5846), .B(n5847), .Z(n3620) );
  NANDN U9156 ( .A(init), .B(e[239]), .Z(n5847) );
  AND U9157 ( .A(n5848), .B(n5849), .Z(n5846) );
  NAND U9158 ( .A(n4897), .B(ereg[238]), .Z(n5849) );
  NAND U9159 ( .A(n4892), .B(ereg[239]), .Z(n5848) );
  NAND U9160 ( .A(n5850), .B(n5851), .Z(n3619) );
  NANDN U9161 ( .A(init), .B(e[240]), .Z(n5851) );
  AND U9162 ( .A(n5852), .B(n5853), .Z(n5850) );
  NAND U9163 ( .A(n4897), .B(ereg[239]), .Z(n5853) );
  NAND U9164 ( .A(n4892), .B(ereg[240]), .Z(n5852) );
  NAND U9165 ( .A(n5854), .B(n5855), .Z(n3618) );
  NANDN U9166 ( .A(init), .B(e[241]), .Z(n5855) );
  AND U9167 ( .A(n5856), .B(n5857), .Z(n5854) );
  NAND U9168 ( .A(n4897), .B(ereg[240]), .Z(n5857) );
  NAND U9169 ( .A(n4892), .B(ereg[241]), .Z(n5856) );
  NAND U9170 ( .A(n5858), .B(n5859), .Z(n3617) );
  NANDN U9171 ( .A(init), .B(e[242]), .Z(n5859) );
  AND U9172 ( .A(n5860), .B(n5861), .Z(n5858) );
  NAND U9173 ( .A(n4897), .B(ereg[241]), .Z(n5861) );
  NAND U9174 ( .A(n4892), .B(ereg[242]), .Z(n5860) );
  NAND U9175 ( .A(n5862), .B(n5863), .Z(n3616) );
  NANDN U9176 ( .A(init), .B(e[243]), .Z(n5863) );
  AND U9177 ( .A(n5864), .B(n5865), .Z(n5862) );
  NAND U9178 ( .A(n4897), .B(ereg[242]), .Z(n5865) );
  NAND U9179 ( .A(n4892), .B(ereg[243]), .Z(n5864) );
  NAND U9180 ( .A(n5866), .B(n5867), .Z(n3615) );
  NANDN U9181 ( .A(init), .B(e[244]), .Z(n5867) );
  AND U9182 ( .A(n5868), .B(n5869), .Z(n5866) );
  NAND U9183 ( .A(n4897), .B(ereg[243]), .Z(n5869) );
  NAND U9184 ( .A(n4892), .B(ereg[244]), .Z(n5868) );
  NAND U9185 ( .A(n5870), .B(n5871), .Z(n3614) );
  NANDN U9186 ( .A(init), .B(e[245]), .Z(n5871) );
  AND U9187 ( .A(n5872), .B(n5873), .Z(n5870) );
  NAND U9188 ( .A(n4897), .B(ereg[244]), .Z(n5873) );
  NAND U9189 ( .A(n4892), .B(ereg[245]), .Z(n5872) );
  NAND U9190 ( .A(n5874), .B(n5875), .Z(n3613) );
  NANDN U9191 ( .A(init), .B(e[246]), .Z(n5875) );
  AND U9192 ( .A(n5876), .B(n5877), .Z(n5874) );
  NAND U9193 ( .A(n4897), .B(ereg[245]), .Z(n5877) );
  NAND U9194 ( .A(n4892), .B(ereg[246]), .Z(n5876) );
  NAND U9195 ( .A(n5878), .B(n5879), .Z(n3612) );
  NANDN U9196 ( .A(init), .B(e[247]), .Z(n5879) );
  AND U9197 ( .A(n5880), .B(n5881), .Z(n5878) );
  NAND U9198 ( .A(n4897), .B(ereg[246]), .Z(n5881) );
  NAND U9199 ( .A(n4892), .B(ereg[247]), .Z(n5880) );
  NAND U9200 ( .A(n5882), .B(n5883), .Z(n3611) );
  NANDN U9201 ( .A(init), .B(e[248]), .Z(n5883) );
  AND U9202 ( .A(n5884), .B(n5885), .Z(n5882) );
  NAND U9203 ( .A(n4897), .B(ereg[247]), .Z(n5885) );
  NAND U9204 ( .A(n4892), .B(ereg[248]), .Z(n5884) );
  NAND U9205 ( .A(n5886), .B(n5887), .Z(n3610) );
  NANDN U9206 ( .A(init), .B(e[249]), .Z(n5887) );
  AND U9207 ( .A(n5888), .B(n5889), .Z(n5886) );
  NAND U9208 ( .A(n4897), .B(ereg[248]), .Z(n5889) );
  NAND U9209 ( .A(n4892), .B(ereg[249]), .Z(n5888) );
  NAND U9210 ( .A(n5890), .B(n5891), .Z(n3609) );
  NANDN U9211 ( .A(init), .B(e[250]), .Z(n5891) );
  AND U9212 ( .A(n5892), .B(n5893), .Z(n5890) );
  NAND U9213 ( .A(n4897), .B(ereg[249]), .Z(n5893) );
  NAND U9214 ( .A(n4892), .B(ereg[250]), .Z(n5892) );
  NAND U9215 ( .A(n5894), .B(n5895), .Z(n3608) );
  NANDN U9216 ( .A(init), .B(e[251]), .Z(n5895) );
  AND U9217 ( .A(n5896), .B(n5897), .Z(n5894) );
  NAND U9218 ( .A(n4897), .B(ereg[250]), .Z(n5897) );
  NAND U9219 ( .A(n4892), .B(ereg[251]), .Z(n5896) );
  NAND U9220 ( .A(n5898), .B(n5899), .Z(n3607) );
  NANDN U9221 ( .A(init), .B(e[252]), .Z(n5899) );
  AND U9222 ( .A(n5900), .B(n5901), .Z(n5898) );
  NAND U9223 ( .A(n4897), .B(ereg[251]), .Z(n5901) );
  NAND U9224 ( .A(n4892), .B(ereg[252]), .Z(n5900) );
  NAND U9225 ( .A(n5902), .B(n5903), .Z(n3606) );
  NANDN U9226 ( .A(init), .B(e[253]), .Z(n5903) );
  AND U9227 ( .A(n5904), .B(n5905), .Z(n5902) );
  NAND U9228 ( .A(n4897), .B(ereg[252]), .Z(n5905) );
  NAND U9229 ( .A(n4892), .B(ereg[253]), .Z(n5904) );
  NAND U9230 ( .A(n5906), .B(n5907), .Z(n3605) );
  NANDN U9231 ( .A(init), .B(e[254]), .Z(n5907) );
  AND U9232 ( .A(n5908), .B(n5909), .Z(n5906) );
  NAND U9233 ( .A(n4897), .B(ereg[253]), .Z(n5909) );
  NAND U9234 ( .A(n4892), .B(ereg[254]), .Z(n5908) );
  NAND U9235 ( .A(n5910), .B(n5911), .Z(n3604) );
  NANDN U9236 ( .A(init), .B(e[255]), .Z(n5911) );
  AND U9237 ( .A(n5912), .B(n5913), .Z(n5910) );
  NAND U9238 ( .A(n4897), .B(ereg[254]), .Z(n5913) );
  NOR U9239 ( .A(n5914), .B(n4892), .Z(n4897) );
  NAND U9240 ( .A(n4892), .B(ereg[255]), .Z(n5912) );
  NANDN U9241 ( .A(n3863), .B(n5915), .Z(n4892) );
  NANDN U9242 ( .A(start_in[1023]), .B(init), .Z(n5915) );
  NOR U9243 ( .A(n4377), .B(mul_pow), .Z(n3863) );
  NAND U9244 ( .A(n5916), .B(n4543), .Z(n3603) );
  NANDN U9245 ( .A(init), .B(m[255]), .Z(n4543) );
  AND U9246 ( .A(n5917), .B(n5918), .Z(n5916) );
  NAND U9247 ( .A(n5919), .B(o[255]), .Z(n5918) );
  NANDN U9248 ( .A(n5920), .B(creg[255]), .Z(n5917) );
  NAND U9249 ( .A(n5921), .B(n4887), .Z(n3602) );
  NANDN U9250 ( .A(init), .B(m[0]), .Z(n4887) );
  AND U9251 ( .A(n5922), .B(n5923), .Z(n5921) );
  NAND U9252 ( .A(n5919), .B(o[0]), .Z(n5923) );
  NANDN U9253 ( .A(n5920), .B(creg[0]), .Z(n5922) );
  NAND U9254 ( .A(n5924), .B(n4665), .Z(n3601) );
  NANDN U9255 ( .A(init), .B(m[1]), .Z(n4665) );
  AND U9256 ( .A(n5925), .B(n5926), .Z(n5924) );
  NAND U9257 ( .A(n5919), .B(o[1]), .Z(n5926) );
  NANDN U9258 ( .A(n5920), .B(creg[1]), .Z(n5925) );
  NAND U9259 ( .A(n5927), .B(n4531), .Z(n3600) );
  NANDN U9260 ( .A(init), .B(m[2]), .Z(n4531) );
  AND U9261 ( .A(n5928), .B(n5929), .Z(n5927) );
  NAND U9262 ( .A(n5919), .B(o[2]), .Z(n5929) );
  NANDN U9263 ( .A(n5920), .B(creg[2]), .Z(n5928) );
  NAND U9264 ( .A(n5930), .B(n4509), .Z(n3599) );
  NANDN U9265 ( .A(init), .B(m[3]), .Z(n4509) );
  AND U9266 ( .A(n5931), .B(n5932), .Z(n5930) );
  NAND U9267 ( .A(n5919), .B(o[3]), .Z(n5932) );
  NANDN U9268 ( .A(n5920), .B(creg[3]), .Z(n5931) );
  NAND U9269 ( .A(n5933), .B(n4487), .Z(n3598) );
  NANDN U9270 ( .A(init), .B(m[4]), .Z(n4487) );
  AND U9271 ( .A(n5934), .B(n5935), .Z(n5933) );
  NAND U9272 ( .A(n5919), .B(o[4]), .Z(n5935) );
  NANDN U9273 ( .A(n5920), .B(creg[4]), .Z(n5934) );
  NAND U9274 ( .A(n5936), .B(n4465), .Z(n3597) );
  NANDN U9275 ( .A(init), .B(m[5]), .Z(n4465) );
  AND U9276 ( .A(n5937), .B(n5938), .Z(n5936) );
  NAND U9277 ( .A(n5919), .B(o[5]), .Z(n5938) );
  NANDN U9278 ( .A(n5920), .B(creg[5]), .Z(n5937) );
  NAND U9279 ( .A(n5939), .B(n4443), .Z(n3596) );
  NANDN U9280 ( .A(init), .B(m[6]), .Z(n4443) );
  AND U9281 ( .A(n5940), .B(n5941), .Z(n5939) );
  NAND U9282 ( .A(n5919), .B(o[6]), .Z(n5941) );
  NANDN U9283 ( .A(n5920), .B(creg[6]), .Z(n5940) );
  NAND U9284 ( .A(n5942), .B(n4421), .Z(n3595) );
  NANDN U9285 ( .A(init), .B(m[7]), .Z(n4421) );
  AND U9286 ( .A(n5943), .B(n5944), .Z(n5942) );
  NAND U9287 ( .A(n5919), .B(o[7]), .Z(n5944) );
  NANDN U9288 ( .A(n5920), .B(creg[7]), .Z(n5943) );
  NAND U9289 ( .A(n5945), .B(n4399), .Z(n3594) );
  NANDN U9290 ( .A(init), .B(m[8]), .Z(n4399) );
  AND U9291 ( .A(n5946), .B(n5947), .Z(n5945) );
  NAND U9292 ( .A(n5919), .B(o[8]), .Z(n5947) );
  NANDN U9293 ( .A(n5920), .B(creg[8]), .Z(n5946) );
  NAND U9294 ( .A(n5948), .B(n4376), .Z(n3593) );
  NANDN U9295 ( .A(init), .B(m[9]), .Z(n4376) );
  AND U9296 ( .A(n5949), .B(n5950), .Z(n5948) );
  NAND U9297 ( .A(n5919), .B(o[9]), .Z(n5950) );
  NANDN U9298 ( .A(n5920), .B(creg[9]), .Z(n5949) );
  NAND U9299 ( .A(n5951), .B(n4865), .Z(n3592) );
  NANDN U9300 ( .A(init), .B(m[10]), .Z(n4865) );
  AND U9301 ( .A(n5952), .B(n5953), .Z(n5951) );
  NAND U9302 ( .A(n5919), .B(o[10]), .Z(n5953) );
  NANDN U9303 ( .A(n5920), .B(creg[10]), .Z(n5952) );
  NAND U9304 ( .A(n5954), .B(n4843), .Z(n3591) );
  NANDN U9305 ( .A(init), .B(m[11]), .Z(n4843) );
  AND U9306 ( .A(n5955), .B(n5956), .Z(n5954) );
  NAND U9307 ( .A(n5919), .B(o[11]), .Z(n5956) );
  NANDN U9308 ( .A(n5920), .B(creg[11]), .Z(n5955) );
  NAND U9309 ( .A(n5957), .B(n4821), .Z(n3590) );
  NANDN U9310 ( .A(init), .B(m[12]), .Z(n4821) );
  AND U9311 ( .A(n5958), .B(n5959), .Z(n5957) );
  NAND U9312 ( .A(n5919), .B(o[12]), .Z(n5959) );
  NANDN U9313 ( .A(n5920), .B(creg[12]), .Z(n5958) );
  NAND U9314 ( .A(n5960), .B(n4799), .Z(n3589) );
  NANDN U9315 ( .A(init), .B(m[13]), .Z(n4799) );
  AND U9316 ( .A(n5961), .B(n5962), .Z(n5960) );
  NAND U9317 ( .A(n5919), .B(o[13]), .Z(n5962) );
  NANDN U9318 ( .A(n5920), .B(creg[13]), .Z(n5961) );
  NAND U9319 ( .A(n5963), .B(n4777), .Z(n3588) );
  NANDN U9320 ( .A(init), .B(m[14]), .Z(n4777) );
  AND U9321 ( .A(n5964), .B(n5965), .Z(n5963) );
  NAND U9322 ( .A(n5919), .B(o[14]), .Z(n5965) );
  NANDN U9323 ( .A(n5920), .B(creg[14]), .Z(n5964) );
  NAND U9324 ( .A(n5966), .B(n4755), .Z(n3587) );
  NANDN U9325 ( .A(init), .B(m[15]), .Z(n4755) );
  AND U9326 ( .A(n5967), .B(n5968), .Z(n5966) );
  NAND U9327 ( .A(n5919), .B(o[15]), .Z(n5968) );
  NANDN U9328 ( .A(n5920), .B(creg[15]), .Z(n5967) );
  NAND U9329 ( .A(n5969), .B(n4733), .Z(n3586) );
  NANDN U9330 ( .A(init), .B(m[16]), .Z(n4733) );
  AND U9331 ( .A(n5970), .B(n5971), .Z(n5969) );
  NAND U9332 ( .A(n5919), .B(o[16]), .Z(n5971) );
  NANDN U9333 ( .A(n5920), .B(creg[16]), .Z(n5970) );
  NAND U9334 ( .A(n5972), .B(n4711), .Z(n3585) );
  NANDN U9335 ( .A(init), .B(m[17]), .Z(n4711) );
  AND U9336 ( .A(n5973), .B(n5974), .Z(n5972) );
  NAND U9337 ( .A(n5919), .B(o[17]), .Z(n5974) );
  NANDN U9338 ( .A(n5920), .B(creg[17]), .Z(n5973) );
  NAND U9339 ( .A(n5975), .B(n4689), .Z(n3584) );
  NANDN U9340 ( .A(init), .B(m[18]), .Z(n4689) );
  AND U9341 ( .A(n5976), .B(n5977), .Z(n5975) );
  NAND U9342 ( .A(n5919), .B(o[18]), .Z(n5977) );
  NANDN U9343 ( .A(n5920), .B(creg[18]), .Z(n5976) );
  NAND U9344 ( .A(n5978), .B(n4667), .Z(n3583) );
  NANDN U9345 ( .A(init), .B(m[19]), .Z(n4667) );
  AND U9346 ( .A(n5979), .B(n5980), .Z(n5978) );
  NAND U9347 ( .A(n5919), .B(o[19]), .Z(n5980) );
  NANDN U9348 ( .A(n5920), .B(creg[19]), .Z(n5979) );
  NAND U9349 ( .A(n5981), .B(n4643), .Z(n3582) );
  NANDN U9350 ( .A(init), .B(m[20]), .Z(n4643) );
  AND U9351 ( .A(n5982), .B(n5983), .Z(n5981) );
  NAND U9352 ( .A(n5919), .B(o[20]), .Z(n5983) );
  NANDN U9353 ( .A(n5920), .B(creg[20]), .Z(n5982) );
  NAND U9354 ( .A(n5984), .B(n4621), .Z(n3581) );
  NANDN U9355 ( .A(init), .B(m[21]), .Z(n4621) );
  AND U9356 ( .A(n5985), .B(n5986), .Z(n5984) );
  NAND U9357 ( .A(n5919), .B(o[21]), .Z(n5986) );
  NANDN U9358 ( .A(n5920), .B(creg[21]), .Z(n5985) );
  NAND U9359 ( .A(n5987), .B(n4599), .Z(n3580) );
  NANDN U9360 ( .A(init), .B(m[22]), .Z(n4599) );
  AND U9361 ( .A(n5988), .B(n5989), .Z(n5987) );
  NAND U9362 ( .A(n5919), .B(o[22]), .Z(n5989) );
  NANDN U9363 ( .A(n5920), .B(creg[22]), .Z(n5988) );
  NAND U9364 ( .A(n5990), .B(n4577), .Z(n3579) );
  NANDN U9365 ( .A(init), .B(m[23]), .Z(n4577) );
  AND U9366 ( .A(n5991), .B(n5992), .Z(n5990) );
  NAND U9367 ( .A(n5919), .B(o[23]), .Z(n5992) );
  NANDN U9368 ( .A(n5920), .B(creg[23]), .Z(n5991) );
  NAND U9369 ( .A(n5993), .B(n4555), .Z(n3578) );
  NANDN U9370 ( .A(init), .B(m[24]), .Z(n4555) );
  AND U9371 ( .A(n5994), .B(n5995), .Z(n5993) );
  NAND U9372 ( .A(n5919), .B(o[24]), .Z(n5995) );
  NANDN U9373 ( .A(n5920), .B(creg[24]), .Z(n5994) );
  NAND U9374 ( .A(n5996), .B(n4541), .Z(n3577) );
  NANDN U9375 ( .A(init), .B(m[25]), .Z(n4541) );
  AND U9376 ( .A(n5997), .B(n5998), .Z(n5996) );
  NAND U9377 ( .A(n5919), .B(o[25]), .Z(n5998) );
  NANDN U9378 ( .A(n5920), .B(creg[25]), .Z(n5997) );
  NAND U9379 ( .A(n5999), .B(n4539), .Z(n3576) );
  NANDN U9380 ( .A(init), .B(m[26]), .Z(n4539) );
  AND U9381 ( .A(n6000), .B(n6001), .Z(n5999) );
  NAND U9382 ( .A(n5919), .B(o[26]), .Z(n6001) );
  NANDN U9383 ( .A(n5920), .B(creg[26]), .Z(n6000) );
  NAND U9384 ( .A(n6002), .B(n4537), .Z(n3575) );
  NANDN U9385 ( .A(init), .B(m[27]), .Z(n4537) );
  AND U9386 ( .A(n6003), .B(n6004), .Z(n6002) );
  NAND U9387 ( .A(n5919), .B(o[27]), .Z(n6004) );
  NANDN U9388 ( .A(n5920), .B(creg[27]), .Z(n6003) );
  NAND U9389 ( .A(n6005), .B(n4535), .Z(n3574) );
  NANDN U9390 ( .A(init), .B(m[28]), .Z(n4535) );
  AND U9391 ( .A(n6006), .B(n6007), .Z(n6005) );
  NAND U9392 ( .A(n5919), .B(o[28]), .Z(n6007) );
  NANDN U9393 ( .A(n5920), .B(creg[28]), .Z(n6006) );
  NAND U9394 ( .A(n6008), .B(n4533), .Z(n3573) );
  NANDN U9395 ( .A(init), .B(m[29]), .Z(n4533) );
  AND U9396 ( .A(n6009), .B(n6010), .Z(n6008) );
  NAND U9397 ( .A(n5919), .B(o[29]), .Z(n6010) );
  NANDN U9398 ( .A(n5920), .B(creg[29]), .Z(n6009) );
  NAND U9399 ( .A(n6011), .B(n4529), .Z(n3572) );
  NANDN U9400 ( .A(init), .B(m[30]), .Z(n4529) );
  AND U9401 ( .A(n6012), .B(n6013), .Z(n6011) );
  NAND U9402 ( .A(n5919), .B(o[30]), .Z(n6013) );
  NANDN U9403 ( .A(n5920), .B(creg[30]), .Z(n6012) );
  NAND U9404 ( .A(n6014), .B(n4527), .Z(n3571) );
  NANDN U9405 ( .A(init), .B(m[31]), .Z(n4527) );
  AND U9406 ( .A(n6015), .B(n6016), .Z(n6014) );
  NAND U9407 ( .A(n5919), .B(o[31]), .Z(n6016) );
  NANDN U9408 ( .A(n5920), .B(creg[31]), .Z(n6015) );
  NAND U9409 ( .A(n6017), .B(n4525), .Z(n3570) );
  NANDN U9410 ( .A(init), .B(m[32]), .Z(n4525) );
  AND U9411 ( .A(n6018), .B(n6019), .Z(n6017) );
  NAND U9412 ( .A(n5919), .B(o[32]), .Z(n6019) );
  NANDN U9413 ( .A(n5920), .B(creg[32]), .Z(n6018) );
  NAND U9414 ( .A(n6020), .B(n4523), .Z(n3569) );
  NANDN U9415 ( .A(init), .B(m[33]), .Z(n4523) );
  AND U9416 ( .A(n6021), .B(n6022), .Z(n6020) );
  NAND U9417 ( .A(n5919), .B(o[33]), .Z(n6022) );
  NANDN U9418 ( .A(n5920), .B(creg[33]), .Z(n6021) );
  NAND U9419 ( .A(n6023), .B(n4521), .Z(n3568) );
  NANDN U9420 ( .A(init), .B(m[34]), .Z(n4521) );
  AND U9421 ( .A(n6024), .B(n6025), .Z(n6023) );
  NAND U9422 ( .A(n5919), .B(o[34]), .Z(n6025) );
  NANDN U9423 ( .A(n5920), .B(creg[34]), .Z(n6024) );
  NAND U9424 ( .A(n6026), .B(n4519), .Z(n3567) );
  NANDN U9425 ( .A(init), .B(m[35]), .Z(n4519) );
  AND U9426 ( .A(n6027), .B(n6028), .Z(n6026) );
  NAND U9427 ( .A(n5919), .B(o[35]), .Z(n6028) );
  NANDN U9428 ( .A(n5920), .B(creg[35]), .Z(n6027) );
  NAND U9429 ( .A(n6029), .B(n4517), .Z(n3566) );
  NANDN U9430 ( .A(init), .B(m[36]), .Z(n4517) );
  AND U9431 ( .A(n6030), .B(n6031), .Z(n6029) );
  NAND U9432 ( .A(n5919), .B(o[36]), .Z(n6031) );
  NANDN U9433 ( .A(n5920), .B(creg[36]), .Z(n6030) );
  NAND U9434 ( .A(n6032), .B(n4515), .Z(n3565) );
  NANDN U9435 ( .A(init), .B(m[37]), .Z(n4515) );
  AND U9436 ( .A(n6033), .B(n6034), .Z(n6032) );
  NAND U9437 ( .A(n5919), .B(o[37]), .Z(n6034) );
  NANDN U9438 ( .A(n5920), .B(creg[37]), .Z(n6033) );
  NAND U9439 ( .A(n6035), .B(n4513), .Z(n3564) );
  NANDN U9440 ( .A(init), .B(m[38]), .Z(n4513) );
  AND U9441 ( .A(n6036), .B(n6037), .Z(n6035) );
  NAND U9442 ( .A(n5919), .B(o[38]), .Z(n6037) );
  NANDN U9443 ( .A(n5920), .B(creg[38]), .Z(n6036) );
  NAND U9444 ( .A(n6038), .B(n4511), .Z(n3563) );
  NANDN U9445 ( .A(init), .B(m[39]), .Z(n4511) );
  AND U9446 ( .A(n6039), .B(n6040), .Z(n6038) );
  NAND U9447 ( .A(n5919), .B(o[39]), .Z(n6040) );
  NANDN U9448 ( .A(n5920), .B(creg[39]), .Z(n6039) );
  NAND U9449 ( .A(n6041), .B(n4507), .Z(n3562) );
  NANDN U9450 ( .A(init), .B(m[40]), .Z(n4507) );
  AND U9451 ( .A(n6042), .B(n6043), .Z(n6041) );
  NAND U9452 ( .A(n5919), .B(o[40]), .Z(n6043) );
  NANDN U9453 ( .A(n5920), .B(creg[40]), .Z(n6042) );
  NAND U9454 ( .A(n6044), .B(n4505), .Z(n3561) );
  NANDN U9455 ( .A(init), .B(m[41]), .Z(n4505) );
  AND U9456 ( .A(n6045), .B(n6046), .Z(n6044) );
  NAND U9457 ( .A(n5919), .B(o[41]), .Z(n6046) );
  NANDN U9458 ( .A(n5920), .B(creg[41]), .Z(n6045) );
  NAND U9459 ( .A(n6047), .B(n4503), .Z(n3560) );
  NANDN U9460 ( .A(init), .B(m[42]), .Z(n4503) );
  AND U9461 ( .A(n6048), .B(n6049), .Z(n6047) );
  NAND U9462 ( .A(n5919), .B(o[42]), .Z(n6049) );
  NANDN U9463 ( .A(n5920), .B(creg[42]), .Z(n6048) );
  NAND U9464 ( .A(n6050), .B(n4501), .Z(n3559) );
  NANDN U9465 ( .A(init), .B(m[43]), .Z(n4501) );
  AND U9466 ( .A(n6051), .B(n6052), .Z(n6050) );
  NAND U9467 ( .A(n5919), .B(o[43]), .Z(n6052) );
  NANDN U9468 ( .A(n5920), .B(creg[43]), .Z(n6051) );
  NAND U9469 ( .A(n6053), .B(n4499), .Z(n3558) );
  NANDN U9470 ( .A(init), .B(m[44]), .Z(n4499) );
  AND U9471 ( .A(n6054), .B(n6055), .Z(n6053) );
  NAND U9472 ( .A(n5919), .B(o[44]), .Z(n6055) );
  NANDN U9473 ( .A(n5920), .B(creg[44]), .Z(n6054) );
  NAND U9474 ( .A(n6056), .B(n4497), .Z(n3557) );
  NANDN U9475 ( .A(init), .B(m[45]), .Z(n4497) );
  AND U9476 ( .A(n6057), .B(n6058), .Z(n6056) );
  NAND U9477 ( .A(n5919), .B(o[45]), .Z(n6058) );
  NANDN U9478 ( .A(n5920), .B(creg[45]), .Z(n6057) );
  NAND U9479 ( .A(n6059), .B(n4495), .Z(n3556) );
  NANDN U9480 ( .A(init), .B(m[46]), .Z(n4495) );
  AND U9481 ( .A(n6060), .B(n6061), .Z(n6059) );
  NAND U9482 ( .A(n5919), .B(o[46]), .Z(n6061) );
  NANDN U9483 ( .A(n5920), .B(creg[46]), .Z(n6060) );
  NAND U9484 ( .A(n6062), .B(n4493), .Z(n3555) );
  NANDN U9485 ( .A(init), .B(m[47]), .Z(n4493) );
  AND U9486 ( .A(n6063), .B(n6064), .Z(n6062) );
  NAND U9487 ( .A(n5919), .B(o[47]), .Z(n6064) );
  NANDN U9488 ( .A(n5920), .B(creg[47]), .Z(n6063) );
  NAND U9489 ( .A(n6065), .B(n4491), .Z(n3554) );
  NANDN U9490 ( .A(init), .B(m[48]), .Z(n4491) );
  AND U9491 ( .A(n6066), .B(n6067), .Z(n6065) );
  NAND U9492 ( .A(n5919), .B(o[48]), .Z(n6067) );
  NANDN U9493 ( .A(n5920), .B(creg[48]), .Z(n6066) );
  NAND U9494 ( .A(n6068), .B(n4489), .Z(n3553) );
  NANDN U9495 ( .A(init), .B(m[49]), .Z(n4489) );
  AND U9496 ( .A(n6069), .B(n6070), .Z(n6068) );
  NAND U9497 ( .A(n5919), .B(o[49]), .Z(n6070) );
  NANDN U9498 ( .A(n5920), .B(creg[49]), .Z(n6069) );
  NAND U9499 ( .A(n6071), .B(n4485), .Z(n3552) );
  NANDN U9500 ( .A(init), .B(m[50]), .Z(n4485) );
  AND U9501 ( .A(n6072), .B(n6073), .Z(n6071) );
  NAND U9502 ( .A(n5919), .B(o[50]), .Z(n6073) );
  NANDN U9503 ( .A(n5920), .B(creg[50]), .Z(n6072) );
  NAND U9504 ( .A(n6074), .B(n4483), .Z(n3551) );
  NANDN U9505 ( .A(init), .B(m[51]), .Z(n4483) );
  AND U9506 ( .A(n6075), .B(n6076), .Z(n6074) );
  NAND U9507 ( .A(n5919), .B(o[51]), .Z(n6076) );
  NANDN U9508 ( .A(n5920), .B(creg[51]), .Z(n6075) );
  NAND U9509 ( .A(n6077), .B(n4481), .Z(n3550) );
  NANDN U9510 ( .A(init), .B(m[52]), .Z(n4481) );
  AND U9511 ( .A(n6078), .B(n6079), .Z(n6077) );
  NAND U9512 ( .A(n5919), .B(o[52]), .Z(n6079) );
  NANDN U9513 ( .A(n5920), .B(creg[52]), .Z(n6078) );
  NAND U9514 ( .A(n6080), .B(n4479), .Z(n3549) );
  NANDN U9515 ( .A(init), .B(m[53]), .Z(n4479) );
  AND U9516 ( .A(n6081), .B(n6082), .Z(n6080) );
  NAND U9517 ( .A(n5919), .B(o[53]), .Z(n6082) );
  NANDN U9518 ( .A(n5920), .B(creg[53]), .Z(n6081) );
  NAND U9519 ( .A(n6083), .B(n4477), .Z(n3548) );
  NANDN U9520 ( .A(init), .B(m[54]), .Z(n4477) );
  AND U9521 ( .A(n6084), .B(n6085), .Z(n6083) );
  NAND U9522 ( .A(n5919), .B(o[54]), .Z(n6085) );
  NANDN U9523 ( .A(n5920), .B(creg[54]), .Z(n6084) );
  NAND U9524 ( .A(n6086), .B(n4475), .Z(n3547) );
  NANDN U9525 ( .A(init), .B(m[55]), .Z(n4475) );
  AND U9526 ( .A(n6087), .B(n6088), .Z(n6086) );
  NAND U9527 ( .A(n5919), .B(o[55]), .Z(n6088) );
  NANDN U9528 ( .A(n5920), .B(creg[55]), .Z(n6087) );
  NAND U9529 ( .A(n6089), .B(n4473), .Z(n3546) );
  NANDN U9530 ( .A(init), .B(m[56]), .Z(n4473) );
  AND U9531 ( .A(n6090), .B(n6091), .Z(n6089) );
  NAND U9532 ( .A(n5919), .B(o[56]), .Z(n6091) );
  NANDN U9533 ( .A(n5920), .B(creg[56]), .Z(n6090) );
  NAND U9534 ( .A(n6092), .B(n4471), .Z(n3545) );
  NANDN U9535 ( .A(init), .B(m[57]), .Z(n4471) );
  AND U9536 ( .A(n6093), .B(n6094), .Z(n6092) );
  NAND U9537 ( .A(n5919), .B(o[57]), .Z(n6094) );
  NANDN U9538 ( .A(n5920), .B(creg[57]), .Z(n6093) );
  NAND U9539 ( .A(n6095), .B(n4469), .Z(n3544) );
  NANDN U9540 ( .A(init), .B(m[58]), .Z(n4469) );
  AND U9541 ( .A(n6096), .B(n6097), .Z(n6095) );
  NAND U9542 ( .A(n5919), .B(o[58]), .Z(n6097) );
  NANDN U9543 ( .A(n5920), .B(creg[58]), .Z(n6096) );
  NAND U9544 ( .A(n6098), .B(n4467), .Z(n3543) );
  NANDN U9545 ( .A(init), .B(m[59]), .Z(n4467) );
  AND U9546 ( .A(n6099), .B(n6100), .Z(n6098) );
  NAND U9547 ( .A(n5919), .B(o[59]), .Z(n6100) );
  NANDN U9548 ( .A(n5920), .B(creg[59]), .Z(n6099) );
  NAND U9549 ( .A(n6101), .B(n4463), .Z(n3542) );
  NANDN U9550 ( .A(init), .B(m[60]), .Z(n4463) );
  AND U9551 ( .A(n6102), .B(n6103), .Z(n6101) );
  NAND U9552 ( .A(n5919), .B(o[60]), .Z(n6103) );
  NANDN U9553 ( .A(n5920), .B(creg[60]), .Z(n6102) );
  NAND U9554 ( .A(n6104), .B(n4461), .Z(n3541) );
  NANDN U9555 ( .A(init), .B(m[61]), .Z(n4461) );
  AND U9556 ( .A(n6105), .B(n6106), .Z(n6104) );
  NAND U9557 ( .A(n5919), .B(o[61]), .Z(n6106) );
  NANDN U9558 ( .A(n5920), .B(creg[61]), .Z(n6105) );
  NAND U9559 ( .A(n6107), .B(n4459), .Z(n3540) );
  NANDN U9560 ( .A(init), .B(m[62]), .Z(n4459) );
  AND U9561 ( .A(n6108), .B(n6109), .Z(n6107) );
  NAND U9562 ( .A(n5919), .B(o[62]), .Z(n6109) );
  NANDN U9563 ( .A(n5920), .B(creg[62]), .Z(n6108) );
  NAND U9564 ( .A(n6110), .B(n4457), .Z(n3539) );
  NANDN U9565 ( .A(init), .B(m[63]), .Z(n4457) );
  AND U9566 ( .A(n6111), .B(n6112), .Z(n6110) );
  NAND U9567 ( .A(n5919), .B(o[63]), .Z(n6112) );
  NANDN U9568 ( .A(n5920), .B(creg[63]), .Z(n6111) );
  NAND U9569 ( .A(n6113), .B(n4455), .Z(n3538) );
  NANDN U9570 ( .A(init), .B(m[64]), .Z(n4455) );
  AND U9571 ( .A(n6114), .B(n6115), .Z(n6113) );
  NAND U9572 ( .A(n5919), .B(o[64]), .Z(n6115) );
  NANDN U9573 ( .A(n5920), .B(creg[64]), .Z(n6114) );
  NAND U9574 ( .A(n6116), .B(n4453), .Z(n3537) );
  NANDN U9575 ( .A(init), .B(m[65]), .Z(n4453) );
  AND U9576 ( .A(n6117), .B(n6118), .Z(n6116) );
  NAND U9577 ( .A(n5919), .B(o[65]), .Z(n6118) );
  NANDN U9578 ( .A(n5920), .B(creg[65]), .Z(n6117) );
  NAND U9579 ( .A(n6119), .B(n4451), .Z(n3536) );
  NANDN U9580 ( .A(init), .B(m[66]), .Z(n4451) );
  AND U9581 ( .A(n6120), .B(n6121), .Z(n6119) );
  NAND U9582 ( .A(n5919), .B(o[66]), .Z(n6121) );
  NANDN U9583 ( .A(n5920), .B(creg[66]), .Z(n6120) );
  NAND U9584 ( .A(n6122), .B(n4449), .Z(n3535) );
  NANDN U9585 ( .A(init), .B(m[67]), .Z(n4449) );
  AND U9586 ( .A(n6123), .B(n6124), .Z(n6122) );
  NAND U9587 ( .A(n5919), .B(o[67]), .Z(n6124) );
  NANDN U9588 ( .A(n5920), .B(creg[67]), .Z(n6123) );
  NAND U9589 ( .A(n6125), .B(n4447), .Z(n3534) );
  NANDN U9590 ( .A(init), .B(m[68]), .Z(n4447) );
  AND U9591 ( .A(n6126), .B(n6127), .Z(n6125) );
  NAND U9592 ( .A(n5919), .B(o[68]), .Z(n6127) );
  NANDN U9593 ( .A(n5920), .B(creg[68]), .Z(n6126) );
  NAND U9594 ( .A(n6128), .B(n4445), .Z(n3533) );
  NANDN U9595 ( .A(init), .B(m[69]), .Z(n4445) );
  AND U9596 ( .A(n6129), .B(n6130), .Z(n6128) );
  NAND U9597 ( .A(n5919), .B(o[69]), .Z(n6130) );
  NANDN U9598 ( .A(n5920), .B(creg[69]), .Z(n6129) );
  NAND U9599 ( .A(n6131), .B(n4441), .Z(n3532) );
  NANDN U9600 ( .A(init), .B(m[70]), .Z(n4441) );
  AND U9601 ( .A(n6132), .B(n6133), .Z(n6131) );
  NAND U9602 ( .A(n5919), .B(o[70]), .Z(n6133) );
  NANDN U9603 ( .A(n5920), .B(creg[70]), .Z(n6132) );
  NAND U9604 ( .A(n6134), .B(n4439), .Z(n3531) );
  NANDN U9605 ( .A(init), .B(m[71]), .Z(n4439) );
  AND U9606 ( .A(n6135), .B(n6136), .Z(n6134) );
  NAND U9607 ( .A(n5919), .B(o[71]), .Z(n6136) );
  NANDN U9608 ( .A(n5920), .B(creg[71]), .Z(n6135) );
  NAND U9609 ( .A(n6137), .B(n4437), .Z(n3530) );
  NANDN U9610 ( .A(init), .B(m[72]), .Z(n4437) );
  AND U9611 ( .A(n6138), .B(n6139), .Z(n6137) );
  NAND U9612 ( .A(n5919), .B(o[72]), .Z(n6139) );
  NANDN U9613 ( .A(n5920), .B(creg[72]), .Z(n6138) );
  NAND U9614 ( .A(n6140), .B(n4435), .Z(n3529) );
  NANDN U9615 ( .A(init), .B(m[73]), .Z(n4435) );
  AND U9616 ( .A(n6141), .B(n6142), .Z(n6140) );
  NAND U9617 ( .A(n5919), .B(o[73]), .Z(n6142) );
  NANDN U9618 ( .A(n5920), .B(creg[73]), .Z(n6141) );
  NAND U9619 ( .A(n6143), .B(n4433), .Z(n3528) );
  NANDN U9620 ( .A(init), .B(m[74]), .Z(n4433) );
  AND U9621 ( .A(n6144), .B(n6145), .Z(n6143) );
  NAND U9622 ( .A(n5919), .B(o[74]), .Z(n6145) );
  NANDN U9623 ( .A(n5920), .B(creg[74]), .Z(n6144) );
  NAND U9624 ( .A(n6146), .B(n4431), .Z(n3527) );
  NANDN U9625 ( .A(init), .B(m[75]), .Z(n4431) );
  AND U9626 ( .A(n6147), .B(n6148), .Z(n6146) );
  NAND U9627 ( .A(n5919), .B(o[75]), .Z(n6148) );
  NANDN U9628 ( .A(n5920), .B(creg[75]), .Z(n6147) );
  NAND U9629 ( .A(n6149), .B(n4429), .Z(n3526) );
  NANDN U9630 ( .A(init), .B(m[76]), .Z(n4429) );
  AND U9631 ( .A(n6150), .B(n6151), .Z(n6149) );
  NAND U9632 ( .A(n5919), .B(o[76]), .Z(n6151) );
  NANDN U9633 ( .A(n5920), .B(creg[76]), .Z(n6150) );
  NAND U9634 ( .A(n6152), .B(n4427), .Z(n3525) );
  NANDN U9635 ( .A(init), .B(m[77]), .Z(n4427) );
  AND U9636 ( .A(n6153), .B(n6154), .Z(n6152) );
  NAND U9637 ( .A(n5919), .B(o[77]), .Z(n6154) );
  NANDN U9638 ( .A(n5920), .B(creg[77]), .Z(n6153) );
  NAND U9639 ( .A(n6155), .B(n4425), .Z(n3524) );
  NANDN U9640 ( .A(init), .B(m[78]), .Z(n4425) );
  AND U9641 ( .A(n6156), .B(n6157), .Z(n6155) );
  NAND U9642 ( .A(n5919), .B(o[78]), .Z(n6157) );
  NANDN U9643 ( .A(n5920), .B(creg[78]), .Z(n6156) );
  NAND U9644 ( .A(n6158), .B(n4423), .Z(n3523) );
  NANDN U9645 ( .A(init), .B(m[79]), .Z(n4423) );
  AND U9646 ( .A(n6159), .B(n6160), .Z(n6158) );
  NAND U9647 ( .A(n5919), .B(o[79]), .Z(n6160) );
  NANDN U9648 ( .A(n5920), .B(creg[79]), .Z(n6159) );
  NAND U9649 ( .A(n6161), .B(n4419), .Z(n3522) );
  NANDN U9650 ( .A(init), .B(m[80]), .Z(n4419) );
  AND U9651 ( .A(n6162), .B(n6163), .Z(n6161) );
  NAND U9652 ( .A(n5919), .B(o[80]), .Z(n6163) );
  NANDN U9653 ( .A(n5920), .B(creg[80]), .Z(n6162) );
  NAND U9654 ( .A(n6164), .B(n4417), .Z(n3521) );
  NANDN U9655 ( .A(init), .B(m[81]), .Z(n4417) );
  AND U9656 ( .A(n6165), .B(n6166), .Z(n6164) );
  NAND U9657 ( .A(n5919), .B(o[81]), .Z(n6166) );
  NANDN U9658 ( .A(n5920), .B(creg[81]), .Z(n6165) );
  NAND U9659 ( .A(n6167), .B(n4415), .Z(n3520) );
  NANDN U9660 ( .A(init), .B(m[82]), .Z(n4415) );
  AND U9661 ( .A(n6168), .B(n6169), .Z(n6167) );
  NAND U9662 ( .A(n5919), .B(o[82]), .Z(n6169) );
  NANDN U9663 ( .A(n5920), .B(creg[82]), .Z(n6168) );
  NAND U9664 ( .A(n6170), .B(n4413), .Z(n3519) );
  NANDN U9665 ( .A(init), .B(m[83]), .Z(n4413) );
  AND U9666 ( .A(n6171), .B(n6172), .Z(n6170) );
  NAND U9667 ( .A(n5919), .B(o[83]), .Z(n6172) );
  NANDN U9668 ( .A(n5920), .B(creg[83]), .Z(n6171) );
  NAND U9669 ( .A(n6173), .B(n4411), .Z(n3518) );
  NANDN U9670 ( .A(init), .B(m[84]), .Z(n4411) );
  AND U9671 ( .A(n6174), .B(n6175), .Z(n6173) );
  NAND U9672 ( .A(n5919), .B(o[84]), .Z(n6175) );
  NANDN U9673 ( .A(n5920), .B(creg[84]), .Z(n6174) );
  NAND U9674 ( .A(n6176), .B(n4409), .Z(n3517) );
  NANDN U9675 ( .A(init), .B(m[85]), .Z(n4409) );
  AND U9676 ( .A(n6177), .B(n6178), .Z(n6176) );
  NAND U9677 ( .A(n5919), .B(o[85]), .Z(n6178) );
  NANDN U9678 ( .A(n5920), .B(creg[85]), .Z(n6177) );
  NAND U9679 ( .A(n6179), .B(n4407), .Z(n3516) );
  NANDN U9680 ( .A(init), .B(m[86]), .Z(n4407) );
  AND U9681 ( .A(n6180), .B(n6181), .Z(n6179) );
  NAND U9682 ( .A(n5919), .B(o[86]), .Z(n6181) );
  NANDN U9683 ( .A(n5920), .B(creg[86]), .Z(n6180) );
  NAND U9684 ( .A(n6182), .B(n4405), .Z(n3515) );
  NANDN U9685 ( .A(init), .B(m[87]), .Z(n4405) );
  AND U9686 ( .A(n6183), .B(n6184), .Z(n6182) );
  NAND U9687 ( .A(n5919), .B(o[87]), .Z(n6184) );
  NANDN U9688 ( .A(n5920), .B(creg[87]), .Z(n6183) );
  NAND U9689 ( .A(n6185), .B(n4403), .Z(n3514) );
  NANDN U9690 ( .A(init), .B(m[88]), .Z(n4403) );
  AND U9691 ( .A(n6186), .B(n6187), .Z(n6185) );
  NAND U9692 ( .A(n5919), .B(o[88]), .Z(n6187) );
  NANDN U9693 ( .A(n5920), .B(creg[88]), .Z(n6186) );
  NAND U9694 ( .A(n6188), .B(n4401), .Z(n3513) );
  NANDN U9695 ( .A(init), .B(m[89]), .Z(n4401) );
  AND U9696 ( .A(n6189), .B(n6190), .Z(n6188) );
  NAND U9697 ( .A(n5919), .B(o[89]), .Z(n6190) );
  NANDN U9698 ( .A(n5920), .B(creg[89]), .Z(n6189) );
  NAND U9699 ( .A(n6191), .B(n4397), .Z(n3512) );
  NANDN U9700 ( .A(init), .B(m[90]), .Z(n4397) );
  AND U9701 ( .A(n6192), .B(n6193), .Z(n6191) );
  NAND U9702 ( .A(n5919), .B(o[90]), .Z(n6193) );
  NANDN U9703 ( .A(n5920), .B(creg[90]), .Z(n6192) );
  NAND U9704 ( .A(n6194), .B(n4395), .Z(n3511) );
  NANDN U9705 ( .A(init), .B(m[91]), .Z(n4395) );
  AND U9706 ( .A(n6195), .B(n6196), .Z(n6194) );
  NAND U9707 ( .A(n5919), .B(o[91]), .Z(n6196) );
  NANDN U9708 ( .A(n5920), .B(creg[91]), .Z(n6195) );
  NAND U9709 ( .A(n6197), .B(n4393), .Z(n3510) );
  NANDN U9710 ( .A(init), .B(m[92]), .Z(n4393) );
  AND U9711 ( .A(n6198), .B(n6199), .Z(n6197) );
  NAND U9712 ( .A(n5919), .B(o[92]), .Z(n6199) );
  NANDN U9713 ( .A(n5920), .B(creg[92]), .Z(n6198) );
  NAND U9714 ( .A(n6200), .B(n4391), .Z(n3509) );
  NANDN U9715 ( .A(init), .B(m[93]), .Z(n4391) );
  AND U9716 ( .A(n6201), .B(n6202), .Z(n6200) );
  NAND U9717 ( .A(n5919), .B(o[93]), .Z(n6202) );
  NANDN U9718 ( .A(n5920), .B(creg[93]), .Z(n6201) );
  NAND U9719 ( .A(n6203), .B(n4389), .Z(n3508) );
  NANDN U9720 ( .A(init), .B(m[94]), .Z(n4389) );
  AND U9721 ( .A(n6204), .B(n6205), .Z(n6203) );
  NAND U9722 ( .A(n5919), .B(o[94]), .Z(n6205) );
  NANDN U9723 ( .A(n5920), .B(creg[94]), .Z(n6204) );
  NAND U9724 ( .A(n6206), .B(n4387), .Z(n3507) );
  NANDN U9725 ( .A(init), .B(m[95]), .Z(n4387) );
  AND U9726 ( .A(n6207), .B(n6208), .Z(n6206) );
  NAND U9727 ( .A(n5919), .B(o[95]), .Z(n6208) );
  NANDN U9728 ( .A(n5920), .B(creg[95]), .Z(n6207) );
  NAND U9729 ( .A(n6209), .B(n4385), .Z(n3506) );
  NANDN U9730 ( .A(init), .B(m[96]), .Z(n4385) );
  AND U9731 ( .A(n6210), .B(n6211), .Z(n6209) );
  NAND U9732 ( .A(n5919), .B(o[96]), .Z(n6211) );
  NANDN U9733 ( .A(n5920), .B(creg[96]), .Z(n6210) );
  NAND U9734 ( .A(n6212), .B(n4383), .Z(n3505) );
  NANDN U9735 ( .A(init), .B(m[97]), .Z(n4383) );
  AND U9736 ( .A(n6213), .B(n6214), .Z(n6212) );
  NAND U9737 ( .A(n5919), .B(o[97]), .Z(n6214) );
  NANDN U9738 ( .A(n5920), .B(creg[97]), .Z(n6213) );
  NAND U9739 ( .A(n6215), .B(n4381), .Z(n3504) );
  NANDN U9740 ( .A(init), .B(m[98]), .Z(n4381) );
  AND U9741 ( .A(n6216), .B(n6217), .Z(n6215) );
  NAND U9742 ( .A(n5919), .B(o[98]), .Z(n6217) );
  NANDN U9743 ( .A(n5920), .B(creg[98]), .Z(n6216) );
  NAND U9744 ( .A(n6218), .B(n4379), .Z(n3503) );
  NANDN U9745 ( .A(init), .B(m[99]), .Z(n4379) );
  AND U9746 ( .A(n6219), .B(n6220), .Z(n6218) );
  NAND U9747 ( .A(n5919), .B(o[99]), .Z(n6220) );
  NANDN U9748 ( .A(n5920), .B(creg[99]), .Z(n6219) );
  NAND U9749 ( .A(n6221), .B(n4885), .Z(n3502) );
  NANDN U9750 ( .A(init), .B(m[100]), .Z(n4885) );
  AND U9751 ( .A(n6222), .B(n6223), .Z(n6221) );
  NAND U9752 ( .A(n5919), .B(o[100]), .Z(n6223) );
  NANDN U9753 ( .A(n5920), .B(creg[100]), .Z(n6222) );
  NAND U9754 ( .A(n6224), .B(n4883), .Z(n3501) );
  NANDN U9755 ( .A(init), .B(m[101]), .Z(n4883) );
  AND U9756 ( .A(n6225), .B(n6226), .Z(n6224) );
  NAND U9757 ( .A(n5919), .B(o[101]), .Z(n6226) );
  NANDN U9758 ( .A(n5920), .B(creg[101]), .Z(n6225) );
  NAND U9759 ( .A(n6227), .B(n4881), .Z(n3500) );
  NANDN U9760 ( .A(init), .B(m[102]), .Z(n4881) );
  AND U9761 ( .A(n6228), .B(n6229), .Z(n6227) );
  NAND U9762 ( .A(n5919), .B(o[102]), .Z(n6229) );
  NANDN U9763 ( .A(n5920), .B(creg[102]), .Z(n6228) );
  NAND U9764 ( .A(n6230), .B(n4879), .Z(n3499) );
  NANDN U9765 ( .A(init), .B(m[103]), .Z(n4879) );
  AND U9766 ( .A(n6231), .B(n6232), .Z(n6230) );
  NAND U9767 ( .A(n5919), .B(o[103]), .Z(n6232) );
  NANDN U9768 ( .A(n5920), .B(creg[103]), .Z(n6231) );
  NAND U9769 ( .A(n6233), .B(n4877), .Z(n3498) );
  NANDN U9770 ( .A(init), .B(m[104]), .Z(n4877) );
  AND U9771 ( .A(n6234), .B(n6235), .Z(n6233) );
  NAND U9772 ( .A(n5919), .B(o[104]), .Z(n6235) );
  NANDN U9773 ( .A(n5920), .B(creg[104]), .Z(n6234) );
  NAND U9774 ( .A(n6236), .B(n4875), .Z(n3497) );
  NANDN U9775 ( .A(init), .B(m[105]), .Z(n4875) );
  AND U9776 ( .A(n6237), .B(n6238), .Z(n6236) );
  NAND U9777 ( .A(n5919), .B(o[105]), .Z(n6238) );
  NANDN U9778 ( .A(n5920), .B(creg[105]), .Z(n6237) );
  NAND U9779 ( .A(n6239), .B(n4873), .Z(n3496) );
  NANDN U9780 ( .A(init), .B(m[106]), .Z(n4873) );
  AND U9781 ( .A(n6240), .B(n6241), .Z(n6239) );
  NAND U9782 ( .A(n5919), .B(o[106]), .Z(n6241) );
  NANDN U9783 ( .A(n5920), .B(creg[106]), .Z(n6240) );
  NAND U9784 ( .A(n6242), .B(n4871), .Z(n3495) );
  NANDN U9785 ( .A(init), .B(m[107]), .Z(n4871) );
  AND U9786 ( .A(n6243), .B(n6244), .Z(n6242) );
  NAND U9787 ( .A(n5919), .B(o[107]), .Z(n6244) );
  NANDN U9788 ( .A(n5920), .B(creg[107]), .Z(n6243) );
  NAND U9789 ( .A(n6245), .B(n4869), .Z(n3494) );
  NANDN U9790 ( .A(init), .B(m[108]), .Z(n4869) );
  AND U9791 ( .A(n6246), .B(n6247), .Z(n6245) );
  NAND U9792 ( .A(n5919), .B(o[108]), .Z(n6247) );
  NANDN U9793 ( .A(n5920), .B(creg[108]), .Z(n6246) );
  NAND U9794 ( .A(n6248), .B(n4867), .Z(n3493) );
  NANDN U9795 ( .A(init), .B(m[109]), .Z(n4867) );
  AND U9796 ( .A(n6249), .B(n6250), .Z(n6248) );
  NAND U9797 ( .A(n5919), .B(o[109]), .Z(n6250) );
  NANDN U9798 ( .A(n5920), .B(creg[109]), .Z(n6249) );
  NAND U9799 ( .A(n6251), .B(n4863), .Z(n3492) );
  NANDN U9800 ( .A(init), .B(m[110]), .Z(n4863) );
  AND U9801 ( .A(n6252), .B(n6253), .Z(n6251) );
  NAND U9802 ( .A(n5919), .B(o[110]), .Z(n6253) );
  NANDN U9803 ( .A(n5920), .B(creg[110]), .Z(n6252) );
  NAND U9804 ( .A(n6254), .B(n4861), .Z(n3491) );
  NANDN U9805 ( .A(init), .B(m[111]), .Z(n4861) );
  AND U9806 ( .A(n6255), .B(n6256), .Z(n6254) );
  NAND U9807 ( .A(n5919), .B(o[111]), .Z(n6256) );
  NANDN U9808 ( .A(n5920), .B(creg[111]), .Z(n6255) );
  NAND U9809 ( .A(n6257), .B(n4859), .Z(n3490) );
  NANDN U9810 ( .A(init), .B(m[112]), .Z(n4859) );
  AND U9811 ( .A(n6258), .B(n6259), .Z(n6257) );
  NAND U9812 ( .A(n5919), .B(o[112]), .Z(n6259) );
  NANDN U9813 ( .A(n5920), .B(creg[112]), .Z(n6258) );
  NAND U9814 ( .A(n6260), .B(n4857), .Z(n3489) );
  NANDN U9815 ( .A(init), .B(m[113]), .Z(n4857) );
  AND U9816 ( .A(n6261), .B(n6262), .Z(n6260) );
  NAND U9817 ( .A(n5919), .B(o[113]), .Z(n6262) );
  NANDN U9818 ( .A(n5920), .B(creg[113]), .Z(n6261) );
  NAND U9819 ( .A(n6263), .B(n4855), .Z(n3488) );
  NANDN U9820 ( .A(init), .B(m[114]), .Z(n4855) );
  AND U9821 ( .A(n6264), .B(n6265), .Z(n6263) );
  NAND U9822 ( .A(n5919), .B(o[114]), .Z(n6265) );
  NANDN U9823 ( .A(n5920), .B(creg[114]), .Z(n6264) );
  NAND U9824 ( .A(n6266), .B(n4853), .Z(n3487) );
  NANDN U9825 ( .A(init), .B(m[115]), .Z(n4853) );
  AND U9826 ( .A(n6267), .B(n6268), .Z(n6266) );
  NAND U9827 ( .A(n5919), .B(o[115]), .Z(n6268) );
  NANDN U9828 ( .A(n5920), .B(creg[115]), .Z(n6267) );
  NAND U9829 ( .A(n6269), .B(n4851), .Z(n3486) );
  NANDN U9830 ( .A(init), .B(m[116]), .Z(n4851) );
  AND U9831 ( .A(n6270), .B(n6271), .Z(n6269) );
  NAND U9832 ( .A(n5919), .B(o[116]), .Z(n6271) );
  NANDN U9833 ( .A(n5920), .B(creg[116]), .Z(n6270) );
  NAND U9834 ( .A(n6272), .B(n4849), .Z(n3485) );
  NANDN U9835 ( .A(init), .B(m[117]), .Z(n4849) );
  AND U9836 ( .A(n6273), .B(n6274), .Z(n6272) );
  NAND U9837 ( .A(n5919), .B(o[117]), .Z(n6274) );
  NANDN U9838 ( .A(n5920), .B(creg[117]), .Z(n6273) );
  NAND U9839 ( .A(n6275), .B(n4847), .Z(n3484) );
  NANDN U9840 ( .A(init), .B(m[118]), .Z(n4847) );
  AND U9841 ( .A(n6276), .B(n6277), .Z(n6275) );
  NAND U9842 ( .A(n5919), .B(o[118]), .Z(n6277) );
  NANDN U9843 ( .A(n5920), .B(creg[118]), .Z(n6276) );
  NAND U9844 ( .A(n6278), .B(n4845), .Z(n3483) );
  NANDN U9845 ( .A(init), .B(m[119]), .Z(n4845) );
  AND U9846 ( .A(n6279), .B(n6280), .Z(n6278) );
  NAND U9847 ( .A(n5919), .B(o[119]), .Z(n6280) );
  NANDN U9848 ( .A(n5920), .B(creg[119]), .Z(n6279) );
  NAND U9849 ( .A(n6281), .B(n4841), .Z(n3482) );
  NANDN U9850 ( .A(init), .B(m[120]), .Z(n4841) );
  AND U9851 ( .A(n6282), .B(n6283), .Z(n6281) );
  NAND U9852 ( .A(n5919), .B(o[120]), .Z(n6283) );
  NANDN U9853 ( .A(n5920), .B(creg[120]), .Z(n6282) );
  NAND U9854 ( .A(n6284), .B(n4839), .Z(n3481) );
  NANDN U9855 ( .A(init), .B(m[121]), .Z(n4839) );
  AND U9856 ( .A(n6285), .B(n6286), .Z(n6284) );
  NAND U9857 ( .A(n5919), .B(o[121]), .Z(n6286) );
  NANDN U9858 ( .A(n5920), .B(creg[121]), .Z(n6285) );
  NAND U9859 ( .A(n6287), .B(n4837), .Z(n3480) );
  NANDN U9860 ( .A(init), .B(m[122]), .Z(n4837) );
  AND U9861 ( .A(n6288), .B(n6289), .Z(n6287) );
  NAND U9862 ( .A(n5919), .B(o[122]), .Z(n6289) );
  NANDN U9863 ( .A(n5920), .B(creg[122]), .Z(n6288) );
  NAND U9864 ( .A(n6290), .B(n4835), .Z(n3479) );
  NANDN U9865 ( .A(init), .B(m[123]), .Z(n4835) );
  AND U9866 ( .A(n6291), .B(n6292), .Z(n6290) );
  NAND U9867 ( .A(n5919), .B(o[123]), .Z(n6292) );
  NANDN U9868 ( .A(n5920), .B(creg[123]), .Z(n6291) );
  NAND U9869 ( .A(n6293), .B(n4833), .Z(n3478) );
  NANDN U9870 ( .A(init), .B(m[124]), .Z(n4833) );
  AND U9871 ( .A(n6294), .B(n6295), .Z(n6293) );
  NAND U9872 ( .A(n5919), .B(o[124]), .Z(n6295) );
  NANDN U9873 ( .A(n5920), .B(creg[124]), .Z(n6294) );
  NAND U9874 ( .A(n6296), .B(n4831), .Z(n3477) );
  NANDN U9875 ( .A(init), .B(m[125]), .Z(n4831) );
  AND U9876 ( .A(n6297), .B(n6298), .Z(n6296) );
  NAND U9877 ( .A(n5919), .B(o[125]), .Z(n6298) );
  NANDN U9878 ( .A(n5920), .B(creg[125]), .Z(n6297) );
  NAND U9879 ( .A(n6299), .B(n4829), .Z(n3476) );
  NANDN U9880 ( .A(init), .B(m[126]), .Z(n4829) );
  AND U9881 ( .A(n6300), .B(n6301), .Z(n6299) );
  NAND U9882 ( .A(n5919), .B(o[126]), .Z(n6301) );
  NANDN U9883 ( .A(n5920), .B(creg[126]), .Z(n6300) );
  NAND U9884 ( .A(n6302), .B(n4827), .Z(n3475) );
  NANDN U9885 ( .A(init), .B(m[127]), .Z(n4827) );
  AND U9886 ( .A(n6303), .B(n6304), .Z(n6302) );
  NAND U9887 ( .A(n5919), .B(o[127]), .Z(n6304) );
  NANDN U9888 ( .A(n5920), .B(creg[127]), .Z(n6303) );
  NAND U9889 ( .A(n6305), .B(n4825), .Z(n3474) );
  NANDN U9890 ( .A(init), .B(m[128]), .Z(n4825) );
  AND U9891 ( .A(n6306), .B(n6307), .Z(n6305) );
  NAND U9892 ( .A(n5919), .B(o[128]), .Z(n6307) );
  NANDN U9893 ( .A(n5920), .B(creg[128]), .Z(n6306) );
  NAND U9894 ( .A(n6308), .B(n4823), .Z(n3473) );
  NANDN U9895 ( .A(init), .B(m[129]), .Z(n4823) );
  AND U9896 ( .A(n6309), .B(n6310), .Z(n6308) );
  NAND U9897 ( .A(n5919), .B(o[129]), .Z(n6310) );
  NANDN U9898 ( .A(n5920), .B(creg[129]), .Z(n6309) );
  NAND U9899 ( .A(n6311), .B(n4819), .Z(n3472) );
  NANDN U9900 ( .A(init), .B(m[130]), .Z(n4819) );
  AND U9901 ( .A(n6312), .B(n6313), .Z(n6311) );
  NAND U9902 ( .A(n5919), .B(o[130]), .Z(n6313) );
  NANDN U9903 ( .A(n5920), .B(creg[130]), .Z(n6312) );
  NAND U9904 ( .A(n6314), .B(n4817), .Z(n3471) );
  NANDN U9905 ( .A(init), .B(m[131]), .Z(n4817) );
  AND U9906 ( .A(n6315), .B(n6316), .Z(n6314) );
  NAND U9907 ( .A(n5919), .B(o[131]), .Z(n6316) );
  NANDN U9908 ( .A(n5920), .B(creg[131]), .Z(n6315) );
  NAND U9909 ( .A(n6317), .B(n4815), .Z(n3470) );
  NANDN U9910 ( .A(init), .B(m[132]), .Z(n4815) );
  AND U9911 ( .A(n6318), .B(n6319), .Z(n6317) );
  NAND U9912 ( .A(n5919), .B(o[132]), .Z(n6319) );
  NANDN U9913 ( .A(n5920), .B(creg[132]), .Z(n6318) );
  NAND U9914 ( .A(n6320), .B(n4813), .Z(n3469) );
  NANDN U9915 ( .A(init), .B(m[133]), .Z(n4813) );
  AND U9916 ( .A(n6321), .B(n6322), .Z(n6320) );
  NAND U9917 ( .A(n5919), .B(o[133]), .Z(n6322) );
  NANDN U9918 ( .A(n5920), .B(creg[133]), .Z(n6321) );
  NAND U9919 ( .A(n6323), .B(n4811), .Z(n3468) );
  NANDN U9920 ( .A(init), .B(m[134]), .Z(n4811) );
  AND U9921 ( .A(n6324), .B(n6325), .Z(n6323) );
  NAND U9922 ( .A(n5919), .B(o[134]), .Z(n6325) );
  NANDN U9923 ( .A(n5920), .B(creg[134]), .Z(n6324) );
  NAND U9924 ( .A(n6326), .B(n4809), .Z(n3467) );
  NANDN U9925 ( .A(init), .B(m[135]), .Z(n4809) );
  AND U9926 ( .A(n6327), .B(n6328), .Z(n6326) );
  NAND U9927 ( .A(n5919), .B(o[135]), .Z(n6328) );
  NANDN U9928 ( .A(n5920), .B(creg[135]), .Z(n6327) );
  NAND U9929 ( .A(n6329), .B(n4807), .Z(n3466) );
  NANDN U9930 ( .A(init), .B(m[136]), .Z(n4807) );
  AND U9931 ( .A(n6330), .B(n6331), .Z(n6329) );
  NAND U9932 ( .A(n5919), .B(o[136]), .Z(n6331) );
  NANDN U9933 ( .A(n5920), .B(creg[136]), .Z(n6330) );
  NAND U9934 ( .A(n6332), .B(n4805), .Z(n3465) );
  NANDN U9935 ( .A(init), .B(m[137]), .Z(n4805) );
  AND U9936 ( .A(n6333), .B(n6334), .Z(n6332) );
  NAND U9937 ( .A(n5919), .B(o[137]), .Z(n6334) );
  NANDN U9938 ( .A(n5920), .B(creg[137]), .Z(n6333) );
  NAND U9939 ( .A(n6335), .B(n4803), .Z(n3464) );
  NANDN U9940 ( .A(init), .B(m[138]), .Z(n4803) );
  AND U9941 ( .A(n6336), .B(n6337), .Z(n6335) );
  NAND U9942 ( .A(n5919), .B(o[138]), .Z(n6337) );
  NANDN U9943 ( .A(n5920), .B(creg[138]), .Z(n6336) );
  NAND U9944 ( .A(n6338), .B(n4801), .Z(n3463) );
  NANDN U9945 ( .A(init), .B(m[139]), .Z(n4801) );
  AND U9946 ( .A(n6339), .B(n6340), .Z(n6338) );
  NAND U9947 ( .A(n5919), .B(o[139]), .Z(n6340) );
  NANDN U9948 ( .A(n5920), .B(creg[139]), .Z(n6339) );
  NAND U9949 ( .A(n6341), .B(n4797), .Z(n3462) );
  NANDN U9950 ( .A(init), .B(m[140]), .Z(n4797) );
  AND U9951 ( .A(n6342), .B(n6343), .Z(n6341) );
  NAND U9952 ( .A(n5919), .B(o[140]), .Z(n6343) );
  NANDN U9953 ( .A(n5920), .B(creg[140]), .Z(n6342) );
  NAND U9954 ( .A(n6344), .B(n4795), .Z(n3461) );
  NANDN U9955 ( .A(init), .B(m[141]), .Z(n4795) );
  AND U9956 ( .A(n6345), .B(n6346), .Z(n6344) );
  NAND U9957 ( .A(n5919), .B(o[141]), .Z(n6346) );
  NANDN U9958 ( .A(n5920), .B(creg[141]), .Z(n6345) );
  NAND U9959 ( .A(n6347), .B(n4793), .Z(n3460) );
  NANDN U9960 ( .A(init), .B(m[142]), .Z(n4793) );
  AND U9961 ( .A(n6348), .B(n6349), .Z(n6347) );
  NAND U9962 ( .A(n5919), .B(o[142]), .Z(n6349) );
  NANDN U9963 ( .A(n5920), .B(creg[142]), .Z(n6348) );
  NAND U9964 ( .A(n6350), .B(n4791), .Z(n3459) );
  NANDN U9965 ( .A(init), .B(m[143]), .Z(n4791) );
  AND U9966 ( .A(n6351), .B(n6352), .Z(n6350) );
  NAND U9967 ( .A(n5919), .B(o[143]), .Z(n6352) );
  NANDN U9968 ( .A(n5920), .B(creg[143]), .Z(n6351) );
  NAND U9969 ( .A(n6353), .B(n4789), .Z(n3458) );
  NANDN U9970 ( .A(init), .B(m[144]), .Z(n4789) );
  AND U9971 ( .A(n6354), .B(n6355), .Z(n6353) );
  NAND U9972 ( .A(n5919), .B(o[144]), .Z(n6355) );
  NANDN U9973 ( .A(n5920), .B(creg[144]), .Z(n6354) );
  NAND U9974 ( .A(n6356), .B(n4787), .Z(n3457) );
  NANDN U9975 ( .A(init), .B(m[145]), .Z(n4787) );
  AND U9976 ( .A(n6357), .B(n6358), .Z(n6356) );
  NAND U9977 ( .A(n5919), .B(o[145]), .Z(n6358) );
  NANDN U9978 ( .A(n5920), .B(creg[145]), .Z(n6357) );
  NAND U9979 ( .A(n6359), .B(n4785), .Z(n3456) );
  NANDN U9980 ( .A(init), .B(m[146]), .Z(n4785) );
  AND U9981 ( .A(n6360), .B(n6361), .Z(n6359) );
  NAND U9982 ( .A(n5919), .B(o[146]), .Z(n6361) );
  NANDN U9983 ( .A(n5920), .B(creg[146]), .Z(n6360) );
  NAND U9984 ( .A(n6362), .B(n4783), .Z(n3455) );
  NANDN U9985 ( .A(init), .B(m[147]), .Z(n4783) );
  AND U9986 ( .A(n6363), .B(n6364), .Z(n6362) );
  NAND U9987 ( .A(n5919), .B(o[147]), .Z(n6364) );
  NANDN U9988 ( .A(n5920), .B(creg[147]), .Z(n6363) );
  NAND U9989 ( .A(n6365), .B(n4781), .Z(n3454) );
  NANDN U9990 ( .A(init), .B(m[148]), .Z(n4781) );
  AND U9991 ( .A(n6366), .B(n6367), .Z(n6365) );
  NAND U9992 ( .A(n5919), .B(o[148]), .Z(n6367) );
  NANDN U9993 ( .A(n5920), .B(creg[148]), .Z(n6366) );
  NAND U9994 ( .A(n6368), .B(n4779), .Z(n3453) );
  NANDN U9995 ( .A(init), .B(m[149]), .Z(n4779) );
  AND U9996 ( .A(n6369), .B(n6370), .Z(n6368) );
  NAND U9997 ( .A(n5919), .B(o[149]), .Z(n6370) );
  NANDN U9998 ( .A(n5920), .B(creg[149]), .Z(n6369) );
  NAND U9999 ( .A(n6371), .B(n4775), .Z(n3452) );
  NANDN U10000 ( .A(init), .B(m[150]), .Z(n4775) );
  AND U10001 ( .A(n6372), .B(n6373), .Z(n6371) );
  NAND U10002 ( .A(n5919), .B(o[150]), .Z(n6373) );
  NANDN U10003 ( .A(n5920), .B(creg[150]), .Z(n6372) );
  NAND U10004 ( .A(n6374), .B(n4773), .Z(n3451) );
  NANDN U10005 ( .A(init), .B(m[151]), .Z(n4773) );
  AND U10006 ( .A(n6375), .B(n6376), .Z(n6374) );
  NAND U10007 ( .A(n5919), .B(o[151]), .Z(n6376) );
  NANDN U10008 ( .A(n5920), .B(creg[151]), .Z(n6375) );
  NAND U10009 ( .A(n6377), .B(n4771), .Z(n3450) );
  NANDN U10010 ( .A(init), .B(m[152]), .Z(n4771) );
  AND U10011 ( .A(n6378), .B(n6379), .Z(n6377) );
  NAND U10012 ( .A(n5919), .B(o[152]), .Z(n6379) );
  NANDN U10013 ( .A(n5920), .B(creg[152]), .Z(n6378) );
  NAND U10014 ( .A(n6380), .B(n4769), .Z(n3449) );
  NANDN U10015 ( .A(init), .B(m[153]), .Z(n4769) );
  AND U10016 ( .A(n6381), .B(n6382), .Z(n6380) );
  NAND U10017 ( .A(n5919), .B(o[153]), .Z(n6382) );
  NANDN U10018 ( .A(n5920), .B(creg[153]), .Z(n6381) );
  NAND U10019 ( .A(n6383), .B(n4767), .Z(n3448) );
  NANDN U10020 ( .A(init), .B(m[154]), .Z(n4767) );
  AND U10021 ( .A(n6384), .B(n6385), .Z(n6383) );
  NAND U10022 ( .A(n5919), .B(o[154]), .Z(n6385) );
  NANDN U10023 ( .A(n5920), .B(creg[154]), .Z(n6384) );
  NAND U10024 ( .A(n6386), .B(n4765), .Z(n3447) );
  NANDN U10025 ( .A(init), .B(m[155]), .Z(n4765) );
  AND U10026 ( .A(n6387), .B(n6388), .Z(n6386) );
  NAND U10027 ( .A(n5919), .B(o[155]), .Z(n6388) );
  NANDN U10028 ( .A(n5920), .B(creg[155]), .Z(n6387) );
  NAND U10029 ( .A(n6389), .B(n4763), .Z(n3446) );
  NANDN U10030 ( .A(init), .B(m[156]), .Z(n4763) );
  AND U10031 ( .A(n6390), .B(n6391), .Z(n6389) );
  NAND U10032 ( .A(n5919), .B(o[156]), .Z(n6391) );
  NANDN U10033 ( .A(n5920), .B(creg[156]), .Z(n6390) );
  NAND U10034 ( .A(n6392), .B(n4761), .Z(n3445) );
  NANDN U10035 ( .A(init), .B(m[157]), .Z(n4761) );
  AND U10036 ( .A(n6393), .B(n6394), .Z(n6392) );
  NAND U10037 ( .A(n5919), .B(o[157]), .Z(n6394) );
  NANDN U10038 ( .A(n5920), .B(creg[157]), .Z(n6393) );
  NAND U10039 ( .A(n6395), .B(n4759), .Z(n3444) );
  NANDN U10040 ( .A(init), .B(m[158]), .Z(n4759) );
  AND U10041 ( .A(n6396), .B(n6397), .Z(n6395) );
  NAND U10042 ( .A(n5919), .B(o[158]), .Z(n6397) );
  NANDN U10043 ( .A(n5920), .B(creg[158]), .Z(n6396) );
  NAND U10044 ( .A(n6398), .B(n4757), .Z(n3443) );
  NANDN U10045 ( .A(init), .B(m[159]), .Z(n4757) );
  AND U10046 ( .A(n6399), .B(n6400), .Z(n6398) );
  NAND U10047 ( .A(n5919), .B(o[159]), .Z(n6400) );
  NANDN U10048 ( .A(n5920), .B(creg[159]), .Z(n6399) );
  NAND U10049 ( .A(n6401), .B(n4753), .Z(n3442) );
  NANDN U10050 ( .A(init), .B(m[160]), .Z(n4753) );
  AND U10051 ( .A(n6402), .B(n6403), .Z(n6401) );
  NAND U10052 ( .A(n5919), .B(o[160]), .Z(n6403) );
  NANDN U10053 ( .A(n5920), .B(creg[160]), .Z(n6402) );
  NAND U10054 ( .A(n6404), .B(n4751), .Z(n3441) );
  NANDN U10055 ( .A(init), .B(m[161]), .Z(n4751) );
  AND U10056 ( .A(n6405), .B(n6406), .Z(n6404) );
  NAND U10057 ( .A(n5919), .B(o[161]), .Z(n6406) );
  NANDN U10058 ( .A(n5920), .B(creg[161]), .Z(n6405) );
  NAND U10059 ( .A(n6407), .B(n4749), .Z(n3440) );
  NANDN U10060 ( .A(init), .B(m[162]), .Z(n4749) );
  AND U10061 ( .A(n6408), .B(n6409), .Z(n6407) );
  NAND U10062 ( .A(n5919), .B(o[162]), .Z(n6409) );
  NANDN U10063 ( .A(n5920), .B(creg[162]), .Z(n6408) );
  NAND U10064 ( .A(n6410), .B(n4747), .Z(n3439) );
  NANDN U10065 ( .A(init), .B(m[163]), .Z(n4747) );
  AND U10066 ( .A(n6411), .B(n6412), .Z(n6410) );
  NAND U10067 ( .A(n5919), .B(o[163]), .Z(n6412) );
  NANDN U10068 ( .A(n5920), .B(creg[163]), .Z(n6411) );
  NAND U10069 ( .A(n6413), .B(n4745), .Z(n3438) );
  NANDN U10070 ( .A(init), .B(m[164]), .Z(n4745) );
  AND U10071 ( .A(n6414), .B(n6415), .Z(n6413) );
  NAND U10072 ( .A(n5919), .B(o[164]), .Z(n6415) );
  NANDN U10073 ( .A(n5920), .B(creg[164]), .Z(n6414) );
  NAND U10074 ( .A(n6416), .B(n4743), .Z(n3437) );
  NANDN U10075 ( .A(init), .B(m[165]), .Z(n4743) );
  AND U10076 ( .A(n6417), .B(n6418), .Z(n6416) );
  NAND U10077 ( .A(n5919), .B(o[165]), .Z(n6418) );
  NANDN U10078 ( .A(n5920), .B(creg[165]), .Z(n6417) );
  NAND U10079 ( .A(n6419), .B(n4741), .Z(n3436) );
  NANDN U10080 ( .A(init), .B(m[166]), .Z(n4741) );
  AND U10081 ( .A(n6420), .B(n6421), .Z(n6419) );
  NAND U10082 ( .A(n5919), .B(o[166]), .Z(n6421) );
  NANDN U10083 ( .A(n5920), .B(creg[166]), .Z(n6420) );
  NAND U10084 ( .A(n6422), .B(n4739), .Z(n3435) );
  NANDN U10085 ( .A(init), .B(m[167]), .Z(n4739) );
  AND U10086 ( .A(n6423), .B(n6424), .Z(n6422) );
  NAND U10087 ( .A(n5919), .B(o[167]), .Z(n6424) );
  NANDN U10088 ( .A(n5920), .B(creg[167]), .Z(n6423) );
  NAND U10089 ( .A(n6425), .B(n4737), .Z(n3434) );
  NANDN U10090 ( .A(init), .B(m[168]), .Z(n4737) );
  AND U10091 ( .A(n6426), .B(n6427), .Z(n6425) );
  NAND U10092 ( .A(n5919), .B(o[168]), .Z(n6427) );
  NANDN U10093 ( .A(n5920), .B(creg[168]), .Z(n6426) );
  NAND U10094 ( .A(n6428), .B(n4735), .Z(n3433) );
  NANDN U10095 ( .A(init), .B(m[169]), .Z(n4735) );
  AND U10096 ( .A(n6429), .B(n6430), .Z(n6428) );
  NAND U10097 ( .A(n5919), .B(o[169]), .Z(n6430) );
  NANDN U10098 ( .A(n5920), .B(creg[169]), .Z(n6429) );
  NAND U10099 ( .A(n6431), .B(n4731), .Z(n3432) );
  NANDN U10100 ( .A(init), .B(m[170]), .Z(n4731) );
  AND U10101 ( .A(n6432), .B(n6433), .Z(n6431) );
  NAND U10102 ( .A(n5919), .B(o[170]), .Z(n6433) );
  NANDN U10103 ( .A(n5920), .B(creg[170]), .Z(n6432) );
  NAND U10104 ( .A(n6434), .B(n4729), .Z(n3431) );
  NANDN U10105 ( .A(init), .B(m[171]), .Z(n4729) );
  AND U10106 ( .A(n6435), .B(n6436), .Z(n6434) );
  NAND U10107 ( .A(n5919), .B(o[171]), .Z(n6436) );
  NANDN U10108 ( .A(n5920), .B(creg[171]), .Z(n6435) );
  NAND U10109 ( .A(n6437), .B(n4727), .Z(n3430) );
  NANDN U10110 ( .A(init), .B(m[172]), .Z(n4727) );
  AND U10111 ( .A(n6438), .B(n6439), .Z(n6437) );
  NAND U10112 ( .A(n5919), .B(o[172]), .Z(n6439) );
  NANDN U10113 ( .A(n5920), .B(creg[172]), .Z(n6438) );
  NAND U10114 ( .A(n6440), .B(n4725), .Z(n3429) );
  NANDN U10115 ( .A(init), .B(m[173]), .Z(n4725) );
  AND U10116 ( .A(n6441), .B(n6442), .Z(n6440) );
  NAND U10117 ( .A(n5919), .B(o[173]), .Z(n6442) );
  NANDN U10118 ( .A(n5920), .B(creg[173]), .Z(n6441) );
  NAND U10119 ( .A(n6443), .B(n4723), .Z(n3428) );
  NANDN U10120 ( .A(init), .B(m[174]), .Z(n4723) );
  AND U10121 ( .A(n6444), .B(n6445), .Z(n6443) );
  NAND U10122 ( .A(n5919), .B(o[174]), .Z(n6445) );
  NANDN U10123 ( .A(n5920), .B(creg[174]), .Z(n6444) );
  NAND U10124 ( .A(n6446), .B(n4721), .Z(n3427) );
  NANDN U10125 ( .A(init), .B(m[175]), .Z(n4721) );
  AND U10126 ( .A(n6447), .B(n6448), .Z(n6446) );
  NAND U10127 ( .A(n5919), .B(o[175]), .Z(n6448) );
  NANDN U10128 ( .A(n5920), .B(creg[175]), .Z(n6447) );
  NAND U10129 ( .A(n6449), .B(n4719), .Z(n3426) );
  NANDN U10130 ( .A(init), .B(m[176]), .Z(n4719) );
  AND U10131 ( .A(n6450), .B(n6451), .Z(n6449) );
  NAND U10132 ( .A(n5919), .B(o[176]), .Z(n6451) );
  NANDN U10133 ( .A(n5920), .B(creg[176]), .Z(n6450) );
  NAND U10134 ( .A(n6452), .B(n4717), .Z(n3425) );
  NANDN U10135 ( .A(init), .B(m[177]), .Z(n4717) );
  AND U10136 ( .A(n6453), .B(n6454), .Z(n6452) );
  NAND U10137 ( .A(n5919), .B(o[177]), .Z(n6454) );
  NANDN U10138 ( .A(n5920), .B(creg[177]), .Z(n6453) );
  NAND U10139 ( .A(n6455), .B(n4715), .Z(n3424) );
  NANDN U10140 ( .A(init), .B(m[178]), .Z(n4715) );
  AND U10141 ( .A(n6456), .B(n6457), .Z(n6455) );
  NAND U10142 ( .A(n5919), .B(o[178]), .Z(n6457) );
  NANDN U10143 ( .A(n5920), .B(creg[178]), .Z(n6456) );
  NAND U10144 ( .A(n6458), .B(n4713), .Z(n3423) );
  NANDN U10145 ( .A(init), .B(m[179]), .Z(n4713) );
  AND U10146 ( .A(n6459), .B(n6460), .Z(n6458) );
  NAND U10147 ( .A(n5919), .B(o[179]), .Z(n6460) );
  NANDN U10148 ( .A(n5920), .B(creg[179]), .Z(n6459) );
  NAND U10149 ( .A(n6461), .B(n4709), .Z(n3422) );
  NANDN U10150 ( .A(init), .B(m[180]), .Z(n4709) );
  AND U10151 ( .A(n6462), .B(n6463), .Z(n6461) );
  NAND U10152 ( .A(n5919), .B(o[180]), .Z(n6463) );
  NANDN U10153 ( .A(n5920), .B(creg[180]), .Z(n6462) );
  NAND U10154 ( .A(n6464), .B(n4707), .Z(n3421) );
  NANDN U10155 ( .A(init), .B(m[181]), .Z(n4707) );
  AND U10156 ( .A(n6465), .B(n6466), .Z(n6464) );
  NAND U10157 ( .A(n5919), .B(o[181]), .Z(n6466) );
  NANDN U10158 ( .A(n5920), .B(creg[181]), .Z(n6465) );
  NAND U10159 ( .A(n6467), .B(n4705), .Z(n3420) );
  NANDN U10160 ( .A(init), .B(m[182]), .Z(n4705) );
  AND U10161 ( .A(n6468), .B(n6469), .Z(n6467) );
  NAND U10162 ( .A(n5919), .B(o[182]), .Z(n6469) );
  NANDN U10163 ( .A(n5920), .B(creg[182]), .Z(n6468) );
  NAND U10164 ( .A(n6470), .B(n4703), .Z(n3419) );
  NANDN U10165 ( .A(init), .B(m[183]), .Z(n4703) );
  AND U10166 ( .A(n6471), .B(n6472), .Z(n6470) );
  NAND U10167 ( .A(n5919), .B(o[183]), .Z(n6472) );
  NANDN U10168 ( .A(n5920), .B(creg[183]), .Z(n6471) );
  NAND U10169 ( .A(n6473), .B(n4701), .Z(n3418) );
  NANDN U10170 ( .A(init), .B(m[184]), .Z(n4701) );
  AND U10171 ( .A(n6474), .B(n6475), .Z(n6473) );
  NAND U10172 ( .A(n5919), .B(o[184]), .Z(n6475) );
  NANDN U10173 ( .A(n5920), .B(creg[184]), .Z(n6474) );
  NAND U10174 ( .A(n6476), .B(n4699), .Z(n3417) );
  NANDN U10175 ( .A(init), .B(m[185]), .Z(n4699) );
  AND U10176 ( .A(n6477), .B(n6478), .Z(n6476) );
  NAND U10177 ( .A(n5919), .B(o[185]), .Z(n6478) );
  NANDN U10178 ( .A(n5920), .B(creg[185]), .Z(n6477) );
  NAND U10179 ( .A(n6479), .B(n4697), .Z(n3416) );
  NANDN U10180 ( .A(init), .B(m[186]), .Z(n4697) );
  AND U10181 ( .A(n6480), .B(n6481), .Z(n6479) );
  NAND U10182 ( .A(n5919), .B(o[186]), .Z(n6481) );
  NANDN U10183 ( .A(n5920), .B(creg[186]), .Z(n6480) );
  NAND U10184 ( .A(n6482), .B(n4695), .Z(n3415) );
  NANDN U10185 ( .A(init), .B(m[187]), .Z(n4695) );
  AND U10186 ( .A(n6483), .B(n6484), .Z(n6482) );
  NAND U10187 ( .A(n5919), .B(o[187]), .Z(n6484) );
  NANDN U10188 ( .A(n5920), .B(creg[187]), .Z(n6483) );
  NAND U10189 ( .A(n6485), .B(n4693), .Z(n3414) );
  NANDN U10190 ( .A(init), .B(m[188]), .Z(n4693) );
  AND U10191 ( .A(n6486), .B(n6487), .Z(n6485) );
  NAND U10192 ( .A(n5919), .B(o[188]), .Z(n6487) );
  NANDN U10193 ( .A(n5920), .B(creg[188]), .Z(n6486) );
  NAND U10194 ( .A(n6488), .B(n4691), .Z(n3413) );
  NANDN U10195 ( .A(init), .B(m[189]), .Z(n4691) );
  AND U10196 ( .A(n6489), .B(n6490), .Z(n6488) );
  NAND U10197 ( .A(n5919), .B(o[189]), .Z(n6490) );
  NANDN U10198 ( .A(n5920), .B(creg[189]), .Z(n6489) );
  NAND U10199 ( .A(n6491), .B(n4687), .Z(n3412) );
  NANDN U10200 ( .A(init), .B(m[190]), .Z(n4687) );
  AND U10201 ( .A(n6492), .B(n6493), .Z(n6491) );
  NAND U10202 ( .A(n5919), .B(o[190]), .Z(n6493) );
  NANDN U10203 ( .A(n5920), .B(creg[190]), .Z(n6492) );
  NAND U10204 ( .A(n6494), .B(n4685), .Z(n3411) );
  NANDN U10205 ( .A(init), .B(m[191]), .Z(n4685) );
  AND U10206 ( .A(n6495), .B(n6496), .Z(n6494) );
  NAND U10207 ( .A(n5919), .B(o[191]), .Z(n6496) );
  NANDN U10208 ( .A(n5920), .B(creg[191]), .Z(n6495) );
  NAND U10209 ( .A(n6497), .B(n4683), .Z(n3410) );
  NANDN U10210 ( .A(init), .B(m[192]), .Z(n4683) );
  AND U10211 ( .A(n6498), .B(n6499), .Z(n6497) );
  NAND U10212 ( .A(n5919), .B(o[192]), .Z(n6499) );
  NANDN U10213 ( .A(n5920), .B(creg[192]), .Z(n6498) );
  NAND U10214 ( .A(n6500), .B(n4681), .Z(n3409) );
  NANDN U10215 ( .A(init), .B(m[193]), .Z(n4681) );
  AND U10216 ( .A(n6501), .B(n6502), .Z(n6500) );
  NAND U10217 ( .A(n5919), .B(o[193]), .Z(n6502) );
  NANDN U10218 ( .A(n5920), .B(creg[193]), .Z(n6501) );
  NAND U10219 ( .A(n6503), .B(n4679), .Z(n3408) );
  NANDN U10220 ( .A(init), .B(m[194]), .Z(n4679) );
  AND U10221 ( .A(n6504), .B(n6505), .Z(n6503) );
  NAND U10222 ( .A(n5919), .B(o[194]), .Z(n6505) );
  NANDN U10223 ( .A(n5920), .B(creg[194]), .Z(n6504) );
  NAND U10224 ( .A(n6506), .B(n4677), .Z(n3407) );
  NANDN U10225 ( .A(init), .B(m[195]), .Z(n4677) );
  AND U10226 ( .A(n6507), .B(n6508), .Z(n6506) );
  NAND U10227 ( .A(n5919), .B(o[195]), .Z(n6508) );
  NANDN U10228 ( .A(n5920), .B(creg[195]), .Z(n6507) );
  NAND U10229 ( .A(n6509), .B(n4675), .Z(n3406) );
  NANDN U10230 ( .A(init), .B(m[196]), .Z(n4675) );
  AND U10231 ( .A(n6510), .B(n6511), .Z(n6509) );
  NAND U10232 ( .A(n5919), .B(o[196]), .Z(n6511) );
  NANDN U10233 ( .A(n5920), .B(creg[196]), .Z(n6510) );
  NAND U10234 ( .A(n6512), .B(n4673), .Z(n3405) );
  NANDN U10235 ( .A(init), .B(m[197]), .Z(n4673) );
  AND U10236 ( .A(n6513), .B(n6514), .Z(n6512) );
  NAND U10237 ( .A(n5919), .B(o[197]), .Z(n6514) );
  NANDN U10238 ( .A(n5920), .B(creg[197]), .Z(n6513) );
  NAND U10239 ( .A(n6515), .B(n4671), .Z(n3404) );
  NANDN U10240 ( .A(init), .B(m[198]), .Z(n4671) );
  AND U10241 ( .A(n6516), .B(n6517), .Z(n6515) );
  NAND U10242 ( .A(n5919), .B(o[198]), .Z(n6517) );
  NANDN U10243 ( .A(n5920), .B(creg[198]), .Z(n6516) );
  NAND U10244 ( .A(n6518), .B(n4669), .Z(n3403) );
  NANDN U10245 ( .A(init), .B(m[199]), .Z(n4669) );
  AND U10246 ( .A(n6519), .B(n6520), .Z(n6518) );
  NAND U10247 ( .A(n5919), .B(o[199]), .Z(n6520) );
  NANDN U10248 ( .A(n5920), .B(creg[199]), .Z(n6519) );
  NAND U10249 ( .A(n6521), .B(n4663), .Z(n3402) );
  NANDN U10250 ( .A(init), .B(m[200]), .Z(n4663) );
  AND U10251 ( .A(n6522), .B(n6523), .Z(n6521) );
  NAND U10252 ( .A(n5919), .B(o[200]), .Z(n6523) );
  NANDN U10253 ( .A(n5920), .B(creg[200]), .Z(n6522) );
  NAND U10254 ( .A(n6524), .B(n4661), .Z(n3401) );
  NANDN U10255 ( .A(init), .B(m[201]), .Z(n4661) );
  AND U10256 ( .A(n6525), .B(n6526), .Z(n6524) );
  NAND U10257 ( .A(n5919), .B(o[201]), .Z(n6526) );
  NANDN U10258 ( .A(n5920), .B(creg[201]), .Z(n6525) );
  NAND U10259 ( .A(n6527), .B(n4659), .Z(n3400) );
  NANDN U10260 ( .A(init), .B(m[202]), .Z(n4659) );
  AND U10261 ( .A(n6528), .B(n6529), .Z(n6527) );
  NAND U10262 ( .A(n5919), .B(o[202]), .Z(n6529) );
  NANDN U10263 ( .A(n5920), .B(creg[202]), .Z(n6528) );
  NAND U10264 ( .A(n6530), .B(n4657), .Z(n3399) );
  NANDN U10265 ( .A(init), .B(m[203]), .Z(n4657) );
  AND U10266 ( .A(n6531), .B(n6532), .Z(n6530) );
  NAND U10267 ( .A(n5919), .B(o[203]), .Z(n6532) );
  NANDN U10268 ( .A(n5920), .B(creg[203]), .Z(n6531) );
  NAND U10269 ( .A(n6533), .B(n4655), .Z(n3398) );
  NANDN U10270 ( .A(init), .B(m[204]), .Z(n4655) );
  AND U10271 ( .A(n6534), .B(n6535), .Z(n6533) );
  NAND U10272 ( .A(n5919), .B(o[204]), .Z(n6535) );
  NANDN U10273 ( .A(n5920), .B(creg[204]), .Z(n6534) );
  NAND U10274 ( .A(n6536), .B(n4653), .Z(n3397) );
  NANDN U10275 ( .A(init), .B(m[205]), .Z(n4653) );
  AND U10276 ( .A(n6537), .B(n6538), .Z(n6536) );
  NAND U10277 ( .A(n5919), .B(o[205]), .Z(n6538) );
  NANDN U10278 ( .A(n5920), .B(creg[205]), .Z(n6537) );
  NAND U10279 ( .A(n6539), .B(n4651), .Z(n3396) );
  NANDN U10280 ( .A(init), .B(m[206]), .Z(n4651) );
  AND U10281 ( .A(n6540), .B(n6541), .Z(n6539) );
  NAND U10282 ( .A(n5919), .B(o[206]), .Z(n6541) );
  NANDN U10283 ( .A(n5920), .B(creg[206]), .Z(n6540) );
  NAND U10284 ( .A(n6542), .B(n4649), .Z(n3395) );
  NANDN U10285 ( .A(init), .B(m[207]), .Z(n4649) );
  AND U10286 ( .A(n6543), .B(n6544), .Z(n6542) );
  NAND U10287 ( .A(n5919), .B(o[207]), .Z(n6544) );
  NANDN U10288 ( .A(n5920), .B(creg[207]), .Z(n6543) );
  NAND U10289 ( .A(n6545), .B(n4647), .Z(n3394) );
  NANDN U10290 ( .A(init), .B(m[208]), .Z(n4647) );
  AND U10291 ( .A(n6546), .B(n6547), .Z(n6545) );
  NAND U10292 ( .A(n5919), .B(o[208]), .Z(n6547) );
  NANDN U10293 ( .A(n5920), .B(creg[208]), .Z(n6546) );
  NAND U10294 ( .A(n6548), .B(n4645), .Z(n3393) );
  NANDN U10295 ( .A(init), .B(m[209]), .Z(n4645) );
  AND U10296 ( .A(n6549), .B(n6550), .Z(n6548) );
  NAND U10297 ( .A(n5919), .B(o[209]), .Z(n6550) );
  NANDN U10298 ( .A(n5920), .B(creg[209]), .Z(n6549) );
  NAND U10299 ( .A(n6551), .B(n4641), .Z(n3392) );
  NANDN U10300 ( .A(init), .B(m[210]), .Z(n4641) );
  AND U10301 ( .A(n6552), .B(n6553), .Z(n6551) );
  NAND U10302 ( .A(n5919), .B(o[210]), .Z(n6553) );
  NANDN U10303 ( .A(n5920), .B(creg[210]), .Z(n6552) );
  NAND U10304 ( .A(n6554), .B(n4639), .Z(n3391) );
  NANDN U10305 ( .A(init), .B(m[211]), .Z(n4639) );
  AND U10306 ( .A(n6555), .B(n6556), .Z(n6554) );
  NAND U10307 ( .A(n5919), .B(o[211]), .Z(n6556) );
  NANDN U10308 ( .A(n5920), .B(creg[211]), .Z(n6555) );
  NAND U10309 ( .A(n6557), .B(n4637), .Z(n3390) );
  NANDN U10310 ( .A(init), .B(m[212]), .Z(n4637) );
  AND U10311 ( .A(n6558), .B(n6559), .Z(n6557) );
  NAND U10312 ( .A(n5919), .B(o[212]), .Z(n6559) );
  NANDN U10313 ( .A(n5920), .B(creg[212]), .Z(n6558) );
  NAND U10314 ( .A(n6560), .B(n4635), .Z(n3389) );
  NANDN U10315 ( .A(init), .B(m[213]), .Z(n4635) );
  AND U10316 ( .A(n6561), .B(n6562), .Z(n6560) );
  NAND U10317 ( .A(n5919), .B(o[213]), .Z(n6562) );
  NANDN U10318 ( .A(n5920), .B(creg[213]), .Z(n6561) );
  NAND U10319 ( .A(n6563), .B(n4633), .Z(n3388) );
  NANDN U10320 ( .A(init), .B(m[214]), .Z(n4633) );
  AND U10321 ( .A(n6564), .B(n6565), .Z(n6563) );
  NAND U10322 ( .A(n5919), .B(o[214]), .Z(n6565) );
  NANDN U10323 ( .A(n5920), .B(creg[214]), .Z(n6564) );
  NAND U10324 ( .A(n6566), .B(n4631), .Z(n3387) );
  NANDN U10325 ( .A(init), .B(m[215]), .Z(n4631) );
  AND U10326 ( .A(n6567), .B(n6568), .Z(n6566) );
  NAND U10327 ( .A(n5919), .B(o[215]), .Z(n6568) );
  NANDN U10328 ( .A(n5920), .B(creg[215]), .Z(n6567) );
  NAND U10329 ( .A(n6569), .B(n4629), .Z(n3386) );
  NANDN U10330 ( .A(init), .B(m[216]), .Z(n4629) );
  AND U10331 ( .A(n6570), .B(n6571), .Z(n6569) );
  NAND U10332 ( .A(n5919), .B(o[216]), .Z(n6571) );
  NANDN U10333 ( .A(n5920), .B(creg[216]), .Z(n6570) );
  NAND U10334 ( .A(n6572), .B(n4627), .Z(n3385) );
  NANDN U10335 ( .A(init), .B(m[217]), .Z(n4627) );
  AND U10336 ( .A(n6573), .B(n6574), .Z(n6572) );
  NAND U10337 ( .A(n5919), .B(o[217]), .Z(n6574) );
  NANDN U10338 ( .A(n5920), .B(creg[217]), .Z(n6573) );
  NAND U10339 ( .A(n6575), .B(n4625), .Z(n3384) );
  NANDN U10340 ( .A(init), .B(m[218]), .Z(n4625) );
  AND U10341 ( .A(n6576), .B(n6577), .Z(n6575) );
  NAND U10342 ( .A(n5919), .B(o[218]), .Z(n6577) );
  NANDN U10343 ( .A(n5920), .B(creg[218]), .Z(n6576) );
  NAND U10344 ( .A(n6578), .B(n4623), .Z(n3383) );
  NANDN U10345 ( .A(init), .B(m[219]), .Z(n4623) );
  AND U10346 ( .A(n6579), .B(n6580), .Z(n6578) );
  NAND U10347 ( .A(n5919), .B(o[219]), .Z(n6580) );
  NANDN U10348 ( .A(n5920), .B(creg[219]), .Z(n6579) );
  NAND U10349 ( .A(n6581), .B(n4619), .Z(n3382) );
  NANDN U10350 ( .A(init), .B(m[220]), .Z(n4619) );
  AND U10351 ( .A(n6582), .B(n6583), .Z(n6581) );
  NAND U10352 ( .A(n5919), .B(o[220]), .Z(n6583) );
  NANDN U10353 ( .A(n5920), .B(creg[220]), .Z(n6582) );
  NAND U10354 ( .A(n6584), .B(n4617), .Z(n3381) );
  NANDN U10355 ( .A(init), .B(m[221]), .Z(n4617) );
  AND U10356 ( .A(n6585), .B(n6586), .Z(n6584) );
  NAND U10357 ( .A(n5919), .B(o[221]), .Z(n6586) );
  NANDN U10358 ( .A(n5920), .B(creg[221]), .Z(n6585) );
  NAND U10359 ( .A(n6587), .B(n4615), .Z(n3380) );
  NANDN U10360 ( .A(init), .B(m[222]), .Z(n4615) );
  AND U10361 ( .A(n6588), .B(n6589), .Z(n6587) );
  NAND U10362 ( .A(n5919), .B(o[222]), .Z(n6589) );
  NANDN U10363 ( .A(n5920), .B(creg[222]), .Z(n6588) );
  NAND U10364 ( .A(n6590), .B(n4613), .Z(n3379) );
  NANDN U10365 ( .A(init), .B(m[223]), .Z(n4613) );
  AND U10366 ( .A(n6591), .B(n6592), .Z(n6590) );
  NAND U10367 ( .A(n5919), .B(o[223]), .Z(n6592) );
  NANDN U10368 ( .A(n5920), .B(creg[223]), .Z(n6591) );
  NAND U10369 ( .A(n6593), .B(n4611), .Z(n3378) );
  NANDN U10370 ( .A(init), .B(m[224]), .Z(n4611) );
  AND U10371 ( .A(n6594), .B(n6595), .Z(n6593) );
  NAND U10372 ( .A(n5919), .B(o[224]), .Z(n6595) );
  NANDN U10373 ( .A(n5920), .B(creg[224]), .Z(n6594) );
  NAND U10374 ( .A(n6596), .B(n4609), .Z(n3377) );
  NANDN U10375 ( .A(init), .B(m[225]), .Z(n4609) );
  AND U10376 ( .A(n6597), .B(n6598), .Z(n6596) );
  NAND U10377 ( .A(n5919), .B(o[225]), .Z(n6598) );
  NANDN U10378 ( .A(n5920), .B(creg[225]), .Z(n6597) );
  NAND U10379 ( .A(n6599), .B(n4607), .Z(n3376) );
  NANDN U10380 ( .A(init), .B(m[226]), .Z(n4607) );
  AND U10381 ( .A(n6600), .B(n6601), .Z(n6599) );
  NAND U10382 ( .A(n5919), .B(o[226]), .Z(n6601) );
  NANDN U10383 ( .A(n5920), .B(creg[226]), .Z(n6600) );
  NAND U10384 ( .A(n6602), .B(n4605), .Z(n3375) );
  NANDN U10385 ( .A(init), .B(m[227]), .Z(n4605) );
  AND U10386 ( .A(n6603), .B(n6604), .Z(n6602) );
  NAND U10387 ( .A(n5919), .B(o[227]), .Z(n6604) );
  NANDN U10388 ( .A(n5920), .B(creg[227]), .Z(n6603) );
  NAND U10389 ( .A(n6605), .B(n4603), .Z(n3374) );
  NANDN U10390 ( .A(init), .B(m[228]), .Z(n4603) );
  AND U10391 ( .A(n6606), .B(n6607), .Z(n6605) );
  NAND U10392 ( .A(n5919), .B(o[228]), .Z(n6607) );
  NANDN U10393 ( .A(n5920), .B(creg[228]), .Z(n6606) );
  NAND U10394 ( .A(n6608), .B(n4601), .Z(n3373) );
  NANDN U10395 ( .A(init), .B(m[229]), .Z(n4601) );
  AND U10396 ( .A(n6609), .B(n6610), .Z(n6608) );
  NAND U10397 ( .A(n5919), .B(o[229]), .Z(n6610) );
  NANDN U10398 ( .A(n5920), .B(creg[229]), .Z(n6609) );
  NAND U10399 ( .A(n6611), .B(n4597), .Z(n3372) );
  NANDN U10400 ( .A(init), .B(m[230]), .Z(n4597) );
  AND U10401 ( .A(n6612), .B(n6613), .Z(n6611) );
  NAND U10402 ( .A(n5919), .B(o[230]), .Z(n6613) );
  NANDN U10403 ( .A(n5920), .B(creg[230]), .Z(n6612) );
  NAND U10404 ( .A(n6614), .B(n4595), .Z(n3371) );
  NANDN U10405 ( .A(init), .B(m[231]), .Z(n4595) );
  AND U10406 ( .A(n6615), .B(n6616), .Z(n6614) );
  NAND U10407 ( .A(n5919), .B(o[231]), .Z(n6616) );
  NANDN U10408 ( .A(n5920), .B(creg[231]), .Z(n6615) );
  NAND U10409 ( .A(n6617), .B(n4593), .Z(n3370) );
  NANDN U10410 ( .A(init), .B(m[232]), .Z(n4593) );
  AND U10411 ( .A(n6618), .B(n6619), .Z(n6617) );
  NAND U10412 ( .A(n5919), .B(o[232]), .Z(n6619) );
  NANDN U10413 ( .A(n5920), .B(creg[232]), .Z(n6618) );
  NAND U10414 ( .A(n6620), .B(n4591), .Z(n3369) );
  NANDN U10415 ( .A(init), .B(m[233]), .Z(n4591) );
  AND U10416 ( .A(n6621), .B(n6622), .Z(n6620) );
  NAND U10417 ( .A(n5919), .B(o[233]), .Z(n6622) );
  NANDN U10418 ( .A(n5920), .B(creg[233]), .Z(n6621) );
  NAND U10419 ( .A(n6623), .B(n4589), .Z(n3368) );
  NANDN U10420 ( .A(init), .B(m[234]), .Z(n4589) );
  AND U10421 ( .A(n6624), .B(n6625), .Z(n6623) );
  NAND U10422 ( .A(n5919), .B(o[234]), .Z(n6625) );
  NANDN U10423 ( .A(n5920), .B(creg[234]), .Z(n6624) );
  NAND U10424 ( .A(n6626), .B(n4587), .Z(n3367) );
  NANDN U10425 ( .A(init), .B(m[235]), .Z(n4587) );
  AND U10426 ( .A(n6627), .B(n6628), .Z(n6626) );
  NAND U10427 ( .A(n5919), .B(o[235]), .Z(n6628) );
  NANDN U10428 ( .A(n5920), .B(creg[235]), .Z(n6627) );
  NAND U10429 ( .A(n6629), .B(n4585), .Z(n3366) );
  NANDN U10430 ( .A(init), .B(m[236]), .Z(n4585) );
  AND U10431 ( .A(n6630), .B(n6631), .Z(n6629) );
  NAND U10432 ( .A(n5919), .B(o[236]), .Z(n6631) );
  NANDN U10433 ( .A(n5920), .B(creg[236]), .Z(n6630) );
  NAND U10434 ( .A(n6632), .B(n4583), .Z(n3365) );
  NANDN U10435 ( .A(init), .B(m[237]), .Z(n4583) );
  AND U10436 ( .A(n6633), .B(n6634), .Z(n6632) );
  NAND U10437 ( .A(n5919), .B(o[237]), .Z(n6634) );
  NANDN U10438 ( .A(n5920), .B(creg[237]), .Z(n6633) );
  NAND U10439 ( .A(n6635), .B(n4581), .Z(n3364) );
  NANDN U10440 ( .A(init), .B(m[238]), .Z(n4581) );
  AND U10441 ( .A(n6636), .B(n6637), .Z(n6635) );
  NAND U10442 ( .A(n5919), .B(o[238]), .Z(n6637) );
  NANDN U10443 ( .A(n5920), .B(creg[238]), .Z(n6636) );
  NAND U10444 ( .A(n6638), .B(n4579), .Z(n3363) );
  NANDN U10445 ( .A(init), .B(m[239]), .Z(n4579) );
  AND U10446 ( .A(n6639), .B(n6640), .Z(n6638) );
  NAND U10447 ( .A(n5919), .B(o[239]), .Z(n6640) );
  NANDN U10448 ( .A(n5920), .B(creg[239]), .Z(n6639) );
  NAND U10449 ( .A(n6641), .B(n4575), .Z(n3362) );
  NANDN U10450 ( .A(init), .B(m[240]), .Z(n4575) );
  AND U10451 ( .A(n6642), .B(n6643), .Z(n6641) );
  NAND U10452 ( .A(n5919), .B(o[240]), .Z(n6643) );
  NANDN U10453 ( .A(n5920), .B(creg[240]), .Z(n6642) );
  NAND U10454 ( .A(n6644), .B(n4573), .Z(n3361) );
  NANDN U10455 ( .A(init), .B(m[241]), .Z(n4573) );
  AND U10456 ( .A(n6645), .B(n6646), .Z(n6644) );
  NAND U10457 ( .A(n5919), .B(o[241]), .Z(n6646) );
  NANDN U10458 ( .A(n5920), .B(creg[241]), .Z(n6645) );
  NAND U10459 ( .A(n6647), .B(n4571), .Z(n3360) );
  NANDN U10460 ( .A(init), .B(m[242]), .Z(n4571) );
  AND U10461 ( .A(n6648), .B(n6649), .Z(n6647) );
  NAND U10462 ( .A(n5919), .B(o[242]), .Z(n6649) );
  NANDN U10463 ( .A(n5920), .B(creg[242]), .Z(n6648) );
  NAND U10464 ( .A(n6650), .B(n4569), .Z(n3359) );
  NANDN U10465 ( .A(init), .B(m[243]), .Z(n4569) );
  AND U10466 ( .A(n6651), .B(n6652), .Z(n6650) );
  NAND U10467 ( .A(n5919), .B(o[243]), .Z(n6652) );
  NANDN U10468 ( .A(n5920), .B(creg[243]), .Z(n6651) );
  NAND U10469 ( .A(n6653), .B(n4567), .Z(n3358) );
  NANDN U10470 ( .A(init), .B(m[244]), .Z(n4567) );
  AND U10471 ( .A(n6654), .B(n6655), .Z(n6653) );
  NAND U10472 ( .A(n5919), .B(o[244]), .Z(n6655) );
  NANDN U10473 ( .A(n5920), .B(creg[244]), .Z(n6654) );
  NAND U10474 ( .A(n6656), .B(n4565), .Z(n3357) );
  NANDN U10475 ( .A(init), .B(m[245]), .Z(n4565) );
  AND U10476 ( .A(n6657), .B(n6658), .Z(n6656) );
  NAND U10477 ( .A(n5919), .B(o[245]), .Z(n6658) );
  NANDN U10478 ( .A(n5920), .B(creg[245]), .Z(n6657) );
  NAND U10479 ( .A(n6659), .B(n4563), .Z(n3356) );
  NANDN U10480 ( .A(init), .B(m[246]), .Z(n4563) );
  AND U10481 ( .A(n6660), .B(n6661), .Z(n6659) );
  NAND U10482 ( .A(n5919), .B(o[246]), .Z(n6661) );
  NANDN U10483 ( .A(n5920), .B(creg[246]), .Z(n6660) );
  NAND U10484 ( .A(n6662), .B(n4561), .Z(n3355) );
  NANDN U10485 ( .A(init), .B(m[247]), .Z(n4561) );
  AND U10486 ( .A(n6663), .B(n6664), .Z(n6662) );
  NAND U10487 ( .A(n5919), .B(o[247]), .Z(n6664) );
  NANDN U10488 ( .A(n5920), .B(creg[247]), .Z(n6663) );
  NAND U10489 ( .A(n6665), .B(n4559), .Z(n3354) );
  NANDN U10490 ( .A(init), .B(m[248]), .Z(n4559) );
  AND U10491 ( .A(n6666), .B(n6667), .Z(n6665) );
  NAND U10492 ( .A(n5919), .B(o[248]), .Z(n6667) );
  NANDN U10493 ( .A(n5920), .B(creg[248]), .Z(n6666) );
  NAND U10494 ( .A(n6668), .B(n4557), .Z(n3353) );
  NANDN U10495 ( .A(init), .B(m[249]), .Z(n4557) );
  AND U10496 ( .A(n6669), .B(n6670), .Z(n6668) );
  NAND U10497 ( .A(n5919), .B(o[249]), .Z(n6670) );
  NANDN U10498 ( .A(n5920), .B(creg[249]), .Z(n6669) );
  NAND U10499 ( .A(n6671), .B(n4553), .Z(n3352) );
  NANDN U10500 ( .A(init), .B(m[250]), .Z(n4553) );
  AND U10501 ( .A(n6672), .B(n6673), .Z(n6671) );
  NAND U10502 ( .A(n5919), .B(o[250]), .Z(n6673) );
  NANDN U10503 ( .A(n5920), .B(creg[250]), .Z(n6672) );
  NAND U10504 ( .A(n6674), .B(n4551), .Z(n3351) );
  NANDN U10505 ( .A(init), .B(m[251]), .Z(n4551) );
  AND U10506 ( .A(n6675), .B(n6676), .Z(n6674) );
  NAND U10507 ( .A(n5919), .B(o[251]), .Z(n6676) );
  NANDN U10508 ( .A(n5920), .B(creg[251]), .Z(n6675) );
  NAND U10509 ( .A(n6677), .B(n4549), .Z(n3350) );
  NANDN U10510 ( .A(init), .B(m[252]), .Z(n4549) );
  AND U10511 ( .A(n6678), .B(n6679), .Z(n6677) );
  NAND U10512 ( .A(n5919), .B(o[252]), .Z(n6679) );
  NANDN U10513 ( .A(n5920), .B(creg[252]), .Z(n6678) );
  NAND U10514 ( .A(n6680), .B(n4547), .Z(n3349) );
  NANDN U10515 ( .A(init), .B(m[253]), .Z(n4547) );
  AND U10516 ( .A(n6681), .B(n6682), .Z(n6680) );
  NAND U10517 ( .A(o[253]), .B(n5919), .Z(n6682) );
  NANDN U10518 ( .A(n5920), .B(creg[253]), .Z(n6681) );
  NAND U10519 ( .A(n6683), .B(n4545), .Z(n3348) );
  NANDN U10520 ( .A(init), .B(m[254]), .Z(n4545) );
  AND U10521 ( .A(n6684), .B(n6685), .Z(n6683) );
  NAND U10522 ( .A(n5919), .B(o[254]), .Z(n6685) );
  AND U10523 ( .A(n5920), .B(start_in[1023]), .Z(n5919) );
  NANDN U10524 ( .A(n5920), .B(creg[254]), .Z(n6684) );
  NANDN U10525 ( .A(n4377), .B(n6686), .Z(n5920) );
  NAND U10526 ( .A(n6687), .B(first_one), .Z(n6686) );
  ANDN U10527 ( .B(n6688), .A(n5914), .Z(n6687) );
  NANDN U10528 ( .A(n6689), .B(mul_pow), .Z(n6688) );
  NANDN U10529 ( .A(first_one), .B(n6690), .Z(n3347) );
  NANDN U10530 ( .A(n5914), .B(n6691), .Z(n6690) );
  ANDN U10531 ( .B(mul_pow), .A(n6692), .Z(n6691) );
  IV U10532 ( .A(start_in[1023]), .Z(n5914) );
  ANDN U10533 ( .B(start_reg[1023]), .A(n4377), .Z(start_in[1023]) );
  IV U10534 ( .A(init), .Z(n4377) );
  NAND U10535 ( .A(n6693), .B(n6694), .Z(c[9]) );
  NANDN U10536 ( .A(n6689), .B(creg[9]), .Z(n6694) );
  NANDN U10537 ( .A(n6695), .B(o[9]), .Z(n6693) );
  NAND U10538 ( .A(n6696), .B(n6697), .Z(c[99]) );
  NANDN U10539 ( .A(n6689), .B(creg[99]), .Z(n6697) );
  NANDN U10540 ( .A(n6695), .B(o[99]), .Z(n6696) );
  NAND U10541 ( .A(n6698), .B(n6699), .Z(c[98]) );
  NANDN U10542 ( .A(n6689), .B(creg[98]), .Z(n6699) );
  NANDN U10543 ( .A(n6695), .B(o[98]), .Z(n6698) );
  NAND U10544 ( .A(n6700), .B(n6701), .Z(c[97]) );
  NANDN U10545 ( .A(n6689), .B(creg[97]), .Z(n6701) );
  NANDN U10546 ( .A(n6695), .B(o[97]), .Z(n6700) );
  NAND U10547 ( .A(n6702), .B(n6703), .Z(c[96]) );
  NANDN U10548 ( .A(n6689), .B(creg[96]), .Z(n6703) );
  NANDN U10549 ( .A(n6695), .B(o[96]), .Z(n6702) );
  NAND U10550 ( .A(n6704), .B(n6705), .Z(c[95]) );
  NANDN U10551 ( .A(n6689), .B(creg[95]), .Z(n6705) );
  NANDN U10552 ( .A(n6695), .B(o[95]), .Z(n6704) );
  NAND U10553 ( .A(n6706), .B(n6707), .Z(c[94]) );
  NANDN U10554 ( .A(n6689), .B(creg[94]), .Z(n6707) );
  NANDN U10555 ( .A(n6695), .B(o[94]), .Z(n6706) );
  NAND U10556 ( .A(n6708), .B(n6709), .Z(c[93]) );
  NANDN U10557 ( .A(n6689), .B(creg[93]), .Z(n6709) );
  NANDN U10558 ( .A(n6695), .B(o[93]), .Z(n6708) );
  NAND U10559 ( .A(n6710), .B(n6711), .Z(c[92]) );
  NANDN U10560 ( .A(n6689), .B(creg[92]), .Z(n6711) );
  NANDN U10561 ( .A(n6695), .B(o[92]), .Z(n6710) );
  NAND U10562 ( .A(n6712), .B(n6713), .Z(c[91]) );
  NANDN U10563 ( .A(n6689), .B(creg[91]), .Z(n6713) );
  NANDN U10564 ( .A(n6695), .B(o[91]), .Z(n6712) );
  NAND U10565 ( .A(n6714), .B(n6715), .Z(c[90]) );
  NANDN U10566 ( .A(n6689), .B(creg[90]), .Z(n6715) );
  NANDN U10567 ( .A(n6695), .B(o[90]), .Z(n6714) );
  NAND U10568 ( .A(n6716), .B(n6717), .Z(c[8]) );
  NANDN U10569 ( .A(n6689), .B(creg[8]), .Z(n6717) );
  NANDN U10570 ( .A(n6695), .B(o[8]), .Z(n6716) );
  NAND U10571 ( .A(n6718), .B(n6719), .Z(c[89]) );
  NANDN U10572 ( .A(n6689), .B(creg[89]), .Z(n6719) );
  NANDN U10573 ( .A(n6695), .B(o[89]), .Z(n6718) );
  NAND U10574 ( .A(n6720), .B(n6721), .Z(c[88]) );
  NANDN U10575 ( .A(n6689), .B(creg[88]), .Z(n6721) );
  NANDN U10576 ( .A(n6695), .B(o[88]), .Z(n6720) );
  NAND U10577 ( .A(n6722), .B(n6723), .Z(c[87]) );
  NANDN U10578 ( .A(n6689), .B(creg[87]), .Z(n6723) );
  NANDN U10579 ( .A(n6695), .B(o[87]), .Z(n6722) );
  NAND U10580 ( .A(n6724), .B(n6725), .Z(c[86]) );
  NANDN U10581 ( .A(n6689), .B(creg[86]), .Z(n6725) );
  NANDN U10582 ( .A(n6695), .B(o[86]), .Z(n6724) );
  NAND U10583 ( .A(n6726), .B(n6727), .Z(c[85]) );
  NANDN U10584 ( .A(n6689), .B(creg[85]), .Z(n6727) );
  NANDN U10585 ( .A(n6695), .B(o[85]), .Z(n6726) );
  NAND U10586 ( .A(n6728), .B(n6729), .Z(c[84]) );
  NANDN U10587 ( .A(n6689), .B(creg[84]), .Z(n6729) );
  NANDN U10588 ( .A(n6695), .B(o[84]), .Z(n6728) );
  NAND U10589 ( .A(n6730), .B(n6731), .Z(c[83]) );
  NANDN U10590 ( .A(n6689), .B(creg[83]), .Z(n6731) );
  NANDN U10591 ( .A(n6695), .B(o[83]), .Z(n6730) );
  NAND U10592 ( .A(n6732), .B(n6733), .Z(c[82]) );
  NANDN U10593 ( .A(n6689), .B(creg[82]), .Z(n6733) );
  NANDN U10594 ( .A(n6695), .B(o[82]), .Z(n6732) );
  NAND U10595 ( .A(n6734), .B(n6735), .Z(c[81]) );
  NANDN U10596 ( .A(n6689), .B(creg[81]), .Z(n6735) );
  NANDN U10597 ( .A(n6695), .B(o[81]), .Z(n6734) );
  NAND U10598 ( .A(n6736), .B(n6737), .Z(c[80]) );
  NANDN U10599 ( .A(n6689), .B(creg[80]), .Z(n6737) );
  NANDN U10600 ( .A(n6695), .B(o[80]), .Z(n6736) );
  NAND U10601 ( .A(n6738), .B(n6739), .Z(c[7]) );
  NANDN U10602 ( .A(n6689), .B(creg[7]), .Z(n6739) );
  NANDN U10603 ( .A(n6695), .B(o[7]), .Z(n6738) );
  NAND U10604 ( .A(n6740), .B(n6741), .Z(c[79]) );
  NANDN U10605 ( .A(n6689), .B(creg[79]), .Z(n6741) );
  NANDN U10606 ( .A(n6695), .B(o[79]), .Z(n6740) );
  NAND U10607 ( .A(n6742), .B(n6743), .Z(c[78]) );
  NANDN U10608 ( .A(n6689), .B(creg[78]), .Z(n6743) );
  NANDN U10609 ( .A(n6695), .B(o[78]), .Z(n6742) );
  NAND U10610 ( .A(n6744), .B(n6745), .Z(c[77]) );
  NANDN U10611 ( .A(n6689), .B(creg[77]), .Z(n6745) );
  NANDN U10612 ( .A(n6695), .B(o[77]), .Z(n6744) );
  NAND U10613 ( .A(n6746), .B(n6747), .Z(c[76]) );
  NANDN U10614 ( .A(n6689), .B(creg[76]), .Z(n6747) );
  NANDN U10615 ( .A(n6695), .B(o[76]), .Z(n6746) );
  NAND U10616 ( .A(n6748), .B(n6749), .Z(c[75]) );
  NANDN U10617 ( .A(n6689), .B(creg[75]), .Z(n6749) );
  NANDN U10618 ( .A(n6695), .B(o[75]), .Z(n6748) );
  NAND U10619 ( .A(n6750), .B(n6751), .Z(c[74]) );
  NANDN U10620 ( .A(n6689), .B(creg[74]), .Z(n6751) );
  NANDN U10621 ( .A(n6695), .B(o[74]), .Z(n6750) );
  NAND U10622 ( .A(n6752), .B(n6753), .Z(c[73]) );
  NANDN U10623 ( .A(n6689), .B(creg[73]), .Z(n6753) );
  NANDN U10624 ( .A(n6695), .B(o[73]), .Z(n6752) );
  NAND U10625 ( .A(n6754), .B(n6755), .Z(c[72]) );
  NANDN U10626 ( .A(n6689), .B(creg[72]), .Z(n6755) );
  NANDN U10627 ( .A(n6695), .B(o[72]), .Z(n6754) );
  NAND U10628 ( .A(n6756), .B(n6757), .Z(c[71]) );
  NANDN U10629 ( .A(n6689), .B(creg[71]), .Z(n6757) );
  NANDN U10630 ( .A(n6695), .B(o[71]), .Z(n6756) );
  NAND U10631 ( .A(n6758), .B(n6759), .Z(c[70]) );
  NANDN U10632 ( .A(n6689), .B(creg[70]), .Z(n6759) );
  NANDN U10633 ( .A(n6695), .B(o[70]), .Z(n6758) );
  NAND U10634 ( .A(n6760), .B(n6761), .Z(c[6]) );
  NANDN U10635 ( .A(n6689), .B(creg[6]), .Z(n6761) );
  NANDN U10636 ( .A(n6695), .B(o[6]), .Z(n6760) );
  NAND U10637 ( .A(n6762), .B(n6763), .Z(c[69]) );
  NANDN U10638 ( .A(n6689), .B(creg[69]), .Z(n6763) );
  NANDN U10639 ( .A(n6695), .B(o[69]), .Z(n6762) );
  NAND U10640 ( .A(n6764), .B(n6765), .Z(c[68]) );
  NANDN U10641 ( .A(n6689), .B(creg[68]), .Z(n6765) );
  NANDN U10642 ( .A(n6695), .B(o[68]), .Z(n6764) );
  NAND U10643 ( .A(n6766), .B(n6767), .Z(c[67]) );
  NANDN U10644 ( .A(n6689), .B(creg[67]), .Z(n6767) );
  NANDN U10645 ( .A(n6695), .B(o[67]), .Z(n6766) );
  NAND U10646 ( .A(n6768), .B(n6769), .Z(c[66]) );
  NANDN U10647 ( .A(n6689), .B(creg[66]), .Z(n6769) );
  NANDN U10648 ( .A(n6695), .B(o[66]), .Z(n6768) );
  NAND U10649 ( .A(n6770), .B(n6771), .Z(c[65]) );
  NANDN U10650 ( .A(n6689), .B(creg[65]), .Z(n6771) );
  NANDN U10651 ( .A(n6695), .B(o[65]), .Z(n6770) );
  NAND U10652 ( .A(n6772), .B(n6773), .Z(c[64]) );
  NANDN U10653 ( .A(n6689), .B(creg[64]), .Z(n6773) );
  NANDN U10654 ( .A(n6695), .B(o[64]), .Z(n6772) );
  NAND U10655 ( .A(n6774), .B(n6775), .Z(c[63]) );
  NANDN U10656 ( .A(n6689), .B(creg[63]), .Z(n6775) );
  NANDN U10657 ( .A(n6695), .B(o[63]), .Z(n6774) );
  NAND U10658 ( .A(n6776), .B(n6777), .Z(c[62]) );
  NANDN U10659 ( .A(n6689), .B(creg[62]), .Z(n6777) );
  NANDN U10660 ( .A(n6695), .B(o[62]), .Z(n6776) );
  NAND U10661 ( .A(n6778), .B(n6779), .Z(c[61]) );
  NANDN U10662 ( .A(n6689), .B(creg[61]), .Z(n6779) );
  NANDN U10663 ( .A(n6695), .B(o[61]), .Z(n6778) );
  NAND U10664 ( .A(n6780), .B(n6781), .Z(c[60]) );
  NANDN U10665 ( .A(n6689), .B(creg[60]), .Z(n6781) );
  NANDN U10666 ( .A(n6695), .B(o[60]), .Z(n6780) );
  NAND U10667 ( .A(n6782), .B(n6783), .Z(c[5]) );
  NANDN U10668 ( .A(n6689), .B(creg[5]), .Z(n6783) );
  NANDN U10669 ( .A(n6695), .B(o[5]), .Z(n6782) );
  NAND U10670 ( .A(n6784), .B(n6785), .Z(c[59]) );
  NANDN U10671 ( .A(n6689), .B(creg[59]), .Z(n6785) );
  NANDN U10672 ( .A(n6695), .B(o[59]), .Z(n6784) );
  NAND U10673 ( .A(n6786), .B(n6787), .Z(c[58]) );
  NANDN U10674 ( .A(n6689), .B(creg[58]), .Z(n6787) );
  NANDN U10675 ( .A(n6695), .B(o[58]), .Z(n6786) );
  NAND U10676 ( .A(n6788), .B(n6789), .Z(c[57]) );
  NANDN U10677 ( .A(n6689), .B(creg[57]), .Z(n6789) );
  NANDN U10678 ( .A(n6695), .B(o[57]), .Z(n6788) );
  NAND U10679 ( .A(n6790), .B(n6791), .Z(c[56]) );
  NANDN U10680 ( .A(n6689), .B(creg[56]), .Z(n6791) );
  NANDN U10681 ( .A(n6695), .B(o[56]), .Z(n6790) );
  NAND U10682 ( .A(n6792), .B(n6793), .Z(c[55]) );
  NANDN U10683 ( .A(n6689), .B(creg[55]), .Z(n6793) );
  NANDN U10684 ( .A(n6695), .B(o[55]), .Z(n6792) );
  NAND U10685 ( .A(n6794), .B(n6795), .Z(c[54]) );
  NANDN U10686 ( .A(n6689), .B(creg[54]), .Z(n6795) );
  NANDN U10687 ( .A(n6695), .B(o[54]), .Z(n6794) );
  NAND U10688 ( .A(n6796), .B(n6797), .Z(c[53]) );
  NANDN U10689 ( .A(n6689), .B(creg[53]), .Z(n6797) );
  NANDN U10690 ( .A(n6695), .B(o[53]), .Z(n6796) );
  NAND U10691 ( .A(n6798), .B(n6799), .Z(c[52]) );
  NANDN U10692 ( .A(n6689), .B(creg[52]), .Z(n6799) );
  NANDN U10693 ( .A(n6695), .B(o[52]), .Z(n6798) );
  NAND U10694 ( .A(n6800), .B(n6801), .Z(c[51]) );
  NANDN U10695 ( .A(n6689), .B(creg[51]), .Z(n6801) );
  NANDN U10696 ( .A(n6695), .B(o[51]), .Z(n6800) );
  NAND U10697 ( .A(n6802), .B(n6803), .Z(c[50]) );
  NANDN U10698 ( .A(n6689), .B(creg[50]), .Z(n6803) );
  NANDN U10699 ( .A(n6695), .B(o[50]), .Z(n6802) );
  NAND U10700 ( .A(n6804), .B(n6805), .Z(c[4]) );
  NANDN U10701 ( .A(n6689), .B(creg[4]), .Z(n6805) );
  NANDN U10702 ( .A(n6695), .B(o[4]), .Z(n6804) );
  NAND U10703 ( .A(n6806), .B(n6807), .Z(c[49]) );
  NANDN U10704 ( .A(n6689), .B(creg[49]), .Z(n6807) );
  NANDN U10705 ( .A(n6695), .B(o[49]), .Z(n6806) );
  NAND U10706 ( .A(n6808), .B(n6809), .Z(c[48]) );
  NANDN U10707 ( .A(n6689), .B(creg[48]), .Z(n6809) );
  NANDN U10708 ( .A(n6695), .B(o[48]), .Z(n6808) );
  NAND U10709 ( .A(n6810), .B(n6811), .Z(c[47]) );
  NANDN U10710 ( .A(n6689), .B(creg[47]), .Z(n6811) );
  NANDN U10711 ( .A(n6695), .B(o[47]), .Z(n6810) );
  NAND U10712 ( .A(n6812), .B(n6813), .Z(c[46]) );
  NANDN U10713 ( .A(n6689), .B(creg[46]), .Z(n6813) );
  NANDN U10714 ( .A(n6695), .B(o[46]), .Z(n6812) );
  NAND U10715 ( .A(n6814), .B(n6815), .Z(c[45]) );
  NANDN U10716 ( .A(n6689), .B(creg[45]), .Z(n6815) );
  NANDN U10717 ( .A(n6695), .B(o[45]), .Z(n6814) );
  NAND U10718 ( .A(n6816), .B(n6817), .Z(c[44]) );
  NANDN U10719 ( .A(n6689), .B(creg[44]), .Z(n6817) );
  NANDN U10720 ( .A(n6695), .B(o[44]), .Z(n6816) );
  NAND U10721 ( .A(n6818), .B(n6819), .Z(c[43]) );
  NANDN U10722 ( .A(n6689), .B(creg[43]), .Z(n6819) );
  NANDN U10723 ( .A(n6695), .B(o[43]), .Z(n6818) );
  NAND U10724 ( .A(n6820), .B(n6821), .Z(c[42]) );
  NANDN U10725 ( .A(n6689), .B(creg[42]), .Z(n6821) );
  NANDN U10726 ( .A(n6695), .B(o[42]), .Z(n6820) );
  NAND U10727 ( .A(n6822), .B(n6823), .Z(c[41]) );
  NANDN U10728 ( .A(n6689), .B(creg[41]), .Z(n6823) );
  NANDN U10729 ( .A(n6695), .B(o[41]), .Z(n6822) );
  NAND U10730 ( .A(n6824), .B(n6825), .Z(c[40]) );
  NANDN U10731 ( .A(n6689), .B(creg[40]), .Z(n6825) );
  NANDN U10732 ( .A(n6695), .B(o[40]), .Z(n6824) );
  NAND U10733 ( .A(n6826), .B(n6827), .Z(c[3]) );
  NANDN U10734 ( .A(n6689), .B(creg[3]), .Z(n6827) );
  NANDN U10735 ( .A(n6695), .B(o[3]), .Z(n6826) );
  NAND U10736 ( .A(n6828), .B(n6829), .Z(c[39]) );
  NANDN U10737 ( .A(n6689), .B(creg[39]), .Z(n6829) );
  NANDN U10738 ( .A(n6695), .B(o[39]), .Z(n6828) );
  NAND U10739 ( .A(n6830), .B(n6831), .Z(c[38]) );
  NANDN U10740 ( .A(n6689), .B(creg[38]), .Z(n6831) );
  NANDN U10741 ( .A(n6695), .B(o[38]), .Z(n6830) );
  NAND U10742 ( .A(n6832), .B(n6833), .Z(c[37]) );
  NANDN U10743 ( .A(n6689), .B(creg[37]), .Z(n6833) );
  NANDN U10744 ( .A(n6695), .B(o[37]), .Z(n6832) );
  NAND U10745 ( .A(n6834), .B(n6835), .Z(c[36]) );
  NANDN U10746 ( .A(n6689), .B(creg[36]), .Z(n6835) );
  NANDN U10747 ( .A(n6695), .B(o[36]), .Z(n6834) );
  NAND U10748 ( .A(n6836), .B(n6837), .Z(c[35]) );
  NANDN U10749 ( .A(n6689), .B(creg[35]), .Z(n6837) );
  NANDN U10750 ( .A(n6695), .B(o[35]), .Z(n6836) );
  NAND U10751 ( .A(n6838), .B(n6839), .Z(c[34]) );
  NANDN U10752 ( .A(n6689), .B(creg[34]), .Z(n6839) );
  NANDN U10753 ( .A(n6695), .B(o[34]), .Z(n6838) );
  NAND U10754 ( .A(n6840), .B(n6841), .Z(c[33]) );
  NANDN U10755 ( .A(n6689), .B(creg[33]), .Z(n6841) );
  NANDN U10756 ( .A(n6695), .B(o[33]), .Z(n6840) );
  NAND U10757 ( .A(n6842), .B(n6843), .Z(c[32]) );
  NANDN U10758 ( .A(n6689), .B(creg[32]), .Z(n6843) );
  NANDN U10759 ( .A(n6695), .B(o[32]), .Z(n6842) );
  NAND U10760 ( .A(n6844), .B(n6845), .Z(c[31]) );
  NANDN U10761 ( .A(n6689), .B(creg[31]), .Z(n6845) );
  NANDN U10762 ( .A(n6695), .B(o[31]), .Z(n6844) );
  NAND U10763 ( .A(n6846), .B(n6847), .Z(c[30]) );
  NANDN U10764 ( .A(n6689), .B(creg[30]), .Z(n6847) );
  NANDN U10765 ( .A(n6695), .B(o[30]), .Z(n6846) );
  NAND U10766 ( .A(n6848), .B(n6849), .Z(c[2]) );
  NANDN U10767 ( .A(n6689), .B(creg[2]), .Z(n6849) );
  NANDN U10768 ( .A(n6695), .B(o[2]), .Z(n6848) );
  NAND U10769 ( .A(n6850), .B(n6851), .Z(c[29]) );
  NANDN U10770 ( .A(n6689), .B(creg[29]), .Z(n6851) );
  NANDN U10771 ( .A(n6695), .B(o[29]), .Z(n6850) );
  NAND U10772 ( .A(n6852), .B(n6853), .Z(c[28]) );
  NANDN U10773 ( .A(n6689), .B(creg[28]), .Z(n6853) );
  NANDN U10774 ( .A(n6695), .B(o[28]), .Z(n6852) );
  NAND U10775 ( .A(n6854), .B(n6855), .Z(c[27]) );
  NANDN U10776 ( .A(n6689), .B(creg[27]), .Z(n6855) );
  NANDN U10777 ( .A(n6695), .B(o[27]), .Z(n6854) );
  NAND U10778 ( .A(n6856), .B(n6857), .Z(c[26]) );
  NANDN U10779 ( .A(n6689), .B(creg[26]), .Z(n6857) );
  NANDN U10780 ( .A(n6695), .B(o[26]), .Z(n6856) );
  NAND U10781 ( .A(n6858), .B(n6859), .Z(c[25]) );
  NANDN U10782 ( .A(n6689), .B(creg[25]), .Z(n6859) );
  NANDN U10783 ( .A(n6695), .B(o[25]), .Z(n6858) );
  NAND U10784 ( .A(n6860), .B(n6861), .Z(c[255]) );
  NANDN U10785 ( .A(n6689), .B(creg[255]), .Z(n6861) );
  NANDN U10786 ( .A(n6695), .B(o[255]), .Z(n6860) );
  NAND U10787 ( .A(n6862), .B(n6863), .Z(c[254]) );
  NANDN U10788 ( .A(n6689), .B(creg[254]), .Z(n6863) );
  NANDN U10789 ( .A(n6695), .B(o[254]), .Z(n6862) );
  NAND U10790 ( .A(n6864), .B(n6865), .Z(c[253]) );
  NANDN U10791 ( .A(n6689), .B(creg[253]), .Z(n6865) );
  NANDN U10792 ( .A(n6695), .B(o[253]), .Z(n6864) );
  NAND U10793 ( .A(n6866), .B(n6867), .Z(c[252]) );
  NANDN U10794 ( .A(n6689), .B(creg[252]), .Z(n6867) );
  NANDN U10795 ( .A(n6695), .B(o[252]), .Z(n6866) );
  NAND U10796 ( .A(n6868), .B(n6869), .Z(c[251]) );
  NANDN U10797 ( .A(n6689), .B(creg[251]), .Z(n6869) );
  NANDN U10798 ( .A(n6695), .B(o[251]), .Z(n6868) );
  NAND U10799 ( .A(n6870), .B(n6871), .Z(c[250]) );
  NANDN U10800 ( .A(n6689), .B(creg[250]), .Z(n6871) );
  NANDN U10801 ( .A(n6695), .B(o[250]), .Z(n6870) );
  NAND U10802 ( .A(n6872), .B(n6873), .Z(c[24]) );
  NANDN U10803 ( .A(n6689), .B(creg[24]), .Z(n6873) );
  NANDN U10804 ( .A(n6695), .B(o[24]), .Z(n6872) );
  NAND U10805 ( .A(n6874), .B(n6875), .Z(c[249]) );
  NANDN U10806 ( .A(n6689), .B(creg[249]), .Z(n6875) );
  NANDN U10807 ( .A(n6695), .B(o[249]), .Z(n6874) );
  NAND U10808 ( .A(n6876), .B(n6877), .Z(c[248]) );
  NANDN U10809 ( .A(n6689), .B(creg[248]), .Z(n6877) );
  NANDN U10810 ( .A(n6695), .B(o[248]), .Z(n6876) );
  NAND U10811 ( .A(n6878), .B(n6879), .Z(c[247]) );
  NANDN U10812 ( .A(n6689), .B(creg[247]), .Z(n6879) );
  NANDN U10813 ( .A(n6695), .B(o[247]), .Z(n6878) );
  NAND U10814 ( .A(n6880), .B(n6881), .Z(c[246]) );
  NANDN U10815 ( .A(n6689), .B(creg[246]), .Z(n6881) );
  NANDN U10816 ( .A(n6695), .B(o[246]), .Z(n6880) );
  NAND U10817 ( .A(n6882), .B(n6883), .Z(c[245]) );
  NANDN U10818 ( .A(n6689), .B(creg[245]), .Z(n6883) );
  NANDN U10819 ( .A(n6695), .B(o[245]), .Z(n6882) );
  NAND U10820 ( .A(n6884), .B(n6885), .Z(c[244]) );
  NANDN U10821 ( .A(n6689), .B(creg[244]), .Z(n6885) );
  NANDN U10822 ( .A(n6695), .B(o[244]), .Z(n6884) );
  NAND U10823 ( .A(n6886), .B(n6887), .Z(c[243]) );
  NANDN U10824 ( .A(n6689), .B(creg[243]), .Z(n6887) );
  NANDN U10825 ( .A(n6695), .B(o[243]), .Z(n6886) );
  NAND U10826 ( .A(n6888), .B(n6889), .Z(c[242]) );
  NANDN U10827 ( .A(n6689), .B(creg[242]), .Z(n6889) );
  NANDN U10828 ( .A(n6695), .B(o[242]), .Z(n6888) );
  NAND U10829 ( .A(n6890), .B(n6891), .Z(c[241]) );
  NANDN U10830 ( .A(n6689), .B(creg[241]), .Z(n6891) );
  NANDN U10831 ( .A(n6695), .B(o[241]), .Z(n6890) );
  NAND U10832 ( .A(n6892), .B(n6893), .Z(c[240]) );
  NANDN U10833 ( .A(n6689), .B(creg[240]), .Z(n6893) );
  NANDN U10834 ( .A(n6695), .B(o[240]), .Z(n6892) );
  NAND U10835 ( .A(n6894), .B(n6895), .Z(c[23]) );
  NANDN U10836 ( .A(n6689), .B(creg[23]), .Z(n6895) );
  NANDN U10837 ( .A(n6695), .B(o[23]), .Z(n6894) );
  NAND U10838 ( .A(n6896), .B(n6897), .Z(c[239]) );
  NANDN U10839 ( .A(n6689), .B(creg[239]), .Z(n6897) );
  NANDN U10840 ( .A(n6695), .B(o[239]), .Z(n6896) );
  NAND U10841 ( .A(n6898), .B(n6899), .Z(c[238]) );
  NANDN U10842 ( .A(n6689), .B(creg[238]), .Z(n6899) );
  NANDN U10843 ( .A(n6695), .B(o[238]), .Z(n6898) );
  NAND U10844 ( .A(n6900), .B(n6901), .Z(c[237]) );
  NANDN U10845 ( .A(n6689), .B(creg[237]), .Z(n6901) );
  NANDN U10846 ( .A(n6695), .B(o[237]), .Z(n6900) );
  NAND U10847 ( .A(n6902), .B(n6903), .Z(c[236]) );
  NANDN U10848 ( .A(n6689), .B(creg[236]), .Z(n6903) );
  NANDN U10849 ( .A(n6695), .B(o[236]), .Z(n6902) );
  NAND U10850 ( .A(n6904), .B(n6905), .Z(c[235]) );
  NANDN U10851 ( .A(n6689), .B(creg[235]), .Z(n6905) );
  NANDN U10852 ( .A(n6695), .B(o[235]), .Z(n6904) );
  NAND U10853 ( .A(n6906), .B(n6907), .Z(c[234]) );
  NANDN U10854 ( .A(n6689), .B(creg[234]), .Z(n6907) );
  NANDN U10855 ( .A(n6695), .B(o[234]), .Z(n6906) );
  NAND U10856 ( .A(n6908), .B(n6909), .Z(c[233]) );
  NANDN U10857 ( .A(n6689), .B(creg[233]), .Z(n6909) );
  NANDN U10858 ( .A(n6695), .B(o[233]), .Z(n6908) );
  NAND U10859 ( .A(n6910), .B(n6911), .Z(c[232]) );
  NANDN U10860 ( .A(n6689), .B(creg[232]), .Z(n6911) );
  NANDN U10861 ( .A(n6695), .B(o[232]), .Z(n6910) );
  NAND U10862 ( .A(n6912), .B(n6913), .Z(c[231]) );
  NANDN U10863 ( .A(n6689), .B(creg[231]), .Z(n6913) );
  NANDN U10864 ( .A(n6695), .B(o[231]), .Z(n6912) );
  NAND U10865 ( .A(n6914), .B(n6915), .Z(c[230]) );
  NANDN U10866 ( .A(n6689), .B(creg[230]), .Z(n6915) );
  NANDN U10867 ( .A(n6695), .B(o[230]), .Z(n6914) );
  NAND U10868 ( .A(n6916), .B(n6917), .Z(c[22]) );
  NANDN U10869 ( .A(n6689), .B(creg[22]), .Z(n6917) );
  NANDN U10870 ( .A(n6695), .B(o[22]), .Z(n6916) );
  NAND U10871 ( .A(n6918), .B(n6919), .Z(c[229]) );
  NANDN U10872 ( .A(n6689), .B(creg[229]), .Z(n6919) );
  NANDN U10873 ( .A(n6695), .B(o[229]), .Z(n6918) );
  NAND U10874 ( .A(n6920), .B(n6921), .Z(c[228]) );
  NANDN U10875 ( .A(n6689), .B(creg[228]), .Z(n6921) );
  NANDN U10876 ( .A(n6695), .B(o[228]), .Z(n6920) );
  NAND U10877 ( .A(n6922), .B(n6923), .Z(c[227]) );
  NANDN U10878 ( .A(n6689), .B(creg[227]), .Z(n6923) );
  NANDN U10879 ( .A(n6695), .B(o[227]), .Z(n6922) );
  NAND U10880 ( .A(n6924), .B(n6925), .Z(c[226]) );
  NANDN U10881 ( .A(n6689), .B(creg[226]), .Z(n6925) );
  NANDN U10882 ( .A(n6695), .B(o[226]), .Z(n6924) );
  NAND U10883 ( .A(n6926), .B(n6927), .Z(c[225]) );
  NANDN U10884 ( .A(n6689), .B(creg[225]), .Z(n6927) );
  NANDN U10885 ( .A(n6695), .B(o[225]), .Z(n6926) );
  NAND U10886 ( .A(n6928), .B(n6929), .Z(c[224]) );
  NANDN U10887 ( .A(n6689), .B(creg[224]), .Z(n6929) );
  NANDN U10888 ( .A(n6695), .B(o[224]), .Z(n6928) );
  NAND U10889 ( .A(n6930), .B(n6931), .Z(c[223]) );
  NANDN U10890 ( .A(n6689), .B(creg[223]), .Z(n6931) );
  NANDN U10891 ( .A(n6695), .B(o[223]), .Z(n6930) );
  NAND U10892 ( .A(n6932), .B(n6933), .Z(c[222]) );
  NANDN U10893 ( .A(n6689), .B(creg[222]), .Z(n6933) );
  NANDN U10894 ( .A(n6695), .B(o[222]), .Z(n6932) );
  NAND U10895 ( .A(n6934), .B(n6935), .Z(c[221]) );
  NANDN U10896 ( .A(n6689), .B(creg[221]), .Z(n6935) );
  NANDN U10897 ( .A(n6695), .B(o[221]), .Z(n6934) );
  NAND U10898 ( .A(n6936), .B(n6937), .Z(c[220]) );
  NANDN U10899 ( .A(n6689), .B(creg[220]), .Z(n6937) );
  NANDN U10900 ( .A(n6695), .B(o[220]), .Z(n6936) );
  NAND U10901 ( .A(n6938), .B(n6939), .Z(c[21]) );
  NANDN U10902 ( .A(n6689), .B(creg[21]), .Z(n6939) );
  NANDN U10903 ( .A(n6695), .B(o[21]), .Z(n6938) );
  NAND U10904 ( .A(n6940), .B(n6941), .Z(c[219]) );
  NANDN U10905 ( .A(n6689), .B(creg[219]), .Z(n6941) );
  NANDN U10906 ( .A(n6695), .B(o[219]), .Z(n6940) );
  NAND U10907 ( .A(n6942), .B(n6943), .Z(c[218]) );
  NANDN U10908 ( .A(n6689), .B(creg[218]), .Z(n6943) );
  NANDN U10909 ( .A(n6695), .B(o[218]), .Z(n6942) );
  NAND U10910 ( .A(n6944), .B(n6945), .Z(c[217]) );
  NANDN U10911 ( .A(n6689), .B(creg[217]), .Z(n6945) );
  NANDN U10912 ( .A(n6695), .B(o[217]), .Z(n6944) );
  NAND U10913 ( .A(n6946), .B(n6947), .Z(c[216]) );
  NANDN U10914 ( .A(n6689), .B(creg[216]), .Z(n6947) );
  NANDN U10915 ( .A(n6695), .B(o[216]), .Z(n6946) );
  NAND U10916 ( .A(n6948), .B(n6949), .Z(c[215]) );
  NANDN U10917 ( .A(n6689), .B(creg[215]), .Z(n6949) );
  NANDN U10918 ( .A(n6695), .B(o[215]), .Z(n6948) );
  NAND U10919 ( .A(n6950), .B(n6951), .Z(c[214]) );
  NANDN U10920 ( .A(n6689), .B(creg[214]), .Z(n6951) );
  NANDN U10921 ( .A(n6695), .B(o[214]), .Z(n6950) );
  NAND U10922 ( .A(n6952), .B(n6953), .Z(c[213]) );
  NANDN U10923 ( .A(n6689), .B(creg[213]), .Z(n6953) );
  NANDN U10924 ( .A(n6695), .B(o[213]), .Z(n6952) );
  NAND U10925 ( .A(n6954), .B(n6955), .Z(c[212]) );
  NANDN U10926 ( .A(n6689), .B(creg[212]), .Z(n6955) );
  NANDN U10927 ( .A(n6695), .B(o[212]), .Z(n6954) );
  NAND U10928 ( .A(n6956), .B(n6957), .Z(c[211]) );
  NANDN U10929 ( .A(n6689), .B(creg[211]), .Z(n6957) );
  NANDN U10930 ( .A(n6695), .B(o[211]), .Z(n6956) );
  NAND U10931 ( .A(n6958), .B(n6959), .Z(c[210]) );
  NANDN U10932 ( .A(n6689), .B(creg[210]), .Z(n6959) );
  NANDN U10933 ( .A(n6695), .B(o[210]), .Z(n6958) );
  NAND U10934 ( .A(n6960), .B(n6961), .Z(c[20]) );
  NANDN U10935 ( .A(n6689), .B(creg[20]), .Z(n6961) );
  NANDN U10936 ( .A(n6695), .B(o[20]), .Z(n6960) );
  NAND U10937 ( .A(n6962), .B(n6963), .Z(c[209]) );
  NANDN U10938 ( .A(n6689), .B(creg[209]), .Z(n6963) );
  NANDN U10939 ( .A(n6695), .B(o[209]), .Z(n6962) );
  NAND U10940 ( .A(n6964), .B(n6965), .Z(c[208]) );
  NANDN U10941 ( .A(n6689), .B(creg[208]), .Z(n6965) );
  NANDN U10942 ( .A(n6695), .B(o[208]), .Z(n6964) );
  NAND U10943 ( .A(n6966), .B(n6967), .Z(c[207]) );
  NANDN U10944 ( .A(n6689), .B(creg[207]), .Z(n6967) );
  NANDN U10945 ( .A(n6695), .B(o[207]), .Z(n6966) );
  NAND U10946 ( .A(n6968), .B(n6969), .Z(c[206]) );
  NANDN U10947 ( .A(n6689), .B(creg[206]), .Z(n6969) );
  NANDN U10948 ( .A(n6695), .B(o[206]), .Z(n6968) );
  NAND U10949 ( .A(n6970), .B(n6971), .Z(c[205]) );
  NANDN U10950 ( .A(n6689), .B(creg[205]), .Z(n6971) );
  NANDN U10951 ( .A(n6695), .B(o[205]), .Z(n6970) );
  NAND U10952 ( .A(n6972), .B(n6973), .Z(c[204]) );
  NANDN U10953 ( .A(n6689), .B(creg[204]), .Z(n6973) );
  NANDN U10954 ( .A(n6695), .B(o[204]), .Z(n6972) );
  NAND U10955 ( .A(n6974), .B(n6975), .Z(c[203]) );
  NANDN U10956 ( .A(n6689), .B(creg[203]), .Z(n6975) );
  NANDN U10957 ( .A(n6695), .B(o[203]), .Z(n6974) );
  NAND U10958 ( .A(n6976), .B(n6977), .Z(c[202]) );
  NANDN U10959 ( .A(n6689), .B(creg[202]), .Z(n6977) );
  NANDN U10960 ( .A(n6695), .B(o[202]), .Z(n6976) );
  NAND U10961 ( .A(n6978), .B(n6979), .Z(c[201]) );
  NANDN U10962 ( .A(n6689), .B(creg[201]), .Z(n6979) );
  NANDN U10963 ( .A(n6695), .B(o[201]), .Z(n6978) );
  NAND U10964 ( .A(n6980), .B(n6981), .Z(c[200]) );
  NANDN U10965 ( .A(n6689), .B(creg[200]), .Z(n6981) );
  NANDN U10966 ( .A(n6695), .B(o[200]), .Z(n6980) );
  NAND U10967 ( .A(n6982), .B(n6983), .Z(c[1]) );
  NANDN U10968 ( .A(n6689), .B(creg[1]), .Z(n6983) );
  NANDN U10969 ( .A(n6695), .B(o[1]), .Z(n6982) );
  NAND U10970 ( .A(n6984), .B(n6985), .Z(c[19]) );
  NANDN U10971 ( .A(n6689), .B(creg[19]), .Z(n6985) );
  NANDN U10972 ( .A(n6695), .B(o[19]), .Z(n6984) );
  NAND U10973 ( .A(n6986), .B(n6987), .Z(c[199]) );
  NANDN U10974 ( .A(n6689), .B(creg[199]), .Z(n6987) );
  NANDN U10975 ( .A(n6695), .B(o[199]), .Z(n6986) );
  NAND U10976 ( .A(n6988), .B(n6989), .Z(c[198]) );
  NANDN U10977 ( .A(n6689), .B(creg[198]), .Z(n6989) );
  NANDN U10978 ( .A(n6695), .B(o[198]), .Z(n6988) );
  NAND U10979 ( .A(n6990), .B(n6991), .Z(c[197]) );
  NANDN U10980 ( .A(n6689), .B(creg[197]), .Z(n6991) );
  NANDN U10981 ( .A(n6695), .B(o[197]), .Z(n6990) );
  NAND U10982 ( .A(n6992), .B(n6993), .Z(c[196]) );
  NANDN U10983 ( .A(n6689), .B(creg[196]), .Z(n6993) );
  NANDN U10984 ( .A(n6695), .B(o[196]), .Z(n6992) );
  NAND U10985 ( .A(n6994), .B(n6995), .Z(c[195]) );
  NANDN U10986 ( .A(n6689), .B(creg[195]), .Z(n6995) );
  NANDN U10987 ( .A(n6695), .B(o[195]), .Z(n6994) );
  NAND U10988 ( .A(n6996), .B(n6997), .Z(c[194]) );
  NANDN U10989 ( .A(n6689), .B(creg[194]), .Z(n6997) );
  NANDN U10990 ( .A(n6695), .B(o[194]), .Z(n6996) );
  NAND U10991 ( .A(n6998), .B(n6999), .Z(c[193]) );
  NANDN U10992 ( .A(n6689), .B(creg[193]), .Z(n6999) );
  NANDN U10993 ( .A(n6695), .B(o[193]), .Z(n6998) );
  NAND U10994 ( .A(n7000), .B(n7001), .Z(c[192]) );
  NANDN U10995 ( .A(n6689), .B(creg[192]), .Z(n7001) );
  NANDN U10996 ( .A(n6695), .B(o[192]), .Z(n7000) );
  NAND U10997 ( .A(n7002), .B(n7003), .Z(c[191]) );
  NANDN U10998 ( .A(n6689), .B(creg[191]), .Z(n7003) );
  NANDN U10999 ( .A(n6695), .B(o[191]), .Z(n7002) );
  NAND U11000 ( .A(n7004), .B(n7005), .Z(c[190]) );
  NANDN U11001 ( .A(n6689), .B(creg[190]), .Z(n7005) );
  NANDN U11002 ( .A(n6695), .B(o[190]), .Z(n7004) );
  NAND U11003 ( .A(n7006), .B(n7007), .Z(c[18]) );
  NANDN U11004 ( .A(n6689), .B(creg[18]), .Z(n7007) );
  NANDN U11005 ( .A(n6695), .B(o[18]), .Z(n7006) );
  NAND U11006 ( .A(n7008), .B(n7009), .Z(c[189]) );
  NANDN U11007 ( .A(n6689), .B(creg[189]), .Z(n7009) );
  NANDN U11008 ( .A(n6695), .B(o[189]), .Z(n7008) );
  NAND U11009 ( .A(n7010), .B(n7011), .Z(c[188]) );
  NANDN U11010 ( .A(n6689), .B(creg[188]), .Z(n7011) );
  NANDN U11011 ( .A(n6695), .B(o[188]), .Z(n7010) );
  NAND U11012 ( .A(n7012), .B(n7013), .Z(c[187]) );
  NANDN U11013 ( .A(n6689), .B(creg[187]), .Z(n7013) );
  NANDN U11014 ( .A(n6695), .B(o[187]), .Z(n7012) );
  NAND U11015 ( .A(n7014), .B(n7015), .Z(c[186]) );
  NANDN U11016 ( .A(n6689), .B(creg[186]), .Z(n7015) );
  NANDN U11017 ( .A(n6695), .B(o[186]), .Z(n7014) );
  NAND U11018 ( .A(n7016), .B(n7017), .Z(c[185]) );
  NANDN U11019 ( .A(n6689), .B(creg[185]), .Z(n7017) );
  NANDN U11020 ( .A(n6695), .B(o[185]), .Z(n7016) );
  NAND U11021 ( .A(n7018), .B(n7019), .Z(c[184]) );
  NANDN U11022 ( .A(n6689), .B(creg[184]), .Z(n7019) );
  NANDN U11023 ( .A(n6695), .B(o[184]), .Z(n7018) );
  NAND U11024 ( .A(n7020), .B(n7021), .Z(c[183]) );
  NANDN U11025 ( .A(n6689), .B(creg[183]), .Z(n7021) );
  NANDN U11026 ( .A(n6695), .B(o[183]), .Z(n7020) );
  NAND U11027 ( .A(n7022), .B(n7023), .Z(c[182]) );
  NANDN U11028 ( .A(n6689), .B(creg[182]), .Z(n7023) );
  NANDN U11029 ( .A(n6695), .B(o[182]), .Z(n7022) );
  NAND U11030 ( .A(n7024), .B(n7025), .Z(c[181]) );
  NANDN U11031 ( .A(n6689), .B(creg[181]), .Z(n7025) );
  NANDN U11032 ( .A(n6695), .B(o[181]), .Z(n7024) );
  NAND U11033 ( .A(n7026), .B(n7027), .Z(c[180]) );
  NANDN U11034 ( .A(n6689), .B(creg[180]), .Z(n7027) );
  NANDN U11035 ( .A(n6695), .B(o[180]), .Z(n7026) );
  NAND U11036 ( .A(n7028), .B(n7029), .Z(c[17]) );
  NANDN U11037 ( .A(n6689), .B(creg[17]), .Z(n7029) );
  NANDN U11038 ( .A(n6695), .B(o[17]), .Z(n7028) );
  NAND U11039 ( .A(n7030), .B(n7031), .Z(c[179]) );
  NANDN U11040 ( .A(n6689), .B(creg[179]), .Z(n7031) );
  NANDN U11041 ( .A(n6695), .B(o[179]), .Z(n7030) );
  NAND U11042 ( .A(n7032), .B(n7033), .Z(c[178]) );
  NANDN U11043 ( .A(n6689), .B(creg[178]), .Z(n7033) );
  NANDN U11044 ( .A(n6695), .B(o[178]), .Z(n7032) );
  NAND U11045 ( .A(n7034), .B(n7035), .Z(c[177]) );
  NANDN U11046 ( .A(n6689), .B(creg[177]), .Z(n7035) );
  NANDN U11047 ( .A(n6695), .B(o[177]), .Z(n7034) );
  NAND U11048 ( .A(n7036), .B(n7037), .Z(c[176]) );
  NANDN U11049 ( .A(n6689), .B(creg[176]), .Z(n7037) );
  NANDN U11050 ( .A(n6695), .B(o[176]), .Z(n7036) );
  NAND U11051 ( .A(n7038), .B(n7039), .Z(c[175]) );
  NANDN U11052 ( .A(n6689), .B(creg[175]), .Z(n7039) );
  NANDN U11053 ( .A(n6695), .B(o[175]), .Z(n7038) );
  NAND U11054 ( .A(n7040), .B(n7041), .Z(c[174]) );
  NANDN U11055 ( .A(n6689), .B(creg[174]), .Z(n7041) );
  NANDN U11056 ( .A(n6695), .B(o[174]), .Z(n7040) );
  NAND U11057 ( .A(n7042), .B(n7043), .Z(c[173]) );
  NANDN U11058 ( .A(n6689), .B(creg[173]), .Z(n7043) );
  NANDN U11059 ( .A(n6695), .B(o[173]), .Z(n7042) );
  NAND U11060 ( .A(n7044), .B(n7045), .Z(c[172]) );
  NANDN U11061 ( .A(n6689), .B(creg[172]), .Z(n7045) );
  NANDN U11062 ( .A(n6695), .B(o[172]), .Z(n7044) );
  NAND U11063 ( .A(n7046), .B(n7047), .Z(c[171]) );
  NANDN U11064 ( .A(n6689), .B(creg[171]), .Z(n7047) );
  NANDN U11065 ( .A(n6695), .B(o[171]), .Z(n7046) );
  NAND U11066 ( .A(n7048), .B(n7049), .Z(c[170]) );
  NANDN U11067 ( .A(n6689), .B(creg[170]), .Z(n7049) );
  NANDN U11068 ( .A(n6695), .B(o[170]), .Z(n7048) );
  NAND U11069 ( .A(n7050), .B(n7051), .Z(c[16]) );
  NANDN U11070 ( .A(n6689), .B(creg[16]), .Z(n7051) );
  NANDN U11071 ( .A(n6695), .B(o[16]), .Z(n7050) );
  NAND U11072 ( .A(n7052), .B(n7053), .Z(c[169]) );
  NANDN U11073 ( .A(n6689), .B(creg[169]), .Z(n7053) );
  NANDN U11074 ( .A(n6695), .B(o[169]), .Z(n7052) );
  NAND U11075 ( .A(n7054), .B(n7055), .Z(c[168]) );
  NANDN U11076 ( .A(n6689), .B(creg[168]), .Z(n7055) );
  NANDN U11077 ( .A(n6695), .B(o[168]), .Z(n7054) );
  NAND U11078 ( .A(n7056), .B(n7057), .Z(c[167]) );
  NANDN U11079 ( .A(n6689), .B(creg[167]), .Z(n7057) );
  NANDN U11080 ( .A(n6695), .B(o[167]), .Z(n7056) );
  NAND U11081 ( .A(n7058), .B(n7059), .Z(c[166]) );
  NANDN U11082 ( .A(n6689), .B(creg[166]), .Z(n7059) );
  NANDN U11083 ( .A(n6695), .B(o[166]), .Z(n7058) );
  NAND U11084 ( .A(n7060), .B(n7061), .Z(c[165]) );
  NANDN U11085 ( .A(n6689), .B(creg[165]), .Z(n7061) );
  NANDN U11086 ( .A(n6695), .B(o[165]), .Z(n7060) );
  NAND U11087 ( .A(n7062), .B(n7063), .Z(c[164]) );
  NANDN U11088 ( .A(n6689), .B(creg[164]), .Z(n7063) );
  NANDN U11089 ( .A(n6695), .B(o[164]), .Z(n7062) );
  NAND U11090 ( .A(n7064), .B(n7065), .Z(c[163]) );
  NANDN U11091 ( .A(n6689), .B(creg[163]), .Z(n7065) );
  NANDN U11092 ( .A(n6695), .B(o[163]), .Z(n7064) );
  NAND U11093 ( .A(n7066), .B(n7067), .Z(c[162]) );
  NANDN U11094 ( .A(n6689), .B(creg[162]), .Z(n7067) );
  NANDN U11095 ( .A(n6695), .B(o[162]), .Z(n7066) );
  NAND U11096 ( .A(n7068), .B(n7069), .Z(c[161]) );
  NANDN U11097 ( .A(n6689), .B(creg[161]), .Z(n7069) );
  NANDN U11098 ( .A(n6695), .B(o[161]), .Z(n7068) );
  NAND U11099 ( .A(n7070), .B(n7071), .Z(c[160]) );
  NANDN U11100 ( .A(n6689), .B(creg[160]), .Z(n7071) );
  NANDN U11101 ( .A(n6695), .B(o[160]), .Z(n7070) );
  NAND U11102 ( .A(n7072), .B(n7073), .Z(c[15]) );
  NANDN U11103 ( .A(n6689), .B(creg[15]), .Z(n7073) );
  NANDN U11104 ( .A(n6695), .B(o[15]), .Z(n7072) );
  NAND U11105 ( .A(n7074), .B(n7075), .Z(c[159]) );
  NANDN U11106 ( .A(n6689), .B(creg[159]), .Z(n7075) );
  NANDN U11107 ( .A(n6695), .B(o[159]), .Z(n7074) );
  NAND U11108 ( .A(n7076), .B(n7077), .Z(c[158]) );
  NANDN U11109 ( .A(n6689), .B(creg[158]), .Z(n7077) );
  NANDN U11110 ( .A(n6695), .B(o[158]), .Z(n7076) );
  NAND U11111 ( .A(n7078), .B(n7079), .Z(c[157]) );
  NANDN U11112 ( .A(n6689), .B(creg[157]), .Z(n7079) );
  NANDN U11113 ( .A(n6695), .B(o[157]), .Z(n7078) );
  NAND U11114 ( .A(n7080), .B(n7081), .Z(c[156]) );
  NANDN U11115 ( .A(n6689), .B(creg[156]), .Z(n7081) );
  NANDN U11116 ( .A(n6695), .B(o[156]), .Z(n7080) );
  NAND U11117 ( .A(n7082), .B(n7083), .Z(c[155]) );
  NANDN U11118 ( .A(n6689), .B(creg[155]), .Z(n7083) );
  NANDN U11119 ( .A(n6695), .B(o[155]), .Z(n7082) );
  NAND U11120 ( .A(n7084), .B(n7085), .Z(c[154]) );
  NANDN U11121 ( .A(n6689), .B(creg[154]), .Z(n7085) );
  NANDN U11122 ( .A(n6695), .B(o[154]), .Z(n7084) );
  NAND U11123 ( .A(n7086), .B(n7087), .Z(c[153]) );
  NANDN U11124 ( .A(n6689), .B(creg[153]), .Z(n7087) );
  NANDN U11125 ( .A(n6695), .B(o[153]), .Z(n7086) );
  NAND U11126 ( .A(n7088), .B(n7089), .Z(c[152]) );
  NANDN U11127 ( .A(n6689), .B(creg[152]), .Z(n7089) );
  NANDN U11128 ( .A(n6695), .B(o[152]), .Z(n7088) );
  NAND U11129 ( .A(n7090), .B(n7091), .Z(c[151]) );
  NANDN U11130 ( .A(n6689), .B(creg[151]), .Z(n7091) );
  NANDN U11131 ( .A(n6695), .B(o[151]), .Z(n7090) );
  NAND U11132 ( .A(n7092), .B(n7093), .Z(c[150]) );
  NANDN U11133 ( .A(n6689), .B(creg[150]), .Z(n7093) );
  NANDN U11134 ( .A(n6695), .B(o[150]), .Z(n7092) );
  NAND U11135 ( .A(n7094), .B(n7095), .Z(c[14]) );
  NANDN U11136 ( .A(n6689), .B(creg[14]), .Z(n7095) );
  NANDN U11137 ( .A(n6695), .B(o[14]), .Z(n7094) );
  NAND U11138 ( .A(n7096), .B(n7097), .Z(c[149]) );
  NANDN U11139 ( .A(n6689), .B(creg[149]), .Z(n7097) );
  NANDN U11140 ( .A(n6695), .B(o[149]), .Z(n7096) );
  NAND U11141 ( .A(n7098), .B(n7099), .Z(c[148]) );
  NANDN U11142 ( .A(n6689), .B(creg[148]), .Z(n7099) );
  NANDN U11143 ( .A(n6695), .B(o[148]), .Z(n7098) );
  NAND U11144 ( .A(n7100), .B(n7101), .Z(c[147]) );
  NANDN U11145 ( .A(n6689), .B(creg[147]), .Z(n7101) );
  NANDN U11146 ( .A(n6695), .B(o[147]), .Z(n7100) );
  NAND U11147 ( .A(n7102), .B(n7103), .Z(c[146]) );
  NANDN U11148 ( .A(n6689), .B(creg[146]), .Z(n7103) );
  NANDN U11149 ( .A(n6695), .B(o[146]), .Z(n7102) );
  NAND U11150 ( .A(n7104), .B(n7105), .Z(c[145]) );
  NANDN U11151 ( .A(n6689), .B(creg[145]), .Z(n7105) );
  NANDN U11152 ( .A(n6695), .B(o[145]), .Z(n7104) );
  NAND U11153 ( .A(n7106), .B(n7107), .Z(c[144]) );
  NANDN U11154 ( .A(n6689), .B(creg[144]), .Z(n7107) );
  NANDN U11155 ( .A(n6695), .B(o[144]), .Z(n7106) );
  NAND U11156 ( .A(n7108), .B(n7109), .Z(c[143]) );
  NANDN U11157 ( .A(n6689), .B(creg[143]), .Z(n7109) );
  NANDN U11158 ( .A(n6695), .B(o[143]), .Z(n7108) );
  NAND U11159 ( .A(n7110), .B(n7111), .Z(c[142]) );
  NANDN U11160 ( .A(n6689), .B(creg[142]), .Z(n7111) );
  NANDN U11161 ( .A(n6695), .B(o[142]), .Z(n7110) );
  NAND U11162 ( .A(n7112), .B(n7113), .Z(c[141]) );
  NANDN U11163 ( .A(n6689), .B(creg[141]), .Z(n7113) );
  NANDN U11164 ( .A(n6695), .B(o[141]), .Z(n7112) );
  NAND U11165 ( .A(n7114), .B(n7115), .Z(c[140]) );
  NANDN U11166 ( .A(n6689), .B(creg[140]), .Z(n7115) );
  NANDN U11167 ( .A(n6695), .B(o[140]), .Z(n7114) );
  NAND U11168 ( .A(n7116), .B(n7117), .Z(c[13]) );
  NANDN U11169 ( .A(n6689), .B(creg[13]), .Z(n7117) );
  NANDN U11170 ( .A(n6695), .B(o[13]), .Z(n7116) );
  NAND U11171 ( .A(n7118), .B(n7119), .Z(c[139]) );
  NANDN U11172 ( .A(n6689), .B(creg[139]), .Z(n7119) );
  NANDN U11173 ( .A(n6695), .B(o[139]), .Z(n7118) );
  NAND U11174 ( .A(n7120), .B(n7121), .Z(c[138]) );
  NANDN U11175 ( .A(n6689), .B(creg[138]), .Z(n7121) );
  NANDN U11176 ( .A(n6695), .B(o[138]), .Z(n7120) );
  NAND U11177 ( .A(n7122), .B(n7123), .Z(c[137]) );
  NANDN U11178 ( .A(n6689), .B(creg[137]), .Z(n7123) );
  NANDN U11179 ( .A(n6695), .B(o[137]), .Z(n7122) );
  NAND U11180 ( .A(n7124), .B(n7125), .Z(c[136]) );
  NANDN U11181 ( .A(n6689), .B(creg[136]), .Z(n7125) );
  NANDN U11182 ( .A(n6695), .B(o[136]), .Z(n7124) );
  NAND U11183 ( .A(n7126), .B(n7127), .Z(c[135]) );
  NANDN U11184 ( .A(n6689), .B(creg[135]), .Z(n7127) );
  NANDN U11185 ( .A(n6695), .B(o[135]), .Z(n7126) );
  NAND U11186 ( .A(n7128), .B(n7129), .Z(c[134]) );
  NANDN U11187 ( .A(n6689), .B(creg[134]), .Z(n7129) );
  NANDN U11188 ( .A(n6695), .B(o[134]), .Z(n7128) );
  NAND U11189 ( .A(n7130), .B(n7131), .Z(c[133]) );
  NANDN U11190 ( .A(n6689), .B(creg[133]), .Z(n7131) );
  NANDN U11191 ( .A(n6695), .B(o[133]), .Z(n7130) );
  NAND U11192 ( .A(n7132), .B(n7133), .Z(c[132]) );
  NANDN U11193 ( .A(n6689), .B(creg[132]), .Z(n7133) );
  NANDN U11194 ( .A(n6695), .B(o[132]), .Z(n7132) );
  NAND U11195 ( .A(n7134), .B(n7135), .Z(c[131]) );
  NANDN U11196 ( .A(n6689), .B(creg[131]), .Z(n7135) );
  NANDN U11197 ( .A(n6695), .B(o[131]), .Z(n7134) );
  NAND U11198 ( .A(n7136), .B(n7137), .Z(c[130]) );
  NANDN U11199 ( .A(n6689), .B(creg[130]), .Z(n7137) );
  NANDN U11200 ( .A(n6695), .B(o[130]), .Z(n7136) );
  NAND U11201 ( .A(n7138), .B(n7139), .Z(c[12]) );
  NANDN U11202 ( .A(n6689), .B(creg[12]), .Z(n7139) );
  NANDN U11203 ( .A(n6695), .B(o[12]), .Z(n7138) );
  NAND U11204 ( .A(n7140), .B(n7141), .Z(c[129]) );
  NANDN U11205 ( .A(n6689), .B(creg[129]), .Z(n7141) );
  NANDN U11206 ( .A(n6695), .B(o[129]), .Z(n7140) );
  NAND U11207 ( .A(n7142), .B(n7143), .Z(c[128]) );
  NANDN U11208 ( .A(n6689), .B(creg[128]), .Z(n7143) );
  NANDN U11209 ( .A(n6695), .B(o[128]), .Z(n7142) );
  NAND U11210 ( .A(n7144), .B(n7145), .Z(c[127]) );
  NANDN U11211 ( .A(n6689), .B(creg[127]), .Z(n7145) );
  NANDN U11212 ( .A(n6695), .B(o[127]), .Z(n7144) );
  NAND U11213 ( .A(n7146), .B(n7147), .Z(c[126]) );
  NANDN U11214 ( .A(n6689), .B(creg[126]), .Z(n7147) );
  NANDN U11215 ( .A(n6695), .B(o[126]), .Z(n7146) );
  NAND U11216 ( .A(n7148), .B(n7149), .Z(c[125]) );
  NANDN U11217 ( .A(n6689), .B(creg[125]), .Z(n7149) );
  NANDN U11218 ( .A(n6695), .B(o[125]), .Z(n7148) );
  NAND U11219 ( .A(n7150), .B(n7151), .Z(c[124]) );
  NANDN U11220 ( .A(n6689), .B(creg[124]), .Z(n7151) );
  NANDN U11221 ( .A(n6695), .B(o[124]), .Z(n7150) );
  NAND U11222 ( .A(n7152), .B(n7153), .Z(c[123]) );
  NANDN U11223 ( .A(n6689), .B(creg[123]), .Z(n7153) );
  NANDN U11224 ( .A(n6695), .B(o[123]), .Z(n7152) );
  NAND U11225 ( .A(n7154), .B(n7155), .Z(c[122]) );
  NANDN U11226 ( .A(n6689), .B(creg[122]), .Z(n7155) );
  NANDN U11227 ( .A(n6695), .B(o[122]), .Z(n7154) );
  NAND U11228 ( .A(n7156), .B(n7157), .Z(c[121]) );
  NANDN U11229 ( .A(n6689), .B(creg[121]), .Z(n7157) );
  NANDN U11230 ( .A(n6695), .B(o[121]), .Z(n7156) );
  NAND U11231 ( .A(n7158), .B(n7159), .Z(c[120]) );
  NANDN U11232 ( .A(n6689), .B(creg[120]), .Z(n7159) );
  NANDN U11233 ( .A(n6695), .B(o[120]), .Z(n7158) );
  NAND U11234 ( .A(n7160), .B(n7161), .Z(c[11]) );
  NANDN U11235 ( .A(n6689), .B(creg[11]), .Z(n7161) );
  NANDN U11236 ( .A(n6695), .B(o[11]), .Z(n7160) );
  NAND U11237 ( .A(n7162), .B(n7163), .Z(c[119]) );
  NANDN U11238 ( .A(n6689), .B(creg[119]), .Z(n7163) );
  NANDN U11239 ( .A(n6695), .B(o[119]), .Z(n7162) );
  NAND U11240 ( .A(n7164), .B(n7165), .Z(c[118]) );
  NANDN U11241 ( .A(n6689), .B(creg[118]), .Z(n7165) );
  NANDN U11242 ( .A(n6695), .B(o[118]), .Z(n7164) );
  NAND U11243 ( .A(n7166), .B(n7167), .Z(c[117]) );
  NANDN U11244 ( .A(n6689), .B(creg[117]), .Z(n7167) );
  NANDN U11245 ( .A(n6695), .B(o[117]), .Z(n7166) );
  NAND U11246 ( .A(n7168), .B(n7169), .Z(c[116]) );
  NANDN U11247 ( .A(n6689), .B(creg[116]), .Z(n7169) );
  NANDN U11248 ( .A(n6695), .B(o[116]), .Z(n7168) );
  NAND U11249 ( .A(n7170), .B(n7171), .Z(c[115]) );
  NANDN U11250 ( .A(n6689), .B(creg[115]), .Z(n7171) );
  NANDN U11251 ( .A(n6695), .B(o[115]), .Z(n7170) );
  NAND U11252 ( .A(n7172), .B(n7173), .Z(c[114]) );
  NANDN U11253 ( .A(n6689), .B(creg[114]), .Z(n7173) );
  NANDN U11254 ( .A(n6695), .B(o[114]), .Z(n7172) );
  NAND U11255 ( .A(n7174), .B(n7175), .Z(c[113]) );
  NANDN U11256 ( .A(n6689), .B(creg[113]), .Z(n7175) );
  NANDN U11257 ( .A(n6695), .B(o[113]), .Z(n7174) );
  NAND U11258 ( .A(n7176), .B(n7177), .Z(c[112]) );
  NANDN U11259 ( .A(n6689), .B(creg[112]), .Z(n7177) );
  NANDN U11260 ( .A(n6695), .B(o[112]), .Z(n7176) );
  NAND U11261 ( .A(n7178), .B(n7179), .Z(c[111]) );
  NANDN U11262 ( .A(n6689), .B(creg[111]), .Z(n7179) );
  NANDN U11263 ( .A(n6695), .B(o[111]), .Z(n7178) );
  NAND U11264 ( .A(n7180), .B(n7181), .Z(c[110]) );
  NANDN U11265 ( .A(n6689), .B(creg[110]), .Z(n7181) );
  NANDN U11266 ( .A(n6695), .B(o[110]), .Z(n7180) );
  NAND U11267 ( .A(n7182), .B(n7183), .Z(c[10]) );
  NANDN U11268 ( .A(n6689), .B(creg[10]), .Z(n7183) );
  NANDN U11269 ( .A(n6695), .B(o[10]), .Z(n7182) );
  NAND U11270 ( .A(n7184), .B(n7185), .Z(c[109]) );
  NANDN U11271 ( .A(n6689), .B(creg[109]), .Z(n7185) );
  NANDN U11272 ( .A(n6695), .B(o[109]), .Z(n7184) );
  NAND U11273 ( .A(n7186), .B(n7187), .Z(c[108]) );
  NANDN U11274 ( .A(n6689), .B(creg[108]), .Z(n7187) );
  NANDN U11275 ( .A(n6695), .B(o[108]), .Z(n7186) );
  NAND U11276 ( .A(n7188), .B(n7189), .Z(c[107]) );
  NANDN U11277 ( .A(n6689), .B(creg[107]), .Z(n7189) );
  NANDN U11278 ( .A(n6695), .B(o[107]), .Z(n7188) );
  NAND U11279 ( .A(n7190), .B(n7191), .Z(c[106]) );
  NANDN U11280 ( .A(n6689), .B(creg[106]), .Z(n7191) );
  NANDN U11281 ( .A(n6695), .B(o[106]), .Z(n7190) );
  NAND U11282 ( .A(n7192), .B(n7193), .Z(c[105]) );
  NANDN U11283 ( .A(n6689), .B(creg[105]), .Z(n7193) );
  NANDN U11284 ( .A(n6695), .B(o[105]), .Z(n7192) );
  NAND U11285 ( .A(n7194), .B(n7195), .Z(c[104]) );
  NANDN U11286 ( .A(n6689), .B(creg[104]), .Z(n7195) );
  NANDN U11287 ( .A(n6695), .B(o[104]), .Z(n7194) );
  NAND U11288 ( .A(n7196), .B(n7197), .Z(c[103]) );
  NANDN U11289 ( .A(n6689), .B(creg[103]), .Z(n7197) );
  NANDN U11290 ( .A(n6695), .B(o[103]), .Z(n7196) );
  NAND U11291 ( .A(n7198), .B(n7199), .Z(c[102]) );
  NANDN U11292 ( .A(n6689), .B(creg[102]), .Z(n7199) );
  NANDN U11293 ( .A(n6695), .B(o[102]), .Z(n7198) );
  NAND U11294 ( .A(n7200), .B(n7201), .Z(c[101]) );
  NANDN U11295 ( .A(n6689), .B(creg[101]), .Z(n7201) );
  NANDN U11296 ( .A(n6695), .B(o[101]), .Z(n7200) );
  NAND U11297 ( .A(n7202), .B(n7203), .Z(c[100]) );
  NANDN U11298 ( .A(n6689), .B(creg[100]), .Z(n7203) );
  NANDN U11299 ( .A(n6695), .B(o[100]), .Z(n7202) );
  NAND U11300 ( .A(n7204), .B(n7205), .Z(c[0]) );
  NANDN U11301 ( .A(n6689), .B(creg[0]), .Z(n7205) );
  IV U11302 ( .A(n6695), .Z(n6689) );
  NANDN U11303 ( .A(n6695), .B(o[0]), .Z(n7204) );
  NANDN U11304 ( .A(n6692), .B(n7206), .Z(n6695) );
  OR U11305 ( .A(e[255]), .B(init), .Z(n7206) );
  ANDN U11306 ( .B(init), .A(ereg[255]), .Z(n6692) );
endmodule

